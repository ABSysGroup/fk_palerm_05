`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PZ9WssJVas3MlCAJeWCr1KO/cAjuWUjxL6KECRzCsWBSJRQqJH8ZqsZaCzmE5Hv6
ZjOcF3sRiz5QMAZRb6/vf73Ek1lGMNSyjLMDxeWy3s0ZGLS3V/Pdw8/78bea3iR0
yyLb6QggaxMrJeGiu4AUsMvx06PdydYHVRc2Bi4aCvUV6klsLiX8+2ujn1WoFtm3
Mo3/2+rCwdK1KG8cn8w/Y+nKCLX5JAPYiTRTYS2rIzjptODMvVd809P097dRP52w
ka1LKxknXXxdRwhusdDkwygzzqMOWWWzZXP8oGxLvTMeWr+fB0GAmwT3qD3DEuxI
da4Z8wBOsdmXP50s1VTHF1/zlMpVDM2tcZFkz2x6m21Y0MzrrTY/X0iOPrq1do6V
zQTMm9up7PA1IfY2geMkRoXSzPP+smzXzCd0x/jrNAoWbPCLJ/MaIs7lI/GXlq26
P51+m8a9aI3XP73QMGoM5r88XQFTfuVXGeGFPtCKPFo0eZ9r6wurwWJX6qeDKy1a
5k4LGrV2ZEm8CqD/U4BvAsP3k/Nlv8Ls+hSiFuOhDz9sRqgQVIVerPLIWZX/8N6u
t7awPXRYrLz388eYG9Tyi7KCqLZ3EMPwgyh4o/dOiet3C0nF8TPGP0FLY1kZkxK7
K1Vc/tH6RYa8Y6QN+0Fq0sa1yUl22dHakVFOz0gr6xLW4CUs9WVpEfBAy4f7/sob
6+ij9xPqjl1bno95tr0OvhnqC3Wj1X5PAJOa4WbblI2XlL5nMxu04DieB+e7ablz
ZT4yUH9xgT64gnJv86BP8dNyQkyFfz4aRy7tw+m95QL71tRZ4xs1PxOGmF2nRGKX
dZEH7hwREV90w3AHYLvgAbX+xumgkJY4oec+3f+4Lvda2clU0JwvWCI8yQnDX6YF
/sm+KbBj+4e0/hQYCk0IHqcu16IRrFRkejYLxD9MLug8YhbzjeJisRuwy35nXfa0
mGqQlsdK3XvoPJ0D0QhxVvyZl9FACMOn+WfrIqH5ciFdc9G92glDQWrd72tvlkIP
6M4cFpARBsiTNOpmWpzAwIk8tRFUqsowGX8cCZ7vRECrR8a0odj3ETGM0SzA63CU
wa4OsLkR0lUStzWttXT4LouqkROfvu6BSxLHF50Dv0DCIbY7NTKMe1UuFmWPufDB
CV5rHeirPTuaJ83vgW2grEBxCI8fqOQsul2I1ZI5Da1KUOQo++5VfT/TwO7WnFi+
GDIK+p4zeL0Rh+fdCbTSxrpBNT7ihF3VyM49xrXIueJ4vNpC4bRIQSM3aNqiU47z
nkaxUuskDNZ4iLBnyzEb+9ORDVni5sKknMvi22fklsXdj68+ywY9zNEP+QGtrWph
hQPbyxONxqMkJpWO7knyH5ZPJ6xhx4RglmFTjh6yuUyfEBaV+/FSpJAufTjazYFY
i0L33t59x2kBJwrfvjjypUvQtUAH2Rn07nmVy8SXJbu9+05JgglJMeH0K/rbsSmX
hgGs4LBbrbQVBlYnrPRcb3TDCJ2SeK4YAGXCSDIT/6nynTrIio+9KzZHQbFgNYex
qzATHVHyzsIb2795I7C9XDG+d6+L/cpClODSwkNbefw+BGzpk1Zm4h4g4d7ffxlB
f2QtZ/QwAOzT9HnCFcnB4qug1NSItJO5c7/YDlREBvx3s7o56AWqi966740Trsuo
G38FX845z2oR1+3d1cpjoqwsgm0Xv/5vc7PSfSnmdI5prOutMEXLlhgv2Lw8r7WH
MC5d67SWj5nIY8uYn706/nMG/x7MxaINLr9Y63xuU/U1w1seuqgupBctfNsvINzW
TNnkD2i7lZKmxzDrV4Zx0LrwBS4i9yNtSy0IgqNNAzabILaMIrVBlbliZvXgeObw
aSbwoovf6DmE6yrczCUWGVFEtmfR3l9JIp7LoOt4wQtMWTqM4n7I8R+5tEKq4TWS
zjT9DLfJ4mrXtDn+/8tt4xsGJTj2qnXuP0UhJFLaQdaguQGFrjXQugpNnZHTjQSv
Ry0Ewa1/utaq2wvX0mQfQytvAc3S0XIZRy6peJSWApQ=
`protect END_PROTECTED
