`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yRDLzx1gr+oUiWHBYWeOXpcELE7ThDfsjaC5JbpVktglBZorCmOMuy4qKJt0LoJr
W7rci+ytZm15sEwZIx0+OipweDTgIskG00bxx6psZECtSoegkFtwINH05tjXRR8I
fjnYo10NPDLvx2QfTdfXZhzkXj3iD+ZBt+nRGIXOiXo6rwUeG6dBywVeaCQ/VDF4
RcqOerQHflRGtYilh0u8RztkZmP36WWUPc+yZAj9DOl/ydUomd6TbhUtIcTvFISH
r+8WihP91skfEfSLBcyYn3RNXtgDl0PAak+OIcJ7BBBncvLC2+7DQwRrthLkWYO/
tcA57xL8R6MBJL3QurCK2IzCfBQKNNe3op9w+kEeqOJh02R3vCYgOYurFVeGaM34
DtW4LRJMSf9ginaheVAyuw4jjEcxDs/pUfCvHGxI6envI+BMoZywzOMAYhCxtmkI
U89s9lJuBE+2S78hlXAnjvifzZ8kP2SW+mZt96AJdWUfzl7RKzmm7qi+HLSUKA3l
b175sazHPB2NLTUxXDzwckWwqd9+9jVdXW6slqSbGDOWjfa+1dMQmzkjVZ67LOZ0
dsGtKvkc4J/sStlI7Fhym05UJU1s3H1nWh6EgFRZP0Zquuq5FfPn1OgiAkaB1c6R
jtM2+CFGHxuRD4zZTpa4Gw==
`protect END_PROTECTED
