`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nowmz4sTWkBDDDya8VB4Mao4H66GyN9KN92d3WeLnkTx7iVkW/JQ3CfRaw6yAOQN
J4nAZ5W2qLGK5j0a0VYj5fUfoY0KTi3o/T1PTapKh2/hDEBlqRw3/JxibCqVwooF
thHyph2CsT5P/3ZNSN71dDsb2axMeXKIWOKFz9vkow5stc+kaDrTYPzkY0Y8flfH
ye80e1nkdb2I9/KiJ4Byq5dqkW7dV+Tw8bDL++rkUACD9J/B2I29CkA6tL3Gkxbq
tH90M2RQhJbrUpd1LQJXqqqEZeNJcNfjekP6wD5XTfT68JXD+z+kGcw+6ge17iOm
th87XEmTVfgDuhSaSA7NZxjWO7BxmS93lDDPo9PFKCRUTpVj8T87JvQiGnk28JvS
tJtddxTmzUjvQr/Ywqm3FcbSoz9gJkc4+nJ0fRpq88as+jU6EXSfze/BWAoDXE1I
/FpzdbR9s0Utz2YWxUBh7kK5ybuqdt0SwYAj1+3cJMCOwhuJTeepFxb1RgnpxDZ0
JW/un+X9D721BpXD2UqfB//oLNJwCcy1xd27Hrz0rWo3wQWgaYMDLbqW8kfm07HU
MpZLflbSYWIRsFk5j3nzWhDQGF9FwoMAFKhT86YX0IEqzgnwqapiwhjCqZW5PH31
ZKzRBPdc9necJYuPwxnU5WgLWP8rQufkDiPtOp5OXMqmcm6NmH8dx98UVQRqrc0+
4Oq0pHCVtBQJI2vt67yVwaDiLXalFQWkr1VjmQVweXklOzIlw8+mN/YC8gN5JXOt
SrBcVnGTMNqKvck4jGCGgF/PVnVrZbKAwOZCw6+Tc5UJCKZlkOGkG1RVFRsCa36+
Lbx1/bX7/ZIS2bJ0I7G72TgWhNxWqCzTTwyyG2u1gcXHlat4shQvm8layTs6/t2M
kceSMYpG2PiJf2Guzkwvslr6zHpKL0aF9QnqwaLB3KUhbjGRXx1AdFwZphLQT5cc
D+IbZLgurxx9NPi9Qj70yeDziMncVlGqao50hI0EG7zO+n2zaxzxssSyEWPyVwF1
2UgiWTLLbl5XrvYzZr/68r4b5MBuXkES8zDlX4LDEMlKQfe4y90CBSA6jkb3BDk0
Bh6NLWnhJYcBNqVgFEMXTLQfhPyivP5HOjhXPH/CuBGxrabr99I7zOuXemEtB2ph
ugP7xPuJimQ0DCvia6kVwf3aoeOsIbb/6fpTHBjmdMWEwnCJj4vh+oL2KfkTTtSB
6TAEArDiqpbjgAZAwmjzt/xcZLsAp0VJqBcax5Iuv+aLbRxanHfOvmIsC9Ypzgcj
qAbsahZA/l1/eNVA80Obx4cYPu6XkMvTuLmymvb8RpXQae2rapQ1vt7q9q239UUC
cAialJ2Mk9Qg0jETKzh5P1Y95gEidJpsf4aWY//pj3ln2w9XC5sYm6SegMZ8/i83
uUZZxDEKsaO4ztljgJ7JdO8DBekd+zF1s9d7t5SORXqlgalbY8X1nBxPAVtPoXYf
f5KEkKrgUoAYEj4lxrIWCTfaYIeBSQ4q5mdlRBZcOztFUFqO+GxM7jMl/qeWRCaL
jLEK9SY/zuuOkqQS+KN4Tb/1HZVNO8sptxHlMjUVkRHAXlASTrQRxufHyYoTPpyc
viNjsXihgbjWzEMGPizRsRZM3tAe6D94all8GVwlOw9q/Ccrshl2WWOTWEpp9vnb
9c+q+NIaDanwviDsqLdz2IULPeBPMmWJPCQngX2O+DtXdLpmFoojMxgmZcpc8gZo
aFZ4+nnoOGV117Iz7p73ptuw+lIsbV8xQmqL35p0i0lc/geslSi59ya7lAik+emK
BESxMhadDTYWJJhYnbPSp0wtdF8gKrWC1IW8figl+9KqZ+oS7UfPxiKPk0uheMCK
4lez3ECfAC6EITA7lkM/FHKhL5hzagpEG9UJNOIFa6dOx/MJZnT0AXN8/b810SG3
e2589YYrvkkfaPAJr7qOCycIr0Z79br/HRZ/QHgpzYldF0whL2vfmOPngdxV28Ls
YiPnJfB1oaYr04qibFQKbYGl2RRuCMwqvwl/AHwrDC/+cy92TLHCWxJzaHzIg8Ar
e4kocbtNZ8f4+d0jBYRvkiKtR5EP1XUr332ZAz21pfaNNCOCBFW3l9DbdHCPzZVj
/QYb/82GKbe5FSKpimZraKc4dLx2XMmvVW+IlUvuSzFoP/tiQe+ofkb3T2u5fhmH
owkzhkMe9kSQ6UiIud8v1aCEvIZAuCXANCidMnl8xCl319+nQyxJRpB8CqR02PNj
ZtcJeAUmtnZMmJD3GMni71ukIVtqWpbfJQaNO5+nIbnG7oTMERuXMHNsmdZv7MQH
sJVKEaBSJf4ixwZO1jdRQoNNvRQ1SIqzXjaa+wqkCwZcsUc2HOoa4S2RDY52QniD
CsN6wc1J23EUB1dgo292VVFw3nkeVQ8ShWLIyNCvtFMpmBXtYi3DUiCIgTFeNeex
Y1c9ADHEFQUE+i6VFZ1zNIbpGcJmVlQJdJ288dVdvAAZpeDipGYopyfzNRSfHlZ8
PFQDim0rccDVwU2am5F3sbX54m5VWH3TNC1O/thie8Mz5G8XIbx5rH/tlhky1t4V
Tdiu1J5SqzT2S8AahJw3EOFwSUnctbrD14g6XH7dsLDDY28yYMFT4BPIh97NcxJr
RClfyzfsMO2YntKBpcln1XdsTZ7E7P0dO1h2RQUVYAqKTZRbpaGssTdCpfqmTIed
Zr1vLUC+ZUx4a/v/N93jdmcq0PQxY9LkyEoufqze/f+Pw47L7utJRXqFV7u7PLen
vl1DtUiXRYSpAfwgXmC+V8p9JedRQdLBxw8hwR+7bpTkm1me+SOe89ZaYZtZNW/I
3DKJf4UROhk9sRvW+J+7d4J0ZoojKnQGEgvlFtH89zC9Ufsd1U5zp+pofZo/Ms1n
g1h/nzGLARIGRzLkXlckKLqoGGhoSQ4SgDYQuFO9wYIrjRU6gzW6NDtUnAqESczG
puJ3Wxea81tme7NP9ZXkTdDpzORuf1hvfCzD2CKxcuCMHVVJsxv6QT8tfqi3fLwp
ut1QSI5DHSV571GlFdkno9UTwXHswcHO/c4sdErCcxrGtR0DFZD6ffizUt84YzKa
a1UWO+9CzU1TPTLqkAMbI/5NZqMOt+RatG+xZ6kaiMa62cf5+W0t7kLipRFUGTvY
Cn1xjYf1rgM+BsaGgtj3Bu9BkcQpdixLsMQO/h1sI88NSiFNh7Xme/sMcfmZtjyv
13DqAA9hZwI6db947vhGDs2xApnxGhHHBQrM0mtWAZw/pLvdooQnI3KfBWEsOO+z
Jq4hzDAOX9XEQSRIq4VNJXaYQDKCHpjx01L2p5tokF0oatJAX6XKcdrNVORlXi96
icyVS4WEbabIFIvo01nIxF6LooL+ItqQDINIifPqZNAcWLQj5shzc1jlclnGkuvI
u5oklaNISGEgTO1VcOifn2L0dZUBLCiMDyB2+8SwDrOxP4fCSFusEWQQ7EYVYIeC
OuNDD4jwUS6Eke93EPMku/hEBAw4y5RkcFrqwuDdGbcWw9XXTiZAW8QIwMkjxLtL
KyVfnfcuonCUQyt6HuJoKy0+AcTtrmtYtcepWkm8DLBP7UCrvw6sNwTd0JnH+Tv8
P8gAs57DBdxY7J+fItnbJ/Ryc/QR4nxg93MXiepsfRHdI64FSl37xPbzUqv8exN5
zwlIl2hZ+S7imaMkVE+6iOiZ2I0qxxPvPhDR3ucBMPoJTDXOyCT1KATgBomXQ++a
kwk0TLfjjcYTfoxyh41iEopet8eblrLfIZXhxG0ZrKYT94CLwAy57H99kyAqFEID
SdbpuV44WATQjemR01xPxwQ7FtBVSovDWIm9ik7H1trP14haSqidcbdsLvl2rKjW
Ke0LjY3+ba/SgoBrHCliA1UDzTep+c58kiE7/pKdflaLY4q556xSYJ6R88Em/wkN
fcASFbFRuzR9DGvt35/QUcT3itqy1N2EBK3cOsQJUXyAfF80sVTEoNtj9DtKoGdb
R4PO/2/PQboirxSZDj/FrYZfapLOzoqSTRxSZa5PczvPQymGlbqzGNGDXlRhFb54
NsOMgRbJG2jMuvGCuPlwUV0M+E/h4vRArUT40BvE+OKAYJWtjTupxoibRnFJHXW8
Wtm07NN5K4JO5vI/Hi6835wKRB8Ynh4O53JmGcG9rbOT/DZiiZvrM7y0hzvy5bcZ
Yj65T8B+YajG0G/ojqeOuriLFfCfCpa+/ijajAIDNA5NNRJ1Ur1hUhx1/BBTDvNX
9l9JGy0cnW/MXy2T/tRiRyuzQ3KWdPXLjCmYPx9EkOQ=
`protect END_PROTECTED
