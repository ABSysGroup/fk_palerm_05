`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U0dWDPicjm+WAB4XL8NHFGM+bHS9eXlAWXb3MZyLjMa+1fUg1k/FZCvN5VvDwHQX
8brBVuISohc5MDblMP59nXXcoipqD7aMoyvnTK/LcSwnjANyND8IPEW6DxFFrN13
DMbNZez5FQbNJR+Sgl7v7Y2qeAgrop41Azf1IG7uwFtYv67/E0pKCw6duJpOlX6+
dXfKk0Ef4iQT8aNc+49b5v1miXL7AkupQ6nFs8N6bXdZClyO5n0ptxARf5DtoRT/
UP4IXjlZlmAzC1bsjxprWVYjtKuJUhWyN2UjAowOH6mHPB76lX4NNwZPIB6pzczE
vBSDD2CyaVZ4eMWcOPnYKA==
`protect END_PROTECTED
