`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gv3/pSIyw/rL/LwKBY/qLOBGVX9pidg6na1oZWM9p+hNwzq3c9+QaOjYJGq8j6pi
A5tEvdOFqJ0MCqOfkrkjPK+LGn3dNaGrV8UfRQAxgAJL2ZSKMUz9Hov7VQmSTAep
Q48ofLYufRxnkL4ysK/HzxFYeyNhBSV98bYd4C0bhbf1z6keioUuLIjlcxt0nH1r
Gammhv9iiltn2cK6dvQyzGzaxKqda3j7qt3zgM0AE0YoEQC0bLyAM+cu+kf8eToh
4rCidOrouWZrKY2n+IvG/BwnGPEWqjQsV5ESWs416lXGDGBGT2PpgIkcfBmRRaXF
/CmMeUzdDx/iiTJVZOmwlqJjfaRHiXTbjXJ8lBkGzPl2qzQHJeF17CH0CA03KpCs
bJ/RN5+qFpi9LWS0O2loUA==
`protect END_PROTECTED
