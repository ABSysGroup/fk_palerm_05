`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xp7KzNMGDpZ4hQCwn4Vk8mA8EJ9dnTsL1gZlPY67HlyRc/lDOIKfGltD4mxyyOij
+oOyd9LvdAx8Bmp772h6s8CTyjEzD1QD6nAxyBNk5KoqFvE5R7c83y+8a7LFINrZ
cckFuzMgWkgNpgADXSxE7Sbsb6NcULK0U7ApEzjP8/ZfrVP1qxmPsWgjHKHpZbXp
Gbt9GEHRbmUn2Tj61wJruUhMhC8xtMvbtf0pzX3+gh7Zp4iSPXj3rY+S3jbUSGm7
WS5Tu+5cqsJKz9p+Phm/R4IUltT7Lt9kH2cZbFAZkovWv9nIZUhJULS3TZ46QK4o
vZ39nEfdT5k5c19Dew4qGg==
`protect END_PROTECTED
