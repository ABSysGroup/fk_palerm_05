`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7htaU6gaK4cy6Rx47Ha3ToG1xbPimfkAt+H4bJt444Zhboy135Ii3JYaFkgOlI5L
GtgrqEXbibm6RaEliSnpVg0GdOV8se+FfalnKECCtPHFEGBfRVtKqD4D57Us+9hH
n1oHNGVkvFP1h3Yi75QNq478Roe0rp9QLDQHhnaeyP2Mb18aC+2vI16IS20ggG1h
0fsOqyThH2Pzgt2fPLxfptwvDKYa/Tz19Z7Cme//u4FBmzuVQ7t/+LNbA8Pe+8t3
u61D1S3YFYWIFfyXSC6Wo1CR9isq0WjFe2zt9GIwgeOXkIhfmvlDUju3GLX31rH9
2ffWVDl2r6r9SuQHS/4kAgXudxMyc0PYspReZ7s7hiOi0bPoyfv/aQ58pm16NCok
+G/vmUJY9TME2OWJcNp6ptgeR9VJzSSEsbr3zRWgbuE8YothHKPYPVJ69PrD15Ur
/q7lUzCi7/uYmuk+digobn9oeVmoPoruTuvYLgrurlVcQppuBJ1+KzLH4tDsmFFZ
ue8kmCGr2m0ZgmKx6j/UxgPeIHcQO5EVequzABtKQZLugpkD7hJbrM7uv2Hv4fDs
Q278tiF95NOTkdeN0KGDz64qIixQwEuQiua1C/dbjneM5WOCOv70wj9tTj9oe4qb
6Xsfz4+M6HgNqfBsMu08LG5ZGYfXzubbwa8k9SGrx/j1g1YqNARW0I6MEJWd5YhD
LXHRnhj5ovCWwVjwwM/UP9znUX2I4FEj4G9Hzg95AM00XTwTPHHS6U4sHchb2oiD
csKwqIzj7pJcsCEh41WoZg==
`protect END_PROTECTED
