`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Gt0OMc7ZRHA3+jz+4shMa9rQv7yYlsKZYbPF6vLWjQikgXUIrd62me6KFO2UCHC
kHoIkAiCLsx/gnUxlUqXhOloczZf73MLkdvFvlz/8o2sicPMrlfH+1seIzejPN4R
dE0yQpEhrjToHoOOj4QvXepa7TAUe/LHfhExIGua490qIQCXrWQSnONl31jDjgWH
hMMQIbJJk4Z0Y2DLrlS7psZHjOqRo/R6gWwCgbUTgR7jtVt8+HYTcLTxQ23Wcdfz
Kz8JP+md4T/AOI2LayxJjcUI7Gl0FPBjPs9eyVQ2Cjrr02rZgN0XWbpkIqaPTA4E
PVU7c0F5tnwxNc0S/DMxi+oxI9BR2N02+EtiCmrfYVvM+jPgDJWX5fe8Njk1jXaq
b17yDfOJi90+bxZH54Wweg78IP3ftjqIqpGrpJ45WrVX0df0eetwMAS5T0uE7IaB
SxLAOL2EysV0+Jo2m0IcDObgY72tebycSiCbX3bgmXL0Y6lm+O/C1HvWqZMR9k8h
skfJlf423noTBQuGrMhFydgnvlf81UNEW2UZ7R5852PLCyPUWxUDOP9BRyrUViXE
POBy3F7nDwhf3HeVUPLwnoUSDlXz0urzMXsVk8zuyqO67jsZfqe3ObAWlMwHchhh
QUEn1qS7vQgQ9R575M5GEZhOcYZ5RRXYZWi5gtErQlFt61HzgFsxnTzPlyDRYcTl
Nm848/Re+VPMoSQh9DXy8lNlKcIBNrRyrFszeLWwxYSGNYun4OkjCvl1X2Qdr1Sa
cWFHWJXBQig5Gx7DjjuHyBE507S71HawdbtEIts+e9kFY5mkcR8VsGZhIOrmLN4z
XoT5QNtp1va53R4j8iUrHjjCQzbgUI70eVvkg/V/hywoV2yd3ULiM+DBiKY3D6G5
g/AbAAVbTAmcK1BYKLZ+02+AfOy3srPHOLQ8wZtt6VztnKblQl1zk4JWup9zJkD6
cGvOwlFpFodFap/lPnOUC+JlG4N1fN5zCXb2HDngm7gWMd4KBhNcar6Xw5HAyFeI
wj6w6BUXfbuJbe2aPRTYG2H+Rn4LcsiBuuNjz8ptUE0ThxyWoQg1rxYWOyx8Q3E2
N7KcFjrk5XLLgdtM3yx+bl19vFq6zpdeKhaDcYSR1HpeSbuucY9XfHtMyG+vHjWw
eoOwBHwuECYhA9sC6wDRsUlGA30mC6zOCIqrfazYiYLaJ29gTWCu6ymHgdAc5zf3
sxE0XeyRl7S5swEaBKqDuEsJz1O+MwCeT9QOwZtBNhXLyNaBiQfvB2nU1Is6TgN+
YDZC41+J7fC1jCzqdyZUW629MO5sLQkNftYd0I7k9MKrhJGNEYy9nyegSGx/4wNV
o/StH1IyIqqRNE9Pg0ncVOmiSx3ZSH5DCfwkhdLreDrKoYB3j6QFv2SeVven4UMg
h/rEVjfOugZ1f5keEf1O46EtuEYxbRcGogc4vLKNCsvX1fX7QHIi8bKlAIJalQxx
6wCDDMGXBqBu2iKMaJy1e5Ejblm1oIDcIKXbzqnut7gDo+YiVzRfYc7Z20lU/5E1
vJ0u3Ll4owcmwawoamP1oE4tHxmBoIliNSlOIUkpjShIj8mzaB4GpWfUn9+Bue0p
ncBjGu9vExirG7UIzWxvbJ7OiymfMa3K4TfF/wAS6ifOCdujHuEFEsFnad72Nagr
tWuxNrbeg9OQhe5anKglnHUyilOJLA+guuk7i5FEon8xWPxhixSivSF2QpNqtBHk
ypYQKwdw1kX2RXxS5/5Hkm7/+ZBjG+Pvt1iE/Q4UcyRtQyCUXJvxR4i/GuYYMAqR
3ByPDPpDSNFH0CNi/VpjvTzzDkU+BlmT6+3ELsdlH2rQG9jY6MW3z21nPbF/lJjD
DbH3k6IlSpwWOw2Jjl5lUnH8X9zMraHbXjIKeZJiSfngvGfKzsZTkfnANJ5b/dqD
hKLSxiv/2B/J9VQpct/lJ79Y0TW1BzVc585phAfZpkTFYo8+R2r75lKqVN2iBImg
n++81wdki4bnLlKzv3RKN5gryMW2Eqyhp51+NOk3kyYvar6JxpGUXfOEBPUbaPlh
s71d23sFuWMb+S8nW2KVdw3Cwx23eQnvs7g5i8rCBg9Jyd9gVO4QMNJCmEr/oB0I
FU426SXbFZG3rYvAEwViHgh6S1Zvw/p09tXQ1XYkWteZTTGW9EHNuitUbkXX/FcK
X8vJN60wAAUK4CYrwF5Qqsx9h1ond6O69dUlffjRUEmWNzd/oLbkPPzl8aBfcaLr
Mq3hjNTMWJ1jHgPBLfxNXGgSXkYZPaoLIfPtaFeM6I+2GzGDxKRLoyCIkUtLiOEE
DhzntJ2kdosEIfDuY3gjmhI0Bxib369ic70C6VBuICNdGmd11vB2X7KZYiwlac4a
9smh+cfNGBh0YR+29CuPA7ji7YEZpSk3YPAqkbOIHpYj23BTrc3uIP6fFOka35gr
7qzsU422Jv1Wa3geL5x07IXs6ejGLPzuKAighN2u0j3Pcjim4EEnb9JCVzSXYyyc
oNXAWpamnkKj06+gA7iPH9BnYWbX8Iq4xOcibUIuGWY03b/mBRbhL/7K5C+IIjkZ
8rtdQYyDvu60o7LrSd9YjhvlxY9kv703fTn9sRqeaFhX8QLH35C+uRdgTNo62c2P
/JLvOPQSUUr95MqLKbtOne6cjbCeNkmkW5O6gI7EauEbqqPD6LFwcpDTtNWX/qE/
AdRG5lrNkE/a/OGaPWg6BWAv17aJLMnFHAoAGCKKLKXj4pfv72iIGbUDL3FcjHqk
FH7vqu6FLYJfFBYsxcoM+5MSe3UlDLG/v+/d0bgUJ4KagJltpyF0Zuk49I5FIk3F
T/g5UZlyrL+gunJhDVF+1YcKJZMbXR+3n4ZvUzMyAh65vTc/r1BtDmjCzny73Hr/
C3WwHNATHXIZLcCX8ruiVPcWbocif5uDAzTNPfQC/k+lPx42xjtC/4RKkxPkOQu/
`protect END_PROTECTED
