`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B4m6BRSfhR+v4VBPTt5YkRn6LD0/lvXEg1GOIJIXoW9RZaivXgJ603yDny+j5N3l
CJssGWjglzCFKx4oMIPF/gX/8+UbzWms8ScSiO8D9GWstMBMyoqLeuRRJT0Bx2UY
86RBNQsJwMIIBG6vIc0TKhJiLIHAUthrwvf6smsRU9AM7uMNI+AvFsMyx8DAFlEr
+bCHpKC/EJAsJy/xJuiC7eqiyd+AZoTQ86Tm3oH4jFc+srJZwJMDCL1qvkBgx36N
hx/nPqVWKg9jK0UWyLVnD9ZGTa4p20hvetPSJUdH1i2yo6KgZJlb3aksqrWkCgAl
vLJ5EYOizuSOTbQu6WDVxjea94DjBmvGRP5Iu4Wve12RrFFSy7vxjGQlaW9qvppo
hqgYS+nTpCWGJ0OXmXy5boW2HofTBqIuNz+5dLuCI2Q1/p5VglByemvQAMcwsW/+
CGszwpnnkCNWib+nSqZWOYblCOXiRqzwFfJzHA/ocojpR9AesgxrQg0hCvqEdU20
Fqgdzzif38QjzG2CYdIZwsjENfvmF7CtQYD4CPmYiQIJValEe4Mzu7Fwq6fSmvhW
yHECEPPKn1FQ2Bsny4RC70YUY3O1j1h0ZpPPF2CF+JCafS9AtoYnLEKg7sBb0byq
NqnGuGGHK/pS3MOUC/L5odzJ16JRz4275zljLav0D0KgNR1FRtUerWDF4XnlHr6M
8C5gptaZQAWTOyf8J5K2j2VvZ1pU8LMRKf4pXYhU6/H8KOytUcAd5SF9tWWQA/c9
SwT/lxmuh0CXDevUaXswIAHFGP4MjdclVRd0YGkwb+n+sigckNleym9v7UFfKT5t
oet4D+N2vp5qVpA4x3yLV/ERozXAvHgDzCTjVSIUg+0c1cGkcKcAG/2gOXv3T2x+
VGr+qdk6He69XufvSb2Br8E3dCPDROXLKWTXpCeq2BLf6CoG3qpxILSF9Va4urwI
EF34qSC9FchiSwIS/7JtWk56fGCTpbo9niXM7ZHSiaUHUJieycNQ8gqUf2nMDhhQ
Faza8Yd+GbxhA6FSXEFlsCVv7hQL1gPwrUh2Rkf0ldYINrVkt3oE9Oiak1JyHEhC
4ucMUoX7gAXERpBbM8C54waHp7zCQYwVPypEO9CrhySZ8b447PJo1ZzWQKCkTF5U
6D9x3WHM/cJhwADt2hQmLzBm/CKLzVUk6B7fcSr0XaMdiEdhDx0/DmPBNfb3kMrP
v6fxtTq9IVJ+WHTaEKT0eUFWYDptrhegt9B7f/RGwBUEeomAGtpRZ9Ea+7fLOKey
wgIdF3AMTntpNi4S2tRgdXI3aUz/t7U9LJY2+eBn3AOKfx08ZU2EXcWJt5wqwSYN
uSnv6YRsTfIXiMouoPhM0be+lVBm5zZ+6+YoqD9ACRtLJ1iXQ0ABubxs6TboM3K7
sj1dYDaOWV5T1YuMMoJ/sEYRyavoH72VsRhp08GsOdLvz60DcBtB6SFZSr5CCLEX
+7oxVX00hWmBY0uqNuPUi9DUZ1WjypJetKC5ggUSokDaBhA3iacbYVRhddLpiU5o
/tdT6It2lzGAe5wRVRm0VouUolomZ7cZZuC1Mc51LJmAJ3Z/GliaqTHnBw2tfrar
1p9mETM93DNxrPTQ2qjydGy+PHp8btzlWdY7XPNjS9Jkw8poy1qaontw0kbMWhKN
2uJqic6/Y7SqcmaBcQWT4sX3L0SpglGTGBChqEQns+HWU1W4woAWuoe/XnLbObeu
LakOgfMuzKfWsSWlUqZaypRN+Y7p6nbHTCdl2TThNJM=
`protect END_PROTECTED
