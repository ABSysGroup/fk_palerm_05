`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZAlT76BG+YpyxdHrupGH2BmOlYkCRHf+8JFPZNpFfZwQxuc18juKnWywX2XdAfFU
tgHyLhmEEce/36Q69MDIXP9Ow15ppQ8nsj3DrE54t/r6TbDYwwt2fXTs2qbDPC6F
C4UDOrbZuwIP6rf92sIfAnoz2ns7hBPAo6EIlQeou7Zd3cq5gZ6iq2MXjOwZzdO8
lsvMNkaQAFVToFO+xGzKtlW00H22EVFh3D8MW2Uet+gneub4eUMP5KWv9N4Kv79o
hhlc9Di7DIDlxg4Cwc1oZ8TtjcgG/vFDKEqs8QZ5PNoCP2u2HLUy+S52o3SSffJt
`protect END_PROTECTED
