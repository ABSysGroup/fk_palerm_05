`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sbGbyiELs9xHgKkfMBs3ZpT9jCINiOHV58D/kbywmrry25DoKTi/ht+kpICXw+ST
K+Hh1CmnPFbsIIjr/JAbESSGbH0+JwhcT9kdMGOpVXQBkEaXePQwCS0qJl6HlacG
lkeuIK4DcodQrl7EMRudA4Y/nzPPDfYR2TYhrVIuB8ZqBcWY3lT1jsPCrLfd3LSD
5pEWJql6swAuzAiErTn03+WGj7hIHVyg1OdqQ3pryHW9ObIGqV3R1bsJk8zA+lA0
xl/yZuwJ1Y73BXUXmURbYFRnmUJMd8IFtpsOE8J4kAttBqLTBWG24L168kfoLbEx
z6KePmvKnGI1rtOW3XoGiLSbonynvJnPe/Kfroo38V/0xetT+g/EBmMnaB993VM8
`protect END_PROTECTED
