`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ER+lFRz+sCcUrbIk/4izC+Z1foUU+W8XZay4sm9vrGi7ZTvvT2N+o+QXma/wihIE
fbVEnMQp+K61JMuUxW3p9f3ZyVwurq2TgltKYdWiEcx8zcHivuE/bXCryJB7VU2F
2olRCAot+MBToLP4/3NxdmGJkw8nRBBRTj8Ak4VFgMuWYrfVNyKE0mPiRrYqHKsX
zFAnwZt0m48l9Xu6Iiaadeegu2byCu40n2kCaqiOaojcD96CF7ntjz5ry9k5z3hQ
x8Ay0moZihAh0z6kiCH9pQTD53e7tqaJTJwH9CNm4Ks8pNAMkp8uvmuZISsJTK+k
dklgRvwZNzdNEaa+UmSUA/U2UW/RXRjmua+YKgAxcjuJxOG6MDEpVU3n+PchJ+v6
`protect END_PROTECTED
