`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZG2BAgywf/hPWiyfap52IXe9fBMUlAkzL/dDkyNjxju/1gln9Jvk6G675Anq8eIG
vwLH6g8BulkKV7r9oYmD+9+Gz9jhEbeHYchgvnOY13BVChfOAw8pUOZC13K1YAa4
sV5Y7qgGI3wWqZNEmpYiw9SkZKJjK1xLKu1VDYn6fJR3mMN5M1k9Y/6JTEiKI82t
wlt34SrxRy9DjB9RjPJJJkUCD3t5x/wCzAUEuDnJ6hVI3ZTH8Yaw3k/YcyN+hgr4
ow12VdDjEN0AFL13xgZbArZgOnNXs20yYDTRRl6NCr9Q7PjwU0NJu/6n+YcR9QHn
2pD9+SP0d9ieTdnx4teX2Y80+LE9NS5AZg25JwQN3EYidtZYyWzxFW5iUD7/yUr9
yo+4IRjFawZTEZbhUWRNxMYW1H3B4hgoEcFn6VX1/72dkUEtKnkKZUaf4AaeJPEL
nH8UwtakrFmw9Ns3D0lg2ndM6i+Pf4RqSX7caYYACCkEHt8J6yQP2qOsZT1W3nsr
Ff7wjBzpKVr35xf8DuLOy8WERbUmXCiA2B2Yd1NNqqpKX3HG35WSDKRqHa/UDFyk
2XNLrocPJvVzWLBRwv7OXFGG5wwjDmfckjMzvzTKAL48lp97p+/HYcsZoZQKky20
WZjxuvULESOBaFJR4FT2+Jseps51CE5zZjsmhhSjBkuFAkqj9vFs9C+m+l4o83ib
0ydn0wqh+XREZQx0b4Wls7zmYwB5cRosvX59hvqc1nUeypvIT3yXenP5xSOpQT+C
9y6UF+jMc95FaVn8IYUqhAmLlLn1P0+LEREJ6I6WqWADtzes06pl9NjZJ0cStsfu
wjyxEFYfrsaoZmwC1nsL2XDzErrf5Cfqanh3e+syh/oXduAP8+ANaEot8DAOuWFG
Rq+zAuXQZUFlvMT5fzYGveGtMgx0ikxs48/Joavootoc6Ijc4LamoekvO9xjOQ0j
tHLI82NlhdadRvWBR8nE8CY14U4lkFHRIsqqnKLmeiA79D4FBG8zTrqg/q3MDJpP
r3ymHDOt2jB+Iv3qxj7Helqd9kbd7fN8KN4lIUu3bCj0UlumL3ZIX3Dl10A2XBrw
HrmSaKVJFXj7CxgYcqoxlBqH9hBkAZzT0hdt9UJ/9tIFoq9iab82TcNd/oUcWGiX
zH5+zJkCdhemBepUVT8nV/pkwRxDUUUZhqurzWnUF29pCk/qYd4K8E+37W7DVLIr
deqz5vhVg37sT+50SvCc1RM76uGVLGDpEzF7OqYocDc9uN4ErTpK5W30JOaCBql3
fwiAbn1PBIB8h4Mhw4P/1TG036L0JBUpbLR+NbRuZQNjQRVY2qozIyfDlw+oZImW
yx47deGZ0aWpdIL36P8WmotOex78N0Gbbt0dnwugr1NT+z/ZB6BUMkfBABJ4+1cP
udKb88X0fPGhRDz1ILsVDV4r4lxcTnQmjBNcxKm+/lVvqTLBPK1rSlqgmRhzJbQh
EartzPZq6nMQcOu98yMlTaSEBbOdmixvmxg12Y7e5QH+pgNJyQp9727ZP+7T3zpt
8Ye6z4gBTDf6wSmqQHdVlOwk8T4WEo0lO9drk038iwUC6AD54jmMp0r3LqK/Rfta
PBA+gwGSPmMnvOiyhBUfyu0OfZYjOjgX0hwV8RDV89MNDAzCw80XkshYTHBITZmI
VvLrQCW6D6OwMAKdcqF2hqx47gT9Fq8vt7/vCFLlTWhGm/yCIon7xfwJE3lJiO4u
/D3luGEKMwqHRPV/2LQ4gF8XSTGjVQGhFi3KGCXgYhQ=
`protect END_PROTECTED
