`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k7lQc9bmdRUesrPbVTN/8TzesUq/alJokgk+iJkpoYU4V/hOPJMYiu04OuvHiBTC
ENwOz9qb0J9stOp82Goo+p6OKx4jms9vKKOUjRT00WWAAAzoKj8JjyUY/58ihhb6
eQ4QOwbZw9eWdDpBA0L6BaCgAwEBHxT7N9og2i+eRNrPSBvaQAzLABUOEnzEw9Vi
APQ2nKe7uMT5GvjQlyoDn/WONaoyW7+VOhppA+ZgW5kGBt78UartY3usmM8N6PBx
WdJQWihS7BYh/Yuzp6CJ3vn1KqocsAjluLh/bgIU2QP7XmM+Rq2OoDBB4/qRlKps
+1JcDn4T7q8fPM8Gh8TWtaxw1nHo8VuaNUmAPf8RX8I//Jj1YzXNB329tzF0+Wc7
S58BrmMuVpcKfid0m45jIvyzJFlFGM4RL9w84ZnL4WoDorr+d7xK7izD+uXYAKnw
S0EWGWTjz9VVOd6Tu4EznT/FdYLB3asbCU/9NLwZQ0oRs42yEJfcZ/b3wrKtuM27
1OmhLm3yQ/tCI9p2WwiGJc2od7JxzEmpdY2qNY9AF0lpGGbCTMLab8siWgErUCOE
f6Zvd8GHwlXHmmGR9H76zjw6IF0vgU6yNKnEVzwHsQaFWt6gRHfYfWRbYxXmNsMo
eHoVoaTGTpx8YSjryNfhua02LvDGSohshVKw8054yy+ZgoI9Okq8gY6/xf2nDlcT
ByUssFg0cnp6+XQKhz5+HkdfLKl/a+zKv8UFEZHu3ndfUvdd90uXdDrnDFkjbJpm
swALZrahgBMV5KxTMkv085FpY4dQccR/4aT67cYSCXv10gnXKG3eGvNhpKt4o6PB
TDXwi1h3gfW3WrSUhKiWbzbGGPfZHQtj/Vab4Wq+/CKnMLU054UCCNVvYdxhBc6w
L9Sh/Za073usqPoYs4KsJ1uZ6Po/5eWoeX7RP0Zc6UzwaaK8pDMgxWGk6By4lvXi
EBRiS2WzC5fWIl4jJYZU+owFVfDjEy8seAKfhDkoZfc=
`protect END_PROTECTED
