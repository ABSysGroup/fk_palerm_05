`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R975u6jAqTgR7hFUyOEA8wLwq7XGeFGQlrj+bDbS8jPgXm//KzFCmFf0l+7AUOBg
uNXNHJv5uzMNZyJ8l4BY41VmIX3wrD+3icOUY5MZJkA7LHlc0xlNldukSoBjegqY
rAJEAbrI7epqikjMKBNgAOr0HCb1sVgFKz0Mq5SLF75WDk8/+sNftK7J6GYkwVr+
l4fbUgkI6H1FF28MMBxj0txSfNC4VD9Z2/g7i28jmqDmKvkbzIwkgO+Ck7nRw8Fy
/Z0C88vqXaEkpnz8d9uNCQRl1JbkpZJjf68SjDPttbo6sq2z+tuFKobT1fCt/tPx
bhKkk3cEzgOk6RcJx9xF3k39HQzeunIPSyEVtPwQ1QRvqvUlPM4C5H4ci3T9LkgP
OlkuczD5PoY3v7ok49MiZx7+vQ9SiDlohN6UAJMb9jn2RwlTtvGltO2wjnVH/xml
XEfglBpw5Xhut8dbtUzUwYyHeo3H8v0bM9LLep1pLtbCxQDQ9jETEJAeJ3HcHVu+
qoTndVGNHuJ+AvFOlUm3GY2fLgXmQLzkJxsOVKxd06X6I/QR5FVznvS2cSQwgJXs
nB+85MmLizLnFsMwxl0toMv92bNAeSl7zqbbow8C/EJFWQRxqrLp5hvwRWXglcqf
9OlvlHYe+g+AWiEMmcIgvKM5bhuc2Iks70QHGItIxviBJeWlXuO5Oo9Yp45pghLl
k3yborvRo/AvNRr+RSRUAU2y2FdlPkVYxx+8jjvzPaXJm0qzcXg/+Ym3BI0tvfHH
CCKLA+D/9mk5fzAZvrLmyJxgv4flz0TEC+hO0Kft64X0aORcU9ms1xYca9RoXuQs
/btQgwMLdC2MtfL8kP693/6dOZ1Vap9YgcTkWlelwe8ZfNrgatqFhkJgaKZVtR5a
qp2b3zns0m/NYjFOfAGo/R5/GqcEM6d0zTvLXeZV2JK4SWFtX390qS9eg1G0Dp2y
4SdkxU8Y4gTHwupoXMNacSeW0aAGhTPCmUaGlWCUdzfDY0rc9q9E6cRayDK2qNyO
3FgoSIx7tlt18QyCSd0nmUQ2Ko6/icKogccNr15eI8eUnc6SasQO94DIeOOFRNz4
apEKOIkLp21En0YgOuhUd4SqoVk3xQNb8eFY6jujNx6VwyX9Dl7v9ITIwnNGdeSa
mrkGoaLSBDr4X8Dgmq9nOUquPbW3/BMywIVO6pMm/xcVaJnkmgpt9Cqm/etR5Ud1
LmJbtA0zjdbqZt/MV7ZVSIAcPfKPpK5KpMT8i1E5yD9gYIAgonifsUtuCm17WpDD
TRp8PVqbLrLHbNWY/WD7D8KMPH3fRme8LufHY7VxdNVPjaDgPq7NTZlyS9rdC1d1
JGnoc69gBVZXc54XkOu8yAtTKnlmJvtYqIHjbxAWFx8ivjZTwftfzN58+6AA74PP
Qcyr6s/jyWSKWpVvMDTgfbTr5ryQ33c4HGqgpqd86O7b3YTqMHeIaXKhDrg8RF+l
R5A/y9IhwGPBh7aO0r9LCddF9SmWXoXBYfTfXNyWdJuTcPhgv/4TgyE/p0k5JdZJ
kYWbpWiSXnMmdktPIFCvm7mz0lnb3XbY5IkCYqFv0Lw2Sr6awdbtywK6qwo/jZAS
0L3gc+030le8ZDV0MVi+/5uuzNBeMF6b0f0dtRmdfQPuKddAnEBBgmmjvBxmXz4t
rlMEC5LQy8EsMorNxwaG+EgzIh4dvusghhRchpqu+VUbAmrGs6m7AtqcJUHpLo1k
6/kGt9PlpBzCzkYSEGoJBxc9a3L0z1ZOru8GFUhKlrOxRPeA8dz24W+sGRSMdkBK
iiFv7r/0gC4kqQPeEjKFuJAj5CI6+tAtOTk3/U+bdOw+td1lqW1Iao8SfRvPdtbc
mG+YDrq1QTmd36kYunMGm7v6y3gYar53t3q+Nb9oDL7CjyD43kLDbcz4a0BPyZgR
67mkU8B0v6GElWB57Uz4UpGzrZzN3rxL2c+Chjl6YXS/IBks6Lpv2iX1qWOUtClh
NPuxrKVZk2TStuGnSeSrD/gOMwg/BL6kN9rKcULUXwy9uhU3g0b4XGrNlKwABl1J
dNoqCn18AifGxaQn3+4M6ZxeAxcuO/2gHYvlR0+Fsz1wevsO+6q4xXQ0fLcXNXiF
zenkzkuKgkGz8+PGkr/IdfFgLS/eN8pfoP9jj4/Jncc=
`protect END_PROTECTED
