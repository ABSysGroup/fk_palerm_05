`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y5jvBQxvS6bhN7rmOpAyao+fq4BJ7PxVCsvHToDq0cP8Ib2cRp14VMikGpknaSgf
3Oax/B6lc5nvydn9OChEu1J1hIoIA/55oCHaJZMrFpeC8KNLZ52nhpbUy36X7bUy
4dO29D7KouVto32qES8//mfrctmKpDTb9qqobwRGUsml/33DUepz26zCtm0ILsbM
RaZS+k/9AXoL3GdlmdGIAjRnl9tlAcf8lEfMNZ9uvMFkDc5fv8IHonDDb6fpwZUH
eCFJ7d5oNAdNeNqMDYJG3nk2XbHboNtuItz1X5y4Vx3D8KqF9fiqYiSRsIQer1r1
s40yWEJixO6UmnX3pOnD7q5cFQ+SBjtjJogx+PEy5xCIfUtnkivXG3lowjcBPZ+l
9E9DKpnXvulg8oWxRcGgoFjbvIQMA9X6J+97f2JyGrwxZdEgsRmYjXPdFkMBLlkw
vdY7pT7XfNoNdjOJ12Ych4j3dO1WYtz/iAi3wGHC5kAis1EH+2e1zyIJfPxwqYIv
Z4a/Bl9rbZFrv2ya+HuiRhU1Q0uu3zFzmHXFLYSFeTLFCgVnkvLx3oU9OnYowuCC
H3fouN/lk2jibusLD6I4KbVhN1GKtOjx/y8/+1AyvFRYKpn0jFomSE4t93+0aNF+
B9Mi43JPgr5mnoPtQWoCGv+amhiqLFtUCsvgX1CAp+IR1+DUNew8mswi6ZzaYUpp
uN3K9tljbywrgO7STFAOug==
`protect END_PROTECTED
