`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IECdIrkIFo9mpm8OsCksBEnrIzGK4IntKNTsuiMw8Ocx7Db4guRXzVqDkHE8/+Nm
hOD2B3CgbtD5kmLhS0UNbjW7Qm2ill2qilPwPPsT83DUP59XJGxQanfXoz1dnjC1
DXN8sTCOvpQaXJY+tTDqZyJ12FtRQejbWOJMhKVD3H0GCvoxfsYenz4hzm2wNlJC
kZjp37DSe1e9IOqXGW6BsdzA5dcZ2rfUoQAS6VEQ/cE18Fnc+5Qx+GSzOzML4R2d
MuNgxibDFH6qtUYgeRZ0uE7l8ARMSn5xM26XO+HLfrjwxYkU1XN4uTrGqxGQGHjq
GbjnbDj1fyT2GCMAfUWmJOVn+8DYw0tNMdYdiuiIBTxVksuhg432zFilIJLCK2Gq
UXIuUB0sg/lry1lW98AvoN+l9Iy6UNaRbHIyz+NmsLI=
`protect END_PROTECTED
