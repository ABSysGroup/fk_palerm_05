`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PP8ploZ2uqWcX3eQuIh5Zss3fFMAYwTsmZu3mv+jG07FNw2UESJcLZhOGAtaR/E8
cgDTwYwqO/7a45+ZDHurqtq/+2OmM8qxzlYyA/kK0InVTlZvajJzYSwLF86wwsXv
lOF0hAzi9SoQ8gDq1Bc2euVq2pBGc6eUEiVkA0SCdcHouK4S8y0XRN4xmVZxfdQv
fa7IoeKjHaUQesyaSMypCeCCTb6Sb5GLmAP4zjongVcRB+mER74ayvqjzlklyGzo
dlnDybFFacfMRWJrDP2+G1zz3+XsmLdxB/9x+/dPtSdpGbgtvXhpAsnbZvAiLV/J
4mFN5rLKEFC1CXSNTSfc8DPe9y5ZT4C2Lxz9oNQAhSLlbNCWG6D9eOCMUXJzL7Nl
M6UL3FwBPkR4sXiLgshEMA==
`protect END_PROTECTED
