`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JDPG+a+2xbBklsY1OowhSD3S161jGeM5birUL5NfxcSY0VvJlDer7b648qQ1Xeq1
r6gukMrBKH9BOmnGpI2vOnJIvmhlg/ssJHvoZSiDuAdfbIbDdlDMaEsmNMFZ32Dk
PafujUYWA34s5oODt79jAFBCV8L7/tzJFVvCQZfsIooAeeKys4bpTirbtRDCEJRA
4jSC6TnHDkGhvIY1LGzHInmhLVASPSOnsLwBx8DRxgk6YITv8Wv20f3LMmU1RfuR
Lvkn7zQYDqf6cdQ2XXOLvNrmwpXfcVUj8FZWcp2oAnF+mPWD88LBQ2zM1WuH/CBl
6qN415IbRKR0Cat7hu1S9MQMJVFzYdww1VsOPWnhXGmf7iiDapHf/myiQ8aDfsMP
`protect END_PROTECTED
