`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
noUhpnFOB51xh+OpFAhJXdRBNAwHR0UI2OX0aCMiFsTbZWIRlTRjuxd1meUlRevT
FvFAZmT4x/HKQObWv39XpdOz5JL9mwfv4MD6MgpBBxX186zsJNDIUeOsPd7oUSuy
1+f0gkNDInnKZCxRrEIA/U5fPYSueOfToyCMMvt0pSD/3Fw4kTOSULc6kB9aQj9O
0sdUSI4VQYgoPDHl8pZVenj5oW8jZj/qlfSn0UFWDq1sbp59gAoe1oauGh8AsSdq
tLeN7O17ueflJW81JlX4Pa5+pghDRG1Z1cqJE9Sxq8DCt0ebA2x7YnXWWOCkOeon
JRUe92fN7jKXdWqmd3D9iiq0/G4QXGsoz66k0EVxfDNPM6wy0RzV2frRraEeDMPx
TQEbPzzdj0Khroc+3HgzHxNrLagiiHi8PZhxJDe9kcmjt6bUEvoQMtwA8XTs5+JP
3m1Ae3t2PRmgW7JJVJaj1YGJ7T3XSRHWN7rXKt9uGes52mP+rQR7Y8leX57qF7Yn
Ro6BSWPpd/tDHbvyrSC1nB5nzMXJc0dnlG6JH9ekXI+SDzAze8xD4POupNmjMYTk
Lg4vEF8xM0lXUsGnJH5q/pYkXzAMGKQn7/e7uTKZKod8m8FzU4B8p7Nf0cL+5b2X
9aVqohnZNfojn73/ezD4mxAhrvijuOHWdKqKgpCYxtIJ5BXZJ67REth6mk8ECwyY
j+1j/Y4pIrSCUp2AK1RjZjG+z8Or9V5wXyAsJIyholsMtS/QXdBTfiUj/MLS+XDQ
dDTdgE1lNgcto9z3OhuSDtSR3K/RkvPo5At7iKa6I6od8G4f+q+6NDwz4PwyWahm
NprBLSPwxEaqebb4X9MyDi4s4HHgxB/taApudYSmufsDHZsmG3g5jYaPHO3bfkSV
6OTopUfzkxWhUh/zXS76RpTm0CFvzT5W+2FR3FNEU22MW+ow+Qaa8/XSjs4Youop
L3kaZ4p6Pqp/N/5rawTl40I6QSnmvHYBCoXQHlP0wMq+wUDNxIzju42yxwdtdnFy
2Oz38ZM5WKBpp4iCHN5d5MQ6LSYVIZwVn7yLWFJ07zAxcEoSowmMF9wI3aHjIFjm
WYY8XR/2x8SU9z7n80tVT1NkvwOo7BHxPi46BlRldn05+qQYjD23DhS64jn3Y661
fN7v7Gdd6+xYBVzgZAv3E9P1tye/7xC/QVeXJGrF5c+n3FimO2yV094NvAbel9G9
YUbhGSIf/C3UU+LAI/B6SverrQtLw9tfubqAqecJoUU3XUdeNEbLbqZpXz6YtCSZ
sCxNMEMfVIdsJaGscnZGx/aifxDiJsU7LEFLvEoX9r14ffTFW7jm3XEsvS5fWRsV
bhog8hvC197j8cNzuG7VgTePVQYwaYrJ4nGhx3tSMjDpZT7a4k/nDBYolnlj6qKm
7xo+U7sUXK3/BC7A38KJMrKu/zjq5XKC2imIzOHY+/riwY3IAiE/dvexjd9UVpcq
aS7DE7PrSM2B9DAwUTZ1VUFVp+6+K5/R5uUu7rM/opoesLflmVxzsr1ItjQoTruC
3QgO5tCWqyvSh2q8C+DcLVi2cTuhXHT4gn7XwcIfJp9ZluAldKsLocvRmnwhaJmz
vQg2Hc/xZglHK4WAWSY/OZvG1QozkVfC+L2rBI8x6UMwrAkPic79PDShSCciWvcV
BlaedcJ5JWtlRoa8nHclQRyViLbwhdrVYnwmpsiZL74yH1sk01pgWaSxdVWZNXGo
NUPvlTUUcQfjwtm96cvAcowlHpMYGEwFZFjG1AkXVBQghju9I+FFe2gAeqhNs4Ll
iKZIFwCxunoxZzFYF5xbPMom7i+asdJmUtL9bvVeQBS0szjkVNdW2UB9dl+KnzD/
WRN+1yVknzEbOLVuk/ROacHpWVTyV57QkkgS2Z58DOgFwZQxdGsXW9bzAZoR9VS8
Xw75TruHknUzhsz9jWTp0X1Iqo2VVue6maZjeWceQFMXdobPdoAqyxRaCyONELfz
YfjpdrsO3CxK6NPZpjVFYIXJcoKj4IT4rnlu/tuHdcLZhyJR19dvyDF3d7QD8u9R
4khgA+0ODvjhJuGt/nTXP03ggilr1W4kgBt/eWnbOLAFlQPHN0kENPylXLSNoRx/
O8ILndEjZmWW91Kdmu0SWiclyYdl8wtlOjkmubu/ZVHDwaIxu1SRWZMRf74qyyMR
0UEIjpWp389qT0MilmDKlFNW9smMdhi7hMdX0Qd9NRKSVqUzo9oGsx9+LAI1xKhw
E+8d6A/y0xgMnRPZhsCb6Et+fV3u5xArjU+zdrHzHl1/4m+Zn8RXeSLxh76/nhg+
2Ubu9+6Eo5/svzaBZlhyy+Wk8O93kzIzmwhPUqjEeR9EEWn6vihdZ2QwA4MedJM9
ac08T8z+hEAHesyYshhhtuxKuIT0cwWeGly3JfSnud2ZU2K2PF3onk/zXUaLaLLy
joWGbV6z5U1xbJIzDlF3hQvdtGWce/ku+AJcWV9EAhzsVC98+2flkA9J0JLBnfC7
CxYXeYl2g8W27sIIQspXUHq3TPvMsHwCtBAaHQpQ25bTYfsVe9zyr+6mMtzRdMkM
sjoDTROHtGFxas5Hx4zBsENjDzD5Tn9yaIFitX4Ob9OHeVkjXYoGGY6BEdfBfP76
iMXhbXebF8vVRvAerRST5omI6qXfqi070AmLcx5aMx3GSoJ3/jOec24BszHVayQw
6G7HOeQ84t+KNCkisV0/kC2Vy4nwzrqbSJj+h1GGmgggeJ8whs+1j/7bHWQPh7wF
XWPyj9EvNqloO86MlM8X2xI+IPXywfYB48NduHNPL1Y6EFqxt1c1uyrPABN66L0X
Pn7/tDOmEOhejLBO0TGMA6ZA7ASaUB1vqt6v0NUvSlP3HX7EWKqfVNYM2og54NNu
GJII0FuHTU8eBHF2SWchwtzbrYdWZIdPGG0DgvdaO1OEAvrZ9at3QPLvIA40oBWN
hfH6I7qVNIZ9bu1+U4VlIZwydJ912jQz8EARTuamYdlZRvidusNtF9tkHsynfM+K
ug2gvY/f3uo5dAuJbgz3qH4UKn/o5NUI/kvK47A6n9GHI4A6W4SRzn50Ly8SuGkc
tpUuUpH8j7IZYnKBg4wmeum1vLv/hAuUp33XjSgXmM4C0EQ/0fkSOye/EpWxrcbV
ND6EloKiGsV2isXA/EacV+TPSkB5QiApZdd+4ISnTYaEcBlCam8UGi0H0wJCHpZQ
MwN4fp/v1h6FKkO2SQltXxCHeKpMkN/CgkBZejUlaBkl9fWS+qkiFVQr9UAJhV9B
7DxjNVdyrs3MaZmcaaB1JMxE99uM0r6DVKhDynFhPg0SYrsMM3TVj2F0Ybz45yYf
1gTY86orQxrMsAd/yfo7NUA5cB1gMHLDwHk6oPR4Uq1AK5ADcK5rpTiXD+vc1SE+
LEY86cNMWE+39p4lb0JDjVdWF2YpvSbNuJNTt+hnq5IdIML6IaVrUtaJpWoGDK2G
2bu+MtqV6Z0vahPt6ekZSascSSf01lN6Ioz0T9EDSE7L4Lgm45psP1V/082bAe3o
gdr5Kek/NQmt2dI10vRh6ktT4y0DPSVQlah58rq3DqeFe76uR6QEKD4IcZwzjmt3
wx1n6MyuxoRs32fM3IVPuEfp/VcDvdjYxd3cSeB7tM1m0KT36w+M3RUUwtio6Qih
u7tN9XfOCYmLCzCdZTr+hnN2Iq3Gc9N/qvDb8K0SV2EZLLcO+0a4pqPIuaOgzTSu
WBmwHrB054g2TI/n1cxdNfxkTOkM0LUFWh1ojwbBVK5SP9B43DqvK07ZHEAUYzKh
8V8W2rt5cwyhHKXqxBz6dL3dVUsdyYPRC1fvnwwP8WqfjTUkf3uZHRT2dPTmE/Wh
HXZWiKZGK0vt45kFPwMK4LfH0fUM8x8YUCgnCOlxR8a9Cz/sR4vvAOTJpXJ9dbk7
YYYvqnzi/MTwzdzQGFubfY3pSQdS/MhqaZqNjHtPVj2NS1SZvIJ/YOsFVRSGDR7C
7cBV9ejMiY0qOs2BC1iLSvzwhSWke/fwydfmhpavH7sxAHm09+o1qtOHqf8wR3Gk
yWPyRouaTjLaZ/csdVeh89ms+rPfPpIii1cyhS0pCHePEBSwbYnvQW8ly/TkLFWQ
Wi9lNajo+NnbULSMrK9MiL6j5LaBvxOsWnuDIjmC6KFt1MsCRKzdOxhZgtXFZm99
coejOC4TmHF/tmncxsLW4LCiB03sDeb1Wga+2GstPg68HsJoi23Mkx9aPUkCju+a
qVov4Tnw+vCoVpbF6fsTk8hSQwQVCb2HnsALmW07eRJvWykylyNajICQqpjnB4s+
bxkxIohFxO5l4YrMFdzjcBtZfMOQtJvqa/foLy+UJqDzGbUL8DdHvCY7ajjPxvII
KZXkgtVowyo/eQsZg2YNm2oN//YS6SmHJ1hRkwCKqGq0+D5Ua3948ebBTVbAnq5A
aYsvrYkuVxd5B4L/OFjojjeqU5Jhw1zVVIAMCLxP7SImmpif4vEBfOjb+W9Zr7uV
zylFX+3wGrYLuCvbhSnRasB7cQglm37n41XLtTqmdzslir26/WdFn9XW91C0v/ls
rEyANTYPvYV3JAmIOHI2uNKPyrE7RQnfqoBcNu7r63gOH0XZ9hS8iXcyAvKZ4ngJ
ijC6ww89197kzK2s9xifycheX+BTXOCrOG6pAP/gPtogrc7cHY68LbaAVfxh89Ba
AAW4pnRYBSR0O2qvv9TAeXICyl8Vdd+tXR9UFQPqbZNTxtsG6D/QvXoHCqRbmPMv
tE+G+eqDfMVnTdTXjyHQs1Pu5DTB1ObCDTmM/bnLLA2UwRCx3puFG31pWwmhUlhv
VYd2fqgyKL3ZN8rEUol7TBJD6SDHajaAtOT9FR+u4cLsR8NXoHq191Br0DY3Pm8K
EycjpLeZ9XOIhnvvJwVqSRno+YJl8FFqQlKiBV3/7xogKbu9cOOMf9SKgJwFTmFe
Xzncqxf0x2FCQiC4DLkXO2nzGNnEQuJrVDpwQ3HwdHMtvnx3gC8zK8CNgdghBeeZ
bUo4Qm8gvzDfYqOKfh7G+DdDCTo0VR7KPx45qPVKdGu/UpoV40y6FZkOAueU8c9N
CMHbnPf05b9raX/T/HlZj3T4Ite6u51ebwO14WMj3LAeOvqmURRx5nBF0xTZ3q2x
aEJOf9W1fOnyP53HTKQWAy/KhMsKxFX59WS3HeAG8fcE1XjbWFg7Yx8TxelVj2ZH
OwrJmAdwI7oC8TqiGkFttNh+ZKi1/AK6BmfW5YOvqOUE1dZ8/M0cWHoxIXGvmHhF
wy2bZnhK60Ooke0CDSG01v7pmCXybnEIEZ6KNue24uwdg3wYauv8riK/6H9Ri/x9
3MteVGglIECO6UWQkkN6Eyn+9aU6wdVrLstNIFOyJVJX8f4CcTwIwRNhsZ6UoWRL
UJOInWcVlpRomAY4rltNgAT/bsoeltRAZmFYp/7o7H5KrhImW2ygPD33SIYFotGc
4aWO/pksQBjwwfVn9EIy+40Wo9DMpBvba1yrjeTIm5VziOEnB+fe5NpNQ0Cako8H
fWKt23v0cnyJNGfg/rzG80BhWAVAwPwnc0BwQeAXFG23dE0XuPulmCb5R4r0gnAF
P2t65STrP3wIVGKT4N5/l5bA9hXxYiO+6ocMZZ42LX1kng2FNltTnx1HORjm3qNG
/yvQigmN+yNpgebpXfVIbXAp1/M2HoRBG6qT/4gcAIVM44oze/owuxMNI4znMgNG
q/4RNifvEyBNsHu5jN+fe3gd4kN+xC5gYM1eKVNNFRaTqJuGiE33vWkjy0y+ZZPz
YxnSe4QEyeGCPnBxKFZ+Z6SBJTeeHUOArqqA7191NfkkvQxpRfCSKjN47nVU+EDo
7DHJxWl+ruujdsZfE+62IB45Wyc0kyys/+8Z8KBiGnDOSeXJF6PsVoahnyJzxo86
daZj5R6G0G5whH56onNj27WCC96Gd1EtwUZEwZW/0aZt4AFIpsKkZSfYsI1pc1I9
q3+kJn8Xvt8YN7+hZJQmdt0enDbmstHSY4pDC1xMyp3Rl1rQLCUzg+RCrjbKYIAV
9hlHAXDLogkuMcqY/SR5f4D5ggK02RCIeAWHWM62SphuN+iVscU5RFfboL57OVQk
K6rCtt9GMLTzL/Vxpb09DZiRTk8wj6KtjFigr0vFODN57oMQAYL95pSQKdkH97r3
z1gzKycpGN1uJ6cNZUJwI/hANd1hh6IVLpib4vSJPgd8x5sNAztxUemWocTbcgvo
NddceQK7KArreQnTpeqSuJutYmOdWVK6CfaWuqyklYAkCUNGHDCz1kfOUhnETjjZ
CR/229df0zWZweUDml4V6T4CuCoGjhOtU3cgY/HO3Q5RWKZI3MIm/dUznPdWvVpm
n0EK3i3vxEtkmb4TK/TWPda/zEo4PB6eSMYjGesMRRaX2u8QpezHprpHpEodhC9V
MN4/KHJdrVrtKIIUHxTTvQQLuFeo6CrSHag/RP/DkH1cV8NcliQDiahD7B+n17Av
QVzKpI6sjlOWAYOvvxcZmUannt+eOWJdaKEhLznuC7JZqhFaPfn1zJGzgGf/KAQm
hbqWIrhnm2xdoHjnoz3xnEnDoRloCMTXdkbpInWs3O1az8WpA0nNReL9H3XOqt0y
kWGzvnRmXi3KAHZpNgHMar5ydWZRvzHZjfICftJzeqUTNYbs132+OAyAzPS0CILs
F9rEosclWlhBtum36x+RUCAJOkECPhbhgZBeY49p6TSUO3g/9ERc79yGSk+vwhcl
u6CRRanijvwUAGCxPs5CGZvzMIhcGtUMccSgB7NEGBYh6KwfXt22VlnhvIqonJIa
iRTBMgA0BARwk4o5wuUo8Ur48zEzZSjML5BDj4DaYsJQsCeknsaY0IZ8eeaVug92
/Ax/aYk2Y3pudgBNU8eYtdOsPFL5u8C2uDhBx9joPoiRbo00u5akvPQ3XQpd0rI+
lM093oWx8Tjfijr4Exe/yRG8h+pAbmhwOzXjYfkSIcqGHZ09ERjb969p3/IP2hlW
epsRyzGP8q0ys0KzriCGZBeVJ8F8Tkt7u/9Mt48jzbsnzUutoU1AIu1qZ3C/IYBy
EM29OPJANdV5U0OxIUME/nJBuAppmLPVPWR2w+tpYmg0DJiBchRvzwX86x0Ni4Sl
BBMK5w1GqjzGUbcXWsN/UepibRh7tfThXgVt+vE4AA1NPnE+8ZxkHsE7qh0ea4N+
EIod13ctZ016gMT3M+qjPwV82UhXT1SXa3tcXKcvSWTWUTWq26exQtlXODHunYga
VM3thhsnp7WG4hC9cVJzV/lVc7O3ULGf4Ru0G2M1NdN0G/8WjuvEyHUFAUkxKTQL
PbX9dOcAJlD6amaR579llqE+UyEWapy3YE2O2oZ1z7InDa8RMm9zjGlFH66Gt+cE
GOSU+wo+YL16v0HKzsRlSuT/nWSE95RZOfGZTr0IoggR+CEvh+8N0Z956F7I0kLB
/8CLyxqJqyyfvGMDiArLRXfL8GtdcPZMYxTZgnSFPp2TxE1fFgG8oUvCdA8QUsBv
mbPVfJGleFt5bcnxAY8NMcmZhXIEnUpHO+o66VYJcC/SIzrv7PCJpLvFTlI+3Ejt
snM34Qem0tTVuaEao3uav5IUfFy6Q5ph01EoM797AiybyBSGUwELWeTxiMfmzVDQ
tdqqF6XhoAvS4tWCLmj517P2IOi31Noc8TTZcDlUQLNyF4dKWigIVnFLUqldwhkQ
O3cEKA5pvmNTy8svJne6kg7ZW8XpSzcd07JuKXQlsJmsqi95qjbIyDS9u+keXg85
X4O7uxbt8mBY7B82MZxcZs9Rmf7lOMx1Cp75DIkO5uoh/31xpalqevlcphfxGkmS
I2Ah9aq3hR1MtcXi+R25bo+nFYPfIXlEfX8ptG/iWUGNufEykQEVY6KswyCgTAVS
6Kbe3CKl6Sx/jjdx+eg74CGI1K9Po3bIE6jvQonJGFQqwvF0Kvhc4h3glofFd3vQ
g09e7UNi9URR85jGLoJegbMdPuILP9M1Gr2S59fNv3Vb7MtbVMolFJaQZHr/rRHN
+L6atfkDi3fH9MunPSomQi3MZs+4aWZqNQR5xwhkYHpQsCoC3krEMEX0K3ynUAI4
F8JNABi1vytL7TJdg11kWKMw7TZLG129kzACy16QpTODyLa2/MqXx8VrqCoQ+dpH
b4MQryw3BAIiICkL7wOABh+xx1ZS5vkczBc72u5u2l+AUzwe3qRV8cnR4I1XibIB
XFN+kfumV9EaC4FojH2cjK2XM8VdNC2H4y3fh9K5lUmxqPDDkrFe8IUY5JM24GlT
WKzcMN8v50zjPOV7rN1m4T5bE8maG63kBBPmgxCge51YPz9XDARJeAYL9eyTA5m7
tBCvKZadz8sT99wyQJEwvltlJeWrAUCIHl7n4eWe5XXQVDRPntEcDY+FW01OaDQB
5giozGcfMHE1h7+a0SBMvaz/rhTTasfojPmmhBorxijDKwJdOeqlrOr2blgKNuNc
BZqGQ98xhVjM5jJt6ot2IMcmyPaC6+W0+P7+XjX7hGwCZWfDrraVR9iEGlF3KbiF
+Kmz9bCgYQnfNangjKbEyWHrXW4do8twh0Qa2iBqH5nrlrHCt/0owohk0hA7615o
qTAQn0NKYdq+C075mkfZxM7M2+xSy9xRtDPbv9kqwMF/nh5T9Jrb8zb0n+ty2cuk
OGyIIKCRdsD3JJCjv7v0wvbFMb8N6HDa1q36leq6Ke9vimuNY1vWOj2+Y88OeWdH
n70B4xzjjIvEVIZGuwftT27M9Uou8Sk4uT7oOfpRADhZmeZFxJL/C54RHgPjF8s/
72zj4gK6XnGvjhCvbm6u8ajtNWudfB6S1z4mU8KHNkXL177ucJQmwdKVWRju/iIU
yWjJo9q35NVs23iJ7+n/l3tci0hmJ9MLKltYn6/HJhamIshuIOnVRp/l0UNQPqBw
sZaMNc1QHMhqc8CkhOkaVTXbbUnkoEsfWnPELNNcekjV0MObeMQYGVXG/di+7DIj
cwWOwI65jim3GoDC8CCGfaCf9eR7Mce9+4eKJKvAVNrgE19HLfhBQReX8ivtL9gV
NxL62vJRR9Rovxvau1khvOieeEClE4Dmmck0xUL2JcoevU49TW8DdUIEAbcjoN2s
f4USQJzArK6nslMAxQnoVJ+v9g2Kuj1l5Ks2qnLJj+L5Ga8GVdHKMkJcmc+LfqG1
h01wzfIYGIKOlh9zvJCpCFWw03FmIqwuW8UWWtQLz8+qyEJLJfLAMMSqv9mvn0Cu
gpAQtaHeOODFjVubZwsVsTZgLLuvWjmRHkZ8GEGRipo008ZTx6+xilqsZqaVb3eI
jNS8IOCtUrUwhU9ZozvNyIHzxVHbjUrHgEKLdn7utDHqGaSlvyt4FxpwQtC7p9H/
dBjuJXpADQXt8EvjtHPwqJszCvKnqGE/IEfsCiKjKLP3U4ElyQC+glb0gmNFtmkR
yipFzgIhV303fkLbPKM4Zv8y5fSReHb7pw6MGvP9g3fKvS9aDlEYmmgX6SPg+Ye0
9bzMkduFcEOxt16y8sQ42+aVNiiwSU9UtBTQ8/0z0cjY4BeOzIBlqwkRGSkS0xrA
g0JTRhqTFsyVCKkxmF1BXD9Efog+b1ymEL/iVXHX+jXJQAjngyrmjnXkAX1uE/Xi
axQWmkJAskyHCskOBydt57NCeFzX12GKGzn4WyiKU931ckzDpo9DFUb91FAjVXtK
4Wp6IRs/Grvvlge6hSvMtwwVs7NSeGpHckIRC7eYW6kSd8SN1CmvZwJpavVp1QW3
gMOQLnuxUkHn8H89cUlKYgV7LHUw+kDDeWY2VuHPQ0LJb+0iYDc6C2md15WKHZYn
xTzNt8o+8YJDQtTSgw80T5rcIUgT83hZm6vmkx6xrz+X/9xPGspPlTmDST0CBqv/
TM4QRwwXQSY+2SI7yAmHXVmtVFrF+Lh9BCwntCUYizi8kKo0IRtX/JfpDn3I6FJe
gtwSbTxWGfWRUD7hKtk9U4mnXAuDRcVGEAqFe39OaiZbQbU8mW1T6AmqVpeJxFk1
RFK8dPkkGqQ+mgBBSwnp7uSE+LMPSCb7tiYD1R5KmTDrcZ625enK6uE5fSPXneah
VNhfX+uyAt3Il01ymoeWXI25VRUk8MR410sa0n5UJcj0XHDMLIIQ/eTNrbZOFZqb
7Bc4QqLePiWsQwC1sMw0A3/I2YtUiw9hpaNO+xBXMlbOpIjwbpgcHa1CWPusn7uB
R5wTzdEVuW3qYZ+4g9bZVFAt+zOoqvcGgDkoqK+pdB8qY8lxZrkDrSMufAb67wfY
+VoP4IZZPVO8/BkNiwRLD4oHNexFTh37lLzG0ob8cUX3Np5gu5at8qelRbMxY20O
58OTSflaysGJq6QN2j/fkKkLTKv/feU+c1ORE24Vcc9NSPZpQwvQ2u2Na95EYWRn
EZ1+0ItINwqrYN5/AhwWpEYNRt7sGwMsuuOzrbWY5jQxYFByZP4Y0zg9gX2+P7yZ
Ts1zZrg7d34h4gpz1wk1NxQNoh7Z9tw4TEi+3DVQ+1kSOQPiyvGf0sDnYwAxURy2
FiwBEh0ZChgZGzMDlF3OjVpNIdjQU5iEnQNCz0kwbalUPY/n1lzUrecLqGwf8IOc
SEOql2mVswQc+h7heXKGXkhxTZoB1rfBUODZuGzsnPprOQqT9MkLkmdAJzG6uyKf
NLJdrYqNqqwGuwkkwFFiAJuDvPbXeO/7C9sc1lA2MTFR+rifyTOWoACXOG40emnZ
QBBx1T9STRj+AWxnv0NiniBp1NYrDrjm/TYlvnhUh5ubQfIfZa9EYzjEP3GhoT2g
R6OrmatqMXBDPEFPdd0iJAYKIhy0Gt/lBRI/JnA0FZk/po15tIA1fAZrKQOYvHUh
4rk14GgsBygoYcBSAL4XiNLXujjhEAvyyyLu2ZEdUCRiv3YE5tvIb9fASEE+N20c
ccC9/70KtdJweLatq0WjZJtk+o5273SKkjQ7baK4mmVf9NGa6lI91B149ZhTAFUw
FYNa8By7Ukc8cXuzrlrzltzN2cpe6HDcq6hsWkBMIfZt6JYFWl+lGgIyQvKc+DW/
fmICTB8JDu48Fzjy5+GzMrPKNqIyk4yz3fm/BTU6P0XjqOh3sbZcYRTO5VVsj9+H
fSNPJML5xBEFjc5CcUtvwBRhB+1zIVdmn60f/vsVmuxOCHZq6QR9bNMlqQUhHm+2
C7X7HHX5KOu9GHGL0gmdTkVpetkttE1THtadj5J/99Fah81UNe0vLLUHXb0r70wQ
lnPO1UczZM5ppYg4z6n3truscMlx3mRLiCP1nwn6f7NuHHyuP/KNdi2QGl5mhkfx
klo9OEcbHzDRw18O19JJb4x++vVaJcT+31gi+z1GQhOETig6DDqz1tgu2HzA2nSP
3WhcxwqbkRWLVdtNo62vE4xtqnw8coeQVO17MzXicgcRnlvGG5bPydZIFmr6GfZP
A80z1OrLL8fNtNz2BfE/ras1FLQW09DxisZO/oyAKFjxUXQCulSkCts1kUWctw0K
48xqE7qzJuQX84fG02xyW6Jv284zS672fnOHalJ9IleoVBARNtzqDDot6eqApQ/q
cpFUEVewSpPpyR90Q4ZHWe/N1VDPmNTr7bXHhuQGcHm9qZrumLFO6tO94rWM35Cc
n6mpR5PYhI81VBExUpcnU9HtpdX0Gdhe9xU+Ng1qgZe/AjsUFprwCBAb090Y/RPP
FmVuWSYRwXNHtMNcpp4pd7oNTOKMtqYuxdbQsb2EFje7WYevub+u30DU9VkJA+AZ
fgg5e9zb+CxY1Pb6es3nDeI0/c+R98twSC9jw2vaxIwqEWEqIimQH1BpqERoX7Y/
R1X+H7gmX46eeDDlS5TY9fnFRIXUtwMi++5dqzK0lIrkz93wXdlmomAsL9pWpYNe
eJnY8AytyASpzHdosen0CwzjAswLZ8vaSGQVoW/Y9fw=
`protect END_PROTECTED
