`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u4BhtTqi9X1zbSmBOZg/EcdIFHq3ZlI+ylCHZMmPKCIeoqXt0QFiLFDhua/ydpB0
9NQC9rSd0v3CaQ+uRV8TQGvgRFO/zamrtC9YvaP2gCR3fxzWWUCPOmnvwIo8fq6W
/ODu7BfW+Kv1tmFIeeWdlfW94+nrTPe7eZYiA/Wkrk4f5XHaS2mF5H1YMVq2nvz3
zNrChJ/KBYxt5qVGkxcGeY5RxjQJmCoWjhbzo4p3DftH1fGlsl7BXRwJjXYAYZfG
`protect END_PROTECTED
