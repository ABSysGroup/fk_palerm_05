`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KFpTxDbMFF7ZiCZw7uCV4Q+aDQzyiFp11MybZ3SacaQEi/WD9cfgY2ucmqFXiE+x
vcSSV4KPUl7SOdab0hyEMv1CZmz6k3+kLUDUv1+yic4e+YMY117nHY9x7pkNxaP6
JUv5o+C0vrTXbc/cr9vK6omm6p7pWhv0BaDEwZsODh8O0KWrYv3PuGBVcKatWYzJ
rRWWOUBA1rQMdPw1x0gIMh/qXhDOgkiPOEVxFdNyLGfRmDG5tEk7FU43uETPFbG9
GtgObcyiO1nHH7BJ3w1zBRZHOyXl891TW0WE9TB7YnIdgVrgc/HTy8p7R1ArjdRA
hi+uQo9JSLsfH/2GYHa3u0FJG+/Vlc1HAUS2xNVnp28Y5gnEhLFwGPtEY10WOuy1
wxg3gRk9VBPIRVzp/0mPIp2XHHN6pKZHPcPdMcAApIelGWWKFmjTYEZM2TPCaRCe
Z40LXEp2ZVzYj9dO+1W8DQw/ZhtMQXirD/PSwfEUuDS3VdGUggsOBqeYc8Sc5tuv
YayII1aGKFqU+GQFdiB2W/mUXGE9YcygPCfRtcmCfqgdzd76Ws8qEsiRYCkVDtEM
yxtKyXovRStofc9b5knuLk3hLy/+xTOC3RIzSYDBIT1FLeFqQWmq0QXe3KXwBi2U
y+JCqOcs5oN3cuktFU1vhdVW07yKUlEnqHNUCg+NU4xPDsY9AAqhavXlfn/dmClm
bM/o8D4YpkEw8PVJCmZnaD4dNJl725ylsHu7nPtwP+gfQ/1JzuPIk4eRULZIK6zw
UUF0W7g35YfXA4IzrVkycoWItNdxFAVmcunirg2IsOB5r9WxmiEGI57kZLTucQn7
vWHCKLjlrWA1o/YvsCNzGbPzxrBTDHXjqE+YOJoUszQBRbVlVL5LAFK5+f6Xp4J/
z0opl8c+u/XnuDWl1iAhPbjuPHgLYCnkP34Cb63K9ZkQ5fLXLoNcMY2yi20mbBN9
CT7FUM8TkSEmA75sYdugZhGGmDbSv5gOK+kmXjg8ARZLYgomydAITiDZFpcbCo4W
Z4wBka7kRbqc2MEO+sXzROD/eK8ZWSE5Bq34W8tFhs+Bsr+43o7o6gMTlAJ10XeY
Nob5gyKTgMv3RSdwSt8Sfd0fZt7AFgGTYNAxAkWo4YEvPBa7E4sRNnCHnAkx93oy
RSu5M5thYL0TkdffM7jxbz0nACnSTHi+c19xEzJvBHemp0XZuh/TAm/1JyRuXjNI
RURZmruN3pwFuN+vbKeYAQVKlpsuvHfAGfEUk0i8W0Vhwk9uKsYp0WAgmXI2LQ3H
FVCrk4k+2KQcWONUpVelDAhp0DmTFw6Zqz8LCquy7DdCi3QgSkhDHsFZsd771gJt
iXGdqVQLCCL2ofPVL5P+2G6MD4f5FiD4c5eI64ArKTXyo6yqqp5vHu3NKLQGFlR/
GnwOhGqT1NB7u7dFQyrB5BCF0miY+eYgxxQq3Pt+rqJlho5yDxEyhoWrJ2GCR6Yb
9c+XqQZOtRytfxWNUHZqP6rTtvm8g5hg37l12ZvDnolLEEO8Qrk2zFylPNl/r5zH
27DQrrJHmGJl00h0HUbNQsibKR4yAOr08uYuCUdrOzi8ghpQUxhsOJLMyJmuAg6H
V143MyaJkzjCD1QajVG7zkiB3S/PkyRM9d+V4ebOte0QxPWwVdZret3mpLgARvLU
XvG7BIZ0MhBOCR2IIpkWOSkZgs1KFbc530Kxj0bGVebhB8eOxunPc3nMgCBID1Rg
X/8HnkgSAsSg1TJdSBG1AwDep5GrG9nAlXjxFVTWK2Cjhm/00qgtDK/WAadoTva7
Z3ve9+W/PsNIYvGbuZhscKls2FthnEkTWb222f6eYV3UvyVSnGjGylPvq8/B23Ya
nykzS7MpcgrdKl7lhXlGdDudT+WnoJGgRMEruVokWWCUT4I+l7ZDGg2aqF76Y6h6
sBRvQilnFU7Ql46BL9gRCH/yR7tcz4HMJ7hY+bCF/jSVAea9Z01d4y76vHKCX7fd
+EtnelOVC+M0GfKXqs81m4SsfLko+PeuVa8fVtXVaHQSwYtWZW0VG5zWRJF3nkSf
Nxfq0UIpptZFI/duCFC84FRVyjC2AxjwuOlI6m/O/Z0aC76+eWxa0AffCSjUfIOi
ZI0DPOA2yOmXCosp5aJnjjl7Q0TuyOHl7tVRzjGVTxXg08DcZh9F5X1pcNFYpft6
dS8qS49qyTEfdiju4mWxK3gLyTJu/jDWuQM7tCj1u2f8jjefAO5RQjdlepYmre4L
qfPOIXDypYUmgT83DWvNsycdkJC0juxQK0Jnf8LBVWfmlP8Bij3alOJtesmmbBj/
K2LEOu2PRD32S/1iXT/cYClYoEkiCtGFSpeO/l8CHL1T4lyNa3uqGouKfbAhhzNI
pZ7dv3zeQM58CM2r0qYQAhEYcQPaIR9/HkMGwtmun5icdwIaIAdNCib8QbnWFPab
uM+6XOxrRPU5bL9hzHx9edC4yXB3IoB6ksGAmYYRTSrc/H3XzBv9n73Qf8p5MDlv
NPr0DB/YHSmt4DP+FYLZJ0SW3qSX//fYLzdiWvkfZJPHH4SVieiX9ZOne0H3Qqt8
iyW4J06AD/DBHFXY/7l3te/zKUjnu5NKgKheRcsKiUliRQQxR3dFVSDchDHAs08o
ZQ8q8jGB4UF5vAPi3q/wlSEZ8D6vk4cnGpDQT03R5HcGGXF+7C72ljMcBE+ZQYR/
RW01kbbPWfeskbVoRQambCk+69PY4/8L3AOWoOd/YCcW8bFbBHzy+eiaq8Si5py+
eXD/75W2XL8m0/9doUnmqBwyED5XTDi3xiotnu/mPSMfUFvc1Yuf39L0bTtbMpSV
fDRKDVaVllhVNShuD/dnyob8YT0+r1oEEglxr0/XBmjvi9c8E8e0uTt0Oz3qyKPH
k43TrVn82lTPASMhHaPfr+qCWvo3IdTUZu2frMwW0s/A2e122FQwDQN5mEdZf0jc
hUP6/qcWrclN8rNOvMkpqc6zhsoJO7g8zPEdYPDiXh2AN8VKUydmVNfGAreV4Ita
CqDkXFN4PHdNsjngTIKAOGYCFx4HvlnwYPLS30q7Mz/VBf/BzZ2QQJbvRMciqfIY
QgDsCEp6OreBiyFaoWx5Z8P3KNHzFbi4b/Etn8sJGkhZDv7UqpY+pOIXgR+nYSZe
qizdxmZ1wSBEXR6X+vR0iKPvjfXMERpXRB70nEjr8DoEYjujxWANDpwRsukCySp+
Y2h+Dsblx81dFsroc9Kv9D9TH3EiP5ht9uKMpb8OGUPXhaEZfC5l6T2hX4eKkghR
fA0Y9CTniCfBSjaTF5Dp969M6OYT+RQraVsadcQrSy98mOXkM9tQU8hfhxmrqeHd
N8nppQ5dVTjRNCzSBOMqaA==
`protect END_PROTECTED
