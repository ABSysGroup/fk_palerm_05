`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y5T/w3RtW7W3zS7btKzUJPMIEjgCzCq/3y85joREoNyvqZOBjOHsezIia+/jZN3n
LIN7fKGGlVpavH0Hcg1Fce7rxDVRzt3QqyRksD9nqIZCu/defXwav0QXUf9iVl+3
d3H1AGvf1PgLwXdkrMMYxUJxPZ7DDtTROM4+oiNmfDejcShsyi5IShaPPcw5Ez+8
DSnLYr27kw5f0lum9w4DtPhiwi6PdH2lX3FLUcjrm2wtrDh7JmA2dwRh/I43PLEq
dcbwfGOuRHyoFX9Zof1TKLViyJfWvQvRiz49gEB06WtnE9hhLd9b9PSKgMbSlXeF
pp6FQpo/iNo84YYeBusjLx46J9tnRd3wJMdfIBKBPy6lJuzuvadeF+8OD5QN1N8c
C3lcJq3SxmPLeuclcHa18lggYCMGs9m5CsFRaoLoON4lvlwa5p0aqd3nAuU6im1M
dFDE0y4F72RMFC8znRpEFJiWDjFJsZwECEAVdHq5pLErdvDuQpjtDmr+kyIIUhk1
jIxcvmgqW+6XjFWe/LZSdjZNrsdnwLXP5hlkNhU+OhEW7puv39raccWfBrCpXtNl
0XG4sSKflq+qTDmcqFxlF+wJV1LGJAcwCjzUAAoWkSOCKZRBQCACyS4DdNUhmSRd
RE1XfmfrnH7Q6ERFJCjCTMxJ4C5E7tDODkRhEr6XCgodYBsTKseESJBA8R9r4jg4
/d0GTj/QI29S0jZxP9IN28zJu7wnso80OYXvWdDKymk=
`protect END_PROTECTED
