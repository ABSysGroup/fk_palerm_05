`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fFyYebvJCJRhfdZXB2bjuAEEcm4ot65iPmoROUA6hzid/mOIwUfqV0Luoulsbd9O
qGuxiUX92weVmVP6+UPN9CXhr948lAWbs8zbZ70ATIJYDamll6vuQmzMovLtvDn9
SmRPCol/xCvH1W4RbaGg5ABza/buhVQnds45FW1/fYncNW5bla9LF08+ZJFbFA/p
fZVjq2TuRJVaLDfjWIFF2yo2AcpbAf4JeR68m2ji3Dq0zUCRCtoNJ058+GiQhsiU
r/pDGFDiHRboucPOlcfOIh0gAuwNLO4hLOwkguo48c0=
`protect END_PROTECTED
