`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UZVnI77PAAmeGn/oGiKtYsR9XdGF/z7nGoich1fx+WXvB3JUOcvbJAjuMjHAwFsB
NJfQ7+gozEwi5eHkJ6XiURFD6OEYwszwX0a4JoNbLrmsaZQ3kNeOWHPkjtHl56M2
dZz3NqT6+uJ+Yl4Q/u43XdkdX5zu3LZt5jTNszSvFuquFMgKpitF+CbfdDvjbVcQ
7bXZDDqtuRtv7NOpfIl1p0Kc/dxN4OpQO7gg7J5H6/oTK5Xd9ljJ3rX5Y/BqQLaD
xD5ZTBWs39T3YSMjth0473wrXUtOT7aZ8H0rBHCaBP84HEWhCGq2wWcDUn8cdgHY
HI2GL7zCZBlXktEohyGEEUFIj/2dxpz9UyGdZZw8Ik8dhaAnmdqr9wwH8n0g6ZvH
4+UG1YBUe9I+lH11EikDPcovVSyY3zGPZPVQjF5AXuyBUvNt9/uO12yoKFqF+DFO
dga+wV+kJ6IVQgDaEgHMQLtWRNzYfoRtTDM6a5g42mSdQcN8fd8U0PYL89QIig4L
MOGn652woP57frgOu85+tmnfvm/ugJfMWO69/scrJJf9HGh0Tyx5PrUp11k8L8n+
IRDOkmkKqvO1j4KzJ5KOv/5hjR+vzCa0uvJ2FHvS7UiwvwHdl0iC3E/rsg+53Dvo
gXM4Bbys0Jno2hgna6v6R52YAGlyQPGIPWag+wqx7Mm2/+FSYnDGg/mLbavMUciQ
6yrvzIkxQxHivceHcy0ZkpuQQa9Wmg6UhJ8oY5dKNQEukRduJ6Lozc0Efgl8cpgx
LrL3/fhZ+zdjguuKsFDHhqWqFDP+rn3wdJS6e3GGg2R+p9ICvBYjYOcugzoFzlEs
ZT0rUkYY/c7kTiNwsMMWFw==
`protect END_PROTECTED
