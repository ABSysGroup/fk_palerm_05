`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zH3thGps4wAnlZ3I+Mz7Lq+vX5bE+s1GNPiXi7Uw5E9Z8esraJ9OSa10F/DLtUS/
h5nPrZbE3AuEtuEZ44HIsJ0k6AruhJFE0QfcMpUyQNXalc4FvLEqitbRuFqmLLH+
iCekf4fKKYACrHPhEO0DdCo+I4VhbYx5DdN4CZBOrPCl5A5csTnxSuMqp/qh4Ajx
71seNVu61s6LEWSxEbENFkZrNkbfDKeZ9WuPluI/AW9z7jBag2LLpCXReMriizDJ
R69DWtDTJvdeFGjECLTIOjGxV0KeM5JBFiBqtCqLi4WUpL5O5W/otbrhOnpWiHPq
0HqWiJKbcSENYFWdbKMJbAMuMYilMBG5dgscrsXomh8pW9r74FiodZPDNbXi0ugG
cKhP8Sj24zO+rPxPIQwQUalxKvhNGF0z7O1lkT7gkccW+zNrLJ3nqzX9S8Dfir73
5OVI80WhEka0qyk+lNyGcXU7VEsLFyEjMFCep9ko8caTjqJwDp9VV4QhqmU0bEJd
4866FatIEOqRHEIw5z0jOZ/gokW30YW6zWwei5kJ6hkRwIUj6Nc2N5H/mTt+iy/Z
xzDX1X4nhsURyz5ZYIj4O2hdBt7L8p/+Wq8J3/AxE6sVSa/dLGLDYWtf5OxU9+rY
k9KZIPwu3DpnHHw2Z6kCGkr7BgGfreSZuUpRoSKbEOo=
`protect END_PROTECTED
