`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TiER6V5urWJlk4GviXE4LHYsfOczh0IPIrrIG8XFiqMCH6OlGli3G76HGH3UCIQz
0xtbQxZvzNmZahbke77XwOe7NMIaYQ/AdJJU6GAeyr/aWdasdYmDOtKIb8/qAbEh
T0VYamuNMZfMu0Z6rTugpiLswTdkh1dXwOn9vMxxBQhLGESOjc8eryD7EEzN+xbO
keU570Fs9KBWL7VnwQCUAOAdmA+7ADiDhKnfYQyBgVTNZ3ysMszqgYgFlY7g61vb
/nd6rvbCde4EPE3DfKrbMkia6PwMhJxEh3PUYUNWWbRXnV+iKi1sHPJ/uiKSe3Za
MUZ9G6JC452M2CibF2UaK/PFXOjB3TBxtQInhhdJ8e5PwCAUl0QbufVxQK2zwiEb
1u+WN0NsWkr2yq7LOBT6qcib+x05pVoJwHF0NgNAaeGmKhmT7k0kmluG7y9lmeIz
utizZiSmj5N/S5AOxx5apnCuzeXhEFUsXa57bmOvgYxLdZOS6DHRyvx1dRY7Yf2b
6kU+YslOyIgPxUoiDvmvXph7KrY/G9PiRIY5CB3hJs2wPXPIpThWjknfS18nuuvA
qLzL2PdXAhraxaL/syQvbHMP7PrTBJ3aRQhYq4yHn8V8Z87d5WVigwZnqoXQqgTf
JkwC/9GIOwOxCj/L5wTM8g==
`protect END_PROTECTED
