`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b5OgSHn26sCxuZyxJz6YqqeYaAIhfMxx6/Mf7esQCfGmRUItI7QMRY8ch0IVGEab
feOz7n3gTr/1Jymif8lOqpm55u9KzN7uT/aOzluBk5Ap99PvlpggOvBBGo21VHWQ
drNhrQvTCiBsk2qr6u6qtwbAVASnnG8J7B3iTo35AVJKQrSvzh8WGWVkjpW04olz
KoCZvQDozbXxGEXGKUu7eCLubmoVqSYWIcPVSAkjmDVRD32adtJZX4wBE1idgMPc
YsweDJTuqcHllnuEbBsCEsBAClYv9Da7Ukm7kU9YgfxDGSKx6SGpfd8EbYSlOLg1
VHGlg0OIjRN9EhYsqAjvfZY97qz+TvhmY82+vyFQDjLDzkIablFGqwY6VX1k2b43
2FhXRgli58vsdHMTfBytBvAJt56G7uDwYegcOhbi/cR73vI37DdDVsKO7oDg9jaP
GUwC5VbMDRLV6x1fAji1Jh8l9ARGK1vpb44ca7ja9bi1V3VsMyrHbvbbfnZnLZds
+64rjVJQhAPp8CvQAO9wzEGEkoNV+AY+wYiad7YR/zKqfzQo4p8EceYGt4EKN5Nk
d7hTsgGm8KGnmRyYs8XYpSfnkIiqQIfaBR/ExNxcvcoc32K0YhjYSouUM0Lf+kGy
yFCXViFjr0Kh2hqgxp1mKu1n0rO+M1giD8VtPpGi1Di1MEQNJCs9DA6djZ4tT+E3
eE/iUzqswXfI9xyA5xTiH7medWhVibnLgf9dWe8D4JMmR3QZtBqfdEcAnzTzAQWj
vVLDcUcMW26gzXloVEyJGQ==
`protect END_PROTECTED
