`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9N5INWMuhMXfH2IIf4C6vm5nLh1UR0mtLolWJuHA5hP92YthQD3TnwLQSpXps9XV
xmhAjmpxtbquupwdCk/Psmrn/3xPXCJHNV/8CyMXLlKfd+HChazp0IH4KOSYL/uW
Q9zHldahnBQqDTzmvihIC4ybHLVAYbyYTr84kGA0w1HnvZ/PJ+g///b8WGNHvH+N
+Yf+MCPzZvWtFqi/jsL54UBoFkKwGz5fpgwWgEwP4Vv4ZWz4muB93Bd+Tk38VY6n
Yn8SRSVKsA/EKM0ee48a0Fa1B79DiF/RVSEEzdI7aBV87aolmUIps8rG8wxt12Mw
ma4bels91+1L3wm82UQaKcpppmRNjz2X/T50xzBmP4n5hpxypZwUF6OPFaqw4U83
JzRvDZg1x30qLYT4BfMSL3288sRSYZKiHjlaNrOqI92fwM48XaEJOkwLFCX33pT8
`protect END_PROTECTED
