`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BOURnAr2Nw5/GVHsjjT+e8nVI/iT0h0Q6bS6Zth4fDVJrk9V8wdpplOhGBqm86ux
eDZajoYx9T56qrrXEh0eJZeFoR9sS4hxYSZQ8faPsmYtBnhUvaGoB60QDXG5ERrf
gdTnyTgy9szgo+uuZzdVHmrRZRgPXAJySkXlCkw9uetv29rxIAEMg7PolcneA1W+
XherHA/QXj20RaLaovdzHvTYgL5eXnGeTs3HJeOwrS7b8qbzdUJ31CoikgHvXpDH
1XdIZa/X1fzu3h0yGkZoQf2mZQE6lxgH/sWhcWRhV9KazvKt10FcoJo00axsD0yv
hBvTH9TwZPPAsQ7HLBUcfrc5bcxhZP9MxLtZqyx6yQibveeRJdVXG6q/UQy5yZ2r
N95ZkHt+5zVyW5t5PO9M/mqBQbhtdT+1AX06k3BM18gEpwhLx/6reKD/gQFYchE7
WGjNqz/ZBwhG5uzc1bKhTMiCd4m58VqJb2wS3JdgYqyzq8QFCiVqlOP3HgilIyVQ
T0qYefqmMhrTv/GWi6Kzw6V2uj4TaC8ZbwX2Ek2kSUCoSPpyo9LrmEy+C/kdOEy+
lE4MMfDaKKPIRtC8x5n+8OVGsVlJnxLFa9gV048LFbpts70f0DIOWl+siMqTsgUD
9lH0m4PV7n895dMkaEdWGAySdyfpMm15PcO/8DANlXKHGvouoLnC2A/oeF1bSOIK
njzTzoclOkO1hnFE/ZJPyLE2soo3TSKCPHmi1YZG1xGWjieWjqSkQ9LWMCXoMldX
w64KjlOtD6xTVyWtvX5X5ZkjLSfRb1H3RAkqsbu12gSwVfWYbGIAo61EBaW6DKkm
ql3Zo4rWoDNb/58PDKfx9WF6QLHursoPWvfBTOgjLZTQhV/dPHMigTp5NoE/PFgf
HgSlh+hAXPqU4OyK3v85my2FUM2R9fHEXtNB1/VXRfZweDqdlVAtadcc6PQzdP0b
HR/sEA0I69pWB8zvGWIFHwqmVmKopmdbMxuaUaBiXMZV4utQdriUgS0hidn4SKAB
UAwCy7Crz1KKaB62e+sZ7V+fYYQdkDNjL1VaD3LlFng59/OH/9ANKuTZtiWdmfFW
6qtmEk8gvc9bhMWs1CUvZa6880f+4UK1hpZ6fMzD9P8oHV4Fbk8cU6mfQLLuFLo7
qXsfVEQSewRGbrAKR4tjNZOqtW7ZeIv66+vc8BtKBPOlo13LOusQB1Tfvid741zQ
0kSewRkzagfuxEnF7g5WN5qaqfWG3gPWd8gnEG46kmYPROne//HK3/qSIXHU2H+V
q+1ldqnY/E8eFWRLmgmbwq2KsWu2vawGUs48grcTyq6ROnqulal4tJtYy9LNlPPl
FzPqOADFKlbV2Y4Qu5fzm5Thizvjx6BVt2WLnjxOVr9ENFQIsKLOLuULiRim9kDJ
WW1P8m0H7MxdY9cTUaVipfYWjOJLEz6n+sw13OT1paeH5ONa7ALQKULiBv+/Y0Sb
`protect END_PROTECTED
