`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pz0KYjytVgR+eni0775A3ayeOydJV+K9V6yfUCY293ybBTjkThGUwwNZLMcm2Vu+
3LuSAfA9Qtu+mwwuwXEMAx5HWZoO+qbwmsgJz66FETduG4hHT+Gh8il7wufDu+VI
6B8WCAanXpWBSXIehkv421PFpxDdG5TPj2gHiYHGB84kAqHZHvhGgOnsbdAwm6zC
q2mRf3ftIhlCBGF6+lY2UuTRS4LjmdVNC0j5QHzNEcyM/TnBfs9FCnx0XH2SET3y
40kCY3WMp3Io03w2vVg3X5EQdy2J/PaBxhlYq04GiBg8+AqYtbShiXDwTqdZFW2q
Ynp+XvYR/wIaQjQz3ZbYLV4YIg+ZFrPo1h3z6f2qAv963ABb/tslOJJBgvWeVmHE
XIr0UOZGtGMYRoZGFXTD7oofquZfbV9clZfIvp9V1hV3FkRBL0llYAknBC0PjYcG
C+sO5hq1X+EypC7B8YSvrPFa5d0rI53X2mmfFbAhN81zK6JHlbydE3g3WCBuCXaE
pMoh6QB5ytj1logYYRtIabqz4uEqdgYDT2TTy/Eddjxg8txbgNlhfLg/tcUM3TZg
Y29dLsxYfZwQTAe9Ss0UIPloPZ0NepO8yQH/MGe18YdwhgIGEMJBJeXwTBD34w1m
FmetaR/sQFF7u+chPu+iifwUy2AcouN20AkXmFIQqUdxPOy3LCojdCpBhPKGaqX0
ubYW9ha7PCFOHymtsorKfI5IHOVWARY67iPveunapsjiBPXhtkgX9570zEdKublA
fpa4c6oVfxWH2hGntyKsr4biq7GeiolDo10LdG1q1AjCsbjNsdsvaJcdVj4xBtpd
M3hLVytefCCNd/jjxZcHMOTpaNTGp/Tmq5FIMmDXxnC+JQa4aP0OEXsFgDyic4X5
CcntSKJ0aGKeIK/WUqMWbaw8cEBTIKj7+zXeL41xpn0=
`protect END_PROTECTED
