`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qIpToqFg2v67vEvsTeJRxwc6/l7iRcikYj6ctdGoz9pENgNYxEwCzh/pcXYSrMDY
TIqjB9oYlqfb9udFzCHr54kL1WcGG47u6xK8K+hcUbETyoyiUNw8KrmMSH1kKQJ4
Nd96Tz2iLQ1HtJ5WHKnR0E3Kf4K/70irqiTx0bq7nM6SwT9r7BZMHxOSGQnkiBfk
ahP3B7s+4Hi8kH+wdQzax8YVkby5ozTm9ihzIvlNIouoQrhx79urSc+PkWwJlRcz
JLvtCRCG8lFMNst46H3ounbvQbhW/OZPHpMAKNQGTpyePago4GgAT7UEQZd8gMIX
f95qBAS9kXIzZjsY/uvaiA+6NLEg7RLD/3PyBHsqxxZdI0tlUUm8R12uaxWWxNuN
JiMnOJ9HM5AIKXKR8iXcj6xEf+OxTpcYAyi6E4vjRX5icWlXpjDT2a6F8Lt8bJVE
lP6SKTC2knUfW0mnzrnZ2phjM9joZrqYL74YIZkjjiqBb/qLkfuu0wRmdyl6Ek8f
Qip/DJRMaC+gbh7bc3WTEhPnK34YGNnxz9Obw+sBRwTzrEzBNxhM0qHlHmRdqFue
3Xw49ZQ4NJ6+jQr00lEogcJJgymK3rVJZF3/sox3SxEGk1O2xUtjJzhaDjUT8YAU
YxV8YjqM88s+TmXiqHShqG9rblc9QLX7biaos4SDZDu7+uqpFPheoeMKBMxcnQ1C
3KCrTbinlMS5nIdR1K31Flfvh+MyfrBExZenHVQFEDILsKpJhQlUkARixyMEi2oo
rzoEqmiBJqGazP9BGIG+AtvCzSQbE0EKDpQifjwCHEY=
`protect END_PROTECTED
