`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3lfN12Y45Xf4Xx3chhfygIIQzdgltn0ynStxJQIDWraEIL6DwAmOfhhlGChLJ5V4
QC71bwxym/w8zB00oYcMOejN9SZT6ntDoqqi7tRzT0lezOatYV+ktbWlT+L84ki6
PeTmo7D/71hFBhxq/9Gt3vXSo/s4L1cPFdLOC9wdxjWlQRAjGl7YSfVwUfigEJKP
kfXxYM58sCZQnNQr/Jx+rSFKVuchvdAgc1jDNy5pcd8anJYJdfglMl+r8iZd5rNQ
eaSnu9COM8zSZoIRncn07BIGQ1aegaOGsHQ6gOqIAYFA5i9wz8NHgXA9JAwew7AA
TnoJ1f0mMVM/hiL2OaZY6O1TiVGMPlcfZ6rOOzc0LfhTsZGCn91x+TnW+A/1oTf6
9lKdnwNAuS6T5JnYh1vuyjdlNCJgrZ79VTONz3gzd81sIGFl6JjArDjnDtCirgX6
OUgI+nNdS7jhpqnXd8p8z/PTgdKroYZSDodFbgMH02b2xigXUbJftmwgp/XLUsC0
Tyb063+Z84LaXRY7e2cTH0F4uieYPHstYN+wOfkw6Zq3TZEbt7ERHHAWCSPej+6S
aSpuJ/ZzuPclkxOntafvxpLp8r5GQTVKUC1ZfGyQM2+znKAqWN+PI3zahZYc13Lf
vfEchof2M/YXdM3i0vLbAb7MMkglQlCD03Ylw6O2b4r3VozRuBbjSDzxVoGLgBQj
BiMam0VxtK3v3XCI2ujDQb7buBfYEaA/ffyYdaBb/QI=
`protect END_PROTECTED
