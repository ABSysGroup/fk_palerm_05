`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KIySlHW7BunAfgjH6X8KwO7oV9yTq5ajwON/pQtZg5FnI49kq6VC2lIEOJFFude8
/eUwA2kn46uVCxJFzbiTCvhqQDXgJsxGj048KuxfD9mDNvNdPH6W4e6PSgRhsQjT
uCOBkk3+5zaCXpTmLnoZBV7ThfLPMN/UrQ0O5MiS6QRNmq+nGTis/ad2CRFAtArG
rn5Iwo1ihY20VJXed2weZAkWf959Y/QFGKIJUg0J1iip1K6FhpuHWZ0WpRwZtnC1
l/052KPr3U0cZdd7NyGpJcUcUlNcPyHICWM5Ih4uc5VG6ljVDizMcZXdKCEqjFd3
uiWBtMYj1DPWFw3ePX3p8A==
`protect END_PROTECTED
