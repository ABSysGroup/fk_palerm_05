`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sgk6PRTqwXwWMnPFMqMKt+OdS1O4VU7Y1zOSAZ/v0Qc8d6mIKHWq2nwAgwDIY5wV
54Y5vrmf3aK0UukvqbTEZAu3jwqma5HuYo8hHzC5T2ojqvvwGzw/NXWlFo68kGRn
CzMZBPDn3x0NOS0adfOhXgOILdhrjzQv/NZ05zUsf0+XE2bODyiv0vVWj4kOBzA/
CwkEE+Qzkoa7hfKU99ifVOKH4YX8YWG6mhphvN57p7OhAuU1Ij7/PKPANMy9slsf
ekXmKd8J3pTwA9pZG+Kb4ue0hkQ8uWzW33S3TCbSL0YKQIRXHpiyGMT9MaWaq574
b+4p3Iti4aKwxEY+n1OEH6lEP5gpj8rwYm1A96Q+628s9BUYsRk8NMhq39k5Wr8T
RQH+QPOO4e3pxs7YlHqbHTzzBY0Gv503RV5YaKIiQ/IYKf5J6U1Kk2bJokBZv0c9
af8CU9/JIURcmQWyxWUScQ==
`protect END_PROTECTED
