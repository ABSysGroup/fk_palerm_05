`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6UGCH1x+g5zeK8KXDXYtZwXaVTQwYi39NHMyYhvnoWmAEtuqe7zAuA02NuM1rAmI
lK6tClu0Prwt98vnCi4x2hZaPbo3Jg9hXXAUfOaCMeohvrBxaG2/cwINdL1axD9p
OiFjKhcu3ckRN1srVxYeH4U8G4c5uqtEz8293gDku/Z+dSO5nnJFNFmv5+lt75x8
TS2FbCMYIl9p4iQUUTy0JnBTORPRHgPLCSx7fY2KSo3MgmHO99+WRBtEmto53GRQ
SpUalEpl8kBVNnbbCprVczXu0lp19qb8CWcntRs4Lk82M/P//fpV0S6QVz6zXPq4
MptQVgCmFhIRIPViRQ2y8GjAKWZT1+KSyOaRfYDUykPdaLBIS4hGzmSyeKDXLh+E
YOxolV/muidO34fxsCUfRCLJAMfMZxlJ8kOTVjjE6aDF0dYyoU9GLYAv7tpShYLU
Dl6/Emx6gMdgrOGELNzwKOXhjdpwHle3U2iGg5aUu3o9WxGp1E0gPe6Eb6KTlcvC
QZtpKH63zc1QG4eCYkl1UjzlLSVpmyDlVzrGEp2JEohfiMCQHJiX7uwC1gRgnera
yXe4Qdxp4e19lzbKQQX7wL1gbTFHa1CFw7pVvtHnSJifNvbsW5KDkTFIlm4lJ993
7TvwdKAxfPL1ps9hT5eEw52BKAKEfgKanGoAAk4r6P0=
`protect END_PROTECTED
