`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
scYNxyYPVb36J+pybLXfYl/lvfP1d3MHPAjAmPtI1e511N3it9c9zaoOs22bp0Jf
xlHEPPU8dQNVankDGvyWz55UZUxzZSI3qHMOCnaiHZGsZy7POAKjLUsHXCWzwQd/
BxxbMRhXJeLDfW1cR4nGvJnGMTD2W9jVVNQAKIKCEZDELcZH6+k3oFxPraxpIbG+
jDqU1EW6IAkRovMo/WdwqAhbEbmaZ4qgqVGuMtPGtOeTxjRvritA0aCanR7k7hES
KEUwSV5YirU6iD7LNTDcu7FOyGwAztLFEmL09I2SwAUBGKkPxWT48gbXB9KhI7p0
u8EUzm6yljHGEK91BJ0dFmVosJtw/DobdkMYCLaf/+E2Rm2iptWjfKIIbJ0DZZt+
NZ2Shg3/XBq88Dy8CcaU24kOIEiOke2CBLj+aPxrhgNoo6chSGjyWYxeYqp6tszA
Z7VO+9buRT3Bt7E4Il05axDCfy0eIeOfonlLmOcj+JcZL2TwJ3A0in16TU/x0t4F
X3vOtEMgRj0VL+HaXc6gZKQJIy+09YzO/cZU7MlevWOpbUoQ6yJIsiVJCZtx88+3
amIi9SrkDTLyiZFEAt1s5w==
`protect END_PROTECTED
