`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SqoS96+SKPC+kEAPfjdseZvGu7WpTkfUHX1RerLxPLHDDavqIVffRX7u0nsLh8PY
qOZcb8sxJFRwxrdkfo1Naje5hi1lhu9Cdu9GljGaJ7R09xsc0cEA7zbqii6op7TL
F5rP/JQKxK3iTX4xVOxf9wHevY+mScnszhSkaHH5OjVgCq0fbhQaTwmqQfmxL4uM
oYxcy+9gpWGLYM2R05FgGQJcgugddl2p8X81uHzZP3F1PDTysoYDhtStcWalymnO
cqIrNGPt4MC5qG8S+WsqdFWXLETw37hd5yms3uNb18IiBCuW9qvisZNKy+9M/Beu
4/3PNWYrTVY4HZgW5Z7B2y163maA9zbT2yV5Mg433dIz8Aymr8yntGktbBhNuojJ
PE/Kqt9Elxh/9EKmZH5aLgS4YAuPn242sJe32Wf7KfFKgSYeMBQzto4CwaywV4zr
phRjXzHi15yegT78AX8tQWTPrg1eWMm9OYMvpFl0mcmWLgmDMJn1mygV6R1zJAjA
E/zxCYrOXUS4VwFbjjd55SjEiWuPXlNNpJQFW1h1TKOGj3YfWOUGYLwMsKpr8R0C
IqsfTVD0eC9rFpD4nwGy/7TGEqc2CzNBIdSluK8SRyT8rvBQBKYAr80HmFxblOXv
V2WVGUkkAtBD6B8u7jWYy2O7JwBbaq+nXpfjyH6d7GvT43FnPlFo+fvXS+8prgtz
MuZloODMGMqab3GwYQypNVKQ7FTkWxj9lzloI3Hlz8fkv09qfDXarphe1doqvwRB
VZxxWH1jFjEPbb3WV3VMWhpukdYsgoUCysltJCv8lycRLTboJBAPG8K7dNYHjVot
CIN0bCHwfoc3IqILk8ZQ+RRQ2614IdFVzz0uFF5vzmSWy4WM93z/4mZwspIipV8c
cdVEonBNCVZIFumhs44uQQ8dFzK4YbRQCZdyzX1WSCCqRvgRIGXtkSBNA1rL4rwM
RerBRuKQBXbjWWx5Nx0/1kZ9sk2IPWcbTeC7wmYgnXC4iKW1uXvz93zgDsTMz4oE
JTNGBnTmMDK7O577NlsoWw/W27/BlPgcRihTCWXaLlEWDma9HwP3PH/6rtV1iXdt
iV2G5A/F5ovYPFVUDoclky6sytzWZbMZcy7HWN0odSNewU5pulzbE2rfLYaeBKqN
/JrVsN2QpgBYLmuQlYibXt4dBRgfJqNuFR9jw2OQ8NxKHcbilMe6BF76BJFnCtSr
mzVkghxs9AvBKU2FLYJ2ESEi6/OGG04321GSITypvu4xJJT6pG1KXAv28fpTVjSs
jrvo9NT3DSO0Ey6LZKygoFS+uNnFs5UnfxZtVgqXKlxMez0P26gMJW8/+XQNbaPw
8EDj8gXce9G2Lhvayo6s89rHlFSkcNs1h/AadDzTwZIfNFtPQb5q3eewFk4dhbjs
FZ9L+jD9KHlNGNJsaKBZr14XkrpNWKP/jIGmienRpv/HIH7P4mIz4i8g/cDSi5yn
80c4U4FuX5XZzZRxrqdvOd03YRAJqEwhteowVB7XM1ZDa5bL0OOyQGpWz5jKqq8b
IHV20/+yIMswx3lmJRgmWB96g2SKsYVr8AA9NJe8Zf8ibv1rYl9Impwa60LV4Uda
fTOe/kZz1LECEo6uc4ZjA7W4rlIdkhlLJmC69JuGFkUzQ2ESnrf+jVdvKi+QWK3v
cPE9AX4SUTG3nhbWldMnghvIwYlb4wwC5ciNAU+EstnlFBgGPnHigLejdTs2kire
+G6DpDkL1xpdS3XN0LMRUbBxPeyIyXjNq24/oVknjodKSb0Df5IDPpe0YPeEuj1O
wPTVFDn8m6ChHU3TgecaKYrzdzGnNi5dRX8pcUadGsBvZgjGYDCzzz1ZNTAP1qtf
8NcthewdHWazcrok7GIGvZ7E/SYh+ruU6Lz4wvhGBkOg1TQ3u38o6yAkvn5EwRR5
psVY3PllOpRXAjjs2i47vtkVEpOj1F4OCNgdRVd8t+sudzeqg8TSHal3p/rCYDWB
kCh0cnZwLmszawTzeAU0T9ndCvunbCPfY3XtwzIJZjwK6CZVfeZrX+iifgLHG17t
dGPsqJoxnQ9cCcTHul30SZye7MxJoWQOYUmQURqsIwBeq1/LyiXdnw+KjufWGqG+
AbM8UPbKBjFqDlF1K/UfTtt6AqLNP/j7y2j5clG6J5t0KZrQwthj5WzO+w1UJcVu
emPZJQa0BiZ1hSxnE97RggVp+FMKU5epORDjH8aa2v7wRDg7FA0X/rOB+LyXucPV
wRNVLzDXI6A4O1aeDO/UTVG/3Y1dpQuiLaDuNWc1iUIcDAqzEs7noP+SD1KLF0pn
pg9jokaD0dBnr1cjb0iY4lzsS3rOZ9esh9oUkubhgmYD+Kwr8z99Mlv7nDdXJ+wU
LoHI/pyzQR5NwUULTvzjpONcvgU7vgzhNH2A/v1n4lMxMLMdzoRueGPob+jGQ9Ew
Rna8SMtshj3Z2nCGklxCuVqYawzWcXDvuvZ+HfzsJnyzIPMbcYKl58l/8uvHayMI
5b9UT0QlPgt9MiJ2xi35jeJYzoP4A4B2Q67bUinF7mGx0vxOEp/I772qhHxo4aYm
mrSQpC+zaGUoBZLx8cmdRyBOhuc3DmxnNvZhKyin4SiqHFM+amqkTr7GInboYd82
D+Iz2byhXEiE8WX+8jEbCNqYeqjpxPM3fKRXa3PepHza5Lk4ATo+oWOVQ1MmhNrZ
hSGOit5PnxtiVns9XdS8Aqw2ibbRwCGFOic59HqJoQFhFIn0dJEGKlvbe2TyA+nk
01gQOcr5jDjC8rd93jLdJxXU64JMvR44pKEU79ttBn8Nt5Crhw6gPU9y+9TAmyVT
erU9sZiDE8welD9k1Fn3+i6+BA5WlFXEIzTtUAl7G/I2H7dzaarEmRLVixjYqVle
bYu9WIdV+eZwz3KFVXfjpP/tGEDkLRei2W84wW3nrIsbLrH5aUuDJhYGJCL6ZX63
JpFuRUu32h81mI63T1QGNBAWTNQIAAMWKSjnEHtitjqjYoEqHV6pN3xQappIf5qt
NJ/Uc6aARTje2aM8a42m43vn+apdwpSVQFz1U59mlj20mtD+pLlEQJCPLcSzMgv3
qJO/bo8avUrIviFljRvcJF0se6anG1H5KzIc1CYV666L8Wth3dEApr37H9sZvB+E
CwoYja5/qH4EylNseb7itsYsR2TIBQlR31jWy2TGOR1+fH46IcuUH11FKYZUOTIS
/ZINP6rKYxigT6JX+/3Zdnw3+tRNe9TU8gUISxF5lOW5NnWXFkWUzBGOSWL2pc6E
NUf8EOUxhp96zWCR0PLRuEdSdD8+cLSmhOfX/PBhVBBkRjvsviRKyWooBDxMcvjM
ROwJCL4ezcnEj+zrG37Lt7eVQbTJKj/VnkBNMYepaKqH1o9kEOsyRjJGn4yEG0dK
aYY2PggYQrneFaU1lySXXYXsW6WQkFWCmPt8jJeiGvZmhvy5muON239xRrQhjNC3
DsoFRA8mDoo6xd10Zb1Y644tvfsyB28QJRJ79VwLiqAjbuWnTZt9QNGx7pjveVFQ
7laSJlc65lNlOwiwR9Pnbc2ztRXYHYBJ1kQyzNXmb0d4GhS0YV2NTcneoze19a7X
gUzecYA2e0d1C7CpM0Sb7h5YnG17XiFRbbVoeBBVZiQ+wrhbubAJ4RwxxIcxiR0K
EaZVmMh1LSraDhTh7dZuKrcujffZotlVGdNAzjUnULdUeuU8Spov6FZWDU3o+6JO
JMKwTvIclJQieILxi+3VCMGNfv7LhjA6uDCrdrERSF3Lj0e1u4JZVel5J/XiGMVn
V0pAfzw8lLji1ihLVKh/mT8FDKE/I0CiKK1n5AIHIDNN9HD2itOvaNO1UkrQ1o3q
Rlg5OsIluZWJrZIE3v86KdfirCSCPuBwh9oBYjWRHTV0GBjoc1AeJUh+MhVTdcjS
7wapN7HpQjIck2JgryBFPagmMmmzsOmTRQ+bmSXGyZmc6nlRu0rv0K6j7fa8Axea
IOHAko5oYmXRIymgakGhfM8OENjp+ObWY0vLqc/MnwIZMZ5yrSs82z4vNEYqUPJI
jC9TBp9q18rHmHpaiW5faWoKsXzW7jx88eEkhnIOcYa+3kQRfQPBstHIgjotksVZ
2l1hKKpP6WpVtKBuR5ROpfWKtxwGJqsCWRrNtPJY/k98VmCjiUGKcJOMHEsSRysz
mNqpizBNm2blNlOBR4eTERT58kjDICW+yBKoJm7ZQTJm8OHktnuz81Tm31HLYCu8
PBTvLDf8qTXIFk+4ORnVxZBHKr+jO8QgvwPEmMohd35MNBHHzVN0asVSyrx6rLc6
fc+/7wH+gdEL6SPmqFAgT4pEBzyhOqZyC7rcH10W4RoNWYw9W8Bdi3F7o0vqA5h4
N9CX/IJp8SNcwBKES2A8/pRGkuehrf/mAa3b8C0HN+aAnVv+nQXcjc+LjRENXNaC
vrhEEgrSA+0A5RMGfQRASEZoi3UvdjNl6mhbljPHkiFqI8UIaeto5WHloyRwRtRQ
R1hVRarWvXmRp7fclAyN551eTkNl09rPqPgo9IXStc/ys/uz0U9ROT2hqkgT31YY
k3EP2oZMQyhq5umjjAuM+WOAICNPOcmnpfs9IovZNJVHERjZT0fzOmVC1ZdkNj7h
3P4ihyNws+c9ru9wCaSuV/kbZPI8i2zYJwN1HKKo5v5fKNsZhtrCqfBpq9VEQ7hR
eIm2W47LdTsqD0FsPesJmgcToDsHLtx9HgIoXRv9N+vOZhoLOoGN5KcUi/p8Sczw
Gt5ATfgfWAyNiqioUFUx+ySPbc40qdCo8QiTB7HyiOOchWqp539Lp5cK4dy/na2y
tCBXNfrresBTZeQE3e95PSouKpclXTgY1ZVB70gpekNtqdF74lAsWI7iENDo8jFo
PX8cCJ0CO9MoNTIaY0Kyf/SFYSdcXXbVpaBdJiGaw+5xQSBIlTMK1msqZIn0meWr
4JyoFLPtazHDzmgFJQyax6PLHBhxyAXoi4wtKZpKoUjTHyqZftvjwfkQodfkVvtI
cVm2d0w+Meiugxxtj3zEyYLJNqTxtruD07wFpfpfrxTiHlr2zWkeiO/hfs7lW/6O
eejbQ1em7+EB/gkY/Cyl21uxhB0rlwCwNetzstZODlTS1HZQvVXqc1tbsMOhRgO/
4yYxX4cuQInTucnYFFlB1rM4Jam1RAAVR8P9qbHSSi5WDPdqRnrjT+X+ah8H8V2R
uJKXSeJ58s42qFm7e3Ou/7wDAc+aXFdvdTWT5jLDEW3en6hJ1UPyyuzV8ileAlvu
0mQYrvN5A0eFq7wKf6+qvGN+yF7SXP6I66BZWeiA0LjkGJ0EIZFiPbrAJc+Kruet
KBdmagwfDBSgWi5Y9w5NiuJmBiLRiYIfvjXVpTxXEK5BpddNGJzbEywCgU+DvY3Z
a3oRVlk3mUrsKLIFy34UD/h45VyEJgxpL/110NCsnQvgCYufI14PhcKztdbPO2G+
OSLkRH4oDdAZLsyofbdOKIxjwQglFprhxoD69z0OYyc6FrixEwmw9qiQxJmbl4zq
6FMXtFDMbKAxI0J/ISAht4WhfdsjlHnSwiggZVOgdWzw3dXBWE3YQ0ReBhO9c18H
ApfzE9QP/kLkCuOWrkLaTC0qAjiz+2sAcJYFggA2SjP4cYkgk8yZCpAu/lIsi1G3
56t74H33h493/QnmNqZ6hm2W377lEfoadDbLTlW0RPfzsa/IQeQdzfz4V5Eu0fQ9
6SRCVP5FrERsdg/puIdcLFAw17gwiCEfbgBZ3gYz2ya6mDJ56FJXrmvd2TSv2Jwy
xZnWE38MWjbrWt5IylOo4RmFankM9C8rLFE1ZxIdM+IJ7jWHdHj5FIpEzuRD6l7y
dnc3ulVPKfU82Wg5aFeW/v6RAYQBMjZiedbM1P7iNiTQ739vV8U555YpUNEs80Ie
/yYGz7ydLkecTeXgGaOSMrOPaJxzCJccOzUHqV8C7JMVk1Wzzq0f4orK1svKtx+k
EtYgwte8QWAfO8uanC5iRyTpEGy1ygZi2gs1JzNbeMnaw2DU6Zau/hqlpneqsNIQ
6/4M/SzTh9Hv4kK/UZdL0BPQb/jn8ikCKycRFdrhkUWKYqge8Qa/oD0LDjdDBwXV
Hys0381fkTEOEOUUFn/ee0UfzcMKPU70mrKFovKg2TBvRovqT7SrwYqPIUon2zeE
A90m1BdVKlCA6YUuZEdQKUIoOk8AdkRAOv8Rzlh6ENXSctxEZTlbhm4d7P031hdd
WOWk78nhzAsCshdtz9asP/ByCrLfn2XbAVH+RFKSYRrOMkVX8voNTDmIHi/snRF5
pMMKHbqyKe6P9FT+/tvCVezi82FFdu/esfypSvpaXzliKG1J051HWUuBEYAMAdlQ
xHDET1TY1iKU/v7FWDg/c2FEWMg5NMJ2gfs3pPlCSRfkN9mx2b8WbKLAZBz8SOWl
ajdaqJplekuI4dmEMfp993+gkBiZ7CtO3XsPCs3udL27TsKDQZDpE+Y+ugVttUK+
Bx7q+TsOyKYnKGnuJylTTGfIE2hcAkN5unoOjVDOj5Z0GoGl5xSyzFnfMGrElJqe
I5x5NR6Xj2TfssXZZhS5U9zV0zESKA7oZdSDn0hWTAn8FKR8SDUewWPElIzHapUc
P2prmZx+TcLZ/A28VxntkWfnKP0E8jo/3EOZWDRqX/zL0+liN5zhb8YL4ynBp1xD
JRoTJszDoLiXlQw+bDl1rgZFfXlzrqj1GawZzkeUU+sVhR2nZrcVD4X9Za+JfKrH
QN9M92Qw2RgbstvF0QY4jZDNEHfDvgz+YCE8+YpRzfWSdIZyOgIHQUzQYTyFANkq
f4uv4vm8a070ZYNiq37QHyzoQMqXl5nB+HQc9YwdXVHQmQvSjpUCzCqUB0G3n0D9
dfm4HBc5gzpjUL+zvhhFA9UAax3R978Eu9vmJfK/wjH9jvbra0l8oDMm9dH5qiGN
Cpt2QVw6GL8MHQSH/o/I3QF1lg4o1h50zhLwAbJu8u3sVmREI/suquY/nUHojuMb
n0M1xD+pW89t2ZW0lxdFkRSM/uUWaY2+FNZ3UReIaRWf9X3A3KyWiWH0KT1tQsU1
TcjMQMRA5/EmmRI7pj4HMOmCgYIjQFc+aTPdZAJK76q5s7gW3U0Tq1AoJOoTVs+O
5bPrCL1YZ4XFYd1FNWvtSsPVwEJf43ZmM6t+X3zFNKpgsly3TfpsXrJnyUSH6qZb
+xR764Aqv2HUqaaYrmnmqXaueFQD5+nkGW26JW9xFLk7DOGBQFjS+ta0XZNQdiKv
dRu0LfMt9Rzj2sc+SFofQtfWiNcBV1rGJ1+UPeoaYLRMwTdVUsSVBkrSDAaRbafH
qGpCRTausuIve997bsV8iIYirciryoOHx609q5iHm/Ntkin8FL6eVr34UAsYod9T
8wfhXzJGGd8Mh9FZg+KMKqWuTd2MGc9sYAPsRV8YLZdmIOOp0c/5fLU99rULYYXs
wsVD8/TS6JMhTxxvCi72ZB81gwv7BLZIGIuAnXfxZE16p26m34GzAIPb8pfVa44k
ebgJmCR2mwvU7ghGfiDGQWpmbuiUn5cRBMziUXA2Pk4iAfv+kuHW9pcqA5mkd8oG
GEps/N8oPCfEYtGQO4v1qzTM0bri2itleXarPJHiFRXy/ovAENyu5X6DBdknfeBo
BQNmALQ4s8lwgpF9f7bVOdSPChyXZB6TWQx/B4VPJ5yygDZHzEaYjLu3rKuqP7ir
x6BGQ7cfpQ7t/q6bnzOmRNAGgDL5L2pCGOWY+Qw96m4QbXsYP5HTvqsI9QFh0BLx
G1+Ai6Ni8y3Zb+GhuTlkn8Dv0D0msT8tU8ER0F0McpP6aOBFCHRgdTNX2hpyE4pX
JJGO9WQbDPAxEtQIZeuJ1eYhxrUZ2+7P1gApAxq+28WMTfkuVYzq9Iqfsjcy/A9S
yDzgmzZ/pEn/YMwTP37tTpvnBdJXHA6EWp5vV5yXrYTfLBKs4inyC5EE2/HKuwPH
OMEdBretdCxYQFn0HcvE4NAtUP3ZpP4sto0Cv1vq3dBsmAhBmQg1xtf7hIZR8+VR
lq51zTYws7fyAZaLjRNu9im78Ev5wK6l7NSC5BjIj3REM7edoty+W87UkqT8G7pM
goTYakpnn7O5mR90HFMP5R/p36p5XenbYWHXKaGyweY7ocm7rJ8o5MPoUkxXCern
9cu1cH0EcGaXLh0rb4eT/3P/BPU03ONRk8+OqHbDJkbLPQI/T/RebhYVvH6dkeKD
iVJ0K83R7CwZJc+Ml1j1rvr8KMv4iARxGbeoBEqZ/tTIO50h7Ttyrz8RHOQuF58C
2jZSoDU3tgTGXZI+5xPmmSJID/v7ABfLVq6sgsa6y8P895EemtjySCw8dgXwRx2h
OJ5XylDIfEVy3c+9uPPMZBT8Xmsw+I//nbOi9tigyxQdgQl55ZP9TpJlKNw2sf0q
7wZ6LB5axU3Vb5zvNk0u5EmPdM4mN+ENglimzI/sbgP+WA4DjOgv9exuqfYhRj0p
KFnUXKZ8CcmoOqC9XyTNNSj24D6B2xIdmIr2Azzry19pw5G7vydRqXFrmDSDRyg/
mPEd5fDWIvcSgqUBdOC65KEH9fy+4RsLYO9BO+BCPWq6tJL4nthDpL6S7g+SHwpG
uYGuFhwWSwF68d/4/47vjMGEuU+p3cjgr1pR8djfhAVK88bNPKQ1m09jQYXya7k7
WVACzTVlQZ+yu2q1MP/hMVCg6xUZSy+kfJBZimgQMb+fSE1BC5zAEj8WJnLWSB8n
8MVXOB+vBfuz+yxZyWWQTz8+VEnZuf2qXjYEpsXDLANVIpK7WVxTgqyuFGYKMCpE
UcxnUAVa0KPJl2gD8uCxkDFGiYUy9oX6EYld1KgWqskQ5PU8sl3VQqdg0S4MwRqv
brDUg//jy5qqTNgemN5lt59BH9gv8PQ0DOlTZb+Fj9wWUdClsefxx9UBQsUoz6Cw
J2Hpom9GASuCud3Ju6/0Czz/ueWbf2Dd5FZoRwtFqAn2lI43r+oMoAFsIwVxijil
/+SVSm5ZSv759MnGidQfmzTf4ImVPxTcXhnessa3xOPIXng93OKA/xwpr+hNO3Yp
9AgUWfKm9ZM6jShe+SMX0QiKD+RXrs4TxCs13NL6pVUHIaLTvWCrztwpESsO74NL
hv3lHxA7abBxGJn3pWfDPsLWDq7mZfCgc6EKfDjiU14mso5rgCA04QCGz96GTshg
NIiTaYdC+mfC5pB5JG1C7kE7HDzx/SiMWw8jE1K8SaCsuA+HXlsxEGsQVDcjxiam
COWhlPrKvlXU3ybq/yEj8ZQ0ZunichxmhjQLsQpKdmiQgxVLDsNlthztTlnWFXip
vpGZj5zCYUtPlwy7CHDYAYCCoXAVSx1oYVDkFiWMopYVbNFT+CwHW7iqLHyUYusB
Cyc3YY0kO7ztZK3yAnqcsG9FMsSD2TNx9jxP1gPU7+gN8egWdiuLIgQlf596olLI
jBFxGLhKfE5GNEuSMJKxq60aZ+xp5Q5E297wqCg3JnPRV/arQTzRaJno9smHqE8x
NOHCZLi4r0fPMbhZzHini8nLc2ncvjHmGsEHWK1wUavllj7wRaCfJD1rgCdlyCPe
YiqbC81L93Q7VbtyUcjsqOPUsIl7qCj6afJQhpz3dXlOeCRm3dRAEiE8V51CAj9H
oIGYsfLuZoDx4GHGHqhLYh1rOBVRfWh0v1et1Vs1FKA3rWDSwrCcKmepdsGUrHGY
xPACQlEJzHkppmqJTWpquut3hYPgUtrxEX1J6qJA/6Si688W0Rvugi8ZPbvHGpP4
/oRYJ9J9SVMtf/U9xi1n3b4raScLJLyOfJhxjrMeXuMUJZhtBKEhXe04jRrBwxoa
PxjbSSwZQCLU+hblXnYrWiFrDMrvMmxVHqVJG02GOhMRGkReKLLQxiiPxL7HcEYA
jPW9FalZ1Gg23afu3p0Oxa8+6CumNDzq7sVE0kIWB3rhHsCwU2rLMEc3dQFf1tn8
3yR6ZqgbAC4CMGxTsVqF/3LcgjGIRCTFoIWLRGRAMcKzbDuoz1qXnnX1qlDkYe5n
dAWG5YKRUZHPKBDxpLfY/7FHeehdgbt+6K2eI+y2H8iRQaTWCViWb8sKKPQto6aT
bVRGQDrtyFma8tYGkm+VfFjMjiYx7LEUYSDgkrCxl6kdik6VbgcOy/sEM0a8jRdj
UPX69SOsA310gYCwcnU8rZngSHH3Th+eOly6O+o5TUgjqYf2SNN2c+xmV99NScS7
wZ7MDUwISf0VhTRvJklMOZSMU87jXmVTK9LhKjGWY62ye//l7aIai9q8A62lhdRB
41AAIKJxXk8GGxnhWeBnX45LM3NL6VeDNLbAjQeGhkCuzXA7cb17X+CdpYL1imse
0uEp5+HbKEsxPvysjFRkrliXbr6a2yVA/CRfCjyJLy+7jrte70oD+Tvj3SLQ7GIJ
PdeGFeWXsBtSs/RieyNAjJtivDokP2uXzUHd59gIV/1vPwPZRHFnvflKLwxLnxsL
LpOJcFL04XRJBGhUZUcLLxUE/CuzYfpQEsaVrGdyi0QRn1vciRl3bDfvsz58/EDw
XYwru1hemtJvMhNKAq6kOLDbXlFbofhbRl31nG3oLhJKP56miBTpLt303EiMRymv
QR98SnOr3gn2ckPjCRrOEtbVNH/M2GjSTEoCetm6RY++C+BVRGInY6jcr8jziSYo
5qYh3ECvf954goTI7MfCf+YNp6O6GlNc4Dgbt+EYWEqBnb1qKkfEWpozSkPn8C6N
oS/RW6LQArwmWvRYqvevMDKlq/g9CplkD/YqkJQkDUMuY0wRyBU/U8/zL4tIS9ip
uXIn0Uxg05w/N0sMVdm78B30ZhHjuleK0lXPb/QcrfiwjtouoytSZVN2qazCmkl+
EJfsTDxetDM9fEUo7ypAeN+8M3f/dYGSEfr0pTLtl1FLHgr+rxSoJsk61DAApWVD
9K7amrmf4mn2pdx6xta1bApSQJhVWMfzk4d0Io1/UZpfvlLSDxGUAb3DlkTZGAi3
bbN5aaN9p/pioPO3zoycTvBbn0aSRP17DbBSWyK1nYd5qvz2qaEfdNTtJJjv3h++
A9HNzLSHS+nZceQo2kGjmE5Ahn1oREmfCu8zi8mb2ozECfq0RGsxoRP6OOgdeEzq
qd+GBEnG0ld2xKjuLcwPqVddIsI1oMqahtWZ0pfna86aE1MncCDZUvz+IhGFsaJd
zwczrV9TqXAG3I3MB6BD8y+ZK2Z880NfEZ6L2+iN0SHsVtRrE8pOyMmhSrOaT2J3
7I1vUzaKgN1WlhukWGwZxYWacdPj1p2BNvoLQAHF3MQbO2MBYcQZeqm6J4CWqZX8
ToTCF304/KHp2qazWW7wKXZHqhF9afAt2Z5//hZE9/YrnOIA9S6j5GAG1WQ/GnWF
BL+pYgfblRoTEUelHnHqFMwiIB0lbb+qHzQqUXrQjb2zZX739STXEapQsDP6HH9W
dRlM1hyArAbU+ggXvcN0GKhuhdtDShzyy/pN2g6kwHA2iBLMZlQGfPtwH/3pKGBE
sUDspQvC/b5tHJ+8FKSJbrri9vrMDrVX5i9x1sbjDd+If6uEivNN2bumDohjObuq
e1MDiTrBDl2zdWdXfZcLRoheYpGqiSjlBVPUdZ+kKR/Kvfrt9TxFeJkjA0+aWpcD
WxYf+8tgPWmvcdPDtHDJMhv8XzIZ6plXHeMOOrOF+2CsvdLAls9hRzVZshVpPoUW
IinVXzGme4Ko//0GSO+99bH/aKi+ePHjEA+PVxduU5nsTjbnm0r6h2FmaLraTldG
iQOWl/fwtOUmrg9R6g5z/ymt3ujl8/lbGxI1jd1jXV27SgBmlhKAGFaPxQbmIBlz
oZeWG534kk6uP/yQSk8GrtQn8FE2RxDAHVJFBkyb8rR7eZlpPlT8DVsg5IyvC8Dy
EUM3RpdUuZIF3U0VMD5N4vvfVrAyNKgDql2zwxerRydu8zGknQvIuRXcMZqmDBm5
VyMhGQJ2bCjUaX0TIjbUh90s5pZrfQdT6loDxhZhdpEf+NTPpHTueJwBuw6NUAvE
Y6gg2XCIeTO8gR7ICgT5Ym4Mh1qCKv0f3wPyBo3KiWFJS9N19mz0WrX9FYKMoXUA
Qk+3+8FGheukNLrFYtqrLViojK418I325m+LvH2MXk6OroafSU+tUspdv7puWCYj
Bce7bq24LO06X00VVbc8qwXPHbNs9FIZVBeyxjkVFQhXZZkMxG7pGAIORHnrO0JK
eopG3HIzMCR+FzlgSTfn4gQoArJ7BZ/e9siJMr/uVi81c9/GpcXm1KHkuGeF5000
9WhN6I7jqJW+ebLQ4av/VKkW8F4RB5hFH7WdqZiyozaaBtq686KP8FbIhNYfVKbQ
9PWAiBPDGPX9VBxwPCehkC7FQqI3ZfuDBJY37VtHP9sXFZNhfZF2WBg9O3GPzlbC
nAXFesYa2kl1sOv36vtlgZXzm2ZZl1Eat7uo9ifOweBUxtvIQzB5GwxF2O5NsHjm
2kEsAJSBMnlGvZiO8SmLEQfNRCgjIVxEVRnu7ro91L7jmgNjqlO+qSiXKTXy0Qkw
j9y8mre+A7X7XnXCGEuGyjEAUJdIcS2ctXtIsTURwrmYNKo6sNMjmuZjT2uC8TA5
fo3yOeBYLwBwYYJXy54tdLDJ2MJ6j4W0MzP9CXWNjxpAfBuiThbVJsXcy+yQYWQ3
xNnSoe3pr8+/dnJKD431xiYnEo00nl4WiBHkhnVLpLAd58VwMRvRJhm4OnwqPFaZ
M0M8voG0+dgoS3/oMLeMYDSd1TYWt+2j//CAoN+lr7NQ4ptm4hD55cOUfl4OSVx9
B1sw483llZ4LMVXBdJOxo/8PcEgX+DYcRAmMhwVfup3VMrA1pALq3kB+CgdHbnn0
Rj3fHsIpGV5a7Fq85pNSh6diNW1322MPAu/mzA4sMflXEs0E6ncMXSZSX3/wo8NG
r09hU1TNKtM7JbKif7QnbdSN+UXu3nGlsuIUA3E+A7WyE3ToM7j3C34ju7p/dL+b
GvBzbo8cxmrsPHQel8dDlHReXmW1xy7QLN2g8RqLt8o60gT2d6CejIhEoiTkPELI
wm7dvIZp07DoLMm6SrmkL0QKmzX83BqTk+ydD7uTjpLHQWFDbfmA8BQaybpv7C5r
EPEpjQ+5oZSjtj8DlrjX/H7CcbhLBraRlpT5YJ/EmxI9pJKrfRxZWthyOqURO9Af
yKGq6rRIuJabHaUqtxbWrAqajCPu3TpVTaa5f+GDHytvuBLrzHTuPRe2dam+AuDq
J//PobAx2lWd1Fss25zEUys/6+8qZeXu6Anzwz3BYExyQD8c8YAktQOrMrfeqRmG
czk0Cizexu/w6QnVRIZIrgm+9NTrxYUslK9dVQ7PtSWJPp3qkp3d7Gs1Ry/YGFf2
B6RRE3BW98wA5GFa+4dqMgKzijA4F8USw9YWLrgvwbQu2kyI5r/CG/zrgziERgHF
Q11QvHWbKeaWbdFE7acrd2+pis0wbw3Wfdg+qZPsFjeKmvJjgZ1Y9srgpR6rv/p3
KRFb4YLM2JomVCy43oCCz+OIXYil0Ol9UBWq1WjqznO8a2Y+46rg9akP3VMLQqcN
GY8itjIii7Kforez9bFESJ9KP71xsNlyzxUss/xU7s1CrGm8HsPX3QTAUH0Bp0Ab
NK88HWMXFQDnWZQiQbvt/Cg831tE4HbtkASSkHIEXc5Rgxf1HnAWh2QMiRdXUKaq
WchGn4gedcJmzHxtOQd247sYjoNZwkW0hwuSF5ihBx5f51rDEGT2IwtoQvTTRr26
P0dSMzpaxUVViujfOIIWO9OTB2xK51312yKBJg7T6wnKr9U4Sr9eBxTMRq1pXwnj
9riBVUyfs6pnV3vCQ7XiIN26WKmIa9oZGZJmk8AdfihcLsPHgJHrDs+sHxAxk9lP
Wv48n7wu/4PmYq5YfuwTGOFWdoD3NDd+pJyL0iKMLock+v8NMqr036upMr7roFsy
KHRwJG5SVvYLU6dlJAenGj6VTc/awU+KdYcMVFI8h+Ad0jAiiEWNrPHQJ1wkhswm
nVngiyHMXoKRwT2qNUVoTQQyDOPCrol0oiXFKlOCr7fu8b7/GY4QYdTSDc7eby69
s2RD25mLd2A/JAUU8QY1BNCcPpsZGM1Nvu7+DzA3JmzlXxqmQicghqYHPNRtXkf6
r0v2otprT7B/bfd/oz/GO1Cj+X71ysdgEQE4OxD2hkrRQHrjPtkYJybcV3lDbaw9
nFpR+Aduy5R73ZjFTv3cBD8+peymF+HeKy6AeRQjOX+g2PZS8M6QKMossh7CM649
oLaYBXKA5RcV+WrmBBiqrbI+0HP48//tUNFQWythtRSoQ/A3vMP7B8VsHsBP6Qmj
DpdoMgxBpULWLdtR2Y28YgysB8g7FudrdfAHhb9pn7i4KDek4n6XQUFeG9vH+jOT
RRFqbfB7LJFL6B5K8zeq3ZKqjCj2A94CLudmfYD0mq3FY2qE5ZNG7r0cXMsiQznd
Qxy20gftEk5nsateXGrl+ejQ1NwhMH9aDEv3kKroYjqN/0ZxxEXq1sD24ubNUzya
F51v/CmBrql8pk4pGNvtpA==
`protect END_PROTECTED
