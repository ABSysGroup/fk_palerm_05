`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lAy7/dN/bzh5pMHNFgMLGKnoa9ibTaofA/EpE5gMuJxkNyvBKf8sdd/xYxSa0wj2
Y0bsDBvJpM+X7aNpegQuM3CEgOedHrwRVTBfkIRJx7dAn2mS7U+r13p4mCaLEL71
G+sOiDd1ILDBFp+9PTT0PhUZJMF1SsvnjIjS6CSnJVs51ettHl08cYP5tebpidKV
mflvEEYoKHZF0ySb9dy+1Dk9YCHz7J9Bb48aG0JxI2CpLobwrSZM88HyPjqzDayC
rddoxBNVOXVOTpY0XnM1aiQ8TJv+mDUfzu6szZDx2ZLusER/2WSo1XxP1dC/FgwH
bIo24bE73DFt2WA6/HOW4Fs3LhuKGCIUGkCNvDGEgj511nL+IFCxJw5+zDC66DuB
Sbrnd96lRAHkz+2el45MDNYPl2z5QK6Bd3GJfwr9LteKHa214gY9pgz20RycTEqn
aMnLwrAqFaAzvNlDYuuSWPi+Jt0amS/IG6MuM5iPWlE2ZYOUnJN+7AaQRlrx0+xl
`protect END_PROTECTED
