`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5j2iEKn8kV0umA4JW0BZKxh8LdkfhZ1Gl+FEj/iVHbAei0TPuA0Ip/c8n8ZJheit
6JDVkORHb9eVqH95afId51MinnWsBFwYfWe6frKTng4ebduvy9ZPxKfihX0KWBHW
z/nyc1teqruXt9yRMLbRIwxXGBW1yJYdASvyTlsX25LD5dt0fEXygL7+zATgINCW
NHda9OBDLUCJZrd/w0fkn0sArn790Dp3lzUDayL6LW8Qzrl/eLJMimCwItCAdQrO
pH1oHMc9rg7BeyKhvmBW4Hi8j3ii816CpAIa4gSGI+duNBzeRsU60p863/26uAkA
aFn17m3G0NPDSU7ACv0ED3FLnZZ3gToHX0GFYUPexONmKk8YXiEfHLP5vWRM0UIP
rFS1PDo/VbTn+AaeCIN//Q==
`protect END_PROTECTED
