`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rgDSNEuhknlAtqhVdO2sjbPgHpDP1Rc0zbs8z+Y3GUQ/99u/rcKqFGVu/PYtBnBL
1Ive2CksYvkaeekodphublU2qlkHhVxnmrEF4M041Bz4MYh7P8Fw6NK2yU3iE7Zm
x/uMiT4gXQJPCKGENFdpIhJPPx59JutgJtUL0AmVkO4ndiHKiqqfpJCGygjDMrSQ
GLIeyCvyrSVdl2Wle9p2/LTz4fQpJVta5XD1AXuz+PDAdncJp37+iev1YfqCG9Et
42O/C7cn6IW/ImEL8X04Qx8vTrxX/+FG0N5y9qDo34WbOcBMkluE5YuSwqaSLgs6
qqHj7KQVTBiJ/6NkMclE/lDTGnwAnS8BhS12siMoUKGzgIQgG4gPpWr3VDCUVW1P
jYX5myu2K2k6I73rTSz2Cw==
`protect END_PROTECTED
