`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kmY3sRwfP3jwZsgGZVwNsfK3L9+usCMDFU0Pm868SlIibzHaxUFga/nzFYy4gIs3
CLCGmaaoL04jZuHfwQWAycRKS6t6TYSAuPO5RDFcCzO914aWuiRQ6/UYLzj30QI6
2CCzlod92EGuVFNGh1tgdf5+t6yT44viNoPGe3RmIUelh13n9P3867j1Wb6i8dRH
YgHoaVE1ffl7ICXVIpl6zv8AcS1VOZ/dNbq6SaW64kKmJGGOTwz7J/wobfdIPUx2
Q1rSNYL1JbgDPXFHxONrrAD7nyttXOzckSZdTuD7dSQgDtTTkp1X5cxwtkYvAtuP
siiMbag5SbUPJiMHZQcHSAelAg/+qzPb71MRif5IZq+2txhXHkszbaGoa/8atrYs
c9ywb//bG/xLGyboQ4HgxKe0CBqQ4Sy2v6wQgMt6kv4WrYD2T6VAXP0/8zzmcXHp
QmRVuz1eLt+t0QFYBG1y1XjagLIpCkX5mvQqOsSxGT0JnWW5ev1E7wZYj80zmXP2
XK46yiELXcD1oqAT9RLDT7i+2/NqgG/5WdJj04tD57af6tx/XEV5q6MHOEuSQm70
JEH58rnwkqGK7v1hvtpBaUCmANqtbFR1cYyhzZamEkjA7xfEYsbm6DDwk+Srn6u6
T0OJtixvUQVxONthT7g6JKrFIu02sfjM0vKrFpLzjHme6tDl9P5KOKQW/D/oHXL3
dBdCaKtIS7e0GHR8B+eJgb2YcGO0eRb9hisENee5vzmjt0z2DDExcDdJJyYoksxB
el8Xin5A1RV7xEaBlsl4iTnRCqsmAc2zMwZVExIs9AdJBSStbwm5Ba0b5mssls1+
OA6JPwkfn8GrT/9D4yVUzpgP7AaRT8qY7V4K1jH+L8ztmm+OG2wsEHIRE9diTTbm
KLMVNMSupDGVwyQXbgngRcJ4Ecja4hZk6lzWuh9pUNVqhIVBXGGQvo0G4hMCGcQq
zkuPjoLzybKV0juZGqmzglwJO63RZgDH4Y9hXFH1Vhil9bDe0mb26CPvWtO/afoX
WIPWEBOtnyLKMv0KIvM4FZMaSN05SWrSfVuJ3WJmU5nxUc9KAz3LDxrHB/Pw+Pkw
Qmh44nXClUkI/ZeiRCuWF6pJgnSpy1RPjM20e4yiYrmddWjrM4yLhxPuRxfpBrVw
2nrDgKzZO9bhGEwjhweZG17G7kL4g517zdtaXUC1vCpFYCDWf/yPVN9coHvajgmZ
MiNqvkmbV0bfnz8DdOaolqzKTUJpI961ttgkh4nC/LjS56nf9neSJJTCvjUkwl1e
jQaDL8dGE5979YjTboeCDdidI0vcd8/TCU0rvpZHG8rkqFSyiSWMvoUO0SRLp8iL
IuaR/c2RHLE0LG1lEkUNCeIhKYrC9ZwING2NAtx4tgIsCYlXOtncuaSKeDO7ELZO
KszcJCIaa4nNt/zruJIYEA23v1EBpMBa4bUVH80jSMx1zqATDelwvgRgXn8f4lrd
XZpUIZ+BpDiS7I6/BiJdG9DVAs0hLdoiytbDiSC6zIJ4YZUIwZ+Jognp3kc7dG+d
zoF1R5O4HYrwEhUQt6N3e5lfvfJSN7flNmXrkoLsWxyLCZnJPsQA8HbuCMT+D3E2
wqEu8MEMtRgYObk/wGGzXpV9XSz1dXJFj3pGEObeA6g6IaQl6FF/OjuvZlFrqw6U
9hMOohbuZCS8YcVzUSbm9dvUrB+K1oytTqNN+S13ViYw4oz/RETcupUAdsSNTEn5
Na/XOhTnxq9VwVmoRC6FW1m6JDmhhXabHVCK5eSHjT/Hu35Md+BfA3TrJW9ES5Tg
IplKiu/s3WkknhOxW0Xk0lsekw19jxrkn/KQH4HsL+t+G/RxJSFIuYwUil6X0sKq
G9U1IcBATV4KWE6Fe7i62WCF5A/1L770iRn6cxROCRXeGLR7eFGPKzloUdQf2tFP
j/j60WXNzmyApH1KWQ/AfQC3g/46k0lDc8txx3A4lUtSsUTLX8SMZwLSRlfWq7w/
s6b6FxYgCeIEcN4Dzao69kM4dZ3CGGu2IKXwh4w6z+8LEVuAme4qtaxSY8mhLAwe
RUK8RGMvm7V1GRmF/DZ8H1rIFydoo3YW9gFjH14n+K72l5U5OZU424nWWpFH/yDn
9QgDZ0fJqBS3hooTwSRRCvUG0y4u1ANTpTvLeJ3+OA2MxNo9gmxdmzlO9Mnplcd2
e+n6OL+nnnydgZYGEdmCrN+DagwEM1raSYEFlQqvG1WiY8OOjbQD+ZPtqz9/8GtW
DN1kD/XOaw8xvtMgeqGiEQ0RGykgL1std21cLQznY+2HARHj8zVJ3utR4UICXnQu
zMa00ewv2SuWcY6BUMHvySKRP3M1kZALKG0vh7sWwmbdxLr+ee7POSxLyIonEPcr
jsCBjCyEF0acw7ZXJLcngVKJM7Zfl9qOnJXhUAQTXB8Zzs/S2m0487pgcojimial
TxCVjI3hD+U80MZC0pRcRkTXTalosRvhqUyf1PbCO5ErHbhp2KQ33/gVTaLaLfyk
9QPAIUN4g9olf0tJozSmkGQriOVICsu+joYLmBozKQCVGXKS0EESdfHoisRdMphF
F3qhlWlYWkNXyeve6QL3cmw4IxIPkAKY+NADlgzRwz4IDvdknyuhQ4k5KkSP2f7W
4HLHxi1YIFWUqnkx65+7bx3+Sm4vx0Dntt30kW3fNl0FRC1bohg5vzwglx2ZkQga
pmMIRjjQf+DOkOPoY2AhoutSXXZmFP7lDEDFQivG9nQmceHkZuEUgM8lDdz0SkS0
+Hjx1tX2xd8vHex3yfEgMaY1kH/zDUu9zwhEEoAdD+Yp5Cb/q2Qf2Mz4fpKvui/z
T494wVNbQrhF7/76M4/irK8VqlEdDJ96IFVDfYm6AfGx9Gg2yAtvWGjdiptcNlZ+
zx5bI+31Dd6Eo7WDtwwT5TQ6RqtRWqv7lV+9Flc+K0rWnzLuiQXf9EltX+wjaBwd
Fjcb6InOJ/mLZnm7wWUmBnvjBvGoa87Poo9SqhE9HePiZOn3zlf1IPY7EVPHDjuG
2yIddyKD2fJCeSz3uc/665jDryR8V4ZzfQD4DgyiLvJWDGYuvCHHuOiiSTlpGSrA
CfiNLx48X26Kq8M5dIK3kXLtkSM/gk9YXLBqHXgvMzJ0qSxfA9P+ZVG4FmC+ieRN
gppjjGjTpTPSa84+y26JI5vLJD21u5ZdwpQPo8A6SgN71n+AX7xNxrtM8pXFZrll
142swyqVypZkLs/ok8VdEjDFz6EC8hJRNJmcQMd7XOE=
`protect END_PROTECTED
