`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ms1Z9BmUH64f0gwCL5GYqxbb/xtSXmXrWhFOCFIxS0a4klbs38ZAh3qP90VoAnRx
S/fJ5sBYeS+vaq6HT8gBqZ9Pf16ce/XEQGyt5jUKBFWvKiW+vVIePE9XFFjxxXh1
bwGgrPg/ufmBDdYvlIbXN1xFfdmGH13jX7+7IlJKgzkfVOhvAABKCffqYp4KsNbP
1kDtxU9Xuwhh++exCqXzxZLCQV/3julwI0pX4jVw79vtdxx+T6+Q5jlPa4ysRuZK
H3W4kqUMh04oDYDc5FOaBhfVEp+feWAAderUNrz/FVn+0NAE5P0XTJ4nJE2oHhqD
ccaOocW4UEdaE6OzHUmHyla5AAxPFEYNov2p7VZAfCsnHfpwMyZdxOuM+AJT8aQ4
r8va42HJ/cTCcXS/+Ibrx/wesjQUph+CIBQTgyvJE1+Ea95Ye2t+If38FVVTvFJo
/0mtnS7nLjJeiHILGbm3u7wWvrX20XJgTdXKNYkeYFeMMkMngTFmJIEBOLLPNlIx
FlwgCJ6haw8WTKtD0WmCijd+13PCgUUdFq+NSAAukWh6KNRSZPCb0PmerWi2jdf/
WtIFnKSeAOT1gkSpUPvpoXDEey3Amah12n8q4CDxDN9x41WZwvGDhVbgyN4PHUDi
htIDFd6LEMieqsioJrJBhCR6G9Y7fudJ3HpWB2AgF3M004l+jKwQ4KfsYH1SHO0Y
bFUKq7UhyARz7wF+Cn9Bg2Nkg506ta95tT/ERu38SBAqjTRrKZkI3fFTpS6FmZfc
kNMxirW20I87BJtGLxllZmsSg6rQOXR0ySc+DmFbVIveIKTk8Mn6FVBPcvqNqaGU
C9XF7ER8fPORd7Tx9hSxiSljNXkiMh00XOwRMbDPg8S/iamJv191gIBf1xBAEG/e
6bPdt3AK2D9SFncwQ59jMVqM3cLiH87p/iT+18THIiIvk0A6pGoWWn+ixRGo/YSi
CFvUq5JNESCdufJDz1C8bJ8XK8VqTNh9lz0jL0+ZN3DxeQGBjUw0tUzraliJHz8C
rzPOURgNtnoB5v1691FEtPwWlkDe3hL9g7vO5WjgaXG5Gdjz+5p+/GZ3hMOqlZxP
zXtjixwPAwsvUqi2gJtaEz3WqiM9hw3DRHTOwG1oAF65ZNFZDCLCKEovNqUZC0l2
iKoUMb1nXac3G9lrEZUTFl/hLyDBnZFsh5bTWubsUCctJiQ6gkKC+6udbqqIUmlD
DZ/VmZJAS7Ttfj300mNRNuXTZWn4rGIHQt980auySGUQzFOyrcn4h1LeqGIcN0rV
/i4pgdIdsdt5VhN0KFz52yuqvH+y36E90klJ6W647NXpKrNVsBBG2M/uz29P00KS
0SsbepdiEA8bO7yA2stgMnGy9AB3TGrDFqwAO56m/mz6LUk/05ktigEeSEeQ3VRR
FAEPgK4eMMjeCLhysc9QNiAygkDEK/V9HKy58woRz4yDZFx5igMhY7pFaEbsttTf
nQ4XFfubXmxfErRgnZOBLC5zsJBEIl66G/9XEwFp5AW8Mwb5HQUfDEI5zVnvDYu5
TBTeW65N/PCSvBJ7g2Y1Lzn7o4laEDXjtYnSfmpWZ/l1dEtbG+CTj6GGJrzFYTXL
e4ERLWNOYfOGOZSQLKZIadwVfd5um/lJZC6P7ey9nRN3e4jlkNz8RCnkpbxzxK9a
ijBJPgn6OLq2HTb1fJVBfC0B9hOaKHJgacA/wlIqMG7mmG2kqEs3mnKRgE63H5yB
g2QEN6EPOadIdNqszwnNd7G9nQx8JIETAZtdMp+sFvERVmKDUbGK+t62NNm1Tjr7
1LTZHpq7E9cgkEMFM/G/9HFYvpc796jCW1FY0mO6ZQ1tImgB3YAm5PE7ZKO5fYet
sJ66uLnx3SiwrIo+Dx0IWgQlw41eKm2Bar8uwUedkkxHfUPs8jGAKB8rfkp58rp7
np5jZ4DBDtAymtipNad7KDmcKyHlH6/xwuNjU/3HFX06uNSpyLkgI6HcPPen/48z
9f0uGGYwEkvyJnMqlnP1Hxe6qeVlUb/DJGkibsT3crK3J6O2rdKXTR7xehoHLS7o
n4LrOhTh5tVmxFFw+giNWpUZqr2HNFAeu4fWfDKnMrFre425aAwsHySgWaGnG2iE
yARVxCYpTZGMYnkJy/f+niVL22l7AbZew6CpsMG7ALVcl7lq/WGaObkhsf8faCM3
`protect END_PROTECTED
