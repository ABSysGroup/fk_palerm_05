`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EomjKeBmgcXLXq853sjaOiXhs5dy4QaLh8fhz0IwuHPHYCrt3R0Mg0G8sYCwtCyO
IPUsWG5GsPGR6E9E21uTM2CvgHOhWTCP7MdXNOTMeVli7yT+PTotn6qZDwJYQbVF
S/TEfL9ongB7l0c1Wwx3FYfZJ0S/GxprBpxOcx9dKb202W93XANrTsDtgzgSt0J/
1bso9RhmMf+4b6n/fdRCc/wLxqCimg29BaAMHMaErjzf4ARt30vqqHiODEC4yu7F
UXp6FdJTUdpoyYoYrlM43Ta0hIp0MEafadvNmJa4708=
`protect END_PROTECTED
