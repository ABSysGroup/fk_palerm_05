`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rW9cuY0Qfwd550hnG/OKBDIBW7i3WHIgAtA6NQRclP4kYuWSX2n+DAGq5PC+mZAN
GeFm0sHeAPnDgQLUkowqtg9XHmkWFxUZQ63fDoE+UezM20Erxn6MHnt0gP0zd//C
FgrOk2ksPxDig1XIPiNrutXtx9Hu1tJuc56nCbm47sGu+2h9m/9FpvPWUHdviAEp
V514euLoCFLuJtCBIhIHSTTNe3PgDVCCa1t0pY54+eP4eLVZY8LSCPGud+cFSYbP
yBYrjmgLyhtEzpweKgS1Zp3ATMjmAgha2YwhfMyIv4VktXH2t7rWQ84vZDABxk9h
zw7fPYpZdE5N1cA8sqRQKqyWPUtEGP2lxz9UJb2KiT52ABRgzYJ1JW1NPB5s6Mst
`protect END_PROTECTED
