`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CrfgO3mBvCIT2ICqBpjsuUK3cv/VgnuLaFJp3R4B/QeeTRIIiWEd55z4tf1U2UMw
y75g+Mzbzb5y2Te2e6A3wx9plQ0nkCuuBMPp0JbVwQgd4SjiToXu1eISkq0SAhNP
Akgfcs+WsYTDFACULkhL2wWIAcxaFBrfxpaW+5HLKgyWhCmqfFo+K0i32AL/aTQg
s0VkTODB+nRQuKMf5qET7FotaE9RMtCGJAGfPxTZ3GpmVsztatoeBftFdT4rjRuO
/EWZB/X/x/QJBE+6C6yzEbF7nFOQpHzR/PL8v7TXPokw4h7kF8fUhPiFX522ymvn
4B2Rrn6ZzoygUpqmMf+pSKuSgSEswwZdd7VJHDNMhk3+XtPexItH9PY9HaeuUFza
uuViOD7dLSiLpFrPAmJ6OZ+iqWs809SEkdeGDtAjWuwnIVGsq1Sgf3lLHTEk1tvr
tNATic+PXwwQ1uayr1lF21YXQWsJnXVFek1naGIhR68BLjw7kvu1nDUbkbvb7kV3
+gmI12zVzeH9uk/qRoUKxLtSzoU04emV0VY3x1RXcrnA5/ekh9Defg4Dydrk2+ZR
5KkeyBrARuritor5r3BzsmWzOx9xXZpz+V2Q9Slhos+hbGAjxGU/607hHSY4EubS
k4qQuqdGdR9pmqC0Vjvge8HWMDTBOYq2mueYrEYn/PaujECxyAcRPblWVzBpYGP2
Wm57HM+0h893Wp57/iRkBmR5lm8lXwIXpSf/ZybM+wAehCBmaIqBXMsrSABs5Som
KxgfosH4WWauHZnOeKiycItqBo3Oh6uczyWcaAMieDBTikb4bRRDQR2sOoNJ0wnh
LfqCldAEgxuXCohYJoonclSNuUHjRFPXXY8LzxhJ3RsXNn5rugicyXWg7OG3UNEe
KdMTFClfuIxpp9QlNNwspnSuCnHzxSjNtN7iTbwkO42IMa8M3HGH2SONWV1hnIwi
`protect END_PROTECTED
