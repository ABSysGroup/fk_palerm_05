`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rnyq6J5MrRDX7XtoehsuhEK15n8ktlQlIdkQ8YDuUf71rkTyEwU07QaMvHY0IOK4
GywNY8mXsM9c6XPu3D5pxM2icxJFTMSVCAGSaQSRrOA+zN4uNAU5LpTuvvSn01sw
zT/+jOTa8o4iAG63k+9DAK66BSAgnspWYSFNoyF4K/7fpVw9HHg7wof6mrlGLQKp
e4aTBAueNOcv0mZXwGufIbjuQqJIP0dHIjLWTjvWKLe5jP7DWg4PCPR8y/MKzr9t
lUJYEAblXbf9QJRwOLQag1Br2oVdixmEiSrPCA6oWJRmTPftgGJuf62KwilKPpxY
wRI7xBzBW66X3CNd43UrjQoYEFW4GVk5G2sLntMfj6FLAaYq6s4UfMrvLAN1rHFZ
iAjzkqRTrxi/gsJ4E734ng==
`protect END_PROTECTED
