`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tg9BR6T36KrCdJ5IP3t8mbI0bqDmN5HjisLMRLI+/yI6akL4UQVowrL9HzVj7qsN
nHyr54sJ3pepyLuouYp0sZLcOGriQlwrZ6yHfcJjlcD5gdAQ7rwm91Zl1navTkII
CHAqwyDxMpuKIxx3bLFBVfVea1LQ6sdSkxqmgjPdj6J8K4ZE4mdza5O+CoccYZiu
I+5wKFb+1S1ohcgqxRYBC1urAHlPGy0g3ErdBPiUah48mZR5s8rSIU7H3eUdLDwT
e/SDGMKzHIam16beCncwv5lNT85BLXp1RuPjQ/4eTVYrDlGiLHe9XUpL1OVX9yXF
kZSE2F58NqV44G9iSU+A2I3x6vY1NnlQWIUKrIFh8z2Qm+/JPClJyXOwKQRTeLI7
Es1XKKnKLPIrPTGLdESp94AGjmrbYsdwAw1DcDqjVI6yP2un4Ak9g4Fy9doHpv7E
c5Uxg5L93SfVdYnWCTkhkhffAOjxxzC4CVLi85ZUtvOmk7NQtV1OK9ogyY5//kQ3
4Ed8FTMCRH1G0Ao7s4RGRS4qW/KZHdXtcemyLZwsvKcrKsLy7v19KI91mUW8/Xru
IQGVScE2NXWNViZQE0YLrKFAfsVQUd+lcIIFTtqcY3NwI/Hc65ykQZcWy+ugEr1k
lljnt6dkWxN8EzTaSzDiuq+1TecEt6gDbpQ51ZdSUxMXKxORdriDX7RlhU5AcjNi
zra8DCL1LEluVweYgnMRPtOOIFaO2CImlGxRdGH41GzJ1V+MQrpEznv0/8OKUdD7
s4GHBW4FV1e5/PZYb9HFgw==
`protect END_PROTECTED
