`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rjRu0OVtGB65lbS+X2L0bnKUT/3OiSv0DEWHDuNnW+ennijOR2Jupmaw+xMq8M4h
D0Ld/ohaKdYqGuaF9/Oy4dvVdEKim5PMC1tZ/bZWAtGjcAzIpWXRN/NfTLrfAY1F
bWTgzNZjwRkxtUqD3pfglKzrqGaAr10wtO1LB+L6a8+ggtwIOATZnnBKezRvE8ZT
ADbMUwdhT4uLJPl0K3IOWErztz1O9JNGk5wE05ZIF4THc16lnkOhbOXf5rsj/QW7
e2mEox0acFtdRkz2BtquDesjXQWdxWF4aP2liYOwU9b0x3NdciD+X6Knp66wGufy
CJ5NnLv7n2k8d9e5oQZR8ndaOAquzaoC6DGkK49yfYeQWtLqKxMyPMYxDtggITm/
Pc2Gg2q5pxycRddwZscQGy8rCQpuR/k6AOAhp30R5oQcaV0GGXqWxs7YtZqKnLPj
1AiOpWYMSB2Gj44rVgMBHmsjYj+UwIOs+Pdal80G8pqrNPIiRhoPegxZB67Wvvd2
tyUq5936tstaT81jfTlcOgqKp1FsE8lTrOBvdg0svWoTXZ3NrjpbDK1u2wP5qODs
64sEmvq6yhCu2tbYRj94jKzdnrznyHn3cYwxw+E4D+ibWf+r+jgpB67HuVVkto3N
P/fDbrs8QWdJXg4T3+5O3Tm2ZqvSjFp+rmH/pjX5RIp2zdqdQFlDKDJUtRQqz3ob
CCxtzKr47q4cUMBrSOyEBGYYCu5rqfnwZXLdNmtfS++U0VTf3+RJs1DDKZmWf1C+
mTDKpHjL666mtm0J+WtfRCRro8XC1Qbr7quJjpMvEFSx1Op/IQgAokUc+bdt700l
ifgPFlnGo8Ko5uTJoI5BeB9gAVkK32hlhqdHftS/0K63N7xmI4EkiBALib3AQTHM
vl/Dt+98v7Wdx5iiNPdNcMHzX01/gd86yjcekKlQGDYnzWlVKyZDQZbOb64d/vRq
sHO2qveQvrTT5GvKj/e18Ot1ye0HNySPTw8jx67osovV42USXImjHtwrCb+iLYxz
OLuExu+9jvT764XSngId/1Nc5NqVzvoh2d7ZTI6p9gF5Y0Al7b6VFpJwKccH5API
s+dADMCJR2rMMJpD+IOnMdtQSSGEs0QmLvFXHjVHWf1Lyiktunsedzrzu5Fa2QZ1
bpBgdZecTqie5cGm95rYIS3VLgHLWroZgJUkh7MtilUgUFO+RnBn97/js8MS7cHs
jWqvIcW2LqIGmdY0j/Cro2DY93uuNelrk+KfN66K1FkboKEBeJtx/xkKmabusPHP
eVGMg6FgbYq8xNEyyYuIVwmgSUNpV5DuW1zaazR9vkPO7SkPP35/aZ/hzJwlJ/zK
VuikUSrhVaffAyxJi12WyQUlykIbMR+VYVmWqjvgokr8srdCq7fK6i/JQPsBbFC4
AGD4/YKud2eFMNmpKD5jS96UUzIeXS6oNi45EhKXsUTpim2Pz+dTrVhCE/Uh3Nbd
9IXzyhD6lS/q7IBBPo555AeY6d8uPCneVh7O3vg4vkGcbrWLVuF9R2x5nfxaRtss
h34lpleTg05xs4fXrgzOiMRbP4//iIp2oEQeZRP46ui3E3+Zm90t0AbtCMPTdK0f
n00fuhu/dk+Us98iGXGX7LxvbCZb2pfd+TxzdH/87ts+VYYlIWPc6AR54fCD6Ct9
K6P7xliCArm0dFBOXszGbI9fgQDQWrv8B6gNrc1JHuP5Z+yM/v8OawZ1NRwxOcBl
L4fnHfKZQeHri8G3+6t+qCDcvsirWciYihSghtaCbbtlkM0+pJcu/G1B2lifcGv4
MwCKNXjttTN6XCmLVmATbDDVxk3kPfUbFS2vZpMkZdT86akMNTRZGdgwdf3ZKk2r
JDe/Bq5/Sm5CaCMEfCvnXrWonYP54zJeZSdJosWLxgjT8k6UKWt61NVXeZSTXm5H
wKcfsLLjdT+fZc4VTW/HqnsI31DtHRdpLjIYzVPKN6IDETzkETfIf9Oq+o8x8r75
XhucX7kOwwDK3Laco7xa5enA+jaCIbJL77sKkEXSwF0WCu17rwgm8JkgQEcABEq9
cm37Wl0f+yRjAuTq2ArEk3N9CujK5sItZ4J8TY5eq2JWLTusmyRmJsUuzmc/hjX/
RvY1qLfhl4BmAyL82V3cQ4OdzNu+qK2o/URuoUf8FooGk56LB2aflBnQjqEO8kbO
/JAiwzmKHHZvmpcq+SvWB0Id1dgg9MVTJSvP4bd1NjgP2gg9726fRP++zFT2d+Ci
SlhI0aMk3XkSUG+yO2ot1aBpeePs/ZSjnEYJLb6Zb3poyDmfNmNuTLwRtnCQQCJD
C2pKsoNkTiZ6I3IIlEALD8qf695DDyVbkuGQh9b2aEdhKDL0KGhbOqB4YSx/SQLn
+VdrJ/4LgOnW9+bMHplQM90wgyxL+IzkY6VkkZFEVhxPJIs+XZKLHBsze1ShsSiq
7lOsWxqUmRgKZFvwaYt4vtd+IZTxq6AjXMTIBBBmfA+TOSvxZhqOE1NyGUSNYr4S
XxM+DtU+gKBd3Su02gqADAWcp26Mh3oWlpOBCp117trMXYJh2vlKjGx0F5FH8LxY
8bR2jb2W2GU43/mdn67vhNLo1ZS64rxUYFV69+wxmSFPNxctWKCTYoAGqwU0kqKr
PDt+rbRhFnuD/2N/0D+GB6Wl4Acr6zGVHa85ObEoYBRRHaK76ARVa5F/ivhIwMRf
Pz0RXZu6VSqVOVH4FvsyQdgMIQIQLi3+gmhlWVPKz7bXhstpLxx8cbcj63xYmvlK
+NEeUpPJXjsZNU+oAbPHCIDKch5lMZC9QGysG3+i5o1pT2wkGZGSjbtZPh1j6nzL
ecwM2B3GYvVBHFzjz9Ede3NI/PCzQbr4ch/Svo0tP68UdEEJRnDwXeYIDB5/J0KF
NeSvCtb07R43SsRTNTFzqjVy1I0KK4Dp/t2AC65rWnpE9iB9m+3CvVz1fO1vJjzk
rEW6jen7iFdO9uraY/2Ag0Hd9YrL0mPsQHE9kSkJJws=
`protect END_PROTECTED
