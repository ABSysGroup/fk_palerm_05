`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SIsfjDxzvFhnoM1z2ndpqVHusbrnrhP1pFlc5Kuj0I+lA4mKuRu0Vw97MXJeoirx
ElqO5nkEBX2aoL9ZRKRKdWlaQ/jvU/0DpomL8nckg9SxUrWZIlLDFPvFDsQQWkcp
BmW/RUVeVXnSlVJ5cftJMqCYGn650um7IE7uJeG81KhKPHSVtUyF/hQLOS+yfRMl
eCEnWpiW9c1a+GtB+SjQNuv68z561AI63oLCm5BiD1YDxMkMhIu2Vz8b3bFmfTAX
DcL1U15UtU+AK8dLb/hg15vOXaBTrlvOBGi+0jLNw+hKldCl8t97jim4ZrdMhF1v
`protect END_PROTECTED
