`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d6oKAfYu6f9IRdChJEmTIEBgkQWDjvgEbDik8GYs55uH1fnmHmSQOJPvCtZsfKdW
L9sVClX95RZ/WC1MFKY5BOdd/weGRwL5ll7RH4aQ6vgpiVdpYlQA7+6hk4jcxT1U
POJMybfFp39hs395MqbkVuPzTp5K2nv0nm1b5CxtUARqaojduPOqOSwNagkHStO3
uByMstYV2hcc2GY6yvp6nwb+vp7GWQ7dpFp+W+wsAPOQvjJgCmLpoo5wVc2YZyou
Mbzq+ertHIW4sKWCt/mdicwjVEOt7BxqJDR0KR0/Gj1HDDw1nHV/H9Fba/cMB2b+
bGN+jLQFuR096F8uqJaFVsO20zu4RDNezImhUflfK0CIDjnexzoFNUyzXw4HK6Va
ERvVmwDSsgehseTGc8OcYNM71DKR82vtGTj9Pqm0pN1FF3TsawZe0SaGTnkRKPTX
`protect END_PROTECTED
