`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a4/XkovH3ackN4z4SlAKn3BH/lpaunZjIYmYzj2VBYt/0zwiP089LZyYkMeFACgt
pJIkWI4PQFpO2JBHBlLfDkbIoEctIeSixWxrDUbhJBNMUeiOl/GjtSi4admZ87jW
sENsxLdeDdAYNW7hTtO5r/FctbiRuq4K8rtgPGx/Y2c6T2T/au+Rc5lqFK1CMIyD
6nzfarlFoxIsRGAbqy38xyybvnbcOliz+L/djm5hvghhddsU6o8gAg3ufvq6K6XX
jAAG5uhDVFvIaXf8APbNWmKiq3o6pd1GHEL10mKH/ie4GvXh4+onOvo4gBy5QfOC
Gk2wtndSnQEo1dwCKSM5GNKthtGRGshgePQ+YsK4gbhsYIrVNRO0PMGwUKIcQkpP
`protect END_PROTECTED
