`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MrsHOn4zuGyQVFXfulf3u4xSSWPtC5v/9Scbc+IVwQOaJjnSvswZqedJxvyOX4D+
urStTaZp0otY4T+/9GjP2zP6w8bdabQp0lBvxiJrH9tPhT5bifGHjM1sTFq+fXIZ
mTH1HiPEwlw0d4pYtnxQHVa656GkeQ46dANz+fQJGKLrjUfcouXh6/kfkSBoY5g4
RXnRSAGRP8j4BganJFbUOV6cJrJi2Xb00h9p/dAF+gnuUqyc/gTKyAXLicFs2aer
02AnFLTnfWfX5tX33lyBJ8x7smEoq5OTLUnkcqWOAd14cpUF6k0vSDMPmQwoQP0O
RiyJuAIJsdmMXQRCX43DF3rv4FwrZO1yB30+0Hu1ZZRGA7IegDDI52NMtPUGgSjf
yBZ1HEWpAI20o/mjNyiv/1yQkqHkkrOYmC2Eh8PWdFpMRQPWl2e7UFl81Hh/w7CY
Ik4pUfhDn5M4hoIiEgUglbrPDpvOf4O4sV6maZEvSVcU+LxY7bpEm7VI0GINrq8b
y9qTCZlE5M9vpQ0sxpzJvL0rDIHYQB/zindCeCCsKAA2uzAaALcSgtKgWCotUpuA
j5abGlThbx70RSqt1LGL0ZCJjCpG6aY8gsNjyljfti6ZOdNGVo495EJGTaHA4noR
eYgQPmYKcAgQunGTEeAvLJatS601vu0rItOy9k/nP7bK57ZZxJSdPrgxB0V+4FLI
HyGJIxEnWidb5+QKAZm4SHiruZaqDl3hxK5O/n/KN4JNH8929tHlLFlLA02lcuu7
ssOTr1QZjzPNHvjcg6pvwGueenyd8i5V0vOBSL999smqHlZA1NJnGwuw4kCbCCmE
5V1Rws9sPtWNfsyz06vZi8u/clIKX1oA5xlZFWVc4Xc1ircb3XbfBbZRtKUBx7JI
uCqr2c2wjMoOW2AclXYg8n8aeDiZMptXqKsCZlFpD0pp2AhtjSHSdvSXtapRiiJy
03vswoCMNEY1zzTEft23bR5sACpLVRnvx+2IxPosGTtfDTyz3++MamScSm/iJJfx
87nwhNURXGey8BnIjtQY8+DDMwy5KDq0GuOU3z04HOPxSHXvZaHWd7mXln/J7Kj8
kEXzsr9Lp9I/nlxdUzhekSCNuMVY3FO2W5rakvYQiM83uUCZeyWHKMDNyVIN7g3i
rhkq0PFw4/ZAJdflcHOkmt1z1oJjlPAY7FEn2BedKuLDXlLmoWmkfD9jZLTM09ms
XA7SDgX0fK8q4H1LE6+OyywWN9WSzkS68Dv9yu4hbl9TLShuHx7wqZiY2zPo6Ds/
bdVv3gwAyWGdH7/LEwPqKHrP2ZCfrPpoQGbZUC2dF6NIuWNXJFkWiJkEgj1Zsv9l
YxG3SgnW1D9+EToIMxjyPV3ZeXank5DBvxqxNKXr+vqIdedsNHaleMQMagTXkct/
xEYKumjzu6xobdC3DntvKNhQlz17L45cVvkhf7B75v0zYDc+Cb8mU9jSkqlB+oUL
+eL+Hnx7/Pb+kH5O+otiYw8yVkv92sKSlBlk6NsaSfMd3ooNAqu/cKjcgmVkv93S
+IxbVobBUXBxQwyfkIf2L+v3D2pMtQw78v+8+YAGQHUG4CM8yz8pKWXP8mwHBbEA
NGm1xl7MMi3DXTUI1tkRBh/0jlzMvCJSZbW97LjH39L9ZFQ0wlpZGfGVzjb+Rhkp
jcr0Vkd2hIxfAhpQdyvzT2ch+23pjO2OiSvilBi52Sg2CWwamaL41+d9q9c8/Xqx
6aF2dA+pSHQU1VHMd13sAasOsw0xA+oQOsYG40rHwFtbvGAZmuHzIy1rMzQ2GWBk
Rkbs04wxwqJYBg7kBt7n/hKXCPkZ4eqcJvbJH6LVrC10lYv1mlGbXAeCxaINWtxt
pMQjRdxoz9QVsIjk5lhBKthzu0KK9cU7731c+RvoXBlG5XmXSpSvD5z9w6ECs3UN
8ZanqMyrkUx19EBqzoyBW6Cmf1aOrnMiyIn6y47PBQIUJr4Rl0cMuGj+1h/ig7cc
BHyU3x/PQIrxI3x3Pev/VZsjjSqZlRResRnQytJ78pHtiQOY/sLpG+7AEhr4LBfA
+JwO2Y0fTFir06mpLibkYghVzlnZ5olfbrgLcfxnTTne/5K2LozZPM6zWh35KcLr
AMIr08lvpeEdS2MRWUjsow0Hg4Zao+W4QhY9YWz+02YIA+ajE7cVDNbD9N1yg59Q
gmxheS5jbVphRtta9oZz6PHPo2KEbCmYRKLy7pDHUn9VHVB+ihRWoi187SlTkuDK
RquCIJHSXheqw4fzVA3rKB9O+8lnDY/JO+v5R1jCHtxhmO4EtiFNTcP1/b4GYpc0
mH5DO5jukERGqcopdyT2DqXJvbWX/0FNu/N9U5wD+HDyd3cRzucKelcyah2vDhPE
zVnDItwqHCd2dYHZFD+gdwzey1wlBCk/HKrlJubaJUWro/dZ3ZN0bdZpwVodRwg1
dphsqRQC1+PA2ilNkxqCF5DpeJC4yp4QBJly5J8NqdAij1JjRZ2ecEhPKzVvJUd+
VpAraR4aCu6wmuMPNa8ZXnWvpLeCXo2ift1jLLwy57g+Eo0EgM8ST23f72IwJ07F
a0fZMtSKYmrSAQKN1ngpKv1d5NcT8KOHZC0L71OnPsvTSyOgH18IwXWc8ubyoQQY
rIN4NTo56ZHcq47cSOujWieiiIrLUWBZ4oKZv/eNOsttZYPkiloQDG+EquFXncf+
5gnL0TarvzF4QyWqUbZ4HHZNbnksi6F2WhCzMMxADJ/2KQaTU2FYfIb0jbc93hlR
OIb4V/9SAsuERU9E/qjSOGIWMhJsRV+4EEF/19C1X8gd7OQxLy9oClN7inqHaAsR
ljsdXZjXped7NWG8mlVr9yphRiBidAQIfHikqX7qZQdBQuBX63xtJ7RpTn8u+jmc
xfX67PmOelqYksclqyVznDiVBYAwsSWPalWlKonF3KnstUqDCvdHHtX83l/7F6gf
SZrrDn+//HNnui4DJycK1jXAIun0MJPiuxNFAkWDOudmf2lxDx6ADyKaW0/1RI5l
3JgNcklJS8iPfvTWBTOH6rUXEWzjF4JJyXcUpoODP4v+cUq426LZpBvDFy2v/4cl
2t+5YUHs4r0vaezLZC5Nh7RrucwkBgyoHME+EKtvJfvnq+pFUjSsDo4UwLOtQIBK
3Ac2J0RVC3sUxbdp+STGnGda7nPrCHSC5HQFKeL40683D7WTvDZiTYVtsE3cP8hi
MkrkEf0wu2ILMWSUr+Qz2qAYE47jOD5AUHRHVjQg9HmNeGLUDUYKNZ5yb+QzpHoN
dT1K7ecFS5PfpRFcuXyToyqR4cr+ffIK+TZYDpyt1nTEB+tRmp0MeklDoIr6+/By
V3vmDrPJl8D35eHRibSRtytNQUvyb1uDjfEb/x/pIgcxQdRtxzXX9etDBD0xqQbu
Fq3rqKBHy+O7XkU12vTx7ig5NEQ11Cj+n8SGzMBks0Io87B9eRTwx20G4ZflvqB9
2EAR7XFnYyIS5WeCVJ5jOgAmLu3gygVMSKzqg3WEKlTpw6HE2V2Fg4ejR/a0DH5y
NcBWnwXmD0dXutesK5KECXvIDVUxk/WT9C3kx6L9r+Fl77fTfTPtj6PXMRf1xFBv
xBstDYncovCncH7h+npm6tYopC/4ZGxMPQpdJ/CKzHU=
`protect END_PROTECTED
