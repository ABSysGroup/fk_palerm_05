`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I/YuFjvPS0bw8c423Q1sQ3ephTd0EgD9MenL5vyS/FOrdWMaV2EAFTgnmx7cJccK
c9Yx9JaEoiAOAjgDEIYHmfZ4COlbmk1DVm5Dsnyf05cmEmdjoYr4gyZTQV7Azt1W
W4c5TI+5rPkQVqhcBEnTkwRBvrg5Wv9r9wV0ux8LB3c4h89B2eb+bNK1GCngQs4A
qzkAXqRqHIbEbd3W/OtgCcgWZ8PPIUjrr6qKR7IvtkGvbdT05uXfzU8Pk9/Tdrwv
8VX3bsq7sSxi/xaW97IklOgqfcvTDTvbdm5wowrM14hre4cNbzWvf2ixLmCd1AOZ
+fZelc5myub2L9tmD3OAwcmipfpGzcTLbpQE2M2q6E/+rc+wnH4mkUT/S9MKAW0m
zxjKDQZQi+K9yxZtGKErdPv1mqjywTUwcnvnpU5u+zHymQNWHroC6MUPoIJfQSXP
Q9Aj6PBx3t/6/J23V+LThDaPAQ9Do4i8y5lylTHPNzDfpVNTBRbMEAqWB4HMgfcN
ruumyvZ5CYI/x900ZPIRXSCiDjF5e6yJlUS7Zo8kOE1ICbWxH5+UFdhrtuwvNM8t
t9LUNvOAm9MAAHnTXvoRDmRlW0LroL5abxss0ZLYz1N33MEjC2rd/CpARzCG97uQ
DuBL4GJ/vhGu7toRQHCfe2f/dFiHtAAquDC3f4VDZjboSaLToWMjifZ/EcculupJ
F6GmWDM03WyojLkLK8ghs1mUFZ9e3aptSMx7okkuTPG8aBG6CpJeR/6MB8PQGGmn
LlEYa7GrbX/OAyx/4ATnRUrcaiJlTcvSJdr3AbZzhg1Br1tUFJRDcoSjVRJvZOtL
bVfFD3yWy9vVcyvYcUhl07zoaL8sbi2WTNwnotkuQByGUksQ6mePO1/VyjBQKIwB
1RYW9VP2ABqXuBDysOTiQLQTTbxX7zDhHmz9hovmY2NFsrlf+J9qc+K09U7hq/3C
CgNkLzxVHZUq+VAk/9ujOi37O1NPp2rZLi/OM9dJB9+gqhJRz+PC4uq5jBp42Gk1
Z/8NUcSxSiFTkZJkMN0emhLnV7LnztY3yBDKiYGRJD6J/7rhkI/NFU2yFug7K9dl
uvnqpa7kQQWh43KtvDcNnfs8r14ZW9dvN+76V2m2JtIZHR5mQTlLIAEMjBybK698
/jlOIM1QPJY4xh/VYLyqP0iC/Fnfte4d1A0VcAqfi+xdV+pbIS5PA3PRhnpxlMWb
0LwnygC3TBc+1ENpdQdBu5sUaLDGXLHmxeauP9jriOxcmzQJDlQquZ4uSyKvKDaW
TudslXEHqSmjW75sD6TGuExCeZ/jo3scOYStbvKGzg+UR2QoNGPX2ilz+ZGw7eU7
xiCrbFIovD1MU6wlTs43BU+FrzdZd1YjlSvc3LV0WeZiGusk7VCV8asR4kVCTINm
VVQ7G6Y2GUeWPo67+lNqHA0PFw//IGDfAWhKn9OxwT4zp62DE1R9eeku54Jmjx1Z
7zhIVrM5PoD9TJlCzXXsaPFX7qqGhEbLfB4HEMLoaXYnYo9shFrdh9R7Dm1fynyZ
Zw73HKsw2HWt9TsV7NnVedlNaRVRERdW/hnHgePKwSVe2vu74nPlqOXilu3uok4v
LJd3LZcG4ZllHjdxIItawjVRHbFBVy6zxbgppNiFC2nabQqaPM1F7hPiPUCAww6m
WTPstRVKMeyKl9ZlavitKknbEM/cw9R6aEgPjzy0VgAKiNTg/TyYUT8G3FBdxP+O
f60ZfeiA63yfVTITxsOcDecCxmp06P8qa0rOn4fcfhDpCE3YSwNOAvgimLB6VuZh
UCZepByxykxgU6ysx1qaucQHKcFtuTylW8b1whKhC9cx6mf88O7hbkcRNPFA+XQa
JTiVPbU/nNccnf1fi4P8TkwndiUlgdn+5AOCNDOJZI2Vp3Ohgu2esLRaTXfDh34V
Zz9PP6631PnMajUXGUHx0RWHfkJV4BEolTxc1GxGF1tcz0QP2BdGlOrHo8FIrrA4
awOjn7CMGhOyEuPA1YQ8CAf1JxIFpExsO+Bm13NmkBHnZ64rrE2fLbcY3b4kqQir
PHR32qv3ggQh5wIG/yXRKp7ZfhTkGEp/NXLimrBgxLTxOiDpFSMRLSHqdius2XCk
TNUorr0M0EyKbamfKnMGD51BMPm4mDOLRUYS9DL87StHfakS/GrqhgK+mSoL9wAN
MO8YBaARQYYZugNPvuqSQ9S83UGto5HYHCPuSZoWvQD+kkJkq/Avw8pOa9Zm8J3G
i0GvZ+Irr2rIkl1ZVYDFWRChmTo8+KS3PcN90OqFd4rlk9PLLawa3gxk45NQMD80
F7lKCsDsSPgZ5g7iA5EdB6zgJlhah5wzGv/wFfZ3m3NFTD8yw3TtJe6/sBLkyLmO
Lc0N/VuSTlHdBI2rOhhNmW/3S9YkvsCBFp4r1Q2h0Xb7MMyvWJ7WdT48oqxlams9
ABUuxKq2vOGFpKaYp0pqTE1zjrk4LogtuiKlnU5vQgjN5qrpfirbKcD+y+hgpZx5
Yte8tVL/mz53LLP1ABmbDxx4Upr9pVO2vCF9K9S9tjfDd1qiqMXdPMsvDtxhuuyH
CWuNX0eL/gEPvLPGSrp5+g==
`protect END_PROTECTED
