`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XmhAaNiZOLoZ+Wl4pj4r80/wWnIKRIVN3S94lRxIJAEWUtI1h4wvawzCmQl8xseG
uHZPSiT5spEc+4M5ZyMZFNCVXAiGQerYLERIJgMFOpY4wUAH6Zg7Ii7mArbZMga2
3i5LVa8xnc6DqK4HVRaKRJ/aThzQD0hNKxBbn0QbbeipoV0N9+qXN8d5byrEg+A1
WplFMuhON6sF8lVWM+cJMsvfe+vgb3PMKB7XJYs1N2N7g7u6QGlXtVRSOAbx8qAs
UkQG3NnE+B0qB6felfb6jYbit8YC7DXilPojBhA0x8yWvmLK8fwjzQNEhWJAFugS
FWdMweZvjdAKlZDq9DfXw+n6/DzLbr2CZfmhwN9D6MiDLQqvVEMU5COuHh3mOYvP
MnQhEKfkKwqprx7aI48COntZGGZBew1WXsfbzI8WqFcneFmtnRtqFjvvzi6y9uib
tWY6zn80SfKlm3enFOQc+g+tbfxcbcwo0vEpOjUBobaWLdczyP0xfAnWrqrCcmnZ
BNC7WuVc9VEx1Kok8ZgNUs2fS4edoQWMM9lQcNCqyHvbYB3fXO0ZdAsOLyyCz6N5
6747rBm7L1CWgQybiCDhs72IvxhRq1hqiCwAyBiFMnc=
`protect END_PROTECTED
