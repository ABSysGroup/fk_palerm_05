`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mJPZh2y/yDAe2D9m3p+kcgpn82FjyMvLAlJySpCCD9X/pAKV/FMJelf+6hb0ThzQ
HSk29M8b924rhwzLw1FKJq3j2JGaMj4AwlDVJGqGAWHzOQxQKgxhjQlNYJgANpd3
xdsx3MO08uhKS+wdO6wy+THrr6sNeUl2U5otNbZLxDtOELvxLq7tV3gyrH+vQBVH
urpqPBcNlssWyg2tQnnE+HOSUxvVaXxG3OtSUC5/gdrwu+5LPsd48xCKmdOjYO6a
fXz9Bhrl7TcJP1k3yf1E19rux5Iwt3fHo4gB6tRJMLHyc16B/G4LrIRkcmDgoadd
5DYH6uHda0aPA2M/7sI7mn5W0/U+W+jVXcvPMImw/Dx9DR2E6s80+Hvy88WQOZw6
QTZtKGy7tta8mt77yH7aQPkVVgM4tT7TDLmrFIo00e5wtnIhy2GUPrb19fpAu/Xy
HWW0sVf48GiJ4iElqZIuIqmuUaozf194U/1elJUcDKHedFUxP12VDByAlyMuKMih
jTnyAFC77f4L0qWf8oZZvctiW+aLD7JqVnI6F8eAUSAWK80mM+iSan500h1erDkD
z/yoY/En9iCDnBpGYbYfRQk5TxO7PwU2PJN/+xB/10m9cOaZG8lZclHQMBH7hN36
wtXezjUOZChZnzFLtwuHBG/hcSj7ArLiXSPwSLGe4LubsB+MsGV38G7dCIuYjhrb
H9ceDEoUuSZyjkWvykdXc4Jfj6fo/KBFN77EKbkp8iBJUe/D4HKGo2e9DHM08k7j
IfOegS//3u6/uctyYGjEvEd/09mop22orKteIf5sAmE1y96kNG1arZSkuwJhDxzY
UBcLn/SG0rYYrfVHsdoY+Xp4U5v0OqY0AdndCvAX6KL9tB/h3MwNbD9lpAMeQF7k
qNhffsmAH1OqqUm8Rp1f3Q/wfxJ9xjkTAw5Vzg+wg675ExFNuaBW4L46qcEhnLja
ttVnoyZWIxkODRKCMQ4o9EyJ6oY75Z9FRXbX59TKeeLz/xvX0qmJDdXUWcLDvO7N
LVjhbmmD8BdRbKT4FW6xxNMDQ+OHEZ6SaEo/l5AJADD/VWIB6wERN8q7NO0msY7o
+Gm5M1laL2bgVlFWDkSQbPDo+2yV+l25P/3zrq8st7IlJen5+UMWkxPZZPbRt9nB
L9vWbKS2d6ovq/73wNwb6rN5k+e1IhUj/XLTO0DC3OtjmUWAewEMZPalzE2+hgBH
tbgDVStQg3YZz6Vnl4z2Sfff1DfuCKG1/M5wyqbp+alpojGbA3/IqIWJVx2crkQm
90NdeUZfkJ5ztgohXSm/QlBtAG/TS/7c6FHWVXSa8abQ/uDphAQXD48AZXQdHqMr
UrfImeENt/RIduyx/rpdUdSloZWB2D6lnreUMYl1R3g8qa3O8mbO4pmyXF5TFojo
WJZ4ZUHot2vUKyR3+UDHpDLo10OtmtEDQvS5FpwwU+SOhgalXs9Xr8VZKlh7f7zj
M4IPR72SBNf6sW9hi/OKUFIPDDdBBK7nY3Kvlo4mZ7o38LROGTYJIjgfDTxPvua8
jbwG+dCXDgVM7a5z9OtHSH+d/mhyTFdHL6Fh4JI8SXM3+DSNAQb6fdGAl+h/5/vZ
bx9NFAdohnOWnLtJb1NKhkaqRBGgQNbbmn6fBT8uAGjgWzoPro1uP7m9asZpb1zE
gzO5zUZXtfczleMhgflB940lBakkiwIj9DuPmuAbmSez2B9ILov4k2i9pYKJ1d/i
uPKtAs2GimIoB4c09wVgYfHSsAoFKwsOpj7r/nlH8alEkaAxNcDMKVWU0fr+n57x
mLL3VBBL4yjNuSjsPSzsD068wGsOIA/2VnWPVoV2OICZlBFCR6h3fV5OsD8iTR1b
G/PHGfNMEq/cBXzHhMXlEQiW45zKfXDa0ZukYX/aDxBpi/iOpCvTDQAxA2dP6ZrU
GHM7XFwjLxIJW8exzWYGrNt22UTtNxlOcfPvVuVYunbiSgPAuXS/I2hlkX90Dx6C
x1Vu+0MpHznjopGZwqZeiIS9IdpZSTSliFjTWFLoGcYU1ZL24DXo0yfoApaAste6
IpwMRNYgsK+yFNM017VBU7pMxpih/CRqz7OppRsyZZD+RZIVtclxgDyA4nW9tn6S
ulfJx6L9r55ckjTOiQZd16Z6zW3W7PFbpi+aq6K4SNyWLHzfcGDkkg7jwA/kB9RS
jiBtE45NFNmXwVDCVSoD413ont7F1BccZcgSGYWV5KEGE3bgdfCZJsf83AVnJBGs
iWPmGEySTbXcPcHErfF9dCzLKMIUSyzMUl7o7zhY1apI66vbTdOIJ147EPbk4x0T
n7EsuWXjib/Z5KiEJpI99MG32QnOFGoRXKLZ81WjA0Y=
`protect END_PROTECTED
