`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YbPqYIZdFdBVKX2eBB4Rd3crFam7piM46DI7gp+bDji8kvGTKjyOahLbq6J8magf
wHUDXnv4uA4MnVU34kTSHK/FLwQM3JhZAjRIy93ZfXBH/r89PiGkqjsYHO5mzGXo
0V1HF5U/p/BFhuCJ30XoRq2JTqwdQ54Yyc9/M91W0GXiOBZb3RHa0AOjLdsJu8hS
0M6R+fWONx+3J+y8rG4b/c4a5QPfnSgyvjhuzlLSMhxRQNvZUGhWRRx1iKl5H2UX
lXD7RiBpDrkF/OQaNoBC08RGK2HARELgz7gXm1kJ8ToQn7LGt1C/Gejuo2NOaTek
SI2josbl1I/yJdXjd47z51S75Hr6ztNvLJZY7MvQ0drfQ+DzjjS3abugwXB8qIqd
CC671BBUFx0N9v3JmgBRJg==
`protect END_PROTECTED
