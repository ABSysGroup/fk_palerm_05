`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y92cFKPa3pTmQLDxwEW9ZR6Ca1TTWhXYPSa8Eyn3JJh3qXcOrimV52xprLnTPNOA
WdSy917PkyfYs2dIhEDHKai+8GmiF19ELKT3fhyFyroHClxCPBSMReKfFNR6sosc
v/tIhGA5vRerfdotdRCTPfhHiGwS4x3/01S3VI5gxZXhMvLkq8Q7+ub3UqW3CnFh
fUhCakX5yMTY2jhHIUEI16PvaToJWwYMD/BbU5heEW7DiSeSPciVFWAbSeCir6eP
erkFZoyCCVSGw5W9ldvvx744OgMp4i3OpkAe5jknPYpT78B8Jwmvcn6vfLI6zwlQ
mg215u1RiAguL2hmmCdi7w==
`protect END_PROTECTED
