`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mkSkuadJ2iknXwN5r4H2WkppfjYkHQraAc2KG7J752Tx/i983Jjzg5ztFvFZXfwR
upSxN/BAd/Q2QyZGUHcSpDF6+7ufIjoxVJJPC7obvSij7TuA7jCEdyCzTQjqNmYq
/zbd1wyyzhSg8A76IXHhtKT9Nt8mj2HuKNT30gvSXlf+2ULrsbbqJk+zAk1ketuS
uYmmHmdu8ACQBHJgZjLNs05ea1jSMGDRcXhemMJ34J7yfQKWOmCRArICRQx990DS
BqnFM/zG2lluzNd+rMdcyw114jZSguQHDTMIz1Mru6BH/1Nux7+XDaprW6sbg0O3
SZjZSPgVEAJCkASnsUjUBfA6f1atJSVgfsoFgWkvrKCyFUyOqKakR8QPd+/uohAf
nbuYMLL2gGbMMhv0wH1W3PgqL82FqL1GcgJ7IMSKiUjUHJuwsNgJU7YLyM0TvBSc
eW0o4z9rVWRbuZ//m+Es3G41LytNoEARmTFu4K5HuRU+qk/PzA7CvVRRuKvBLPnH
3ywDckUyTFsAEfYYgMy7GwOc9jv1v7WBho66VmkeiNHJsOItyM+ESDf10ye38XN0
`protect END_PROTECTED
