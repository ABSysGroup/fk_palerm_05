`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QWMoqApOPyzTpQehjQc9CeEbJZgbpgESV5Ppmu102/mYCBWi9pHo/jvZVdjXuJSu
a1F6BGgbc5yurCH7NIbcIwxHLmaNgDz8N7r1AogkWqJXOSk2oS1d6WR8Qp+FSAdJ
QdRoZRGjFbUiMImucB7Kd0AY1Af28wY62TMt3Rh6VphZLEvOysmKQ3w4rB5jer+A
YHhCcnqwhCnN404mmt0Z9gw0BGNBsKxke2AWB295Vk+Rz2BEH8SylFGbEiRk+9b/
j7ceZ8kjbI1ImD4s/apqsLELZhzr67onwTbRORZC/ci2/JdqNKheSuw9di8LQFub
nQA3pd3cmsg1H/Nqz+dJY9Mpg/47AkOd4s9A1iDtpQuEEyEU8ULJeFsrz5TnN9T2
Qf6sojZuHYer8y8pS9jibyM35sIjiIF9uCJNGzHP5dYb1Y+5bpX/I5AtWmpXb13a
J3ngAzffKnlj4b4XHN3mSlRQQxtsrxmv062wN0vXgoNYIV/EaVwOq+LvKbEQ8v/4
LgpY5UiLlgIsSCRnNDc+hLumehY+OvcZhw8jEojgnNIt6RZVTDO6mEWFWQv2deR6
mIj3QXvFRqKqu4XVjnvy72IIBhQyAQm7qE9UqKFPXz/xbPL/Wco7PgdBRx2pyETW
fsH+r8iNmwJ5sfdTvZGDajA2mp6wuKARRshKAiApNqOLrxjbWtuptuzPFzbzx3ys
xTL5pKk32Dxi87J/ICP9NrJTQD9fjSXK5/DE1UtREXKyedWDw0x8EivtRgPpJUyw
CRDqcGyldkMmrh7nIx70EyRzm+kOeQBvsQXl8M7GzYqGHkch+22zeG90vmwC2Hbt
xb3oZ+0TbWm8BnzSkEn9/eah+h1e19HFYTaiSPUzRo9vCLT4aD/tasjp0cEWHUKx
nUY3ZDGPMgz5GDydGqpiOtzLofNuoR3+I5oHNDNu06b9PGg7j3n2F+STvBpqRQvy
t2nU237UZorh50tmxofjucsbbzxo7lm9g3Ty54N3xT5BJlU/kIThfzvgALPd8KWX
`protect END_PROTECTED
