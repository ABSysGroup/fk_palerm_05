`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XyU/wIG2I//VosaYAsl1LrQOXH9H8BqoLMswXQ0VYPX9gdl14r4JZEfMZ1h/ZP/o
2pKe45sGeZ6zVW+GWxmJVy8GXxHA4cfM6rgO4t6JGEqRvVXdWqJLSvX0NhUvRsEj
BDlX4LaBnMv+j4ygV0Foq05KHigugCfNNyubgZhQY8zzahPhkW0VrA6JCP7vYA/b
t1kTYh2rTa8dq1x6Y5Zq8B50CHWCWwuGkp9pi2U93UjBbnj3DqdlX9a1/Emw/WRC
gj8+S5EgHR5jJB2uDjnR5vl55owYMqxEFGkRoMRiuu6Ky8TlDaII2SazQnYc8oG+
bgJVx57bmgnfFWCFBuDJn5xwoznuyByrDNxzko6rzhrr83nwoWbySFze733PLRpC
JPwRjmFxFjws7dnrLVu5WrmJHQHSAQ9Ym9HolY80SIYXqAiOZ6RFYXM9uWxAmyDP
MvZLKud42m7FF66RUCIyTO0e+Opahaj9QsDD9RyO8MTDROJ0Fbqjbu5s9Uoc6au1
`protect END_PROTECTED
