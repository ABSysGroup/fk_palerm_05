`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e+QZEgHaB1ZHRfO40sed/IUQw4OsG7dIySfRlhUn6hHVkYxXkqXTRjLw5sbcnOJz
Q+thQ0/rdaJrbepS1L7FAO5UMgRRIENK6JeytE8Gc+EPd9MjYxfmNjvFhI4Bz5UM
4CjiuqXxFAAhJZpHAVwmWKJdnVv3IOpPRhsBKFamN0ETqLBxUdBQ+TXG79sph9M6
jxpYkWQLWioEDiZo9feGXNEnUblxIT2gxPyfgn3CjebrF3Y8oNOp3WUqi/hfG2pt
z/Q2JNPZDpgmAfWvU09NrYNjVyPSHOLsXp5F5QzIcMxnvRKE9sNm+YLSYppQ0rhK
+Nktzvu1i+PjUxNxEJeuOBHbw6upasRqWcLiIVdE4R0w+Odgfio6NCroEHFbN6a4
87wqbEFC4LekeruoIU156hb40q8pntLLZVrOp8mm/KD/FVhB+lXKgVnbO6Xlzc2s
xrSqkwYxBgDeeJQu2lN35g==
`protect END_PROTECTED
