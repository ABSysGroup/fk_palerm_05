`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ucl3hbFyqpEuEgMkAHs3qfMAClY8IDMnGKSrQjwioBduX2qAUbCwIPBpCKiVjJ0m
GsTIfftfCLXjAQc/Pb7ichQgQxh5+TdFiy2/HsDr1g4BjjI7cIhoU4a289zlER+9
cSCJ083xXQMEkVDyMBy/VoPyzNlPXm7ttugAAwkEp8fmEBuckTksahknEeNaB07+
ABVnAmvtgp6Pmq64tEQI/LWPwE/uSyhVSXkMIaUSlh1/QsGXiddvFHm2Dm/mGWdr
VfYytgJpYYwLYol9bCkLd3wBMEOxuEshWD/xMyDHsMyKIqv0hL0zFmIVktTUjdWV
qr1QfnixegIgE9vauTaS42eUaaM3St0NoZUTCtCAvJpQ43rrXZcrqW9fDQECsb7S
iypvWmWJdM3Y+PsKuNjZOB32/gNjQ8OS4zk6WcfbNC9P/4NznPk3ici6hcSKiy2C
QUub9gVLu1CRE/xuRdjKRVc5l8MeAgFvrqVUiMsNt4w=
`protect END_PROTECTED
