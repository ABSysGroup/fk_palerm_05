`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
quyFc5n/XdqThwthXQj68bnlIB+G3sfa4k3vAL4i6c4PnEQzw+yoZjhLWw892K7h
ebLErKVd1MfrnRAtsDge40nI/LSDk/ea5JGJZ4bZPPOyJbvHaUg4TluxRvbClglo
LnMZFpZzmgSQQM4mCi8z39EVhl+vU/hYauw4VhsVtYNpSbALvYyAwZ+y+okHoQ4g
Oqq4rHjAp4ReOQCrkxjAcdrxrjQet8d141qkOGcQOJ4/DvyWDpiixLM1VuFwCv73
/EoKU1H3tobrTfUio3lGJNKV0PxcNpBYlBSZLzEIdFE=
`protect END_PROTECTED
