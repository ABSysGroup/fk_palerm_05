`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gyfv0yH1z1tJ5yFMG3AlcSRti1NGxQlQQOwRFtSfB5YOFEQS9U698w6eDlkxgkb2
fwWvjv7OPUcEsIDJ87HBrx+yiHLoIHZCJzqVIjbkmao/2tzlePUuO5nkh7w/hVAt
qLS0VWgoZF9w47khDUlyPgBcyWrMPkPWexUZFgLnjZ5rjFS0PrWJ9JJdcR7bdLZN
9p4HQ673L+s8dAMIQ9ZNbZ1LRPVwIYdqv6StqQ8uEBhSZ4wQU4AGQYc4kuRa7IFj
qgSxJ2nqq1Whc/kAkZJUOd8ooBq3ZOHNzIxHctq06N9ja6bSfbDmWbbiaxF4qdRc
SoCcRXfRGmHrw4eqQZK9KB2PwHjm1jiN3x5myfkx+rNMs2yMQzWoumy0AseVP/I8
`protect END_PROTECTED
