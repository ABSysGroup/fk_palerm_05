`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+RW5aUq+a+LofMvEnQ8YKY3Ixkb5wJWOFJTdKHeyazQvS2AR4rorFBuUPEO7YpGL
YasPuDIs0zetvb1HBlAEbXU/3NC9IlDwtA1j83wGRiN0Pp4dgpA+9q9mj04zpoYj
MON3Sj13qIyejS8C9syr8tYD5EqRzE1F8EUtIzOADFAJs9Pi9um7vlCR2IQzUSoY
I14laYuN0K0Sw801+XUcC85MO+NDBbzUTh3aKkjvXnEJPAWZefkPwWp0hJFh33J8
ci6Nek9Pw7pN2FNVxUto/mtDlyc1/R6eimcoAKfld5eFH7Mc/AVVO2PuTKDVeErE
oBjKU3VKY/VhZ4YbtOmcZkSSZnGCEWu0Pv+huXaPQKHjxUHmjWa91zhdzshtOqHF
`protect END_PROTECTED
