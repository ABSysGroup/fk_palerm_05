`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yLuPtYmcq8Id15e9rWy354FxsPRtJ2aj5Tc0fLVAZJkJd6ZhzVDWIlt4K23XkZtq
xVZ/P19PkqAHLzBwidyAQ07vvaC6LzxNcCoCUelnVn4y17XBWOQFPW0IoXf3wC5c
/pEVbJ0hWxbSj1U+Abjlcuhl8rOJOzOs9TegbaxdP6FhLyCg+IXBByKdzwC3mm4V
6XNgXiiTGg544pihCoW6goKsSgUbcttDvJNDmKc7yf3qvRhiV1oXIXAZ/VNBzYln
avPOvqBVra6ZJLpa2Yyu/xxzhQioi1peEp/u38+KiJm2/lGn6LIVaHdQEkUwZnrH
p7K0JOUZvAGo2/EhZd1ONqJjkKkZg+Q/HGdI18uzva1JI6sj8NtZfuIafrcj6f0d
51Lt9LAaYDu9oV79BKlZ/iT5iWZqHFRK4I9lobP78U7pbwl2LW77egzYNjjwuPe1
GdvOVg5OS8vFZ3So/yUOPDow+CB3h7azM6DUis/P3kDBNrodFAmjlCyJR1cjbHWd
Xbb7W0XpIFyeH88JrGn1NvQBJxosJMwOBnEbjDwCp/tqfGioYR6tZAQ53zQ00Br7
YYw5HKiuJvp3SJs2UHQTKbGJyTXLuL89Sm38LCO6NyduISI6SmOQgxBxsWgBJIln
Xhl/Y0mDTqZ3UG+7gKKH3gcaKrpLVXZn3m+q7pZp14q4LnHD4nONTfp6Qg0yGdhg
b1bc9PKEQYf2UK5xt3CV9gKUAAdpf5xIECiCbGt0M3k/d6lvT6EgUy0KUHW1MITt
67KsgsW7NiKE7dU4zL8rh4bIvT9pKOqAz5XPWawREJeWKl6hBlh+YRwNBrnzfuOs
QzKR4B3blR117WdZMbRjXe4bxkkKkTuslGgyj+mqR0dCZ0mLRAtJJTL8AOMRfFmi
0MccrzPQ7NvKSBZhHKQvKjm9XcUkFvMIPAYLdNZIj5M7gTR/3XYRUZ3CFCBecrrU
gGORXohBsLpCTORiAMBF2SOBnSLSlO2iv1DgJGCgRuba/0pEn1qAVuAhtuo8Csyt
ILSwAXL2xfdEYgmLTO7whpCgj4mFtZIdT0FrnePZscMa2gey0hufMutJPWcmJjx8
Lo3DFU11l2RZfPGTCVxBbZxRlqixPQVzHwBUcg3hhpCwOhGV4FvXYk0W3VpD++o9
gAqFxAyO20iS2Gx93Cb5XDsry4IfzhKhh13XW9a2PwISzbCPJPpK03VIa2mHAdk3
0inZoE4vxe2Am9sW+1h4twI4KpGfRaO+6lrtxayEK7XSEFRq3CE2XCEG8Cbzzr+B
Xrh2FiEQYZgReBAlW3ZfascZQzxTqK3EM6plSxJKgrU/p69utGaEVP69xgl40ZET
R7GF09DohD39Zf+uOIVuNOZRXjUSYciR6ow00sZWPYMW9e8aaSlnkcTadk8hC6iF
jhODqMGThvqxolmW01yXAmuNC0K/MRDSKE96M1hxX4jiZfhj/PM/NvU54begrP5I
bP8854KLZydBr141ZACwaDjEKZvbL7M1NqNeAcTqc2v/3F7lUtAi4Rny5zYnvqNx
k9q2RwWuEVDOkW8L3bFlkKHdtm1ubRUyw7h2+on0GV132TnZpft73xc5c9042Y/g
pUXCHMwnGslHe2wYmcWv6pSt8LUEc3SJCC3joQeM2SEzE1YluYbrFP9/1YyUd3lL
+p6J8MENdncQiun6JYunsw==
`protect END_PROTECTED
