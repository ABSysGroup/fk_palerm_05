`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gmw2KUOMX8t4tTELNh8m/wy2NVF2CwcBlF7IhJ29oIceQWQGLpbYgc2GxbHV8Aui
LF8odf8p7Szh/kE6GCLFv86ifnqGb51V4BkFbVvOj88b+YvVhiadEbTPJtmA3mbQ
AakxB5mPc7Tz/5kNvOMLwxCVx0Kbi9SmKTpYqx12sBUdhk8OcpaycAwNqp6ZcfhP
nUPxIFKM0aRvyor7vVKayDEE2reuRsgmPkCSSwC3wQtvfxS/2M3YEkNWqD1TWtMk
Sak/3MRD4PrjLP9aNtHHGRSqzYuP22/RqWAMGHhgRZrFsUElnuY4y2visFpA345A
V7UIVamTwL/+HshPgyTOm4TxejA8EZm4+ijBGJ6QNQBAorNvD98VNM+DaQCuwzuc
Hyl9sJUHEcvVvERJUtsYdo8sxlbvyYG3XsZ/j6bWKwItb40evURaKZ3Z19zamIYt
MVYNPBoW3QyT3KUn1LRQ8q8Vc3jVwh88MOo6RIdX5fVYkQvA2Cta84FagynBOJ2B
zoG4y81sNux32ghBpUnhqwWXBjzUQO1FDiQE06IKAtcmXvGu0gztI0dXtCQhGYa0
SMCyXysk51l8lc9NlEgmL4aBkS0X4xtxyp9YpSZbsfiqN/snvAQC929Id/Nir/zG
rvmkJfVfEIG26RlbVs9yt7IQxE9hEWKTiA9zX6ZUrkpGzHKERqogIFhhh4zguhl3
aiT/MRE7S5ZSrrvy9yMu1ENFkM3QsUufNwn2hYq4Zkkqj9eMfjKS18Vu4LlT4dJp
JauEgfXfUk3WRB1L0oaiGb65sqNz21HgPqqjHgWr4DC83VcsdA1Z3yvv5Spe9uvK
N5IObOz+wSQP+v2M8xNYHsB8DVGRvOzABBLD1SYK8QmxZHZUJBNyPLq4yGhrCBjr
A7VWvbOk8XzqWv1TpF5SlfYOW/R2PF4FG246dj/o3ZfWd9JMjf/y+ZdhofrGoWK3
2GcqiktrGGVza+nwGZDssIpdC3eLWjEygjXadPdlEFz3catORUd0bjQViLG81DY0
V4dKe/qveBsafv+QvXccyYDdykH50eci6xUNnbZU59YnCMwdfDCZZi1quAF0L9qE
feqATIQl+x9FlXqc755n/xA00Lh9rO2W4/JmjQUwd0VNDEdA3IWdkNbZs1BXnMHz
yEUz0OvyiswJe4bexFg3+XxF/pMv9ADJYNqAWiHNvAY3Xh1tmZSMFCNvgeFa0aXv
fLC1JDPU400fAMJ77DJujM2b3Pe7buw11WBxWQXGMWiqJlH0jLPTNDS0W+GS3pMX
IlvknGylcv+WM/gBiTDHtHUXG/3RVcl8xW5c4LxRpEVqGuIsGLD5oBHzMaKXSIAd
2NotPu1rQXu78bKM23CP2R3pTsw8gJQzzCptFrWCXXOjea4WexnoHBs0KcY+y+vv
JZjL9RMc8E+G0PvQb/f8uOVVYSj7EmoX5RkA6G8HljdG2EA7E1sU0UgaRfddzhke
FXs29cJqYlJ3CQpHEn9CT1JCeP9PjnAXdvYugNSmlmzhrK6odYS0uGz2LNylIjh7
Tt0+snqEINWOT3fp8pjM5zr3oSY0X2UycYgMZ2BwwlM=
`protect END_PROTECTED
