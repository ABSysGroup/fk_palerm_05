`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ptIrLZmY5CLhJXjKk0X18LRGXZrKA3IYvyNlX3zvIuyudFKqLdSp6O48dqICcpsm
uEx5xCWL6ZQKUdQRUoqjwlOl/57+anU8gq+oAg45qO/HbFj1U2RNQPa+liyOYCTH
qowLqgjY+4GKOpWRqBPhdmGOWov5FCjVmmGBiGd4XCzz0OvwQIoPzvkELNXyjn94
QuAiDAaYlNr9oyWHVZ8X2arrp9MAIgbf8rXjMN7JCwcwbvYMCSpOjTDeh2nvG+70
ZZHkbX25U7wydDe+elMMEdYZlgc6oT7oDpwGtAUuC7Y/3GdhZk8ZnwcUPY0snV8B
cZDIhx2v+EeSFnOft0WQjYgvTk8RHAl2xrb+VTz403CIl2y/2A2B+lVxOIb5zrMF
pA6+gTyLjgGV+81LOEhdLdDKn2GkEOzikv6ya5erxJWu9j7jb0OexcmlwFQEyGDY
8WaIDgpYutTv6WGhRIFKhjj7NLqTtxVKge+7ue8bA+s=
`protect END_PROTECTED
