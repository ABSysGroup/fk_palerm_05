`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B+ayo8PMFEMOJzzVz8Uj3zxSxQkhl6pGpM3IL6unYzDJsFzhSRxNZj8WNwKPD9Eu
WsO7qpZHTNcON/uiMIESoYUcOVPwLxR2wnOydyLCPHpY3q3DRhG2M21AboBgwiQC
Qg43VsKtv+2TwHMSgtTtipZceMlubWoMpfJkBGNpb3z1Zpzbwd+1eny07W5VsZlj
P2+HMEBkcF5f9E9j/6Q/13PO539cA89TPKkeX6IV5UI3Re8LtHErt54MkwSrE/7N
np1hFVy0yn+1xvPvaJw36zTPBSe6OdI/mG8vUIU1ZKyLrM8PXHcXcmk/1yW2ohbY
tvxgS0PxvTMltwaEXTHUPhO8DMG0HGgrRdprFDqImt1mLvVmookOC3qF3wivVftY
L9MFBN0eDalz9rE9j2Q+b6NCYXQvN1hcNoAaaGcLjYVFpbW+p8GDKfGNkq3eiSQR
YP5XTHwj9vS4H7c9qqdfHpbCjKDhQX0uHMNNzUQZdZc0wBArXd6/fmR7cLobyK3/
gWmX3R5bThVJQssMB6t44Cm4fDoDySy6Y/1cLNfFiCvysKLqkPRLbp4Cu+Htxq0H
oQegfwMKZkwJk80R9E8g/GmQ8M5o/l4PpPug9fFEzR3cIXgezSl+fam6ymOV0JkB
q6g9Dgu8WKU6B8osPPZ8LWZi3j+HfflCQxPnrra8//IxGiCw3bGpRuqMVnD5l/PY
OsXDnIHqwPBZWUAfCFovIjLpW6Dz/3PewTqZ/HwirpHlZtyxZLCZahIkp4vmzQNO
fTxARH8xcaEoUMTfPtzfyq/kbXEXsdKG/lYH5viTDrpUqPX1iNIkc5sgpgqU+J8+
nv5U/aM9jOLpsppkoktvu0gnExlEDEZLxMPgAfabZKC1kZjB4C5kkTUCQnpElY/r
NPfqvFMRyuIYO0mwbcDupWBleosPETKwJJAXdSrRydf7Txh9+GWAYc+XIgiLzwwJ
97CuDviA9yq7Z2e8snftOcGhhe4EFla1aIxKdOUG1kxRgtAiB+R9UDOzsBJBPMcb
LOdkUkxYdt+lAbt9hsBmxqrWOJ+G2uSpXq1ga98QKyzfAJIKjKoJgh32XK8TyCOa
KncAecBqreQRfT4gKR1xRv57E8AC4cSLg5OLW9/9DXX0Uma4WlCmjU3En3IDCMJg
EvzSDIvuEEvdLNHV9lV4+GSrs8B/uxU5aaNt/CgjAeo/bl5zd1z1QI/bDv0S1TZa
LWNIFqxUARG7YYPlUNzlLwBxdCEqgGCy7XeVCmcb1zhYVm12RWhZeLXc9030+m6u
T8rk8LBWCOJdm6XkWeRfyu2993rqSN2ED8V0FXFhj/B+r9eUngK/t0HJ7pkvvH6Z
rOXUU52clCCiLar4zAlT2XRBnF+QYHd/XsO93prYY6SbCa0SV0VF9lU3DA1ESyAy
H4A0hck8JVfxM9OiK2pLND5587GStRhZhXO2++a49bViqkZgsHChlHoAV+A5Inc1
5OmXkSNjo7HiZxibaKA5w8dtyKlmjYPg5UhbaOBufFA0yyvrqjPSgWbdhKGpFbwy
lyd2mZJM82nmS3mtNFVSkIiKNWsyeu2cTlV8Hv0r7xiRQbIEFRPoazWAUmRwheNB
5vKZL95H+h+2RozY6KVtRRItP3G9gVp5FRGospOB5nlhzL1LOB3ZYfroFlnCR1jJ
W7K4fn2UWRb35TxtHDGSFSscuNWYJ30a6Dey4YY++b+J7p/AR3V/rdqJf/p3n7rp
w8iVeQweQZv53bW9g6BdV3ecto6qFPfAtYNFnKUedswTLqIT7D5hrJDMheWwp/dR
pUuqxr8PRHKqCWKzqrEA1peYgYrxnqfm5OSijmAf3+EljE3jrhb2jIErQUlGNPQt
7NDfk9ep09EevQKtMuGheY1N17H4sP1PKVH7ZQvY1PSNOVKMP3vog8zmnCUEWJlY
IN5jHEHx3kt01i02+2UMzSvmcTsxXBlCn3L1qzJs3yKbzNgu+oHn6v2HxWyKUB1L
YcD520deypRLJBdxNAUunTR0rS5x4gvjDMH7HUxF7lU0FSytLQ0eM4wmGkEL1CgX
TDr3mhsV8GMq4HmCWagl3yZCw4HUM6X8phxHnk+ac85R8nO1b0GxGGEVuMW5/Yl/
REOpkK1zuWrh2gTZ5kIaT6MO1kJkd6v1BdXFkWDrnuQz7Cu773K22plLYBabfYET
nffUmeN8FNoisbOJFXtEwhPKS1wxj8QMVJ3cX93gBzIvSRfdWlygz7cK0hpEpfzv
5ODf6xrmhpFYgM+/aN9HvXaPYUqmJB3WKheTUIQ45Z9O3xL56mUQCZTy6gbGjCcQ
xSGJ461KYhM91mhtuOWumkTwvJbx2mHo2QyHUJGGq4HaAzNrx/UqbNCaProLsDhK
Te8yD3Htn9ME7holSrDIj8glHLWehJx+POSVW53UjLarfzYR3rewJ8Wkbic07R3k
Ufe1y26HyGY/6vFStHHjfLwuWl4x8TTWW7mq1zcsu7kAJTi8SXGdyNxMA/n3TK0h
k2/xNR/2qmAKQ5khvAVKYFWr6zCY5DECvNuOFgM1XIr4rGq/NG+I3J8eDPqLTXfj
RjYGGGyYn/dHzNEl+k/wpnoMKWv6zMucTwZKlyNQfjseK1HdBir9YYM5pVW2N+jq
oyPBpAnrvQZ8tsx2wqxZf6HML1z5vcwlZixahfMnqMi+uY8ViwfbFP3NIcnAJOpg
v/qgSI8TUVHkHyW+Ek6VE2IgzqqaxyS5DUR9oAB1MPpof63PV6K1ypqLgXAeU951
Y+/f7LCjquCr6fdfD7lUKCGNQEv+HPHKGnILdDg1uEJm9RylJUAputwnzAR4GUNo
GS2op3iocz8x1ifnezftwMB9xNFIytAGxVUqJBrtTSlzJxe+0zEWpm4QmLu6Rx3I
2HSPUh8UaQwF8FR0NaoY2hSwh+J1DbaOP9xhA9X2EAVTVZMDmU5PwgYNUF+BWeZC
3JevlsuQ5kc6FGCNsd7oK6/oXuXNJ6VYNFPJovHs5SpHRF6/R88YkJ2UkQ1NTZCQ
LO137PsMeborAfHcj+RTKsF1Hx7HziEsMpAJtc0EQE2OFJdT07WmzogV6D+5qH+A
Xfs7Q9OxsnqcENOFFix6VtCriFoZLYSNbQcfj/wFSfABVkbY9K77xSvKiflD74+E
CHOgJ5UJqzrUnKJDPqjZd9Hy0xOWHl+ni8gbi/Oyety5vW6/sgcdnHBlieuMPqwO
PL4T4E+ARcEaGTRhiROjuU93y6EENk5gTqBZf6WiqdebWuE37+QWb+llGJDZzNgZ
W9kuCzHJoBtyNCLV5WqXukrUd9eY02uroTGcPsvDoPIzKKyFNBrrkU5VJYczQ0R8
V25PzFxj9vsGbyPYzdJWPdfLaYwOL0c6ALlQRQebioNnS7JJCOgVSW9eRdAYK9gR
FbjdAP7BHOn3xpadfgmLRSw79x3xKslLSahZvOjdfyho/BRv3xTdtSkzyuUo1RpS
iFqk/GdCaz1IOPFnL7Wmi8VWV0MJ5UhIGJ2hkV69xU/SNX1QPqq5UesbXHx9dUbq
/fIRQdD2/YEIgf7JRvVy1bmNwOPL7WpGzW4sPpU3cgncB7iWO+pDhQiqYoEoz8Sy
SS01ROCW45e6dCU2eRorQfT5XjgUtv0R51IlJsFA0ERI/hn/zoZiVXH51vqAB6nT
RW4zgqTnXHBUnnTOeebATTFIC9otQgYEg/AZ4RvdPYXD3Qi1Qtc5c4iKNazRo+Gq
E0nOkesuMhgs96+ZthC/BrioBqnWAGiotHtNczvJk79j1fSMmJB5PpeFskVBpiB9
K9kTHrwiJ0Hfrm6t129Fc24KGH4bHHArXxF1cymoe+q8o2CaFRhpGdL+UWf0q4mn
QHGAZWzPlkXj4idZhD9k4iiCbebEzdjhsxPVHbH2a+auNbrngh2AuyKbbTjuD+2x
MyH+sChW0Jrlp2jdN02Ly9Dp+5u6cTd8LZ9+nnZ8UPpivXG8P+1Hy6lIDVbpqYQU
flUGS61gqKmXs2nYJQn1uRgOk1su5ihJF0LqNPyPXN1dvrIeVNJ0Uye7/4MQHX4n
ktHMLL9kXBFY5XPgDR7fJ8FZ3KPYi5v5RGzfPUc4XGkdHMHEAIckm6X4dhysQTrA
PGdFZqmSn1Oq+ASd1h00OJTRYyWkgKYxoQLd+PW7oOp28VM/nJZ2cYoIqfPoPl46
WuvxbkE79U9HC/sH8n0kJhNUgAsP1gr6ePErzrtoO0SK3Apng1vKbKfvm107FmYW
6X/Q6ptzuuh0YIl0wijfjLVKvKetX+61wjB50hE2Y6nPd8yQQ21DSar2WZ46O278
dizTaB3U/8WKqwjj9MCF9nSBRijNlav0M3V2vnLdsICFeqI5hTpLf/40++kFsTYi
4tZ1Cl0CKvHcPs9FfLYDyhhl1kH7s7XW0vPhQoAdFGPtF8zYQa6WPzWli4P+U4CP
W791pyegVgiQxFMEtg2h6JtEYpVYIXb6qGOFiR0UMOsSCAevdDUcm72+g7MKfsQG
qvSgds01p588ywMAKkrjCXziCz844CT1xeE8zGh59loYRmGB7hR/EA78DSiP62CM
M3sRZxV7T+l56sfL1//6kVgXQbEbKtdk95il02AXz3RY0pk4pjlvRAqk6CMl3/eQ
nRTCCYN+SC499cucwS9WLOdoj4ckwBGC++NSqPb9Ztkg20uSbsXCR991gHGRzUb/
GKDswtNkDXSn3TC7qPoqiaVO6GD7uleVeGOGpyQWF738iPcxJK0aqX1PHhfWHf/N
EYVIlR/qQzUNIV+ZIIqDDdYj8LjCz77ToDPylKbntNZlY8TMxBFfCy+ZcoREvRB1
ArSbfgiGWsEsHEk6nPJfBkaa2xXcwetpJhakjH+iLoRg4gmb85pvWW/M0CjwkPNA
ASULsLZg9cUTdkZeY8STa4vQ7q63HxMWkcis61zBmdN66KwqbgtLNn8sEhf43XFo
nIXt/Tlv5LNelCgH40cDqKOnmzboK/OJ1beoeo6CGDmt2YMB9MlbZIHM4Z4Ub5J1
+LRC8YumFDoTB8Cblsiwc51oi8JNZDsLgQDQnLqfjowqQ2m2UsK07EwWjzj/mECG
mxHJb9nqglF+1eOzPK9EBMpw4I3OOvcbyOth7W/4V0wmItDo9axZReQrtK46lApG
XYvtlwiwsm3ifn2HTwxkJy4u+XBMaOZQVUR/oFDFw2781wdnuFue9RY9NxziqlYC
J1APMbCxaV4/aZaOg5Tl75zTAyP270Iga6y/7V7eRerKepXSnHpQZ0ppHjVcW5oW
21obc4lIty6n44TWBiFvuYakUNpQYZ+jHhDHmm8JNB9z7jAPhiM9P6oupuV+Ujfw
07y2iBNMRtQpp5QQSHuHAQktWOcBxQIGrbAvIZ7WN9ErybHa9A+3OVuie0DQkAMQ
zgGh6fptpXk4kHAKYoi10STlVm3xR9Quh1TWqiO0qYeVuxAcifagSf2Jj6xtltTn
XX/EOwjW+Y1hl5s7w59/nT1q8GD/9FBxAgj7Tfni/xVUgfeRoUf+WLXw4YMz+ncP
wGlGuCsRxcrSvP7Lk3iPedbLCKXuBxkXhgg5eoMTgJhhcWEFCXbceGDoPgQDN9CF
20sQkFVpC8McIQGRa3Dci4f0dUytP9afa0TXRGuOvSvdEaOKqjmQGVPkIT3qDb2U
o455kzlW9fGZe/V5WawZu/p0Bre0+dvG1t+/oFJBgp+RqQ1iya/VhNAzwwbI/GGa
WsLuFrFSRIC7JI68klR+AqIAp8+HCgmo2ttN/kFQzCVl9dX3u0yesEVJx0AKzxhw
WLjYc5E8wB3gDnprIxKHUWIajk9TFmlhLj067po9KnfzJdTYrSNJofnHGttO3/bh
di/pT+Em/U5IdlM1t/ehbCMucCKfkq+6mRVZrX3Dt5aYaJuMxzWewPbZVl8785Hh
MMy0YHA0Tdtk8WsfD6cQ1ReHlMhnVZLtaH6J1oNIp2L3RHJbkqjpl+IXdQ3nftlT
aVkxjVkq/TEjxae8Z3qpxB8otuD1xHv6cEgNQPbwLNAQ8ErsuFrk+SUF2KmKymgW
AIFuxxj3eFWxuDYjruSuWTcUAPCxEYNfUHOGHzrP+nzI9ynimDX89Zhjoz5mDAG2
f2iJZHMTXp7o05FQnynfmz3TIib9cvwPmkrC7BbHcX9G/RnyOTbRzYObRWfWP6SA
5JFIATB6TfM6dD1THueD2cp4L5ce40Q6UCrBS6FPYxDTcitObNDE2pOTf7/DrHZp
d5GOG2fnhXO8jw4j13bQoZ2flYeG6+kYem5AGVAsrAw++8/cit7anNmWcxDemJ+9
Up29Gjf7sYYWSche6Z9LSr3mioMYkMSffgtDfrCBwv/jnPuHoJFqYNnfLF9oHG19
bsPo6jfRlz5aoFpujKo/HLOWmDuO/rPSIhgeHx5PCdeSPfLJBeFaBwUqo1fRPfo8
Umpj0V2/AmuZWaqZrVQu+xYyFRjgvexSredZ1HP0L89o1tiUSHUgdRwxuROcKT+X
9C7csmtzWAyhliZvcNgXjtKBBx3MuJXBDuyeA4cBvnvlme3ekPfTDpVhWE8UDTHQ
JNGEt3o6OR9sm8GF43dm51i6TPed2y6x4wmAJMRsrF/L8rMeRCSJ29PZSPp5Xd8w
Lb19etnMf3Bi388qLuwDogUKVJXr4iYCq3C8G7BhXH41aheHYzapwds3mZuhryA1
yz2Xtt062dtPDeO6GiBL/uV/cwgKGcSBciOCahdMCa0qyuscaOXgoEX8A4JYjk0B
D4n7hWvROHME1bXhft2yRu54tAOExN8LeaJ50sJAIgMEitAodqOIvvNjYwCluapA
sdZutgd5xXhxzYrDUdFVB+xkYjQo803sFvHL6wMqHplHvcHhuESAdlqawEQiq/tS
eAZt6kLIe4rqnRkliLl3inmeLjX69QOBWKgHo4fHwCfuP/qqMhXY2OhljNFSymNR
8ARsFZLprXaxqFsDhjbQum8Tcl9HahbpdgMV8L4M5kJBMZOUubm7acwm0LsQQCxR
2Jjj5CoOF8LP8zsJlOUQk5HpBDGXX5aFpaDus9eAHCH5DvusTEoeSkfri/Aq1llF
RN4VTe7d46m7DIIsL6MYToQH2tgWmn7MmK3Dhv1DDsHB4DQ6RsTWc+6V/gbQExVx
1gXpps+LtQ7a1jmdvWYoYNy6MlufG8sjv3JJUWLrU+zaXP7bwhL72TtLQBJLy/wP
k+Ev9McepVwugmrOU6ZCX6BC8mUE3IdBhbtl8s6R9+MzZE/hG5bu4ySOCVJQFKSy
KVAgdcXqXzJ6vTlBuSejcoPBxfxkfrSGdMz57AylsC4cBg4l1ZzLfrlG8JNZZbup
pNF47G07VUYj2nFknR/08V/BraLPhEkTD04VXhy0qblWmIUZ5Uj2URfP4DvH7BmK
IbH9NR/ztSHmzmZ7BRmUB9vJDtVkLhcmUC1QTcMSM4txgWa9EbD9vvJB7e0OVErI
2/VmmTRU787ARDWJuCtpUAfTOR5NS3htbQF7bbckgbOMK2DJIuh0PjiGqmS9Fz5n
7UwG5vq3FxVgroPO6pxWEaVfncGyrxEzR9lzCAPT3UpRqW2rCDPJAxpqus6jkhoH
Sjej22+zv/STWh4dHdLcrPsSH8vfAueaZiVm+Yr/aaUyhXlLzj/OGgJOD9hJ1o6T
AQqlVA5uBrAEIXoP/PgEbclcoxF9eNPmb7frHU+fDaW+ZPsubf+bKerHJPuMgYwR
wPTVzJ71en3tuYVQ3iMRSFe/EPSFGplg4YYBkfEgHYHVmAEtA7JSf77n1kDDqOut
OusWNUzRoJIZ1jsUiWtJr1O0xgdc8UcVIpDmOjkXa9/HJTiQg63WtjnbMXeDLaui
GhVIBLO3P3L24vNi8sa9kZY2laQDUVSxE/PuyImERve2WRfdRLP3UdScTvHbsKeu
VFx+RF5IW278UJ/xKnEQKfiKhBKE1B0tsHrPGxDPOTSgp+2lmnrBvBN5+ALOdJ8C
YOVrsWRlwMWlhMYleumNVq4G51u+OfpzNuF1fNAL3HUbPrjK5Ckp0r1XsdlsYw7U
ojO3sPwbe48CHgVOBp2Gp3HibZk3FVTXvNr6dcxd5axamryZnW7+3UjMqTqDRbgm
sqEyGwXOJ0NLMy0S/6VA+FHlCPr7yIDJt8ZgjrF3xq7qYMa8GB2s16L4fpiI16U/
yqg0bI3wpko7Y6KlWeoqzPDpjBqfu4M5M/lhCDidecbE/2199Dc0fABuU2V89u18
jmr2w7ZV+Ew+ML/DsML4xcOAE1YOdMLfmz220HevS1AWqJg6QTI7ktK+2g5P5Qxw
5mW7lJ5nQySrSRZUYvZulIZUcgNbL2SvtjJHibSC3TLWFSCWWOCMgxtuNcwX1yJv
lALxnbLG/HqpfjWw8cq+z6NEm44cvu/QQir0Uu1nHI9sfe+HrFhxn7oueqTw7r4S
KzBkTNYM/sluVRBX7b9feJ27tOlYdzONPQOqyyPAsEUFHNs5GiUwbM7nxDyh0gnl
+Z/jMB3sFRoBJkD9m280iy3R+5erlR7gxRKYZFU1s4B53hfuvtHGIPcajCAUMooG
GiMWU7dljCSvR3JyqZaP5J3Rk1HGBEkduM4U8v1hwkUh8aYHowFvN6d6cUvsCbJD
3XrqtR/kul5pZ4QydFHKgsMeYhE4PGQKp1oY6T0UO9/ALCRzjc/mo99qOlSc3x7Y
YRxzEJYn3+td6g4S+ctmYswnF2MsclsRgJc/eT9ZLcdJvu+O3JjOw1BMFN8WBKjW
Dr+3hv/0VXF45G+9kkIUte9YIhSATZG79j/zWgBXtR9USVSMNqs2WuDbrH6+2jCU
Z4K4hLkQupWQSDQ9l53ZMcIcgTI1EhyfE0bOWM9SsbIoOD+k/mNekTDTR90ENvbA
gnwhalY4xb5RKy4/jZwNwbYVL7O5227+R4ebzXfh1N6Q+y9eOzxKh+DYgfomKb1k
i1ymmlXcgaQNhw8Na6S8YaP+sPsH6dJkdecYmjYgRh+bKjMpnJrFiVjGG1vmwvCi
WrtE8YSCR4pg2dq7qthtBfJ+zHFBI4fYMqt92BnKgW2AVJaYAd11R90ngiIkf+9H
zjcjfe1pMc2X+wKlgKE5C4bqUDSgNEuClLnapXHsFft/4Y39W6RFY/EDjjOCNh5q
gA/wfSFVBf9H9lM/4uUW8fZQH2Zlk/ctwgA/WRRxSYD2wpk5otRLfXv842qpqt52
wX4ceATpH6LTXg55fwNb56BRBbuwBEi4kmn5GrVBwSZlKst1T1PmgIcEHQi4CF7k
KRyda5x5pgDY4GUV8gSNY0Fh8QYjH3PEGS1g0WJuIu88OO9Rqw0CxBeVCP48DOwN
JHOOUXC4y/Ez2yu0r10P2zq5vCRVM14ARA4YdRwOyYzHIozfR52eUanFd+/bJ3J0
/coDhN4iysVJnqB7Xva4BfS+K4mleHYrSs7KDJQPYsjm5optgoMdQ9P75/nJZbgF
iG7z+i5Jn0Bj629nXVfi43RY++yh7DWBpbCamHw0/X4fKt6jwrNR82kFYc9UlA+m
gI8BDvWvYmJNohmo7DQfBwxqsr44HYIrb2gq8t+GmiOEvbbnx6gSi6RUJXJ7bJh1
mkAak8kkCVQabV5VdqejhJ0iCUXqzSmCmRusz0K69+ZBkNfJ0p4tTAg6QTt21nBU
xDIRqWnauRz2VOOsG4RhRiodFbXN1CcZNEshz6kodi0bi81itmjfNAbGd9qjUFxG
xfMlnjlLTp1vyV2P7wW3RtDuErVwIEvVhJ/9efUoXGycZOA1tmkpbksgQsiWIlel
WIxt8r+fBzHP9PYeNbEqUiOHLmdeENraxaQEM8t/ZuOWxGJXvT5ujdvzIvAyhFTb
5ASGJe5VaaYHUwrWOfNl2XdTaaZstu+j1TmGB0Qnl3q/45HYv6BgFl+skruZKizT
uIM0eu8tg9XDu/IClE1wMfwuI1ndI+bkQYefWLx1V5aRmg1iHBJTwx/HNQi0XvfL
A7j3RKFW/zQMweF1L8iz60jRsf5kvn6rf6CWaFaGB3xrh60dpEMRj5FT/2LKn3m/
Xus538HkqA8daLaxln1IrHBakbZi6Y2ZRFizMQEnxpKxTsmNa0f9XpYGZab+3GdW
ALachVkwlj1wT4xwApVtZhOvag0b0lXZFo/wsAyGteJ7erPPHfPIv3uZxKAc85Fo
OMzD8rda7eopalNtCa7LI/EICUQMPs2oH7zCnK/TQibflo85bn1lBuPGvHvNxHln
264WEVmxINPI++S27Sac9EdRYqvlNmll19nW4azkpx2xm7hYrl+4DM1fchrJZNHB
AoIMTpSWzmOXDg6A4WkjJYu7UtrsKvXy14jDGrxalFwn9Ffo/0NH5YSlDs7Ag+FX
IOcrXV+5UovnhLyqGZ6sDPOHH0cuSajDviOsEL+878PqPy8AtlYo2ulX0b02kcrp
9H4Pp44pGXY3KF2byiz6oNk5iH1lHsxzVerRD4NIwLZAItkmWcVPnyT7CiLWJ+dR
YlwWkP/5u3afOjVwC0ONKHzMWzUaA9MKvTtuWSXJ5cpDMzvHcinMxUlJrI1GmJtK
OIBh9WY8LWznoq0tk5CEHomNmoWineOz9Qn2yRCqNV2HgnpRvfXyM9X+ibb80wZA
POru0pBcU2x9rmDuJLKtJUjzxhHbAQlLl0PJdp4FUusbJy9lK7zRDpbjDRyBwaq8
+JXAOquqY3CUdklbF0c4ruqiIBqRQdmg0zjAqoZdQ/lKqDCTJdHZtdQ6dqRzozqj
2uHtVO9y8f9LVsXTqA2KhTL5Egzk7DBS/4WQvkApLq2r/UHxKNXpwod+WJlIr3qY
Pxy0xi5PQYyQGexSjnph6yqBI/CfJ2MYOMrGfBApPZq/pjdGNB4THHKeEFLFiioi
B9FRWR7Y1+z8qO2k9bmU5W4v80Rx+uY06LKx8CkL1dDmBse0h5/Ba/BHqxSaFCs3
f1nW5ioYuTdb1aVpv8u5eZJrTC+UC0TlYT4cyXfTjf5uDwdMOtM0Il7xWgRJhmxY
CbQSBfQwfglkzml7M6aQ2GAGsooHsDzBUTU+p4oJxvHKu3BlV9Z6xIUepNVGxORk
TNRS5QpzocGyyCHP0BR9nkEwMgoXzVlo1iii4TRnFcDNqIdlMoxOmfT7GqnPbJTC
QmIa0U2xrwccm0O5DPBstWNQCEkywAlROOMbLHFDoPojoje9B48NUROabagLb27d
J3HidGwy5Z6rLPLGBGe9Qgql0J23cvMzH4ZRhZ1UoXk5e/o2eQxPEXQvVJwkxIfX
dA/XoekYMqyKOaDJu3I8RsPc/S1kfrWlUcyDwBl2CJ8qCZrRqrIMMwiqIzKCHJXp
DYFLOnBP2KRAqEYBwc2maV4E926q3xde3vzwR05csMyXQRONeba2Cmc5labA26/2
JW40KOoU76gLT++Nld1NGod/yY7iuswfCrFPY7QZcRSExz2mhBKfTgWjZHLlNxRl
kcA7bAi6YiKg0ym6YfSRPLabMX8OzHrn4GsvyRX3OxDi9wRuZfKMPX9sLNKmHG/P
WK/Ynyw2mpI9vwljtbA26TafRQR/uKeb2jJrAos6sBs1JT5InGGdpVxYH8An4PC6
vBvsRXPP9AExr4lHi0MR31L3oZpA0GzXqcu35oAc8EAIdQu7sOYkgXyKAZWGtY5H
d/OsrQMpkQEcDBfjSVFCAAdmGEQPi7HWY8eEcQ6SqjLQQ8cAlV/LlLsI0+e638OO
GUMSxAm7/3ORJF0nMgaTNbkH3qhOJaCN2TkYgSrP7tSamYBdyZEW05CT/9bPQGDH
3Ysuc75j89CqT9mv6zv3cL1S6tZ870R3K6Q1HIQZ5Bf4IURgHzy44hBqDpqBgFye
whZckP1RHdxCAjS7THI+m93J4EQz+180oGrksIlBgE2C4dCMl0gjASg5KsiGa39h
08GrskxFWVgX4jA9e4k58iIPmsGuO5RoJM7MShkHm9gfy3kCGpgx37gBbHh5UzaU
Axzt2eP1ZScBbfO4rxX6iRNuTqH1BduKCca38+7D4PIv6cjBP/hsDfqD6k9e7qQn
eVvYt+Cknwy1Dxp86I2PQ600FXpPYcXgwSqdbrE4m4FH+mVzMpKTDRS3xI6NXKUk
CWSnAAMiepU4AfjNoG5PPzDkl05vrRqzpk35euFSdEjB3/lkKMn1CK+O3a0hoT/e
tRkZwS+1PvqKaPTIR4lOnfnzgY548ACotuZDA0dcyX/P64CdnqlTiIpWCMt28mv1
QDiqm3Qs/jPYbCeMSeSOqK58lX2d9AJaYBTdh4hd66vwRcLHBIJxjhY4rk3XS4Ln
dS5Q1ckOZBfO7R9/dVQM/vqciyCH9Es+lebKbozc5VmXYrPr4l+4kqGLNnMLPHr4
sqQbOLJOnT4t/Z7w8NlluJz0VVFnzwRnFL8rKkNeYapi9JYY9DSNCD450+vAsfwf
qzvrS5+UPGWuhjZB7QSOjEW2XJZkMPFv4lYtazlrPn1oWPrneBiDqbUszRzqEzBf
g5Tt+BiAd8+foEFnBLV5CozxzVtcpqaKfi6rO8YiUCvgDX/z9pwW4fTnlEbaJDVK
/+oAvTeTHzD8BojEYMTqV4Ryg4PrMmAy885q1MEBBkmQWv5uSYgQ4VZ4wT94H00H
sORhvQd8If7hMU93dSFGU0sXBVlRvis8jg99cmr7nzaAWPg2rWBQNFpm/5j85EHG
QYQ6zHSzijnesoGm36iNwlYNvWsoOH9YDlHjZouW8+PyPNGVboAT9fyAtmHx/V/c
uh8lnFJntlwnDcE1hZBJnwHcp4BX4NOWjrGzoWNUUCPJiSbRWQLee7xlXTQ3hATo
ffH4DCIS/xK8oy+WIdle8RuA4vV9ocy97YRazk5hVokqJWHcScykUtxJg3fttbpE
CgmSiO5KWRUuxAbeVKfjDWrPiyRjoHcDTmDRkCngJtR9KrYNsCL8EMxeNszM/RQ5
F8Q9xC4rPSdG2Jq4sx9wZqbA3KW7sglJxY32KkGyTbPvnylhCmX/p989BaTzyQ5S
aiq6zQ+AQlJZT63KYNYn8ckhOPKPixB4lJvbLlSCYyuFlp/vLajruS96RDmOzY5F
G8USWRaBd20Ryn5M5HCMapCk27puM14tfBXm/F1SoCUnmtIlYO7WrwLO0LJ6PR+N
1tDV+rGdcIZqP0IsMC51fSJAD15lv9LO97xNvBAjk+gFlJsfwWPPgmwVUwM68/Oc
voKBermM4vtDg3pnNsk9jgi25/tjmu3xWPbbv902C6SmnXWzGGJ734T0knBOQkye
iT0+ptAoPWiBC/LiYJaqvRODNbCldqbZS2Q67vR0HKi+ESNRn55qua8LBasDjHQC
FUMOnW+LO6fAzqlyLdj2ijKoBI0i/nwQkW1A4aPTDnk3zErUhiTAPfhcDBV3EeZ8
3cfGw5XzIG2+WSr2eico/keqTuGgcM1GTFESCbv6Te5xzvpwqmYeMLW5S7oZ1e2t
oYlHhNpmbWS4QxZgnotlNsnSEGQdsq8tNu3ybO8z3Rzmz9Ys/NYs40jwMx00KnVA
Pj9jTGvwrJdlrz0Oel+7cJg9DDsjvS9oy6vcE48ZV0u+S2lP79RfAidmRW0feZN7
e4jCWSU9eJTzC+gK3psYwTNpIHb+S1GLVjNLWCRmP02YUiQJlO78HlQrRoribk8R
8gV3z/c6rPoViX0bgJFZfFOVPmPdyYcGN5vjj03s2T+10J0+CW5licZ1IeO61if3
BTEmjPHSsatptN32vV3X/hKl+Dccuzi7C7eM+xH2/3/2O/mV335fx+n5wBJs7buV
HCkCHtQbnRDL+arX3a/xRY7C+j+r3mL0xBjjqWODr0h5HQNqswgn5nthDa5bAB3u
L8ZGSH2eom+eie0trxnZIvxdSVexnY5FMJJuEKtVSRePvYJZjJO96bhAqj2kn/RT
+y3NnBa0WWgKz/AnL6wqztlcN25gp9cc9RolxRotKBShgemzYXLetZ+YYE/aT4z0
KL8Px4MvxXAqZYc3Kpyv1Vnrb05V4JoKkCkAVu1WyDkFm+6L6CELxPbvBlW8J45C
/UUUIV1jtzs2MI5Kx6aXoLAoWbfHZHf8ZRQSDW2owRvR/n4NKO8uSBnzuFxawAd5
yJBkweBCc5fVl9hn75zzDuYI4LiGwj47hx3Wentdp69Tlm2qsWNGG6qdU0kkFvbU
jzuTkXXVVABFLh+RFQIVZCajRTmpQwfzu7yW2VnECdD1/zxdxFdt0gbHsEeeqq/n
EtYzKCm144HWZyWVnS96jEB1uLf+oDNSlX0RuzvCRTM+Pt8CFF3Aj360Cm4Lmj2l
Ci7uB5PHPlkr1ZY7G8jtWjcamX+hGxkK8wrZZcVWgZxJpH0uhhCl/YeVuw51tYfz
bypOBvDjAyO8JIDZj1/ttBZFLwWbIIBP/JEqPyaa1qVAc7G4CUxSKTYCQFXO3G9q
riSMhiGSK01vahUYBRHS9rFfgxXfdiEErC+3ParnLDWQNXPBtle3QoqPXb77yMKp
eMMpimxJcSrSvfTU8IhovAWXHSmXwkXz06aKXRHziqkh5pO8sT4MOGLNAZnY+3mu
xEEMCv0T6iZr7jGGAf4m9oQANnAapVeAmd5OiMS57wqUsZmZugkpKFfeArhw7Kf6
XMN0Xf2l00soiYQWilgvkjLpOQbZPnMtl2EIWefpzAl5Ov8rlkiYiU1HBk1E85TZ
tdoaXmf/xMqo+CbhiG2tchlzJZLba6AJF0j0fd5KAsd6VLVm4dN/uSAGRM4sD7vb
cC31lRXrvXxGNeFW+v/He90L3Wt9vp4bs9Z91QYPofGJB2Fmskz9lmWfIdyipALn
MLvc1TFlcA7Q/Tyymfj3xDLv4IPX7Vi+lA4dA1IouTOjQRRfbdLq8FPPWPCKwMzM
k9tGr1jyMisQJrpxkgxgDbPyGxkkyAQbPhlvHwTyZkUO3maWYCwdw41dmr+HJQRn
A6UEM5MGBqXlQqqgVye+NhxqcsYPJ743Y/2eUQYz725WG5KhVtUhue05y3MvwOTA
zlC6DHrJIhBNynJk9BkhhTdYw3rc+XRBofKFsJZwTMNWpaFTXkUgIkhlQJ8CcQ3O
STvPBQo25lS5ph3ugrtdHabYg26qec0vLw9HEXLk6l0rfgLTgFf89l71kpAPUF+0
P+4OpIHl/2E/BHghNUZIyIyufsFjgS1wz7Iwfq/eIpyBOIXUsH/ZJRvvjKm8WM99
AtRyFd1xsSRJTYjxZA635/FZM5RKaEJDSrHOzYn5Xe65aQuJVP8mC4nkmCChXC6u
EdSIGL1Z1lkTnR0D0esz2dMnAxZbLEo2VyZJGiUZqY8wbeB9o3Kw2vrnfxb58KJb
C32ZkeNm6xBMmjwbjTi9VIqs5dgHxiVUt12+r3gKMmOopJH0WRfJdzr7w7M70Cq/
kR3PSzwy+gYQbaSnR524Q+4qSQhDzQeffEeiqPdOAvaZ5OkbctDJMeWwgirSsxPI
M5wcXQ7E9IvRfuE/K8rfYo5/j/Yqg33Bwd/4Zm0pacu2Ta2wjcJKdS7G5Ysa/qzc
Z7bsCATq+Cgz75geHQxvdXzQGXdzJ6hlpxuGI+Mk41BI3sopg3ai4hp+J3Iq/AF8
2hOTjGHFntTuy5PMSA6iKTfBaTO0Ba6102H1OJDG1cBMXDrWj4p1b8FARqNNnjjz
X37f1AffY4DwPu6SRvTFZA4yWVhi9AYjcXjkAvLafPORRYqKTxSnA80g4kfxhK2e
`protect END_PROTECTED
