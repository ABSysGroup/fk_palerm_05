`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jVtVTPSlyIyjvp3zq0VXD7RTGa08OkajpTLSI1XGUzbF9+CC4qyyG/42FhRuBCbX
zA4HTVlhFwHCnRivVLyLzYTUL++x0vpq+rMXrMYbr81ehJKtt2glvsVC8EGRBU62
h+1OBqRMHgbGdM94ubtkn6sXiBJDCo7XSlb/rZj3FZLJYFIC7sXa0wOd/T2dcZ7I
H485NW0xzheEqcGbz+iQveHNaRRI49mh0+hktH5TT9Oq6R7anoIx5Ow5zQHMqAjX
pr7Ri+H8aTeJImVwXi1Yroo/rwEM7CfkyOLpcUCQGhphsTC4duCoHAusRbw9sRuU
lGaNJWGgrj41SvjYyAV+ZnwsllHflrHjy8QR6QojeI3qqPGy0odKAbDzwpo4Mdvl
Kds1bbZ9s8CY2tlK7sJlXH41rPL49xxrU4JkF1qtQWdF+hKvz4VRs43xMOg3vLl8
lYdkhFlj2yWimbEr75ijU+jt0zTk18KWUUh67qSv+V6FLbaA346MFVQCKwlSUh4C
aUWLQtxJCLvQsUuXOTCgD0xmy6Fg4xsffxNckiDDxScJeVlX3FXqBhYf3Hb4HZqJ
n5DTF7LvYutsXmOUPdG0lRJxs7igxJ4wK0077eOXl6hIVL001Vv3ijUxuEfuTNMd
rz7f9W2fh4MAjvEkDkwJt4ySp4U8OqKKdPDDycGA2UB0SMlN0qAX6WXXnwwl0T4i
uOURnJkgwTp2xaeeizuzAl7mfwW+vNVGg56FosQ/fhdcjZ4zBV4zKU0o10LzW/zF
LNuQWPKAYeePsoggrsSTfiYis65F5cQiXzO86W52ld+j1mMywZmS8UIygno1nuAT
597qZpeNEat8sCewErdnpwG0Lu9RZZSGat/3FwO2vL3Uq1CmSayWPSc9iOoAJLyg
E5AGidj9Jjxa5ZV2oEbGxrAnYi7vYV2a+Kudl0PfZHuKPi8Auga4vSM83Z3572Ne
oCIgnuesnIMwssba6TAKhb0OqbpfQs32bKUlrmXZ+j1NrQgizwbqIRhEID+U07By
N7AGJz/V4XqVagLV18smn9LPoGxIV+RR+IzVjuYn3M/pqQMIB6ChaumnICG8WF4p
hBuHH4k2djsVLcftlqLkn69GTsUBTT1wV90rYUH8042++3S5yWdKJprz3+5IcrY7
/9dfa/nlncSHwCyvOA3o5PTHERJmzyYJNxMaETzHEYPRGsQzp7nYoqkWbT4OP7je
eMbInZjEwab4RKa13YOJLJzeVpcAoinFqOmmqcEWM/uvlY2FBPK1dg90N8sXUExE
6Pe/kvAfcIf9P9Pn2Roz6vIuATFXneAAYVNSw8lxKcKqGRw1aqM8WmOGK14NC/34
UGu6kaLhcSST9RCP0vW3e2RH2dlzZDlZS54Fftapk/aTk1QLak9gktQPN6okJEv1
VpBpi31FjeeFb1apoN3NElwQJRamQ9S/dnwDL0nYMag9BZ3BSI0r+rKTRC/RvvMj
uWwxZswo76Ak9xG7fOjY1cvsAXwlCKIScsRGex/WNA8k885wOXDflqiMy/qS7lGY
s57w7/QTq4lEaaZMsR3HIDWNK3UtHHtX6zQdRJrRUCh5F6iKkMK1svkQ6kQYKH2a
rBdSZa27/mUqjI+FTyz2mIA589fi48MqMLs9uw9kEHHwflRxeJ5rB9zGUk2xabnC
uRYzrvDB3bcyl3noyjUlR0IRNJDbS9iKhYkWIuwL+BzAxzF+lh3sXovlYlO0UFs8
gxleNqYD5cJ2/bPSTc4gej0zaaOgtV+Kp1Go8unAJ+bSN2jyAjCKE+o2Muf41mo6
OrVnbohDvKZwoG4cNopiHw==
`protect END_PROTECTED
