`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IJ0wMAksm8Rzb+0Gkwdx3g+iD3L/lqSdj7DWAh82snzr63zfgWNucgOVxN3MJAEs
PmKfUoUr2KmNXtg9xv7lUjnLswJs2f7G78yo/IM9SuRMIMAVAHLIHYcxlwMkRFF3
VSbB8SJRFQoyTd4+zwBGSRjsWf4oC1vb8PTWZK8SOS5+X9PnlYefWHmnLGfgayNY
Z1kzKyV4g5mgFXV673VKjV2n2V11yEo4t1oRKConATw+6rQzGaZJcxQaCI4+0k88
73YcL3aF8smMcI466MNTRiu6yk3flVehB4z51V5H5cxdFyWiZbQMCnHNuw/p1fDV
kW/CK7Uv9In0HdKyZnuZghaosT9dZMe+fpdn6xclliwoDZryIuBaxmhnrTKLOK9n
4aNa7cYFd7xiDXPouZcBiVwaDOAyCHcNZ5qPZsXbxtL7Sl2uYXhEAIGAAPuPeZdD
4hZNhbj3c+IHDFuB/fDjs+1pAIiaB5Lx5EeFxtUyjNuyDBvBQaCXJ4XKHIFKRNW+
R8pmP6Zsvpy31CzfQS3zSFs15U3wXBvZRu3FTVXeVgWagfmfrjGoea5VMc+6tqqC
Acoh2/2Eu7YS8Zzuq/HL/GpmZteJwq69jyWFeEoG3S5s0CxtVlJV0B054rzxDRcv
hl9j/thuwDChmcRcPj556Qy3Gf//tjpFBfqXeM9MUElbHk9P2aMmbHco7mpRj84I
RRuH5z8+uESZCnkIANXTodEPAqnCiLFLz0IwzYRHCZn7N8vNegG+LHYLJPIcZ/cB
sK+VFhnwM1EBDVUK3kerOS9VlAr1bmchTb2ENs7fOOmNaZ0xOmjb7j8w/L1sa/TA
9VlIavrHHqFYgBZefDQvVfruX+jv4tVNvdo+iinoQqhsXGQQZibEuA4h2ZHQBrwc
GGfBM2m+Kgdll4Lx3k/GwJPP93xahko2Z31BZL6eGe0kGRpw96LC/pDXuiMlspMj
KIcpOqsORwXNlOuqWDbOX3amgpry4SXDyR4Ig6nuSlpM9mVbyamU0lsMX++Bl9dd
`protect END_PROTECTED
