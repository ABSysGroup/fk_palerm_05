`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DH59n/slcgG3SPK2XwmHQLAu0eALcgKJ+hFaoYPs/SJw6MNB2NZQ9ctzcVPKKvBb
bA5rx/A0Iiiu/CySAAeFuzU2E859xn26lrVbhcvDpA38T8I7SqFOjSvIv+bOpTSa
lZLT65GkfeLg8Pmk3kig9LPE4FJ306lL/7VZpTsT/03IsivL74zsPcGZSxSg8VNA
t501lvEudWHP26pjvvC9DD607zES3wuaSO5fuGsdZuJr2KGX0HyLOhYazJKTVELS
t72olhRjJ9O8o5rN4aJ1K3jXMiG2Fo9mrBUP+wHi0wuGv6lR0xgumJlT/WVwsjNe
daVaM4LzbmT0uWv5X4PBK4zx1h07S9AJroYxy2LtuyQ21EQ2OSmq4LgTQ6GutLjP
tGGJJfN+GziRQKTwOLiP1XDwQsCC0/B/T8T+6z4kJ9O1qEKRKMxCAYNBhWHNC9LS
HZdXfzmqFRLN++lhLX/7hcjbWWrcpV0yHFmkpQCQqvg4usHITp1kX/HHqfRMf7RT
wJL2BciJVdZgoM6TyQ/Coi4pGA7YuWmoGrDtOU/PU8DYCqSeSWM4HggdAAeitivp
YgI75VkIACw7TIpqiPQP6CgZoNODOYuak3Hd4V45Rx7SSYmr/TrVrLOemVqJ09RC
hDtCMBO5skZvvPWW09TJHihsQey9Upet0bmQv66y+E0Va/LasYXPA1KN697u+fsW
KBv9q6ZwwOAe54nYZgsswguP4TQX1mB90FZwDTj8enlX1nl6LsjegbEIqOu2FOUC
+2b+za2zSzCWvkIzhoeSP/F3gGQZq32FAVrJMJySZN7SCaZlZnSLg2vksY70wQRp
P1WzT3PkoJP1nuLF6yMtX9njo1nHNCCrK8GnbO748QlLSK83fHz0uQ1ov2NsALA7
ypxIloPskpc8s6LROlek2eP+1T9pPr4iAI7g167npEZdUlIwy5hUf1zWsJsfyD1f
wg/CE4RoqoXyqMRgEM2R3D0o7XcuM45kRODX4eyUXhjEr7XcdossNoTkzmFZAIEh
AFt6F6M0g2FhgfYyiVWpd8gPwyVRoZG3VUsJZ9IyYQePC5stFm/JyvYX1enlYp1q
wfqUdiLj4KUFNAdkll0b2NyNlBMAyGoPoASsNPUSdv5OxawwSBbYzccqu/gLqd67
A1ENvXFeg1sVILOsqYZGsVpJZfAllIyCFaFPe7JIt8Je+SmSrmIrWYyYqe1DPLkN
ZBabtA9TKkSZOGI8asaT0OmO/pdnTidLwZWwrZ07fUZctVOlJrsrM7l6TtcsBIxt
+SgL8uxtiGEeuQdWazodBBd5m9gZya7e4WAcq+lc7pQICeGdHvqhoWG3CJxB6GWt
ni5g/Zi+qiZQBK6xDpN0qO1BKdKNDTyd2KLvoP99yOFYFdlKILCjYqbdLWyYejda
z2dkPfkfga+Kft+IpdDa5mbWfx2gvkUjJAamAziopFFkfcQ5DHdtV1y49aXESNNS
0IPqgMnZ3dQ2N/HNPpdUeekeOw6dV1wPwtLPGExCxdjyBSCNPEAtuwqRpZX8M4AQ
QowjG351W2f8XwkCX4NMumJLKNMRPor6UX2LGfaQQI4vzrfm6Qz9n9ExBUj+PC7T
WzE4OZWbkwps8wc6/0m4n/FaTmDnkzkKCRyjTmZ6KMzjIJyF91Vklu07nwQqgLGv
QzBRGB1vuVNOHKFjbQKBVOnIQE06IjA7nWycVvB/+WDjNkKkfdWbJwn8NvH1q2k5
Pw9EJ1FZzqgO850oFItZGevmUx21xc1xbbcyWI8ipJFNVnLjku4Vx8M0mO644z3p
tQl12Hyv9YITgYfkTxcFgsxee+oJ1yC/FaElAjg/xFGyUrG/d2EeBLFfVBAQVJM3
IHojVu1KC3bcit2HkaqURB2N+6ERz/0n7zV3CZhGwSGuodHt222FC/R5iWOwGzD4
0xD2nFI6GQa2ftn9AYJEn3QSlAqrgRE5Rnb7hmaN7Zf/7yD1r6PRFE8CegKrVx8W
Den/LrxwcvaJNbyKkWAeO508c59KrVYlWjCM19L0XG2fugcOhT9oEqI/eutJdI69
`protect END_PROTECTED
