`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hYFiz97HY6Ulxyn/DPWvaE1Su+7Ndj9B9re/nTKTW4vD3phHMExnt4oJ4v/ouyvm
hzlyCcsaC1Im0LjdIzf0gg0XHoaaNfU6HX2mGNjjb2U7cI8xRRZzxlW+/Vo/h/ne
5dPOKrxEE1iekpnvkQ/xrpPuzricWVHrUVEqArBaVWRkEKbYa4vb2immsQEvjcyl
/LSloHRQ1MaLXMQFCF6/FOXyH5xso5f1x8RYy9owYvvTxBqR2Hj7bB4WYWUcAP+t
dg7zGuTXItm2t8l5xWDa4p8tLlvnurHer4/daOWC0ZjAxSfV1fG7J2ZT7K3z8Rk5
+qe5iujdk806E0q2zqeVTb3z7oh0wJHyCrVQyWthDUlIBZ1laSUZJ13St78YxZKr
xa/vQoT4Hgvbow5ikhcZFRvwxz4G7uXRY85m3/qM7NqIrg2sDt5CocQT4zgg7Uyw
0OKcnntqXqHNTu8LhTQ6+aALvZ5XNX9UGHfgudjsGfk84JtfH25D2O44ZNazzPLt
syddogJA8V3Wxj8sr0Nv9zYyLkUuMqnHhiU3hzGnVb6yoNJM5xDsxfxX0I8tlcYY
885Ogf7gSVczdCJsksYKDD1/0XlU0T4byZfbjTxtq+FoFzeNb19V979ZRIcF6DbD
SoFwSgNOxT6dZHvUcn/n+1ubbGZi7/gWydwpg9Z/5Drs5g0IvAxqD4FgDG71kBYb
`protect END_PROTECTED
