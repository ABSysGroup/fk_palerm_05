`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SVrVPVE4Kj2eLTOpOhdvzlb4DRTZyWrEZVQJ1MubHRAO1dk6aWSIsaZzUPq1r8GE
bth4sTnXifyTmTCOKmsf3OQiQp+nIdVb9WNHBgsJzxz+czl1Sn3iql3k6z45+skD
SlTHsfaM7SI1zWNCaNsZF8riOVsOJs8MiLu2tS2oZ0v/cyd/dF0FKSPDZOimjJZ/
Hx4tKpc1MuPFb50ybZDITwjD6P8SLIIx/mMRbEbsdhldgd0dx3zYKN0KvPfy5YQw
KPUdgkdbi6/vZOjpij5026YyBmebyRQ7kCqpo/TgCvVNK0KKN7gyfC3NZ6ec4B7P
jujox7VaWpByu5LdwG92Ko/ZJfr20jI8A+q6DTZPQAVlVF4mkGKo60YFMM8gOEFW
akMOEaIwJH8rZEk7auTb2BpjKv0cduDqgWQqLw3lMO75xQmhQC5pSbDwEnK+SHl2
baTJXpq0mmHpIrlDzC2Je65n9Q6Tv8N6wnUoSKml7hl10yuyr2G5C9LVOmb1Fymz
le/vBY+J9TOPB2qAQq1Qyq0jltmmQby9MfpDWnhrLASPSEbKzdAVkkPDaUhVKeor
95RDbPhz8eEhOnfAxYK7l9ZP8yYa8xcgolRiSQWcB6QHCvE+7VpaxTn50KNhWxzy
xUMNe6EjKXOGd/F6jM6V49J3N9GWnrxVa+97qUJXF6QPgTWoTJds1WTRY51uhl+g
oADmLD8CsqoIbh9Tispo8Fd042pMd6kIA2G4nJvRja2zZyq6jGx5w5/fzRdZHl6U
sWbGu6x+sn5v5RK+c6BXT4Jwj0NSCfMCpT44XCB7sIh28Sj1hwE4hKjMokrGgSu5
zGxTWdAUFEVu3e7A2jwtdMUriEPl2k/+K3r5LMABcj9Hg7jg4wFXw7//yAWYFtyD
TiWxwN9EVoGfkyyr90hG4IXd64mYo8NlElFhDHZXkri0qNnHHTOwhHl+Ot5c1H0k
5LisYt61edBs9ko6JEyDPRv92LgClizv2CCaa7i07gJcJLuvJAaEDoUCZhCjH6bY
zEe+daVK6Su1XiRkMFqW8gpkfJNrY4magahOTKYLBCObzcYkl4skoBfcwfZC1OI0
36unq0reRZHvj7Z+N8h3l1Ip3OepSbOUGVE72DQqpLQ/t/dCYFXMOb8UuT/7F/qo
tou8weonCPs0s/1tKvDL210wh9rLoBUw6udDx4KjRZ/mlAlT23+MyK38jg5eM/FQ
pb3/VdRWtBD34j1WcNmQqa7Bgy3WOqFEd+PDEvVyYsSPkFhrWWsn1o1FipSlyS/X
7krxBFKxw7bLNCF8BqSa4J1xq6ydBd2j/zL9YkE5OqQS2A4gyLHDSm/XidysTaP8
pa7WrT4173l994AtT5gvshfImw7v3X/qRahpfpMWXxuL63OK1HOd6FNTLfwKLHAN
bfMHW1Xnr8zH6e55aSIqZpyMOeo0D+sUCVJk6js28iAZvg0h+pPWFksP3qGz5r+j
iaTbJcFuqY9JzLRDMtyIw9uBw/62WegHDxxflYVQECA9XEra3hwRbsmn0BdMm4nR
ahG/ZWOH8SM/AT9e0vvH+DhqsHmIK8l+llyATd7q3LGj/YnKCvLBrJlfobWWVChq
plgOXBL2g3NfBnnq1eETgfaieOAQSHoKqOawBuEJywP8WAsFOm/uuB1psoTVRo6e
XreV8N6NhoITOifZY4oy4P0DTztW1IZi9ye+50U91lwgR345aRkmxa4AoZZQoYCk
brerQS6QT4PjnWDlQNSIFglrEc3BlKdPJreHB5nUbAPAvuxF9GNaDVEZkkBzrxep
X0FZSmmSu5UReAWdKGoS9EEZSROHreGykfIhK1HHJrG+pmMc36vpdYoNybXkGowT
ZikwkcNdsyKy9mievARGxXTnWmCj9h2BquDbR8FcJCdacYYwuuCQsj6k2YF6opHp
3/cX9cEmtEUUCmS05xdxvMbzdC7gMiylWm4LiDaA68XMX2BudPZae8ggsXDmidsx
2FJRavbjRfAqQIBOWFIV4mp4BS1v2NpP89an9yqDh6dmV2KeJDl2+WWu7frVepCF
fvYu/RnU/2VXfp0OGnUVwFIHtucNm4xnmTq6sCIGBRQIbQckMPwSkS0YiSrk66kL
zBlBmOH9GuNmef1miWf17CjyyU9WIdAlx+EqgXnU6ikM4nJ6wbSsBJCukgXZ3vpe
O/43YG8UV/sX6EpaxJSSETniaDF0DjPes2hr7mHAYlnoL7nGlLYqUg9JnIDznici
u8SJ5+B2LVrvlc25rAkCRGJNH5E1dZu2EUy0MRLXux4zstGdjUW1EzfHurBJKnc8
n8+sKLYNW2Bd3esdvcYgMV3rU7q4j6JpnhpmihGsWcDSis08cxsTyTNOFFmvnXbn
9dbWRVzYvkGMRHqdSBvOsvvzXQ7cJaU76ndP3zE/ypXbKMgqeZgcu2r+jnLyBN0+
BBgJQS/P3ZYdbzC4teKPeyJ1ResU2UaX/a0bOh9Yr6HN+PJiOX2cjnbBHNfpVwfY
hZUjANbS0Dx666juxs3xUBqLP5Tn/rcEYUovAH++Ck8PQcT8n8J36mVNCmLz7cmT
3Z//iECJiNZLI+u2kuH/JUQRjGi6C+nEnRsP+73oVCaTjCmQXzVF+xtXyfpn0jtR
nLqZkDQ2NPSrwUqEOVBOs5jvwGeAf2SSZmLK70Q5UhhzKB0YY+dOOPBzdLvLQIT2
yBAsUUD/5P40tJi4c7BuTf89kcmwWm4P/1wu3ZomIkZfVT2Uq3/BZoWfafgqY2we
a6abOsjoxCIQ58ZdlRpJUFX92z/4LfqLojo5Th1n2Q+wKKmoqqA04Imv2zh4gejR
MKd3KbMUPzZn3zEO1A3aXp+3NtvxnIQi56ZW0Jmyr9/NKK/HJI/7+QVvggRS4LZH
+MK3IHQd3QPgzEt7WxVBYbo6cltZGoCS9fuHNa/i9mgDl4gi/pWda7JB1Uhcz6qJ
wQqAkVz5RvbzvsYjx4GhVApHi4AsCboSLzqg9ssoHoQrSZaOKbwTOugr3Z0HUKs3
5PnTyKMPBLgUPJiacyMTXTahjljG9vnWcWcxpOPqths0YEPXU8dwC7FKM9Xl1AJa
vasNoDvXyPk8TH1NHN17UOXly+jztu81R9V1hM//AvucuCimzh51RHavXWYxjb//
E3zLMzZtk5J2AIsVBaRLuZvQUrQwnXFwoKWYxOSoEcat0gXVy9Vk9zImlgpDP7q/
kSHCewt8ZgzWmfT2xnLODfx/ezP64bPl6h3sO3IXUMTwHuGgiS7P4ni1hkODCQCO
ij+uUfuLl/a5KcrkcoVn5S6QD28ebujtn3syb5qdeSuY1UwQUOfpRLgHg+KbQ385
a3UI5o1XA289amcEk6DXTJEe+8riW1kpQKFTcwvOr0b+3BfKbzeVH09+KmwHrX+J
bEHTRO7JKF9emfKYHFnYdtmyPY/XLyJ49YNac4p8HcOSpsvm+Eb+zxxELALbX1vU
BfreCfpT1diG+rZRpS4ZDmd9XUUneb99/Waj68MI/6kYHN81+WQdZqjdWpXoSo5k
H7nJUfq9dE02bkFA/lLuAoLmJG7MJg4JF4+5gN18UgloOE/nzJ/huUXLQtTqDNab
LyF2kpHKdxvBC4no2pmeh1D3BUCIJuB9Ig0hmkppanWvpGPNEBeclq/GE8IwwtNS
2Y4dHkx1x/4PW6KvGYIisDatPUZProXTyc0kdz+NAc27d74GgivMTWzTEigwjsv2
F3/+vaeTYcUVlutZlq3e8C+kYgNqOgtUOw5R9EBlWQadltNv84Hnf5Hb/BTZS/0O
0OeXBRu0L2q5LVBv6F5MRvIUqNSy2uEZFlFaXM+k+LkVe9YlckLkElaTw4Y7Jjcr
aEh+QMukC2Sr3WUkFZy8bRZnbJM/MZVoygL1jespzkKKPz3OHu28Aeyg5LL1Q0cX
5vCNLZNGJ4N9+PPHQmb/nfbjrc3L4VgVWnKGj5jPaL9L16pdLUaljWUEXrh9j/e7
dFBfbyM1vKaQECVvyGnl+4nAjmaVKYy6L69tPmR5cSnb6NWVR4oFDHgWzVBDMzOS
QMro67x07PkpzUo3Q3vqpw/dsptv1D/JedQzLTW012lGKObIrOi8K6wXRXfapO3A
fjmZc/6/OzQC8xnuM033CQ3ZaUnKV+081XaEwJsDVmGd6pvVAkFNTqH114vGxZkO
yrUzHSjbg19FpjEx5Rx3vQuoe3ZEzjJnao3evbWrJ9TRH7EZtBVai3RqxfQesaOc
ZER9QzkahgHD5oolxofuVIJAjgGGsBwuWeeHO8Z9/z3nhNPrNqh7L4X7WHWq/mTJ
TA3bECdopXoKrO5MFzIdeFJR8FJxLfirGF/QO024jzcy91XwY4tWmBhg4gl2MsuS
Heo5u1OY7uZ+6PYzDtEpevfnCvoQql6Ch60Ik4RVk59ChipSA6UYfkCINTD5mWIe
TqJCrt52ZEAAk7gUd4fSAELbBBatfsNvvWTzgMzklnLA9WnE6FAnsue4tl7CfTqI
lc1GyHJPG8p8bZybt45CST1YrQy+IjPgmL4EHkYw+MA1mSTCn32zwe48GQg+zuUY
fFUF1uaZ/0HRv64Z5IUQwpATohKvZ04p1qGgTZCjoQ8PbGLLxeJt04ykdRh3uxxn
yMZ/EHQYTvPkM24L34ymDdJKlEWB1XOtFlBx8CDvp2XPu2BTRuJuyHB5LxQ6xWci
CTVMxj/AKn8F9UftGy/7vDJpXwOr23o6pBGftYAnTHVcYh5OJxSGY0s7eA2GFjyI
XaQEdrIIKYJQefiQfDiS31+lHW2VOOTBDPkPzsN8127/Pepn61QmBRWuDDy2jfWy
gQXV9SlVc+R+9Pn/63dCqHCxDBpjX+tgCejFrubpbR7BMT7MMKyXpzx0qU4TjqC8
jpT5m1jNlhPoj/LJ+z9reUaECS/DftNfbNtQTnqKH4hJr5+LWowxowis4/BQ40CH
zExx/gyBU8Fcmgzc74Pre1VsRI4juf/1yxY1HmC78eayBNRTaRLHencBp4CbcIm7
Sefq/KgMmvTje3oB7MjEStFmuc2KL1ZqCFtfx1chMczm5Sg6U0K/ZAQ+tSGx5SnY
wnaqvuX/7FWe9qeS0UL2yPY7GbIlZYMrvulX1KOcXAzV4dXUnE95feEcRphyVrgm
yfW/GjMeDC9/bFAGOFNjFdVAywqmiP8sBdXafTiy4D07KBjQB0Az0teJJU8WTNQa
XODJmz/Hf2THex7nJ6RU6kh0Fxz2WfGaHRMih5ZhLinDCPokpfW3epuDtEs9JWrg
bpGShwRVi95QPTwLHaCcBwNi9H1CoSRiSoNKW15Ls+PunoixRGtfmfr5o41vDW1h
IWQEvApwOGeTTs5mYJXRoK7Sz4JEhNZQrdUIYzbV4n9H4f5vnPEUf2dbS8Rl3zwP
MCbpWKOX/4bpxBWpKe3Q9tvLWgYodM/9d/8bFpI6jmdQZ/gxnRC0F1pKNB+87dHm
IVucsb9x/P3uwebWTtc+SCkW4TW6O8pE9Fr+whKYbZ9JBpRDxc24wlNn7WyLZUQo
J68sxQGoDxRj2VNX6KRLinJaAR2Wk6Smoqjp96Dl4p5I5Bw+BU7F1d/S8okr4QKh
uFri371S/1VxTA8iZsPfY9Pe0s8RyvDpleHeq7HUJHt02vPrcZVntzHFb04f2p0D
uHM70GNd9aaekpaecAzbgUMIK+SzFhGtaie4B4oP4xxV551I7iGaTnUf+DfzKoAb
Wh5iNjXOlN0i/34oNYYNF9LnZ7vR3nFyFiSvuc8T0fHJ7/XRHvi/q/Gke37mqD2r
kfEpvl9cJuOElkk8XTMlnUnpmlGJd1Pu7lJwCOVbzTZUSvUlscrdSpj/+jkNL73o
VW1VEz2Xn5XwnoAr+m03zXv+QbQvqoAa3rPuo6sx2VFa97vPfNKPt5JbOiTq7RaH
nEBpeZwoG4jpnMY/ZxEG4NWvLzcQVfbcxA6ggsTXrpxnPmkCDQ7ZZ24BtzoL8Alb
nm3KF1uvw8nyZHxZUyNfuhbUqFRjcND+GXGnymeqVRP1BehESiFzIOHIFNV2x5MV
aEbf7wRmzSTVP81dWqiRRy0iTZWE8Y6O/pzHW4YUKwBzIUwFEy6uoLoFUordv2xb
BFp0RE5FsY/0I6n+sv+4x7g0yjibVN+5Fwm5vJ4H1vTVOccHq7MxGmoGv+Lk3wh7
1uNiwFO9VVSLJnVLs26tXHu5tJ7ptygn8tj5woNd2wN1sj/WlgSXcKBfdBqChnxw
0qMqTvHcCNBM19sCgxPVzOcyj+afUbdCR1YXPEaGyEDJfFVQa888bmlXKeL+E+iq
Q6RJ/Sq3xYqGhty0A0E4pX1H7Y0ZB04ymMA0iXYdlyR1spPMzcXhzsa6UQNVQ6Jp
qO3TaEWl+Id4HRkegyiM7UPTC1cb6PjZ8FJZ4frQ6Uc9P8N+9XSssvo0Agn8cZu6
JeptDmV1TXtsC6Tt3VxH13K+Np6g8IeSKzHa9pCaUA0CqiqKwZTc6KHCBFHWdDLE
6qE0UzXhN50Fcx0svGjlquuEdQxoCI+yBAWBjWeiSDwbtBdeuou7xjIn4LQYVn7t
QoaFatrFsMSJdNpxLHkLx93FoueNHA6+2v/w6Ym6sfcsc5IlaLDCqcIJS7BTrePa
uNAdtjgIxLAb/8Jm0R8k+NE3phmlceDuG5M9Cchh0PRd5uIi0DG8meufvhB9k5wx
5kocZuP9luqVizoj7xtjUPY4GVFBtF9ji26KqdF2VCSGQpJ5dwAqAtpDKIeFZeP2
RqtdzzptdfFN8erdXLHArgmuhqoaR7SKhdNWh9CotvkagVxxlZ0tHRzo1p3VKQMC
6l2cZLwfR+clvksr7DsMs/SkfS6LpQIlCcTaMU/OnCQPn/6DwdU25kj9cFn9UFfy
PuB1QGT4oTSgFM4KBF7/W5QNDq1jlZqEf6bXSA1Qc8bu6gBiZB92r/nMWNzr1bPs
etEofVDPuHoPME7yqgjzOsHz7GKfgqTBqcZUZ/3W7PhDrdskG9THcSgKh2RW8T+W
mtuyLe2j8NYfpm88Jbxeg1662fJ3cxLaIIX3/PMw88huUYakVseBxcrVEMeV8s9+
8j3JZ/zgBp9GQzKDbLnbzUkwWNS/2qgUcUXbc19sNLBOy+2BI+iERV/zceZeWU70
6D1pOLP3utKcRSfY/mWKYqT8airRBDncqFISqgr8YNamxPz4mk8/z4sCspGf4aXy
seOp4NDgZ/fdYXfKsyysdCmQZw4hvPJevcJ8mmXu4lSmWjjeJgrgw8hOSAydItDw
TMYaVRUs5vm0H84bIiBXb+4p+95Fi7qE+DeXT3Bq9fx4ku9q4GRqMgURmoGoQAM8
AECNnMCOVvFYi6w8wNf+G91OkrewT5Z6QxGN7i/4u7AapmrRTh56k7zlZz13213w
vs9+JUqNw0kUKnNn+Vx2F0hmreagJLph8Eyw3lUwqy+HLUdtFRvWVXbX1aEBaO7W
70coFYzOaJSy2C4SzghvMWL6l4rZywK1nAj8K56Y5/OSO/7Xwapo9R2/lyh4CwE/
EwEO8dmKatzZWInrNz3SA9R5oyTmNl4ZzVViKDCUX45e4Mipr7qhhhw/Xs9iZQOC
+PqgmlS1EnuS3YlETv+vJOIQY33hsudd90EZImyRfGz0+GCviHsXeiHm0oopfiCA
tBhZ3L+wmT/EfOcpXCnDJHUcazcP8B3wRs1EQ4xMsAxHyfqVy25DiHW75wUdw5GF
3RTm+seIzz0lv/mdafEy9OiKg5B4j5LfGRTrqoYDf77VUVz9x64jX8TxQWbFwNwj
6hvaJKkXbMUG0yDMBRn+2y41hN6m5IG/5wL91tEEo91oVuIUg9JZgvKxC0kn9kK4
B7lwcDUZvt6ZJ7URanJnDX6z2dTNOAbH7d02ZWQmJKpjB2SpqveUjVvlw2a6QJ2Y
waVVzMY6POYLu0EEbi5f5zmpbLanYtfuppN2LzmML6wY+TXIO35rMzGGfuDa+bcn
bGPAuOBzA+aLxoZ3LsdcWeQ0V8RQ4Fd7N+OtKeqgzU/0CVu29iycI/zeDlbun2uK
OiuNkh7wHPpJYz6VZ1FnbdEmRE+1VBHc+bcLaU7SEjc0OOsjBCzdiek43EOVYwAO
lVrKzxFty0EEziBIySoakRGyNHUzyVnEAyPdztMk4Q1MWOGeL3vxBG63s6McOY3A
jkZTSMalBgvlR2/3GzyQV9jj/RX4FmtmDP/CZZH0arrnSL1UbQ7N375sFwQJYBek
j/710Y/dhbmkQYp+NPDL5YT1bRgJZMygAEPQa62HoZe6falprMyKzHSqld+0p/rB
Z40oElb8OpANsFpxw8EYBSOLjZAdKJbvE05XbAsxxPzkVJg5yZGRg7kELRVxWNxr
FIs2Zpu1Y2TH4Z0xZyJgH+oOw5S/qxmXrpXD9gOPzS9B8kVD5Vm3Bzji30OV3EJx
PVCNOAu5bpz49g9DNAP6Rd96GKFUpYDZRn8KGZ3fHLpmcASE7DlECnfJX+uccOaQ
7vmkDHZwF7sVTIk+kfef7lBdmiN5nkbJdbmrAUot8bqB93uG2UdEj2vOeVah4QsN
MyzVssf348VBcwiyMq8IjtHHVXJyAHYtHI3V3liZZeZP5huOD+xdIgEcuVkdFbG5
nw576VQWG7GIj6D4CZdozqT9ieLkO5quxJZHlrgODOtVp6ZZwCP3nxc371UJ6D+G
7g++D8jmN/qlR6dXmqjx+NDQ5G+PO38Y+/TVRJ9p0tfiNkcGuBGSQDNwfeJvrRTc
luhLKFbG3QKCcwDV7FjkU4DAMcAbz0NsVWcKmRH1yFnBn7d6FllwSwXFzZaK9fOj
luERu3BwknovPXA5c/3S2wcQkYuNIIG9Zy/5CCbHvtVeTx2IzPMItRJfVsSnNsRa
7ijtrnByLlgyWLbwSsQAXGOmdXL4GLt20KLcmikZ+NsFABU2II0EbhwzVSyGMY5f
dKIlwt3zUEmpIpPujY2AkCGLM5mIxkqRXUeyUxpqd/yMVgmAHWELf47MUujmOsLe
ySkBPMZJaJfw0ad9KltmgOfJhqpTwTHtdXquzfXcMqGFkCjiXYEUX+m5i6jSCTYd
sZR3KTKpkfDTAfLheABarq8mTv4+Uy+u/dlcEz7YEXgGaLH2q+F2yQ90kv1AhLbi
/PECfFtpNH2XYFS0y9rjQG5jIdZgBIC8thsyVXfYI3r0WGFB4aH34k860c2OpJCN
pwEA0gnn91D90ME9yQt33+5eecBAerOEMOishkQTJUmemu9+MJZGMJnoLRH11rAB
eiXVwCHRuIYS9NHTgQ2dOEHWsRLqXDBRpYxMDtb4BBOB83FB4OK/ygaDIl7cZLFq
lEoEmksIGnDCRzaqgL+m/ZQA+4Krf5qdEzTdBGJjY+bDxoZNovHFO0SkOuViI5E0
4BkiCGUexS0wDG483C+N78AmASVZ0Pz9UVr+4BKLchFqaVsramInjQOAlLnqC5t0
VWuyeH8BMHBP4dTIh0n7Ui1PtE4ao5tgfsY/xcveNyvvbWbe/2mvwvn6lr6nZndW
ZpTElmGHqQqnQIL/2zVsbaaWPNNHEbxle9pnjxYz6HIlUQCZFTMcvEtSqoXDJ8lI
QHuyw1pK25H1TgaN1vodZvbyEm1NFfUeebAguHj3i2JZxZeHCbLYRPJGhJnN420c
5gwoWkRmzDW+ixMyVBdcYlAZX2a5gSnbvVffnVzOVj6akdCRxZosT0MaT8qzkQS/
hAQMdtVljjOxrS08r2OZLfsEqGDnBXGtrk44H+bhWkj+7RP980JS9LwrA092BMd+
wRSSEUVA8kmjtJbR1lTTmgpykoaglBsDcFilYg93xo0qocfdkFZ15D4N7KwtogMX
p82fL8brAXMfnN9nemgSLAI2hu1zQn75ucqumdMrnqXazdpK3v+RzmJA37gPtNx+
DnwRyJQkYku1Reg3EO/i2Ti9xsqlszMFzhsntVM8PUsLbd8ATPGo6NFKMO/rffZm
Dx+efsX9sEn+dKyPbjQ2g33yUFBjLz4mDrwmNm+BIdgbMdiAPqPAfAaOKvlJ//gM
G9HGtz0hh68gM7Fegbah/OpQOmZcZ4/6jye1Jc4R/yW/vjRaHo7La1mw7fffgjb4
8MLD1YOh1TPbxk9NUXdnOqB5EMoQt8v7Rn7wtoTjy/IgJZ4Y/7+MreAn1GEKPXfN
VIw39J5ekM593tH9H9lLDl4m34V5iSNQyzfupSALBX4g8jAMqgjiPuJ2kaAkdCYe
ISxoMPh5QawkLccEemIgxGoVgVSEupm+6DoiBp+TexeEIS8qPfpGvOGB0isz4+Ee
II2QzqmVK1L5VV1qQYDUIZ9qQFppQN0q2dIBKCWET00NJsH/auW9dnzDhPOSkKDH
We4kEfLTdqfRRURMy/+W/ncC5FXwx+5h6vTyCIny+9LFZYuMuYrxyU3dOeZNoLWf
LvWCnNnkAdmRqSlTLPNdO5zRS0q5UBjQssIozig9LtM6iBTAp/C7m5BBsN+oAVdY
HCvkIMSaDg+eKYhgNUlGqsONCkHZx+pxbHV3eCYE7NMn4gL8/jXMJ8FT9NMLNiU5
LzK8opnVAYv+yvv5POEUDDfW4JaJ1S+pvaw/P9zc2sKMjgl6880nEbW/bG3AsJcx
FJHsgMjfDg+IkyEnyXL8PktNB3u9sEXJpNd/KOfF3X9vU4qaKE0D8W2abP3Vfupn
8F4H0991A1UTuDL62AqQL5650wx4ftXUtyE1v3ZApU184MVIIeT7HIaCPP8M6bvh
rBEpzzZJpiPLuoaDgQUBEC4xUEOfkasJ2ECXoGxr59PqgtqPA2xpGc0uUHa4qkeX
p5usK3TXIDKSfrwZRmK908iG2r3bsxp07MirEEjvwfRaFOGvS/nKRb+AJEKPqRmE
1WV2F+Y3ZcqmSNqFQ9jUNlCrtu0U59XNvJGuyAdqQd2mMZuTzend0GnI8bm7vaM1
BznfLch2igNB1UPG8IISvVb1TH0+YgAv9a+NE6XQYdza40QiEL4Rcxt+1/4ACCan
xehxuv6y9AZhSfptuBLO3eHGLxrDKf6hHVhTMfnRm+k59ofch/TcgN4WU9bIy93l
tnU/DVaEJIV0kFQl7AbTLG+OF40j7t6y0JSZrDakYyR0FGDCwD5Vt8FSt/DzZx3W
8Cp/jcRyNc0noz/kVc2a8AJcTgPQ+jVbT4yl8p/cucBWL6Cr/HA0i0Am7V0StXiH
rqFkFTC4RRnAvX+NvhNR+gYMvecv/PJjpB16uyAS3ftG7+jbviqvKFZi/41aPSVr
+VeHpYHIcoR9b9ccEm88tsKKJRFQtYW5YkArOB8wxG2s0F20bSHfBJOgehjMolIR
3ga8ozplfBlxF7DpDrnFpD981s9EwePs8TSV/YvFAu0t2p4WJB2ZOmMdT7ZRGeSd
0Ahm3yp9qd49cks3KVl4N1IaMu7AtQYB0IL8SBaYnEzj4I0IXm6F6H5YLseO/4rW
XchErC7qaxdv9S9I8n7a0bPvRTK0kDfNoOzIbweYgBRG1jgttAa0EQJ+UnPY9eRD
3ss5QWampeNBPoODADqMWzlad7syBHuc2Cv5o10dypKGvfWmCKjtxE35uUa8DPFI
ToH1NKcja0zCFjhS021esHybQqm1/ncfulgvLliK4ZG/n7UXdIiRUe6F1oW8ylv/
87fEMbnvrmDdQ9QqRCbvS6xnHzOTFVs5uUg3j+Adtfv1A1EuHOo3BrxKQZyFijnu
GQfR90egsmRDd7in7Nv6bYA3IUQDN7V6mwlkDTi45tnxDWRwhIuRyloFeeDhM/+K
Y7VTgV1mBqqj2LjdDNrgYwV9bIA8ehax9KsxA+15KbhtXTM5bQdhchwCMB/jx5i4
a39GQMdsq7BmzCFEPw/Ob+sdH1bHbMmZAScXG1DRPg+HXMesCuLF7fzfAY8EHEkd
k3dp59TennSa1zeWmQAxSdwh36cPh61ittbWzi6u1Tx+X1xkE6bqM8tC0ydYNWNX
c0VGKPR3lLR0zPyf3N9TMDyof+ykIEpwuWTnlGxTBYQoUaHP7cXEozNln/j0J4Lg
k7rrM+86YZTbaCOFABPzoxSjrAQfnZH/28HgYAthxiIeXtdx/+4VFbkibLjxZQ00
dkpwSXJxrPVQafuNQeGN9Zcy+h8paAgambvrV8uX1wvBn9NKgMdwjiqLu9zKeofg
KtAJyq6o3ELyn+D5XfMENNwYyXqW4QJLV1DOZj0nrcv0cV/45Udr/JO93gLuAc5S
0XJisNrIQHDXmdWPL6jZNRhPGIuBn2xWVXd0l5PO98f2zbErpKBD6GnuZbRtxtCT
8bW+PaRP4ENtzmRJa2P+Ue+3fkUjO2Uw1xw65SKs4lKuxGae5DueR5UamfSJ8JLY
mFXc9QcCeWBUClVkpnBYXQt+folIJPRa51cRLhVJwitHRf2jNbKo7sOEOYHOFH+N
M09lTpJecOXmISYQq/uIx9GiAFX00eX9rGXs4jFMvKriYFK9AX1MzwvdQsYOVNUU
TVIcmol1i0ZSus/4xZT2K5d6J4n1KU606KZWS6EIA8bMaWm2UPqiDTrpFR9bDOTn
VAUjSxA9RWaG6octfr3A1MOM5xDZOR34BHIvu/uyCHRka+oNuKjNj2iw38+cbt5p
D90q9uAlPMKqQGgIUzpfFaGusB2W8BudBiOKJWZKkYQY2eSOd0G5IxCv/4fsyxyB
J09xx8G8/r/RLtwk1RWacHld3LfsOQUiMUxa7FCTA1COBa5FAd6bm2ApcPrs6JUu
IlQqTFgP169KqSCQeDceXj//bygdsxFLpvx3uixYaWrDPDwRYe+rOWCAy9qtKqq8
RZWY2GWpdfIo75aFpxr+e6kdGxXk0Z4o26pX//Q7Q01bvs7XxohT7ej+6435/AdN
9ENTsdHyGKgPa/41ZvZXzQXPUC8MkvubxDLVxB+2z6Jg1S3MUHO6q0JlUb1dv0Z6
F1FUbUjWwdyB8JEVL1rEuebapnmlLRW6Of4zS+ZkAzpW+hfC5I9emWzv1aOWit/y
UTs/fuNiT0XACHyoqnW83nj+v3ffh/i0g13dxsIUfb/79d+oDTJ1dNNBc4CVnmsT
XNnl/kh3yLipTfLJHWumEfWdNr4+pmfL8zmSKmCiG27TbAlzCETvuqEm6JbRDYAT
Vwr8h5rfga2OOEVkxytNBU828RWWf3N9Kq1Q+djQlHBQYvDTRoskMOsoCL/lmZv+
xIfOyeoYZU5UXG71SvkjStGqT5NAkAgDfR7oY2dR6vLZY3oX7IPo3GHPD1+2pteK
UpZwCo1vau1DvaFsx8bgfCmXmngYsjHN+BVz3CbAoo9H0dOxC6pZ1tY9eeJHf/Mk
LL/xzKI2IfFlGwjXH2skRAXT09T934d50tvGsSUUTz7MQFlqCnBhRk16gqRNKsFh
M+9Ok4+nGxLUhgclmNJXqxARL+y/feW2Oyj1/Y4Ng6UOIF1ANpErBfUk50qyjinV
na8cRxvp5S3xTQrowies4se5PwRczGquGS9ZNUP6u/4bPaH0fU+SbBzKZrqffhQj
dvTGKIAdRg1MXZWisvpKI5nviZrrNiju3TaJOMJjJkH2k7NnDtQzVMwXKgf66M+v
OomBPgVZi0JR1IyOtro4b6M0X4Vt+QdbBhNrqRRKmobtxl7W9FsVytXq4X6EVA17
1H7HRhIFaZUawJBGKqs1cjo5Y6W+ZxPx0Psg5pg/IfU5lALAY9uDLHZR+kMrpff7
1qvFBtCgLu8p2zXvImKCvSmH065axCUacEtvnUZGYsgR7HNrsofsBV37R5exO5j5
AlYB5+uWG6nAqMqbAXWn8Sm66YuDgtXOTwg9Lrqhk+szVcwILq+dODUtWaEQQqbj
QctMlnUBOAj6hRduCnV60M4OTBy0Fg2s9zv1Y/mFnaMFNJasFPmWV0WgLWMYWdXF
YIp9j56VBilcFB3hhIwLXTQ3wc+uYDq551t7jR99oNHIzI+HARytaFBc1KTOxLji
A4gTHs3A/7cHyQqnbjRTpT4LaxEXmxTWTkcN/1uMlAhLkFAx5zg2XYflmoOifmos
QbBxmV3yaKb3V6k/JlVuSRKy794FElP8+NkwGwDl9IxNmHlm21Lf2bdBsYvDVTjA
lg2bFiN5IG5KfAK5c9ZBdMKry59qULBGl81UFRr6xZa0aKzvIPdVd7WqDlT18deX
skKVPDfEH2F9Bc7MknY1pLc5VI6IRYN+Es8DfSsJtFgzcivciWU0VRVnUFiTjXVS
teaW+mNlXVR1JCDnexvctSiLcGQRYcWsypsmkdZq2NE198oVQj+MGunc0S43OTkb
Pjxmv6KoCkBbprWBx+9XMv/Owubb+sJvql2jil/O8m4z2Eynx8ZjISVAMnNBkbUl
5v4lFKRj7h7xPbcxPkhYqo/2Y2CQXa2IRZUPrLIlee1M1O2DepJqBTdxtc1MxaqX
fzbuAaB3G6MOfUVu83HXjXN8mwu8ZjcWH1cZ9eSNx38g/L+E6I6XiSWWU93B9EQR
EClIsU1BYgYJyoldWLRVp5XrpODEza0RBXa7KpxYfhhzJn21m6ccbVzVX+PTVLFz
wnTUYFbe+T6wNZXw9AnNcOboy49KJeUjGIsl3sgDM4BKhHu60fWf9psmx38muIHX
EwuH3v/CU0Qi121rigYmHET+xhV0F8kiHBiH5g/a5MiqZ4cHQgnEIa8u6RJsXv5j
/8ngNB8E8mA7Mltgm2OkVoFZmq5omnjC6jIMDj0Vete0C4qf9F/ellbUofCdbFgH
nAmB9GdSbd85W81d2tM8LDo0ndBsJF8xQqNT7qpHmrqQlFQ02/5S2qHMDObD2f0N
GkPrqnR5H2vup510TQTjeMXNFFRRwaMZm/UToIJ+78R1cQ3cdQFa2WdeWmuc5U4k
zzRUOQjT4gDXJa13j6+Ku78TDg8TEAakIYBcpYKxnSNw/wtOu+nE61xta3LPjM+p
fdn0isvMd6uLDsirkxFu1YrEaB+AeEkPCTfnToMhPocVVlgZKnSjvlxQ6M2I2yTm
RNV4XWxzdQx6PNMpEMMuDmaPIcB0qio4eqaZrUw31c6MAn5GAThVNXMDQs2Y8Ge2
st10JyKtlYolLAtlBfCCvD3rdfVntWnkAoHCB0hBibQB07sm2Seu8q+FCfncKkZ6
ANFG2gV/OrsmbmU5x7oY5PzZU4V1wKWhbAd23eUMWq98r0mPTLaBfLi4JuF/EMfy
krdeSAWzB3ag/9F72/Nal6bZ13WiyBCRgx1txNVdkkL0VNr7rOv26LXuF6v/d31v
aVSp1H3ZJfcnwVUxcjWE6h9fDI+Tg6tP654jV3WPnluoB9wF2TLvq2h4aBcP62Ql
8EqecLXfAgwueytcvXD5TgWkrIXwS4VnWeOAGfaF2PPgMd8T6mtcCZyIEzN4mWId
/uNfqrYNYaV5ptrlv78U307K9eJElhyXs8y3PaY6ohBboZ3EXMuvhbRKx2keoV2q
T1p4+RsFSWRcI0/+1WBTNOWy3tC0syb+MTPB+V7tmXilG8z9lY1ssRqgr0Ij0Hs/
ziz3ehel5lyQ06h9uxH1JEWLnU5c17w5xD3f+DNEuHN+d5FOU91/9KoSGCBDRMpH
T58BYEJSHP/ZDWI8S+kdHeW4fdEYrBwv2czRJwj3zz4TPmaHrUbxVJk+769qLl3h
/7eoB8hM/qU2+HDzW0VSYPxPmj90MmtzU4dBHpjv4BrvM8Ua49ukFxHTsA7XrlIa
uQ1Mv0cpOgyRQPLRcEDVslhCPqmrJFQ457SUhaN4eicrwWa6c6KyXWsrM3DyiTZz
xFjQUpOzVF2GICOPdsJH+b0PQBZD6XDEPHpIvDHtu8gi7GcdYqA4iF+EYDSUp5Ws
1PQ8PgXLUPmG0V3la0/+ub2CVpye9obxkJZ5vFI2tETJlgRBVEhlMVTn4KirLa8t
sguFGuAXzONuy1+xn8yG7mcG2S5AY0IzMkeLmiAiOsz2gK19UN2hXtTcWLT+SJN+
Ul8+Co3yCNGouX1dfN4P9ngdNSZbJ5dTbJ2A1dIxoUr9U0K1HJ2rDzC/2iV1QpJk
KCU+fOb6H+7dx4kCxEWiRXu24QM8GSu6mSxdcwIT42L3DLTApP4xI9N9IFRI3W5t
wDGv4BF8R/pl8xl54ngQ3SmSA1JCnhy5tY14oTVNN6S2aeWiKzvUk+dgTmIbFwhL
whohLZ/HAcUN7EodWEnDQAy7ScFrgwYoq2R7H7Tfzumh3Iq5w5+F45/uu6AwT95w
acFNSEbKs0h9IEgU6SACyABIIRUm1Rao1Lmi+k/ArGChSOGFr2GxI/0xNAbkKAf5
AXAPYgV9hZrsPMh+6igE/rg1QEl6y/kwr0QF3gBMPZ18IEihjYWUGQpkElRPtKdp
IzXtA3+vXPc2NnbQl0IHd1mh+Ed/Vu57b5HkuP4KHyo908I9peJA5C/7tNTI9Yt9
UJ8b8o1DdT/TWx27d/EymMX/k6pg3KA9n8HGIEEoCX9gDG3frHWm83e33mfExjNh
/ZatmaqlV48IHe9KopD5vm5unKB1d9vIYpBvkZe93+fbsntStLc6nLp4Ls42ueX5
93akcQtSEliqeibUAkdwbBhhsdLUkIdteBQ35HxGe0yye+lZa6K5HQiyWAknnfjK
Ino9N0wzAVmO+YmKgvQtEqzwqRFHjZRnwVuM4LbkPewp7lr0QEZwBTp1Kf97AKn3
OqcpgZXfMdTV81ufMVpGjVHxBgrWjWoEUG139FK7UKW23jfZEVaH5zWUJGViOYha
0TDSKA211fuazWGDKw09/CO4tA0nYvs1OSOsIg5yiIE8sLCnSmhZXTnHIAx5vzKy
fUl/zPf2OeD0hx9lWKPJnNfMsJnUKkL8exeEY1ulx2E1ECbAAxCZ+AF578oxXkSs
6NpibVXNAFneqojFTRDByNwcAnG60Hj/O1LQMhGLBfax3yrQwqsaDwFmPU4j5evC
RKh1qJt5ZYPVYBQ85EkgBsXzVvFirjLp3csoZYzEcmW+4T3TfnzAvJpLakfV/4CH
nSXsgdjp6JjYBn+WYLolQ2SIsg7H8S+UULtsQHNDm12wSm5nTKoqqhtsXOPLcdVT
USJ96WO2w0K/8iceJEIzBHwLV+lUWCtqKqn2/CNxyBM/lrg6DpHo+UNn+K+wASI4
wY7/c/JQclQJbkUqz0LSWQVvR0NNFeI7NspHz8SINce5EYkwX67uAkbDGtgQjziy
cW0E3p/ghPHvNlVNb6HefGab2Nt8pOHIw8D6PHfBWB+93AfYxfEnyDDIu3gadaZb
RY1a2IFCQadXl+ndKSiGMPLhE3c5ZDnoPBoXjlXhobKXLGFtI1DFFHzekGZAlGMy
vqKRTCr5itROZtNv7Xo2AuJdgFcsV/iUp5E8zSdRpGP5oIZ7IkE4qOHsqYbhWCQg
nmv5MsXWATwszIrLXm3GrmVJkeHzPs/upNVohib/NmWOxUXgLhsgLHynLlYEhEH0
uhyb5ilzEiUf4tXd7hcoEWN5fCEGuBaNuyp5wOjsxjOTxvgpVcmSIpSUuWBA5do4
cDPAWtY7YeYbti9ghEGqe0Itb9OlwG26VfxcGTxnNQysY7Qqi0ycZl5qNmO1K8O0
mv1TN8mf701ntQe5attytlB+9HdBAIeYmQaRcaM/rCEpk7OfKnPh3W1u9Ol/mMhu
ay638CFsKZcGBvWtXZxmz935ew5CZA5FMICBFX55acNpJ2L2iMokZ0cSA+FLT3/5
/pENkSzBxLwANSgdzgw+cuF9t7nVayFy0/2hRSdbhwOv6lSfbpdYeooJjqONlyd9
7K6jIud3dfxSlmUrYWVA1uTsZdMInXS5GdpFJ0vFUEdq1R4G6q7jq1bbTnkwjh9M
LHrn0z9fAASLPBEReBeTRt+T9WzyiNsrsRHQFhG5FRu+wvivd6Tq/EP31dWF6fXK
+xTtjNOf9m01v11bWS2H5rDAt20lM68ZyyIl3h6jhFCgpZPFJ0Fdw967QOkj4msa
6msQHHOhvtHK+9346kDhxutLOtAjYiz3rxA3fYduaNXzRGdh94gDnFctva0vHivN
EMH8JO8P+MmClbkt5AlJ2oGt/MP9VNaRpnfjrbEluYaeafwebtK2ijEoZcwfJSb5
OxJfQe5+hjju1JOP/BEbhHmHaiNOMnVrOrS1Dh4rnknDJOM4sSeyBWe0IPAsfScN
qSEJBcVRROpuL1TslXmyqxBkAA9JiroHxQW4ABfuIHwwstdUOm/ItY222hivVeF3
zwXWZaj3OEegfzCTTAAfur3odBDP0sVPX85J/rxeDYnjkygyDj7xBGX7KW8k//Rs
dh8Acv3gsRWPUsrSZ0GXHduX/5kSYzyh7IM4bGSlWM8l5Tvjdc7Hui4QPi3Y+Bxv
yUHKUiyx6PFnyrDyc7FKM6dBO2epgL3leAMOgPSgD7PZbYnNUzrBJeV2G0hJEBIU
mkSVzqMtyF/FlE0ApH7qiQJcS8oiV5N8JQhqyAuKTa6kCdiNFiO0MZctdapZaGC2
lUHltJsoQq6AU4W5ZUN329mjagSjPprhrFI1qkNk1C/V3u1oB3ySBj0to/gj75OF
QQ1IdqMaVvVwquXVwD/i8OvC2cPeMdRpBvSo0l2eIhkmbH1bKG57pAWpJ8FwCc2E
UP1d5rjlHCieF9sgBEsc9Bw58u8tX2p1MTm+3gS+W4M7SYBtd+l2OKSbIz1CY37G
oZA9+05kSXWNTHJ+HuT9Ixc4BAIAbaRiynuLruYfRHPNDCKYEf2z0FfjnkKuuzeU
mzeZAF/ghAaFk8GK8BoN4FtdKbAGqKgeV6DcR1/WFrqIOIyD1YohWezK5TECSHo0
R6znilTnnM4ZbYxG9AIJzhZ8vfA7biYKTi/UP8y4QlL5BZtHgAmxqGVBVdCjvxQv
x291HEHsqaEbQVid9hz2W2EzcH5XYg9sBM5tVhRaOj85tGu8eSlJ1J3pGi9pTrbV
2/RsfOdOzhZpt5qKBaQaB8EAzMFs5mvpRtS838DmczZOmlhNsuPkdnWbbWkaJSaZ
CK6Sh82hKb2onEpE1O6jBg8Bdy2JAUJ1GygYqFSv9JOZs6b5uzRsd8DLmNKNvi5W
NZUvV3STjvY1QHje2vrqzg5kq2GDXqDyopBNgGKdKkXgH7in2aIe1LJ8l4G5YH0s
Vo9sWEurvXrJHaBmAZ5H7OGQPV74oGZjxTVcJtXdmzTUtaBAkD6iBm/CEs3evDLf
SCFz1R5VsTjSwwklG7eGVLwB2+k8mc5m54X63VNS72CZMSg193tTjQUazcQMpwEQ
jJtEqyxVjl73OdBz7t7UXYdmI711NW+1Mc7ZYm/9+zLK0XraQLH+eY7mGavcKorW
542VeN+dQpBBqeawYQf5Th/n865vpUyc9FFgEbg2dhnWU2AWktkDNzQNlZ4QEy3B
YPffYHmw82DK8LM4jPY3SnYVDa7LkcYcRYk4/1Yijyxu0t8uwj8qIzGbgS3L+cGJ
ZuNzsKSrZVrViE+voVbuLPN9Mwnp4uNShnNCJd/lwQOp0C74B3MjIGwq5nobuZlB
v6Xl5JXbBe/qZQSuHIXaZM8g1lKZ4i/CtE3pYLOqoH3Pcr7RhW2wU0lfYRp3Ysqx
skMiQKP5KdPT8IQTzsCWtGUe5cetO1NFViR+enTqWaaKAF79SZsghh5iehKj0SzH
eVch1ey3H5EpJsZBRGXAVnjNxdr95Itvd5fyk5EhhwYPf/slpNWwqJebJVU0ULie
VozCvBcxO413yM7+mxoXgA1WP7+lEE9ZWUGyiv1oPi1/b+aVNRF1ldro/7yR9aiq
yc3qkvU5QI4SG6eO0GGxbtSomtKSdjPTAbFeBcIOXqlbN8Lnt/i5AdQ45QF8s2NI
21UwA66L7exqFR6gwItxgsacz6KNSeNF8rSgEiwzUrxO6edMO+/nppe9nGbf5isF
LJQQIlQW6wuw7ISidngHeA7E7aQ0jha15fD7/etmvvi7kOn3jlFChoYApeRJ2XoX
FGtxM4HWnonhDCKXmKOzF47W+A0KsTm0SbMJky7qVgvTZMlaJecNyPIVveOKPjma
S6RWHRdQ44/zGsCpRLDXmiTpclGgZkI764ZSoJf44YY2OmKsetdaLjQ3k/6iUcLA
3KlVDeYWgFV9GASJHizg3GLzB/7jaDJv1aE6LElFUhYhxUgJrEJPJMp5JpsCquaz
bp4O1JCz3jXzm03AN2WOH5UcJkrTcBXmCOYjSeXOlJSExTE4RwCJ9m7dj8rn2Jr1
jQKNoSB0b1w7AcVguDHQCUxqlH3OqJYqAyk0l9NyeRhPOfUIBuFR25gZ5AjMf31K
QxIxHC3JieeMiX6XI1na5Ztv0tEw9xoXwoX6qwzXQoy3GLGlkD1koU5yAXXOMU0L
lXhhFbBoZNHPgHpEshecJeyMzzedxdUEK7qRuvWM03ybw8ta07S6fLJDTnqnKVJC
Y2OKb9GEpKZ/wPIeubzz2oKYDIwwcIGxatocX0cqCRu3KMhfXNNyDd23pcBC00RR
FWjNIrwt+CxQPRDJdZ2TIhDetNSLhEklUfpP0B97BSpB9gWGWcvQzCj1HF3S2Rfa
TX9vt/kfDYgJUcpkx1ruHJ/neIspE+3WPPC/VaTKAQmIAkdc2CkFd53PbmhGw3qW
HPKoO0gpsFuR6Q/qiDXTDd8Ig0D1rrG/kdeEH9JL3Z2k3RZyFkJNLKD9yhfGZ0Jd
kVZkrtwRZF2BbSn6+Fmpxf1QEgsoh4nQkDb5vK+gmfb91kzmc/IiEBvlaFyfiGEP
ytFZ1C5/C6eJ1WD/wUNlJUYZN6IMWyG+5qNtj9DlgeUKbB39uN74mgXfFffLieKK
h2HcpOmrQOMjdUAcDkVQKtVbhM7aeuM160wbA9RHTCTu7hOGVELVUQaZLMZdzJJt
Rf9XFrapURhqxT6BsfH96ypr7idXXhq03ro0kXVhwmvwquCIlA0Vbm49c4H23q8t
BDthRD2N/KIcHtpl+RvPre5TPQ4m/FJzGTkRmMVLjkTPcmds9CzlEE5miUTKDVgx
w2l52rMCO60+RUPKVnTZfjb/xB5Ey1aLvqPCx/hlVfSW7jPyX75jbEX7mp9Jl/11
yHJGkeAxny94S6IF+OgeWmlOEXuOtPIgldUnBt8cVwi5Yy+cwQyEq496OM5FVI1f
WYA0m6nECFwsW9TYHTJ5PVWVAhXiMNDF4jciNwjfht+9wS1gWfJpSaqaEvdUqT9U
9p52pCoi3UBSplU4I0k4uYT6GvIn3eZpX+nY7YaEd9jKFa/IidEofvlA6jVjQbtq
AlpkhuX6vrHiPD/235ulneXyg4GmJuMP5ZznKXRPSN74DSHsMrKbUDdxBxviUt0t
bTrR1S74br3f4253xP0Mo+JVTCY6ww4YXTlrDX9WvP8JdkWP70Byq4wClZceiOAw
G8rWh97YJzyrwaTIPC7ESD2ZfLBMFs7z5u+5l8SXIsv/f3Zry0FAJPhgHCUdEBTx
8NLwhnwoye4xUEbXEpvT2S0eobavNS1yEI1KXdUmpI0+7CeMAp2zBnwCdhCVD+J9
FyGrzX1Fsiz6tfXTRMbrxNkzTjVZW76ERBEqpvlH3UdprD85QXlMk0gGwWc01yHI
jBOxRDQab6pNEl/mr5Nj6hmbyEHq9oYzl5wTAhFbJ9be5t7ok4cC0DXPplD8MksU
Ek4UkSx7StZtHpf5JwUmEzRIesZMGfpfT+z774KnMDNnpKZTSKcbhNLK/HjNez2c
QCqoVM44qLjcSWkWF5zTmKyO/VV1VrY8XwDM3WSo3W1yrk1RYkvH/yB3WZpIcw47
S/bjdq5hfR0BnLvyiZ8GaPMcJGyvoYgy6olqEcQcNk5kcpm/4Edhmozu96bGeBV4
B6NPwSBBu/weasOeXmGUsTdsJAa58CDgKJzoYlwGgehtSlVjfrAGnU4ORBdO1KNT
U9oeVCIGiSfj1aYcJVDlRqZBXQivmy7p57gjuU4TG++fpzp3/SN7NSNXsSJNDFTb
Hz4UufHNsTTAQ1/HCLOCfSoONw2t0uCUN1yHANj823FM7k2ljS9alM99Eo+7PRBq
556fvByk+VAEMT/hWdhc2CREbnIrJ2RZONYPCn5yX6aJRStkG/TkebtHxOwLJOXs
DWfsZZOPgdS7L0kEDs5WuftM9GFouTO/WfsszEhns4Ie6blTSQCFcEg9aw0SP3l3
XRYi9lCC3ljGByyQk8LLR7PkiIss/4LSyb/J8VTeMgWSN+BkNdUNgxaKzLwwXmYk
8IPH8qBz4FXb3hSdtXtRr9BUrX18wUEIUKyNPdp5kHWkCmYXshZa/ElpYSTiSsGR
fMmAknDXEmYjBmd09fHgHfNhhdHeMYWHLmYXLZOu4MH7Yy0w9xC9V5NCzeX4nNBN
Ri+XTc3M/QexJn7+7byXjQhpIFJZ+B4XsfDX0Rv8AUtBDkC56MmpqbZ+fD/VLGbX
mA3gB1rkbisOgTxtzFneHcDb3WlHMgSZ57/I1gpuXerkNGqqm9Z24p0LJQ8S+xQP
9A/puJx4YCgoVqh//V6u5OyHq3Pd+oDWMzwMicfT0rq3queMnXP456vPVp0vHFaG
BkCD82KjRoapX70Rp7rRBHU042+CssD/bCSpl2pfLStDDDLTodaaoyS2rhqNhPyt
uXtPDCg8hWRJoyA9SxHuuF7ri9+mIGS9+nCslfHdmSqLfz1p6IUx6va/Os5hpxrG
COzNiRw1aoCu6uPKFnZC4cqMSBpHtfi9oczseYfZhYtagBn/Fn7KFWwwZJ1Nj2kF
4rtvj0Z4Dj95JM0PuoUR7ipBRNI30iSVO4t1a+67CUnbng1eGB/vH+DKx48CWh8r
862N1vWQEBFcDyA3mK9TICv8noDVR5sVb8Q39cyUFhHuOASf8VtQpb+XgYb4XlBk
IIElmOrB00PRJWF4oyP2fJoo/dktlrcuTq0kBFumxhrib8S1RnN3rB8NjnSN27Zr
VTACT9REvkcXcoX0ZR3WFLWwSoh5zKV5doACIFaKhQGShXFaSgNkxxSAuryXlFhx
Fie/sV32f/Wg/bUexgj6+Ukp+B2I1TxmhBxz31828uw3qrxnI6QcCaaBWt/omAm5
0F4xarfmxypIaGqFgEpr2R43RX+ZK2sCO95hAXSez79Tioex86c/iExXL3DU22KA
sZWP7mQmpt76AQzDTGEBByeknUjyC31gpbyiAHrdT2USmH+F3PmdTRYMdGouIoiv
aSDYe5LZz2fNG0nQk4h466ZesiuoxAFVpSSLzQmv0Ky/WcQ1pyLWk0qoVQyjvakm
H7RfpL+oHEUhD3VvHAbNEXxzkVh+VKmFHaSzX1lTYCv4qzWXl1B5BoYlDaAsxSdr
c/3679sGnptSlag+eiwtekudn/0iU0d9hH1ikn8TJjeVpnKR+poJjT4x2yigfbJ9
qQwtLU8R/q1eKIy9savnurZXHH8TG7wB3ymdkc6s5IqEF2V4PXhcaEJ6ee2YhV+p
98c9N0GadABCHHpCUSPE211DJh111Iwlrkj2l89ihIsYilxr6wJRrK5ktmVgrO8p
aioBCNUDSt4RNWc2dMKWiFmrkc6MT9bC8oUCCR4Gj/NGatHefWBUBTAEtH+diEJ+
yjFpSV8rmDM7abfDrwIOsliHLwsrgHOsRG8aq2c9CdIKU0svc7cyzE4tWtx2aL4d
ZZiQG7KL1Vo85xOYx+F+IawX1ymoxzuMfxyfLc3ejny5Aogquaq5NEro1zo4HcJT
O/o06wEU9Thv5bH9KOcrwmBWNCodqxh7+x2ZqYdYfm4xrUsd5TPjTyMfHzjpLzqo
nCDTE+D3n2SaSVf1TjOcaBNHJTcDcqtMS8DZDcRBeHh7OFUi5P/eonXUTrwanxBb
FKJre4kCj7lvl9NYcb/JkD/y6qRZfAlAoPOqhpuutI5Sxyyg0fuNCPG67EpfC/+8
sezpofWAmiL2nZO2HgfwgW3rXWFOM/3jcPBI8tHarCt7V0XxonaM3UHgGt4/oIMi
OlENKq8l2fZoImoiYH1N2v+6RNFx1hfKSPO4E871NR4lSIOCpL11yYnGKdc2N5aC
O3ICgirQsEt9RGXYIVIgj9z68bNDHizSwuHEER5roVyboorjSdSngoxKEYgHPbzA
tQnARm9LplWREG3Eh3ZhyFA3SMjl50PS7M0YaLYQxbNyyg9zIV3isRM4me7XMh5P
NNwwuZovcm4zm03gfV/XkAsEwOc6qE41bab19SSg2+Adrypz2bRpXtOFW9tzCYL3
2z8vUmhkqZjR6L9Eqr75BO/LyAMdslg46nNFnLKWhbPoXr8C+Y//oqgo21tcc/ly
VDQzQfRw47wGX3KMwVJgRD67EJAalR6iSo+D+9j/sJt+/1t1uNmT9XI5/60zlNsw
sjdwiXavnVPHDc/hw/vwYjnfiS0MeyplCLFi/jNqWLlsk2yMiUKAIQEgiDAk5tkT
LDepEL4Cw1GfChlj2mdTTbHGAVVMVamkF9mX99gHKL5WzOtMfO6xcmClncIlMSQ1
8XdKQLEww9WmcHQZ7RGPH1BB6+0PG2kNThim+IBJSkaNy2Gw6rmD5pqg0gg0L4qU
iWEJy+oc2t+muEyRB/kbOon3r7ar1i3P2jQWlAiugIehMkRNpJQHkw796H7hIc6e
PXs+LaVaZy46g+XLd8eb83CBygCQg9TdQUFtckSb3BkBEo13RLWmL1GonntI3vGg
ojO9/PjgW9I7jLFbfXS6IH1k2QN3c67uwcO91XNR+tcQWA2+6p9cwglUcireYAdq
yDexbfnQrDD1PC7Am7tE3pHxYaxvSxEu75d4y8WJIOGgilhb+dgiz5TSUKOTMGxc
LPgvlqGTUlqEyr3fY0DwLj6XRzpURpuY0WWpHK0AwjIWZJS1Fis2LB+uCvfBBt+8
brrpKa8fk4XsJtmqy3+TaaDvytVajGV3HmA7ZQY4ejqQw3sDOuYe3M3bBuxBTdPJ
eYtQBjvpAzNHFrFUw/K+mJxg74H4zbrwRU9oABmxyF68rT8zvRJ8VtQX62TaS/tZ
BuqGaf3zVSIxpT0/UFeKTZ9O02YTzjM+RT8erlsZwKCQvnWVQwMrtdMRppTkJtBW
Ik/gEt1jAeSNt8Etlu7wc0+jyXXtpqP8FY7V03ULGigA1aMrFx7Ab8jjcrMDhzXv
TDt9telCCgbnD/IOcnIS/iqHR1y/DfEt9u21TfGePm/pBWKzNpp1BdV9r4q5+4K9
JRCTh6qWwOmChcf1nMuJHhImP2vR1V8NlDgJJkISlx6Pa2PIb8wiPi4KYWUbo/3P
awcMChFZJ5YZTJrM7XIyGI1JUMXlTh4gYAhb5Z19lJk71f507tVJPsZvWBfY/BCy
DS6fg7YT+sIR/I1lUACnwFOBldm7w1zd4qXeHXY22ETxN6Ir8Pqx+HaSsnBejrCH
+8F6JWP417lC8QshjREIe0ebMTKpdD7fhyh78iUIv4UaeRquhzavkcJ1vI/tWwpd
s5y/W0+TVp+gWDjLaYWrDZQ9jaioXsHt/heDNlsHpv7J9kdGrlyNMG+ekXnsHu0A
8qwhn/B/6Hv/0PzwHpRnFwnkifwg1Z85tWVzn30SKtBtDVymF2jRqYjCnVPTc4T4
pcnHJ2+1ZJfwgsPpgZ6P9zaXmuWN+mb/kNnwEqmAIhrdLw/q2adOMpBzB0jg2O4f
QVtZ6iI/7/lTyPw00vyPwx/6r6hmD/+nl8zMf7Cv0lOcw5P9zQCD6TEuw37aV4M+
o0kuGW6SQfbU61ufN1L9cdZ8XV7e3oMJbgwZb6p4iAQYCPkp9MExJmhfy2ucK5xy
a1mscducVfeFZlZfcpkG1GsDJVoC/wZWXnh31EoYk+5knLF8WZYIRidbBmtBSCyf
mnNDr312eYp602aRA/orYaw8U8Y5ZWvDpb9bsGpi0UyeMmiwuxWHq9bKutNtjxwr
4A7XDv6spgdI+Zrg7yLWJgUHbVQCnl+UNUAc1JSQs53L+8rGMvPkm3BRxUReVfn/
svEXzyzSSD4/V941d7lE4aZwr2+DWgUusJgvn+7pEVEBz39iIOWEumkmJ71+r8Fu
j3D29vLpzA2ltUxLAaevVy7a8SZNnc2t8WOao+JX5j6dbvVWiQ8H8K8pcFRMhRXD
Z+9WKZBDSF9Ep433H4uz3aFf2EtFes83kmmWjdak1k80HsWea7V0xSeg6cY9E9K4
1b296qQHFox+bUsyANQAJOWZm1I1ytO25UghgNmV2jBT0HVmZpyUgpVHhAlHHLVp
Zff2/45bjyB5qyYtAV9RcicU+9mvn9bMY80GbwN4M+8JUjvR2U53FyNiPdsgkL7Z
PIBm0I/aEF498hSkGP1HtrX70IyJ+TSYI7ijHETfiLdBDBMp1vCT/k4kwWqj8kga
eTy0xGU2e/tNP7vJjhHgNpgl9OxGmTKsl2nLkH0GBaf9/NT2BOdSL3AmT/uMLoBr
pi4KM0JqJjnguPSxrF2jfWDQLryMxlzihutFunPYLNR7ca+CKA2VKRXmB9or9aRm
qwtCM4Iq96KG8UyrYRnbQxk6VlJ/hA0w+nvrrlTYMilxngdjsPmPhPuouEHNGlYw
MBNLiq2tfqQu3ziG/TKwK3JeY0kEXSYvdQGlYCW51IG2oMWK7XiogUF1EY3j0xmI
1RuFzO/GBjHu0RDhv2pcEu4VyKpeHeVGsGBelxbLTpdAXFZJz67B9IwX6mU9WU2K
3nHIeHplr2KAgoE4K0+Z39G+gzJciB2by/2jxpxajYzxTBdFhRyzaeMDix4+pcn5
ZtfVhLmvlZAW/9GZbNLXxs+0CvzwVX+lJ6BtAQBZ0wyTT7+GPcygX/Nqcsh+n8yf
buFH0ew2bkgXgwYaJyKP7P1CwI8fVZCCHzOXguUn+Fvog6S/yTALBXgKaKSPBVal
OJhmnqNxOlj7Ckt2bNk9mUSwyFrsSDGyDHX0FLkdvVJaJl8ZSrGh8bPRf9G0eRE6
syQHsY1NQ6eZOWrqR07a/6rS28h3BwcIsH7ZnXeQ/H6Genf/gvr2qhUV0ly9UJv+
Kw1oU6uuhJ4Qew1bv0AYC8U9hNYA5YvPi2OYzrqPHBwJuJWC8u2/6KJQ4ublU+Gi
l3oZ6+abZQ+eJ7otNp9hJe150SXljHUD/WuEsQ1yo83krehp9sGuRc6xUUy4yYaj
GBiFYBFAYfPGXUAsDvxgpHvkiUrUwhc8loL9bm7NJ4QjiTvRtPDu6ZcJQyrRPq3W
sejD2GUbOeMaZ1zTE/0HmO1EGUB+1pN58TfcOqfLge/u6uJx6OZy1z+KIgtg5B0P
B/29MlQi09vsZZnTeXK4kdv32CLgoy//XSyLzfsFP7wKRk22+64vFEz9O06sbZVL
Psgkf0BBfdDNtcH86VgouqknFFSmYikS5LkzDtsBlNhM6aufGefKbtVM/kbsQrXe
e7mBbznqi4Cy3scTD2G8daxuip3pGB6/EGyqMsg3y3VG8f+VzaWYHE4DuzTaJor5
We3ZTay1BcUz/Xy7Ls+AIG/i43LHNeB/q/pxSt8KnaSMqj8a13AAOSEBs+eFUht5
oMpFFUqZitWVCsFs0CFiyS6xOMPkDV9phKBe7nctgYMJDtLiFamX49VlBNK/wtta
nwSVEMGfQnPIbsM8U1YJ9HskthUel3QZTcDMMS6phv3w05P2R6B9qn3gr8m0mCW5
mDb/X6jKQO4/euSbdcaMcXCarvFvP5TrBWr/CvHKzrKUTszftnKnV/WF8wKNQXvu
CJFoGxQWZSQVm2eZark/tRKvzEmEDxwy+6Lbk4/R7YRq+At4vImKsh3lUCsnoce1
OR1xYE0ETCVUwWJMR5D7CYblxdpC5GluFzaXoTC+eqkrpoEpmkbKWuZRGDAF0eqb
YVF6L1acxIVzTaVCGidIxeYostFR7m1FkvS6f1uCszdINtEWOhwwNjUg1yUYAAq9
jTgjFZdKFhDCsWthHzrmVM9lP+LEUIRZezFwqKytdRKb2lH9jLFYcjSD0D8nm4z+
3R3gtnzVml8jjMU+tk8lU5KnnXOMzfxKIvoefpWT+e/P0/pnIpMDl6LJ8r1/C+Bv
xq7xJJD6sYKIh7Gx+3bGN9AfpYZUVmVcH3qHgDTNmzlb059nwDUiyRgCOmQjQxJy
FQTr+6xrl1WlfeGs0mpIrsl1zHdQ6ICU7eD1up9Cv2lBy0qZHmQqxKxcEnSSC49l
uz/S+09/lIWv77CVx0Y9AK6OZTkp12ULPUnG97lPjoTRWeGjnCKac/ZDzp9It7Ff
zPiISBwgZA5ydXiSz6VuWTpWbz8v+02vNGICcs6SXvt0uQqCe4pyVNmZFBy7ouLj
LfmEN250AlggmbB9lbrwSXhaliCvgv31aqX8w9BFLCtNrWFl//4atgUqY3MeHcaL
4fI2F0DEOXrvju2nGHBeLMlDme08eiE4YHiLJZ9pyMHcd9mT8k6uQ7Cql1S53Jh5
4IZB/xVh1yLxwkehNG/f/a/gkuJzz83o2cb52eK714Khn1BnWVz/O/szrVVnOt1L
lZB9f4JMvo/R0+cvaQYSNg8abg3KeSm468DxFac5FHYinEfSDwNYvqfmCRQCEWHO
fzD60kRYzGKg30HF/65vuw0i+O0IpY+JysMEGcOkVpQbU09C8Ap/I19+AEQfpSsT
TzA/khX7OMF3fIe7h1d45a8SLmy21ZJ8VWjdr85MsBrZh4ejaNQI7duld/HJuuPn
8pHHfU6uA84GOBhz/niDDlSjds2ZEqhrSmtF77CoVHV80bNVmoDNRVjtglL45U7G
Lf5tzuph3JG9byeUpMSCDmBSymL73q9QpBPxRFk+aFMkQJ0FaAYilAFVlVUgTKND
YA10iyzP1DM4MDUbjLVE7L+bU+GVQKU+WtybX0wnWQhHWa1HuHyY+VqTCwD6eigi
HvmNQsFyO5jKaBFD5IFteUKZCIwYjEpYWdrhVe/K9pNJC37Qz0wHE141oev2Sdtv
D232JkInGaNokEawm4H8nsLkIzDz8OuKR1xh+plRYGOZn4r9cfqzwp981p0c5JuL
QS8V1/X/ptEz3wrp3A6j1edPESU3RF5xZlyE54YX4EsjQoKzWt8krrDc6XnE+kMu
CBcr98Hm3x47wa19NVSZODQ/duhxzPrqiRfj9a2R81C3LPd5XDDSiwyO9hYahgbC
Ssd5S/x88brZVnbjbcMaQNEeynq9Qfco1HcvnshNiUmxbRLyaURKy2JMZtaUhRgc
sBhd6TjKdbXvyjIGZrD8Hc6077Xd9FLGf5veDXidAJlQBzk7J14fk/WjFQJ9JRwe
z89TmjpHcYzQ3/fkm70Rc73uKuTagMKLYd13NdQxN7LxbGPjWVv8LT+Sca6sYqlf
JD5YVaIMDz45wu/X3Ewv2kDjlha0dKL43YXFSbE4NLu4ihfWLpz11jGcchNWgAgr
+z8EXHwgT1pPxzD08xiw4hgiukzzULdr78e3zNutQHp7Vyo+D8gyT/1n8Zg1idtV
hr+f9yc3l1U6t7XhLtXSAzE55Cddl9fq4taOTocE6GxLjlpR6ckjRo/16DJyw0e4
uXjRtDsuS9qoOpeZjxWHE4bQiDm55tiA3gOW2Kb7vq3wrQa3YY70jG0iKBTkvSQu
3gkDGJJyb92XxkLVHk9qNtzZCLC7pZ+MXrWGF82qKMNECVrwgaHJz10vhVE/0wR5
1hXH6FLQ4ipQp4oXP6QG4FAoWhCi81ANx3PAMJY/MXnkXXiZ+AiWVrBIdgsBTlWe
V+Ob6S7sgb0wJJYXOGnoDPryt2i9PW+GbV8Ca4CmJCxwm1nQCvOvOYZ5wTG3flux
6meclga7XDi/gAqAiwCqw8Pyr/yUqcryiLEe+ZT2q8YQAHUQmOKpVE7nqcFQvEQ0
PYkn/+jJ/iBC+3Z3hphPC/UhEwg7IBtn5AcGjJkBmFkcgjyblCHa4npTxrNNzJWH
Iu6/5xBXPP9V/CHiJpWWEh3c1yR093BqDF97BsHHnKucKv55A0YvuaMc75CMzUP8
wf7GDy5J2rX74yu6vJKRcM9W8v1GOM+omTVi/042uyS5DljbO4DaxkOIP5KBLcP0
7ANiOb/4IUkz7nkVnC7xbBfrGKWIAyqGMzBmxI0CXtfAsPvPgC1DYHLJrLQRAA/1
2WW3g5U+zBd2wGiyMjE8RdGiZ0sdWSlV6Z0osStPiQIxk1hUzxup9oi15W9b/DlQ
QLNYHn10VG3nA5zNyxR1QC0O0+hAlAXc9ve24QFMPOrD8WbiwV5GjnQx3j15AZUp
N8U0QMTRzeIQgaw8IOT8CVd+f6t0CThEuWBLUi5kCGzVAt9aUb32WQEs2cE6sW/O
zz6C8IEw3ktPap+PwBMOUvMaIdyFXthbHAeJQM80IIFSteWrDxOjVOiedQrrvjxB
fcYkUzPuCc0JoJnN+tGBcdeiYfiLOc3cXmLFdp9MYo7oAIiogltb5k+JcOTTxcJn
tT+bPgWxQ9gqs8hmMWGEEFKiUObf0zWO9yrxsvSH+tBJ+FRaV66F5f248e6QKIWz
tOYHTEwuo6JYAsYJs9yBbvItsdmtEZM+gt/eQfjZpoIcXV6RRsMEWiHPIp7gPY6Q
B7AictH/lwQoGwwZMBHnAL0sdXAdB6A2Uap8UvY6BxznJoIIIWFKGPjElVYxr6dk
8xtfVBDfPSyf3KLL2d/SjnIJ3dnWW/ZGup54lL1A4RSG01hOdY73m97eROubgzLn
d6ZM+mB8bN7Lyu21xq7tBeCKR8VQ+anZkxh/FWw+t3frvdyOCyvXvdP3BLKZnIbh
RhFwwkzBKDw2AGskrm32uwf84p3j770Rz7OfCl8qyru0SU9UwH4qL2xYYPZwHfdb
7cz51qDI1ItNHHHwm5Q9NyCxzZBT5FuGSgRav6jQVyTBRFLL3b28io7pbRxZfcwE
bhtSihn6un3UOdkji6uB5b3Ybw83YZD5HOAFVoFnGPDRj5TKRkDDAYlS9TF2kYs5
ZjqZgJiegWM7cuBaUHXMtKr8wrjmWnvxn/3IbcF7zChPhMwv3hbe683dbgYjVDfc
t1n1fTVaeXCobiaFRkqmKbvkoBlOcu5hcSHXUhtjcWwFfdCoztXeH7TkyFw4eALh
LI/+NGRjZjZLHL1JAcyu/TufJ7v1+lwI4jsOihmLeuGuLDYsSbB4kQ1xFEvzKHhw
qxeGMG+E3L5g3PNQXwCxsg7vevHBYr/rh0+DmBcyQ+u5PCVd2FsC5qxnhL/l3pZT
5cJG+b/at7AP5/psn4Z6yW9Wn1X4l9lzxZu+H4WJdSIwbW2ThFWBfeXxplOqoJ4D
Wwrp+LdqkdZF76digOh1IHKeBIKwJK7hsiAopkZGTmI+mbi5wvtjw2E1bc7bbkQ3
oBxmW0ysIz1TfYl9mtMfM9NaNVgBstThZFIEsRswdhw51OIW/U3dcwJUiRmzy5SX
7wAD7fPRI/CbneZvKQqKh2fZdKRR2ZtMzjdx1G344hbK1nmN+XNnA48sGELgDDdA
xKHrft8TIAQkv1BQgrc0NPpm++vGEjYitnFQZ6IWpTW9R4Pj4fGKbT7uKPWdL1Zp
+lt5DiBtvGDKn29ckAHasoE65SbaAw+9RAIE0p/0qb5Ut9y4uu5BlMo1UcQEJokI
jqujBFGGLOMhxfn2eae8U/f32yA5jwbd9wRHwqgrRWyoI//sbKzxaw6+zhI7zVQX
cqFtj08uAOCKDGx1gvaelkKkEOHz6vpZ2YCYl4JOqabl9t386bbq8ffHyFOvOVwr
Wf0l57YNy9mGmmbLqvHzqR9i8/jDXmwp0J2Sgp8glvi7+P3Fwj8GBGsCGf3Svlpr
fSR4Lx3m7DQWVUZ8YdV2yMufB924NYU1Meoj+AudU8wlYb6R3hrXMGaNRO+EwPqT
AB+m6GUczM/0Uw/TCcev5ViDdxB4FV40WUFw55V+w9D2ZiZLYzAxPsxJqHC+ql6j
e7PlpiHZtVC3EUy8s//ZT4up0fGO6PJdGhVGL8HVjiCDcZgeX8kgaBpGBo0LwVDj
0Al/hFSZzmY1lItqvelwge8CYvQ9CMu1+N7137nALGA6l+P/C7s0AD+bVpibeR9Q
e0DJW6bVdwq+N3eT6FD9NwzKhE9bcuAmp9zwLFb3lFNNZ98GuW1FnbKR3R166tbA
J6bV4vZbFxFbhKw1I+uSpIU2GQpeTeMCcrXFNVjdbSYX6Ir7PO63UqzYrOqyCdPI
yVsPK65ccu9cLKh6E42C8Suuze71vrF0D2Mpa14K/2AUjw4n+rmkIu3/I4mOpGNs
GZis12Qcm2KTnCH5QzOUt5+j3T9NuWyA5htNXbH6OspQVhd2oVp8OIldZKbrgaDy
GrySwXHaluETPDWblnhtumLD4BH3dfYNqX213bpe0iYkbwn5A7kUDkogT9YlvXOf
g2i8upUIyPPynkt5lol3af9f8Oa03gI6/+7Is1B+QA2SbezlLlcIWDCM3zcgMxX9
YP0dXWNUEXCNvR9NctI2t8GkT8jnJGcLBpvKfkruGANBm+lXVbJ9bUv09wjZVR0W
/YN/OTxfwV92asWSuBDprRz9fFG1jQd+y57B8SAV7Vk3BgnxSRPRMbPQWUrp01Ug
/aWzZK+tRvewKZy/I9P/5NKQtE8HAGBCEw1WMNzBmgqUderWZWiU/Maeno74oTHJ
qKDfvtgvIi7bXo9RAhsdkoWP8AfXOPG7niaWuO8pEwSq6/jX+Wt4GxZN4zrtTwNi
ZhG4HRjiZdgYTVnSVH47hsb8QIBItEcOQsyhVWDOGMzGw+S3oWp5/4BR3KPQ9S2m
BJoWOKuwAisvlxy7PsZBGvKrx022ikth/b/GetAJCOwZMu/uHzIZt1N5llfKbY7d
ZvY3gS0Gu+cr4Ukt+3soBUh7ZBkX+e7n3ssXcCP5UP4WSxP9MU3yxm1WxuSQgd+P
RlDIhoDy+4c3Dg28aehWPrFpTtoXN+iAgU5EIF2xgaBsQAqNWObYEt4sLuiB4Q0N
SjMydxgCRDWWVc+Xe16SgYc50d9azebOycTFqlKN16fo8bufAdc6v9xZYr4cvZbz
GB7w40AF/YUJFXeAGZB8zI7oYoZAtV56vWm8IxP9+ztQk1KwQmg9KehoQdKW+tZ2
m/7OTSy65JX80MGj7MZgTsniiG+vgwgXRPwwgoJAYuZIuvkx68wbk7tJHZnpaQHb
gJ42BeVjcf/NP24aJbzOPEMUid2PXfy/ivyivfHhWn0oFcqvIox+yaaU3aAob/hC
RMcjKfsuHiLgZHeRnsl+EhXxFBz6QQB9DZ0R9ilAsO1joy1BOutbxytGnp+UsQ21
VqUCOSDOEX2OgajYNLjGjqCdRso5b5IGNgO6a3vil7vfyKPam7i7NI2bfQZxGeUE
PUBCFOK4+ZJfiUW8LaDsC8rwgPhlKLbgx34cQmvs3hH1trDc4E8pJnTMmpCEH+9s
DS+Fyfzkrqo3COkfXnW0nJQ2Yzoqqfx85cOMcCtJLDEu65zFt3gxIVgjewJQ6ahq
NqoHk/1fHmO/gr75HgqfVQC/QHwXMZWscuMx+SIeXZUDOK18/GFQsqX5lcRaW4G9
Vg8TqKPPBT9TMEKq069XOdbzLqmkiNt8D5v3TBfHo4aHQMIqOuiwk6Cv3khfjTom
RkRhno7riAL75PuJFmQqWl0RwPEeAYndkW9Ldnev+FW96rr2EYy1JzjQbjnBnWAv
WldVnEQuCS8va8nlgCK2AZEMmhe2DOUzF+dYRfrBNh9mWfqlp4LIkz5TyD4ClPwo
DfQYMJeDRM6qBaAJgI8YP3+Bpl4PbNEV78XZYKsW8T9okEsWkQ36Yg3K9DSrmPXz
GLQQWxs0GF2Gc3dKMY0wi1077gFAANT61wiMKw1g9aXYcIrX4ott8+BsUvqZG/2I
MqXmfQKrnjTPV8UKmQyw9Zbsjv3gA0wX52EGngKMcybhyzdubswX45XmLoo88eFB
ZFY0OcUd59FhjA7nN7uRyhnuGePiCbZLjSoWE3/yZtbUZYA/Sc8wJSnpQtQmP7gD
VQbYqDKtehGPz7I9TGe8F1JDpQCwLh4/L/JFe3Zs9GnrO3rQfUmihCxI43qSejLb
OF50pV4DWYWpmK7lGCy8qq8325hWv5W+JJ0aXLvWrDPJdHpNhSyUmUBuKQlAnPzN
siDFbIJ4ffGOJJm4+OdlLgr3jfR97aB7PUoSR+ayUQ4293G4UE+E539xvHdYtJtK
RwuQCvleXxr4gxA6uG84Ct10Rb98oq1lswVl+Sk7Nl6Sms40MRzf3BftYwuY39b8
hNWEoplMbSU39EAw9qP/cNHF2U+fKXI3rcA048aKuYYzQwZHlvufVtf/een05voA
ZAhx8nkHCdGilalOo+aeuhdNvZ//Nuk0LwMh4LtKINn9zD2fP/r0FeKwFh4wAX4k
iQy4VLy0g+bMhQYlJOxCuU22xlYzx49HmMs0PFaAdvHMD0ISA74vrVTbzBLlbPmK
RItFpsOU7WxqCVMxEG7ufnf9sclMFDoDayXR3AEbG6cuj5S+Rf+9Nixhs/5DlzBu
mwzvnsxGZkHSxo5K3SV0VRRx4koQAkIQu1Dc2o4Cz7K2nU4yZokLTH83CtOJ2o7Y
Du53ItAxyVsQ/ogSi6/RPFOPL14x/0Dht9fyOpQ3plDz2sdQC0tJCD8vAf8l+X32
NE3KcfDddkeLBwQftyobWg3UXK1pLpTIcEFsRdUhHvX7XXeut37fNmnzYbptTmmj
VNoeAwkUyIV6oQauKCs8Ca1IiYBYNv8rSf3D3xzNM5E43aUieCiX75hDCdyQb7RL
5kY2+BtI3B+Po9SidwoKkblazs6ZJfDIpLGmXdiYKD8PKgAjYU0EYZhj2KFtGvJI
WpLowEHC4PY2HSgF2hufpdZOzHj/SFbtmDH5yvRLAyj8jsT1YAGjoPa7riNSatmS
+EX1+QRM9vPeWnahV7FPY377/nbVhduQ8Ot5jtMd/m+bDRTH0WGmk7lU1cggyoL4
7rh5/gUlJFQ30UdPLde483kRZoNUcBr1gt9UMf1BBFdLGgTjWsMQuVYM/ImejyZk
0kQMCwMC7Wj9DWMNQ/hxhIVGIh2OiR5ZOj6zGJ80VDYJ2txAjG+VksPGmTETU2pP
QIihuz7Jcf7OTwB7FLhend1X9kxqC6uKhUuADeOypTpKtvAeJWYojEoJLFbvvIX5
Pzhvc/mNHDX8hLqP+2b1O3dEchta5dn0V/bq7hs+634U5yy/tqzHzRFlfYmCgwD2
Xkbs0jDcUv8FrTZEAYjMyxwvzYkstrq1HTIfyVa2AW4Tnxy+/44Qb9uU8W+LhhLM
oNhsLxW8XULNZ2hVfvcpSfeKFM6xQ/Yv9q0AKgJ2Ky/FwyETsW0vYenE8mx/vRKg
zYynY3vbNXnJ7+H14l8kID5vp3+wC/FnOVM6t2dA1B9bovrAMLb5TNTXVurGHBQH
3+A2LG4FTTYBYLfzay8WJdZlqwvjSFb/uCoSZJ2N5SJmiyBipOSOkvvrph93J9d0
P4bwyz9F0DeBjyZ7GV/xai71rzTbCFLAFCQZCYcji3z1E+aXOUGGrcoowWxSUwJJ
oxfYl5rWYCURqJUYmA7xupw3JuO6pN3EgnNKtrMqK72rq5HW2yX6oK9RXSfmUbtL
dTI7f5CziJzShSvng3VTCmxKQwoptSTySoIHXGd5bQNrCfDmuK1hj6kXk6ci7Cbn
G5zgE6YJ2B166iu36UbIV0oTFzBvjPRXfNW3lwyuIWLuMDQNgwfLs0GBKxiP8wV1
e/zdLCtzKJZQ+cb1fwOjUiYCK6IHoxGoe3PwguaHTHEySKOnMY92iH/pnI7aBgYz
XfoCw8s9kPArJM7a3Q07KiZkGpgzFN82jSIQbDkEduiKrx0sbgHKh8W09gfXM9Fd
l6MPDnLI0e1y/Qujfnh/FIwoSW5js9ZzrcNCW2aOyOJkMhUuS4j/MQ9bzNwsv8sq
gukLwbwY8kISfm0Uivb8ScL2XYrG9gh+MG9xEGYXuWQq47Mg36hIqiVIyBDEE5eq
9cu46ZamXHUPHPxdh713IcuaSbVDBQ2lE0SykajtGSBkN3cSxmVbgztlHGZ9zitL
omiBIqHnjBucSnUPlPHpY6ek5x6eFrxW718nOPiFKGUlzOy5e1q7nACFFU0emdh7
0s57+LYM1nUdk0bPxi/IuYTW8N4Vg0/GIM42TBTxgMY4yGJddIg0qSW6Tk6qeDc4
5pfPuNew57+0hgDPOmbSEkx7p4F1eTKFylrU75MD6bGekWzyvpzqgylb3B33e/nF
WP6iFoXSRqlXLrU36A8NkSEvoSWH4vt2b/Tgxzr0gYTveP6GClnDRAz0BLdcB2Ul
XdT5m1XMQQ58MsuwfHKKy9pzEf7qkd75WJ7tGz0iPS/JeBG/ySjJ+Z59U9hK/AsZ
Aia5Hpd7Oh1zbb8931wECMtLL6v4lBY6wQMNtRTksUa07YzpTaUbSCaZXWiNgze/
ahNrjj0fItcDZ7TtDrbyE4+rEnYc3S9bNFg9x+cpOCVF4LFAUSF6JPpyj1jen6QQ
wuDRpuKKTPEM1lPZEDvfpcBZ3t2ZYnLysqf9pisHlg6Foj60HFMyF4o3ErPElMaA
qetw33wSs3/IMWnbR8i3xu84bprH4zyb/s2Guuwt1LOtHwsUvx8PUOWCClWVfefJ
GfID0dycM78DIqp7P/uhH3YV3vMHfiX3n7cT4K6/51jhevzAQPWJgU2Grzd/i5pX
xIEQY799oJiuvdaCzRWNYOFXlysTJZFZ1EAvxlvScvFO5aWo3sulGCDrHLrxFvea
EzB+QBIEEyg5wnlhgKGoTmhRJB2tMEcE+HpRQwBt/Bz90d3iqhwNDsL3BVD/4JRu
exQ2HGhudeYd+K5Rba5UgRkUJV/Ar0tpqz3DgCRzfamdt443bVmIt1O44+x73AI9
tiN3LWdDX9cb4+IIVnpcGPLyiC7pFODthmyezCMzgaB4jpVNDLc0Q9r/mcmMSyrg
/f2G+5qAMuCsz/f1vxUebqKeofhl2LwWYkHdq6fsLRZhJp0sPRu8gF1htFknxxBl
fOTAwtu3vPqhja2byg8crGYObMEoV8+8GIae2eGEnbS0/92QANEu3DPPOhEU63WG
5BB9znQNzeg3xjQ6zn1o/61nJnzZqZOw4jXoNMTaQQfz2gAPCRE6u9lc/v5rxjt9
cyuypL2pC+8EyXsvrqMaQTZeGxk7KOcDb/DwZCxtkQA7aY5XfqTqoed3feL8h/Og
Crw2Z5CvjOQmdTUX1ck+CBexPiaktX8tLYYofCmUwhYqRV9t44V/7Tur/9vIccjz
6n7RXbyRfGZ0abuIjn++dsjXHQG8SkyCpRtaXU5udpyX2UsyaMCDyL1Bs1UPtTLf
xqBZaaSzj7CDrJVSraFl/rB2+6hv93DcSYXZX4tD6suFThUiehXYrJwHT48fDJAf
K7Aaw1AEDQQUsfZWq4MsME+2z4m2RvgboDNf6RGQuByDo24q/AHEenvYtYwBVJhJ
Mq8je/8BVsnjpgdzvM3rfvYoQ9P90p9vQsWHcHXrZPsRziRqp5P6Zuf88hb3hZF7
Q9com+UtExSxPmkoiwrAoHhOzt4dP4NyW+RiCbN1kmSvKgNn6RajoWVL/cBxVsXR
6W0ert4opXa67XgS8raVr6ULCZ3P1B2VW4iTBt/5vQjOXCCCTll/w/3ND7ugzM+x
/aAcM+tVLLzST1zpmMen9N2eWYiZH2UnLXdRY7kx39iZgj6Q18mHiRgvkWcbBt39
2IDOyga03xTPZc4cLEvKs42CTrRrZ27JMGgkLOD7vsnnt3P35KHETaGAVyZH/CNH
/flS2W4Gy38crhE8Mc13cS4DMs/MIV1/EuFniHuoaciPe53VtFtIHP0gAqFuh7TV
kaaoW7w9/sqHTXp40Y6cx63GSYWM96GLmPx7Q4dcLpL8sTGlmd27kQndDK8krcK3
Wq5cIJ34MSyxADRFNTE9R089+UKid53e5EsaQ02gEWBaMdtu+JsYIofuef/9y/OK
YW5hz9it0m8wVbPysTe1c2o1EQE91cG5PII7ba58y3lKrT0+eyeaz6FBLSwnI8F3
/1hA7TZQrvCIwZeKn1z7MoGADvZWii60v/Z6zwnwWwIE2v8OY6DUcb9qUSiL0CWS
TOuVt+73/Mwni4k1YvjRqgaNQXPxpc2dzutXrmGTEa972/fecp0euSPJjF38SGxQ
0HbikA16Rt/Io0Ce3g2vP151u/vs4+IdOfAvHTJjO6UVkcAyIziWPr+RZu4B9YN6
0Foo1bdP5KCH1rNWlzbG+JUA/CvwCSBUfyDq3wTIMuRN+yTT+ZXahEar9HSRUY1k
SiP3Gte0dBJENvKSZTRgUk/LKmX3als2subbUdwImXWyYLtixEoQIGTkq3zB3sMk
8n0Q6cABAkeE7Cm4119YjBCj42R0UihW6OQ8/quXEdbui/lPylJNHlXTi/4V3zYe
DDYNu20ye/Bcfbum+gjTIM8xGRaaOAnkI7RqN6arElZ5ebvtmD2KbMbC4p8wocC5
PuMujni6G/elVNYALJGLol2k1v4GcyVMJzzZ4KB9d6VY5huaWOJUb5a/uq2KlNEw
zmwEpuLwU1tmg/G6CCeDZZNMsN3YkpMN8g3ZqrRCHUlvzFuD3wQbtLUyiMOVo+t6
iBZWi++z7gsIz8T+poiT1paow5AEAE96zAyH6q8CC0ahwXX6J0yAT7+AkffTUHXr
OaLKGZ5T++q/yFboh94Sw/em10iwa4EN0q9VNt42ZnD3OTuOIJgAfrzisbTp8Vex
cYl+/x/B3qaHeBra9UenC3hXG/0C2tI677BIXSRx4Ph5KKq4v123HmYouxnLlfZF
+xUHov3RF3ZHmb/jp/CAEJVdNS6fE6O2FW48I4eWpCWamRIevKtJxB1xpVKJLi5+
PG/MgppnHWGaxW5rZoqS4gJWXtb5UKlOcpziYVMdqqEcCDstg94sgu6pIBj5ETFM
XAF4/3EmojItdJb91BoJZqcZ0qwOxu4/V/2DBYooNqrEH9bIbnwuQFHo/911I76i
aLQy/EthqrenQ+nKXrkwad5Badi5ge5pOoKRidxD+x6KHrZr6r/peG6rq3uDZ+jE
vQCsDYBkv0ojO7sIz0bxxAqfBYdYlBzXK3sXQgYfDdSDsqBmI2MUh+xdQwvyRYTj
2ubkb4/NMHPS1KcZsfKbWZJAUBl3MpMeqRwhZfsnwGLi5xtsGXQz6OUtid3p2LTa
3zL4u3YP2G+4+L6vidVlqyRTJlZgq7xJCs5EaQsPoeG/LGA7z9pKvuKVGaL92oST
0qqaMetm9OAOcKXVDpPCIiYRxlnrkW5yNgAuUo1H9nkmq5hLfHiaLdEo9Rw/m+36
hfNNjr2Mli6PudlawNb5Ap9RSOui0GbaSLH1asxe1ikPyPQA2YhzjUZ068HG2wMs
EVNGgG4qjU0tji2OwDxGEytlDsaAQWsjmVpbojbgTYOMVCT7jgkpMudQ3H1o4Vq6
AzRxj/8TNI6qN/gbTuIz9hSPthOXE2mJWz0ZQ7AnUbGHeYEVfgvuDOXrqya7XESp
TuWbe2TKIdgyGG85kT2rQ0YSZujww5A6+/EmMrwckbgRpCZHKHKqTvlDYhLZ3JjW
4PURDu1hkUUjL8l27mGa8aeQqY9j6lcqhvyNtVwNdCKlXao+7JtRrjuvAY/rXaEN
JyCPMDuJ9WE303Y5jure12aopQ3qBDx4YvALeHtVyErUOX8mcsNDJ8HPGwWQor9X
CilkyNofRS6tsot5cD0517BL0kYcdssVQhBw3Vip6RSFmWnGSgdPeoCvurlSbUdB
LP9knFMZAFxTXRNk6Qhh3qwRQ17JD6vHSI7acCjpPcmqq06qsKUknK7p4FDjn49A
X0nVrwQq3Y1kWjszjy6XrMlfFiQYqabjok6TwL6c6EH28l/hxxcKKme5JpIwnSGb
TtWcLJII1oVXwZRraj7GqC0xxbux/1fK1GJGBxE4J5UaPdI54yB2PHav30o95P83
2mEqClT3kDnAQ7I1U08LFdfQv/QeOxM4JzYpGRIYpsLZcE5HWAPSZC1MBoK37LnF
C382S9MoDiQBERMLWE0WXp+45dy/+x7AIdXxiydpB6xE20X5SoUphipg+6qVY0Wy
Qks3TrPQkxGxOOsubzmfz+GbyzFRSJYGvrLYzGSBySWXV5oMHWz4hIIzYlQqSE9i
MtVH0vKVvKPErI05X7oof2ZBt9YA8dOllV0cXbfYF5gdsJz6dA7TEng8QP9mnYyl
iB0ohX9y6Oc1EuxzNjSuKAWfIxpVbO370A748WrYE2PZ6H85GTz5fqgcqRDtIFST
+HQn9WSpQ0znCBOyTearIDAGKiRRdrILjHGOGr4/ksxeUHulf0j4Q2szx7Om5+HG
ehizCfE+yLSRVT0VrdbGUbcoAiY4tax6TUFSpNGVAL+bWDGunqEKH4/WMP0NmL5R
EPVmr4HMyFNLuqJadmBD4BXLZvPlEa0/cZ2+AcMMbA4iRREhzyz+/7YFbmnnYhzN
PDMaWP7P06UrWz0tNz0Z5mjMRDiZ1l1ROqhxwz5fYIP2hYqoW7g+m3/CjKORFqjC
7BiAQ52lfKGnBC1RFwSGWffqx6PJspP3jz8qVYiR1RgN6Mgo+ZIma6Q7Z5lYzBOz
METpQtmQtDG/sspJM5T7BiZsK06DDxNuquynJrhtR5MPps88f33Dt1KbLJAc4kUC
t+8Bk7nfvWcaoMoGDDALl2N1zDhaqlxdNE6qQUt1gedsJHD4LE4bjJ3bTP4qRb7h
speEqgv+Aa4erORamDmoxCcKOX/z8Qir3EjY47P5IDFvSs3xPLj+Z17iXF683/rV
wQdKLIHAwGclTKFkvte2bCwHco0HoBD1GRNHb1gQawVMOOPYsGqIFGJPeb1ujEvU
l4RDs6V+8r6e6QJrzAr772rEkTJWhJf/JCn8bxJsuuPw7kXCzy00WAd6Hp4J9L5N
4s06jdctBqzrgG5dYHRoNvffvJ+tBlD+tWCkCt4R1m1sTaqqKAL9eAR9gxRO2YjF
Hw8XDfhkI6B8d2Y9UlJ7UbEDFCLcdsaElZ09wGXD0nWOtEE5exdKKOjnOEMSzfSG
5WhND8bF6XVH5yQpZhjPsWlSsZC70s/nTjj/a0ELmnY733kok9DeFRihDGVyRCRv
xzHUKBMXCRBecjoAhByxVn+IjSqxuAvRYTTcxvTZAlfYd/LUUfN6ihla9ZxCNRBt
L37OpfdhABKtya4+KBcl9KvEkYgi0JX+xVdK7giPGpFqr4dsWE8sv0mUXLHgyY+w
zY0DLzT8LqzvvyAcGGYPaFK9bdRtatdmuuSVNhMfEPUgSz9uNJ0kLeW+5jXcm/Ye
q9ZiUoH2AxdxCyRFvKtrYokvaLabuFEMSswWrTkTR/+1CH/mQLKHabyp9u/frFrP
0M570Wgfvh/KKLmtmwiyWGqb46eWFWTG9iyu8u/QVW8WCjtdCzN8I/GF8ZYL/9YD
Vtfmsc4HTjJHG/2A09zMU/nVy4h91FoT2PSs7w35gRzaRYjzQZ4KjYZW1Z4D9mXv
ffasPp2kzpjIPTshgwfCFazdGDksQe2ojxaVUlA8S9HxlwwAu+GHjT9RIENyMHUl
87xpD5gF2XIP4lYnfnsJ6/5DTUzTfytlJ1bqL/n7IL7rrCfYmx3+KS6rGfMez0fs
Sq1thpIioLcw0UCX9v0Vc+YrvnsLVz3PhCeu9f26Kk2E5xyf2tcG/FmaSo4junbK
4WcOevhi8U7X7V4Z/8LPtCLaogGbMPcLPKMFQcXG4kKtqAqsk7xftx7Ej5D6wDV8
PGLCwpCi1aJ96zA5iLirVj29OENLlkVEB4VUu67R2uyDzsrY0W8R+NCflAq++zfb
IUT2yEsfD60X1Moq/9OvadyvhLH/BS2+Cr/7IMSAgZNWKc4kCeY/hhAkH6WxV1DD
exb3Ii4eXuILdU4LC0XWQuxZH4nyzCyrt/QZR1oWSnxIOYTcFFRbuDs2nFC609S0
9nOJa6cNjZjxsNEYEwJ9TFhk0sYIwVkG1jTer4W+MZS67MImHqORf2BFYImIPS4J
cN9GX4phnvVGbuQxLnXhOXyEHda092qna0ULp4vQuNtoximbLzliMa/9qXd+vtXQ
O1+cM83iZ7DKC5n4xKnoai5YVW/Ot/Fna36wwUSIVdd7ZTN+QsvsDDYHJ6KxVDFc
BPqqsJqm2PP0LubdVfg1Jzwrx49WS/yBOmULVmfDZ9BO7VS310YdjPP+tzbIcr+E
808GfykFPV34v7VUr7mQczh/+hJuU3UWGxBdJgYj5w1HMl9DzWwDvsHYqOQqiTD4
nnhfooL4FUOwqq8iMbtz4erQj5/fo979NtEw2eZcske7sRWjLWaFBlwdhyl4WM0h
Tyi5LLMbX4EtobRxEUNzplCC82PXCCprENSUPODAdWeXYEwxGX2EpEsVVlxGcE8a
wtVpLb4unFNutktwINKgZWjEjKjjknj0rgaV36WnZRn/5ABbY0FbPfNs/MHnKBx3
mTCHGd0pAfD5s4Jy+oZp8AGkom7W60Lj3bcMmbqdBP105fqq9d2+tkPwHHJzBQFs
IOwC1z8+RI9F9TZ5wzVUrE5p3zdeOrZsPIw6k912JiWVqlyiAOVY+EHGbyixM6WA
dtySIZureZIBJv+licLTJMCs1USCW2iuRCfv+DugokkX/ukSOl+HSWV4minfs1Bn
QcKBJM4VZU6OmnsLVwArt2NCMtwgKz1sTT6Yq3TKIzvlsT2C4StbStYBI+HONLBu
DjDl7bdbbpqOenL3i/4VyvI/RHGukxbb63HJ/Ea6/ukUMUf3YupxYwmRw7bBkDdh
D+m+LCLQ1mOeF+y6P6z3wsuSVAzsjigGvRGkVypCppH26n+5EtpVGqqfRYmVKsmV
FRjHMDXzuqp/9GGl+Sn5c/T/Q+OoT+gwmP3s0yF9fgDf2+Th8yyudB+dAMmv/T0N
xFskK3nShuG909xl87SXi8yudTKpFP/3AxacpwDnKoQ9IL8CHneThhmBMSiZ27Xf
I3Ha55qO4pfqecovhiEjghoqtzw7ipFfYoyk/kWIF8qZt92MDy0s9aXjqB16KpiK
cG9OGqy4JG752WvR9UPTrOzz8o3m+kkigzlavUbBXgyiywdZ29e2H+MyCro3yWQm
E5ZBdn6Rq1elHbJfETIxDvoEYrYal5z5mZUJSKHMVfh2NkrfxGOrZZhImAXgP4J5
HtoEXrsBLtfAgM6FadN3p1y6YjIbco+ZBpQsCqcwC1gSG0tp6DYJK0A8Avr9AHEW
tPjuDvKHDVr0PW4V3a6L+IqKSTdnhHXTGBCN95/Z71Q3yT3jcZ6YvEClSb52JWzP
6R8dWKGbrgtQPG1WR/hINZrT5RQrWwpIvRBl/ZyBD1CCwtyXH6feh9JBLJsNFjIv
Ay3iyuf3vciLUK8ljanAQtQuA2lpINtSWOMDsM4Ax0qjjicSw7XbnRpes8fqoXOu
/DZ+hpszxhZdqLTa9LM7kN3fNOmShAajXxVoksLC69u63lTBh29lUaxNZ04o/tRN
+jqKAcmfX6OXWcx5dBIHUFbyV8d9C+wCSe4bIUsual8mBft8lc0ipf6LvmPvRSEh
z6jfT6kJpVULprsRlpOW/U1wEus/MhkE1Ait/RSLGx6jhQNV4FwbuE2zIlGf1Px4
bnR3CkotHGoTppHz95gggVVVAVkDMDwoIhOCMbaUhLjLz4YaBe27HcV80cJ0WGdB
uvpwKDg2eBgbHnmYgLFOykB2GqfpmiLqkTWoxeTlHeNMXnu2+xhI2c8AlyWzjDKN
XeVuXY7tviMH+AU89X+yqEinXiQWgDxW+wo2qBWPK/O7Gr4jtQYLVg02M1pvIXez
KVzpi+jUxjd1eeoAr0Yjay0rzlMBhARn33FxCgNMhLj+93Vs4WPhtuDfW7aefRZv
p8PPEMe8XBAhBlTKgzgSb9iMcVX2Z/XlEsSFtaZLqqXEkPB5UMYHYLiIei11buWE
bI3b7HS76RPNdmtZsA3B2umwSq8mgI6KD/sDpeRVf0lofBxPUPFjFrcHC5tytx3m
+4RiS4CaxIuDFQgtiaA9yb1Wgf9CqphYI+w8VMtlLqs7GE7OgaTWdZ9W9lr3yC4N
XWYzetWu0BiPj8nFCdbjMQiuuDW34/GmivQ2tOT2iKREWyGTnTNeW+3h9ObjqKM9
QzDcGYXE5VaYbfjJ9koo8WXGgrNs0mb2dkhcjT1y94TpyluyLm1iT+OMxflLUmTn
t9QaohgQHhUYsqE6O0RKt19ZzSuwKhvt5zPWR76ERMVfCs+rT5EaDAK9sAV0OdUh
KWaAhdVndzIEwXQ9Zo3x4ke2NmR6LterYEbLtN1QO2aQ+LqmGzLZvS9sIzoD/3zM
4LbuMhKQCnHFrDFbPH0WKix8t+zGWpQpDNTTbnWa9EA32jb6KRWZllW3A5GyNElz
Lz/PXB1BErszdPzIwCPnw4MKTX66hBp5n7R6PWU1SdTL/e42d3Jio9sp+hAmiBqj
9flwYhij4Bz+PhJvwtqDSgovgxQwXGkLAz382Mo/8E6iUrr5Ar597B7rM1iKDVm0
CC9IyV/UgJYeTRyqTfIq4vsb1qLFhJPzZktOBWlVyNA7FOXz/ZvYlM+55sls19yx
jKsNQc7b2a9TQ6SOdJNGWu/xhZ/xVQESed9IYYozO92kVyDgLlhXLnSiZfD73D7u
ySEoFlwul2NrX2pI0QMTElVwjgqgWG1fqD8AbfmKRiORsZ9LABTCPp5Z0kH7omwa
xS1ZuLHiYNpmOdFdvhuIA5pEs1BXnJ6EVaC8VSpkefuaW+VUJAt4/gxieBoasqWs
sPu8Xd9ioaJ+rIdIMVQWqLb5n669RaRlClQgamK7zNvBBKtt4ta1otyI5lCWTEC0
65FiOlt57yL4Dwn7LXENmP1xCHbsWpnlKSEv3e9om9vsnIJNSxkR6MfD9FbCbrXh
u4PfGoOf3o5+lo2uVTp0wQUsBl9K3YL5izCWDkCg+ybdIAhKF25wYgErpp0A5p/j
2y3YbU5t3ryPpx4nnThBaY01BjzzJ7rje/7BGOZmxyejlQgSFycCSnHF3JODWtsF
BpkNuE6+3JcxlWEnpPxujMuPoo4C8ZoNtnB86em1s/QU91LEOfcp0iP5Zy0qSDbh
IrkW/rONtPgOM7G/cBnmFz1oNq371kIHUfeh4httgnzjQeJ1ZpG9yb0fF+B1kgNP
lDpNGrOdUQSHhGRXpVwtg8QG71LzfELAvB8IiEfxo9IAnScCNt/gcVQj71Ui+oVr
xgk0n1nXrG6BRGFOAfBK+PEj9BfbZ+5+h5qle1gCqN+nx/ZuczLRHXYm/wUCZR1h
wWr5P2N17HDIc8OCPA/ZvXSC22fMZ7INa72J4dyCyeoBt8gDe377jx9ZKiHHiP/7
NE9vtgxWgWZkyakGe5+/tf+IQ6OgbamIS7GMB1FRKGK0SAo9tTdjvukmoc1EYaCN
2mMWOVLQsMITzUZn65zJnQJhDPD0MK1UFbVNz1CKTQSKntVH/j4kvSjdyVBJk1M6
RmwgzX/S4WzYe6wHrX8N8OxHW7KqJBYELdlJ4mHEuXDnrSr3ddWTIuBiGaed6yO8
xkImWwZQ+OwvAj8GmCPLgcwwUb5eE+AwQZLZZNjmH0IXF2ZEyyKWp/yFz4HwxlhA
mLsTz+A5ZRsfNUwSGojF56P4Vsjz49BsxnHEecdPpa51g/7Mz9xKYBDGou6P3Dh5
R20wJlQanydHCHFpVVeBkbRqhUwu2uszPhL1bvkcedadr16z/z4TmIx/Tl1oPJCB
5ly8FvItMlYWgpI2M90ecYJh3ANHTMJDzAtBndnI+YjzxW+X6vmpMx2TFhxdaeDW
Vxe8eSN/viwe9TmPaekrC3ow96xIHbnwgq4V9Hipf0mQOj5Qxy74+x+OuyovvBVb
lJSsC+PsII3ZpTV6nlQa22eb2reh99dXG9/Rvrkg9UOxj2LITo9e2irOZVMEVDwO
lhjja1IPC0mjbmrmhBNLw5Qk26y9Xru0ugGfI9ScaNrXeNu7N64o5BAKMxOEiTe+
T2UtfZlNsqE23gs/+dYJGAJ4HHWBX9bUlMfdoXH4qRpmBRVhl3D5vK4rOHQuH1WI
d1OnXpGJHwF6NhsNFT001k0g4FiR9rvaG2rqn5LjQldyWj3rGiK0Uai2EMjDv+9X
++K/eRwfzazmGr35oFXbksdTNYVqUALmfRBCVySrdjx/WWZP+KneX/BzRhOi22O7
LAtU0LIlN4vzfqPKvghIaPiMkWfvMsgLG5VqTsFvRvEBWCK9nsUPJAuwuEzZhvgx
lP30YxbPFH0MvKk06gqdQbfA0Lkeao6gBk1fs5VEweTROs8AwK/4yvTHd02VQLhl
s0Agb8KkT/b2btqBGCAkXGxcASJSTAFqopn2qWrdAdaTHg41O1s8/TNbSJSfvRgC
CAqPLgZDkwNBQ0ejqMHJtM+yGoncrAmhWD8HdoQ4/nDq3ebt2KR5RFyBwz1XLc/z
bxOTIIzG8+HokxTT2k1R+nCgZGaWkMfway1EYfeIfBOBpQyecwVWOB5MAPks+76W
rT6l8MzFpEkZpOVkvYekj9xCcWTcJEqBatYhKVzA7RyubaGznGpt7HArqmPjewko
R5UoR4uua84+vRyXAy/DLA56swmZ0o6NYsc6cPlL78bNOrn7vB4cALLNAUmsHxg3
K3h15o3gRRukkgggKwZOcD24PHfOycOqRyV63suKYvtnX2pPbTcZQ/49o/ijzVCO
dsXTZOoHi16J25O/W5CsU1wqHIg+SmZBG8E6EIsgyNet2aMXI42XkmovrjlLBEwp
z7K05wCqISpKylzLypzrdOSr3aL9ePXSDdP4fHlJa30zRaKCzHPwESFGBxRs59er
IHcj2/xrTQiGpugWuHHiC2eEuqJewFqbXOj2+0dhJGtXXAgvPiqwBIQaRhCSzVjw
KHmc3CpQWdzcS39VmXt6dTRNxpRwHCEjZncSA7a2O3Msb2UF7vqdEr+wzTRtEbrr
vd26h246b/fY+9pH5eI4QAIPArjxeSRLjJyj4HER1K0lZ2NggJt4ojYA8t/MK3Zc
mnWV7bumBs7Huhg8Yhv807pUIBWen4lG+pLlMc/QmtwSCaLtwk8vaiiApOK53kws
4Su8ABiYGWiFT861jtez0MlGUWSzN5IYvPdyPuH6qusOLofKhV6zf654ZOd7cell
qgKN0WXaU2FR2qSUHpunVv+ur2nSCloKTT0/UgZn1Xfo3/L4r3eII5W2cMdakkXb
RWtTP4PRzSPo9xPX3GtqqyhSixQHQBecxVzJA+Kga2cMWvtH9AAWZlNWi9zr5DqJ
N9kLtCYA2eV3Ye052KUEbseW4p+2WjZ71F2raVaHVAF9KtiQ/IWB3OF3QmQE7qIJ
I+DrSEufjUWH0G98hHnBkvmzckyiY2pnLngXDg3pxXWuHhLGArSKAWJKHEJlhbEG
o//4duJTFHMI9HsVTQFfjxdlVa003Gr6clU1Ek7glObktvqtYFqIaMkXWYU/bVL9
RKvhFR5jQHEfOntxoOpljpovvVN9D1UZ8thmKblCwgjf01Jp/3Tw6at4qcYSoLXB
0LXhUi5yssv58LKC5FRsovJEZoPZVT9rCcFwR9vMyvhv1fNzJZ2bTOOiQNpolome
FJeDYfm7hFbNxD7MetVTAadXwhGc/s6G5SlNXXQ+U9zbh1FC+CHMFM22OTvH1rbT
RWpZnkFDcfpaK0AtUv67NBrSMIT8ZTJrXYRJ3V4He7XwQOQGVBDLaQGtBDZ1POiM
U1RL5N5Hd6ex5e1BXHGA22/oJ6cmTwSnJnsSB6mqrvYUVZwoifdSbtePoOPmzEcj
8dCU/wryJxDJMvRgycg/dGQzQVMTOnNuQIVlaPvMUPUzKZAounfo4o4Fh6esNywG
GIITPD8iR6uGPLc4Wc8Kx/5SwVqMax8gq+7q9H0re2TleQMlcmali7q/1fh9T5Ho
5wPJEgJj/hmI9rLY9wiAAwXLJUb6ZWKeFmnc3V6ET7DMcj9/F0DHIKeEb6ws+Xba
q3RZzCWm9tjo2PKEHKGrJ2/fAG2P+qhfpBySaSKPyFz+nmR1w8ZEF7O8acHa4YjB
cwNFz7kvMWjdwxSSiUC6yHRhZZf35II8XfpgbIUIEpTR55GeQ/tIoqPo53gjjopZ
qehd0Sh8ya/SAEnO0t7eLoPWbHYeesmWAUx0LrLUZR1KJk74pkNYXbsogv26gQS0
v4+DRXbapINuVPCJi2RBBamGVce90OiIyMOnxLhYAnlbjoNMYeNIruoqbH1K21UH
+Ai4YOCn872NRGp9Rkj+dR+5RbmyrycWCIrqph2P1vYLWULxNWqcgVnEHyE4A7o5
lfi7jGDNf51ovG5hcUtgozwiIH9qsqWzusKdgncbnx1AtbBCghD81PyWjo/E/5wO
MjJiwU6wcXo1yiX0GJlG3N2KAHivjd7qW/g1Af0nIz8rCpItMFc5VfXJj57z+ClB
t4lyVTZnOpOW9Jq/v6TamPMeASmhtbz4qjXBkCCq4qxcleHJRg/AmTkhLmIKeEfg
LoxjYoxAxYYYGWUAQ/Zedr2Kk0Kv7SQCEG7eJPeWkhIqexj34sfnnYQfkDX+y8BZ
BJDhlLx46Ol7riqmJdnq1GP3pGcwi0RPgs9Z9wycvAYyFP+DhxzQnzUq9RRDFeLS
yc7K/0cYIEUQcT+UBUZK8QhoF2gJgIvqgfE0uH1kbkA8zgTE47fEM/e2s2+AuIB7
8fhJhKLfRUPRw9SEAc+5rJuKMsb9+rodlWn2Bg5Gnp6pSGD1aUIflNhZdmKIFzpB
X09z3SV4JJuvB6Jp0l0Fxq+MoGBA8+XSw4Zeg17kxgIQnf7187WzKqR3H2CxlHqk
dkNLziBqbS6u+A207L2s9auV6eG1LJIwGCn/CLufntX1GqZQxANDGFXdK3QpURV6
9gacfai420daieXKNP3a5x7V9N2Vxtm33z7io8UOSKjLBxMR2D7bybnzaGrlgvum
CnmxDgFDUDgzf2zEfOrjTLXQ3C7ew0XOkExFU7ytRLNWnw2LY+T07djrc3gnthQC
/76XsDpYMT7uvkrUICZjCSTY0PJbe7GQAzEEx64wKSjlKzdYb/c/n5jsQpqVHMNE
+JAvvYoFObMm4FHWLwH7vqKDnyK3Tw6Fu9KG9XYCUq8XLi17Cl6cX19E+cxwkxYG
J7MN6I8d7h7qO/b1tz5TaO/hrfFr6cYmegxgPr6IJ6J1cI7LfoygaZoBmcWyUM2W
AsqdW38nof4NfJ46+pq4g9k2XC9wLfZ/y4f8lh2r7yu3NEavGPxnUlDuFtpBZNnw
WRMmxhTZjArjRn7QgZZBPMDQ8Gj0sXOnYSlrnT9xlzGLsJ+6ZdDqcXAsNBZy+onA
FeOG/meC0A6cYSLzrldjYgtm6xYUr4kz3wcLkweHPnWOzORFapC2hXQVWOgQ/aSq
Qa4R4xrwi9DSh8jsCa/m4z7ekUoo+BVAoHCv2qqyFBreNB0DxiVZeZ9Rbq03DnJg
fCA3EeWth28N/00HrugtWZZwH2eGil/+j2dAFgsM4hjY9mN7uNhgYtG4qpPWaHFJ
GSdKl7s04VQwx4/rCKl9/ZCbz/UR3Qmt1c7ldb9UB2PlmyMUfyISzXRj75grXXeT
0GGG9xC12qSn6OV6YVz0pS5qmYXk2RFXGOAmjvJLlVR3+0UYSQHLtSyv9lyyRASE
KNm0tIOPtv6I7X7c+8HaoDI/0I69hAMqDEhvLZlJDK8NVYQTr506xeFZK2c3Mqw0
kYyRaGbps0dkWJr7v0mBbZvpHh5igX8NcnNuQbds39Ziv+A4K8WRQyaeaE25tdDe
J2F9wsAm6nMtfpy7EEfUhu+EagBU/pKsvrcNnHgLpKidDJRSxrJa7l2A86ay8qKy
M3BU17MEpFo0IpgzB1wmkjG1q4zGTgg7KhAyvCKNObe+ko5JXf7NYoMmgJHS60Jz
Nv3VtUBbjoZMOBXmAnZstt5YbRlFUvOPRbbFPRPPZIgRWlOkgtQ0B1Vh9U+U4MTB
BGTM+AG8oU6kC0PSJplW4BgpgnbnisMIVuxDjclGyECxYkoEmBe+dZI7ztC3Cy1+
0CD+euVexJm0awowvopePTUmuH1p6dl+yZj82PW83Gi1LdcVkFUpA+4LKB5kL3v8
flwlqKu+hyC5w9Po8SPhYsUWXXLAuQKVxKZB3DBTAAMQtmc+0gs1qNbI5svyRMJb
JeR3H1to/x4yqu50h1T3GzrWUwiK0sL0pX+APXKiG6rpPKtdnGoMuW2T9Q+5l4Ej
zaTehxECgVx0tuNz3777kFJjOKDc/TknPLOIPMuLvTSpKjRKAPczH0PcelqRq3vV
s7MIdLxrGQbQoZba3UAvDYxvQfPX9P7tM+IXP3wp6UGcoKvS1e+ZTkyVgwwNoiM6
G+G75QUXgj9/tituB8i4XnZGajFunDb4txthAv3Rdu7lM2KDi+4HlfwHs8/fk8+M
gTXJP4l5V8kfZksAciQ8tXj8iXfyLaxfvObxDoLQspO6WWHXAEfviSczxsQ+QQMu
vlEs1kM26WxaGuVwRpPHrTXKmnSWJFQfoPggxwDDR4TkLKj1aIvP2JNKLK6HuoUR
5jTcZ7nZRReLV0iXLHVyQpHgtQPi7ULL0ekUvL0QLH0pvc79Pm0z0Yj5OwEGkn26
g4PXRstpddSeMHbNL/y5yJ39PIewtgYJTmaq09WAcUmm/VZnI6hoQnuciLLZpnQw
CREn8zaszT1KQexihsbmS7mQ1kTSrFJG9uPoXmVb35Ovbhc9orSNLDe+gN1gFW1M
x4w/iD7+hOXdeTn2ccyAE+pBmkfUCIHeP205QFsRB5pwyCZZ8rbRu+uyg/Trrzxf
c1EcnHN9UsMtCRmK2arrXmpjwaiKF1cm9kr/FJd4NvCzjD1g4TW0e38VKjAuMRsf
BYCFFnKpp+4q5HmzMmCZHvfaGNmo/u7N6hKDDzVdysHrFkP/WV7rrYIfUxBlRteH
7WrAqUKyBweR88+jikEcLRPBzrRWtdP3OXBRb+8L/kpJwKqhfteP1h8cYxOYQWYA
kbltQzwwdEtYD33WIVIX7f8uQj1jIhbjJjs5JpKeyzFq2T05Yn+WGz0lKt90HAc3
BC6inClFaG9REgsseOd7ERXZqJxP9qrJ9yWaxnJD36dqgHSfKxgr1oAY3cZN3K9A
rmetam5r+QMx5ZiWS7hL120y7z1/pa61PipVgxzBy4sEnWHV5icf4oiXbR4TbsTa
r2KyzW5Oh+DTa4638xW9/gJ9iIISpyF/AC76n2falNwGG6E5FF/6UhsM7EhD24Sx
irMr4a76nvKp/35r0wuOW4B+zHEvUI7Ry2GnermyI2VrzuZdJKOtzPHkiV7U+Eub
OXdQh68CkD/yHw1wEqA1sC7jtN6EJ2gnLoUJQ+NIkq/+SiXkh2qc8J1jlV+zgnD3
DYv1O8jO5ZMBJHdMrCNr308QNOZBGqFFgYbArQA1WE3euEoOhw/V/+yi3QewFREK
bu6mAYlIKg8NDnPzsEP76oMDiAUWyhPiVAJSYvz98FrFWCfIs5B74n4ZTo/P+ql8
SXdHO+TGpVV7/c0wapWoSBwuAKpy1gk8vm8UIVKfoVVrlmw83zMoHaEyzZM1Jnll
B9dCLU+DkgUKzryrRJ+S5fqEL7VzEkrNXCYpeHGddqcjTzHMtQPgc1fJzxzGMzsD
HISoCt+9zOIaKlw2iyYVJ2ZOnBoRK1Sn1S7i7MVD9X39RtGWRb0mibxmlK7BO+jM
QgMgIJXz2T47LyoAQ9YvLEvcKWxVKml3api5VvehOX2iBp68hGaYD1AQT93TcXeV
0jOXvNynD/KmiD3/DvEujykeSwm07uHJ53VzOPrNTrerFrtWV7VCT7s/yGBTVFd7
Yzu/2Iy7NVZT5Yc4TvYfhpIeqwpB+ylUC2Nb48xIRR/43r2k2Ry8RZpBNerMyfWh
KjRNDuG0YfwLU33QuazzLQQRgJ+qYNAX+hbpN1rqXW9qO3IiNhpkhrUAhxxqKMrG
xjnQi/YqEKEYFXecEkz/LmZQ52OIwe5Bv55JULwotEnfXAITxuXawsF6Pxl9CDMn
8WkoUfm0gEBlqx1mua1Yiokw0l8XFBpeFvWnbYMDQJ+kKe1sFn1hzfutxfyVoMZG
hC4tDbh7X5bMkqnp5ukeuC9OPRBE6ZtPR40zkE2XRZU+EESqLSWjJC6MwlLtYGSQ
vH5dHQfZl/9ypXffrtsBh2ivMn1us4Df+CAzC9CFbBBicdPC3HOS1b96aMe25hWf
t8e101GhC3dR8764jkF6otI6ZrxhNNzWpZTf0Kd/y9b7c8/Vusf7vKN4rOp3JjOB
lszHf1YUfPhTnoaV5lQENx40/YFmIlNoL1e8lQ4qGf8UL5Z6ZGfPO5A+hn3N8Srw
WnW9pI5FYSEFhUDJG1BNS10KbiscZeMbPed3e+NcxGmMppptwRQL9LnrqjPtublS
OA2ilYUxS8bmLimduDra0H8n1q7gDJ1DyYaaZJr9rbTc1tg1scg7AV66ryz81WbG
o71AnUePMxXbSDDt6QEW8Mnst0puEl79903el+HaviGjieVSd0YBsGJe7qGaqDyz
aLj5jbpWOlIlfRblSBBrZrPGZgzvGylyGSCGJQFnSta02+wdReW+gjBIGJ3ex6/k
v6ZOV/0QTb0Wa8njZdId4hzZqxx7cMph1uT1Csh6yqt7RnxfraQEK58328GJhsyw
9AMo7zOqLHsjcxT9Ya1U4GosFWiOHyoO2+RiWzve/wr+Aiso75pc+ya5YmPvHILr
JeE1WdQecQGsK5n/rlfkzqVw7YxZiSAxYrPkXZvkG2ZnsJBa1HCt9YBbdJnY2wJJ
sY6cW/RDqtC6lSIrIJ1UgkQPYoJVe+2cCdKG7ejQ7jSImHjtjXC6b81CywX2EbyF
1ph9yJmPiYp8Lyn1qfjDBKTabKx4ntPvr1eXZ7FaPuV15d1VdALNeUkm4C4upLL8
3R6ej+G+f5KB/xEIN5rOhqWmENVsJvcOCj1mZOnM6mGtsgfqvIlM4WnmPpKrB7st
UgbHbU+08iq/kGAHTQshjEt3zR798YedJJxac4iSky+fLJa31084U1B3WDiVIX0W
QijAwTLnXWrqJ/y7N0AHxoILL5zWb9LAcuFyqq5ULG1scWIMn0767GmGYp4hLqW1
VWKP0fxN2gMAV/iNpsP+bQc5XB22TaQNfwLPGyJeKxFgYKu/Vd+GfpCwDqDMGkhw
4KK8wXBbeZO541WxVcdi14cwWcsNgWEmQqLZyxQpOuHAIPOGVUWzFSO1Ry2xelQV
+3S+slsILqIQ3JmUtSrACxQ6LL3Rj3yhd4gV8phE0C532x1r1iUXaL8liqfkyZzu
nBKnKFMtqwFkSAGnnk8GkXConQF+h4dgvq5V8XkOnadw2Cl9OL/mrQYGZtGvLvcL
V16+Ho4aXG10PATbYbcvDGktJAA0TMbRXy+p6TPIzl6NtOyCPT2qkp4yTNxyJcE8
ljLwvG2AL1aeuC0kZ7w/UWbNEXHS4VHCKgqVaZ1nSfFbJHwUQaIWODYnrXcn2FXI
i2ftGrwoMjmBti8CrgV9n89vGFNX3H6vl72zldDk18197+Waq8vV6to59DPOR4rh
cDXFB84GlLeeP4TOCjdUEJH+/kKbyJyHW+kQsR33j3oh21LuDMOrD72cCFp19MMC
ZZudqCVkbA3h1P+tnBk/Yn4U+wpbdhvPde4dWRqfFeXuVempAXbwimFOD2L6MRo7
b/Daz1jda41LJX3Mp8Y5aIWa4XcQteAZpAs+OxMqdIRedXoXdz0ZBODcLVOQBYVy
3Kb1Maf2C8qjSKCbhipn2VxNzmZf1gJsuqNE2rywcMPFoyZOQ4wnPdX9TUymxY8d
FemipZA3xfhD4kE9mhQYzaAN/F3YIDMaTr0tUBNay6sGjUkO92ZFcKd0DSqktyFE
PFQRWfZKT9Vw/NQbqdUXguqJYVBTVQip+SwzU9nt1/1PJlIF4GJl6kO/xr58WIKr
7/K1ZehRMs/aerdo2ZEkhzKQ3V8rnmmd5M4HKGB+OoqQWJqXqEcs0LRijGtGALip
R8INEzCgOa4COJcwggjR0jDenSQIbl2Ai97zYrb3dMKrNFDrF1JyCALTfHcr5+ko
o78P07qFlvuA91t9Oo613vBf3ZMHaHeK+mGTDWc2AeZXIZkdEr+gxg1vMoaaLy7I
1IePgPCYOOti3mwV5v4YBvgWLPkxLUDHRK3irX35gxg+MAuXxWzZKJMJ3Jo2vb0H
bbgU410ZWZsePXnzbMfHYI0HDj70YAko2ySaAx+ll2vWnScQVG2F3jKt5eMV6G8w
fpGpDecnCwlVvrdmfpIzQcz2ey2kh09TcmDJmzFGzB7YtAaH+79StO5mEf9+IplE
9pY7VJYDB4CocPkAw5A6AXJF4N6Pr6pr/r7eTuYYFUQqFZz17yxBUxIMmRvol+Is
SddK9uwtJDk3srZl/FRnVLRL5LIND4YBD2Y+l4ghwKcvQDvA0dZ/BOzH+133Jukx
6+DEwnZOcoWrgkSX0UWjimCRsZYiuTicVHUpAU1I/Wk7yz+ofGFdMEC7kfusaAKT
cb2CiJzZv+Veevb+9Qt8Hb0fcZaKoDcOS311wTpyFxBRi4/tJL1IPMtrJPct4Mpw
sxxjbUBen+oBo8cIpOAHwisC8sjFNMvX6y7ziV8x+ImRmtbCuMNpGgloUvPZr29u
5VsZ5gdJijtIxYDWdqRyyT1WBuQ6O/1nHQqjuoiYm7dMm66D/KRQNP0tXtlX4wpO
K2EmaOx1uZ9G+VdH4ZO6MHYSDPeY8+uQ1vVGdq7qnlvJqP5XY5mqokbt/f+No6Uk
5ws2mCZPUkKAiU5HaBIm9fWwAM46PNlVAJNLIw6gjMBjwg6Q2ro/I5YjBlUt9qVX
k9ITyzImVCArKxe0OzF31+Xb/ILFsYie5qPInwiovz73Ux2FAR0znXYGwJm1zX1b
NwoH4QM4j0PrzBipW+rPON1MiwqOOVCm0v4Lqdnk0XQ+YoOv703uTz83REUOMLvK
0idMvdA/pBdSkCNCHmFRlCdFFk5E3Cj3f8OnkPz1vd8p/Itn960HjNulgNoHqwP7
HMeOUH9xvX6mX5TywDu1yU32tEyFJSbVmNhgZnwayXDDqvMlKBW1eo6jHgpnNghU
6Iwa+vJzbvopm3esHeeMhKUxxcq0jm6+zMR/Bo7Sgursgdong0mq1aEMrJUDFpp+
vVxO0/X6Yij206WrNTk10cN6bj1OPxvgsJMe57z1P1oPgRItbTvuI5prsJwf8eJ7
aq/7RiEtUYCDZw0RYvEXz8/cBqusB037pAdTLXjcPlJKqZFhymnlAPCBaGpHEM8p
l4kk12VzaUNfihhLXhlswnjJzBkn6Rxc9i24bsbEVyjdJ322ZpPdX7frl4Rv/t4Y
4g0uwsPoaA4w+iEoYpWn8iit0mRugsromLG57hunKr+fKEPs7WVM0taCIPABB1cA
aKOUrkdNe1GYVDIYZ1wdZZO2bVVzkV7zAygIA4LZCFUqA++7Yuk9sS+eFW9gCahK
X7DfSJeGpcaUFIo5JPvgCUdi38zFpyqwMePz9W8CkX+IcZ+iblEU4L1Obaq4ujCU
/3CXKmzLtku+FYyCsVKC5JfftJekjsW7HMa31E2GWS0T/YK0mUnGsT+2yWhGlx67
Y1lkI4WzIO2QyBigAzJ5d2+9xquqdcZntaigfkQCSceSyCiBQW9+J0uR4CZUP4JP
RGWgMW1/pCUCX1mwqQ7aySFcwCP1N5LVM5kqBXCh8E0u0U3siz85zsn29G+LfcPX
UJzRCh8qV75vyzbIzH7GQRgMvQzii2NlmFJgQpBFczlaTLhRLQ8zqT0XGvWES+j9
A+zxHI71xj+jMepaBefjdYWSbwQ7WBJuaOrIOvqVvphGw1d0ooy7Hf/jCefUmFR4
F0qwKV5ORKU8fUclaIMNJzvhtuMeJta3drWESENXHO+kFDSfGkmbICxsVKAJ3ZMo
0aVIJmlm8/sVbof4IRRYnR+o5DbqT0DuDwqSWhczc8ZLBGuTVWsmm4wYF855bzxa
H5IsUgxmp4sefwcgQ5Vq3iwTElIUMmeAnhQNUV3enUO+HTBVXM8Ln3dOcVh5BUio
Kg3Tm3A5hdIYAjJGBLyXGplQp8neJ68eSgFzjxZsWfm9wUjdZ8w5HYL77T1uLKDK
Sx2Dli7/mEkQA1152ERvFgeALGRx19o9iQJOUiMAKakhxYO8ynxexS/DPfij0RiA
mQ6r+DcsgetfRJh6STBLvxXkMYKBXfpXfzrqVx964y5Lg7RptOagazbTXwHKzFZo
XMapIKw2iWK0fWyqYbdUvhm2kSsRy5R6fxOArSLtA2ZQOhqgDllysTQLnSVcvf7e
J8gTsFVGEdBCYdmnWhUUtLptJK5lkgY7HfMD85FhRCzI7NKtidn36fOOv/M/XpxY
bLydL411+9QtAzmOAZahWJD8Jm1vmlnHRzWymlUATb/WABTJ7T51hqKUZKHRCFN0
fUNVXJpfa9rQp288lG7PLQfKaZ//TDT2ytGK6YbOzhANa0ZixXEZFctaekQvhZnW
ad95TLzTjQ7KOKESH3JHSAeJHZELwPKxa6+FlPWzBBlLUDvg4rQlgNS7OhFHDsfn
6HIjtDMWtwGsWAc99BLkuLh3hBzeEknMEkXtGthFrg7Syrv0yzZiuBXFHKlRDzBQ
XkyswdGYKS5FKM80pNv/7Bk3AjRhv6HfLsdO3G65NNUkpDfxeYHLpsYA3xYIr8BI
rDN8CYmeOj/zUbO3eeNg/Uqb90uZBMQttBWc/ls1bg0i/UH7XJD//0xPr05L9d9J
GI+L0hbnbfS/DlalJqp9TCilNFj+mbIDuruM7RqfvnOLAmoFOzXt8GbLiifqPKeK
kUk4cllauuzYbNi1BhnCc8AUv5AOC3lpcY4MFFoAYwoO35WVi1KYKYqa49232nz+
+60SaCwU1/2LBAov13kGIOA8LfZcr4G7qzP7CVp9AujL8ElXuzwVrFi0NU7UJpDz
0lyOL+9xYdRDMo1l+2+1kiNOOvz/P9qHMEnb1cJW6fXYcHdTZ3Hswu5uceKFDtse
/CSFc77vJAU//9NF6VZQe3BRVqxbilDaFpL8xpB+z4vBDbWl615TJDDNmtw0PC84
qflH+IfNuNiLD9c/5c+3SuZyHJifH6rFOyU98/EzA72rAhzyUdZwJoVIA6vJbxEy
qRnZ8eV5DOXHQN6qAqBEFltgZHofJg2TJ+i6p0ezbH1yzWs6TVJmOEX/ocHfAZ7t
CfjfPyfoT7KbO9dXDhu3Pjk99lUuN1RVYbxl7x8+jExMCOXDbGnJ7b1PbN5G1Q3j
xd/E45jS1cSC/jXFjflfZsY8LLms3owDO7K3aB1fzuBIJ90z4ozivuAaiBDG3rcX
1X3HK7FLdmjMaCLk9PKopvRZnuHvD3x9lGjbn/WxWPZyOrsnK73lR+cnVlP3jyEw
AefqiESvvlzPrXklald0H2JWz79WNdENt0f+iT1P9qLA7d6iqrca5vAzW6ZdSbvG
99eAYvPU7sBb0mdDDDs2lVS57i4cqXPss2bhYvhEiYpCdp2M2a1oXiTDLp49nCnu
X07bFzRNziQfdycrvohRqktqg65qf0LeTjmivQBKV/+nmYUEcr9kAMk7Qmgy8yuv
PDloqeYWIyr2GdCjqh5ZC8kUUe4q1txhRlEHpu6CmiyhrPXX0jaq8SAklu1I75rK
t1DZ3dKMDFt6IrcQ0/b6Mq5MHdaQ32utdl+KI2L341+8QLp2K1CzqaoKcHSijUhJ
fF4TdJ3pkJQkuD/opeGScQP34qxF2dFuOsfVIRHvwPynBDoJNqk8ov3LkjDQYKKL
XGiNPop1q3ftu+BgqQ6xn9uGUcj1miTK9w58UXRm2djIiiIGKwDVQgZ2DKLgb8qS
UlFm+ypyc14DPWAs1PWwTx2qtd2gk5tCuJ/L3tti3ln5dsddjF0DAMIZwKivNg7Y
DTrd5SaSLOMox4CfwuzpB3hHwn5iW4/HSaZ2wNQ9+ljBfEI0L+PqZwdt9uqcyPBW
T8xNHQdvRGv1Cu55WtGO2frlE3svpCgQVZWPZyNdIPgGJK36YR+hGZwtlscNy4NF
tucopuA/8HNVeUBtXBHr13X7QyzvIdzMZ9HHrnYebomJbxoFfMcxAfSRpwTB8Rxc
TEX+ZFNLzroyfM13cTGpDbabuWB1Ytc+uZhb1YGxzd7koExXklfte+WoQCaJGr3k
BT0J8OKujbZFouxds3SOdYJ/F4ivRwLYGvJA206Ms/2MIWb0uGQ2ETHy279yb6e0
EmZZrneq1R3A+5f2aRUM7eSMoFBZExlsEjvp1XfT6IOYbUKw3Rjscvca5GQcl74f
iTkk2jusN3rfa81ivvZ/dFcfJC9OC56Fg5ZDU2/77X4m1wNdpVgUFHWQZjcQPyT1
habfQTSSXmUpber6FQVKCGgOplzy7d/6ib/9vuudS4wGYz0t4wKGk0+yoHz3LZy9
x+ILe+P4F8m6AJPC02C/T9WqLvA6uJb+ikJe2Xv3d5MvAXDMnnA/oD3C1BxmBrT7
emtEOPjHNlLuA3Y9ko3UuZUne4Z0RwJpHBkTm0foFbDLJOUSOlgYmaKovkEUfiSv
7l4DYWMrzVbx6LadlT7Q8fmkAFmsqe2OZaj2RdltNbGFmdL9VRPVnvbgFi4RboRa
/p67ww6HXTAlcYqLwK3MOqVl1fd8wAkom043/yh4OopXjjKi8On66VX9LsLj8lhv
f/uli4+YCRjkxdCRSp0kzr4tyhuszRHnQN0O5kUe367Mml53MbJji7918bWkxXSm
tb1Pt0brah0hAmy2ItbIwnLjPKvHNqLvt4ul58+QVmb0uZD9ImgGt63y0sw1kb3U
N3ndROuNPB1A3nN5kaKq6bgLMKTSojzFQizMREcn+fw6vrZD/1wP3DGqBkDa0DjC
RIbG0o3jYVbYo0VoXVy3eR38qsDT/J6YlXwfs7eXcL1fsZGJb+y+M8SbQX72rGzc
qjfJxjWiKBvb/5cP9xFSVLqeErgszXxRXOF3t2z0caLXzz5wPeXV6gJOyqBFVhvQ
pKaUIYK9pxwp5tq/gptl7F4wdkZ39qlOsXC3bZ88FkjTpXhQyDnqoRfDX7vZthni
I7YJXOuGdXJHmfkWQ2JzytBMnU0wqi84wtFK5pcr/JLvVlXx0P8kxC4at7CBz8uL
m1jAMOt/z2icfoV177WZVc56LYMDiRykT32dupApraxHpEaXdAVF+lmbIOpFMl7F
3+PptYOx9SDz3XPjZwi1L0m3IA7+5Ms5XPA3UH/PR94/FlSRQ3qq/kkrg90ID1i6
CDDVSUG4yO88aoi1xSLiFpONfu1MNYYT+GKR8vMdf37HE780nP5hEAAR/8xvoJqs
lj8/f/buRoWs76XHL46sCL91s1xP/LYCYLHcpj0IHW5fp9txzGT98H6oHxTZo4F9
7BG7B52/plIGj5BtvbBbUy4X9/3pqEHnm+cTLyuO0Y9u67O74rxI65sz5j9OiKnG
0ORbqXdf+kPGFRdj/9lLDgQArxvUAFKNVfeR4txZbpK2+BWoHrJCtj0JQtWnU18t
atELoyxXMphMfqsRKEgq7cnS8tI5pzX0KDZWDbmJNNzmOZ3h57XU29rn1+MTKJEj
kpxBIYecpi50pvdOMOoltiyERP8s7QflfNlWbZJYVTeHOO3/JS4dyEmRLys567wD
na8gQAaPa5PvPv4IJccv5LpIJqn4GKkIzOhwr/KOJyz/mq23kW9zak4wK4zZOc2u
pN9m1oi6Mz77YVLdZJrcnXgwJUOXyeiTdC2lLpNX0McUyO86K6y8mrs+KJk+mB7/
mVc875Y1o9Y8aSyMteosStgCfvGn9Feo9KFOV2Tuqyy1rcfm5UrHpl95hpWNW5g0
FdRowiPiSIsM7oPH7eO2opAjFhL0hx7yW8YQnXaN85+qDAa27uRlL22YTvsLJoqb
gY37tCpLfbahFZzVVLs9l9MtmL3ayOKDP5tJrV8yv6geWdWcRlPYSLYfsd5g8jfC
vmDY8E9GQ3ECExXCimtD8KmidBbXL4dlpXohozGKm1TbfihzTMsqQ6gx0ddvQxEt
L02b5+nC3SDZIqJwmzyeOu6ZMw2hPKVufvFSRyhKHIlHzemwal84u3h+qouP0skX
m+GC2yC2/tjxTMKbExcaIJ2ZQq+6Z1bdzkwsKUncDRr2M1KuH4rMke98AqP1XACr
haEUrGkbxgml6QQWYUrftt16tJFt56e6F/qMwDbkRMYVgJAxhLE7rvq4PhHDwokk
lrNoVlsZ4KZDpx120/Kd0Mwax6mpwumvpOIi8WH2J8ZjiAXlhf+e+jRVsZiF1k8f
GHMNOsm34xDJkzJ+V4P1Lj4FYqwoUg0Oz4PBU9g3TYs4mudLPUf6wTO7AY8zJNbl
fr2avizT55YyIto0VEv4/tshbmXHlr+1FVF/xmw5VRq6bd7wXEJvQAPQf2BgG1gV
S29yueYNWDVLMkwLt7V3SYVmMhDy5BVRBmz4KMIgwNx87FsrqLGXKPIb/uHQMvng
shvmimk5JMbWDprAixCz328sYq3UhEgR0durszzuUperOq6tzaQp/FaToJUdlzTf
YeblUkzRFomN7TEOFLumP+ocq5kWfiaI3Z3KOoekmX9rmyBMdcCBLEDL/HC3b1L5
FbyKViuI5NV8WIPtytcVNbTLxUlTf/k7lgT8LoQzvg97LJq9lXmhOG5im9mFB1Nv
jd3qT1DM5xBcpe3NrlQvu9YrzZJhVV0VtSPF4lk+aPx99FXn+i84yfpLTbVq2mRF
UbjiKn1Q3vUzOVKQxLDSmKdhCHIS3r5n3sekRi132lAbPNoINeOy8EilFNCLghcI
lcZ4o0a3irnSFbPIDKmEokF4DWdAsYrKcbhPYvXydtUwpW40MQ6srOvMiYRA8NnS
RdkrPsnU1khpCS8gWz1dHRRlqYE31baYhGA+yKi7ftueDJh+i1y3fEnGLXc5xYb0
rLyxxerEdFLVItMRX7GUSZlPPkrqFaW90j8mEDwfRD5Ti/uSaa2vL10UULfhk5Nb
y+aEkJlNNwchQjyk49Oicj9bkjRx87FuvUXQSuisEeOzCITkcvlZZBtPoZ30DSU8
ODkoaAnerwFLgg6ykNZ+OgPW3LQtXxJRTh66x0tKfJlYN2nec7/0WRrC4YaymHVa
Lv7nFhiS4MJWddrxH75dsTiikrg91qfnFAVWkWzgOdY2sUZnwc33fOSWXMkBJMZi
dA4nT4dqKxvgdGqFJUcMDsyg/rxpPdFfW+adeLqKuvnzd16SkiHCqQUpMiSUT3il
wE7pWck4XFKr/xyzmjO1zkN3FTzgW1NURfdRLYnHQsLTlD2YnmC6EMxUZy5/+eQl
8qaajMb/hPCfuDiMzfv00F3S4nAuP7xgsC5mmZJZP+p48IkKjBysDM4GC9CnVYSN
hHolWGNI7F5nBkzhnjmTQ3ryaRq/0/PGPyme9RUPJez6rMl03z+1roI76TfHbzC/
02I+PRCvtIdhD3oCRZgcD+pVwweo5LFpqtqXS4n/HQDupIVI5dRuEeCqI/ipeRI8
bt/VMd/NB/hiTILoCvIS8cON088RXtiyuMiTnua14mlX6kGMKDp5buZ/wSzmnnSE
07pyUHYsak4hKNZhV10PDmQRt8+T1al9ABbidWSYsg50L+9I93p66HEoeeTuCnhd
y2AOlcZ5Qyi04wWkckD0Vibpmh+mzv1spZfhX8swmTdRBJxZemfUkin+XLwuU6f0
sIPvV07tn2Yvd1bvei8bGpX3H+7wCiz9A27Qp6Pafz9ji1A8Ki5vLLNcsMeOY+2g
vuh/Lj6/tdGZFLMJZ2fw+xFiRVHwduab7hjt68dlvdC8DnJrwOjNmyYYlremqNXF
3mL29Tdt6YVh36+I2HSSQHzXCRm4Hp2PPv8XHG88M7pCPD7qYQr3BueSFPWx5Rxn
q4rGcLWSNs8OaxvJyy5mTVoP3FPJW4dQPYfau0bNd+ggbQsoWyMJhQ9kspINJszE
YhRIaz2KFZe1eLI6ZlwbUsyIZ55AzPGI9C5F3Rxvw+ARP/4LwtuE2TLZdQRgIXFI
ofK3JHHipcFPB/UIa1CfnzSg4YvZ+IetYfhI5lI6acDfoWffbsEe+ctvoWAs3/5J
40HkPRe4LSsfObOHHd/s96g2f5xxYBxuUmjGtYOeOSqy2g9E6Jmv4U9kpdgDdRyQ
CRlcohAnO7FSnKkhToJ4wDZSZUJJdadCBD6ppHZcga3Vb7vatn3+GemdmW6r3wGP
eB1wBM+0HK430/ThYsskRwiJB0td9dmv1li0w3T6PEdyot+G4WfRAyUngch+BlQ0
2ht3qOVSB4Fdjh2ZZdUl/knpKoQybhMfxV2MR44dMammYbFvqCmkGrrmhtL4iKYT
YwM77EQf8D2htdHa1Pps1lknu7GDZWkBsL8k70NQ86LUwfYwzVaNf8F1QFu0wO18
mSWDkKKCWh3koAC9WIj7bqAjy56CDV5Ppf0OhjADfuC4tX52gi32e4+Qwn2oYCRd
zMLOlL60j8DjnzrPKJBxAJe3/YUSncIsaRD3m2kAyWrJJRlNQSX8I1wjS7f7V/xw
/JiTtW+nl7p5/Duy6CWrR2xPigwIkzuLOVg9xbYqzanTa8lusRB9GSFGQCUF0CKb
5vOiXd3Ew/nBGm6y+MqnRGttWHc8kEOgTNbERFuRMCTjaaQWEwKuO9asJwE967eW
mVWiXUA3rO4Ay27PNd22I5W+JcUed4CGCl1QEB9mlBdJaXwPA+VhflGhE09EcuXk
XGPJKm5E3gBcGNciOw3+mObNtv19UialbfRzrmOmyDbqPH04cuktfMqzeb2/9Jj0
Tu0M4kFM9ts7MQ1EUIFMVFJekBUgFHlaH7aKqmaS0cApYKxIjdH+KAmC59BA648W
DeTjnn/oYHMlhQDnMTX10Bj9kum8WJShOJBgWqxL8pzednuOMXuTj9VM/eLYoEAk
LbjAR6dPve3L38K9uleLitqgjpeb2EWxM1nqo4m/tlGk5KCJY9yVUH9vpADp00jR
FoOuX8aHY+rk9vTkshc4l89vhDDb7IHc9hRAWeEK6Ug8iiQzBsXwucCi7zqpMeOA
VIs52y20RJ7NTOY/vvccwdgY+vavlZ+nVhizahq9RSK+XtJD9CnV4yvyvzoaJLUP
LjTkpubkoYbNDw57ez4GnQ+7f4ix0WS9AB3YiUygona/NY7ltRA48/Y19xK07aTT
7ZMa5absWxcw4W7kegOu/4Y88fiMmlD+DCA5exLIjgiuLO9VI52RzEBTY39IZx36
6UGRT/W0Qs2/7XnSbjre+hcSvbdW9IP2nKw8iftFxw68jQJaS6J9Pnno2Ck4NU/r
Io06z6xc5knzdYQbtUNc++jOgUW+qbXtvko8H11mP6C7C46DHqtitXcTHNhRVDYS
wlVqUZfVXsDmcejt8np8omcYVxfFBPRKbGHGQ2OiOPSP72ge0UhmzYr3LBNFSJ29
Bt8BuTN0Pz35x7lW2beu1vyIdAOGhwzeRqQhQKY5mWsWP+mug6dUoJM28tx6eQy2
QXT3GkYH1NXF7ICqTtqWJ9JSKwpjmM/Rer7GdYsGOhx36LYm+6A9D7LnBSf5OTZS
/Ufck+mbvoBLS9B+aDlgwp4QcPo7QOpCGZvfciQ1Jjw3axCrCxb56haesZGgKiuu
Ztndq1I7uQhcywwQfSbjCtVtlZc1Xp8rHoel/+VA5K9KEAIMmozDTPKEANIH+7yv
OHShro+ql4DW/Fyk7rNQDYSmWDmPEHVheiBvO0Mg2wo/RZrvxXGxWSJX9R4mY7K9
o956xz8aO//tIMFQQtNaVPsquT+hbt8W2J5aRAmdDt/Zs177l3l9PkvQWF1qGj1R
E81h01Ui/2mZrf9+ilChSYsZhSxtRVwxNsHSi2xJu0YANRl3Cvt3pGx2lewOhLfk
zItg/qxzJ/qxHdshSVz6O7ZsfpJIm0Tm+DPHglXzPEPu++6Sd+LtAXyTC4dV/ibI
ZOVEkVLMwBI0pOunL3XPOhxfEssq01iUtFf1M8Py8hizXy/Y3Y+/SkeSts5T8y8u
DZZim05giu51zkAVFcUvsgwLYdsCaosW2jmpA3kpt1LQ8Br6udf1Obh5w/cn4xhr
Wk+jzb4Osr7QUvtAhSs3Y7troOCsUprOPoRnDHBPRAXMC5BKuCn51Qcqa/hMoUUx
JsDQHYK+hrTgYRqEwJ2FSRfRyKdv/Dw2XDpNHJy3c6qvWsgc7myc06xRYkvtRZU0
uOGWUkLgncESPpXGGW2dPtNFw1pkJdbgMQl/xhH2auTF+ueqsf+l9P4iG1v/nAfh
827IbZy8E0VhjrTFXWRfCVwIWSD6Ha3B9yi6IftLWH7LPfR7hDnGphU/glBahXYx
F8qtjipmCHimdhKQUoEiKmIwdU5lcpn90U4hJ+C0cPfuu7WfFi74aAnbHOLvxU9T
CWnA1VIbxIWv3aoGWsLN8tFvAsf5yhAT4mMVifHETpulEhAerH3zDgsckh/ok6FH
sUg9jhQWHiH2bjPnw6qRd1vPjurmUP3VDf6o2mVI52cbbM/ug96d8w4oxzHykyd6
iX8JQBlzNZL07/tDcaGBPT/HFGrbzSlqMsiOg/vwnWXeg7mVU7e58SUiUaLGBOCw
pddntLNPPx6f+KWkSfdk1BQXU1UZQcVfqdszPd0YQEAiaUH4EfjdXcsHYHump7pz
Fh97dSklXYUeJ/WC2W3uZ+6Wb2ccLQPtaOZdY3S1bRlxaVhgCLcJ2fj3oDMGFYI9
XJMSN41LN4z6LrHG0CCjr+40umQbb0SAkt8jI5sMYMGQSmLotCXTpwSazOzHyRL4
HuDSpg0Omgs53jTN0MJFCMGngX6D9bTsaUIS9b7vREx7mxLWUQJCI0FmHkLtzbxD
vJJJBkPGJCPS09WCzrkzH5cUjAzSCC6vJZW59N3S0iPIa1LbzYDvcECedOYuEz8J
YTLdsu2o3Y8KzxUv0AcENJLgc3aEyRR3tvjoR0wzxnH8ypK4MlQxfGyrOh9gyRE3
PuVX9vveio4bCLcuhifOfBrBByzVVUDQ7VJ6Oq9rO6bb5LCY+WeKiD7aKEdZeLRv
x0gZsIyKB+UIGjy96Rppe3/B8P47n/aU/NeaME0xYSIYWN3WqNCg7zhEKG1Qbz7o
fCcO41nGDDX+i11wtUxe0PABBQ5GY7l6854U+qEVyUvbP7iRezjUULnNEhw+nFw2
1m2yB3xDD7lMW/GN97wZq7wqvS9ITTZ0OyI0IundkKzWWMFR5Y/dSByNQ1+dbd0w
zjkO/d/4xknrmZDeA+DrfQ+eW6svI/Ee6BgRy4GOkOaa168ynRlcjEUuU9tHyqCk
m/zAQi8cgNgj4aBraxQ+xE4vtvA3tm13A7JPGYdbu/gDM8LPhctE046OYhq/o3Tk
7sgUfmSe5zTEKMro+r+o7zP6hzVlvar+Xq8iFkZ9YvdZo9jBl9wsOY5D6NhFHPBK
bV8JVqNohOTjMt0JaOYD5D0QcWajw36SWmVJXDmGOR3Azlzo/bu1t9pKLOzwaXH0
gNKNn/+niTU37it5tNUONqjE6+BqMTKKibe02C71v79eicR2n4bwoRDHsVlMzgYS
s7CctbWjX2bOR1ypHeQk7ppCYlQzY1XZLROhaEJTT4OWmp3IinSe/1Dwtx+soUEZ
pHVNUF474QxDgkpJlGMAAa5WFjB1WBpH/hXRfhgG71fBruJErrUSCxdPdnzeKVQH
9IaA1CoF8yKadovy4fRx8Kt8bTp4akc8mOhYHOShNaCeh3UcyW7HRuj/jjk0Wlte
r20i7pAD7ZaoJG0s7buCODTE8YfgHnvDIioOQvcdfOAD5RyCgEefH04+HmKAN1i7
qV0RRjuF4hcqDdPu+2Jxd48XGtTTMdDpC4gae+wpOOMQNwtWDymWBZJNHAr02DVn
ShPjd2I5NcUF9T3UyOD+S07L5lVy6pTvR+LBvzdfamlywAiFZbFkYK8N0BMfnVuS
lIbTPfScpljN4+1C1fZ27sPSyPVRIsTZJoPNT7bIbkvPeXqM+VUTGWgDZfJHTVtx
x3w6HAhDhwLue+m/22w1Mqdjj67+NIDwNe1/UH+7CFgm6nUE9GwuKNnEPeNt3GVD
5yWGYXgodpvv2mj+ovFX/1Be7wdIVsfMSsvb42Rye/A0FzOLELTE/5L/43KK6RyZ
+KJUr5FS3AoPPsyxijKM2qjCqXrw+fP7kvXTCeewxVSPPrY3SCcOIeHpXhp0wDQe
HZabu/pQS5az3J1wvBMlegp91gGqES47Dz0dB5qSdAQPuy66gxmeoTt1BnyuMTNJ
svDeAhu4dPIuZ/tJ24bKtiqSBzViqlf2BA2RxfnJL1P8r3jp1ixa/gRAncM5q0IG
9q4N63EFBG6Y15MEM1ZCHxWvzZX2O4dUPnslVNlM6Vvxl5O2dcfsCuGvxaIjD49y
bosvKx1qSl9ZSumn0ZyVxHjZd7XQyQI/EYwF3kbypQZWRdSKgvENgv9Yy5JlUmB+
ORVX+NgLVWSG/xjwlexydivDvk3wP7X5yRumk2I4sL1tPIaJSFDEri2sq88EgU4C
Am8T2Tr8HTTmIvTIWjWw1oiG4GAH9ANrY4AgS44Gty3IO9xPAVu3fNwdlRmmwLMc
icjTbRQe/6InuyRGvodFHkT2Plg1R7rQgMUlcO5HqNCGF1DhKvkT4Njdvc9EX/dA
pIyLProgZ1s5N7USyX5pzGJSdBLUOSyDMSJqj+efisRIq7+nO8WygMOB43d1iFZX
BzbaUsS8m1yNeHFnJqNCGjiA8ttdFbhXNglkznHWC9QJp6jEMLXLXEDf4h+lFH/1
Hj4YQxJIVZ1WE5Ro28KONJqrHY5Ue9ICh2dpGfkGAaJmIbfERkNjuouaYaANNBtX
VBesS94Vo7sYni1iqZPZHQq008PLZkp7S8QhXqBssmoElv8GDGZ3sLSWV4eTynW5
vEc37rZ+60i93wbIEkXxD/sDyIx1VosZKWyHp7BbaqVOPyugKFrBLdIPmbPjSU9X
qsOvU08AIvyMAYsUklSCO23Qi0liUtcZWl8KU4dIIo4WsynktVqRK4LKHOgU72IF
7tmZkQJGiVK3W9+OBrlicxpBKqG0wkR/Bt0kqge9U5oZZ5HoHn5IGIBYSBXgkBJ8
fK42TphoorLpnIDoPsU9Ste7LKjf/7oTX4+j8av+vOtGx8befyPviAUAdnqj6Kzv
U9FnT6/FRn0EmwEjMYOYm9dVIeEEYVT8vRVyuu1jJVVGbYvXYW2CCN9l8tbzjD5k
qUS83VwaaXPpx2ob4+NRqoMI8sMn3mWwroHhOt8/eD9fiB7Mz0cf/3MFmSoQe2+y
BDot0suVwuyeVW2XWzhmb+AWcWKneZagxBd1JYMZb1o8OIde8A79qswkeBvvhmrp
03s+n6GJacpG0mLahJTIEcLkJKI6w2MYfYxcaUPLL+iqDMEt1te1zcrjOXTzqB9h
8fXkUmeFBrAM2LUG5Paj/AIzJnVGL/siWS9+StQ9P2agb2JB3r0tUt+ZvW0ScMIy
gTHxipnHNFDcrpyyZidRFkbYu0YgJ5MCZBO0mfHENxaj/cl2sFhM0yMqje0tXmGU
WYj0o8OjhLKrGjFlvgKCILVhDY35x0AxEwA0+s1SYFwjztrdoUzT9hbyC82uVjSG
iEW1V3Oyhrg2Tqs2hzeOvixAUQf1CUkt1sSc9Yr9uMQh/QWJvure/vVol7dv0Mf9
ANRy+TPsXDVH+ymn14hmEhRVBg/JwUFcEaRbnNTkLLdTciSvoFsjvJeeGnGxj4xc
RlSC+DIwADYJuHGbaxbuTScdoyrmrW/90xV9tqMr2S5yEQPXPf26ftpZ/puq1MQr
VHNq4MdJNmoTmkahPTT0iHVoDhKwmBzX82vCs4t1NFwSJOY2M1XjWrei3oyl5x60
xZfilxfno+31wk33mfHMjkofe8fGWH56aeI3euZGgsGAhpG9sUomJqwU5aAU41kd
9mXlOe5Lw2g50R0pKnfeMdKtYQrC1KQGLqJ93maVwyIuG7UKsvtgcGjxpEw15IjA
cViUXpt6RxIQsF6isdtuoHtZuhUzsEQD3F7S6Edh6e5D+ksKh3lsKdBzZm7VwDAD
4/Yzr7Nj0cW9aiYK85vDlA1ralV5MRs4YEs0N+TEJKCJ1PsIsjVEDC0+urrMveG8
sjh/9Gh851p7C4SEY0uDuJ3PM4UvfLwOaBgAlDYilfvvuAaziGnkJebjEB4diM30
gnCCNOOOPO8KEKtjCUQSuaklQUCbQ6k6z06HPtsU9sUbZezYkKbojI1YpPkYivIf
qxTyK1EJHmcxJcNx0e8hpJY0lv1tfPzajmy9vUqRPCtmemNJQsvadBG+4saaros+
gJlw2QGmIPY38kZ5L+g9NOUNwyWLxn9j96ZUM8NVvLCxFYvrq34TqaTFXHyizWfL
zE4NqEYCm4xmq2ogJr/hw5vgw1aiYdQoGaD2y8zbYN0EUBE303Ggik6LYRCBDJ2O
TSrUdSX3uLg1jZh9/tsIi00SNhe0Ccpndnbc9mBehi3zYaHX5DkCUjOj7YY6j9cO
HsoF3loBcNH5YK5EbCvcbZezbD27NCY0NlSdVT4BsMqBREfUubMmPwRwDSt5dz93
bL5M0Go8IWeAOUyk2pZOswsvCEpP/cSxWrDysRY4EQje3Ck3Ie/G9yA9lQ9vGQkw
eCAmr7nscUAv6Zig5W7K6WCTxlufyIbW7oRmGPTYcyphVtv/wRi8QDYj4f+mfh9v
okb27HLsfy/d1m+M3dV/yTjeWtAKU4PXcpQFAzGRpds9L4Akzdb04IgqMEgzZwcn
7VOaWJ0yr3WM3HfWK5yXiSesc0Gyc4NC2gp2xL7ate87vPGeszBfu6RGqj17Ju2U
jbrEMSCDVYJttrinqsw4mgCOJ103+7sXA2UEpJEaFwS8DudZKqWUSiw1aPA62O25
95OsED/OpJXmzIVeEb2lCXm+6faVpWn6GgdRU3C98jCajyPxbfhk9mg1SRSaLAX7
49rc0Ckany11uva3ZxCOcD7mfQa06LlpnwUeNDTgVIioLe8yLXeYHkNA7WrA5hds
wAhP5nauSkTmvmXi8ljnEMNcWryJswBS1wAQXw48T/w43e1G+I2LumOAiKMMOOEt
HKPEOVwPwsGhZNj/oseaXlXsWL2QpxPku0WrOgRc+28fkiaH6NzktmtsF+mCrCl/
XSLl7eeiMz5ICCyGQ4TmF2tK356hRQeKxLr69TJJ3zlmi99VMvdXPn0UptyNEvur
OoZ+I+NoDcqdmBoyrZosTdyw7U+glwyCuoz9dbzxB4V7tWd8GcwFwFiGZVNStC29
OGO5JvRkTgpvtmGJoB6h9LIlJt+TE2S+lVt8f3SQOruFPV35ybzIA6yLsaXJDBxb
uHOjGvfTjVCtF9NpoT6Q4P8JwCWNFgJePuCtmgOTHJPs6YVGjLrGonm5/xioLlae
35s52y0jgbMWsQxkXXeXxdvNvj3HF1giT7t89bBNvWa9CM/9TDCFt/FLtb/JDFn8
poutCyPnPIGpllcysfI+Tjl9AS0L1ThnjUAHCJNIw7UZwvHcbSYZRTZnOSXFVz2q
1RR+qf3LUWHz08NhqTKT4ZizqofF52CTjHwIvZ0qYm/3r8CGI2YxGGZsuuYkF7a5
Db8T/IghxKQ/du1VsUTuUVv5znK3sIc6B+rM3FEZPr8Jal55Cr2XmkSN3Mg/wMPY
EALbKwlcd93ueojMuwiXkB5DCj4OWy1IPB3ZC9AwMsHBHH4UX+m+oHuR3stWzopn
XsFsfEMpj/cJSUjV1LAnmX7sFXFvtthTnokG4gfx19Un27UU1xs0PyPrOrU663Zq
FYBvRPgNMK7Nw5USF01pXY9q+26FGVQHHG9wXQ+LlFXy3ykNoXTN8Luclej3mNg6
iotjdVpNKvxcuqpRnsmFscMpXB6pLWMQzX6ZF48w+u4GaCfRc86IaIAgVi3xNEsU
Oa1Se1UhvIYu9CWI5rtN6nB9qvzWZXybGLyDcnCqL140I319gkAbZAKzx3Z5ht05
DP96Mql3WWEFBE5FCLEOTkNgDYf5wHvoRE3dNiBmc7W8pl/BXyRmZ9bJFPM1b+uy
spWe2qZ6I/a2DQkT/lWA0xWOO6twRTY90ZWF4X3eh2ch439evTIvYwjPBvfxwlFQ
+IeOj8Iv9VSNb5Zet2Tg30BmMmWwKANJb/lN5L5xLAd3mVkmx+A8OHBiZscvOmLS
eV7F00PEnf/qwySnrkGvwAcwgmDLfTbqXIvRhuhT4o1nm5E9idCfxvE13a81fx9Y
2lZswTQZkcrX7DZAoyg9ogsYv8yqSYcbqvlUmt6L6Xl8C2x0Elu7pSz9+5jZIo2v
YZ2asg3i6m9I1SS5JHeadOuv2aTchfkW/kiEMzK75+m1SlDL93QQExHiqKAoTxjE
1xNQS1N+RIyZXE92/q+Jmr05JhPqv+nk+Jie71XTNOvJdJMlVFk51fYYZiSPYo0f
jUIBAP5Hxa2Qghf76+z7ZjdjkQpFmTdEIi9pzMm6ZmHAO4k7XJEmTkyHEW7QKEGn
XKq4r93HPfkO4hJhuP6yILteztLf6whNSW495+JghxU1/0xWaPK3g7ctyCDmB3ef
ihIpNU+CgGSneK4LZvPa43r/8IzApmLhJKlhzYhIjzn54nX1rA+zo+vzg8Bwoplw
8QIBFpM7nBLDSpmayTYm3vLqDVkIc9erGYJoO1gTXRVAuYKho9Yw63ghV+WA8JnH
5B9oJWLHi6QiKKTiirnzk/wRf3e6m/F3yCY45OtcDdlboX1xV5/KJjS5F4eHeP3m
thx5XQrPwL6ZqfXDAr5pmUh5OHV5GJTeZ/jApfIyWZauaHBjUkJN2P6aqq2enFdW
wuQoZBTL5pcOotSNf3gA9NxFLvzOqDWqiWvlxGV/AyLuWNYFVWI7ugqT1OL7SjPb
59Skf8KBAX4yL7p5LfJ5H4S369mcmVShxdUQvBQpdFfTRj8uA3WPmLB+37lAJ4TV
ceMhT6eqMvefF88ddMQ41nr2IuHB8D6mDvSYR4giH/rO83+snEyOaqNxV1Kdjv/Z
wxeLe49ha9EHgfBTJPgGRUxu6qVGzKeTnmzt37kfTgyC43zDtwaQ5UUa6dJLgoUm
/dBp6Qfum9vXg8vzMWTNJwCHF6oFUUD1vMK7Lu1lpxK2WSMWftFrlkb1Ux3KMsNp
gr7KnJ1T77+Ir06yyd0JJwoeatuXX8xMFoftojnEHqI0dZLGKtJ5M+Hm7LXUBSwc
nuKezpBd6QGKNM+HBVs176A1d8BjoWE7ACBS5gsSFoN/wZyliKC2Nbc1m3ZTouTz
UjsbOkajeqfAw3JZC5RLtjUCxDN6VdP+lsrm+Ui8ypio5We1bQS6TS4GnCUBU22P
GJj6IkxgYoMSize/OshJyKBDpD/uRRCuAl7jUUsRIOuegQuJ93cc8EYHrg2ljrFp
3kfP9N4iBHXKzsJqkulGOOiZ5V/fVNSpC4rHLOECt9qvtsaJduoC8eOfgXjgtpyV
Divrt9aO8qGQXgE5QSZB89TXIVuZ0vrCRXcYGaQTVYBz/PT8cRjgET8LEOOtfKwP
C2fAPL4acVFZGJhLS+HWoB2bVXyleo32gOtqA/KkV125YOAHa/pdFl++sSIIVa7O
i+lTJzQdyA8Y0Me5tgjiQpxJrHdvbjOvE+nFda/oRcyW8GV31cb9Siq80uCOfR+F
M3OL+mWGcvC9JoyaYiiNyvxKe3GGiQGQ8ctGTRdh6sXfdwVbqfpYUi+aF1Xtp9Ey
p6XmmIOStUgMA9RlKaglKM1qmU1Ft+r2Yzm5RerTp+en7DOQ33X+7PBG4ZNEHipj
n6SsGwxAHKjbxNkC7n4L+3SR7lYlWy6dkZjamdNBIxrblWpVcv8Xntvk182B4TP7
ofGcZggvW1J33mu0u/4kYHeAD6cARVG/31WikXnDK+kQKB7QLFtvMqhdvG7+ysSm
mifZkx7QoSzd6iw7FxTgMHBR3c/UeVEvoNQYMGUuAX8KJJQmlLor1DkYLhg3vmxc
PWhYy/1ORRkS4hMXtjB7KeACxo5+YWq1L8MNVlvo1SgwJdqsjkm2WIn8D/BlzYat
dNVfWomMTP0KOnCRqbFMFzermz5Z9+B9X+b7pYzyLspJ0F4zeVvreh9ahWvPAV84
0EwOIpv+SUwIBJSkOW4c9/r0ukxQJZmvn3Glk0RQH/2YyI7Ch6L2qc+9k0atjh1T
/MLgULwfXUxH4RwFSNM6aNCUhC2J56rnnCUnXsqxx1E1KmtCrfxfATqP1MSPi77x
sjMaA5apYeDwW96WepSKZw==
`protect END_PROTECTED
