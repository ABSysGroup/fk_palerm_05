`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sdXTsKmWRfo1/5M7TgTX7RSDUuT3CEhaSsuxPl8F47BtApMax/sBsvZNsbqZCgaw
n8yQCgbR7G5Jgi9hje4KN2yJhByp8PYTHvvcssrn+70/HDK8Fhmj5s6ITKtci+8u
M7LfBWr2ItTwzao846hXOOIhKNNVGtAjANrQEHrFFFaB9DONJ2QCVCyWJJLen+SO
tYjRDtCQ729hkMHp0pJ0ChZFaw0JnB9EJDcpirAZkIjzgJ2ZPqv6yJf8JndAQSQg
IuO4uweu2TTapIgl4BhLSmv5HfCq6y9GvEljBgewJmghHWRF7yMwAGoyz+3AGq5D
vkSNtD7/ZQ+hOFI3NIV6dFrUtfl5w3y7G7VKa6Vh7MysaauF8AgbOAFxymzSrWcE
8//79LrbchR0P665RJTK51PlQZPecMG4iK7/U4n+eJ6IU4eaN1mxTEHYIPlSO2NQ
fOOCAGqwZtZml4A8/ZSqNhdRS+k8bQUtlGRNt3HOPfTpZWhgpabN+u2+8k8G4WFz
OjJ5C28Vypo4o4muVdrnYe/lK/OuoXisMIpA263f3Iu9tX0ZoPoJcNk5H9ORXDcG
`protect END_PROTECTED
