`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nr88zwpG6ai+stbACgKVZb7n67DC0xKJCLnDMHVD8ZioVUSdnrZXfOA5kVhDcChd
gERvKwXU+q4KEGidq7zR3qTygvLUIFlDPabctNiR2JBwkvnaS84NJ+2V+S28MxnO
97qhj0RLF/WgMFix0j9Dkqz97OKb2Y0qo0FdGm2luzRksKfNM8WlBjG38iqAfave
BmztwMGEPfWjAmrD2C2vvVFr6iuFRb4EO3ooQHEhXjPzvF/a+tQa3I/RABrN/Kf6
oBTSGsO2EgIg547KZ1Jji0tC6tlT1tOUYFxFBtfNIPhZcI7YpqhMuvz9+EEtaJAd
/O98X5DhR8BXbZxQ1qZkPzdfqrlfNCgSBgrTfoF1pdqlelssXGDnJv8HVgZIAiEW
9kqR7JvJ7YWJMYE+SuxDaQ==
`protect END_PROTECTED
