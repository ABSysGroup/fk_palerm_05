`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gDyKgJPzvRGTZzMPrevjQQjWa7cKmeCV37dCeeMNmgi1OcKsISZzaxG1YGq5Z9ER
4cwpGTIqXx4KDVi7VbGG4uweBGxtgKyvKLnnObEHESJ3n70phi1Dn/2pKK3tbHIH
IYMRIdFVjIM8UZMiVSMeOgxkbzz3NFefsK8qSMhzVxzSZJYqGmoj/jvTKnMZofn7
YtCVICZ7pc/uUo6TfUQgsxL79O6j5cYlXJMObHt9zj8B25tNg0sKLPpX4PihLw0y
r+PP9yACmOQ/uG7cJ6uvwmA1jiwZzqD22k61WHHcAfmPuyVe01VWryYHV1gC6ZBu
Awm4bZ7FkTng+X30V1IUd/HA3XS64DymNtT3mqrDk8yOUWYYRKSTX8URqVRz3fjV
ouBtwPM6OhvI9+hyzLwysILzcbREF92bVg3bHQO6vGoWaVhoDg35BmjSpgRfansm
E73lapivXyPOmckVyTdoVJk44VXJ5quGvFdy2tJ0CJOlVUMMU8XQZkERIae+a9TO
tl80npjrYaFVYKqnvqRGCIoHvJEsoqvp5Y0U7Ey73uc=
`protect END_PROTECTED
