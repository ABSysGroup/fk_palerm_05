`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XRLTA9GvTqAXLleZnYnBWCfprw1JceS28RR53VH5a1iJHHXn2GPFZkD6xG9e8Z1C
64rapm3MB+2JjCdK5yTmNVJwHcmgfKupesfZT2pDHELQlIi2I8LOvedOAQDCkUKy
9RpSttAUcg2x6CaBKp1rE8F3WRwffgi4ggXrSm6uuEz2EnDQ5pRVcCrPUibbAJgw
zz/LW9eH8+E3mATmM/4jAxaQWCBYRX8gKqEFECHVx7z4b57EUcGrhDGSeBWhTDXK
nkbRU2DY4NFNBy6FuGSFwmueYbl/qrOD+smq5UM2K271Hz1H0usfeoAMMx3mesdM
yZK9RBjTcDTTZWpqqY5ja8ZFeddKZMpDq3VEaGx8Lg8ePXwPZzEwyAC5UQzwGsdy
Fv8csPG3aJlfHIOIYmf9PgWwnBmoGjkeFqUe5YuD/hgmb+IPrM3+DEakBiMJ7RaL
0P49LDxTOptv75DR8tBsn2CHjmDD+2RWjurEl6cFDe2Kl1trmb1D424btDIWW5TN
0zKYztYD61wVqtGGYmyisWd0dA/q97RajwtgzNbTzxfKjXgupjLgalvR1rPEau+h
fY0//w7lTM5mNCePoalC/EqH0Ixj7lMt0p4ytRqOBn+4Hz1M4FCXCIVLvwBD7TQF
u5/WPyLauHjM/ejELV3g2TKwXul0Hnujzqlj0KbRmSks1rt/sK7+x5Xdpspv2AAl
0cNT7CF6h+jB6yvSKLES8CDpzOpScbQIEEL8yxAVTCiPaZKN1QI8JtoRl7dD8XlI
+Qamdx/AA34/pp8nhByLig==
`protect END_PROTECTED
