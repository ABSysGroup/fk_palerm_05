`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Z2K4B3LG2ABRGEd9NL1CnFdkJLvvJkOV+vQv7RbZhgHSxBNgQDvnL7Y2SCVvqV7
5MinPvxwy7F5TdAsM/Ek2zHj0R2OVGdb45xpXkne7G5MmSJDSfnOD0WCKtNyneve
7U0++8huwP9zFQeY+y/hOc7jj9r/ACQfY1pu44unuz/d6dP/ZY6xf4CSikz9U8Hy
1HcFciO9lN19Ez3Y1wApLYY6yD4blcPvGGaEZ1EvYSLR7J0AmKNffPezd+wo0JcB
F9vzK5ysqEmnX/FE25Bl+dF6sT4cSMuq8O8PonEWtuWpCU5/2k3RD5TYqoLhE0U4
sR9WA+aY6lt/1RR8YLET//j88JB8+Ixm5T6gH0f8yyS2B9h8s0v+HtNVmYprRrUW
8Ysg43sHKL0BxgxpVa8oaSAnbOaB/E7mgyiGJwYzDEEtC0ph9AD3XNukLdAxRjxL
JiuyhTV+dlojRcOzNI6KNaxRZNXMhWhvgINDrGGk3GrHIyr8nXDbjF0Y+5CbDUVG
dGLerpxIS5QYHClFWv/7BxmOUSUKtr/8CCaB6XcbKh5Xt8y3cMCX5gEvAKGt2JqF
n7em3QhInK/lAueWKFo9qoOn2er4kCcjFblox5ftX+omwXhiVOiG7VuzRgs9W93d
n8NVI8vtLBgldwIGrKI2LCduuJIzcjcvdLeSWS8n9b1EKFZ3HqSj+Zm+GDbiKYVU
tpjmYEMXLa6P/smaQTMCqhdF9QY3VPh1TUfoOi01U3/MjtPgmbJbimGLVeqJU9ZT
e1eCpakgU7f4uJskmSB7coSBfKh4DqoAlTcObI3TI+XPtD55fiJx8dg7JCpilSnR
gdUHjm2QmjVRgclaS/2clFQ9FSYkOgy8bbrkuQ4nFxWovHxA8ErUDOQfxWW6+d1Z
NVS04MWq+ZJdW5UXxfLUPnj3HQtFUj5+N8H46Cnf34v5Gw5y+mF53+bBJjo2EAaz
2ADoCH/KghdxNZpmQvz9EXbkBe4jxI923UMdv8KYONk=
`protect END_PROTECTED
