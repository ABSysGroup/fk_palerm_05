`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6OUlPFCnrkuA6FxZPWabo5nHH9KVPxeBK0mWv6rvOfvQAkCdHeknZo3WCSJKij59
NdIFMiZWb5Z3rqvgzmaJRw2c49QxYT96wdfIr1Fk3qm1BMf/6nH2XR6oETQqHs1E
Azj7d4dWutXduuGZ2L1I0MT2tQgYvDjaeVL237upLNL5IdGs4uP2RH9Ia6TDrHRB
JYsFrATQ0L0lyBZCpGp29XGRvB5Kr6bz+FauZE+VNGNfcYdflWI49gJnrM+RrEC9
3g7wlp4kesT1fioGpR2MJsTR1VH4hiHnrpcs60HcRsN0CVbe99gUBzyPBCVXmovD
jEEn43pHU+IIhQnJRTcXio5DDVIYyS2IT8jnKdEuZU5vod83YIEZmJ8il4X6tcsP
5/BDQA/EfotARDbI+PQqB9/aRZo8eYz4aeXpl+UEj9Z/lSM33wCwwyhTrIZNj+8j
D+yhd6MNFPdf4Ah1c7fGNowl6DEpXQX+UTQjci4pdVE+fxwUuo+oFri1vQ1nu1KN
QG3kewXJvSx0+cMdmO5CZ51Uf964z541Dp16qQP2T3jJoXiL8GVAk0A6xtWg5fft
5mbhIeqdqktP6D2JBwKGJNHUxteLuOk/euCejr4fRUZho8sEcgjVN2uf70tQtcpO
KMyGKLwqmLwErmjAhPzV+ExoUpu8OmRFKGV6n4axAnsII8RQN26gB0SEzcfTL+xy
RRBlJVFd/lQ0nW2MIxMiLcF82He5PEu+ApDzKxFiwkzvV6s5kNuYBhM59xu/KSpd
sWr2Q66vxi69ZsON5cJ6IhBv74cjKsZdAr2Ooj5iKHKQt7p0mm+qECR/2QXAphMd
WgHgJlIzyHG+tsvEr2JTLl+KZwvY1P0n1/6DMTkGMZ0Uq7Wgjah15tUFghEntC5K
TDsMRS2MatEGcJmwK1+fNLbeoyPuKEnCVPN8Pjae1YD8LG2Dm363QUCbOFNYep32
qDqRhtx7FAEI9wYYWxKmxf52Faoz+U01tS0jkZURVRvrHRed4xRR6LWWqL2br4iE
04DdjGeOElPgcNZLHeAbEzlTWhDIdtqCi4NKzvTo+UazvDjHCVnFAySG9oEU/KoO
XQ8G62eLc12RR3qFz8WcQoLWHwEPXS9VKRwVrGqBxQT5+rPx6bM22ehMm9x87aZt
0R+GRBU35XN6hy6Y7vlOrgTEOPx3CZAFL9JAuqxC7HIB4NVnKRf5ahi+d3TCVjCy
AWOSGwZyaenulMO+fw/SYtkPkmS24GKCCVlJlVSLn6KvU4NVZibJjNmr8e5Spm4P
qfmZlj8/MKRo4yl9k0Zt0PvxERBe5Pp4DON7FeA1Y59XxXTo68s3eK43ZLa8Itar
EaEumfSAr5CyRnP0XSc2hvzzkMspAfPikjHU+L9MFJpgXdlLsWttf9Uu9beqccQv
UX6ei0KoVaxYXuP+hxyvPVGCfIlrQsDLGzIuSQOi7C4IXvVwkeKwlaNObQjsctnv
gB1YzpJuzB/1jMUyvt3dIkjZ3+atVu/IBSXHmiF0/UIUalznluTu3rr6AKqZDKee
Jqi/ccdcaRvyQ+61YdykeW3q3BAuiiO/Q4/zxhPtjPxG4Mn3bOh5YAsVaQQ3thz+
E0A2lxnkCaGXZ+krzvp1rAcd3500H9VcS3ikY6jv1nbawvWhBJHCBsZ/XedflXVw
uzLkXJt11urofUBM3WFHPm3glFsn7OnL7QeHY1+qMjMdUrGhMsbtuijio3wyfOoU
Fxs5k45+mys81yu5SWbVlE/BVq5jg2oqyKD5z5YNdZjQdY0o98ouF65gRNXhanst
Vc6Wx/6+MAVhAV63o8lVbBjEyaz4UYxUX8NeiFMKAh0SywZJ7kFjN7hBZ1TrIEnR
9m6kS4C32y5cK/G5pzicvoFqUCc1iq8lVKv15JBmM+h8fLDfAEldGehDDEkHttoe
8O7b58WsMLnC234/shG3shdXRT8YwbBf+c0tDPlZd/pPfVxXCwDK3UbF3jqJS7PH
x3Us5mGGE75PpJnL3bnSpiNs1klNj4o7EW+/7Hrfxuv4SU2UmV43Vt6qoUIbK96V
fKZuI8s0CDv3TupqdAmIoWe2EJC89TjUxPpR/GrDT7b8Pib7acjUNf+yUTYDDyO2
53esea8UtXOOTAFq23WOYWls6RzzeRAP7VKD+K5sopHGFVWxpQReHJDbP23Akm4J
OYqTBbWtuonNJzCje3CpFi89qwwTpvBn90aNYf26S2QvSLRGAbkxX8nxkPI86+nG
27e/EYJ1T15jhmciCi6hGXshKC8oPGkFXtbLU6JI6m93uxA392gGLlOHoFz7Phlg
dP792utNrrztXc6hsgu2GvfGEM/XVakpqRP4pGy1QDvs2EHeyjAQnewvMEsrvz80
S6HrSOyQGzEDuHiBS9KGrsgXeqUBHY8pGWJ13KE/ZnHDPRXiF4j+aTUxJZrTht92
6kJtIuII+pXkIuLLexixSbz1WyVxV/PV9cMcD9RRCQQPRA2onqWNTFWRCxyyQEeO
DCGXOJpa9CiIBNhu8avwqdRSzUPQ6YQG/I7NkkiG06cnwFeYGk/WqkaKsiVKgn66
IP2gru+3orfdcji9/DkVtiez16Y+HvckETK1LX6rfukCvN1fI0yzR/zcvo6H0S9q
iSAqBMYZoNXurG5/3U8mxLRcVCA5+ReuNNKsds0JTLxJ28LLIwgFoVh61KNqVZ2j
E5AQgQKqZN4gG49rrZk6hcIECKWIlEXaSIFRErHP6Rfhi0Sj/GDYlgAiW/jcNDAT
WgBXDGYyMTQc4bqs3ugz0Oqnj8WjopLHEl0AVpvkHXGuMXC+pqAoTIQMqxsvroyc
VFkjZIkt8TF13tWzAYlj+/svAKU3mHT1F+Unjuw3KqeqzM5RaTFdK8l+BZAgG8Ye
z/PD/PMdgavt3TA/zRaC2HLceihxqT+vX95lKPFT66HgjivdIuqizHtJEf68yelh
Hn21X5NjPqlkZ3D+C9NrHmbKlv8VQHB3etxNt/ICo4pxX27NwPNMx/SNC2lxrxLg
uGRGAWnFvckZrM84LBatSeb2oPa96J6KrsrHiHqrjoFJfKg6Bij+aUmCsGCIeS7z
P55vo57vtnkuHDjkU8L01FAq4ZK0gECPySGE6ZNjgNKyBa9ntanUEIIedv/+wuiV
FBwimMw4z2u3XkKyNxQ6FQ==
`protect END_PROTECTED
