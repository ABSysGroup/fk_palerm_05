`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zzHYI0JCuyyyGiFkopt2Hyyp4udhLhK4qfXTWsw4IvobW7Vbi1XtwkuT4AaDHy2L
oJChGbGxErlhI4oilOKceUCLd3Z5Za3bUjtxzuP/gwjMdUtJdKjqHlSo7R3SIlj/
YeNWloG7VQtakezqfBFiXC/7C9GXXeYxwt1W/D3ItyatuBjiy4f8gIG0gCweH5QW
VmOKxB0fuZk7RGQe8+pnLCYr4xaE97Of0uf5wOct/mYNzCgtrDuLSFeeWXsrvoNI
ShsinzxZUX/y4HtUzmVu2kr+1hJl0Wz7MW9Zb75LLlCKB4TvVOrIBhdfs3BkfZqD
5ttmyS5NL06Lcr6sb79+wYxzenAp9fC8av1iAdXB+tZqnASoWK2zPGkGHSuNwpQz
TBV6y2Mnk6vM/7I2Dva98aDLKwtTczG2ILFfjL6oKCwmGrO6zrxoRQkioXC5V0SN
YbBeYNJ7KBwNboUUOLVXt3RlaC+gYcSzWV/2oyc38+rkjmN/RHLeW0XbShxvq+is
20GUelpbYNIKbpjzlMr2yuiJBGkkyvrkSUMk/DQ3W77l4Ju3tKgVKhNOIFSTKZE+
lky1+ywYNlodByUPacYymYN+rDrd87TfVy3rRImyEbt+3yuvOH9fq65fsNVxHke4
BdNlIXvVnHU97JPsGoepUOxXkU+aBno3LyzLhyvIvD8spqKqSKTbnBwxJWRNqiYi
V7JduXbJOKsc7Nfjhb4xDs59hP88QA/3AWfcvxfDvffVywE5sgXIDcPEw2y3WmlN
dbqeZ7qzYkZ822bAlg/uaPiLW1rt1NJ8r6u6Y7Puye8NGwoAF7+fCO/VRZKPFksC
uiJMzLV8DLCaO//eaOqHkNsQLj6o57MefGmhyAX/QJGO8EPGoM3KLyvrDWhNdQwr
nbCEeOKM1408ER8n6obIzq64AtxesyDPYC8QSI2sUxdDNI10peL5qvIdF8t9Hyi9
CTCXUaCYnrjY0O+U0Kw7lE3GUkC3FocmgbuFOb2TiHIyJQ2GaWBUK737G/30X373
DXC15aBc/DAsVW8m6AnH6XpsGDBC5QHinzzb6cGZZOVVBuVRbGx5FJCAKxe8QIAW
b1V2oenYAD8RtlIK0/vRTm1Hj6g5jJUJZoD+FBuqyQ5FSruHx7GIVjYE7XzXyZXg
05Klp/7/6dP9qPuOk/6WVT0alZQeq9v66QWpvEMqhwRkRaZJYM4SVFOxo/iJY2g/
LYlbAJREm3b4KPpJ7kRUJtHosLGgj6Os9peba6JieOQWEIuW2w3cGnE16apk5Sq/
K8uLIye50HUqX5PZSn1p/yRwRwY+KDrxUxY9wRJUpRfy5qlSvgnbe9CLksXBjXyf
x8W9HGxHG6IbDBekougMxOTtuBnqdvvFiHifXbl5ihV3xFg0I54dHkNUMVQqQHBN
z5SEGtc51u3sofLF4tW5qtOwtPDDmg0vo+negI7mUfmnWrrruE/9+pBOTAaUwUIl
dxa7KLp6hyV7G1GQrx5dLfVnUYwtBvCZXd2onkOyFjDcOS5fwGLyaBXcgjpMV0Cw
7sFra/f4RaACC3QOlvFZjPZmySKzdSK55c+AnKBEcEhcyF4kMWk8Czag/kUwOjEe
xKKoXe3346ae0dZVEcQk4bJRoFlfPMwIUXL1BZQnC4lUymYLOiwUeuYdceGxEA8K
iF9Z5IjGiYzbvVYTlLEFZ9k7eOFxBp0hx84M+kSYXv6jjxaSS2j2nclw2Ikv1sbX
yIpcc0S3B9w8xjK9qz/aqMNyRPI3UY31gmUa4OqCOP85/hY7gzkaGUMADbOn2FAX
q94dwawypomMLW5gNQuJTHLsdieUXOhuHgfH21V5AvREof9vVUHBFWvKpKtt2/Dn
xWkuCmfqGUiGw6yrsf7qWb8K3AS+VFRy8VBA0mNqnC55kcmT5306fZN9GKx35YWx
sruhFNSFCbo6vJZO06J0suGl3Ek4KY2i/7fWYTlyp6iSp55IWMEdHobnJYL9rd8y
ydPr1SPp/cMzYpEGyVLhfEVm5/5NdWhk0LTakRitTEXJlTI9LPK/BO8RduHnbFnu
pK6H1y1PWDWvo+tPqNoPoA==
`protect END_PROTECTED
