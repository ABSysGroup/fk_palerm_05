`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xmtCcXDWcP9TWT8/r1cPTCMYAqay52adfGgn8OnGBCDEKzW3+JYH1tcOHhtG8bLa
ylMxufh3t+2tgMLof4CQXsKvC3E44ZhZ9wveAKUZXdVN3EvXQ+4uZCsP7KNkP8Dn
2PFSR608bWuCuxqfUGiENOX/nqhvXHBXZREXPH2ThV5pLoXVFs5NFgSOX2JOUfR3
3jsXfkxzecPYeVCT8TW9UzbicXLv+KiZBD4A7dek93+ZMl8+37Ed9sThCWNQfafw
BHw+OJNqvGnIv/h/knwLCWiOPHaPec7BX8CaaGzOIBFiTSPGvAlC9ptyBHhv8MoM
olgZaXs33zrKrMSGmVPcG65OgOfVDIru3xptnCpAkCQ13Mjoh9YKxansWUWoAqLn
mo2wFQaCAeqrNagjyAERzg+v53PtvX9bEhrQo8KKSRJi0lOJIcDuVFZkxnbYPrOL
R8t3dFzRRv0lLrN+j4/o9ixVXTL5cG7oaDRv1i5jgJZVsYfuLt+9AYzumWGCKhFw
8EvHYAuM9X9rEMn3AzC+sh8P562UPd7Sirwh5FQXRYFfTXoSggktxCj7TfVqy6lD
tSmYnAgqcPqIGfm26qYdFZYtjztOZCPnAWoEBFmLE7PmR+8aj9THu1cKmQirYHHC
AfRbu8nhf3NjjGjdh+zRqwW9+juf97O4Sxk3jGIN8x9ehcgzIMi4UxA2dYDYrg5z
zW6LH/D30YyFjjz69I31FVFzVKLjVHM04fpJPWg94r+C5XCoC3f/IjFs4GeZHpCX
JO5LrI2kOcvELdNmphYau5ISFf6gsuV04NHjFiwX6Kk+F2HNc0ujciiSizJrnxKe
Fxzt9PIlZu0TKcbl7+Y3638vNWM+obVQenorRimDEphn7avXOGJ4TAOv4mwcrj0m
PQJf8rv/QLjt2Ltk1+2+woKVRV9FHAKLW+ZC8U5vHjIiVcacngaDhOOf8u+rfY5R
gkRst/xSZL8GzZGfHYN4xH5YtWwqG+LKTidcQxJ4Hdbv+hRG7bm84To6ErMn4L7/
PjBNTpXp/A4pJceRNcdhSDOHM0+TZDEgnygwsCO34aX9FF5bGOIiKIuxMXY248ma
lVwEwhN70N8wz3QC2W+F8CU4cHUbN9AoLsI80DxEdqzQ1DZstIyUmDl0K/pUtHZ+
3q6DNA5Sy2vfGq0H4yJBbc/0pMAxvVRsv7dM8tQNaBbz5ErddVt8evcVe65vutMc
N+RdZKJfCdTQA+C911Z0NX4ViXn/jUe4wje3rODCab9jDEU/rS3djD1u2leX6wCg
iaSwNmcqEPm5JGxqyIuucpLuyOgSRCjBQNlWFa+OHTPI2lv9Tuo9nxL5YGqOwG/9
eYyjtdN5VEt/I8ApEilDgxIrbMUJDre3kUnkLC6Mn7PN1gGsbqYWyFzW1enXXPPN
Ygj2rgc3ysNCDCCYggfr333ZOtf4R8dVfdODQuFGEJjR8A2SqljF2srdNBnGm37h
XHo2vcxe3GMR/fc/+beyx3BBmv7YgN+LRo8a2bjcmQpjfYPItp080b0UJSI6lik7
Wb1/KXX7BP6PNJ2vqVk+FyupuPXPH90mr8oALNtnxEfPeHuaISxozf0C2M56/i5T
f1lfXiR/fST71ybbZ5pgXGo3MEV1UVgQFlLFniYICRlC5GuHtxqJaS68bMs3Qnlu
JJhT92SYyTlLXYOvReKJN7yYGxf5gRC4sFvtZJqBLmAfhHaEVCIt5PsJRvKk0+NW
+Cc1ZK71/EEDG8YeLUHVLwrDLVvd3LC6Dq7sMJ3wkc+xF7a8vA95nmqKmVmZ7Kk9
pqhBQbjUFHuuhtCc4TYJrz+kq09I3ZwCZ5+1B6zYRzQVeO9zfa/7ZHh3qan9BgTK
jaZQugTOQ+d1OjUOXKem1IvHwM3Kc6bLJVIwCH0WY4GsDBg5rj+GTtfWq1e/S16n
Hdka9Al2A3/vTle3okhXjv+iAaLxdkIKDKdWJ6T6O7tn230zJwBVrPN+Gbkl2meV
8ycaEfZCwKH1/iVNCgyG2xTptgR6RTgf4ozv/WJvChXL5fDpqjBssRw3Byqk/a4x
8NiIRF+B5ThJnQvOC5xQjMTGgu8X7aUBICQwTj+2bxlp/l+KSH5G1B97ZV+4FasQ
sJ84CGLblKMsBLcPrdiieuWby7HixXavhbC8qycUA1yLHvUOdp+p2nRgO1PCQWTQ
I+D7Uz3B6tlkSzFUH0O98+Y1XWA1Eg84secx7tnG+JBlUub/ti98r4I280dtNHpD
FIljOkLVE/HO62yTJd+CTjSlSYJ7pjAp9W10SsVCBlzU3EZqgJOLPT6OLs+4MxmV
ZeZFu0aXu4qWLTTG3XaVOTA2mG9ySZmCtoQPQHdJwEjTGjX4Y2IG/ifszKbbQhaV
Huphd7nGA5z3yTiZ7yzLNOmFxnkZB2VJTuEbY1xtK3lO89uIbSJhNE0YCXPkK57S
gbV9ab2YCTlFBBlt9s4sz8MXr+ED3gaVeCOU18Ul/GGl1k2H5ssqxtJwAM3w+nzU
azChZ89PmUySF66koz0IEt0pb7mS+z0wDw8uP80IJpRc8gEyvfQfBuEENt/B93y7
EGYSjCSWrGrstrZ9tt+ELfJQpqcSixyO2PEfxmykTabEF5XAa6hbe6F9IeWCQk0p
ahioyZYvJIv/N7I8CmIXf+uupgGTQ9PuHtfkTNPuQ9667Z3QgaufAifRsOaE31bG
weMIok5D8OGZjL7gQNoT0kdO35F5NCZWPnOT6fuh3GAHrPsVP36f0vVQQSbjzmyt
+zzRMA63Ek/tkq0uCceaCjZCjRkYU31HRWOUE9KEsE0YbUJMKseLpgcrdAKlgBB6
w24QDdZRJ74NXZwyJqQRmjDbcAipDnMjgIVIN4vJsuZelPD3in4KKMWkIH8So2C3
GSOWB/e4/P3GDLdFGwkmFiXVfkE6vRujvF8FATs/xg9YCtzK8lo0alm3l6b7oRDk
lNoqbmrrftIYWNOT5437/yu/ZqM5Ln1q8guMVJkjHonyCdMcqj5vDlTFDlpZvKFU
D5MQDrcwKZiZOBKE30BpSb/fAkJK5gGLiHHSkzkR2LF6ToAU4C/dBOjoVl3ShGU+
lCOTVr89HVoquxA3+/URoO4OvuRK70noiChGHRoQ5Hf2uu5057o7oBo6vF/Y36Rr
Bfw7aSZGRI5gMYHkjxQ4NVdLmyl7a6wZFLQlmlIPgx0jjqbsDQsWWFn3uplL7cFS
2tRD4IhJoHylB4PgaHUc1JDbS6PgWK2NnIu1aRatU2NoxP5Yaafg8wv4LbBN33Bc
H+npjk00xB6yDqcZgF42TY6VHvlnxO4JFJnCf165lQvpUzcpyrbBbuE6Q8XYFTnt
jI7LlnbRA87OA//Ym/t48+9wlRMlT7JeK1zMsZSbEG/TdAPpUjug5X7ovOzKomAI
HQGkn1BP6nIX7uhOU/uIJz2Qr0As+eCNVfxwCyBovWD8RrF46PfihYil6ryqLsqv
FRqOOOHrLAF41cudv8IV6BuL8T9sURQvhJ/JDjS9Oa+rVeExqgqTK4wxJeA7BLIw
UUzhnZA2L2367dye6U216/jYtIABGK26WLKFIcKZLKcNFl2K+G7ozqNR03/eosCI
JuEzJ9dtIbvhabh8cIYznf5v60SDnChTZo8v3CTK6toFXw7FcIY7rX41ssuPDoHp
dGclfkmzTFiciKsWJqqwq3OFg/mC05RlevJV5jZlwz26zIK4VRbLiXzMIHkHYl4R
v60fpLxszcfxWJsvJ8jfFKedOujRxbqryW1CGshwUxrzAWClCib+vXMr4VI95Ig0
yXKknPxhdrtBGKbBTnIOUtTXwyK0CTME2X7ajIlqtE/JSasWG2DuZ+GHGwQUOdT2
ouJVN9guBi6yyyeEBAMXYXz2KJi3GeYA+Z9vKKI5p07555FYtIFNmItKUGrpnCJI
rrvnZaWCib3oEhemafkOJZduyF7gZNBxiZy2b77dIXuZL/5Dz4VAP7t4qmR3Gk7B
NuhrzHG250O1+NTrR+L9CSJ27u3r26bTO8FElOhIPD9zr0RG1csmwNOm6i0H1iYF
/5Ud2qmS11bbuPR44JEsv2Wp4PBdIBxrcYAnjmqWCAuonoKH9H0ey6zES5N7GWKF
+0ZF1hKjgE+zNHjGNoSBjYAKU8lMvvS5sgR1InAjGTyofIB92W0bCa+mNBN4X8wi
AXY7jgoB0lBAd+foPXY9wnuB/WQrFCgb3gGRxsqHhRRCPwJ1UIV1qjDg+BhQ1rb6
faEZ3NnlTqiUDw4rATFb/6LxDz7DXBfOKFC23l/GxIfmyQFF1msS2AXRTBfFQf9a
pPU6t2mpm3dBukwHv1nRnpMUQN0dKQ4O1CRnYvtikcioue8S3UNt4uQOnV1B5tod
UybSoxdwHQPkjjdayeD/vU0viHsJ8iAyE1wF3HlaJ6mUgjskPIdc415G+0mHkmZA
vsLsUr31nBwy3ckKNF6WRGnBAmWAL99bZ+8gh1K/2ftFFTt9nRyJFol+niiESv7M
Nby7tyHPEd0a87ZokF917lImAFBsVPA2fZDgukGhxRfxeazlK5d4UpRUIgZFk4kK
7Kt7BTSAjt0SFfPSs4S+kWkDBNZAjvbjvCxrznprPbbg1dlyiTnb4EVL42v4BYx2
+kueaNeufMtKyNCKp9EeCuqhHQ3VDUoNSBb2SolNlIDhYMOfAtPWUna5pEg2ylnw
hrjv4yo0QwfRGMNjmZC1zOOXL+ctM6fVfkpAuzUwymZ8ezkGYr2HI+s9a1DGQwyV
d3TWReEZC3A9/4lSszereB22q4/gXfDCP6f/0XgPoEEPxlqLV6ccr73MxLM7ybm2
/hBDGjfoU9xstw2VteU7P7NofxB0gqR/ThUXt0fr7uXEl5sLbtgYatGPau7Aqwha
3V7oqZoS+nR82DoJ7BS+0mbPJ6Q2mxGVLZ0KhR1vXYA8Dcdfgpd4pQE16jXcPmGL
y6/4XpL1T0JsG3V/pk5Zl+iKluA7ZVJJ0c8dRveZf4ZpeE1rK3zh30syZCWMVLk7
jObUwhPgxPW417xL8UR9q3D8/Y+J/ZqMjh3ijpa1hU/QpXtEZ8HS7QykQKUKn67V
aBTOTQcwoceUy8HQqp9OiJ7JWuhbB87gEosqP9cMsNQQX+HZdjI2U9knOgoGVdwv
IXveeh1S+VpzyjYRSxq42sv926r2cbkyc2QABOIS06QpsUxzUxrRQxEm4OiPqx6m
taziZrwcs73gjEJstRVrXKiK3iUV3v6OmkPoV+JIH4dpi5leXfl7ExcsbL5i2Ovb
pyXePjGHlq++TVNsKoGWKdbVEg1vGdYU6cuRDF9PKcxMJDbcU45w4hpO1+4V4feu
9SFzGvVL68Tg2mD08dfR5o5iQ/tQxoGQ8i2MlgdwehcC3b6gp/rW3ax6WrnVwPDF
p6ud11tzLbOer0NTzK5n6VgDRKqsnLsk+0LEyJUPzwIOVUnjoqImMXCqO6/79Eqd
sNWUihxw8FetgRMieDUGuQ8dXYhJtAFHu84Nxt9gUPR9P3BWimXmevlc53olcII5
H11zjy7zs92ySM5q8Ztzt5PTOqw2veYTk4srddq5oHmbSYEzeuNaDPWnbbCyaaTb
VwxZdpfAcUu9eGUSa7f2IRUSfLccRsz1xnrmQHqlAvpdmy25kA+cMcZS7h2w86mI
uZiSprwqLJl+S1JLSE9/4frBnfWQ+8puLsbNngfo0pObIpuWkMizVguup5+s8CJd
ADTakearmLVMyKw4NscPMtohJVrLku0KhUtwR4Cb112IbxB4jFsLfNIGn+nMVmcu
AjZTFpEIKPaHLLdFVfoXoabCEq+6rpuWVA61Kz5mkYR25X96MCEVL64oiEUbDhPF
e53gZwaT4LiumxfpybNGhD2ysCQzCBDBHwIUCP0Jb1idkSx89D+oC7tMeZDk3JMG
rDF1v/i6tPkTEIvo4TyA1n4ZacMpRasQM+TysWnad8yzCiBx3rxF+ELg9HCvV6aA
xQQbPTffoYXxiQEzzFQYho4WxjQDkBDdbrnYMZ4d3ux0rFr2z1XY1bMU9aVcxSnG
0ZHrhH+P8yeko/x8bQouzodpHq616A6ouuQoZ8G+daw+4cxaMzZGSIoMbnKHDg5g
Rcpt+v8SoTGWXwHAIOmlAkfrA7Y/4kTA7INlWtwARtz7bvnxHWKXgDftKgh2kAN8
QoQELoLquLKuvsPLG8ckzc6o1zvabSYwsy8Y7kgEorteXd1mIWdkCVCEXZk+KcYc
EHY9LJaXbyp7NPEI/IFm6yJpHVV4/IE7sIKHKqL94IaWaI1B2vwyJ02s3+vBROOj
2MSg7GuCmB88iPpKLbUuzPQxrD67mRqoL2VdTUoZRV2Mno8SDu5AmXXiOK2n7OIw
dteeKEvS80r0eL/Lf+0DIvHZr24gBRxMxMoBcmJOTvE8HbXFLatqcI1oXeTyq2cf
Q3An7qdy9uMZMx2pd/lCaeLl+rM2XnoG1xSDKWcO+ysHBBEwipoSwzOiZH4g5btz
lsGkEYx10uXdLpLQcoHMtZdIYldcxsRrrjpKYc3rjcmjx+G3tw/Zn+z/QAoQsyMM
DRlIpVlOZDc/2ve54vfTTYAlMrpE006dlcHYS/d15OQTr6Ww2fujpCrkINN9rb+w
MDaji+c8bkfcIWYVekc3T6QZemWUOgyI00s01w9eX63cv+IIQhqT5iwv6fDDt71u
dFefVin5lae6kv2a4TZUTLRkoN0hGmrcDpLND1m+4SJ7r3UA0k8Oi2lQvIyfPFte
XHCx1z6pux0pJT6319rtWhJQ82C14k32S0htD25hTdTebnafo8jNs7HRPcynAGLG
/JS2Q+CuHdD3wrQxk+2ZuoA5ub6QXER4wrgZ6EM+2vBxIXK4mqXp6SQ96DJuS6W/
Pn6O4n5f0VO8VNbGeZpaVKRNC364rYDKeSw08D3ZLKJ7ar4DlVYK5KhXqv6g5AwB
oiT4R2rrr7ZMG9rZojiSOy1Bi2AnA24tFuvIlRdMvER+h+nb+x1P32gz6zlM5/Qo
Rfz5a313JRbrs4hRgMwXJc54q/QoCjr4Ce2lqjzgrOiPov7bVcx8vngNHqurbOP2
0InAJ/xPdrE3L2nGQXGtKu6ZfLOSP9VIO1ZUxIYWDVWY2XKOb5jDzbnkJe+DTKMq
Kkaj4nbc2mUYhiRYQVQAzUSQE7zM/SnOcq6PaB1YWkuvAt7l50e7vwxIF2cEXXef
RZJBm+yd5pFmKuCNRhEX11NVRYkzfUF/tLkGH2LJBKzMgXBbdPhC1XyQYDuufGWR
DXAcbu2ZstV2+cqK110lX/pU7Bge5GvYa8QMuH/ijkkISGrQd0KmnrpUKORXTDg3
qOlHIWmuIP196aEPJumk2iXxo0tCKHpZ8CSEtTBM4wgVYTzX4BIsHBDdMpe+FqI2
Ad0rpxNn+V3pmLO7C74Hv9n8Otn10zmNRkpaADCz/I2gTjM5LRJaNcupA6uzuFrL
k1FjcxWlzCLj+JVcNrR6Gb3Or+uttgx0TKKSNv/8kaIXbPdfqh7J+sUYwRSrm3R6
3j47FpDGdBDljBthOSB5z46nYWqeyMzq+IjFpSxwA0AXnVwecvvRFmiQUiv9k6sd
zQhsgpQQOXgIk0gcwL40J1yqiM5jY0DJP5ciTXKXPoSErIRaod7BLdeRb6IbI6Uu
G74hs6fnCZ3XtEGLnfs52gYaBGZ4d1RJgctByPQRuHJm5+ElW3Vm7IsXAkhOffVA
7VPYJGZrK5Vv6J0hdSrEeic74rzwIiUe1R9TAKFxq1YRwwC92kUDdoRYHwrU7/AO
/+jGNnTUWbhaJSECojolKYCYG6dqqfHbJiIC2zHTdNQsk7e5MN42gXuydLCTnjn9
GR23kWGmUe9delieuwq6S8kdS3DDn4yeDBJGxl7SjEFH4V1MUB9VZcgMH85J2UKS
rlJREoRr34yPI5rrltq3lan5z84zgk3OuadlwTDRZOq3K8BkEuE3fJM9UdpipRCb
25TINWWdly2yml7s1uP9mgJxxWDy3Frasj9AJ2VtgPYj3X8KrZEi8yC6dTZ4REEw
vGKuByWxOysF1myv3Ko+tvtux647sbR/I4bmC4UnVx5EwC8Jp3YgMSTRwjcswzCL
ixjEgL1IfHdl04bkLV9TF8GpaY195vvCD9QQZfZAgDwfcJdDbP53TZfxnjDulJHf
zxjJqduHFC9QGYuxsumCBHIZNSqR3xH7SUwu40aG23o4akS0oTQ+muunv28oDJtK
J1wpccrfo4KeDcn3x8ZyJQxFi1hGGFBn5jE+w8pY1gT4VETw8GymvDm0GCWExM3G
U7wdNMlH1+aKIzG68ZAy0hagl6TBPbEhjtBc+Ftr8YP/HQA/Ixg8pUP4WPYziCI3
gKH6b1MEujgY6ug0fSwOlVCuannLpD57PhyyUpe1qlLSAxkILtkrg89sregb1XkT
DtJXaJOZoZ3weEa2npQiNCOMxJxFv7G0V4cE775vT8e0oXd2x2QGZOm/SGS2uVCy
09DM2dPGkEq2db8aQc8jCyJzaqMmtl9wdq0ZUlKAyFps+feaN1K10K1dnnLOf4kL
8jirbTXht6ZoOEn84dE/QytDP5S31AM8G62ecI+SL+dqrdR3fjJuhHy2jYnhKLK9
rYoChCfK2zjbh33X1L9YODUB2+BafYrxp5ua3WjvY7WUi5TroE8vQwm05ZomS1lS
OtyhDZHZYDXApP/PZwkO/RCOy779+LzfssIgYjOAnDR+pGBHuGGpm2wjSb/b0gcV
XWaiPKjFIDB2B/xjJDHf5yzx8QptNAlTOWx1l0xL5ZU3lDBow7vbaAlPAmNPMBcQ
b90hV6ZuDDURzxbthtXdhx7OtqrEi35/XhifwnabZaK1pHPKkNR44bK1J3p/K5ej
ZvaZ+guwvXctFAVQy4/TqUf9Tyf9/XeDDcpZ18nGPa30IjIK/dNfl4aHf66KK9VP
A/3C2ZCSHvh7J3SoDnxfgnE5AtwztwSZOa5yJbXMrtwwH/JI2k6BU7/3k6LzbtYP
pHPGqshVzVORw5ZP6H6doAlt8y2e75oyORH6ht/4hIPPVxySPPP7dGozzggkXKDK
zbydEi5v4+t526O09lixPZUMvk7LfV8Bh11jvUO585ntG8iZCJml5OVTW5l620CC
EOUWrpAiEoTPgtv1coCekIplt8zneLpfu2Z9P1P1bpwAprHt1En65OxXSHmECVzO
MDZs580ZQ9Ku5RepWD2bXjpu8Gf3yba4eL9Awk6gBKnQMraynCsIQ4pIBtrFl1Ir
BOolUqBjSdL+pxiWH239ZEWw4lVAPd22fIc5OUyHPHxwvz0jhQBVV0PGHKF/Bplh
zXSWc4jpwRnmDhQdUL7Q0YnZHM6cv6JWj3CADewmMXMrVO6VKAwbJwfy7/FrowZD
7TkXiKKLIvjWaXB+rzoZ3QNO/Wp/rZjqOF9HKloIRHVQ4WHKnIXs3Epm76k9Fclm
RQOWG1aOHta+Hv9qGmqhNBQ44Gbwourg8TSCxBsA1vHGt3x05L9xjeoOKfNyJIzK
n6er+Z31V8c7yD4k9lxjprtpyWUDsSm1omk5xCr059HDusYj6I81VNgglGy6vTgw
NFgvcJpn972eH2Q8gc9Fgazcxyn4JhZP0MaJTPulQjc6Hzo1ikPh92WT0FUXCV2p
y4Qlli/PzaUgv+dYsT5tcPhewzq6AzrSEq+XN2klaItoH7uzo3eofvQtuLdZqdb2
9y0vHitb1dguMby8iU9KEH4vehaX9FNFn89UMk6Gf+ZCN+D+uNai3WoA9XyHkCy4
Ip1kolfttweGg5/2NOhAmEEtSAOqzsDyj5QsW9smt7/yr5hKVYYRq20YFQYe2Opm
ZR562Mw5sZOgJtBvd32kZBe1qMsCgzSJEGNNB0gU3E1UvLUHrK2QlFboAmysx0lj
IQe501Jui7yEQTEHfWsFH4Wzn29syI5gCgzudT58AEGLwX0dqueyseJ/LFl46tJ6
h/EkiuHCTKnT0LsFioLrh86Lxpel5xUx2FqQBcUjkocTKEiPN551tO1IxRjqO8Wv
GazUR8FILGIyF/dfgfjMkdhLGcHvSphpR0jhPDSu7Gx260OfI+cf2WA3OhKhmbbS
lTRr+AWFoBCX7vgiTYTKwez2f9r2D02/QhA+q/ELO6bVEfUOpNCFe3su0H1X1VUQ
3RNjz5TDjWbKIjukSY5BySaBP3Lkd5DnTQ51TMWaodfb2S+7QVcfCnf13a1SpWyh
sdfS4hq0zizhdRAMVKAx8VCVfAEg5hIgENJtf64P67tG8/jNvo1ew5zn1Izlor/1
DljVJ9QXHdAUA+gDM3LwKO1j3l/vfiBzT5eP21bMuLYVUxkUQ9fjAlgbVCpWuq2q
bxRXjYaIz62EkV1mY6IT5x3AWPW9uTaIZymOJuc79O5LTPNU2x1driyG3lVtpW3o
lYhTcAd6AfAQdtTfhd+AOFLpKPUN172n4jP8wyxom2dns6buB+Au2kahCF8dhtuI
joCNaimMNBYpGAdvGLf1kgywCb7viqmgoOGSC+YuCmtVc6DiWqEyPLE7lQSunAb6
kEtAT+95kyRr8yu769vPLcnA92ZW7AsqJxRD1sYSmO8Slu6DnVAaKhAWhKYSerph
LVtrXiM0VK69MkPytzVAcMX7e8nvdQhZQvVPyOSR/0KOMLiRfBPwnwUZ6VjoOOI2
0ofv4lSG/QbSg9YKGmE9ib3IoifLhXy/4WTd6dXjA1nbULKMaaJrZL+bAsdmPIIy
Y/jMTQ59+ti0bcFdKl3X/438lqb4qIpTe4BrMbfUH6useFEwXKQnKxUUMgfDeW1L
ZOet+QJIe3V+//1RrinZ20McZESjdpmMdvxSr2flYIGIOSVVD86lwVtlahxj9Ejz
/SSg4iL0oh3bcD8BaFqgiZBYklP9EB6GcjxXe1pHnbUKKYWKBhMZ4gHVxHZtx4WF
7YcEpeGDzU7EIflam/Dfkc1LBanX9nw874MlTEkvkE1d1pp3XuORyU2jWK7JIh4N
W/n+Avt/1mQI8oXf5DD8YfPxNKLvw136WrLT7n+WYOCvIIHp7nfG3/Cx3RQgTp/s
AVaCuYd1154NJvUsqe8DX2ev/+31gqrTNvxXiqEy6TKCRjUGzx3zydSzBO+W59cx
D4zjuW1rz6v1j3O54gdAtNAkzKaTIgMh22xr+wfC0MlhSQwwYAU9LX7QsUYnve/y
wR5lmXOhSZ+nGz6REy1/ZlckVTnHi6a3CAkR0TxQ3MpSU/L40+07KhuC2mp5TkIk
3XqQ8rBedz2S1PSQo09nTp4vZFoUuaX4EBu0VSN+jDgBbW9H4vCTqt7V2U6pQURC
IcC7ER0tRplCFj4L2eqkR7ACkGmF0QDvcBPyc2ZlF6xWA5rVh6Jz+yMeIpZYK0B7
7c5ST03VZyNmFOnYkOmTfnAHbp0Fg2S2yqLHbvr8Rzrc+Af+URXjFHowP0+rkCpB
vEfJfasKZTrt/97Z/uuVV4g9HI+kgmmPQFu0kFxBtJfEbzo30CmdP0z8JfG2xano
KITP922O3C5fJOcn9oBfKsXD73Thw3Syje5+l0+ZNnz+/f+vmjkC3HhWo64J6lhA
aFqLLV/1If8GI8V9YvX4j5qz+dmQF/5B1CShHDtVsP0+7W3167qj8txWKUKp0NAQ
2Xp87YqcEzu0c6cV2B/wG6yghYfzukHOO4XzgJLtGvFMCIzt6CcObVDOMz71eZrM
0XtJ7+4MkaUp0p8cSm8+ZwDTCQCdhQk/ki0EM8Xf8+oePlCATc86bao9zaOsl0i4
bA/Ar5z9usJzFlA76LjGbfss9fw7RGN9hO2h0TKzZ01ODS+Gp7+De24yDXailBgZ
IqPreAPWJYhBqaOx1QFLsEGAde2ZWV/uNurgB1RvIBOUipu2nnV/dcyiMiy0ICgO
iK1eOBrke7YE41iqgDPe/mprGMu1JboKX5l2p8lcjya3J3tWwXU6Z5lGhxJDDfSd
dyzgSXwrXQSUcdVmlZXXTgFDwx6jvVni+ZJyMb/7tT5tOj6uh2adphXogl0Qd0Av
e3s+I0FDinEJwATNGqC8+vX6yXm6nCzGDPPpBRqwYzoBWAW2I80xF677MrMwGJlI
leMe4uKx0ytU+AsCoFusvlHhUzKO/v4BQAqyRVfg/Q0N6eSZiWVKkuhMz5vPMpWa
fxzHF3CWPayxEPAhxVjnMUAPEgNoEaPgbWLOmVcc3ZSqIgJhSLbSRzdfPbhQdyjC
PmJ2Ggns0eixhJrHDyT0X81nXxH39+crIf2IYDRwUEesD3amZsoicG/AQLlchU8/
O/V52eMLck2uPLZLLNDVPRxCPminAt+JIQTlYf7fg4pKpXK3yI7s2y/GVb9NxjPA
Ovbu1i8faSBK6t2wElTIgEPS7GplbrPkylzJL/F4Q0psHAkjvaT1+NOIsvKIX5Pf
1Ii3bz7R8B4NYXYyomdHryqRkGQLtgbXR9ePoAzcVVV9j6TeiYFY1Sg9j59q76D/
SIWGU/mNU5rtmykx3t43idXrh4FYH0q4OpepcfmUMHXRhBGRmSZzJKd4Nv0a7lm6
QDGD00ntW6R3Bm4qAU4Sg8VPfk2KB+E5OUB1+rBQMNafvhCQhbAtiRTochaUqXJs
63IyaN2aEyrjJ+har4rBvvV3RxxYz7yKqsd1fWFL7rjbnqKf9hPzJnwlRPvohK02
t4aff+Grw1RtDXWGMQ5kXE6HfTBVXnNGzf1e86m4+k/7GtmD2b1ltq2CGOgsk95o
Fvmj9N3AfeoOQgo78RL26Rh95QqPGPPllk3UPp/Jw+nY6ygaGvSk1sZ2yQqzNrUU
emujOhOnGWRzLX7OsFzh0FawfiZvQz1aUmsecabm3ol6ljtN6yFqh18xRg9BQkQW
/uQUwO2BCT8DwTFRvSF2LUzKDriYk9Y8MFKJKZecuTsNBGYTct5KOO3bUpcgT/ql
j/+8YvFNf/fiwp70vSON945p5y26DoN2r8XeO5lvK7UmTbYlsHjBaJ/pZRHb5CTJ
vdnHc85quXRIVQ6Z9uynStAdeF9PdPiJqLZc1YpmpEFB7ycRmJoIKGw15SzfWjN8
Hk/yVeK5Xw3Isy0mG9Y/yM8T/V590tzJrf9sSYnsK16mzZb3TKOYuRZ9nZFnYz5J
Vzo+FBNfOYof637j64Aw7OzlGv03+9sOoofFQpihzLz6yG3jaxvhR2sINmpM3pp1
T8s35UN6XH9cEfRYARFy/NnEr9pxtVTk3lccp7nfxVsJ2W3lBczcEk0hpi34/uiP
6FiMMZeC//n3OIJSX8hwso5eg+Ddj4haYHyvH9f8jHtEEfXLEsBOd5tYn57COBEr
yKQkIwyyPr1QEbrc5UhjyiKU52IhywAUSIRIW1igQkSGebGv/BwvYqjySUCYYNOX
cqCwyZcog2LcxCee+EPKIF96L1NsaWDaJR2XyAM513JD4l5RYEdEaChZkxQXn+TU
lUVLKyS1Nhwi8XZnBTbcBeKyLMdj9YzEqdmpHyfb26oUxZ4JfPoQ0cRZ60JEhlHt
FnIkDnO96vXE/vxrxKs4BMGDXl6T9KGYLFJKFuGH1dCtiAg0YWADcmOo2FsDyjC8
hk0qGfDwPeGygFO1MxB2MliJUSCharEdEWP3h/R0fu6CBSvlC2MWvTb9Tb68aWvn
DOFQYMHxNQApydFTHM7BVsYZMJSOPh8fYgN/XaleFkLaqhRuqf/yR15JO9JTNlrB
LQU/wwaHOT4kGfYdIYGeUg5e29qoFttQvl7yqttpV/9onq3P9mm43Ne+gCw/YwtV
SPalHbV5BiUTP3hMgeydUOcgj9dIKO5R3BxEuEq0p0WvnF5m7fjfndyvP342idYM
8LZfrC0BUs0/2wWYLIrKKO6fhumvfbPaYrHNu5SuorTHWqwxk7jHNh1veiMGBRSe
1R2MKQxWxTel2sdN7yqCFrwWP5U/WG59NLKAOIkPZLLGioOPl0CE7u7rkbiFsZaK
SAYRs2kyeIBAGXgLtKWxf1PWPRCqdwbl2ZJn5GBayi9PTOkAPpRMrtlKHs8pNdY9
2YyMC2u1Y0ZjRJn6DUUNWFEgHgNUzrGZKBB7gxynUhIsjIRF+4Q9+1Cr737u3zg0
FEi04/c6CKYorsQjyrQxO22lyAAguZ0PYTSHQTTe0aG6s+24/kWzwEFUWgKb5Jtn
PBSf//45cQ3NcibLl/s7Qr/TROxop0dQPD0vu9XrqF+K+nwZ1mtyA7oZG6qyafVr
KcPX2cafJRiaqTEw6FBD+neTqABDicNcLx1TT+rhCBvXYYXbzAmcWmz62AdDiCC6
uVcoqL0bbnM4WnUdywIMSfOwIo84TpcXhobO54xUzKdhBuVwyMW49/1ytg+aLBX1
v7VCPf9wHAxFWH0LxsDI+TRJgdzc4biEIGkxr5u34ckpl4XJNQTPRwm1TJqElXfc
BXsyi+QwyPkuhNoxGEcomFrK6b2s8Rwt3duDpuYIgsz98C/1L5PIRn3VGYdvhg04
7xbR7QET4s5x5Tknnjrpb/G6fvMjI2wgfA06xJTwaFLWFFCeE6eu32icQZnO0C47
cFXpKsxvdh4lZRgBP1wUviDXthVsOR027RBxyfPDFU94O1Y+shxNlAa+J5jolWGZ
nVXyof78tJFf+w+yZZi7SwexlN9MjEjiROdGs9qae99FotVdlhh3Px60lBwXkK2f
HKl1SxaoNpRhbqjBg6dUEp+8YTXh3WME3JA9VnrPTxHicLhfmfv9AQpCy2Z160AH
qyekg9OE/n3DEoV4sQveEb6hr/b2qOm5ya/m9LjMS1HxHiYXxVlr746isIs7Dxqq
w3pSJ/QMd/BWiZMVV0FyK4wo2AQCc19RwKEy9hOrK3Sp0UzXjEiKa2Hr6a9gq0Gi
V4wNUM1nmN4NFvRZiKh2DWaauelhw504LCKAZrZDUyqPuVWm+hOGgg36pVGIwZ3+
gPnWoqV0L4hD6uEmh1+GrqxE694PTKrWyKglr2IALoKKCAzfnoKmQmKUEcI/06ci
ce78c+9Huj2z7RoBBajM32YzqwrUEVZ6bj0bCK7y9tFVXyCbUnOs9rnVcsU9yFLi
HHpAQc2bbsZRgwiEEXY0ZMM1iBdBOC1obVHbUVJYx5e74Fj0Fn2vCFs7e8//AXY0
EGdLjUjVeMBt86P0zocoaCy6WzIPxO0IdiBtBvUD9qQ7eBmaKfTecDQilM7MABVZ
sEEClQmzxE24qdiXUbKLaulkkVyXnOv9WnI4gqC9DLEH7pGbYOZUx2YCptpZ+ljD
TWLE1sjavY+pvfSsmdhJOTN+vszhypnMakjDEht8Y7U2giZW2qoBARV5d4dw4ALz
gikdj30y03lZf10g15yBEFIcasuHxRD86MEubPLCi3JNsQmVxs4cySJBSqYwaJb5
f3Pc4wA7mzvaeVw+KXAqFnuPsbZ6oy1sgWmS3VLPG+CSfG09fg58cmo/VDJt5rCk
eNXc/Ngec8N/357nNM3eVPlOQeaRBlQllP/L4nDEaBXE4WHZ9EYni2ETGOZI3mmW
wru88lfSsPYI/O8aEDhH8Agwgk4w4ypsSPMMNVbcLBGUgCCXn9Iwz1kMZ1N+zb2Y
l41suj/oOnWK2yPGs0A6ZcxbCnhqI69UnPZOEjKFK9QT2d4yFd9mukap+CmMekwK
H20rnYOPrG6wEo+DucxEdmiedKCTWYIqdvIkGmFkFToFHOb5M1RxhdUH3WH1H/6j
4e2NTy6oqUifMhSGccvodkEFKmuprj83+S76PXeH+1n88Vus1/Piwenhj768aWDG
1LwR6VM1M76FDNINQEMLQDQTkmrdMWs/KGfRA8ovEPNL58RXXelH71Pl8IBmd7PZ
pF5o9WXTiAvfQ+emTYW6ZmEZpOsUcfGGFNZTALSR793AzpYExxerVTozUnrak1yg
HXQ7X82DNAMebpERerVQ574Qt7naVZWBOcxD87aSMbbie8EcywKmsoIwkWF9MDsA
Jahny6wxT7rAHz85dOIv4Q==
`protect END_PROTECTED
