`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qViWvHV4+GG+KsupzsLMDNYEUmK8NoWSz9l0OM/NG3Ed8qsRoZPJM1TgM7QgGYV1
QwyjffWD6KbefDTbI5uFM73GtUyRFCBNXL7rxpyxnKBkdws6zjfqAxR8rgOm8HkS
D2udkYxNmVmBfX84pjUiOCK4VkokiAwY3etrDU3ErX1nky8kZGY9iEKYxf8dsMZp
Y5lClDZYyjDrCZQgS4F7ztHK8h0MZVg1PZp/ipqKltXhiyruCFeTyyTFljhb/nSD
RGhVI40NSAqg+/u+ZCZdwixfI6PJWXBqBVCssPDPTKYH/RUNw8DnEKBqne/Lc+8t
8k/B6fR+F42VsqHJ4eoHkn409zEoR6xUccI6+XJegC91fhOqTlS5OBi80U3HBLLv
QhkouQzqb8e/MTkLCJjogm9Nsv+9BTqyIvWcadcj49v8tgdMVS5AHaXoODcfIzJE
cIAdmfnZ5t2rN7V0IsRvJuJkE9bteej3q0NLYE4o5jPper1kQtHfC524V0mQbqqN
GZRIy78MwpV6PATDneuB6awAEyGpPqUAq2JQZlc3xEpAGFZc648ZqKqfuA+IWHhq
rS8gfTsCB3oivS6ivXkoimjmDTQYNtz/5glDF91HTqf1NRDNiTQlGvkwHoSSVxuB
JtuCRoD4ENnB8iRhCRknDhGxkTWfMQASEoNHy9NqQMxKsxQ/b+Jle98SEPOAYziS
ggFDJLzriE4fvvDpk/qLBRT8v6o1egPIKNnZf5t20mtUThzrYzH+nReotgRHZEUX
POcb4cIv6ahxnjm2aPfxxjJne8Sb5mPXPN3i+217cPvn7MsIV6S5E6HaooC9au6X
V4I62jK8mIikz5nzGjCFgF8A9JWoAD6tcMGTDP2cJ0j2iYqUpuFyZQt/DitlclH4
BZ9wfyReiXweEqsWSpHE7U4WegjWSTgyoHIUqjlTJmTTxk11rvwwlx1atiwSW0dS
nAwayk4l62feqntQBQxRpXK9AAoZgun6sIA+dWv788UIpew8QmtQWEHFcZnwyvEl
hSaRxpEN5bdtR93NX3u3LAmwjaFR1m5XATbyifMyyVIDrZ8GFaJ+RTj+yW3m8X28
V7wUyv/8GvZ2iGBArpp/YGYNYiMeao/b4lYf/rCh0lfP6msRg0v6dRIaACeA2Rh1
0Gq027bMRP+RmEbalO3xgFOiL6wQTvGJA5HjMRsFakFyKUt8U5Nv55+k7lqyiDvN
Tbz3baLjPCjv07GoD2YD5vneSMGvyp1dGPBwP5LGCpflH3DVwGcfGJkXYLPR9FOT
ogfIanLOf48J/YrAp6GXwI5URNsEQocZfseJ0OQ2ovNjj+OSEYBIT/AiKVKjkPL6
NYY1evk1Xo60TajXYMsDEH0qxv5Oig/bYJ4528DCK2Q0qgEwuLnU1K8ec/NvsXuY
3q8k+cf387e9/6oiund9THoXzxBkS6pyt1Lxqs2BsU1xKltqYcX73Yi8EjNX3zCG
qkqRAouL/w/nKGLaGFu+++u3G0iK2K2STSH2pwrX1p+6cFA3qxE7p6goj3Gs2sEg
Ibi5rEWrkyeERoURV751RawszXLGy+1d5BeA7qkc1YDL/zP3KmW8+/VJCvvbHio6
252/N8HkSf/U+sjP8n3E70EOueQJko5j31vuUU/XKgGkQLQaE8iXM3GhcN0TQkYd
Q6aBFdRpVl0ahM0NyK5PKCV7qCua7rkAThCdIRUzlNebjrHRJGh80djXpBbInh/w
9L0KLb64/aWu7Z6FHf8ccn7XvZFBx+MsUxasquuTxcoemfdnPZpRUaIifAAgPOSY
yC8Dii9YiJc7lHu+exZjxz9tVipqKbjqixGvdUhgFbFDwonCh25//zqk4CQyyMrZ
4eaqZh9S7C+UzAXOQLYo2wZ8ZkehLuHoTi2FrZjfnrrx/1ARPoqdC974yW2hjyI/
Yr/41fczzFMq2X66AReXzOBNIOJRiUvd8TKqe2DGCkhPJSQQ5HsUDGYwZE2YRwpR
GS9IGNLVkzyREcRS824BfJWJ2+YATdLFJVN6OmgpUhaKiBPKrSC0g0MRId3xvQw5
ffsB7BT6Pwyu02FtznJzlsvfJIfw+2seX65o/rQumcOL/jMyqjGvNmFhASAm1bb5
K9/4AaNKWyft9R2xc1ZzLXfvbdpM4gECwSgE0V72ZpXUo+d+80MKUzPd5EJvVfV2
Au1o0gFL1zSNEKBomb6FnE/roTnfWyyBIlpqWJmd8yRb23Gwt8HLxzxlkWP4uyYH
2/AMe3FPrAy+FmKpIa9CJA4vKjHysCZy3nsV2W+UkLLxwDGO78MIZgI02fJPUukg
xrsEG4oid3VCJnrzMvEt6mIRDM3Igy/OTZnBIMODWvswwruZndDFs1pvpUAFQn0v
vni475p8rUXu1R2GyADRFZYDP22NhQol2gYvoK6qNlCnrE+y5LMweojgUV9H3eW4
txJkeFB3ZgFEWREHzullan8hNaeStr5g6C+WMVLdDZBQq8bPp2TCcWY8Gt7TEMJl
OAQ+I1ulTdW83tJ3qbpCHQM0en2ErDnh1IwIqBNI5XEfX2B9fqVmGhKWeUu015po
mI9VuTF2Lg5C0EeRX8nVB4Fo/8Px9fJMDHJKu3mBnTxK2IWM8tKtIi4+Kb+WC/2A
v1aoROd5T82+k+43X1GtyY70bYE0ZLZLxQN9Yrw+zaEINeG8ee926lHAfJJukD9y
zoAPXkf/4VHFvY+yOV7gVfnvv23QrJPznKBBEQdB73QxCXTmvqmsHfZXwZ8LXMgA
/yytwztvFq5S43T7QdkInG9PFzTyYHWJIFYlVN3wXka+nTS/gms2ZgaJLbqnHx/6
5g1yQoaNyzNMoDmMC1pL4TyaLs0GeCvqW+HTDM4AOxdMQfHETzC1iDbLGOeJWm/Z
humagifLENrmE3htZS/Iu1leVe5vfhS9jUAEUb9KJWDeTbqxfgZ/aMiBV14nD/cG
LrBy9yf3DGsQ6NaiEF6/VdW9Ytp0LJ4iMUn8o7eFhZPg5bmjqoMs286kdcgP+9sE
R6b3IhpKcBL24EHqBJk1jTQTrV7dvUyZ5e03HPf6aCukBDn6nJ5uMfc8JUpyWc7C
7D62LjpoEj1rlP+cf3Z+7eBkgaNh09cC0IFZu+ShET+mKRsT5FkMQtfiotsNDyAx
zcP2e+4fL6rmyl2KS4QoGDtM7iUryae1JJ+bq17q7Hehn3YtuqbdxazjnbCunjc0
nD2EqvsV889cMz7tjJJ+2G1dmq8wxdllzS5D50WrlrqB/HMeCnOIEBsgpbJVfGiv
xNKPw8nh4XdgrF6hicggjGOp15DbV5v6cYASIXEVT2mBjkcDGcE0JwByqaTn8aTa
cYIdG9UHMQFn6rYhMX+Oc8aSCMw+HnXlBcpnhU6t3PDeFeiD46/HAuW/kE5Q6spL
c7edzLCKvZcGnAG7hCm62ynpJxH2WwmSsijxblxef+clLbOM7dMEJvC6KTHmFaw8
8jb4fo9Xfh/xjTvg6ZMeKglRIgov/uf78BH5s6E9TVty++LWVuyCUhFm62bFtj7s
COmUFLEJPx0AT5446O7ABeGwJfrGvO9nrCE5S+FH3X2lHlwOIUdPAtxIiniod1xI
YnYqxZn/IEyOByRV65Yoy6V1xMomGx9ZzHN7GuNaE3xO8n7S+PNVNUgEX3TiB9Rt
i2NDBVC6gsBYKEsgrYHMScw0JIo1rrOsAJYH7R58O0TO2g1k7EZ1wVOXy0Y4pK6K
wU1904vaHW9VmP8YBGzOBUgEL2FaY/FIIVyF7wZi3NyW1LryO+oUPro8Q9n8gJpy
Uzg7vo+hiyMhInkoqVph2jYdikWkonTwdFy02uB4K8eM84OguL3pMRjE6pk2ylbu
1+ANm0ZNVr64dPIunYMV1JUQQaKwrPpxseOhZ7qzaBBdbdIo1cx8VehV11jCaMkI
0dNQNoaJ+6zMcPPM7hxpEdCFqCeoKYX+37HCJrripSPl60XKBcjNUpAWiree3Vb4
miL0FS1/OOWICVnA1NXG1SLu6ZoUU1FighFBPmrySM+Ve7vEbbYBJ6oy1Ejig8MU
jiOPacnTelIcqrokKP/RlZqRVFfO1XLjWlKrDLyxEIaK10WN+q+jh6rRdgnIHM60
eXQgmQ06w5l7UmGbJd4TmrRDIYZq+fVkQIXfzLIiT4koFsjrhcUXBYs1GAymLgaz
dW4xlVglpyJjrgySOpE/kyIc65iazbgQL9UKj9CykSxntZu6ENCHtPgUjkT5wFYU
0x/BNJUykWvSuyGmvfn2ri0i6DS4gLqk21E4Ky0+Z/FFl3ACPxnJOSGXvZwKkO9+
SLmT75ejPSyID4thgf9Ld/C+f7WN2H4yl2mY7Tur9rVVWFMKGEhpBnjwoROGOckp
drEMPiZUsHCbafo6lg53V3CMlpW2L4myaabqHyI57h+YhYF2KjQvgaLFZNCb0+pY
uLjXYymbo5EWB/9u+/wq2R+8ZkrLJqVt1t3pajIR09MGFZ61e/ELls5/Liuux+yU
orhePFuvKSFkY8wnrGaGs4gP9npVi2FTOiSnApe+7usLT8pC7KShU0rs/j7VRKsi
nmgcKu25qSOFe3BY4f1ScNSF8h0KbDpcisbbtvhpk2SQuRYfZ4TIsa6J3A24aNS0
D/wWxeqeMqmzESzeLdCQ/UvgKemk2P9yRefTrcfHpPfkty1oDjJftBoYX9Flo5+K
43xmSTKFlsaXArqQb/qQ+jQ0YAAOGWWz/QA8ZPzu+fAHtya7NCP70jlF+5AFgpn7
z47JZE397oS2w7EnhIep8UENEtIgrduqGnQJIZfJ2xFjTzyEH8l4hFEYrm36/Fce
ST5ghVhSwMkBm9tmRsdTW3H+71x4ga4hvgkX/uJ6oiOsbXrVfNkzDYT2QnvpVlmL
wHqdznJE0tLQqkIqDnXNEfSJtM3VKEWJBMAEpcyMnHrwfD7NCKmy94eHTvghPN5G
KByiG66H2cItwWqFisCY55QPTi7Ei6ErOmVVaeYD/naikm0UtCSvVwUWaKrrYMn1
AgV12DPlcnC2ce92RuL8DgHcOtuAq7eE4yoeaXIEZGwRpPQDoYwMNk9lWZ+hk4P8
UsHa61MbtKpNdUkbY9ZnwfFithNCHmPlpVRnz8hh7W/ZwIUWLS28DaDdVLA+ZVZi
fLDJ+ULkBiewQ/ytTM/Zf8loH2p/PBplMG6GsWZBn7oKsnJBOVTxGFw2yAbdcjY7
dUcVZxCL/8qXLdlXxnr4imDN4Gwy3y5IDuQfWFQtav4GBNUWJKDVJ/d8eAbIw4/T
4kNDqsQTswiXPXJ1WzlNVxazkdAeTgDRZRrXnq1eWU3QWmlNrgK6eQ+MEsxgTCsa
SrtmiwMmZE2swoLYoRIFHvlNQwX0ctTvy336zgI/3dkn94n1FX1pnZQk722vInYn
WNWbdfHIO8kEEB73zbSlPjQuqAJQ8DDca2CvLhBcDVYM0BLgaZEJ0iwve2vmpvUV
XngxG2hq25IIjuJP4Kkhd1QKwYwFvUZFNXA53o9VaI8wJYEa4OHpYxjmg4we3vW1
ALoZtEWRFHiSdwDeRK5qZ9WV2VZtXcnrG8Etgi58/DwUeRoqsGNJQzghzJT0Rdfa
BHXIQ6H1GSYym90yRUOl46hLl+GC8W0ScS6AboCkp4+3vUiUwTqvvu3anNfqf3cA
jfW1D+FFxz+TaG4PdGhxudcmGwlhb1BaOwyvUvFYzmg5KSQgyqhRgfQlarKlmcFI
sR8184uCS5mxz+qDzUxuL8W/uz+dsdaVF3ULdNHLs6briAOiOQ/Y5nED3Exisogi
geD2jx85Iv/I8LRxmV1CcFoi9meViVuSpMGKneiEzc/1eoehs5hGjmcuse7CjjUs
rr2Ud7l/An/2tF0RuOUB76WtcxxfboAzSIHhzyuHarxFFICjIj/NcC8arRiSq+ZP
Qo5ZtE7eYODF/H1pKd7tg+2qbp5IdxsxsNoh5+ZjOCwP8Wt9brMysYEpDBKd0NSj
ipRIkEIoepQp0zTwPrjFczvg4L6RMUUbAud4CcTducEm3j3ScMG2V5zDen5mzt9X
q9yYJT32AY9DOV4QEB9AFxjVfeCE8tCa72gmXPpAw3I7RoVK+uux0rKRIQunVdjs
S9jFyReLLZOhUVdTwQLiMBry4vqM64Ri5tVTH8kvX6M7RISq9uFbSvf0CGPEp+Ul
zYXJUahL7M7eSgeGWgaIPSoKDbhYtRMIoWEr2QNQCrLhLr0oAKGVQTVqHZpTv1y5
hb32sjqfLluqs7HMg5hvJk6oDqHEsckYRZu/nh6bf+RMuXXLj8jZSee1ok/d/vWL
Heg0dLj54qythpPmJK1HMeUYcHaZ+ryTCz9Fol+9d0gSu5q1iNiwp4W+CJAleLqH
rI8Z2FYYC7SdLGzZD1CS2/RNtSelZ4FW+05Gt+8/3/j1LKBG4tIjWFgpd18IosnO
pBTuSbEpFvvhsxBeGB2SqQmiwty5NedUC7mjryZYqnTFQ79JNPQDohPgcSo08jXQ
LWTI8XgPXuBZfkLNEceq92IjRCekZYN2uVGb4NXODv5Hr1/AkkEa3TWD6KtRTotv
T5uYKPA1U2J/geZ/iGzpjats+LSyhV/YNkEl/3Rk+siQS7xXtNm7EeWWGodj8Sah
ymWD6nvV5hN8Pu65IOvRPdpDL/TkV64HN1+mmuG3nBpGem3eTqJA4VdqM9SKutiE
eSoA2mjCkDBRP9jIgjkakvJ5fyOgAGgpSgQMqkbzd3kx0FlkL64lISqaiJCEfty6
J/Xnr0ygFPe+7NeeJTDGfVnqgjmvg9P49JJ1Yw9RU83N7eiNBrqdwqL2JSbi1BWC
Kb20NIUDsPUJ/QUes0HGbTzF1hu1lo57OsD01c8kOIFXxx2sec3Ngp3DQSwmKCd4
23/TOv2smxVeR/Imf025gzMN9/RILI1v42J9ou8htNvCkcPhRvNl7vZz3YGOIb0Y
aAhmJspIh5HQH3M34etXxJBz/+Fay4b5bxSmhikp3NUVqH8/x3yTbJ/3xYvpAQQK
tJTdfUeGgml6EOh5WN+u7PXCTNzolc9vkrFzX0vqK5HTBYobIKEcDRz0hWw7C+yp
gs1zWfu3gPOlYgKEVNCXeej52T6FRl96mOg6zr9HaPUErQL2M26xhuCvq0Hvnr5L
l4G1f3YDGG2KrsJ0DLKn+Agg8CEyucL73X4mkxbYruAH/TLNFQEUCNCaMyq8Iomc
5nKmgaVM3EnXiEJf4j0d5mZKDzBh0IV5CcMnJIvWuozOYt5Ossv2YZ+9D+M/23hB
P6bQbXoZcn/x6OtZiGRRPydXyDwz+EEx4gAUNjQBPoUqgaCJCjwnQhmu2P6uNI73
TIT3v12exQciMF42g0/v6pfePi/c/YKH1lsSZDds9PtraDvVYv5LrukIzInSxQRz
Iucs3Ey6b4x6d1Q+R6+dkgTdxRUjIzN7lmNwuB/CSTkjrzsgZx3aI98SymJZDpbU
oWyifKucWKsb3V9XzcfRmKAiqmsAcPVRqo5ADfiuczav9p7O+5xfhx18Wbq+s6mi
DANJ8CRKa8+lAC8Bxdn2Q1H/UZ/TnvCQhMksPR80TLxomu5PoF77e6dYIrLdr1LZ
BdEgm/Flo8NNtNPpxQXy1ckRd7XihsU21z+IjlOYyEhXHIas4E97yfF4GwSfSZqT
XuGZYPYwLV4Rm7GRxAf8VKl5tfrPHF8YQNPBT1a3Dm2EYaE1L7cz/M9D/8E9xhLV
DUAjDaEGS4eDJDHc56rNg0ltWNDeL8Xb/IJhE4WRd77ra8bwKsgy0GY3WCE4UBnt
VDwW1DHlAcVHDy/rr8yTd4CiMs5+1+eMR8QCqJ3lNddxzrojJ+mByr+cVq9IpNoZ
EPvsXRkvIdsbBKEbrO9d9hxSYODAgrT1Y3mwXJpTnTq45CO8ZFWM+jX6PO99Un+u
LBrsIQtFqXcTPj9WAlO/6EhVAK+UO03aXY12eSdqqFKSQeaRsvg9jSbmA2BPTxAv
mg7ibImiSJ7bzH1MdohHZqMISVeOAK2XXArjIEhJFrPKZQH+TJW3jVUZwiRCZqoE
IhuGgMH8z6gM1EqPhCberZgoZUWu3S5QLDUwnTeyG48w8JsnIxham9MY8CwoHbis
lrxjytWNFsmshhevIU1hYKNhYLNBWh4MaVmSwKv87Yyw+l3KUm5A4BexzQ6ZhnZd
yvn7ChJjbRKr6C/Y87ojGT4KWCqgy4MPOGHtlDLJ2qzDsrQsgBQ75KdBi8SZeXpg
NdVRm2Avj5k5140yzywceYfQ9U1FeQ0emHP/To85Sc3p2j+XImVrH1GfrW4jvj2v
9DpLLZyOobRNqQcnF7W58ueTbrlSf3aEDovgdy4EvexnTBNYaw6VmwO4MZNjgjLf
n7+yOKFcIsBE1kmbuknvmiWq3YE5z6v/hO0Rv5oEUqXkPq0iNHpyln1Zodw6CLVr
peSxidDvuoOefOPURhchfuQNFsBNFFNFovjKOCOgxl4o8KfSqPhxo07Ty6EI/lYc
OTnz2dfnVK8kx32ogHxP7oExbSZW/HpOfkToSlXt77dZS/bByfgj8pbHpyiQUV1s
tzDdp+Rcl6mnDvDkJVQEgHhp6IeKvD9crW3h1Ay/wyV/O2MVz5NwIuR2L9PcQurm
ALjC6F1rbn4f24tD67gY4eNSaokSqGLiPbGNHTT9K7NeftUpZckJC8X1vsr3I9tL
XlPWpd1uI/f+2X2/9Jy273RxEwsDaJK5KeSDgjn7K2FYWJtgv+JPi5dz/sGKvkkE
L4xrmrKnAljaTnRpH3ohspbLu3se8Zey4WPAhIDA6zdmQ4gS+ef6bCTo9cbZ0fm4
BsemQhilyzDczC0fghi36X2Brxw4iuAdClmvBaWTGc0OQWpAWPD0KGA/9xZB9EXB
6d5woi+fPLmZNMAyzCL1i6SJZOmiz438xzs68W6+K/sEG21PeW+UXzGevBu2OIbM
aVYV+3QvbF6tEJRyGc2REJR7mwfcKQG+KKe1iev0CXxvgU9NT/CiIJj4/Hqn0wN/
4AZBC66WKUFtV5J1Vg7bV7I5SjFuiiQW7ne1zI8ike7AZO7/HfM+MRSAaEO/Qc8M
B+lP7bmzMKcXil8sjAOdfjm/tXqQM3HVCvVy7zIYoz05mYfJf/dOCPfO3cP4lWeJ
TFY3wW/KCFAdIZLYFjpzqWhLnqo2CFICxAv7qGkCSW9GSGfjBiLfbsD3nCcvqyAN
nsdTLXukZgdxn5oSs9OcR0ABed691J0eOkoE1VJ8XmyxLdub3toLxeez8thMU1wy
oIrJ7uVEB2GKlI1qUVilLI5hQLwjUycvOm3q2nDaVE1dQGcTYACHdu6ItxbZ2NzR
XYXTJKPGuNvor+fuGka0KnqM5SUgBwdBYKDC7ZrIUt9hoXRJU0eHcTYiJzufSpm1
VSXOkAwDUpPXibwh8/uJ6gyUJ6NAdVwhEjXVy0urkobMdP91xXMdnvGjEGtpzu6W
YC1uGxVQyBf+h1EISSV4iVMaExALLstwgOhayHXF7Z4upW6xnFG2/BVw3u/0rQZx
ezan7k13LU+ZmxDo+45IETpYdrtIK0iLX0AvW9j0Mk1c2n6rb9oRCtxeJNx0SpiO
+1k/S1lF4S8vY7jPhvUwulDXvbOAiQFwHzU6Xt4h5bUAOSWtP1b/zL/Xrq9sfVrQ
3r3NStS6GKY8ceKMjUQ7k2ES+9V36g/1tGuwSxLHec2JCWnmtfK4/VDLjCyQTYJh
A6lXVREiteSAyD5Pz1jSD8+/ACZIQ8/yohpTgonq273CUY7DKP3anaH8dya4Q7Rm
FcB9XzfoCx22E9/hHjCDjNYsqtRbgB7HL7eG/FeL0ArCqaiQWEKG7SYTbgBeoDWh
ekKM3kpnklB9Z/dYg3zl1CHsQ0Svwapl6fOuYPbV3/qPiFjceEY0kccHu6ENclcP
xUY46YjvPoSLJNCPO0hg6o6PL+wayOtAu0YSz2PggrwsolFnEBomjTS/j/YpMnN2
Mj4ArHBqK1aRKZ9LW/8lxW7EdxDVhj+sU3puk7CMYJANACWUFboUSUKu9eF33ujp
jO0LBVXkUl8h2QcixCruawdcdKdO+WXFyHV4KL46QzgWgynroJZcil0iq0gkHv6L
glxRqdJT8XwmRRHOm0bDSnZgsPZHY6997taJaWpsxAdtYdmHECq4GXdjLeFjHJeF
VxHyn+jo4KafhYgGKP2keMZJJPj/BolpUHhk8psn7W1tceRxIKbp6g1PQDQ4Ayp3
NW/ipbN3PYRO7X2IgjllP0IOOBSywL+TBiPoJjKW/MwyEfp8ZV/0sE4FkL29bFNe
WqkQubp1GI0Xajrl+kxiIvVU3f5iPdrmoSUvPWYfQgm9oNOpVf9HdTZJvyuvaqmy
TRlN/LKa5smFH/k6oIr+PotE2UYz0pfyJhlYs9q/VhRymTbWK1ABqHTCfAO1wXBQ
lR8V7KRgyHmtXGCHQCytPi1DK8ujAi5g9ZAPXlnOzJCUd3eK/n1Od/Gh+vLQp+On
L69maH4c4qSWbvM/ihK5NpmWMSwS2IBO2T6EZT+PLg3sD3oW1C1NZIHkXiwP5R61
KpoR1ED/qGHx5sfXD2W9DWsOophnRB+3/p/u/Giv2XJ6x+4YPVTOzoyGbAGme2Cc
YYspEPI9NZwTz3E7rbW7YZIGQAigmtkfQKr6FTvWW1/Ft2Bhhc4ZqPRMgzOpRffo
zBYFsOvDVefOWuYNYweH/e0+A8OTvUprGtzCMs08H9M75diXs8Hu3JkCdpleESZ6
ZsrLb18CWTPT4OsFrbJSamuxMQO/FLxGF6i+TY+Lw27BjxLzPBY1RdQH85mnEM3w
r7W6TCeftcs62V/w7fpMV0BzA6TDZ9NL3cVSldKyuCBB7dplANdxd1B+oErjF0RT
gS3QzhR50hBXKDysEXa6H5ZDmEVyMGFDwfUGly9jkuvpDYuX/OThvDKoXaOPqyR9
WHCLdEMWu9jmYElat+6vGmu85mc7W7zmgEOhH6DrVqDyQSBFufKHR0hqOyiS8bNA
MzwwA4hTe7WnoRs+DAhQzBBf7VMF/5/tFT5lfLASZ7sw60gN/Rz0+QEj6EtP2YgV
1zWBcuyo7psOXA+VhJAiLbOgpY0NKrsukmi5hI9CMX++EJzNmOB4l5Kk5m2JR18Z
fnsStV+f4jJf36J3NkinolMu8dbxmRZBpg72TQ7UaMfKcb8qOJZtchf0j7/mJ6Hi
+bBQp6fPRd4yK8uOlOxsuUROZVr5Yvx+oHl6DMMkf1QyjjAOI4VPAUo6Nn3chfit
MAWi8PNirrdeJDsBRWlH71jcfWj6eGpgaRYMUsuI2ug9+YZeKOfHgBleoKNuAtai
S5mCs25WtWGP+yWXKf2v8gK8EYmMlTBRgVMYIQRh9c6J0qE9SOsNr1oDJ3h2V/uK
YrJr7Ouv7wtl40Y/CyAeYf+FC12XZf5+mrQQqS+oePOvVzfk3/u9U3lGiPdKL4nZ
f9vEgF74mi/r8E3gbMLjJHr2H89Ox0uSCEWaonL8HLNV90F3D1CUyuvSjoqlBRv4
nTyWuZYt7Pfl+1XihqkLWaH7k1tlou+Oux+FSw6O/8cTSi18/mZMD1ZKNGexKPOz
FxW0NECIV/Fzdf29Gpe0TFMAmAtz7DMhePLrMY2kh0HmrtrVhsBVBM9HtYQver+4
KyqvNRrVt+TzmZTV5hsUXQcb28xnSX/yObtj1Er0Sg4CO/u0kdlksxX9+npY8fVT
QJ7icrLpW9aQsaoJTsFp29qCi9vmsxiWERePfykN4QqOnBB/6fsqo2rimh5oMjo/
vx75xIJuzyUvz/ub6Kv9AWdje/qxlaNd0AJ2zBkuyWGOwaHQekJf7VCutOB15R++
yLcfwjkZ6COAZrD/tDCHxhd9sbof0hTXVPiAl9WhmKa+2wZxWV/5CIVdiUzbFamZ
ZH90JPBjKLeBuvgHYQlHYFVabFoEGFyDDbKxq6AJys44dEjq81LQ6kGeEAGlSnSW
spBkY4xw00qYw7D315UlEzxP9WDIMqtM6+EEOkBTUKwtCcdboMZmlDYCdcogSe2g
3SqTExBlxczeJxAWG4Zha43uQUosRxaLH4DlOlrCdFtfiPrM5Z/haEaI5VtvD/y8
aKRnlQuAsSjWMUxkX4ltTVRPT52i/T0bDXIgiEWl9yuVhzaL8sZv7gFjUpETWPoW
NVrBqwDTnGfuX/o0H+v90mPOJoNKp3NY21Sr/aNewDHMOOiVTpPQ6zEE1lkYGjok
iW6cUCi6KowKXb7gHiGO2M2+a/P1qc02s+SXGC4z0FvA+ixVmy5U+xvg3BnZwpp3
EAqIixaHkjiH047ioFGSHFEB4itFxpLls1eT4gznp4k7SwVhbBuZ5cn3DTv7nWJC
WpC5ht+clo5LeIeQsgxMc10vcEZqtBdp9FHDVL9T9tiE45RH9mIpnKPEDRBPcnmY
sz0GZDctDJ1Qc5YPU6SFKlTdTltDufKL7t4weKsKd2ItWpTN8kfCA0LwTd6+rupc
vDRVwRhBZ3mpsSK1/DTLtUE4xM+40oSOz3UQfgddTJiDE8FQCeQTfGWuv4sgnAKS
kCDbOEyR2xBShp/o7ihcNSpoOVonF/UsVjEf6VVxMF1WCHTzMRrYUF+lRDtjGS1P
Vj9Wn9oMk8gEiMSzoBbkVwXzFcitj7DYfGPle5eP0zYis9ENfMTAlf/+LsYKRUbF
g60jv1KXfCpsZQOEn5h7sJoqV53Gy60ztiMJUr45wi+YjRa5d78TzUZDqAZ0DYS3
SuzyqRpf//6wl18mgNjWh0OQg6gn6oGy/TII3m33t3eVHmCw8yJGf5xOUCj4mWx9
/SGYWdXX+hdAh6lz8tB0jsoLO0n417uTLH26CjfYWK8A9qm08k1OQoVnzwZ2IeEa
/cOzDANbQ1n7UtfEev1rHNA7OjDKBPCultUzMtS4t2qNENp1bY90NIP/G4miAh29
0U8d0u6BsH5lUwi4ZCYUVrT/QnXhk5xgFdIJwH/9f7kdVQvxuXPDEvoKTrTO0lNC
qOeN3VIWaw3D2uwhKDzx11nGPpYMbnpekUkD8UYQckTEca4eyGTdgL6voMhXe3+P
q46rvwH5qU00Cgq1t075wxW50os8Ufn/cIgF7J8H68IDSTvaSSYFA+iMbhJx6Maf
Vhej6LJ9DFBnTJGmvQktEri8qGMsEjr5MyuSDcAglewunG+NlziNHhOXKkkYqsMo
CUlw7lmBwvc0CMOPt2s4x1OwzOs+74u45KgZW9kpyDR6KkT7RB8px1eSaHf3xZLu
ZHT0sIKw+zAZkqzDzOhL9hhxXGgf4ExfabAwp68w4Q00iBItcaKiQqYI97gD5RVA
HZDYcJwPQNdNoaVLehxe7AD7/M8YoE8au0knn96MMWO2P30y/VvP10hvxZe9bSk6
wNxSEhjZtc3t2jCsLf5FZGWzWu7eAXhWVBFxmmFmUbv4mYYmujZqEHrof7SKMvw+
MezBddgCGYaL9jaqfpBGvXG17GqGUymoqGeLnozO5pwQFNf5rPhRUujrDtZNSzvQ
G1rBm6O844kr0fFSWTFIYJ4m903wJBriFcWF1j22C4zy4In26iTHVWmkoArFiU0z
Paa5TG2R0DlDpOxZLgE26cnMbYbuu5t0a7KH6D3kF8u9ulohVNXJHzRlfF8WhKvC
KcYVKToyP3PCsstVT/B04dh6ocrltPlYv9m40yXub+Fn3bz6tGYoatXBHKVt45ge
hfl+XZeJwVFwjpzaoEpB6Wd6oW7xhyT1EmI4HfWl/zwoT4HbbMIyKzzfgwT2erN0
a/ROjkbsEAYmoZW9yoYkp3vQZnl5FNR6SRZNn3qC/3DqFroxbRcjrVnUbHu6i+uj
naMsxcGMWlI1sLt5xVL/LqmLaHNsHUoLCo3dJHN61sIXSFUcVqir6yzTwZTrlcXT
3d0w4jjuht4EgnTzFko43piEOYwuit0/KjJuf9D8nkVCxLR1eTbio1r2iYNI7Tg5
vSSGv1AASSet6EknoOnHX8x44rtRApiucnzSSRB5s9uTQr0RaaGlUT3BjTwsnkpC
25dKLDQHtWbySxXQ/2xNtJr16oYXYkkkCYSl0HTwelSoUO0gM9dz2Lunx9KkisnN
38wtLniBCUkoasiKfgTTL3Xmt8SjJbQcJBe6W9tRW4yMHhFBxGxIj1HOwR14bHA0
pZn52SnewHBqZ3hWtft/GpuA9W9cMWyZj+F7MifnYyqgcZrvur++d1/Nw7+IBuqa
tiH+56l498eoNwZynETzp76FIHnLGVaGZmPiihc1lkRQeejLQhnD0gjku9UpaF6Y
xkIksBb+gnfNHLDvex2LRCKZ1SmnXH6VUc0Nb4dyKDV7CeWWedPz9PLO9zadEfFG
t+5VG+w5eWsJAmdH2D502I9QcwNkAsj7w51BcnsxEdn117F46e/Z3S9Oeodc7Ypu
rXz0kpeWhxhBqkF7wVygL5jDQvf0azT9jTmIT21nxjdamQ/dG9HQrfYKt3ZX5AMQ
+qcWYkhpyPCk1JV4FRlQQI5cY7UkUvau6ydO0PCWDUKm4PxCCfhULcAtODT5KP7w
E4RwCJG/kQv6myVRrya3lI3GY0TpSfDhDYTtNDmLYSSXvGrYO6cQzix01Oq1LHF9
TPcZTSYBz1plwOi4Une6l2tW/C6Mi/0P4YNccR0tbFDi2qTzEH+vTCCZRGqZm7tx
+s79BslBOrye2mG9cu/+XnAdtO9PVACX/byYcVquvGwEu3VS7nN20BT60UdXgNtJ
cY6qMfJsmgVDz3+W5uooITEpANXzkFOWlNrkDYs8P6AGrJEJyXMjb3UPOkWWWZfx
JxylhSH+X6VB2mNTLRvmNN8bk9DbGx9a3CClSMN0kR2SePqvhcCfdfJghZ0UR/ZM
b475zQLh/bbRfUER05bUz2fN+mFebiTS+VaKjUqi3scd+p+0di9IPlBX7AwDzfyL
ukI5ueZD9Ge+PW/IgCwDLt88t0imIzdE9tQQXPmXsU7LoWXUCswbYqkdqWXjeHEu
BZKDzi4Kkc6w52q+vPfWUwAxMvYjCnjHzsRb1iaPFCu0eawT1n1Vdd4HzlJxbZiE
xPAGysUgBBT09ZeiLhQgiZjJnGDineB43my2Be9eiDVLfFcEf4l+0GYqWfW0GtkE
DGT8kBFQGs9ix0qXt7/31yKpRPDS16zRVEbEPeK9sNe/9+1dcBOk3nJbFuk+u0gw
G2kXMbrI0Urlr3WS3U9D7aSeOhmlfqF43xLXgD5rXLva9t+hDSaH4j/S58jhyQy7
n5Y9G62npn/LA4Vpa+Tcijk3EEjkJ5SzIbtmmsT0Q0a68W4Ck2dRDZ6OHcAmYunf
xKVt5NokJJrMnBzAiGKgrRGtsl1fgXovx0PRlGm4AXm5xuMEZF7vYwwuWG7kTE5u
KCxtkKSdK002H4Ha6Cdic48SoDHrCOxIa5PeL4+sGLJEJlu3utKZUudwUReOrUCy
UM/QGIv0r+1AxrND5NYT8SfypxxaKZ6uUkeXl6whrtlL56EBQ9ZccfxWZgT42TcA
xGt/ksjkoNm1eb8fVmrqKo6Z9wIOMsD6Ypi3SKQkAWLUAWhr5Be1XHXS0AoI188b
OfGI3ZgzZGhS2q1b042jtvZL4gn0h+0M7gvZPBaZRiy4UzBjDNzthi3W2UmwfvPB
66DlCZ6inzxbM2dfMIKIb8uaRdo9png/nLLZ00ych2d4aJsvv3xTZBlwrK8W5fbp
EZ1+1uVilLjcnPndh4PeSwxd92sGS4+EcZUptgQLowI0dKu8D1BZSYX9xy9Ofihj
ap00th9XQ7qbWiYwwBcVyQOGL8hvkldUn88W2nklRw/sRyjgfQAWCSPJGpiUsUXd
LPgMzubfmvCAY30JOsJe298Of2YiechA5bTYLNYk/bs1GjiRloNhWbTMfrlSt8+Q
l7gJQOTCwW9bsBOCfWDrerIc1WlbD9Zny4izH1+icOV0+UxgNf5pPlrxiiLzSnk6
9Z0XhtP/Ifno8vvo9TozLq3oUeMxG0WzjbcUoiJSTH3gpsQmv60vZlEZD8OX47n1
91FKP64B6VLeFBosMB37Ah2kZ6Qc6ElA5I2rVYbAiiKVS19/lb2rx7GXR8SvxNoz
nb7w1Ezj5/BMFdh3q+Hdlzo8jF77yxfbp6NLGLV+CHyNTQXCfF3M2Hn3JnNCT5OZ
VyiFij3rRmajS444Svv8PKM9qUH/Yum9pen/n7YmHdrP9ffASeeGV4Pp7x/acKQ2
qpG2nRhJojL9NW9avBRAh6zsPVtLuYnhfq3dlOe4xTQwaeIxUXH6kcsf62hhzAwi
HeLG3o6+sQu0rEOsiPCrk1BINIYYaJ/aPfdmOhp7hVP6fiWdhB9Sn0ygMBOsYMxM
JJBvAiK7crj6U/ph2VUGXnZVkQgfnd/1fu7R1JmxmTxfHrc4rJUgxuwtdanOhj/l
0l6eFdCum2o1gXnlNUxj5RH5xXZd6kOWylWl7EzXvSrmVDgUdyVTNsrqGzA/REFd
HZS6G8whe7JiO/bUWP1WTwc6hskhoH6v/umZ3f6PXdf/zTkD2ByDHcG5K3IZ3xHW
9Cb1S6zz7AfQttU425EfPtBGqU5NxKpKHQZomMIEvr4lMXyh9iOIu4n3MsItNAHU
3nmyumeTqHuAzn/bmZDq0kpAn8h07K+MsewhqZzqXEp+hdGeygDC1HCVe7b1XzW+
5O8F90hRVlPJFzGZL730cqZku5qUxaFjmgLB1ar3wNKjSR6GrO1+yj5pO4KI3HgA
YLzyXgaQtrJaIXjK2HiHGfs5l9ebaIqHp3i1tGtX46CBtOgzN1M+AVqR3BRpZ8S4
3VA9HwxUJ9yzOnsSlOhvQqE/ms9aNX761sQnsZCDUtZa2VRWZbUqJLzvSrgn8y4l
oC6HksJv64S1qVe2LD4l60/bm6PK/9QhoUsGXPxGVSD9YsIYftp8kcQwYdR1sZmp
ewAd/OG0MsDnAGMXUDTR+/++mKMGmdng1AgulBmsdM8N7PIby9zqzDJA1iuiBS1b
76w6GGAfoqj+DbTGtqEiuC6CFRVfwHSePwJJ8xBaWyKrPNWDvqwAtvE0A4RQ34WD
QdEVQpDzS6AQOt6/NbO5ROSqaQeXc5n20KnYOa1Yk2EqwyizuU3x/1qMKzY8FZtE
nQS4h8DLpzCYKMX1NuLgl3L6+SzDgLMmffe4cD4oAmEAGIrHatO44p4goD2lMYPt
QlkMdtKTsvTeKJNm+fDHdyXn1GGaqCfsrS48H6qVcRN3zEjXsXY2qjVMxXpkdyUQ
fT1HuCAmPlZ7v4tgx6TWJKzoeG72WYusnlZtYi9iPp2OLeMp/Q+GjdyZ2HlEBeND
7VrfO4oaIeS5E32LC6oZYOPyAbG1vDUdfZTH2ChZ2fOZ+n2CK9XVWPgNAOnWl13G
999s4wrYlkaAm6W+gn0ee3yMUszu8XTSqlIs+Pgc6l/yy6vZ4w26KOXC7ne5e7/K
gwwF5eSEi7loB+9ivIFfrp1a8dooCMdOLnq4b9lxCq5UgyrtwuYagWVw/RJ3iq1C
3vmC3jzATsqZu+mmEOWv4CfvXFadaW1KUPJApcRisiaoXll5oDYGMOF8uuMXPhvd
ZCCCOdaVBTZMCcf6334IUKXvaswcXQfNykEf78vniWniOOTlsc7ebHUJTAbwzabZ
ZjFtjdQVjq3z8jBT2Dju/7RoNWdbEug3hSyU3HrVTUMOKGV22kTAel6QzTG/3Cq/
EBSTN/q6WOEhP2GBwuvcXNYfUs5LF3lLujVi+/syYAzzY8kzokYq8ay0Tm02kWNG
uSte/G4YBVmJxcN9jqiqwDAiICv3JWdaYPp04plkp8BWQt+S0yknB272wPR518BP
EF2EYME0dK4b+9gJ8gHwYuhfZ+dkhWH1aW10VRvLmFg20hnI/mYdluKzflVnQ2t2
tm0LVMB+4oFeIBHUYA1JyKUf4Y+L7WMmEFFu9H1sSAhYwf+0V9VZnK43mIA1/tcQ
Y2nvCcloIJEjlls7zYbR+enrA+i4ifGnMWd8mxhzMhRMMLbXPYHAgldzpFmR0LBn
UOWGvH+IVj9JCbtRGXQYg7QDzYGJNzigD+KsK5DBXsbftBzUnSRHtWdJ8JPDLQjW
uNO9A6Nwq1YyC3N4TF5S0/3U0TR7O53CQzfbOUM1XoeBsNrzVgfWoZffXC4AAFPv
UZFwT4zmOJzVQTvzbif8RYCwRuTdbLXmVH6TcAFNd/fb/MJtFScRqT9/cQUMTRrt
ZIAc4Uoy4Y5gzK9JQSERRG8JnE0zwQEVRPKzybkbJj4b7SDZehCaTQDRNBU5GVgQ
joEFKmeYzJ0CXnzCCXKoaAei9MjWzj4wSXh4z48RE4aGoIYErAqwewpJr3644Ied
Fuzjhx+4RNPmO43IY2eahDAA7mADJoOXSTYM+3PWW8WYnqK9Iuv0nm9bwxOAcbMZ
cCC6qk6yNU3NZcjhHbYj4lVWNS+4POkjm3TZ+3ZjEUGcauJapp4YGVuwq12+1rCh
WiQP6B4SNB2pWpLKq7bUwl/Q8kfaaT+6v+BMe++TSTsqDjwMY30qI1+/ckEoE5sd
4+0TbqE8KymNMGCTMY8rC8zHEjeip3E0ImnFOItWrCH4IJ/jmzOYBLqlKTz8Ryga
/IXXhTExL7ZkzJcOzFEOT1KPoOd3bC0oMO1slwGH8Rpz6HZzztS1Qajygq5TbK/J
tfQYWJJPRG8Oir6Utp9+c059O1INu7+QgmWEJ1Vy50YNHRtZQaJuRM7aI37edT8H
SX2SzU8nVxh/nWoRIXZHggpafIcaV6SpVHdpvPkgRuQol/VtTBVCB3PqSz9NKhK4
tdzLIZD/CwZG2yw4IG9x8wLvfgIuFMDrA4cbjNkq11fYDn5QwfLm3/hyUTXaAnDc
g74CMJp3ORuuKuwhMYJUEHiGqDzrvVuScRqXM2alHDWjqA1zJre/VibVB7ZtUTy0
zdgBLW/UaHbqKCm3FY44vfyVQ2rEIZvoLIo4YtcjKhYJPYdENRWq92aWWrQK922q
mVofWdNodJB/r1QrS1rFk8cdLZD0Xnk/eZtCke9TyPF2JUsX6iCdTMLuwETEbEqh
19ZmwYlcPhJMe9EY1Hv5nIA9aQIXsITEHg68f8IsGnkj9B/A9+J6O9EnpSbbJBJw
q+QZduVxbVf0uICUv5MmEZyyUDziliz/gPLCewav3VuQOShCjto72OKdN3eiBmRf
7uWCB/s9H7KTPanlDmVsuawogNieZXTHPgvU6O6Ln/Xvr9TuA+WSDxuM29Y8AKh2
Z6FnXS8x74t6MR/1O1HINlpSZX8aqLgsl0zoCe2e4LvaGl3vwUStazdqxWfwZihL
qf115kjyvYLC8KVvCkWLj54gUnOee5zkmJ0b0iT/8eP8Jj+czGBtdv5v2QtpSuEE
EMbL49WANCVE0XPWIpHlauaYXPSJLf3fa7XabgRFwxN3Qv6puzRwhY3/e9g4bAgj
QhF+4ut7IRNapmfQWLdCQmcyEtHCalp9NA0Xosiof7eWWbQMzCqEYpElm0xwsyv0
KhQQk68sYnS3zcH8GTYsw7bHHBZunIrf+4aiduhjSriQNhI+eisITUCEWHLWYXGw
GPtmswI3fdXfE4CuaF8AjTmHKNWnuaR9tZ/+k8AXBY7r2rkQ0j5gVUjPfnyCXEXD
gCzDZV+9jU1hymLG7OcTfpLfqFMHYk6J5qEsFXYzfWDEdDh1uoCJrg8LJB1HRrmQ
l4JRenyNegbFr4XQWvF4C7+hY0XUkE+SybarWrSLd7D8zmCeCaqmEmYR6jUULNoL
U5TBWVdRJT/JNPlp9XxvUU6+jTGyNtNy3udbQLAqhS+RLKsZOucpGMZw1w+s1AmY
LIUBMzkrK/9uFuliik8imA1KsJUDFlD1UqSuuKCJBDm33TIOlAHLx8cucOUAA4lm
Vqh8uTk+9tF9oEbVpukaVE8t9GbDAY+lhbQRRJ7It1bfrg+ugSyRezdKy/hbD570
flyK57IZCzfmkVtwzJFK04IErTcY9ZTbS0Aw9nhmrjEorlF4PeysDPjyJGLzWe5O
5RiJ3WvnubyQJcS3C1Q19a7wqUO7DmnnMEZSLm2X5BOF4ZcS1fZDEYp/ltLcGkk9
hh9sikHE/XlRqYzFIRhOccVstC7H0RweV6X0GQYp/xnVeNStS1UhT9zhTOn2sG9l
xoozb7k7cmFP1KeY3SiivXuN2I4gYf8exOWj+92Brc5r1LZmF8D4/hkaHHE9+bQL
1F15OFtFVyJRcfEoeW+i09/a7YQMEokcX/qP1nyuc5cDwlLxiOTIdPVIxZgPaxTo
pPS6kUR8/viWt3dWXKT1njPk/r60EmAn+MWemfqhQB2QCrtvahqUeC6o659cC2RI
mppZmjO6s9leUXUse/s2F46K1i9tFCH/0VPsIisPOcXO46xaWgw9UJ7+KRysZR42
IL53lxI0RooEABpOE0cfdIHxSoZLl3qThGO7K+RtV2M31arke8c9zbkZj9XB1rXP
je7yE1mr6EvcesWDk0eOf99+Ft+WUdY7DSG5HZ9LxEnI9yZLKfzUqU8y3jtPJiT6
MIeQqX0XYIt834tT5pMrS5kWg7YlcB2m1oRIChzsKdlmj3WJM4/w2w4ebZnvL/Du
Gu86rWEf8+MdSdxSrp9Lq4qRDkNGBqCAIrBHk+GrGQBAS9PyDP109FEnF+FhRA+/
OYO/8tuWGnLl8vKJRutWVvSPYuG8dGXR+B5hCxnmpFkv8JYVQswkT7RQOqKN7OWi
6rG8CPvnCmt9rop4QnUZqK28UtFkIWWc4qCCmFUCcn30F6jh8FeugkMD/c5qD+Zw
lkNaEops890p8OLIG07LKvX9YjGfXANSSoVqm0PtZ9Fl/EhvPq5mnkHgp328nsjh
R3nPe/ErjiodIfyqvW9Y7s8bSJ5SRkIjK5emhK6Bi4AAFBHF3ccOYfWjHhzM+DFL
4lVsgWnFEpaBRtiuG6PXPnvZaEWm4SpdGXtzH7lyGAeNBnC0QV6ymK+3WV60v1aN
TDuX3diOIlls6+JExq57ZZMwEr5SIxCPHCtanuioP6TI44t3j+R6OIRRbJbKFCot
dcE8kPQPvE7Yt1DgUGgB9B3Kz0VlaHwR4ZwgYqXCvhzb4bWkOsmFR+rqvSVLLGnC
fZyVczOLC3jSn5H1WbyZFY8E/7zSzrWg343Y/+TewnEaUf3WsWU3aSV2Oufc63SA
BZCmjC8jCHB99UPCFNEjUjQ48S4LEJ8BAQMp4FyLQKR0b+u5fM5wyprtkQk13y90
+MEYEnEMz3OpPqyi8OwOxWuGzd52EW0nCUW6hxp9b1j9cWWXpvVO1CoRilFK85pr
xRw7vVfsSha4qysJ/qh9sRoaMdqFA8ecASoyQhKrHN2Vb7ueabCZnH9RxdKEYvGX
v+Prb9Ars8SYCCLxAEUIAUBs3p2QqVHAPWXUmsNVlkoRKwBotQwrujX+63/sbqDw
mhbNVy3/oCvGs9XsQs6HptTwNyRwyqmd6oGwfBmbsQfWjn09rBbcj2yHUAEtfg0R
NqJYC1hrwoY1OozDcVVbZZHscmnRNx1NtTTSdQNMAKBEjtl7EDM8GFWAWyreQEEm
ebGH3hiEdkvRRRLJCQYUZfW804eqpQHf+CHLiMd5ZDjp3XtYxOw0O0mCNfMJ4b6X
raVTXxz1sZvwb0wO0M2K/s+nGFxoKWfbduwATC1hET7CpXe91zm3vukIcEfqMkBG
utTBNa29sBaUTLyiD18nkTlD+g+XwS/TR9FbLIKbD4HPaA9zxaaxf+HURcOSGQqw
DNaJ/4czoEAYfHIyUWVOGaQgPAW6p0x17cB2IDynlGxyNncJ0poAl7X8p33Qv+q6
2gIShLBDu3HKf60kMj4QeKY8ysfFOiXsfxS5YhB21C43S0lerw2nPJj4soYWRVKy
14QBZEJIce5lGv0GRyMBAgu7ZKyUn7yOakih8vrEwxsdeFVw7BlDPOOidH2AniKU
IRtb7MztTLd3nsji+M7P9jRvc9ubHiKOS1RH9m+QxKWSFqnLj0m78yuvydWODKKw
q0IJAP+6lP1vWrE48ejI3JfRRBC8aPDVCr8/I4nqCmz4e7pvuKpqpFGwMNH+sDZD
LOcST8LrnLc0L3sKLDiKpOpwlhxTXuCNsvjA2OeCtH+3PPCdYiadqQRMm6wUswuq
NXL2VqTNcURRer/hBZ9qx+C5hnPuyJr3gf1tYfDz/PB0u7UqD4C3KFXN79cZr5Yx
gKeR6QMbnpCW0xbJfKm9eobmVnUrDdphR0pmt8kP7cWH0Ael1zyOUOtwoBY2opqV
hq3n8rGdke1A+AiYTGOK/tzx5bs4yNSSUITk+AcZD7oNXpmyaOgf892NJM6wDQQL
LjsRGU18knN4RJaifUlje8iDQevqCM0bTpkGoD6ldhC4JpQq5x3EZtj1NxovFppi
V2/ua8PQ3E1XKL4tz0AyAg9MlKpqTsixbDsyHCcHiOjk8WCU3FNP1G3R6dtzUJff
Zaz3igubxanBnslFyWi2qDRyTwXRiilz4461cMRCvEA26eTTLC0opELTRjzjkqP9
fCl0AbuMhCWKSMgEIrs8taJMsTVvJZF0TRJYMc4ZBsJ1vLkdhFeQi29CUh+0CXLl
vgUr8bzKpfn8CEvkCY/AkLAXtWPt+WGDAByT3+EC5PgAmFTcVSetUAHCK6pkU0KF
uL/aTOZs56kBmKLHkKgQOzT/rFI7jN7zgeLW+iI0b3puuMuG1QiMtKYpzoJIcobV
mtezTpgB002yLISICOSYcnBqy2q4bLO3dLkJH7EJYk3gW0bK7rC69XWIfetnLGE8
4ENyK+I8y1tTpvkygjlvHgPg7Sjw/vermUo+2udsvwzKjTnoIxcyI4SER84dBYrI
V2F+DaVl5NjnNUzW7WbYC5FmPx0ucwUjWJkSexoXW91JkA1muAof6wrXz3Ue696X
jbfg1NurWSRBh8Ft/ixGhC5JvfsGwYIrcHc6w5lkeh+hmqgFdZv7zpAhm5F8+tSs
EKpiaQ6W/MwELA6q0KCZ67njlJdtlne5TuhithjZ3T4CGXhR0aYGG/3W+seS5wjV
5oEO7GHTvVgpZx89FXNrAwPVTdrGiMUmXn0PRH6IIuuoEmpVxt1/IGTUOJpUdzfN
KBAcpBx4ciTEmmsohYgC95qQYcuFsDqXyv3H3f4jQWtNckEb2PZfFZ6+Tm9Nykrg
6s4KqDNF92y/MiQerERFzPjPs8cbp5MT1r+5xmPurEd2Zu64vO5cMIb7fDhOnFSa
e6uyysRGiUjTaUfi5yK8fkFiAtJ1Y+ofX6EL27oGzF2W5uH0FBxBkMavfB+013y8
wnwGSLi5m6ZV3GwWdkPw5D6ieT5UmhaYtWVGciorTSLCmiInSPbMUbo6gtuG44bJ
zXOrit+4rfbblPaky3pa3NpENvhNLhe3A7X3e/sF+DvHIMF8trJnMxDduSI9PKl/
FI257xhBnwnGZj2mwqn/7RyOVamhyfxO8dJiPj8GZJmyCtNdQfc/DNS6aSi/XMkO
awhLri3xCItFB4MVKNxOSEUiGP3C9UnGC71RCfw7H7dSGFo2itARH56ixyVYYPPx
DWW/h6BmbGvnj3uRLS21AJfS/7TUaligNabSB93epCXr0Ht+ETpvoMcglTlo/QMR
LsmFjjmvMXrI3qQ2fxCRMu8SvFKoMuZR4xN4jX4Yopx1/PvuCqvwTrGjLXCz4e2d
OYDAct7e9WOPgwI8aHFVW9EyWpXu+OvPFtlmwGwLSvTL8JCnre1JgAQvDAnjpGMV
GK2RRd3evP3c4pIstY/hU6QWcZRz0e72vqezW6g9JkoAITxtRqYcuLLZjGrJyCvC
YXWyDD0I17lDBIIoiM0T5ljfSWvesywaibRF+8aqCtaarUGL5Kn99tOb5a+GumuF
MI1u8NW/GA3SWKHgLYTwCvMILl8iabcyG0le+Ac1wV2DEaOBBTRf04PyfTGQ8juD
HFWfedZzXX8nk6XFQxaK7cwauRSOZ25/rBYJE0P4FrPzsI9IGf22J70R0pg2Vrr2
75//ZsKKYyfxXIUsxySKQNBkwRLhyIeJBoU3UHMSTo9xVHQn4gINtw9GWd3UJspg
Ay47+9scOlWGWU5DnW/5Dqvg8x85I00tf5QrcI4U2T2HLxqOXRjZx+eHefaKE4O6
wpJ+De8jIRCZuThpT8Vz0G47EIvjvZNPeFLBfzHAqe2dRNNBDlqBlsvFe9gBThB2
3SgqteM5q1ABKo3y9siNVjbU3l3qvgHGmazY3wOIMBGPn5+BnAKHUQYoHOus7yXS
VxuEMtkrQ2fNlUFHMDiI8mf3elLu2xyNqo1yw5RhKmfjdllig3R+7ofS76IG2KYA
qwxCR44AFLifXudSAA6rbLLWwRuOiFh2sFQG9pBtMvPPFP7/ni7SXu9udNah9Ps2
AEzS3p7MZYZWNmTRD3AnHNLoXlSiSd9A8EOytnHoX368QS1DeSYsSLqpw60hcoYT
OCpqLoMdcQkGeL1Jyj5RI0AVLS7GS2QfWI7tmbRQnZlP6/bQ7wHKkfD92+NvtPzV
aurz7ltGT6CoNaVgL1yDwWB1WaJbJspm5lgaPQSAxMCfj+Lvojc8mNI2zkebGcyl
GEDPP5MHShrkj0KXZnL6QQJk0yIljfTiBbp8cvTJvi6sa4lThol5oX+hKqY/Y2C0
GprtkrvC5ePgOUgxz79nyn/7cRK3KKK4M2l988uX9AnMzousNCwizGu9aTWl/xr1
G7jyOxZRM5241gt91R1vtGOC+/nHCjMmlalDBDtQGHLlLfDjvbCwxBZoK3O0SjU+
C8v4QK5At3PbWxd0rsgyd5BM7t2zrDUZiaPd5Yv8bJXPumXE9uHV5fhdM+Ms1ZnA
uzO+R3ilTfH4m5aVML3Q+hQ8B3usJnE5+Dnz+LH6f/ARG10S8m6J5QkjOBb42Wbr
LIHBIbo/8m5UyVIWRzX8jWrhivjgpeVOzhJ4xCqT1Jmy8GApubtJzAmSyRw4JB/F
u9gejNUY4Yo21XM/ZQjrqyy/tlTWXBPA89RcfuPTXkPVldX8AcuwMlAd+uDWwZLf
LJ9vUxFtPy+icv0erpIAC06WL5pVzlyupyHB5O59Lbl1IwjkL2Arh7Yk4/UjOBYq
eTnufAPADh8KyfyKC3qhfMgvGGdavBgnGt0RRVwgqMP3A5dGr2HLMp7jyNjO5oiY
8FgBsp9ZYN+6WLcnIA9C07j5Yj8oA1q397SnKTZ4R2Dhg1h2iZpfyKFvF2xDwS2S
Yiq0V7eFDx6DRdSGVg+FPalhvUKFyJzMdLiv+xPh/uvxPA8nNfF9nhDWXDjMKfuq
ApsVkw6KevUiW3RhFCTybK5S6KoywOKc10w+BrtmqZTkZevovjq1xtloM0DJ2Q2n
06u3YdgGHeDp9GgfHpNXde5QrCWJXktPhrJ3b4EXOwcCOalvlV71ELt96D6evlJR
UUL5cHdFpZi/MnuSS9Zm8TKX/uRdqA3B2Z8K7iZfViiyOOxkSIlJXqPh/8JBuARO
YgCQ0l32ws0OOkPSLJWKIndicNf5GQI8Cz8v9r57z61A00MjrdQA28xk56t/baKO
Tfk8M7maXEgNdCXmQ2VeKlTJt6Bw4xKbnM33+hbGyGx6kg9h59ku0nsuMRgItWFf
eoNL2FOBLDv08RagKcMtmRQGDqJIS+4f1VUjgFHlocf20AIoc4NT+/M9ErJ7utp0
4UqDcba2U4pDxnwXWz5YrBUDtTKYjb6uBDhRhOufdV+d/xSUL/R5dJXjdHdUDR9z
7EZfKwR5/dLIsH3Frw0Sdg+ly26VdicxUdmP4+7WOT9wAELZWyj8OoDntK6GvQYm
qpLdny36bWUYOKOAgUm9BSxsrKAhgADcc2kXvobCxEJbVV+lx6dISSqmm/RqXNkj
6z7hkz6xneY5tz38QRRgfYmwOb8QmwT3IBpjBbRu4cms2sgahy60f0qZerwrXBdb
29JyuJ1ST7wqIyemRp7/wVBYbvOYpjV+1XVnbAhb4l/99kQZfsOrmY18mLZ30hog
WUUNoioy3+1DCcXh2HMBj9vtWkktzOxLM+1t0uA7mrmT6LHWnnNbCou57eomuwrU
s5Nj+tcLMxQBOmcIdPhi9iqyP62Y9pyF33QVctd23TDTPMjUsOHRcdd7DPgUZLOI
Y9AljK9AfOiQPSQh06W0AHKrJxZSEAIYYhjqqPVo4fYR72vGVQ8NMTZYta4cxsgv
n07n2MAdN9Enrdmy9TL9gAODtATw6xWhBP2Tz15m6FiWfVRVFBucaUrABHk3z7i5
I58cA5tCqxt7UjqxJ2oHt8r7kAp6uoy/XI9Ozro1h+EjArQ4qF2o/846ZtaTO0Gn
xxZKYzh0t5Mgb9MOSkJmOdt6rdQzWrT8FvrUG9R+vWVzqKHOE5NUlHENIUldJhYs
JAL3xsLstUkB41HiBH14h2p4W+tDasKrruCxb3G2B6UdoNoo1lQK2eNCnDCgK91x
T6/MZmEiwikPfxl259ychUBABzSqNPcdUjrsvgRbHHc732QEWBMCIfd6Qt83H0w3
GJswYgyxd0fG+2CFvvmJprzFLd+dcpmppq2PV58ktuwG/crByEqiBXNJnGuEuQSn
EwHTIh13ZPi6QTrDeoO8NY9AecR6A1RHd7xCN2V4Jmr5Fc2GJIWUxq1VfYvahVEY
zCj2AnXTO33QpcH19O7iadEXeu3f16IwcmntLQ+vpbeJQelJakgj234xe94iyNVV
LPm17x1NBG5AYmnObBpxpYalQ+6XT6nulHhLIP5vEW3QmnuVqg6H5H7gHKzws+BP
Kgmni0pNRxeEYKxfh9zzZqwq8Biq2LrA3dbi7djrzEVyLxgKSasAqR02hRMUPEzb
bJChoWi8y+jsfwE2kYcoadNNqDz+vaVTFjX6xVJi7i8b3DohMJcAIRarVN57pgXp
ld6+44voHmJMV4CAODz4zgQlSgDTzNft5cHiLlKJoDnBmoa5Sk+SOJvoRwFaIUqg
mF0SabDuLplh4ZkedL/hvJ9dYDDhELf6UVt1JN1u3FhXe8G1F1yKj0yG2UgTzdoo
yW+nMyHmD4rt8tObgZpyDUmWc29LsA41nFomU6WItvA8Yp41RUjq61y48X6uS9Sx
mBiDpDADF+xtuNXmdmniRCS7YoDBOVEYrOaSX1QNnoIo+029AY9DS2aZAG6Fpst7
CrFwpeikPUleDJ7qFfekBajZQUmLJUe5imuqt2wK/tV1lynTMHq8yyWfYS+VH4Pn
gQeaGa9TqpW1+m31M6d4m7myRE0Z5UjjtwlQBpu9K6BG+igXMEQ6M0CmcugYBqoO
YaepqDV9GWFGFMqKG4WB41ma2a4eaaXSc3WEsSwXIsUx7MkEs0TnIfA2oMvgwIgN
JoP9CXwh/nUAC+vffYw5YBzs3QVdmbGUyyEw5G3IEWEzqP+tXzqWsxTuNThwfZ+9
5Uly/E04AI/PLZ/e3vIjEfF1/X40dn+6tQ4udfOZr/CJk6120I/tun0LzLbi+Brz
xJ2QWxCcKQRnK//oO1wZsd+E1/A/J3ozjhTFeuY7T6Je0DY3cSsJ6hGA/a8m3cUU
WdsO+H0q8YB+BgDUndyfsI/MDoIZ22QC9oRpdpzQpYO5/LeLhsbGZbW0bWNKK0im
MhCnMqE18JEL5cT9/XOY7Ep3V5YuA4eG5P1YzApNp1KSLudAuDa+Nb7QW5elcTDh
QJwPY0UN2TIm0ZSLqX32C+HzRrnWuPz6oidOhVkoQLwxZUgV2kvDiNTLgxQADfX2
a7eqb3rK4LBbWAS5AQwo2qBYkOlsS+FJIBR+ldqgnfvUN1NNraPpd6z1hBaPLODr
JHs5/2ZBypXh2ogF+EQxhENNG4p9nqLv7arJY7/tMo27kVPPjbr2s9TOCby5LHbs
JF9pNN+L0dPZBHF+72zj4ZmA6rywyKjqTuUjX+Iq9MEDUS0utW1Bh2h1Q2W62M1U
QhrZvac5TGV7vyMzqFqoklVANZEO9wLwaAaN8AlEIE2XM9Db8vjotgukwJZgGYs8
2k8SyUkY5E7R2e2PGbG9zbYhn7Ooxs6gC2GYAVcvlA9EybxD1vctQIUH1aHcg/B5
hvpYLyhAGGUY5NeT5rPGtg2QyH1Xontzk9KsVjBRwQE9ProzXGNXlJ6vT6Yv0xBW
kNuwKTPyAzgaJftknh05nEvPlRJaImjH9TQcpk06gjjodY96FCJ3/eix8fwKiYLw
FiLtPSeNt1TWo5BnUCd+DEEGldJOktJSYCZNXkCWRjU1TBWdJq6TZlhLy3z/wMul
dnat0Yklpmbik6VY0MgTzUGhadRAgFPMsmNfWZnD914IqhniqEUVDLDJwaC7wGOu
6pBzZf1WAcHJKAcR+7QP+DvBKfxJMCYUM+XfNJWCoAgt8FtxQavmtIe9K4tilxON
yFSXK/2eLegsN0shKlZlnFSCtUibcQuF98o5lE4SsRoynWHHYftkngNwXlm2Nmck
O7a+E2K609RO/+2RDPSmi+u1AeOvRZOjTTvzKWMtzTtUkAljmtyEs88S/joKpaWW
BbZ8njgNFXye0jscM6/VMn92txfjt/kVj7tCaXdBxdcTA6iKhR1DbkHy3JBBrKMb
vozfkiZWcuxyXaITz1N9djj35XVMdSZBEJhegx/PrwY27WUt3Vqk/sJWACJXlSBL
Mr5jGPt+67aUkNkNpm1JpipOTAZx0mRKeP0xfX+hqGCyTZiK1ZglgqopRYVqazl4
Hs0EIHExWqvbjr4oQlbJih/cz/XegZLbtUEJuRpZ2yz6dMWR+IkL9uiaIhxGr2Aw
hmdtGcoEP/WkU5K970EU21fA85DXG40jJ3mgYCpzZLbWKek0mO1nSLWQwJ1VTTNU
u0WAzmd1pQvqcwpBPryFKVc6cQiAR1dxbi6geGPM18pwky35nOw6/wo/Sd0zVIHc
guOcq6hIUNMWQ8xEkGgTGRg14YqnzQCXsLeFFj/G7WnTPJDcyU4QYar875UpV9II
yJLjh2mlFieMtGJRk0Gje2yde5Zl0GvdFGrAdYJ5nR5zzGpeet91kyX24xlz0NF4
K8hAkKxuMeYVWdI9zOTDMEh4FrjRzYTrgP7J9Go9dnks3odiqHsJh31Dmn4i+zFn
zvC0bxsyly/I8LPbAHesPjKkx9AKO+ik/KSYQiHFciJWNalHNLoCtUlqNvq/n/vd
+g1t2Kwqc1PEAzgwH2UZj8kJen7+h5mrqVndlWE5w7BAAbZpU3bhJjEHj+4nWYji
Wo6gQ0AHrHYYs66h4/PE6v0ycjUifsxXvqe3B1iVA7UXH4dH6/nXW3uekF/yfKcj
aOcudAWKr5uEf7Xto2Grg00YzsmxXBLaTyDb+ycUUh+zRx7rcrp53DPvAD9UDQ50
vbA02eybx8w0AzXF/234tjh/KLKoaLlFSBi8mATXcCxAkV4dd+g2fVfLI1VYQoaB
7ayCQ+hCPPXTbepyKw2l1diLKK05sSa44y+Qw8kWsLulGmqlBVBEkjowkLPy0wYu
Rpa4OuyEEJ1PbjnNhcYb0xwa5SZqhlV3cctYlxt7ejgJZw/mWTParttV+ihuLWcO
dWE+5FQ7PTvWG4I3fSezBS+TiqF+bTJ2MzVmmkp8YKsAjUwGVmVdjtKJGDshLedw
ioyzUoZEef/xuaEy8Hr6Yev+GjtBW5A3N+77G75EUr0JH+ZDU4AxLylMjMudBvWM
sGL+kpoClqJbnZXa5Kl2siB5cIaFnLpJKUXXMOJSG+OC1uQCUgcFMomAm/+bV7YJ
Zyh0ZbFrUwqxI/1N4BBmRSk3Kb+fo0AAMJVBgbB9uGJiprZt0G2CJdcu0JMgBur6
w6P8q4UoR5ubhXE0VTHDpbz+jOj7+i+zQ1DI0rrp5rh2NeeQmUQq928roOtRuJmj
Tx/cAQuofA4Ynfhw6Pdxp1qxkZmZNLWNoQCxBHrY0s4lFjfmX6Kx1MvTnwOKtLer
uIKIM69kCJb8lte4HZav7KEX5HEcPs8hbqJ00qZIisGUseBCjkZtzzSfTrIXFi4a
j54MP6/Mr9IKwiOvzHVSgC2aEw77zCk78eXZfM9CrPY0EC+7ExkPER54uPYfEfBl
cIZxXZ5RT2seQTEBrYnIH9TH4vSam2Q12nGdZPVI9ns/sJ9kr0hzVXgSWqV/BOT3
5UI21/aope0LvPQCyP7v8rEch4rGFlDFmo+SXK6T97lmoOJ/0Xtk7jfIYFCtnzXe
E2XZ6LL840JgsuOIqgf0hTrsTcnituZCK1J0SfrX26+9Xa4FDwCBPM4iZuWMokHZ
1Y8cSuMzVePTc7HYjO4g8/D6CVFscF4j9tDchNROO7bY/MvNRoVsv4S0cJVQ8tzt
aGlpdJuuq5uu3Cu5xfROxwpiEqUYlO4v5RwFisE4IAmU6iGYwxLaKFOpo5IHGgpj
Buhp6A5eNHNprmEtbEpn9NOZzg9Z2pbslwi3imzxIpexVsOcNzAWY3wlDcqd4Bid
VYok5UbtoQyk7FWeH9/CaB9l0FumZ2bljyqdbvto/q8f6E4CzxHMerTMOUF5J2UQ
J+9ARkZJnHFxnwtCluts4f1cY9Hygg9m/Tt9Mvj9F7RikuA3tK2PrE+TyEWZdHTQ
mqCLVBAp7V4Q1ZhUkgzhx1it1APo+pqv1qlq2W2kLd70KZM/EwQWXtR0mqrg3lVY
4sDPEWoIEQjdqKABudV/6GjOBYTrI15PbkSZRZUPPv4avkEmKKOXCvEj1uJVm13H
TCsi7+i/V2J6UoOGg0ZAv/fWQvJXIf9VxzfcacDdZhRVrgzle1e9qgFDfQT2NdJS
rZ/PpBBHSNS7QSrizddzXQpFXiGFDwjTlLpi7lBQNuru+/06HRABjIzmdpiEyrIQ
y5NEP+lfVXGJJje6s9Whf9AQiRztXMElXOO3uL29caCul5lltRswWX6Fu57WtRLc
7XuBjHrD+v7eHjX/RqSzyfkLJ08qpsmZRQGtnSsn/OAwZRbc2hnNIbWnDchg6N+d
kqDFXgdhK14N8iGpdxyIxUVZyWUHaBfJRERu9lcE9XULUYQErkDYWmGS6fZDP23u
bSscCTO0rdq3jwkagHMaSQXRw+9mYCAtqsTJzxCMr2wwMvEr6C+G8I4WCyPtHyEL
7VLq3x5FvWvhYF69TDxUmMpGLhdXkSoeSutZ2CNbhukybqMoJOqTFuzEpzPND2Hz
HU9rn0iI1MW0hy00HWEG6WmRbrZig46Kt3KQoGeXQ8b45Cfec5KpYyqM2QaPG23F
Rn9h+JmiytCtAi1+ElifqWyRf3/yyy8fI7cai8650ceepTeZgskb9/B8kmfC5ZO+
coX7h0LXEnmdcZPQBhQQbVdhPqkmNt78CXWYBc8GySFnBdFYivIPsVaMQJ85O+WP
XHA+vC+eJjOlVpJ04HimDMVH4wmypGqAoM/MyfTRnOI4jMwo22LpboUpchcQphac
zEReCbgWDD4GF0hcaIgBo1EZ4QpqUlTIuuyIgqIgYK3le3HDqxiOAGJmjcVH8D/w
KLZ510jNlh9Aa9JNpOf6zTbhvl9GWvvBYZwXE3YltVrKbk+qDN9BsJzQvDCbvUxm
r8Vmsxg+YeRQ2cgnGR9brrQJTsEizDz3zqdUl+2+xaq/QWkSd7XQMGbQyu3nR9qY
qH9uzvmzaYkcVL+UTSIbKpGWOcl3ihPBRCnvo9ZH5deTZi3/B18ral37MqbrvwNW
x0wRq7VorFzbPPyw3vzCvH/asyPY3iSrs2aJ0rcD4eKaeR5Ke6jAThi/EHThS4W2
pXZLs6U50LIH0LsAXdgvSxzMy7nVK4VDngyWEj2JWKfHzQl8nGRnnrbp13kw61pX
7av6y+/dSvvfzDA7JclXcUPReEOgUouni1shs2mvzwKiRTUo3ZXTsOct51A6wE3e
2dD5xiogYmjOQIPswcOW8kN6vzjpvCtzmqojnP9Btdwjqx+5wPobwq2FUjSj0pb4
Yq54FFY9GA8JtkH5bPtkrS3mdlgZEqAMv5x6JN8sm3YwalQKh6jRmIDTI9NMMpzZ
PdUgVlWfFRkrHT/FMACD41Ft9KVhnufoTTgtmda0HhpNCdqhMImQKztZywZaP2sL
0uB8HdIQgfc/FM+pEq8VIWqZLnmngWuPCE+ATMaiajlLqhmJIf1cduhXNMlNpHNR
DAjhDSoaAj0faq142FRwOTiDKVk1UqbClP/VTuNxsnEPHzQ1csbY1xoaY62uzviq
1jVIGTY4FRq1cevU5tJOTJ1MnBlzJehg9CP4kAIOmFo28NzPdEop60TFoVg+oubQ
Eu55Qc/utOzdNmLKc2Q7kG1/c3mTeDIbNpyixKj309j/jkRBDPSJTlvsJJB4v0FK
6aLp8PtbU9wHXBpzM2+0z3bI/+1YhYNfLKxXflat31AaYdJqqtFUXJuhbj+JGDsv
N7lMePrWm7Ofti+IH4Q6ke0ggTdpWLp31vk3I0nGMVHJhUWB8reRhV94HciBCXx7
KRoEe8h0dGLfQkB16B4sELy/Lzr2oVoT1oqHadohVAtqpQthPJpmSGM8AUxnofg+
puLXx2pXZveJb8fJ3ABbQU6z01K0CAstzczsEvDRwPxZJppcrwgnKDHDTJwKInYw
Q1y5H6WcaBrUkFGuL4RWEOd37q/m+EouvqSr1X2ruBBGVINxM2LHMJ6LX+UBLXlU
pWz/kSgDRMtXHOsnYqhRGORXR0juwWO1KKzP6sKDEwMU17LVf/uVN5GLvdF6ghqq
Sa7z0B3PVfpCQgEPWnAujjheDud0vDaoqrm8AOIGHcbE1s4tnvtSvYb+gU0yx6ir
RD34MNQuxwn1UJZuB3f9cpTGC5fOa1v2aTMPOH+eqsAK2WXbOpmT+3/7yMopYcPv
Mr03aFEDweh6/UgkoMbVLsbCnLheKCQRr12cQBped685TWU1Q40CNAA6GgzfhJs5
6lRFpS+yjvWaYmAPNg5TDnCfOAt9udusp9WBydh/zF/CImx837KetqS4ejAsm9Vc
hD+ANPn5GWl6sERpXA52LQugbqR6e+er2EoV/HHghJU65Gdpwf8xh4qzF+JCl2C1
g8Zdr/ZEOU+OgDO0dY8qg4SKoT0h6XHtZGk3ZvkL1gQ/ZEhHBrjkjh3ZPej7XKTx
h1+UI9ge4/YM3QF8PG7Rmm7+9E1r7PGbF7/XcZoccr0JgjMYta3nSzESs/xpS7gV
7ASjEtYlzZ6DZVcXZg9EBcfG+3Ox/l6csHeuo+5cowCEbeAajk88SY8gOPTyEQvM
/xMMSKC/OhwbIoWfFioPeqWh2Jwv7VP1B6VR2Zp1rHuqmkOO1CZLkk8pXWzbalwq
LnupGpSq1pUt/H19ssJuK15YwQZ2wduJ/eD5ekILsWvebPP9T2ZipaTur8j//pk0
8CL8U80BjLHiiA2AYoZZu4Rvyvu/2OKHikpK8lBKpp3i+OQTsRDIpAAzgW802Hkw
QNXtG1GPTnNEgyEvaL/y0MVR424us2kBM6dr2mQVCOs19K5kNrPwXwJNSlDewKA1
C73Z0xBTto2OOOr9IXhBiSHew21EpSFwpZsNI/+m1qew0CAjHkmoI7XtZc0i2v0l
rHbA/kVmcQroxz+bpL3k6FYS1wtEVMI5VQWkPq2wP0DpULkpwU8SPMTeQsjhImKG
ZYYQ7TrWnvGZXiGvhO6wUsYAB8O39CVSDtkfEpPL4dMDCFpVdHbGPaB10GlDFHi7
iTuKEV+HBb0bj70nmad5AM/1qB9QR2hiagQ1U0TdspRWJ8FE+EYAQ9prKAgr8Tuh
c1M2x9+AISQfnmWgf8m0ssbCvtSv/e9NG2+3vO9RW6ZRxbzb7WhOLhgxle+ONZZS
jrzlUMeH13ffzyOAP1+MQH8CAl8yw2E1FHe8Nwz0J9+zI80GTTOQh+pvMJz/DXxc
9ep+1wNgjps/Kn6YXFTF/xjygUagtk0/HMKnFA6093ifVyejDyqHEN3BEG1tfxxd
yaC+kZ+Y4U+qoc0U0ojZwxuWa/omwB11dHH3I1GXO/rDSoAnMFBN0hGKgaNss5y9
bzngDOrT86nRPgEaQ5yUW4DfRhHIvLv+LibM+afblSJy7UJCWyOCAgbkQMadgPgA
03AkXz4HFNAbqOvdb9kv4If8vDNueEnfjCqmm8d03F47UC5fWaEUtGIak06KSxTR
oEBqoDoy0AqxhDLi8vTv5kUQEVIn7He99H0653haG/aFrvILM4/96YpczkDr50WS
XaNalEdoeWY/3Jpyn4/LRpcxGPcTpSCFoh7SAXPkDrIm4EyH+pmMNRUfWClHEWd7
AoWSpEX11x3D+8jUowhXdQqPm/pFBaFXB0hp/GQTIyamfa5i+egehgntF4e5RcUq
yoyNQh+tFIuPR0TS2Ea2CEVNl0cZyPYUAmGWs9670kzFZwZbGQhyk0U5QPzru8tU
2zDNkWp+1CdNOAsc/T7xTBV2pJMcNehO2c4AH/uQBF+tsHxmKzbvNNhbQNHw9FsR
/UIvoYb5/HAvu/4ijrM6kgKtK8zszsmfp8zMqL7ZUWPyeu+DLDLGCCmwssj3VVaX
2caStPpYvAlwGpJnZ3lFj2Xw1cj+cOl/UfwnmXydDG+p1vFHXVHd9hFRcGyJ+VXL
32n7iOGM/DtlTF6q6CSpBMNVDpIm4dGOkQd39SGZMD6YoYq+CIYCMyjLGe1+Dt6z
8xEt1zb4K39O+auDNppky3DHLD/h2pnkq7f520Q9LPCKWyNdOKl4Q0RjHR1tm3w+
ReupZz5VncG8GOfQQH7ase3+DrkhmlMLGHmMTLOvs7YJqXb5JtINdLkWZ6Nj2vqv
pf+8LgpSvZnfLMRirVJvkAa300B/aUP1HiGL+YlM7tnJrTIhi7KtG/ZY1pUF5aBE
I8qzP8F7qoTkwvjcloXDc8kHwPNPFS1mXK79V2qdoRnhW2IYJRBviGOG1CVZ3d99
Xqu/lo3y+EZs4V4+Zv5dTGD1+nkeesL3faYy+GgLhLPm17zcyJpMEPoJbgpAZZYj
044gVhh5rfYM4NWf8IjOb8jFyXhwYuIlTBt1Clmw7NtavLO+HyjvVvzGLj9rtyyo
uqGdxGNGLCLJA81dnVfyPnM28ch7CIozYixl2ThN7aWNu5dIkWau2coDpHAlmtpq
lqZT3XQRM7gdDixWXAorWPCR4Sxj6XtZsW1/dLEzbTL3mjsXVJIDoMccX55EK6Cf
g/sAZ0yzUiXhbAJQfBfF8zfuMUFaAueXc6xKO2rfzbERGgRRnU10knhPiPr3euXa
HlLJczoBfUfcgpjtsMv5DUr28Q2krCQ1tEyKA9YaKTYAkn9YuEDutUel+8jFZrBI
IXxyhbsdi/bDrn53eIl0Z1GbmJ3fnBxpyRq6eIEVBIKOVu7R9bRYWgg0wHSye4ah
7A5rWq0LW2PxpEv8vTL/7SMBFfMMO+rVGMdIgjx240jxeXPTjGSHQ++nTc2+CGnn
rhR7Jq8MyWtmEsBjb+/3pCjjTpX2+tLB6FXHjSYoXQloT7wJAncDPW6y4q+heLaU
9R0iVg/aztrXzV2RNHqrUSOTftAl/y/50cVkw85UIhglDCx3J0anm4gPmxQlfjiB
FcJKZAoDow3D5uHX8/zLmih4KiAEAvECBj4EQGLnshvuOl729wptjZ/5P83nT/6b
pkMlSfd2K3kGtuHkVANVF6Nv39+bBchkGr8BOVWKV6o5+4tlCL4LYnOJ4Hxh+4r3
4G4cc1Mq2Fsj60WOSE4uP+MlKQnyVYAFD6FnLne4/hzGFbnbsPMe/R8aFzgG9Wmt
Y1kvr5NMyM+gGqqEZQkX0mdzBkJAzDf7594kW2vr6T3fPbvFlPv0kaDc4O43N9jp
LzNn6hBZXXCN9Od3XQAeLKbg99Pit77XB1OSJsUxxv+8wvGfBnYrrIQW9gEt+KQi
NnHZG/kFqyw997e/aru+DDVedKwxe2QnxhIGMw4CumownTDLpZpezdFmKUY8hEnO
CrkTd/EfZAaDFaMzvHT0K9tRQltdIHO2wfTvDZOyPdjPSMDJt98NCWeupx4r2kOR
q7afW+0umHuG1REJbpYR+1N5K4VqE/P8qsdur/gKwqGtc3/1NntfkybcEMgD2yDT
2UIN6vMp2p20BgXolRFWUiUyAKlKY4IlCAmaUfcdfza41M33clJLq2FG3wRO2ljT
r8FluK52badAixeHHBzdn1kns4tV0z/q8luFc3lB/94LV9ZUFDkSqzzvkSvpGOd2
+61WASV4XAC80PL4S6bfoNuaEgJ7l6y/OGT+2su/3lviJ6w7sJ/o8RMt/712sPya
Kpa2ayemADeoV8mM7wA4UXwtncIi75lMTZ01IAEf3e3ZUwbvlSss+/Ixms0uRe4U
f4w2nAy8MR/bvTcNN6620BWUObdBE2xIEinPYn+3MWNs4ZYNL+T174RJo+x6bc0P
Jb1FS8+o8morCn0CDzr+gcdozNplS0Wl2ukyrmZJAAvamZ9x5X6FcxvsstMqCBV5
8BnJZ7/IcJb0DRIEcink2KYog5aUqfLqtwn3cNlEMLsVnodptvaZdkMy+UKtqgQL
mRfPUbGuRuSr0+A9cx9Cz/uVMFWorP9qV3xpqC2CCwKWCbXSFU+ynYbuo2nS4Fpt
+1VjpgcILQ+ujuMXYyfPnOst5BO/26SLYZgVUey+v/PO/xi3o49awrv5m57h+4uW
m3HL5iniTdKZWyX6FIdp+6CnIrzVNE9S4sxZtDLZ9kDrFetjjjvDQhFFSIiBsBVj
cQ5ggw1qCt15wHMiYTZOV+/9+m2B68k0en6s4ZpS75I83Zw80EZpbMydnEsGQnqd
tYhj9X291sXfjIuMk7Ch/GUnsWZLVPW1eqDAF3SyOcSFJhUsiZAEioYupDbC5xpM
KFoJc3e6zJuvrtYxCSLjBv35dCFIjmGwU6Y27TM7jhTARXzgCGqZARLchDWaYhOV
y//QH3GSVEg/ozeahTSw+v3dRglwUiuEhU2GTT2dGh2b4Mtdf83OU1rSJOuBBem8
QQMf0meNpMYkM4WJQ9mR3LXAmmKsxr/nzxmohl8ug/lb/+sQo07T6MVKuVXr6u53
srZOA1O6ufwkwuamJZWnnCq915wb6Zsn+HFbsDAen6HrHnhWQIdEhHWM9BTpef4L
hOGriNSCMJyF6e6CLoTGDJw3WqoRFkm7d8xvVyCv27W+8sx36qLRqmV/3oXDy98m
/78X73rhGMAj2nxUBoZ0t/BbnZw/OMK53Df87bs3T6LQv8yxaX23Bff1GSQu7TAk
xg4rMeZR3YIBOgZW8j0by6NzL24X1VO8gRlVpDNYiEMzeZQ2RCF0wFwhKenPvkkP
DYx3F7i5DXoBMCwXo71FGmsp+2zxleWbk0l9FMIyXwSZApXJeCvzzcNi+00W823f
mKPLbpvLZBiLlPNYwhJT7W7tZRb/+YCinagbthO6f/gFDBu2GU8+XAabjfKJ9fme
szwJ/oyN62QUkWg9DHeuPaE1pVK//xaiQbU+4akItV/wEAi2TY5r41cQSI2Hc4Cq
waQ+vCKij4rhF6rb2kERN0j1YmvXo1BgR5tQ1sdsqdS1ry+R2fBE+vSYg283gPxb
sHYWlrv05AFi8qX7OGPbSM7OCVg2/0eYzwXeOe1+ONm9MJD+Hb7Rn/9oufLHOFCV
Ltn7woKU5sotyEA+Hlr4/2aPrfcKhiuHiYbQlu0x/JOldGPHuKrt7oe1YPgcT6aI
q7ey+pjfkP//si+sKpQXYeQW6omlQBuyFuvIJYimkxgOyMHzly9wQsA6zHQ74GAW
hWJT0m1nFzwSQ4u7PT6G8ZFpGQKVvODyGaGindWuc+fV2hj4S6Fz3GbQhRiBP+s4
NI06jKbj69h7PTBxsJdZOmBf+Mp1Yy+NIWRCqs5Bh04IO/KL2Yic0/alB1iAYV0O
QGDmLkKbQ40oyw13O4WuHIEC6scyDLVVpp5SNAtbzxk/4ThSJQZOs7p+Ff7+7Wag
Yrjl961L4HzL+tm04C2x39c28iVM2sNQLteGqNn+ou+a4qWmPE+RZ0D5N1uzPpO5
wjT8tNfKFH5uhQZOlLnX1dnHXiL+KwNk3SFiRlhPZRCPNtixAURxvz2fuGRlpzsm
FMWkxW7zXIbw52xJbnv5JmzwT+vNjD16N5wklKNCIyymq0HU+T3LPVlPmCUUVTil
9SguRZhSMB2Zpyc3zmGAXr43a+gGKVE4DQG3pledXeKRa92qyYEfkqHYbqKG9zjK
7tmpp/Q0jhqEDc2CvPEqkavH90qA5Ys2nHnOFNE/eFdqzCOZ6J3BdK0A4BUi250X
bMnXRGqXQQMcPejzYUPsuOJDgDF1W6KqDTK57oEeCbvIQWxD//+DfKjSxnBjOwgU
9dft2bmjZN/cmpn+slBYZ1WGqDTKjmBGsYJ1wB3k0V3X6mFhrEC0AwN9mg3rjgX6
EiLUdUkfUg2leJdZ8aJTWmKpWAhstgj7pEUcqONUvU3YCyNy4Z4LhkLcOmkExy5B
T52cqv9pEst6WRaqZPw00LRBF2Ntz2w4vSBHp3LsJ0AjdRgudDAyyUPGMeFuCSyp
dfYXDdBT0omhNab4k3aJSax5WJ73O3X8Lgu9Q2o2FA3slvK6c2xWYuR40IokANXt
IPYjm/H8E/eyh7KwWqSwGkXytMqN5vj09A36RhnsGRXGUofnpPpYTvrGbtse/BlG
nTeXG4SQxoTxJknWtot10m3zmL9LxWRNfTJRow8mnkVUrdOfkjxNKaH2PHcDhynT
VPmX0nCafrCU+Ow4NZHo+RfSInPg2nEEgcAau0Rg3uwN8jW0TnXTkGmNfbAGd4cy
K8n0Bbj/s8XDvKePscMDQnfYu6hWieVhBqTU92ytnHLLTEGhBW+7oAYOLpu1gWIo
w52W46xRk5lGjvQ9LD6j83S/jINbGeFCqRcRqY1G2J+wjq8Z9x/iCZxSgw7KT0zP
HIxs0uL7BhCy98hBtbWG8/5LVLIoDkgSM47FoN9HVnTSrxuxvzSC8NN6jwv6J/q/
GtkkecURz5YQT1roau0XKaoF7aWOcwOVHakp/Ng0AG1h5JVcUhUobhuBWGIxjtAg
mEuZEwIMZvFr8/9rna9XcUPyoV+wK0r7hmL7hRtcwcrKVIn+qeQMF+A8KPLCKDNX
etMsEYvLFr8kYh9Oz/0H5aaCF3sabLFv4DOa0w1oPJ16SNHKuckqUfc7fGqYDCMA
15nVGnaDRj9d6HNjyNk50c7ix+eoz2GLF3WWSljtXydxfbhZ8CYOTrk0KjKMtPVl
2yML8NRsoP5nSvjZoGNb6rDFbRdbpvJmBmHjHbxUBW6RhJFy+h1JW9RFzYz069HO
fmKhOWBXNPaAGdqxUuqMlAx/yuTFuo4FFhFK/5CFqp2NqniHzmomrV3ndnMI96eY
0Jmr0g4zdc34N73Zq5rAIpEpZ5UIMSuQc1CbEnl4l5iiryKdMs0S8R2ujOI2Z1Fb
cjkIuM4/IFXg2ybao7hFWdCDj8Jr7rPGBnuduoqbuwwqQa+eS9Y1ptTtfb0q0pMA
rg30+YJbzK3AfaLVf5O7gO45AnUEfI/cHRKIvPZ83SYJr5/kyIUtQ36H8BJY4f/m
9qUmxjtrCTkp0zTz/L2kzNFyvaQEFLAu8RW0aKq/yWic61uJlQ6eDblOTeG4NfWd
Xql8TGOH5Rts8EUVoAmsI2cWVtNnypggXGSnJyNBt4c1iMnFq2TnotiNC2iFC9UN
vON5FDQDiaicwq7z/pPsvtAqpeWSsE8xXtEUtcwsFspH34KUgE9MvqyPnBeIwPdW
609OS4LZrAWHoXlv8PADBvfcqfVmABrNHP5UkNZi9PnD+cJvdIrWLzwW8yiO19oe
AtRFcHS0tYC49sZreUfTwnuxBoXMEoYBCKfX/W8UAMKQExFBxTfZLk1WbN+wmOdx
ax1qeKiQYIEhp00YNTvtwlezGpwuAplLQlFtzAb4ASD8iVI2MyM0+ReEcC+CiQhp
uuLoYxT3+tqpX2ofC+F/bvSOQYj0niMMFeo6R2bgPiE5K6hjvTIKxuMSVlVAwtld
4KCnt7aPwlp/U+rCi4hC2zq/jO/kywCl5hNXTfo6UMJ+e+4r2eeJd3VgiHhnIcvh
XDllLrNS3/MOWjIP5fs1ftlnQ/ApjxfWtesg6YDYwCV1RqGmLLmowY6yDen/Lx7c
Yab8/UF6F9UhnwQMYhxY7dTzbrbz6KHfnwowz8JXUBalgl9VT4bwOjtg1X0dyub8
+scF9JzJkP1YD6fyxCyqyHnzK3Fxi9dY23B7B0qw6ycfOjvePg9QduEuh28Oxt09
gmeoyfzeLYXWzmYCnctf1xrqOpiQh778uf1gE0fDGG9HENetz+i2UGTwFf0DP/7s
trb5/UgWI9MCEze2TLky7PkdDivAGZuwpsDc/nrt87LKNCSDD7ujJHzTEHwTtkav
5EKrapyVVHGXDcmyYIS+lI3EJ1RapsIfQW2XxOoWuzAR0xusuDe3jP5SWbFWjASc
Kah6Vze7yYHrxXGHwS5oNTCjlHkbBMzrJE1ctRwp5hh8NHsz9wc7f/X5e5/Ax94b
lI3rNc09yzkua6PdPlaUkIyqH+wG+4PbLXFR/qKnX7NaIZKzYfvYpgp3yrOOz9vL
C+GKu+7VImFOrR9MUx9Lg//LKobxypBhlWcGgQ/Zh22GVDVjjjXktNcrzwbsY6N7
3IgoNXB0BzABj7uASTl1tFelvLvvX/8WwSHgUoo/c9cgeBGsSJMtHS1UgObgSkdh
P48i8S1mPziMNRmTaNL9lPvWOcZhEHWzdjRk+JGN0s6CWL0MRtCSMnjOwaW3sn1w
wznM7Cc6oCcrmsb4MtLypXLF1/XtXkExkfv/9q9roi+SxXrhYjZzK4P6nGbTAugM
PjisPj5zuKYWQNsra4RXofUr6UJE9Opa+/n9znV/woFOweY0Plhv/0KX7sT7UoGS
9w9VT/FhffX/BFHG78lFeNZUeINQbQ1s/apeGaxVqxNONkCF4crmHxGJdRVrummI
KJCrW0GGp9M8tuGPVvlIiCEXuQFypde9MLh6y7dnpDchYFqqAqFj9EtLAL8Q8bUk
HF+FE88Hm69ChCrxEollC3w8GynfB819KhYt32zYmz326Vxm03aftl5UXFTP8lxD
L16d/Gk90nlQOiC1HYlVjB1d6sVRCSa0U7oVYI2zP88nAzXi2I6MlcWnx9abWQWc
bDWJul+kCUCLJCxIcH1YDwEGr+d/VC0uP1v/oj3+JrJJE9Tk35SNGRbWV22YBdij
rHLcq04XT1kL+5W+irWS9gJGKkB73zpx3zsLQDZpXJ+PAYC38PQxpEWqHoJ1OMC4
Duq3YWea7+2P4mOhaFJkp0VVf1zR2e5snOc9Q1dc/8Ng2CfdU321mmmDM8qpADJO
CrzsMZaTgA0+SL4jk/27ksgTmnpzVj1Hh+FzZvF21621u49JbiuTiVeG4bk+vWMW
ZljX67FeAkEQ8o3uFAimOjTEOiFsTfWLkM/iWwk84sKGuCo6u7xLkV9vCj+mnMXF
W6yu+FnOIN0szhuOQDipGxu39pUi2igGFI2wfv0OI//NLo5FWaEP0TNqP0xRpjyv
l81L1JhBnNl4bQpsZNWsmYSuosczXtYlfprjsXH+EnGVwejsEaYcbREO3TEm9DNO
nM4rph6lGrt9K0biRlozY5yf2jXDWpNLlpqJk3MzsjU/2URNyvXmoq/TX3nzC2pe
51Sb5qROWfHgOrIDX8HU+HSyiMyTvuwihYFfXHCV8ujqSbTr1csai42o2PTVWIY4
LRzv07G1CT63XAJKvH64nyJcEqlNzGHxLU2TdTjhDtr/tfnCkNZYD5cuTipKZ2sD
HzzXbl+TY1cTT6A1iDYIlvgaBKnqZWnufIkn0bx4Zo16UCF/MqaMZjrcPfKTs49s
xfbQ331ybcR8eADmZ0briMzk4yHgVJ2rBwLRr/9OJ2kt5QiPZ4T/4y/MDVebmCDP
MohiZFa4Di9YFNR7+KR2R7QJy8VtdvXU02yy1lpru++jUq8D5ToScjAKw87csJOK
ZcZRab5CydykWeFIQgGjLKvnjYIxZhiaCfqfha2D/5rbbQEheZeeFTZRHcQq8cL5
KKnj0rV7v4PDhR2a2QiIuEj7iEWikL8i6z1Qr4dJAe7D1x16LwmJ4SNrNrAz1knk
biEV7Rka+7cK/IFpkch1AYu/Zxy7TaFwVS0mn+ake4Z8I2XSNCMo/SEQhmBMi86s
vZv5kqxLr5FP3qi+zRiVjrJuopBJS11sLUrgiY0FrkMZwAzOcVMiWMEzp1t2KADj
u2uwt9lTN+X/8XGWM2wKYUMy454WlPHMkrXdnkRl654mNvWDYlEM8TteA4Y5gd19
YFdxHkM0VR7tbKp3iTibw4PR5JQKvNXWh4jmNs+FeEOeU9AjehO1gnNpkcpFXLNH
vXTFoHTU2Xj1BHeVU1ddQqqtfC2PI3183oQ6DL2ziWdYOcfPoiLRzyyYNaTd2eC/
ZSriAW1UwFem+EpQyOXgudilHfsu+VM3F7MfiExgMiGlK64hzPDnxVx7qVllnhnj
LibMhoeGqRa6qL6xskOKJtYyOPbynsID1RiSzhMY9We/6BX5XbsBGqBZ8Qda6x9a
RqMbbOg0q+H7dbhptdt41Qy1alMecCASSkXzoAfLwYUL0vGSyqvZjRFMNXU04dUa
Rc0x72HOoZW4iTcEBCkVKbR8yBpFp0XEHP3fnAYQN9G7BOBGGxOrJwl/ChO0dTS0
d0UFm2HOVW6BjhfbDDaG8pPQU3qexkKYbs1XS6kF3DvOb16uSWMKBbNxgpfV1Pa3
MvnN82WtxgwKIDPYX56HspeJDBqWmXgh2CP2GofWoBVyqBGVSXZpC8GQPBnw2yW8
ULWZNzdjQV6MWU6HVweAmBITtm/XISWN/9M3rVpuDKqZLn1lz7tYYwRzUl2OAtsa
bKZzSNOB93NguYDvyUdTv1kZOzSFjzW/70TNbinxhjurYMiXqhPRnfu1EhrVIvgn
wFLXTJKN5ZmmGzXgX7Ky1paAwpyDdGw/D2LI02afQ3rZnh/4Frr70+z0R47yGL3C
RzyJnDXOnbXHFzYslgmihdVfzE5LkjZj35Zf+V+fh+hZ3SqeyPV31I4YFjivhOWy
xLqVnCC+sRkzziqkxb3wtsxws8SGQC0dWhgWpv22blBaEvc3Bgl6rBO90pJIvpL8
/iGKVhKAvURc33bdMA4Jd7gczMKKqbldUhEI3Cl32Ug86vVDfIi17Tq9ThvUS16K
taSOmHAKRAjaM+/wVAvlOREZTYUO8TYu/irPimnzAWFqzP8PLffj1jW3ux/xAyTt
qMAO3I12J9RRCnJkUcMrk0Qol9M5f9VxA/VCWfAg2fGH4TlRIETG2bmohD4ciR5I
VEn/2siF+gNrYskdW5xRqD3pZfjvSNXrpU79YcGcXxm5+y5pQ7o6uJbMQv9R1BFt
ubJ8PQbuil7BbdpyDjQkZUMOUId03mfYOKsQrZQnHl1VWdHERLy4OE4PM8U2v9nN
6kC1VLTITgdcqJWbgjQLoG2Ln68Nl/QVd4uC1jq6EAxvEND7g7xTFDhzPzgnLecg
166MTS76DKZXHm1eYVNOkHH++asCTe4Op+UBbQMzhzYfMj6daPAKOyOw/CmQbz5l
`protect END_PROTECTED
