`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WRJ2RrD2AaeLv3nsJ7+01Br8YZD2vl/2d3r5s5YFR9ykswUwq791H9JyYzwhVcKY
/h1uZI8JryJOmB8G9nxh2g4V9FFVlmTITmYAnCWpYpyGygMlHjAg+96bqVwpRK9U
eSdXWcgL0qdX20v9QndJN3qxuAgSzVTH2cNi1/jxIHpvw8fBQNFaL63WaNZaoYu2
H3L/YJz+PIWrGEYTem19vjX20C4ouBImCKQZQ24xzkcZTUCWnVGpXbFKjez82qtY
j2xlzvDCeCJAaTKexHGv0bJ+F7XBLG3eAfkt77uWPY5vVFbntrjAjxScENv7vI2I
1fXyenpu0aXg4Jsc43Wq21dfVrh4cjm7cXpELeTTpDrfBWARdyrvmuBNPU0qSYnQ
FmKHcuAnTORx75T4Y8n19pZEzfsmxiqmW1EEehhvSdnm6xA+5myTPK1pRkMVeQWr
XZ2GSCDM6ycIDo5uhxbPugn5zfK1JO0cdrTksLOSeWUB4I8GynDuWVv5GQoa2Tz7
Jv42uR/Ksrq2jcOKFWK4n8GzItfWXnzvUMfEmVgvxYGPOwle3QWg/IezGxx0eX2R
dwsw5SKNyzLvD7xFNUvOMq9oJRdx4aZwIth2O192wT1KijKNFkOqOK9XlztYc0Vj
B4xljgOScdJw0jkgaZmRFNFu6lUUrjrIsZZfPxhOercR4AeAKBZlht1cDOkhwvDh
8PZjKjdjT8T+zbjy8Gf3J38q0mzHM6i9W/Ye1lHiMm8Xr4oQxp5fPlYa+7b853gZ
R+PStzTXSWSrA5RvNp5d1+OKN3mSWQdlAWkiZDpwLB+GmZelAbgo/B/ngcw1HJjU
9WfOHwnvJF3MRW1S1PnIE/LZ4MEecL2n7DYUX3GM9QUmj/G99Q/MDZ5kmDQJ88wQ
iEGfyHuJ4NH/4QWBxGIDjdC3+RrdZNjCDIfT86c/lDdoi/+doHwIfBcGeWJa9mHN
ZRSw2RycsYESA08pudasiOg00//UyZ9ulG1Fm4yXe3y9d16teBwZgKHc6GfEojKd
vL+m4LaH3fa/eNw9uMahLb4d8Jy5oEBTXtCAUIk6zFM77lhDXmtZWS65gcosoU3l
hfxC1RLcSW1h+cTgImB4+PyUid+i0j2S3GhspI4y2St1ZUnvP0QwD3Qq3Qj4WaYa
7UHqDn08CunTny+YLx+wQOGSFTFqpphmmK2JYiXNZzxNKT8+5+aswh3Kyr47a65z
btLgu4Ql7k6L4KiB1S7HtbsGOnG2wBikPSVrS8zcr87y4ABJZh5QVLsyv0q5Gjpv
wRBMAibHa2k0OweEDl0bhmkFHGdGB36rOAaL7H8Wu+DJDhf/WcVzQt7gM6YZf6b+
dM+zbQbxEAGBa3hxvcTNtROXyPlMNSoWAOqL/XzyU+pgsMUypU19hZsFU8ILwrfA
dibcSnjVk9AYAnP8+asSkc0X16ia57Qq2JzTTL33mZneht3xWE/Sg8PI8MeFsj94
rx/LxmPyj9T+eDpdBZFTDEn9GkvSdqrBpXU3DKpgh22HnRbR3nIyo0Bo7uwwjaYT
3tTjo7tSa3tPtNWw1t/LPq+EnLEINnnvKzsb7YJQ1Z+yntr5C1AO4Vl/NAqFV3b7
ou5Qz1Klq9TP/fIkoAGw2TKSaSRCK+eIBiK11iabNwYzoQdOrGzDuUsZOSzO0ynu
bDw3GPRzBe3nf6e+6UNV1mPwEUZBgxkOn8YB6FIPEaNuqEIMfrsgigDE17jNRMjm
Hfsbw1Gkcw6Zz+UFncXgVnOrO8Pd4ZX8ExmPrw3Sfw5T7ErSmPNYBc/3pAHouYqI
FOUFNywxnxT170o4Gzm+VM4G4JZpYzFZlcF96cQcWbc5jnH//HUfQboa9xpo9S10
debPNZfgJDfIQmE+ugM1hUJqsMyx0bVigf7DMEOcgJMb8e64khOHOpGYO+Jf4v9J
ClQl7tCQ8IjYwmc7Gsa5O2sNxJwvewpnRW9OeOzZLL8ZKx0tj3hOI7Lmnup2jADa
arDaTl50n/ybARWq2yVyTHU80TRsZlZJoFbuhA+7nXYkPEM3cTuGkxzKkdN6fjxB
/0JbDusTsiRejzRW0Sl0jbqDPbft/yjMjJkYUwvTmGQf7i61389QsRJ4ZqP6RoSE
tq9p3SappqYfA1IES6eWn4yGqWLb43gc2ckIcDO18bGaiMpQk7MPr6l3XzKkQpQZ
dpXhR87KTFoHmeVVZQgIer4EvP4nP36ylEBlIJbEyKe76C2YsNQp0GB3yqwP6Q9c
phbNlZ7ggDnC43IvehbaTmpOQUsiM37BVJFgO5nsZJd3HQ06fJbwlDaeZnGRZMfl
BVYTYTTqbzIGYqsmYUm12Zjp+HABOTaMxhAP12zHrdlLn06J2DAmCvxjclV60ISJ
4MWxp6iLlzasWGKKFwCMN52WpntSmeZi6cNycO/IVo15vDD01l8LR0M/aCLyJoHJ
6OOHzeMI4cBAKm3/m4ytn0FyOqCw2oN751ggRtlkFBGqK2gVeXcrKGb5GMWrBwK/
0ZC1JiVPQpkAQ0IT9YBBgU6b/FW9v3y+Qs88jUguw5wI/E/yF7Nx5NOUanXBleG2
+f0ACoPjFWjuy6Qzkg2hYFowWo+RW6I6xSgfGfC1jwXqPGUkVpUx3kNePhM8bTBJ
BjMWh/sXZkyHrpwkFZpayigQ2uzIwI7uq8B+cXOGRK5Vcf6ugHsu+MUYjGn8z9/J
0NTDAs6pq5o0J3RQHapSPyBYKAGUMNAUWhoHlALlglnST3NXog/Kw6Bf3kIU1NKI
PYSXEw5dkEoI99ioxSOLNFBdM7eW6r60X0I/JAtwAVXXXEAKmiyU/fLzleXq2HYY
7NHMnoVXHoUGwR+pW0pBpLRd20Qp56O/xscXMC7HYfYZB7emuY10q5Kbp7sLVjrT
OYWHzEOS4aH50F37Xv1kiOsnXAR0anMuwmIa2RRfC9ydid4rMH53Uc94j9LN+uqm
NybR8L62Gf2OKOKo4kCYGUiFKyfVZdVg48IAzAEsr5U=
`protect END_PROTECTED
