`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5v0PGzycxdnIqmgtT4QQe5Dp+9Bcc7nrgq+aA6zNIOD7r9wB9L6wK7JWFVhU0FIv
C2y3t56D7dE1Yvv8QeKYDEdf9mDBe+ixlTMS0919ICwqorMDlHhGnWybgWT5MbbV
IaDf+Z7x8Z/a+Lyt2uGrfT1R9Lyd4Z2y6/lms/nQU6HMGDpl9UX9ahkOgYWzp1yW
M77X6aYScpLJ7NWTyd13mDUXzT8+sq2G21IwbrMWMI2Cy7m38II/EKt65VSOfYZn
P8GE/Q+93zNUVXPW5BJWdlI9y34B3ZdTTxLYTX/PwuQBn/qo7hGM/2d66uYGk95w
mhq//XEKFD9qp9LisX5zrfThm0dSiUpl8UaYyy69KkVDVrumyoQVL9Vdfo6pBhFx
//R89ZNP9n0wSBvK9nw8fmR/rE8PtqMp9kwz+n0swStSWt+pYjPJG0QeQE3U6d25
7agO/m3Exb/F3qQUKyKBXQMRPBPGjGO0pk+85pHXI/Yj+Mndk58fP83pgvulS8lT
Sm3aw7DOK0xh7L63vGVD7MIDvmTn4xMJCMHZX9gmniwRTb6lyXKS0wQFmmrLyquC
ykjwFuvEJr9tbz3Ts+Yxgw3JifJVG5B4wUi8SDtMExlu/GDbkDO/729hd+037qbo
1+6j5fFhVif7Rg0yiKg3QBoXx7t2DmglWHRqOt1kosF/AYJTJEWTiJfSi10uMQV6
nqR5x+/r9Wk0MuAlYvpk5cH3ZZIkO4NH/JHVMxE2tuQ3qyOJMLKq8TuoYEQHN0mQ
dosrJ2FgLgjSt5rftcdqoK5X6OLYTnUxTdUFmiI7se7ooIcqtJl9mh3SYRmWYYk9
S0GU7DZrfjqs/VBaqOAtZK7XiGr71g7zzPsi5+S1QXnSUASu1D34FLZyc2BTFJxr
b3m701cZCSnhKKhk175HcXlwMRM1T1ujgwkGANj3f59FIhWnbpJitdLqa9f+4iwJ
p7uLYcFX7KZv8eDSswDQAA==
`protect END_PROTECTED
