`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tsiL9CajwmuS9u4bpramV71pnzJdXcehaI02oA3x4mxQtvtLAAbrxdzX+XmCywfS
ROzMrVH745iRwq40Vjl7bpvECcN2Wcg+/HwEG+RGdU+UQazXG32KzVHv/+JI244q
Lf/LibJ3j4KLZzQAaLevVD6iwaAchQSyQ3H92NY8s9e3jcbxswQONmpGoFzAVdXV
7NMsxTdHDsY27OxN9k7nVsSVKCbWWbh65Yg6TmwlS3i1C/iWDj7ZhjFpp2mzr5o+
opX4KLZbBLYJKwPJmD0CwjFfyoySp4TKRAQBONpaoLeBWgDZEm0XY27FQwLKQAQf
xyVQ1w7z5FN+G6LeCwP4XNPOWR2EVgOuKeuEbP1C+GXnjWfwk2iZesGc0RN6yds0
Aeg5IR2n10jAQXi9epx7DawJBNVl98NBbHOZibdHDKOPFejbWJZRYcJLu4l/pBrV
9Um7ji4Axc99dY6cKXC7kA==
`protect END_PROTECTED
