`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rnNN9vVT57Y06cKWAZTAQ3yyRuDqn4pOvZRtBr+Z5W42AnUAuDMJ3z+SIyMz2y6j
dTLWBstPl2f1AtALwz8pbzlj7AT9auNA3i5k2LDuS/BMOmVeUG22Iu15mZU25Tse
GYGu8XM8CWM8uWhrKmDX6zp1vPnb7K8EReeUUl42tp3KQ0ppv6LN7PABJKuqYaCf
oqz78deBwQpzzWuHZEzhlt8iHpj7YWS+jA6eUpBsmLURPuZQg5o151Xry6n08DHl
L01P/KWQiNFTm2w0+wJaLUBH5qOQkr8Dw85l9lyChAGA3PnbFvjUmvYs2MZp2z+u
R2fgYUZW4a2zE3jWhrhnYCABnxyBdA28D5mwriKVQeW4nXl0seaaaF7AIZ0mZ4ny
xT/MrGmmQVVT9VQ5A1g1Oolfbownz6m78sM496TVKN1RkE6NX5lSYKLAPDnN+CRP
jHIjbaO9JLBxrLPTSoj/NKSKxaV8bOvDFUDS1FH5Lmc/u0CxF2saX+w53GaY0E6w
Gjjbw45h1eZYM+up9ZMsAJGyANo8PN8Y3Zj0eLDaSqXF7T28Zspdhi/ylnFxZl6h
1hErrpR5TxrCGqhFgflPJTEH8Q0qwtVikD3iQ57NfKg=
`protect END_PROTECTED
