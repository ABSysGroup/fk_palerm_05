`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
28TtyqRrpdFfzfASkgZY3ua9hIK/rfcc2K2vc3zkgGkDi1OU6WiW4y+PgjY7vH44
ruUNxNssbC5LEt25Q9obuoAhS2MtxJwEj3/GzKR2r5IE7dsXIHhBN9BvE9V4g2ll
NnYGe5yInegSxlVtMLEk/yXOIYAv52Y4JptIwdXlxQYn90YeGQ4OTqtj647Ce+Pw
h9LQY+caaXGvFqJCSVgPaqoVM+Nkr2gHF1sCeQsyW5lX08ZeveXcqhvMb2OsEccZ
2NhU1EbsINTDjoPwF+rkjHbbSOD9rSHNaP9NofoSLO367NVmvjOszYqrE5P5Upgg
6rUSqjEscmP0Yi3p+OvhtU/wm4F3t9fGXhsjZ/lxAHscr3+E690+ygWY2QIMCKn9
duHj7NCxlbqUZ8uDPzq+kQ33ikLbuDxf4weQXAc6an7QIZttLSYcAacCjTRxIooa
YXkdnqWixuCYypxJcrJmCSF27IdPKJQSrESm2NfBa3OI1PuxZTk6xX3/qsTg6u7H
DFUYT/+cJUpd76aUM78/mF3EULlXUiwd7UEoJJyHdF3b9q82fpDFdy0+a1h7vtpF
4Za3dLl8FrjTvO6/y8116eoImMFFcpURGxG8QYCGVZsY2aPLKHVjiWJ2IEq++5L5
Em0CRKNwyWcoHo/PSeAAE8hZRJachm0S8u4ep37FJMQZtazA6IpOmwFhMr66LmOA
HxF8XGjyEXp1yFu9vFLvncK3qmyLv6h7m1FN/4+wIttB9jUv8FJZISF0MA+uwbpH
6rgbiwx0qPc0BsWw7Lz0KoMZcIC+SWWu02gspCzvcdByoF/49DcwpjOZqCKURF5P
Tw/uz6Za8DkN5w/6iEMSdaMzpr8POSrv4z3QL47RyBl73C6cxyQfIFRcC+dFSj3l
bBGT506pLMkzTv+20669dlWt203UZ7nZpxgp9wszJD2A+MCScx57GHoFw/GhANrg
1LVOvMqA/yyH+dwmiBhrVIDf4ZuoHbHt3+Mej7Nx8vywR4hcFjaMM4Pi3/yoWUcd
vzsVBkqiwxGwgGSbvsQ7igdHxE8eP2tPOKyYeOycSKAqHtiWhuvRq9l89xBN/KAC
CvIQsc9Dk8eGxH9Z/FP6J9NUXa2fyQRWOQlMop2RTWvqn63WGk4zhGTr5/T8iRtQ
CC8hjU99PSyBTfWlW6rHXHCImzOsq9oGKr0kxxLAER7kNHAhHE9gRark2IKHGlRm
UuUvPugeO1OPSVauY3qSZCWXHpLDgD5+XSRpxhVJhqbYHkE1jOmcCARSQL4ruRla
pn+Ne0RhOxBo/a+GmTqcQZqY3wjcQjAqwfvd0ilxZ9keryGUhNWGPOJ0PhJPOc0g
vl+t9ujd2TERVxOk90mgfNUNo9Jg0x3j++U6lpd8PpssRV4vQG4UDP8HlfiGT9PG
yjXeNNVVBWXeCs4ngy6HSk12cA6ax+R7DogsYOK1OuystpT4rva2ybvtPqvUjRUv
2i+SIlk9HQgrNyIsuiofuZGusMAGOJOQgaX8A+L7rT5jlyjL9WSDD5q5uEy3j+Y0
o8RB0TvmYReTXpSKqzBD4QvLuf2Cwr2BlBD5SwuyoqfShUQql7TidfgL617n9Ve1
x8azLMwymGj0zx6ceE6V65igokgVhXN6tlp3OBzl995m7EVkOkExvwF2yj9zlR41
vJUrAQ9tWoGc9HctrmUClOoSk0HXj59IqmQyH8V4wVO0ZX2/eO+cOX0cj/ypMSgA
pY+f0pvCvcV3/uHgoTZKzGBCxRnNV7/lFcY7+PYgpRD+v3MwJfcdX8M6EZfPevyk
3aHE7bOwk42VgGzU7RDYLu+JXdrOVH+x/qocmsXiCFn0/wwKqP70vRW+YCQqDBf5
4eMPlsQcxxTMOynPwv7Ag6IQRlNWumBQogDXLUZoCFuXUsyN/NNkxwdDbsRIL5H5
6M72CyhuRPfWCqrlaDvt0dk4gS++24I53uiiOpPdRCyy9AuDV4JxjPytd1Vh4Elt
MXWM7bXdgV33pJovMNdbRB+Ty4+btPGzEtDhi/98WZPO7J0lsZ5WxyGk3zzFcvMH
+mSIgMK5rygC+Ux4ifq9QfecNhNkO1HgNxzlx/6NimEYTdWE/OWbrU7SrPyqRzzE
tYErGAcSLKG8ltZo+1KImn9k1bPnaRR2195KVGQXMi5eatX/y4NmKLGrkw7ni4FQ
4pRFab261HLhfFaMZvKOfTsTlXlMo6xgfBihHUciIw7qsJx4AF5DV+GOf6RZDQcM
kJvEZ4FfUmM1MJLahTyPqGqGcIbhSCrsRqKzzq/vEgXBwZ9F4F9WGOw/p+tj74dc
AiWy5oyy07M93QXOIAuyx44hhtZnfPLezwu7UCnlRJQVt9i4XnV/hoTP3EZzVzpb
BMlhOl8S+iNKKhEAatvFhM9xAg3STTC/uLGlEBuYftMl1zuflsgsjtvJqeEYR+2q
m9oIqSa691DA6NgoQU4gLKi1LiSrh70lAEsbP7QxiiRJHTTg9MlWO7cBQSCX9Kaa
7oWKSV9ph5EHGGSjZWsXQSMXrUwOHgDwSn12Y+ewwqEsvK1c8k2gpCBEclyxaxtC
ejhfxxuzOFdVzaoKaLKbQVCd8MJekrX+oxDiLTpSnKI5wk5zgK6/QQLtUY/kqI3M
PsWY4lseuML3Wyl2a5blFNh3gvcBhfKFJhxv/MIcFImLgktQXuTDMk3UCo2pcnV+
Rcc/adjUCHr8sXBgx+2B8Ab+MbTqjNvHEnqKsWW8lq113TzETAofxze9m319a6jO
2PJvtf0YvLUa6okA0Tqd2nte/V+MryY7sYz3mrD45r9e6JzZjGMdIfTKk2oGbTxL
rrsKFRLaP8+9rrsIpeY5QXxjJH8H0I4QUjHiz3tR1zQ=
`protect END_PROTECTED
