`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S+1HLRz1KF2fbytYoikBi+J43kuJpHaa5OttRiC6T8zf8zz7HKZMFQlXKG8eW9hq
UXGMkvrIHBPRYPskBl7kGDmwrDjY3cnSlqlWmfcS5PCJoINWshqhUXXILrczt6XZ
3IZbZK6h+wyKmTLCL2CgvmGAk6y744zPySR2Y75aoC0Cr6jF6EvLdqbASpvqabfa
0rfGc+cchRrswNOZlQets/0diDUHima0slN+KVtzvTvQRTfEZirFdUU/cp0vK087
7BgT774cwAhsLslztyyu5I518+IkjjWcCPW+7RAg14Nw4ohpPhMixe+VsjcrqTjn
nHHwOjTWKGrUltYiqlwBiTttSnG/gzSXUbBTgm9ppRkac9aR4/NujalkbjTWjJwY
VGEn+IJmFUkhs102AKM7spieEjuSov996kxO7reCmikedUeedrPugSsxXRcPTgbq
eXdUoPC1x55iy5fze98cRqefXRbVcNbTPYmcS3XtMQqlKcps8bae80Lf9cldzfXo
o7V11sFBwhPTuJE8H1p0CUFkWeMwgu4LjG7Ips81S28=
`protect END_PROTECTED
