`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YBtLhK8c15nV9LxDfs29wFLMLlY9AFR8m1YEIeytpG0KgfnCG8/E2j2vwNF3c8t1
1hYMKLPD4diC2vJznSMw5eD416WXV7MIUc6Qbo3euOtkNvWKnnpMl/16G6cstMvX
te8QXeW69AwJLriYV/th/qeCpPvt7odnugvlbHmNu+F7mkmmk488Xc569ucQnRbs
2Cv+8gG+vHj+oOkR1/LDdQKKzlpP9yMgtqmcTieJiZEyJ+UpJuEZCWTIGRFnXMGW
5mPwxav0WrarqJFPjmQ5J4qKhl4v4CPu8UV8wGbNvazTu0RJzAZOSaM8LEbW+Hoi
za6MkffZk79bM8AZvjtip1bLTYwdaFcJs6+dymyK99L2gYin//429Egc4ETMlPqK
JwjTvEA9Un6FWAE5OzkDkXNhSZUSYWSVYMQ5iN+8J7Xm8/0Krk9MlJOlEH5gf+A8
9tXXMeBr4RsoRZpTPMF1pVAHjmXh7633e6igas7Tg7WSbTT0yvEEVqkBsH/7XO6r
MiMkHtV+CHd9wPYCmz/KpGcRAU+19nhvNRz32VAoO+tgaA4aH07N+8jHe4L6cEPp
oco1vrCbo9gYJ7zTs9BLPNN2/nlr+ZPGraOKzC7rfdmH/GZsk5Tm42dluPPX4I8+
R0rO1nEjhtnUumy4yK0WBy0J4Df4Ef27m1btRvcgcBtsQrExIQ7pl8uSpar28hWx
XkrSfbF9ffxmgusC8chaIJMLkLxpGD7rPqkzwbD6JS882B0caQrESZ18AFz5uKvl
hLll83gEs4MTlWiMeImBM+tRW8nctdLWIF5QUUcE4f7lewRi/DnwYijTgKoLxoSy
482+59HDyQd/I5ImQFzXZ5r0B2EcSkBya9nd195PLh5GFfUIagu0SV3EVwLeEH/e
mplbNC6Rtiuvh0K7ihlm/X0El0bgqdawUrQL51xijb8l51loUWo986hUu+dgz1dg
Ea0Kk7t5zEM+2Qp+disTnSoFA8a3W8cKcj0X25XO8Xl/mKjauiYJvdXtR3v93xm5
o/uDdsnJACdMpo0L7fKwz//BuQNT9Y9SAjkx7nQ3pdz8fEBru71g/rz2/nUU+36W
ZwLnRpZVxhVttCJWL9p9dxzItWE9Yro9Ma3CziBgrBlbEygFbDMj2OxgzluOMUdA
8B9w0M+xI2iSBo0TLkd5n0LiWnKsmZs1gPKaU7iG8UxiS/bBgwz+JDPmRNz0ISVt
A5o2dDTw5dtp0woxKJtBNrwZ5EVqJmnDNrK9FRd3GWH4NmdG2lq9jfAHJvoIAvVX
XmyiMlJGwpxUnDKXzvEwqMyN24rUr3Ni+G/P2/g1rUWP/cLBHDwCQphSO7tGy462
oIKk7bd5dxkn1N8AW1lUBIQfaz5xeYjzcAPquL+t5Gs0V+XqUv85URqeRy4RKc9i
PeRFqP+IEqLN/wE+XeO1lEVednD6z8HcoAsD3q40LIpA08VYbvEa6Tj2vFUfKFEO
oAJ1jk8E258z/f43Ywm8U1k09Kx3ncCCn+bFE+7FiofjTY9nWfax4SvnmSQTwOCv
bBbv9Xfc6LmOuqxVZl44shXzaCwe/Lc+Zs/Q8vc2/i3scI9mDYvrdPHyzCUvm8lB
7JalTjI8+I8EQWePgcfxY3NxmpU/IrJw0IAktNW0EBDmmvJ6bbiFCde8yMobayF4
887Q1XXqXtc67GVKDKgeX30VGwWG+Leh51pK4XwhKBZu6Bp9jBUBBvsKe/iF3OBN
HJ0mOcAIcM3ZB1gJkbN03pwL5lB1o0B2WpcL8B0aid24YMaPS51pzOWC377CvUeO
ovTBP+Gk34IZd/uRDcB9KJ2XcpU1815HsrgaYyqTNQbul+s6JwDKnu+c4R544/Q5
HLVVn0Njd3FUKtzP3OTOYXuzU+9YBtPvVlNleCJbMuTwW7sKo8XuvnVE8o37SjZq
08QvEnE8x2iTej9nR1HDYGFMdRCONOmkqyBeNg00K/QMaCOJJr7FOBYgD26IMYwT
Vvd5jyaIxvuN0TxXxPlz8eFsC+ETJvhSmipGHDc7ufDmwyowNODLUAc96oMUzabR
J5ZLYCWWAXi+NvPFX2x7SU4FeFzoo2KQbmi5ShRjUO4jWJdibeZ+JfMhkUrLjWTi
Zu8uRjpG+MCZsgSsADz3LQfnEe4NaPkjbS/V1r+N2X70ynvy5FT13frfJXSLncT9
zEElkFoea7lDK+cCxc2l9Gt5t0dOdLFQFxqEYgyjtqGCkf/H18Ff2MXIFqhYAy8V
A3UohgejyTqQXYSn443fBnOKAs8660Qj+b1gb6wOwhgWnWGnVSq7/Rx4oefJAYGw
2M/gvvDQwRZClGqd4SoEYc+yeU/WwKD5lPRGRGrEDLaaJAztRW3Mk0UoNZsGOeN2
1B/2a42Cn/MP92scWdutwJCDvUZvOIuwPgf+J8U+eZGDePuG+m0KlLyszucfLVIy
Jep/KLJUa9XNn04m7zZ0Y77fPqCTGDRN/oQJOcQwlAzqBFOpdsKta7nXN3zjoN1Q
2N54+NkutdPCgcHciY2vB5+y0mfjaXeEG2MdOdryS6nMvc0Yvyg2xsgkfEjDTic/
d25qeMIgCWHivkdpI4BW3WqYbmUWTZBEpP1T1+HD/VlsBa/hPR1EkaSLdkY/IRWA
HNiUEYTX0qjRNYLLiZ4sNrhTsFjlIA+kyQ+ooRrNDqiCsuE9P7AhCMXwXHIMLmrr
mCq5WpnJTlGuyCVdyQFNJx46OdCr+jCmJtuh8yvWStfgU5hLRlHgKhmeRnuIG+Ne
BGHjAru/yPKe2dE/QbCoN6qMKqRl9TaRzkPKkdk4x3nM3V/iILQkCWY4V8NZBhuf
EUDA8I4a8P00hl+XOxfMZPZkSaE+1J4xxugiGRyvTUmorckF9WaqiHkjCV2M8F6Z
9TWTf+XriFE5iMqvO1YIKNzSGxy89WJbyXNZszoDWh2VT81OdFeixVFOBgRi7spB
i+A1exPAvFubbr1E1Nv/bTFuOKDx/S6LWEHeBKjwncjZ251Wg1hkY52CtCwCqy16
EcVcO5bjN7MLQJ/gKwsreFoBMrcv+XmGweBKOeWRzEujHIGo9Isaylmv+Hp5pjdp
cHgJI5Ukta3B7y0Mf9pRhSCvvwYEfREQ2uJcLussB4nBqSQtnBGq137KC5FRw5cB
yEr3F4HfxiZMeUKBmt24YazE2X+FFm3KXHkIUJkELVBfbbjyITHQNKkW7qKkJ+ox
HTPadXqQxVYgUdAWQnoIfPk0/Xp8pvCzTsAvq492Q9Y/dmLu1/inHS4qvbJ75CCm
aLprvxMeTEt7xXoPQ92+1pk8iS+6mJ+nv7dFbTufeGoPkcyx34ObmjTHj3AKhnG8
JcQmRSWZC4H+rJi2q3v8M/JM8lu3RFDZZyx/Jq1iHExnrX0efAWRzGKo19GiQt6M
8GDngIlW2vs3bKRIU2YZKLAfpvCGB+6MqYSZdD3t4h3WrL/6yvoq2IxNL+20lUdn
x+3mIxeCPTPH/LhBy/bdq8j41g38Mlu7oXzt1rLlXQxlKTxVamwP6l/q9EIUa8MC
icQQvxB/BbHruIvs/1uFXHMVqYJhtBL4PhihLImrvQL/CvbA9dVzmY3MZoR7N9gy
aSvgEZbdpzVMtq4FWuweIAHui9fyfLlV9T5cFh3GjU4ZLqujY/dXzyeEtyynYKGa
lUrX6eUpoHm64rINDk13opQPIC3TxpxKqWK6rTZJ14sxSz6pDl/pKjCVhfuwyh9u
8aYU8APAXJ3eMJUuW5FednrDu52XMp+c+RpR8C2HZ+OWQr+saUIcx7RLNWEKWSja
XDC8gXqhGv9lmu24ifwLgePpCdTjTT9OrdmdoVUZcTRrt7JrqWAKwDg9A9HVUXVu
n6V40mF8Nr7BSemWOMB/+EjPoJjvrkX675/Kp1sLbFM2NtT9eoX9AMjV4Bt4HO8c
jU/QlIHBuztaeh49FiZrRllD9btO+XAbaR1vVaRAtj7pFm2UVI5vq0YtZLVJO2ZU
83bskEK65bf0cLBXG9mF640VnVhj1svZ5HBGE1UO5eP1a6T/ILkts5VzHxJlgir9
MVNF4EJSdLXf8kom5d8AFdZ8odHr4+5D9PZ/Eypb1ENG39MP65tE8pqn/lsWO0s4
CKzTnUOYX/c/q5Hb5zsS9JMacd99iUw4kCZcN+WgIejNo242Gv20z8v+kVj+sWAL
tOGMZ0Crkwfco+1+cR2WRWy/ya0rjTxWgWVKFO7RnOFnuY2DOk6ISRQBrPH6dxSd
2CSDHTwMD2tSPtMCM8dj3P+XgjBUCGzr7lX7znlKhYtLzEy0YQ3dlNL2NiWDjjy9
iYYUFJGoDkQvGRuLz+RAmzURvUWLrVm9KBVOgBfKkGZCTzLNtJhSFRQe+e/Kb3He
O5nYUuVHSZUYPdmmUI0gBUwvX28T5TUthqUmVFcCbGYom53Oh2fMBgZBYFdzwG9F
MI+VNMAWsXGJW2TRvplFIjeWkEHz16rFF5qS7+aGjY9mgnwBPWGsNl5y68fRRuEj
NlBilGuGhBkFAbZ3DAgQlgWgSx/DG8b003+DUNjZ+rd9/Zuki+raQEbTy0+6Rt3u
seIwCpVogcmsqAYObnkKbMEYYYmZjTe7AhDdL11JcgDMRIWvgH17dfMvcYe5upjN
p0FXX8NI9KIufMaH2C/XQ9z6UZyjmZ6KC2BT/JGE0RA6O1CTyustNfpiTYgxRKaV
CxO6k4inyrAgnNON7n3BExqTaFLEFODCZZoiblIo1HwsM19IAZdAQ8nt9G6KTYlp
/gzeQXx1g9tZr8s0RSaqMyXtn3kUapnrs/wMc2wa1nnNj1xuX/uiOxJqs0ENaijS
H8xkXzDMay2QeEB/RlxKaTiImKiORppkNbEmJbtdGBTNLFUyF9z15TW454CrgfdQ
9ebFQ6kYw8DAd/Bll7W3Zv29P2j0N4Xr7/h5P6j1Z1PTJSb8c2QLd4+uBY0ljej6
F4BdcL6/oJUTL1CMttM7HaYp72uEKGsVAAM+HdsbZzKoaoW+50LzG1WLcc0IFkvk
MhTPb+914+Yv9J5yChwyTlnZxfdU+9z2o7cOJP5OFp6FoMfax8lXHjRqDGXCdCKN
I41lSzVvJ83o8eESeOmCLVidW/VtBAv4EMroeB8X27LYLopaaTMUby5QdclaKKJB
hMKdPiVbyMhRuVXoxjkYRp36cGJ7gEzdjnf1dLPJ3BYGD0TXjodeEUSfrDFzfEsh
bBLYJ7iAEfzZFtb/Q5CSHVaNrauZrAurwp2VokJEwndWx072sAbSWcmqDvfPrJfy
9nb7zPwa1d3Huts/5+Id1ItWwvvTnzl/kAyaGDILnMDlvz2OI9L8HqBtZrWUoyYH
asQOpy3d6CPAB3jmjFTO2bCB9F9zUQuc6qTk1XJzZU+gL8+bot42urusk6QVxcQA
pNaW1aGIaoQGrgc/DN5d1BxgJ8TXb40UkTxUWqcBPIDLL0Vzn5Gj/lXJyHBaACCr
dglHYPOZAzisr0L4aYVGSgGzchLd8kwDvXOk4By+HaGN7jBqtfLR/JT6qT+8BDsg
vMWbaRJPxLbypgS91w92Sg5xK8+pLbS9mZ0pQwBz6OEzbQA8tHu10phlj6Ulm8Uo
+x+VjUOkji8ntoL9P1ogrI62KY/vvsDKwxh1kiyQK/3wUlUMeacPFOJHMFvTVs3M
1STf32hWALKIdjL+OB6gnBWBus78UBxEPZwcVZJsiQGAuTNbq+J9HPrCLsEG6q74
yLHMMp3vaszNpYPH+TzXLUzOfL2yhkC4qVEjTK13aGW9q7zk/O26C4+IaKIq2qJ4
7uVw1e9fb0LjvTXGpJ90h2f3Y3L5K9AovSCL6v+NdJeWc1i5tY1sdGHddCJ2CTyR
FTOH5MmPBv+y/xG5t8CBhfLr8Vzwf2QOFkostebSFO9K7Rii7v3/2KPqHG4RH0LN
kjOMETkSpbxlmhVwdbfnikbDfV1pG45IpB+So1SoSpEdP4chlVgZwOZwv6Kl+ERe
tqgHRX6dUG3JZ+cL2GHgIA4CFFdO5uexSQT+51h1eK2OCRFMILMRIZo5MS14hBfg
Un5r5SbFTPZ1xzufFjCRoeuRE1xnxUjbTQP+2BNxriWbnRG0LCsXu+agq5+CR+Bh
1dosWYm+OoLF5BYWGE54ZbkgHSLcanF8h6e84cuL6Jhp1RgMG0ro48CxNoZwuBwX
TrbvjqTujX+9HETiLPv593XQG5FA7kCYPNHzqpVl43wAtjxPosr5vl+0kxKKm3Eu
na7iVDQ2hU1vt6e7YVty7GcxzfuxnkXOML0+DLPpXhfMyNXyiNFXVqhCh8aSy+xz
uynbrotbXe5wyhba//Obb9SoRzdfJ7+RNwOkUrFfUbg6U0v/SvAXvYNjP/tmet/J
U916LU5RGB7UH1GwoDzJ7aD9RV3gJAakERpTGh8vELlqU8Us/dCHE2y1tXNywNgL
eO2njTpMBkwI7H2hgWObBF7USJAdzjf+CxnX/oGaBshY6JC+jqbhO+21V45Utvrn
hzkkUXtV+11+JhMzBlcQcGYjtUdPTCFuNBjkh9BxqtUvV55d7ntkh+Yl8/V7sdtU
Kti4bW/A23Z+hAa3ApUkEmcF/uuvVRRAlbvvesRb4h+YJURj1P9SmEGd/bp5TDsT
wwBJvliudjpy0OdbCJ0lmF/ocSdBsqoLoC16xyQl+s5X7/EXHONrW+Lx2zCkRRn3
n8K41N1acD3PX8dBhfYf4gJnnyJTbnFcfeip3VZf5mKLaXLNwuCgpX2FNsxXNw8J
3Ei/SVYJtiy+iuKtakSSVnTtoR+wHda8LR29BYqQcFdpDuqwUPGPTFudAd2F8Ure
Zm+Fxn/0FOOYnbMJ9mt5kyNpwuP+iPxftjQxIiRTPLvEQeXr6MiIumWABTD4Lt58
bUxcNdDuHe0ArdOREKvPIu2CEkCq/Wa2OHrcxoId0olwL+cxIi6HOp82t7AP+pM1
X2c9JbVoOX2mSYp4l2LM3ENCk9j+9RiZ3kO4luBEiwbaLEeLhax2jQ4HgTDzkJmW
Ed7hys37+LB9VDpDdtZJL/0lL4niAlQB5gpIGpG0CzS8QN13nEcNcbU/8y817IAH
TPW6d8fyUlEu+ntxTTx2XpBlxZtSY45hcIjmgz7mqeaEqDJDsNhbmG/iJ9PCcFta
mtOaSTM3jX8IfMrtldXblSg0RwpJl8Xl7Q2KGlEiE6LR0soVf7Iq0+OKC8NIva5y
lt4JGZ+d+y1KmcBzPGRmAUiE2iV7AOkB6tVYbv3cpd8V/7fr1MqRw8DiG8+dgqdA
nQ46WCV6Is4pywORf4gcT4C3oRD7nPqvk3DpCrmXrfDKWbdvSxp+795mGXPIvQv/
HY/Sj/+x8HfcIG0lRZ2mWV95NknS/hovTMgxov42UYelRFpyOY8PFc3IV0Z/8D5d
YW2pa1bO0YJDJs3mHCujeLkGzZYw63Zhsx8O3Z4fF2Ku/rMJbeM9mEGsJredZ0mx
wvwngpg4VWRQ26oUeLpOzYJKsAtQNk5J/BVqnli4Zuk/FrQ7Xsqh5AUPAp26sCzc
LvvvK4g3UxM1W2U7p9mQuPVS4uTn9+Qt7x/KA1nGAUfeqx/vduG+wPVmJwH0gSfK
BrnBjNJiDFzA+YGie/1k8TCu7lcRfAOWkXUZ9F6btdyicGLcZDm8cUubffa2FMAB
V4tH2vrSROUtbS85/yW7J1JgvnVjPmn+JntMm1kgzpxK2lIYKhskf9R5/ffdTkTo
PJbo4N4x6bb50BfM1Ta5T2BXq5Zbe6D2fyZYKGG+WJUF8HombOHoywNZ9R2OsnlT
gGNC4sKKDrYERQDQMT4UgZaybyX6QEsVHWinjuxHy4zQCJW4i2LzYsO+maW/fNfx
67fXe5S2yQgdBAeJutjsxeD/eMombzGiPj2cHNfLwVKdaAXPMJYTs5S0kJuuL91s
RO1z8/2bCaA7o5tKyv+YkhBaDc0mS2x5E5jphT5gZo27y1WIHRi96TlZi7XbhcE9
QI8a/B5CPLuRqCx/3Z83PCa1tNO0J139Z+1f6gCKjGIE6uBQaoYk/ExOzOiqNRzc
gDI7k91mn1PTXMTfMhhfy7QABa8iEzBQFdn6bLBO05Y9jvaEO4t93vdv04lNqy+g
v1bC/+4uvqgx0sr6Bn3il66SbUUWRKt407smApnJLR1NI6RS+FtD0ZYMkCZSMCGO
5DPrKy+1ytKl5EWmtE25ZOtde9gjcKrXkDYHLna8Cjigp0U8mj3wGG3z2UtSK9w1
rem85FT1QVmC+mswAnnjb4jpyH9SouxRHuU0X8bXuTVIGaYSeNKJwc4ley7dqLBV
p0zLwHYVI88foSCbVusl3gM8zkFgW5lpaDZmKU1MqfmmiUtLzj/ryC2E25tuSTeN
H6+YAZkl4tVnsbMtvDyAluu9ce5zj9qd4Rt8l9v09gkPNNsuvcgwAhlE/ctg8924
+5pgjqDxh37Suvt291UBXDH1XeuIKr/mutbJDfPEy2cMAi8CgXjSlMHLQKjXcP88
/afUfj2vh8LMCXF0G5C/GMLnbrwhXzKTrnXxcZ/YQeCdA0pEBA12MjfbfsQz/Zfa
KRM1iWEbkE6cPfBWv94RbufAcRxXHVs5lotDcDWS2sndl/dtV823Q0kJ/VaES/uF
PlRxFQUmToHKgq1lYpUr/Cg8nK7XnRqueD0sCfr1DTHverbbyLrzmSPcQvCi2bkp
jk1hbSF/XzatwE4SGSoiLI7q1Ecc3JqfdFvavy9RPQxP1fllH1pnGh0kDJNxPS0f
ZHSJGKDxZm30ZRu6ZILKSA96fLCMXtZ50QnK+7zcJZkpHTzrVrQ5WpgKdwJcMK7A
fnlyOD5nHRGUkbhve9eQPENFWuHi/ASH7DmC8mOJtB85UoKs3UjGMy12JJWpskTV
YbpiJ2/nKABp5xwbnXaxXdSIl0TTOGMJnzD9CG94ONp9hN2s36TW2yVt+HW9W3ZC
AkFOfSDxVjeqo0ZE6VFahxEcPO7sWrAridR6/VSChQD+4h1htJL5IcjOrW51EheJ
AGmny7uKE4Sceds9do9VO0nLU3yrbi7NgHTtSza2+M2vQ1Nlly5B98yDWAHZMvlD
c+YHVs9Olwz7crF47n4jHVBzvtmRmn1CTVjdG4+RaFvQQgLm/R0nSvfzm3q7kdLO
A9jOYxltPMRxb70Qr269elr+XMGCdgJa64FdPlrPXuUgnLpMJ93tRvBdfvSfzim/
PSGKQ27VkVF6xsywbFIr6UGkDvGUDPHeOVyUDAegQhz84MRWxC7lJeqbhxU93tjJ
+T5boVYlfhY3kxLvPQwB3i8XZmHA7iG0CfsO3l0MxzM4nHJS4PCmdrFHPHA78wXn
SMOsvErrWIUGGlMch3UzfIfnG9vqbm9wTCF/ySirr8wVo8okYMvjD8rLe1JXmEuE
AtWFwq+9e1GvwbK0+BTr+hw/aOH15V2VM1lzcuf0yxhALJjmvbcVSXNQH68YPNYJ
nzkaaYr++mcsr6Gc8bTn1GFFpe8WDPnM9jYFXeYqDvTf8mTcmAffBeLa96Jke7yM
lFbCZ8FYOMscmTFW43a3X4jixsQbKhz155mdNYwSGerBZzsPrfPkeCoysdfRqOqA
PYLMDaIo55Vk64nCp91zi4gxTZ9qjgoyf8Zjqj0Ie+xuBjF3UN9kL360Ax0jrjVS
vvcHC606k9pFhDMO7SpgKyst3q+h4C7gf4rq7wgZj6b0gQyh/++YnkAQzjnMSrtt
plRMcsEBkmg0bWuxnrLkYhcaJeRN7/Id7nBCrp1hIYePIXXEFwxFXRCTypEq3sfL
jCMfGAyqBp6tPTG8811S0PaRhWqxv4fUUo65rpwbD4av72z4cEHGMmzVc/h4Hov+
yc+z5wMXsiEkzU4urZB5Nxy0Y2seZIJxQNiG/FAbM68DZRNBGhfxa8Qg7YY7b8f9
syuu0GM/c5YJD1pH28rp5AtJdF8HwuhLOdeN3VvFFqLph/ZyRs70gYqL0otLF153
RAF2WJrz4loScTpOeRAqYtf+Icss1Vb8N+uibBHgKwcDP7nlVsF4rZulQuCh+1hk
bpvDGC4RS9w6BZYnYgjWxfJnrb8D+2S5uTYwH8E+kB5djo6OgE5jAGtXug3ugwVV
u2ne3LoR9EzcLx7wKQkE7qMZoz/ncEwUGThqcGkmhnnw8ZwthGYlLNCKnkwfKsDB
qQ5Vzrf01BV2oHIVHiYL6Kaf+/TiiLxcx4fT0RKcyz5CyAwMuFk1L+tb4YSoqqEC
Ol295OMKS7ZosqAZzEJiTdqnLREMmfAueiPAlI77QKDK626UIDYyGZE+c81x9OUa
ZxCNKHuFY8g9aj5hDHoEcbeGy4MHkdLFuXqEB7107+0NXNCOdOgGKOXxC+FLgi50
uV0UoETes1cireLhUk23YiP0W9Ay0vi+i80KAwGIAhyywximR5dUKbsvEmLv+RhA
ZcQ5w4YRJzCEi0oTFc7eHOxkno9yLbfI5o2yLkv4Ek1Tne8UD9Bso4Qx0ktwaZWZ
/NdhScZjlb6woELSuTrl/vcBTXOIBX1w/ZhTrkyH2BJJ9AQDIu64xL6onxv9kjxq
JluUmD+rMgM2YYCN/fCrGxbnOBz82Gnbp9cMpXN4hrh+csLSFaq8Re2k413jlfqW
akjFSCEOjlWvV5Q4GzlN8YHhwcddWN+RiUThBWwbN0nwEIEC1GSDbqptPIpxGlyv
YR4Bt71+R8iyReRxHqd12HZZvTGHZusY3fL6JlrM2qo0xK1QcgVOnq3kF4SzeBC8
FDeqY59VhS5+KunyPgIWXIElo8va993KJLbcsYsLf5OM17fyonNmEUsEM3LzEK13
Yxv5G1IbOO/W6ZbfxXiQeKCg3Ay/WpTnZdMQ0Mk3P7fq4fTGtZfIlYgGOtaY8aAI
L+FNCcujPErkWBi2nbnPHK30aAhyP/lrABsZh496rabhyQOW32X0fugmAbBxn0ZQ
i508Wlxp/tECPBj1nGTk1S9fkby6XkRW/NdSDvr73Wpho0HW/C0/+GHetXN5+AkN
fgWVSNPixdycyOnfV8nakmkk2Qz/xcCOLd1iL8kilDrXheug8Gq9OV+O0YPUvCGz
dhczotR8N+GbqaGLJBK2+HpPPRjwqHJ23xl1H5tHvSjR+xzgtrozc88KWAnLSz2h
5TxZTqxSUE5b3MQKwNB3WBDK4r+3OzfnH2DtGj+nweztnfvJkTHHScwjSDvfgrjL
yZa22JdCMYZIzqyXovUvB96QndxJTsCmvybCON8JtIZfAY74kc6YTB6Cl5RCAEu6
LQzIS/BLvDbaljD0Zf1F2x5QkdAs6XnHKRMdr0CVbD0O+IRiosEl1tZZv+j5AXuG
79/1lYDNDntyXnuDMwAFO3Rg9ROGr2lOzCGuIYm3S5t4Gsj79WvL0Ds2q1BmOq0U
K3PM1ePjPfpfiWZuLBs+/v6yCbrkk9mv7DhEyu46XSwDmxGoQ3ePk6zT7lLSX1Ki
joCMqb4iedHoR1rQ1q5hRFRwta+/6swAckj2Z6jqOAap5WG5Q3SbSwGp/9ybWSFo
Zsimnp+XvNIyAyQGUJ02hkoNOXge+5losbeh3vz61Wb2KSHK+E4anHG1ZOJOpebC
gsfhfbfJfpZFLOp3tIWwCpgJuWgjw1uxyDxCm28YjhKtV1gBVPu0zUVm2AM4wdu8
rookpAUYk+I0Kg7r1UFONwLbZhxtN+lWk6wNehMzHq0st5Lf9Di2uTKry7fJ6+mV
1dCPHdrGe5ZRAxTyCA7nKjlYhxGebTqwRsLwvFXuHtLwtlsILYNRx9h3MgIU+gZ/
AFnNClIUCrB5KG94X+kZU11MWe7sHHCxyhJ9TdndlvOxMJS4ciHvPCWlLCKzp/c8
VBFm3gTC2RI4NDgGFUhKbEwGPk8cbRJQmuLwQlKheIkG9hHU+TdNimyISmrd1GxK
xivnJaiSWGHyupPaUH2vOzIZCbFRPGaNBtkYsmLRIFEXOoZXAAzVkj4+ec5e3JK9
uhGXheOkUjN8/hK4v9wEJqmmoVonelob30oBpCwL5qPHRBqL9JLN8vm8DyxaRj2y
HL7ruhqSvNvqsyRODLl1MUcHTG551A3yuE2CVSscN1MbShRrE2S5bunElnYjp761
NOWX7CLYf8kF4thUnyelAO4KgvUac3V9B5o+Y3UNY7fqZfV/KcjLYWAWmMiDPy6e
cYIdkV5MOuHERu6Np2H/K+/W2SlR+pwhlVj6y0w2Xer0ZXqr+4TmlSQpbxHNu0LF
WueX1zhHzXUo6TUvhV85Ez7VE5T8PgpegXSRxUxiqo0Czcf2yqOu+Lxp6QBTc1mw
btvPV0YtcA0YA0fSZK36yE2x08xKutnxQ/IAI+V3M42orDK7dcpOJgftrlu0i3iM
8c3brrBOoI+PV25x5B6s/vufo5RG/3BbJCf3pq5YBKdBOMdTqq1vKbkuXxVBFi14
ctEILD2BdPhWU9g0Dn5QXfJCZf0YgPtvusv6WOt/so4V67TbFhLN59ZKzzgoUGjY
D+iygxjJgKBKrpD0dCSCt0Hg7erhIm4gkSn+vsy6UoHHOGIp4reSnrExdE29ujE/
hMSMBewTgleWvKtCZo8Bg+lkyAmwWsV1xNLYe8vd5aOr7LWy0pIA3ixMQ9Lb7eJh
hWanI9NBoiKJ1ksgnzOEf3MSP9hevB4o2b+owNaLLq6be0ae1s8MHR1joSwj2Gcb
R2g9rDmpyd/+biLntVFvlSrWSWIOt1zE0dVYlwUk7OTns4O3xjG+4jsWazOTZ5nL
PuiO6SUuFIa8CXOoVaytMYrGKpr0aM58c7TS83LnUH2K0kWnbZO1wx29GvBTxJ8Q
PxhR8RFj5SOVZekKdj7MSmlpG7YtjoBQDcI8aIB+0OdQ7NSi/T7kfWOxHKxOE70H
6UiVTD1EveOTwoPWjlee//z5mxwbI10WAsmbUAbL23qYK5Tihyeyh7vJ5OrCj//4
84cEMI7kQEgQA9nluSS0PQhnQe/loHpx9r+icc5m0+fxDA6MNOdvHcMvPd+FoDYd
FTFG/yQ7QLzJQg3HedOVk4JZ6Dn70Wcy+5daIe7Lmg/HEb1QsTCSx9m4rX65vHzn
xTSxRQqFrW5QFKBbPxqLHg+ZGM3QF2HNEgnZYwdC72byoKlC1/w/OmgrMVFY7pGH
MRqXGFNsq1x5N4+SfMD3u22VJjoNqXr3iXFSCSIfQzec+vCZI+ATIbHq7v0JRspP
UgejJwVDOxHRQnuNi6EnnU+TxTkhQ+wOnFT/hPBeR43I7h4m4tw19/kNYiaKkvb/
P30jUT+pB2ZorR/SIKZb+S4COCVpAiEogaW4bWh/bQ1+OvruqqCVaePo4RrLiHoB
dhBWtlK7SemcrPHY5KJzmeqDvTRDRiaVu+7I/YfLITfpEaOz9UR54Aw9G/ojHwyN
qU4gvwEJ0xyHpFxcCCEyDSORMcD/LUbpqABsBxJ88/WXrOcp03hhiiQomgVcaZq2
45wB7J8mRf4ICB0TRyujInJgdDXiUGckW7D+B91edbPNTyWa+rcnkKkfiSHIQDE6
bGVdwAieI5SrssoflmEMOHOuTB+EJW9BMcB8ewNX+FrIWdAKTeO/KO2vec8fwUt1
GaMs3B5Tuw0q8WBZ2t8bU7N/iuuFd9O+nHndK0eepW5rSeC9iU+yyumQAIUKbQHo
KABqosaa9p5AtDkTk4d4N1ZRUzkdohua7T/PhKQe1IN7ju1YQYSRS2ahoAqSM6zu
O95Veq8i/NmzUlgQhhcKQe3XxW5rs1JXDXj+07xQ5ac5/ugoR+MN/HZOZmhgcCNH
zFxU0Q1yXSz0yCMEHhjE7uM+u6364iaOOv2+YPg6xc1ZAiexeZTZXaBpl3NTGHFJ
9ZF7FLnh5P1mQeYhWsnFIyTXaYBLCNVU1H3MaVJoyR6EQHC+1s4SRjWUYQN3dM7u
EDcq8FP2003oyKbIERu57sR54pT5frFCaG03hkVk93ocPCz2rlTnjxL7t6o8P2RM
/JyWQbLDE3YD/HBNwBEV0pQYqgX7XxEIn7HPDcZOU0WXIgbeMyvVSxz4jbJf/n9w
qvus+N4UPv6ttfwkMJLIgCBYPgvyDZebf7Fo4O9zKGHoYa/QET18leAfoKh1xncH
UciCUWABhtlF42WjvOCeNElKc4MKsie+0ykXKb91+jjfEjx+t8rcqQcXWu3WeCXl
lhK5OfcvmvhHqzA/cO262hpJ8CQvTfxzScirtL5Yz4nX2UTRO3sOxwUrontP5QjN
B+phtXH1f0LxMKWrPToz6WqASDRtagR8VdDWBDSw8s9+F2eh0Wu5zfVQkDz/J4DM
JirXP23b9SWOSBNTOzecB6NQ/p0448JQ3WffQB4Egf3WRbRusapVYOtG3Qs+NXlR
CHWuW3r8AAr/sCcDd5+ZAs2rYwVhLgSAqbbCFj9XreR9J0xgXxUKBhzzGPetehNO
ImPldg9hBXd2RLsi3OzTuW77T1CNrlU1eK3JJpycAsDoJV0gTJeKsyAvqA53Bw6j
D+0d60k5UgPO8vH4yqMjB9VyDxToNsuWh5egKSnnudUY4UeSbSsSOm9Q7NFwxlj9
tcmS11HUZwrzFKV89GQLJIy2ek0yIO75nCjNjg7Jkgp3L8KmxZ4Yu8QbWeNnnXYf
5CKmmp0N5R46J3EQUykLsG5f/pSCw2KL3dqvRn+bo9gaPDC9EVfiHLpWGloHtKA+
eXCscQcZs9vpt18hLfJYGaE+UBArKk38bl0yeHgPhwbTHmQnG4mRyJiInrLF6Kiy
jJbHdX12Aa90yMQuJ0q+tXYI4SThCizGzFv5Q+11OUNyDAPzq/6BrJCir6zqjS7u
bHpvnTCUSkGslwyzvHCsoqK/cK9Y8hbM/A2T+YtbDNoQzcdW3fMdGY7qEs4HHADM
SVU6KPJ17kqdR/kVw33Q4a+TCmJwbrdBSPUEN1igP5gFIUheyztUqftB0O5yoptZ
P+FKSnJecMKiJSctH7AzEbS+7n7IFqfzPlLm8l0fQ6nCRVarDEzacKByVrdjRznS
fDqRPobi2SnngRg4Zxxf1Y171VUmo1yv78MF/lCsSQEHPtjVXYLjsRD99zeRdu4m
y6AmvkWV5fh4c+wvbKH3/4UFmbbq3+dqpQvVFHgSnKNlsdTCOzist0TZvxYbK4hE
zoKM0FJytI9i5TAjh0K+OMtfc+PpTSxGMqEum65F0w8MDz7C17M/NVwftvkNaFhw
e4cEQMDqtmGfuaqGwmr7WU+/Lhjlbn1Ivwl5pqXZPyJfZD8y0mQgks5SrYbuzRpP
dEFL6noh52CPGWYrB+Ci4OI6OuWaqkUB2BqMbYZu/Lbvv307OppIpFTcONK3hsij
rKS96SCK4gXEPmyOGUrGuJ7m9jbRdsfmlsHXYq9Q++kx9+nYqipm77+YaiBnEmM+
YgFdLupd+RAQp+08YjGiIWI/rrtTiKAkSPG7lf2QU87n0ezc7sJt4/XkVZJmrK6/
11R0KApBIT7y9hqWt4KMMxSd+pgmLNqKq8/0Fx4EdQYBjaLfploWtIYNjFnOSc5+
ukOCEDcSQm1F3lsY0HBAskDMjGHlbWgmw8OHQw59stH5l6BVEacqJll0CFXdRZHe
PNrBw6bXZGXovtFqI08NN3tCUfygNnu/eKjb/JDOp/uBYwzkV6HLupCZjvL1hKeV
It//GkRboM0dE8uV+wDgcjLGBbI+98xCyHL++kAGMvMM4dfFFu2NTlx6N3RxwlUs
nQ4HXb7ZesoMlC2mhM2UTOtc424tgpXO21Em7NsS4gvu3GGDmuikB7BNKBqNhD2l
JA5GSVKNxoaBRSShfE1BCbq5fc1Mgx6O7BatGjyKppSGTieDP7cZ51aYMGtyab2U
AGFDiCbxhWOiQ74MqGDGOk1WZeIiGAxul8XIsi/Wn5sIyPPX0FUkJHfvkxS9pfZE
w23b8+HR8X+9ivUckuY7ve3VCeo4m2vLdps6vxN07oF8xgv51jYNfhfMWh3i6xly
w5g55tBXtcgogpcAHbbrBEDJnNkyfcKaFHaj+pAFGe5JPoW4Yt4vdB0KCsjDBUFi
Y4z4Vm30hASs1+KlzJDO5MUeU5WYea/iqpDbR5D9Ustlg+T+Wv1Kr6ruaqFG+k/Y
u9QkOwL4KWzNUP1UkCk1KO3MezFoQG0DGVpgl7VuKn/7zkb6XjXojgNRkcwUdwaA
iqhLceFifrWKoEKdrpTtH8S3hDLzhi79hLRJGwz5X5pnaT1LfzffmuUmBlBRyphp
f7GrfoXYwUtQyfTNkc5BNXzgGYXIlcvNXM2P2I41kqt+iJ5N7A7A+tbozMMltUtS
qGFbH4L/EejRcb/LEgeewl7Ntd12A6qJX656dAPfAFvxt/zHh9JIyRmRfo7Pry8p
OZYaX27NBWmjhYKDsn59KipA29NJtPuJVbgmY36e7lUDVBRN8FSJbSrUmrTtTqTN
U4k1h6U6VUA/M2LKpPvcCUuV5SEHvq+h5CmN6++7zGXPxw/6e46vHam6J1kr0uDJ
AorKswNYTvWZo5pzmnT6Px3QtuRG9hAGBvOq09HxZk+kmOHPuHvQVtJ5lGQVuQeZ
/Lv6ywhQluitkbvFytFvF99OA11c5jHnhOOu5TPc2ytGZwLUPGuo9ZEdAN6Sl0Oi
julsV+1IqXVOt3PB+owUHKQ/XQcwRQkpfPzhGFKX0489CF/dxlwMhUmTborMbcp1
GXoaaLY1v6n434RorjtB4uMw5FrsubBYcO33hYPXlXMv8315GW3jux0S8Ez280eR
fSfneA0t5XGMPZAMUpUnv212Cu7rfWDgpjH2vJ2IaWF2osxssxxDID+CPCuFLFly
Nt7PY87Isq4n1dpvJhcU+LZcZ00OpgZ0Cjf2dnq+zBqQqZeGLkdoviB3i9tD2IPp
EIp+YHOnnUSCpA/e4nyknQUaCyVbIm2mJi9HyYOLc+Mp7HjC1pt6kYX23xHJO0ZF
7K+OYvK0kLYzwJyMAa4Sd2Lrd2J1U2Qp/FG4MT+I9AtNb12txMtYj3SKUWRdnZ+F
BECZr8PxtFF3669Hyyvx0ah5xRFxr6u22coY3QaLL5VZM4HqVpalgDZ4hgpvV1YY
qcbM0beuTbgKFHyYnNVFuw7pSZ0EgPDVazAs2J1nnZ37jT/Jj2o/pKTkF7CnORc6
RbNa3pTP5j6R4dDjPE5W8VMM5HjliDRpdFeck+pMcctnT4efvVbUWCTqFbNk0Zfq
1751f/bsHja8uaNvrqHapMhE/hlIN3wqoVSre71OEkMolvIExy9NQvDPLGva6R8k
AaGjwbdK8MZz5zG/vxvAokWRiMAZzglgSZC4zJZwOVm7cZGi/BNVH0yGv183QHmc
0LeGZPmCEMY5XAqueXUWULtSu98Yhk5XjhsiFncnvZy01YzbL6gQzbqb9/uXMIeR
T8FZvtzH/dzY/fLzO4XT/u+wmX+/xLbKFwIo0TRz73HPHJlx5X4PXh6m8UAFR+jh
juINjboNW/HEHfGRSFw7CydMy7ua16uFb3bGMmcMEpA1EcN7RLqQnMRjwtZvH6Qf
j2F+8j0rz8y2XgBDNTyS1V7LcAVZty47jK/3ZCoujtnYO7HSeXlGYvwrA4ktTci8
C9SrL/xh1UzMHIEcUzLX8zttbtsJJSE/ryu5Lw1Oguu9cf+ELJjFtNCktnwBDd8o
uG7HtM9ojOiTL2nGIhL7DMAnkz9m6tTcvNqQtaFpAoYGKLJ+NMm8zcJmOAA3JtYa
L8YndjH1T/PVyE4fD9TCLi7puQpZcFbSGosHkZlrH1sLbldPAXWuOb6CZlxUskL0
E8zNmPuX3Zu8CTPlcmuwLe+nByQv6nqKgPpwOpXttTNmfLI8XwAiR5MXpj1ZHVDW
sRSlzn3te8NRQ7TrjdRBMGMm0IPteGily+rVjLGSApIifBcc7BoqP34sFmMj4q76
Vzh8We6juZR8jKbqmSlyLWxZ6dnwL3Dj/qry1Aid6ylyuFMA0H5jW1CkMtPc6iDZ
STnOPdUaO4LCYyV2icj8bu9zl5bhH4bYw1hpNrH5MMR40f+2ADignz1G1Icd82d6
0neryJwmxAhUxInLwfqsaZEzhDAuCV4qokvJrUc2DmjJVbPGvLiqbRpMpUWQdqxU
MaVG3Fn1tvloNh4IyT8zV6O6630kbwlfh1J9SkXB9x18SjehkUFdRfuM/03cEyan
Fy6Scexj1YSFiNaDnvM6rDP/K/RbGuKgjpmfrgOrkjwkhLdPGuNxrPU/vMYjF56c
VXXh+FbWcGGV0wemJKR/bmqTciecnUabzQT/6/iK5QYH15ExwpY1haICNt7+xg4E
3it265EVDZAHMmPnCzrcjxES356D68l4VcjTKVgeUcPlmTxN4kIPcyBmo/SBJki9
/sk4o7Gcv2vW4c/njVi57aJikVrtcwdQ9a/T396ncjKnj6k73xyb/7X11MpMTvPG
5zraia0qm/zbz8GDrdy1elnOcqOnTHJrowS0PMFtSdGDaLPoC9bPalCYuOeZxEjN
B9hX1VfsM8xBg1tL2ohgW5tnD+XX6R0PKZveHesXITcsLCvV8Q97n3IjGAJkMdul
gd1MrptbOLx2weIzCOmR2SUkufDVAkKMPuj+jU+m3Kn1hL/xFzL9kW7Hc5hg9/7r
XhJiRWBAiA2HQyzA9Jbqavp+KkLblqsZgrH0qnRhuT/x8NaxWcTATuBLs0jdTWyq
NfBQ6GG8NRLUJlKD8TwL7a2Q1kxZHwoJo9f0QfbYg/KOzH/z5ucu6981wwzWIwlx
z2PWH0iqFA8WTghbcnfgQFcaw3lo2hW6DhncgbmLi9dKJ0ZipOiUeB2Iea8vkmfa
xcaqClm+c+tM7uXop0bx+/+RlgxJ+3dOGmP7L68BzrMUzFWOXglNw/Ew0rcavbEi
ppnWH2NY5awSITo+ij8kL59qb54kgDxs1kkPddI+0hYDXQ8CqCJSZrxAWRTSQG6+
8cvDoR9WREBIq+J7R9ec5kjc8B8R6wbMCIJujryCLY21BJ/EDBGbHlPW50KJZyx8
SXl6oTEZnp7T6rGyWGMOxPlJgKlca+vt+JqU3iFE2mB5dwXNPkg/iQZvmjkc1QtX
Mo2H7do/RYwlVw9VhLfzVTeHHz4SzjvV0MbKHWWdQWlGXph7hjcELRBRosX7Rd/e
ragNGZYTqvdBYeuHGj/7S4glJeAnpUs0XK2+5dV7ZWNV52hU2QNuKsNtZ150rkaH
DpRAlvKCk3cDAMiS623cYZU+ZHmbLRwp9d1JJ9IGdE4op0ZTwAeTKf11FXY0YEJn
9goMeDQ7WQedCMF1bsN0Eg7Xn53ecVHvO3xcZaLSKS1EtRBGRs9Ys5LDZU0NpYIx
cM0hvnyGCdS2TMj3/3tKv6jQwAAHBVQA3M9y2Pb+l3SNcZCv4gxIYrLpZ1toNYkZ
zjZ9nU3NLJRmMy4RKtGSVng9olXUlbIsVT7bl4oYTaONxBAGf1FMh/l4V6HHN03u
wutBCrvdo72TcUGNRRQn7NO/o5TSQS6Fw6FQ773XyexwUaaXr3+ZLTp4qv0oQ8Dj
fjoRdPiTWNy8M6oSAZGb6Cq5g0tuytPh+Ad3suvgR0P/g2ah+CprbZEl0QuWw3dj
7fSTiBiPqGWdlFvF3kmakp2UG8DF1KRz2AqJUCXy4CBw1nZI8LUNcQx6pireRyvo
aoxua4S+unk2Hffbp15LymTcGzzPt7nDucC/fmqmp3D7KYdHEelRhwUJ6TBbrP+K
Oe0cuTw409BCjQsZoTYrhmREb+B/P79cSIHQsrFWKZF08I4tkXF0CCc+k8NywKbI
BbYBLLtdULHGk1XLfwfSTVY+rNNl/nyJhWnzy4+4T7Q+3U+IPyKyD5gvUGdBKjxL
oL3Ak5hJelgr13AsGcUfzPGykrKRBxLLQO56GaE3c+nFAl5H9KModQp0eTeLpHA5
gU+afJGOe4mKBByDfio/nvuAuG/OY9JfzDpnTRsXkeYOokNHpllHbHbHG8hApqLb
xp2b1xaYYSSm6jYZS/mDQM0oOx8jiBDTmGnXdxxQl+QLw4GAhkZNPWPC88qHTkWW
0XIT/lqlcB8HMYr2bTb/oUblZjNndwG7D1+dodJLlilPtZc3yUInLTqsrVz815j0
i3MJMcLBfg2/r4QAhIzqcDq0mX5eRnM3fAO4m64XZgFtKNH28ejqlhN8HU5fsQb+
eLwtQmt4c+gODgTDdEMkAasxpEg1sNCdbR9DhLxmPT2pxN+k1KxPjD80e7pl7WMp
seevexbcC7xscFLdBh0elckKyyfOUwSJRDjvVTSPUPF5LLmilAsjo0JwXsGyCWYJ
wXxqyuC/rd+WxB5AjKdRPmI+FM1x+YNBhXUgJbVuydXxEJedAMvZY1qjW3pcbXf3
9MZyq59sslEpal3q968LEnRGpjNilQYHNACyxh8qiuZ+8g0IGvGxn5nt/r42DVb0
3RdIKzDByvat6/wfAzFGnJuvG1O442ANngZJFq4rUhS4ZDe0SvmLdViXPs9dql0f
qkhGANxOpHxfrEO8K8rnqD0CX7dEH8lAN/RtuMmDaRAFogrMrR7c95+Rky0VO6m5
FbGnPpDRsEcECC+6p+9nu1Olb8sXBoxgqo55dAIiEGEEvRAg43bnlDy+yX6EvRIL
XbewlwsRE6zj3zIySIBFujCG+mM96naOR5vXwP2xdm6Dd/sz+xR0lTsXJCLHODDz
ly2qx3x6KZL4c2usTEGGZTlLRzM2Cy8GaiZO7W675PtMLmxGVHq/WkN6Y32J8KOk
Yh/yBCniMvBzzXGjfxmbbeE2/i+0W8LAUY20v5HJN2AiMZcVSg+irWarUutl6hgx
RQzZvp9hjulBs2bBuW6oZEjN7wbSMAWR31aiwoXUuSbV4+1CZN6flpfVzxAZU3j5
x8sXQAAblAP6m1lUV9SE3VEMqdPI5IRGo3MIzDeHgLRcOl1mHanvqwgen2R3rGyG
0wNAcrCChBOFKMzS4PUB19dC5vy3z+AOz2DjxrfQnXQ1DHedQJe+kL5jvuXedMGb
ew0qtTH2s4L/CdkWcSdknHI3SfnqNPURY4giYmj7qvJHWkk1VFwCcticaUgwQ/4T
JIsIz9Y03EucpjeKK8BT7+qFEieWgc4uoOU49CnVYd9Wu5PtyDbgXeInEVRY6Fee
sREGKrgPAOA3CxKdOEDMxDZVeyLc0lyESc7EKIx9XDoKkIcCaepHsh5heyvrOX47
DHsp3uCw37VZFlulPUdOG7dtpJuEjkM1Gqr+VJMt2MSamGfgChaOk/mmijwLculB
XEL+FmzObm1mtoDBylZzvV6Pky5FEGW8WluxlysJciQVDv/k87TZuOn2ko6NmQt6
tEssFq9QzDnqYhVmRfpiIGGYQooLME6Yc75Oeuz6RMWH8/3ML2Nctfoj88hOPDiL
qXDhwpMkm32rd1F59ypRQzwKY5snILBf5yfrv4SGVw0cAKc3BsRVfZx34B7Z0+gr
sBSbZzQdu5/I8PVxJGBNF4wbAEJHdi74Dp0yM2ndiucz5YUiFxT/QCnP8n2sxbDL
6qsPv8x40EatheivO22Rk9g0QvyT3bFSiD9Ifudom9VLTeLrvYdEwvnXyhLJhLGt
xIDwqFyIuJp0G6qonJzcu3Z/fYP1p+XadyKJaTvk3dmo5JJXWzFHlx2uN8cYcaRJ
6E3KMuAZik1GwmfnBAAB/MLjwgLoDokmpN4Pwlr00Ki1kQIz/jxOUwgeu3glnVOm
ywzJ+vHMNWdJ9ewt9JHh+V11a5FGF9pM8N9Mr/QE3QdE8FbChI7yWV8oMaPHpBFw
7uKy+hn58/LJlzleSUx1fO4hRPfvn48d1BNL31Nlb4BHI2/a6YXn7TnngPMiNoHy
+0hX+DgLGUtP60deGC7M91dcw8ZkubB2q5LYdG40GV/EJoF5meflgkn7zy4PwLQ7
kJrRsK8lQqthY9LW3PMGv5/1/ngzzIepb3NJ7KkAOX4oD5Cz6L4+1G4RZmLaVPqP
kAu1TDdlkMByN5Ur5+LSDt8styL+QxNeW49pT1B/CFN4j6IXbnf4/bOtP8/iNOeI
any7rikdLoM924g9Tzi7UlL8h6dV3Q/ol6VozBJTsu9G1+xuKoq6yRPBaqSctJUY
9eRF3ysIGYgp5k7cQTz9JnPX/Z1wWtjgCg67l44XdDHWpm+WfUyVaEFjL6Db3Gz/
I26wco/CDCpbudHsDsa/tcgiicbIH4Xjr4zP64etgBD8DsudsLiYVZNVt4Dn3OYB
/dmzEQV9ESv/6KeHN7oq0V5MaJa3K7F/rnSHG/p6vNOG5c4vphnFgdNo1xg49abK
5qnSqyrDCBm3dAVQEKy2KyKQOPzGXs4zheV7vwSZgrTS/ngJ8eY3h6Ds2CFZIrwJ
L8Bse2iXRqzdbvbzgLuqY0+GgiGA48HAAKN8ylWi31eAgBwodftLqVV6EvoUl0qs
dZEYzhoZ/l/nfm2ItpTyGFv543u6Hrpb/ythFIpAidXg1YPNPnKE4oJMQoBtexhQ
+nZkdTFIl9gg8QUmUK1V31S7IBPtDdTb9ubKIB5DB0jtzrOWqVezIwZPO9jEJccu
AJ5m8Tk7tLxDpuImw7xd5mRdpseVlha6sXx6PBgdW59ZcwXQfos0fz/R2PfnlW9D
5NwkFUIOVXnmkq4jZvNieWuQqviX03Psv/Wi46eZCfgq8tLETHpu9YO7vnkRtfe/
CR1QHXgYbcinstK7CWQ035t8we8nFckLO9ZPygwCn48lADWvFU35cR7dKc9BM+Zy
FgB8Otptp74ZrocUK60RSLpp0d4+LnrFjJOi0/FOIm5i+LVRzJKqWAzbzYLMeiF/
q1/qpZsm7ufb3icaGNUyY2wufvF6MGzQWLIdEyo4IXAZeH35cMYx7g6zZlCyjvVw
hhpMQWDsN2KMU3cIpNKu7D8D1lIaj4k4nHpyUFUiIfP/+KmRhcOv3lbhJcERSmWR
rgzLexcl7TgfQIaHeWhToZi7V+ZG8Rn2x0dG6KN1d9pSiEEpoGfMRVWRhNOndtKg
TtAj/+SVmYijwbo9+LxpjqbpdXxVeZVeg69F9VS6aWDh3fkiXdXHjYrgcEuUY2Kr
2rO0AjfX4BHQ7yPgySZ4Z15r6cUlD4+XYWSEHZJtiLnD6Uv7etrqlspT6ngs2Hzk
2ppgbHDKIx8ljLn0h92Uf3ow5PkQh5pgfiiu/tSTR8/lIDpGrP3uJwyVEvs3SBKp
XpULim6Xix4MQihN25LDflXHN3Z2Lwvr1rsnuQiUxrQj+/tgbAS+D6b2S4jp24BP
9UvYQUCns1WQHSRfK9o+GNhGgnkhZYbYmaYk79ax958nAzAvbqul2GlanvccLfuU
jLM8MkzzQ5+R3CHzQybiGs8XK9dZhWKoBrQfxSNJ5AQ+VeePr6P8BtwAOrjW7eqR
A3rFsgPApRb+qmIr9lOU/ldk4/DohD6CVvimNh6R6NNpteIXsqFpzhYKQbwM1DjH
xJiIg1l0D38XTg4aydVDVyj8HgVfvE0Dy/fdLJTdk9p9bggZ6QLEiTweYo2Ijixf
diyv9MeT9hO5ZRX1B888dYM/kjX9f7q3u2z4JQ8Se1GxBNFdhqBEoW8jPO4+iLzN
x4ymRcZwss4DS/sk1AzYTI0nMAWxDs5JqYyIzEqzz6cBZ4BkopVgH2WEpf1dnEjg
owBgx8HmP4l4oPv6d+vRZjEaI1DBVXEmgvlhmuUNT2kcgteaqPFXeImtkcb7QiCB
yl9ju4DbgpmB1kkfhx/ejPrJ+ikbmggsPBVrS1wSJL0g8MHAeqmVxkiqKxn9VeGo
u0Llz3u9G4+6+Oa17dIOQ1G08hDDnRLULBD38S+dDo67Z3FScuSK0QM1LA5bypmI
qXVCEFABXNYUOz4Xflz8MSXuTIohg0B+Mz7bk9dunqMsGabHvbe2MT1kQEbLnqyW
GxkYXoiJuJuisTse+2wRikyG1rrbLBz06GcPfMuQeKBdFdby1Ol6HsBpCHgZDgSe
TLYB+ZzSNtl2mwMdtxPq2lElQQpBEMwe4XQjSNwqsNqA/bREertpLjqsLWoeDWLt
/+ZDjeJL786ipVd/9dgBEebFVOyhKZDsjWKg4KQf3m3IL4er5AxkN8FA73LBZZ0P
+BTvvqy+zRnEDZU8GRU3OpQ6Y/q86Nqebr1sW6utsNZea5jlNh7p4gjmrrXa0HBm
cpTwfdORmQ1fjtLwNN3XAmdqIdkTHtjWXhmcbTQ2Ck5lfGaBN80Yrd3L8WsmzbIG
25DxphyZ9cEd9IJfFKyYUJlYWFK5xL3TWbdXQSha1BKYCgSQq/SvnQvLDu+BmbdD
mcbLZHvdLslA5D9pHpGL/3ImxMhzXbe4juUxs8KlcEPzDyQwM7H25RDZ1Ug646pw
TQquDLgilTuh67hxqraH5Qe2POa3ry67zdhR9uH5DetdQiDHSnEVM7yoZHKerg4X
nWiTyJqzVlVKFOtRaGSXoHNldG2+f7mLHvzIun+6ceF2mbJIAf3lhxP+N1C3rPwC
hZ/OyFBNcXa/gPVXOeDXco5Yy1JTG9lJ33+dL2dzAgIJ1zFHfFJaVqT5pJcay3Cz
qDPvqSHOL4QxZlPbjAzw/aDgq2v3pW7T72+PSDeXqkRBy4Tj3FNT8ZVWjebJ7SRQ
hDB6w1oPC7V5mCXE70hi2TRa5JdCcUDycyWClF+OMdB2umOlkaV5oqBoIOT4iqUZ
dWu3yzRthulMaeDU2w4LYi/V+oYNJPXkuXZzhsvdor5BhHKzsYDCtFRQfz7JXKnz
4AMpSwKzm8Eh1SrJrmIEUHiB81zly65/EcfoSrHC2adVLCnPVW87rTaJQBi+75gM
gPfQ9Op4w5Cu+QLdTsIc9iD0L4cHYh65sz17lhsieHjL2ZozQqbz06NErz5cbPGr
KJu1/fPqM1zIuP6kh2M+iXGWtp78q7HK306txigw4mD1so82P9D8zVG0HtSCyQ3Y
Nm4yPT/sWm5wzH3DzGhEJ1aIi7jb0luJh8y3E7yoO9SnGlGsOJG6TIQ+plyZWhL4
k4/ezOS4oMcb0Y3CzRl9Y+tSMBN64mfCaaORcyevVbGrC4QcaI8gUddqYbU0adua
mGK7j9vtt5JPU1/ZJ+DDWpcy6aB436fHZOf1/UdzA0IpkOwI/Ff3sx0HJaACIGrY
GzJGY02irtfoQHm/fhPt5+uHOsCAEcpDE0PnjlIC0xoZr9Oc6nnfVOwrkgOqi4xk
yAwLrIHMcHYV/0HQLi5CLacD0oGUQi+dbRc7bnZgUy6GxioIDpPeia3nxR4w+36c
FwgEkoyNTjLvG8TPtT8+ljXK+Cs6Z1rED4E3FtgcLeGLuEGPo0ZV2soQQzA/Facw
QFNzEP7SAAQSN5+Arzq4zueX3FwLKk105omwxxkghIJmTKOjDD/niVdNyHVqNDYS
XjQ/PCA7MUwmIsHXap42xLkmZTz00WLF3hgvsB/Yqik4NjRZnlpYe1ttzPgsMm09
x5o9BMyNMwKyj5jstRDJXJgQ22C/EE1n47ZMcBtQVqDVUqIz6dpt2ZjGErxb18EZ
bhE7DyNqpoQJ0NZ2gsP/pBAVCvpxwKxTEPGRBWfMon9xHFmJCyqRXvryJJxdyeB3
wuKN8nk8g5j2kl54agkpIFGXtw3wEJp/xUcjQcDBZm0HV/ae9bz7tmgZWi90Uf1a
u2tgrbpOtYf+yiE9YZFHoUsiMOGL+oU3Tb1JH8cALOU42MB2BGQxtuUjbHbboK3u
mHK0aoZhotniWvQjAqIh56fPkunUDGX9nw1MSzdabaRPFHdU2sHVO5bEPwnp9Gse
MDRXB9tELRDCzkebjViAa7A52i6M1LHk8OcaWb9Vsln0EuhEu+KlB8iVYLEYlXcF
t7Z8VLddaIelzSTtHMdqJBWPaQeFMkW4PQEsn+sd36uVtcSEP/UBwuwFnqTPsXEe
jVqNatlStPeYfCsY+rpjuOs+s4lOb4UK3URQ2JiI0uuV7u6NfIPHlnLjIkKxRhwt
0d41QkF+bAg4DtNcIQ5xDA599EI84IMmnjyEvLSrZ7RrJ/JJJJGrBqa/63pZjv4C
rnaz4faulDcyFJhiT1SGr3tjNaem5ntUPElG3fXY6LxoFw9M/+vJdy+cvgFE7L3f
XX+6Gp0wMgJbOP1AV0+SX/QYMa7ccAZojIDxqgEI/nwjlk0iMpTvVAXruEqeECt/
kY8nQTPgGrb39EJUsFTZrNfqFXuF9OWd9/9gG9jcueIbuVTZ9CzG1JJxs42ZtEof
o6bCrf9PoFEM61PGszZZ5F+DX39wQrAG+8U07HW46xg8jn6hSh1Dz3oNm3RvPY1F
bw2XpZxG0OUsOEBTxqGnw8bnEdESa1G51NsY5hYetV2BpZKfGmQ0kRdRXKmBSgpY
MK56f4FZp8CdPKA1+00hnn/A5wsCBCQhWmKEPA8WTCApXwYpmIzhZ816uusiaekf
H77Ddyozc18a2umvUSTv0WPZzrka34H/gbW6qBav6LXgRD6CkEkUzFVkj3Cz/FbS
Ha/Fk8Xul25XD0DxM1mzCbvgVOl1k848/mlLc4xl9oleGVxZEA14OPSwW2RCccbQ
0IXGJMOLcQqNYQXLXiksJHDHUCdZ1exbERvtCLsOtcTHFpBpRDRyPmZxqr9D2rHC
6IpqjdFN2LSC+B2qxOqnKSzCBOceXy7wBSoB9nVO7ASnRUpTdpavDdG88W/d/dcT
YVeVEnrpImBYxZ++UACSX9aTj38Yzj1Rmweestx20/lqhvrqt8+HAIvTnNrgbdYE
STQc0yxM9TGjL5PsXHoPxh3iRwb1nhFgh8HhvGfC0etE+IntDUnPgYuudHLyONIv
UEVIkPpSVP/w+ovdxUvsxFDAdGEAoGg7tAPeHOJ7u8NcycdUIioKYZPmDTdVHL/Y
pGavm2537fp97nii5kUe/uiZmyArZJyVh4VGCKVEb+IKe8P4NWbvzPBduS+lrxDO
KN6swduWIL5DJ3Jlypu77iQmOxRjF/waRHIwPP9YSFTn72pL3xfRvNJZan/GZ28a
5B9MHTycJWxP5q5wHz7qBKR1KzOdt8oZYNBXa/+ewp5KfQkUcbmWM0SFTcZh2LrM
2dRrN8fRSR7f+HXOIFYE3C1CzHi8PjpnoC1uUp0GWUGPTfl4des+2DKgqa5EHkO4
JCUp423Hgg1H9zyyfAftUpfwzpL+Ghwg0DarXYu7nTZSQQMtU/HankvIeMrEGvsm
KvzYAqcD+XLfXBWJHDj3ARTTLkeXFcSwZJHNvJUlYRT32MxT5SQkcRXwdnYdCuvE
Kx1mvmeru3Y9NkaA5yMs3ih7jLRTC9q8nP9xw6wWH7NnWFvdKm7q3cLIUaMcbeqt
PFQt68VRNXoP3pC8buUF9itoqqtn2wbBoeVC39vKpRyUkPa2dNtO5pvHYE/99Yxg
c5e2FLKuigbX2ciScSWgf/rsc0V40kwQks7AfW6JrmluFxi83Zt7s0xlqA1rNKFs
W2N7L56Z54tNilxT2tw8TxBQ7Hb1ApXC2/vYf1SpTruTEMnLrXp8pBkJZjY7pmeS
1RKntiISNxkIbq/ytMKKYz3XUhHLz+XhV6pcY3LyhjK9cvxQly32sboaA21TRxED
gR6y5HvFcqnSfRDp1e+O44wfoUnS1xgSkad9diGbAJjoHw/44Lup/JX5iBPbGH1b
iLqqweH2CK0LW7m3PMD3KvbyOQc1jpVBCJlKn3aV7oP+BR9vWOsewUkHv9/ioCWc
r1Gb2C+EwQUKreK2zers7ymNljFpRbzNOQN/Ix1wTTWZrKIdtcJosiuJuBC6vQ2C
hvg2vl1TZ7QgGxHrEaPbeKEeJNoWh5OFUTMO1Fl1LDHAEeCXtjWBBJbwelJkrymc
BBhAbD228BV/oiTqHTPq7NQ1gWZu2XL/1/QxOGAm2CLdkCFsIsrG1+anh9+l86Fj
Xrz4j/n7JIFQFmb3tKQK76xzejunbTmFH5lqpkaQTT8gEet9zQCFOHcfnPU6yjSA
Wpxmq4RoZOcLd6o+CeHgZpVqoZhZa4MrdKUHYggdOclo8fEIw0T/anmtHOpXbeVr
2YbBgwwYdSoP0s8NLs8eR5k9ZHUXCj1eSfOx3MM5BfBrN/8ZkvUv/i7hsxbrt1rE
Dfa/vimZZVRYPUGnrTXBG9O2jYym0ZY9vQ2p3ryETUYnI7K6rBUwDssw0KAuRFN1
Sq19GTqbtXA5I9aY2WHOXGaOHCdG3xq9QoA9RvC0ifo7ELkOs8pT3LGo6Aab8HQq
a42+1iLmR5FipeK7Ymv7w0vfthcpE0G7KBF+IiEAKk8+O+S6wnpOVYRRhfZZIqrQ
RWUJ2kGcTHQK1WRcCwPj1sKpgoQbpT2+idzuv53HyXDYI0aHCuFPwWEUc2Saof9R
I70daTtkQPCkHnAm72FQ48ReJNVZKnpinL6gqQ4AnZyn2XbfKhG16Pa8Cc1MT38Q
I3zl4ZQkarqqkGnJJ2c5JJDKW4S5l3cJ8NR6gReZhyfggF+0cMUy/bWcfXsEe1un
tDTnT7N4h4oex/8Xf2FJ15Sr73so3iz+SVp4dljV5IO32ZG2t9tI4OCAQkMMd9xC
OOqjIIbBKrz/c9wwVrqed0LviYgizO5bLwUU2ZLev1Reqbm87RAef0ENGd0ahOJ/
p6MPYT0NcoHA2RseIoehrmahHg2Fdr0apH+O9SGFiYz56RkkvuhDQc7WrNm9+tRh
pH1dBTpoVHoUKERTR43MoU4D/0e/wGjpqqiAG31OVAeu6njf1j1cKstL2RZsbpD0
u4o6xWUE8uq0kUxmnndRh9fwa4GZevFN6yf5FYsyLN/w98GXtIWd7Wm0p8jHLwZQ
+Z9RcWqkVKx67AnB05HfUvqVcZVKL5q5eWPxPg6oSsVXnrJ3a7y4Cxjvl9SSpMEo
dWn4RNIJsW62bQPSIf4Df7AoSwLBMdm7X2gW+r9L3DU4OM5DUFZZQ12LMGnS1BMA
g78JSCzd14MrVSBWBkrx7T8qvawicshITnPjQx861rJZ53hPoBtOcWfrI4d4QU28
iQeGyzX6lD4QOoRCH/WtIMvj3ZhiEJV1ddXTxu0h/JsN3VacCKF3B/BFFXzF2kLf
cj7W5lTGa/TwkjE2zSyxRvpq1B17Kwl5spPMfmW5s1RTGzzPcKwsb3jSXxKY88b3
7NOwGlyVtv39sbVWFD68+tQkjzQ2cCcCLP6IqpEOe4fFxz+n+8IjVhQCf+NLLw01
raYsF+xlqVlqkxMaqBbWaZDbxkfRTozoyE2vCtLRqLD6w5xWDaa61oXGyIWykSDs
n96vQa4NBk35/DubOu9Iz9tvhFiC5mE5azstJMiE1X9pLpBr9Fsh0VLkh9Esgi0e
kiAFli7C3oxx+3QuMlxAJlJ4pkDupqpAX/gihMg2SmM7Bid38V9Rqson4L7zEclb
jy5UICULxV+CCMQ/TG7mQtulHDlDB7tWZf8e6UafjFOJc5fdwOE/NXsodO6fqZ5i
BMbymE4AspYbIbl1SrzlybVTXajVgkMcQY7jGpWGFHKLZDSgaTbIy3sHVN1ME1Es
uXwnDPo8aVUAoZt71WJ94P0KqjfuPGXDJjx3RK/XnojUPAmAi/rLouEQegZOVPIu
zx7c76bpNrkxbEKTn3VgyhjVay+kJwLv4ucG6ri7JPQYJD01Xaq8alLZoxuRUGD7
167iCL0EyuF3BvQy5QsUPRNSveuSPTQcdx2rK8FZnMwK+QhxmxVRkj8/4bkDETVy
lO5bf68TuFp7rb1sY08gCX0UtsmaNtITlUuLJ2/8pbxL8ckGAWDIOFclQHZKzAwo
Idp6FwAyn0a313fSEEzwPZ6CfAQuUkIoezp3m0CcsxnGmHsdmwnNXY6xYZvOYXT5
MLnAgkjnK0R6+CXbkhUbWEVnkEWrl2XH1ilvsqXvxXNz5R2vv577TLmv6X497GjU
Tit/nWx++xt6F7mecul4kKN/SBtvAvFvFMAWt1+hCCppAmlPtSZJHZwHgQmUDyRr
1k+Bo2f3D22B317EErvTPTcOgvrYP3lqqJ07OSV/ZlgjswG3Eh/zUgs6OEGd2CML
6bvix9kG9cRWz/HRH/eiM//rn7LafbK9XLngvSNuSUgx7Ob0Xuw4YCiGJIgWXwae
12Utj8R2gK2cmWgzBT0ql1bDvLx4wNZJeetYEkFQbWoa2sNMF5igVFFvfkMsUMY1
GVAYX45wR2PKraoQq+w8F0zedhOc6CfEgt1GvXjpvTe2qdP6rHO/5I9gQoTzJaN6
vsiWV3PYdw+KI4Rt2ba4BmItVe5MPVPL2Y9s3cZ4r/Yge2u0FxaQ1zdQaWEcs0mJ
XgnDAJEFU4TxjMLVfHIE6ZOb0JFKqIt3KZ0upbz3Oc72hYaEMYAoEH4cEPVYV0sH
f1wDwNGtohdc5wy+/bVYzISuNLj2A8O5qItzdp1mCBs6bMB1iZHguRW7NQB9Bcbh
qjHtLHT+uf+Djsoz0osDcnqrxOHe4KU1ZmcEUI7s4P9eykb6zCJ2DNL1s5T6xjDw
Ot0tZqlyzezusTYzVwJ2IyYyMWoytLHhDLjHfKfbHupMCW+x4m5+AEw668ykmtDr
HXhFPQiDHpGDzIK8f51EombSphguJRyqQ5/2OnD7ZAfZPFfTneRQNOTHx/69xW4+
wVbN7ztOXuXZjJ2cSrpJ0mZz2X+BOq7uF/emFLB3ocprruffQreTje3MOkJfLnTK
xfC7TucihfVW0gBNtfRT2OzD4maLGQG34/q7QkXeupLHJxg/WvuKqeIWoz5ZrWXI
R+G/yjsdbZxXTVVteYb0pyf8x7kNsJ2HnKYggZWEHxeAD2ntd/QjT48B6MgxjD+U
wr8BE0GBcif1Sd2rHKNVjUKxZaFgsWD6Fj2DHJx597AdOXhKrrCWW+6eKyUV51QZ
DESqpmvRgmvxW57J/uME30zxHPv9Ye5WF4c15+Y+efe0tt7uiqzmt6iDBMdmuz1V
n9ZtiMY4AkEP9UkYZQstKJdTudH1toKqU6SWJ1eRxoiO3KKaP1UfRGMfj/oL3Rb2
EhqMU1BY6bTy76Fw36PFXGo6BSER0ahx5KvjI0FA25qmmIAE8vKAoxNMjiKxeEmV
5d1PW8KFWSY8GgQxngNW8WcZVYFq2Fn4DezN0Tj2JAGmexi2WpG4y4GNOQ285Xq4
yP6DlKFxWTt+Tn/C1g5fvuEhHpJPnsFUaQ6lzkUeG++XhgC7pQsXUKnIY+z0D27M
OYnA+I5UWlM5kIe1D1sY5GCSe5usU/aMYL+5NT5rimvOe8a50pq2kdibyItdEnsR
e+8GFvIdQ3Fdzq2Nz+tsB9kdQfJrWagCvRFvm5nCgE3S6ZmoxMB+/75iKdJYGCF3
6Y9cE0iOdXT58k5ipTqNzbdu47QvRJOcMqkLXrm1uuYjUXPNy8H4kcrTM//zQzrZ
Rk0T3CWWQRVM4VrqQxKUguDMhIHcYf49Oc3+VLk5U+9RfjdZc/GqBej92t760zqg
AkCn86HUWG9RXRoRkXCVAPZTdg4ZlyBuQFz0uWPU8AJH0SZjqPtbabA9WmQw+c0f
6NBbB0nPRfu3eNBjuGABywvMk4hVWPdtbPGaF/AtloiS4fSYHwipZ1SzFBzdVGtD
ZjmryYQqg+G98ul3+okTZnAh+bUdqnx4DRn3hQUm1l5QewnCaVOqjSa8b6BbyLF4
XuK3G6KNel8l8EWCUTYX7iOUBrYIuxcPPBuyoQBPJvyptub3t0HZA6isE5n2TtUc
RDVACxi7K6z1OtVeJbJAbeltnByYgw86WLzl84s43SE1qI1GGB+OMiDNNBbQnYtB
qREkgsK2SfH0ot2v1gBgrCz/Pm6OrJRH+LNWMYA+qvpxzOG5uIIi7808Uj1o6Z2A
YXmhfI3hr0e4U1Lm7AP6bMKcH8kyRbDM/kAgTVdWXsamOurB6uGA3zwy6jqfeNcY
E2SjoC/GL606mgi3s2FkTDqcJhs6sUoLuF3fJQ4z4XbQ0U5Za3KzUeeda17/Khro
NMcypZYbi+NZD8R2ksRVR9+9ROnHcK/hAbwp31wNcEovU324z57hMAG4WRN2Lzlr
KerRYydxeaMq6UW5SPQUVPMQT3C28GdcXjNvXWCcp7ChmF74aTfl+X22L8GnNkcg
W5yovJiy4JGRWGklhIi9z5dzv7mnVsdQpo0ogawfL39UhCso+WaWaQTwKl6zFdWG
1eyNBhYr6pxbO3CBgadn65SJKWPJ/V9qPF1ZkkLllzNxSrMPy9YnOnSn6mYjwH0S
GHaie9GlFy5CqblvY6Nf5pK1DhjuMsmPJFE+Bg/FzW9BNfOQL78UHIXkfsYRR/Xi
HUZ5u5fqw5pluuMaGt3qKxuW4ZKebmuQRZp8rV4JIWw26bB6ohybs9p08lG4ad0o
JkGpW+bqD8qtbbYBd2+w3BLPj6o6QcvsKE25GpSg6rKXi8/K4jIdfwJdvgGNRoBg
D6ru3qGyhG9rMxSd/3mhhAlAYmuAVE3iQR49IZAn7F/kjlDJfXINMYZydQS/PsNo
6SS53g75lJw1u7P8f9q8WwV9OGoXJ/poy8zoNP1vRXTloSbpQ1LpfiIAnu7J8kyM
LLkKfc71ETlDCxvFO7W+TdrRQPklsEbJaeAZs6iPHn16H0iikGYB++ru3wYH0jcm
xNa8yxB87Wt3RCFZLBcOp/Mw7aIBmZc0UjN+kHbCNwjxo4JmidPXibYWiHpZ8bK1
+g3W6B1THgczQyNBrxldlNfcMdZvvS0R1w1jmTvRjj1591sBOt9hGl8ggB/GKw0s
cumc0BZWsIYNcbdpzLL1spdOEiXpuC1z8Cg82IwnyEIK/2OLEcngDIcwlwWFeWDP
TXptQiN3se/CLE6wgsMQigWaYyFODqv+IJgZDIBovwLeLdFJha3sjWPGbmHo2lFG
F/TrY+3GILIxYky16DFLsivtfghVNbksQoT/zkJPWdZlE5p7nRLpnDc2IkieWv2D
dYfT0ikMlIUYdyqziM6VCY9H0mg/+ed23R1Dt9ydXtWXuJiha6TetGg8eX11jKad
dyhVgC2+cu0uxPgMqZjmtsbFDfaWGc3uVWobwLeEfJ70K4HqU5Y+QkvD5LUJ8/9k
UnDOFKebC0TnF+dUyGqf/EcWpZ8dyj2Zj6SPXKxlcXjvO1m2e3os2HYRp3Q0ioWF
Py+1bKuSNIJuUxlYgfW8MFZIfhCLkl+nQhx0nsJQbxJYUnpXllwrIrE65q3EWwpw
zW+dBvyAXKag13J9T3mMs+prGPA3tfmkYK3f60Zh1FUW58K/kVfaNvnrL/SIr4eX
ZhsGMjvw0U13GV/VKIub/UVP7m9xOxC2F2Xkr70vpw2Ynp/qB5Qio91jRQYZsc5S
0PiIyigCsCgaFg5HTDhYdYBzvgRBQNmjcnRaC6n6nJdq0nB7VoqLEDLcEq2o/1xR
irYwqTqqkbcM/I8U9M20kA/NyqiaL8iL65GmBeIghFKJOR+4dNF2k13DlEDj+MWo
gNuYaJd3kU78gyRYb6EwV9PG3NiuBfKUD1x4wzqibzW2blA5yAdnKreOs0fQH0hH
GC8/1u6feHl1o8XDaTdLxhb0T7Ril5fle97UqKMVNgecvjLyJggKob4VQa2IRf6y
EeMlvOdtjRJN2bzSftMP2CQkk35UWQe0qwFal/IJh1k85Y+eUsWe2GBWuBCIcSbF
mz8UYdfsKQ4JCOGsTG0qBT+5oNPmiKXkOddzOxix98BYi0LTG2eFhB7hEjA+N8/y
6WKDw19OPQA8hR+GwB098bLiIg2LZeGgPFnHABofmWcW68PRkEK44bdjBraVKyfv
0wFifj/9LDExd/xrDcspfaS3/GjVdE4LbvhDq7lOhD+wiOHVU1Po7O9RMaznvnsb
IuGBGDiLk8MJcwtIynxgdkfUYiJBKfRs22NZNgYdUCk9P1LwTUwKBItcLnFHf+8r
whu8xLfhNQ+HAG+IxKP4gA+87tYAQun/LYcnP74XxGXcf8HxEpDUc7Etg+6gfmuT
J5htGmhrjRbJEXVG/ORXCA/4DLFpVbMIjA2FrzQ3iJLfPOqY7RdyOpy4u//hzCoQ
5/xQh7lT/k3CcBLSugFTR+NBxq+XyvdHJishGI+2A0s=
`protect END_PROTECTED
