`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WFLjLCjFIxJqPDtzK1hslA8FJgxHTRC1FTDeF25iW15cqFRlMaT23pThNsMpTXmf
0Wm0JScqWtcbusk9a4OlhuLqhx8QPGozeWDSumb+rJTTGRULDyomLQGs4LkeqvCo
k72VKAPO/rFfpR2aH9jd6za6E9yTQzNyvb0b/pD97O+GQHdrHVIi2OnfeXVkvYDL
EkOGl+w/DfQmzWyVtN6nltoq6dzM0mmtXnrPzrBcj0OCjyGy4FWBqqDusW2n0aIW
VtF2dAdaFgsr+a2XFUBTMJWkYGF7NH0C4xfSWHqXVz9mRqd9qXs/uXydDeKqXxYT
cvvAg+OOLtlzFKAL1IHPDW9bwSz/uwn2u1oun6g3GMiLWJEBOJNmC5kVOf9ymgna
ArHPs0A3BtOhL0iMXI3IpC1ku3PVheMk8eoq4XQfOL+bVofY+tBQ72K2e33DLU5M
FNMV5x6GHra6oSs0W+Hk8g==
`protect END_PROTECTED
