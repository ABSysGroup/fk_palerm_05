`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8mhmxEXrHb42WzGsU0kVBPZz7QiLjDm+JNDMecHkia2IEqzljM1h1lJ61kKe1qRK
xcQViaLt4jL8OVjMibFS+t/SpoVHvGNcYK2SVB8/jH67Yj8sZJrfE0yJcb94+wbd
wN+yUFmm8xMyaQ732ioPX3xm6dqYX6XHgPFh1jp7+sIHYysLzSeLINEN0QQ+3oww
O/HIqpQH0ZE0fTFcS0c6UFEd3A0ip8j++fV8zB8wTg9/F7J+HZHdrbrFzjGycz30
pkkPsBqyNs7UFwohCIrDweIaGy0Whcr0zgTAmp3w8/PulxYmY6GKjuYbDJV822C7
Q9wUfsL0EccfWxJ6y4SsLZPdUa06jmRERsu90gdkE6gaL/fCsCU0NePhemjm4ToS
3VxBSpqBvDszxUC/Z/liGuFt17GmXPjGBJ0eeZqq/5rdvtzVrNXkKZPdIw0tl33C
Q0GEBAbYp56FYvE9UmeODGOoeKXEl0VBpc1rWJwbSOYuvTRcC/RA/PzuK60M2/D4
OW8yGHEGf0gKMySxuTGptEHFA7IZ2olQsZXEhXSpCHIVybIMKz5J93OXRj3MQZEz
rSyNnLY/j2b9qlZoLxzB+OEPAhwuKWZaMbKTo3g5Ek8da0IqEN9H2Nakt1yzjXxr
2ghxQPue+0/DDYBWWIgb2QuvPNSe3+MWeAhYBiU5TI3NJIdqpiUlQVbOcn+iQj+r
KcRREMC8b1BIUgMh7zq7cMv3Yk8fpeqgYU15gZPIjWsMGlA/njZ5I330TC5Bss2s
+2/7tJWbiQfsR0qD/m4tpe+bgIVujzocQsO5XtxKlO74XECx08UC6jyGp16owSZk
EEkdfn/HUzdAAbKk5zT5WXVOFSSnbxzFQK3SvdxBUkciQJEI/U+X5es0qaD2qntY
HdfCPycI2Paw12m0jKtJjZ2bZD75PTbckpkxgTAhYfIzMfY9pvuUfg2Xwhv9Poe4
Yuj0+9Ce0HqxTY/Ql+QHG+yKu2JpTzCCkJ9g7U+caQt6pZ0rjjdng/5lFUnDjuKb
3qXZ0pvuMtXdFjFgIe68MZIg/DlJj8/L26E3sRDu5mwlewEasbseeRMkP0k6afG8
5eEl8Q7bP5lweNeZGDNIyic8ozo0uUStOO839CmzgFLSlLvnvceGeQne3NBdqY4x
zLQrEsyLO4G14hr4TJAD1ukafr9uc7dZi5NxcqdJrbF2KAO+3IPz4AtEOGQ+7dLY
KZxoM98dwj6OJaMNM2RgwaE+ZRx6AkbjJDIUGjs9FNqLkmOx1z1EUCOm/WazuxSH
rJF87SP2bXZH1jdWc12ER6BFDNqbAOzMsFqNQ0HALT+bbC5r7jR1NUB6+tVm7RwK
F2G4KSO+BJiSYPnCkyoJ1q4OAV+7Xl3wTTEs4ZJzZZNZ/tpIx60C+cqqvzHEUwuG
CQxtsOeVahyXEvE2AQw0C8ySO5DosL2gzRWuDcU0R6CLvWoYYY9nNGqmH3+ZRSOY
Yxu45BsT6Q5SGFWdRVe9O4YeRGNzFimqZWB47ml+wW1PhQPXCFscNmNaAubfKcEj
YvgdORshBoBCkweOhL9vTfkJYOtrI84bBNId8nIc78NZ9XmWfh8VR+54wUUFh11x
a9KYslDUOoekB7roh4+WVKF57MBwBcgxGuSpMrTzECRjOSOH+IcynPcgzNV1n5yq
PSoiPut2lhVnay/RkuR4vtANLSnPl+b+rwAHCEAAbBBw/DzjozBS6wxKB+4j2gw+
0nxerjx5A50OcKcqtzdKH6FX7Fm4GgexO5keorpkCQqM2of3GfiO9xoENqjSwDY7
D/ud06CgHbmNvh8f4mfOE8Fp/ioFma/htLkg/qNnBlTUi8TXHYLxXVhjd7n27o+C
9+LeVVumcSIpnXB9Jm4KElUhp4TJd8Usrufv4PSWMhdq60jiOSTxMf+srePy0I6g
YuDEOUVFZPtbbCovpW7ZDUUG/dbnOZaRxIpVCVmzrDHR9bdWnSW2kMXPMPRhyoua
7nkRcZCXd1kdcbHWRbPMLXlLmzPDRigwyBrYhi4A+F/V77HJ3zDRRtz8cL4lbVGF
Rc0PL4/caglmGT35bQc+cKWKO4dXz5tOXxBtq2EJmk4hiAUV7+zoJ6XyRUx3L5Qx
aJRYzU5//guU3W4MQdwZuqUwtegYxafdWaB2ZE+XXCO5mTuB3285TdyfyJQvRlNi
wiV7jXwElkNtc6Z+xmoUImjSGS2AGAL07RgUBAzoBvrZtNpHl3IylB+HteUXzNww
XLo8pPJUfpphuIMvztV8AneinYKl0QJtWSkEZbi+5qVer9Fx/uSbPodR1Fvoqix2
FWj+Nt9+kA622+plMpXX8u43+OuVJ6tQrVILXIhW4djQsND1mCQPzCsr1MUDFNsP
yBmi5ORgEq0XW7uoG230Bwd/vN60YHJupDMfcw3yoqdYeGXJ6ofHMffTrwRqIhX+
1g8OkBba6sHr/UwRpdXdgMT7mzhl7O230BZ2RkMzkXyxnnMJ1t54qtzxqX/EjgOC
PCNlxRxwzujUpzyZbj43HfVqAy+hYLVtwTQQ+6fzl2fk6lR5RLax+Cmm57ciIrEH
DpFysJ08l4aIqCaymEOsi0a2UvAe4/TfdG5Q3deQ/1w9PAkca/RfVzD1sjS2hDUT
VoD6RSasnkWSvJO+Ly5qIuNu3EFXeUr9QSHlseN0Hur9cSgki0PyUjAn06h0u2sM
82VtFsZ4L5ZHfenMCVz1bG18WyWgZm8CAhXI2zXswhO1G5W8yzgUIs2AbEC7NtRR
rc9eq+DZrRSOOpzxPCNuCaKBJfaXtgGzrv4vMBFkJaLGw7iTLxsvKrliEph3JQcO
XqG6D5tnka90ts9fBOvY3BflOaSymbmHHU8CVtMQ91Bd+ZEWpst996fstASeVEQT
eB2xfvV1NkRg8HqY1X/OrzYNkieehC6mE8mFmrO4HuA4Dt5TwGZDPvAJpk0vB4Nw
Zg61Pr8ZtG7RaIZ/PdpRVrc5dX+GqgJFaZNvFnBpeJygvj5IgGg18C8LSr+QNGyh
Dn/zKVdwIWUV0oOS8ex46a8CEoO3Aq3i0ynbIOQNNtEm8IUYj0SjDk0prKrjUvyE
FhNQUKJgrL7hwnaTN3Sr1aJZeYArrsQIjDaS+oaCwTvEI4rhTnPSBT+jyLXW6dqE
uJ7yrK6EV9c5NgMewnO7hBhjklQRccHMJymqzBHdg4wqyWRgG4HwoUy1yTufEJLt
rQRdhsG1qHHYbcIPEtgaBn2jGEfCsUJvcHmt5bJ6PH2IyxGlZzc/P3eAVCH3btrX
Tj0EA1aZHsboD60xfQYvKrsCC8S0UEEOeU6P2wqVkJMxiFq4uckLx07hi629UExL
E5mZAYmo5hK57g8xzUPANiVplyQLmyZ9EAkb/bt8ahy+IQlkvcSTlRtZ8+tZe7Y3
vIcyipK8doGFou95EJ2Z+L/PCVDf6R3dc/jEt+LdXOPk+HKpBwg7CpKTzEIwKTln
ZEap5ZH2MChSLFXkcVZzf10khD47/tNM9+oKshJVpoCxdS/RlRwAU0NlasUbVtMk
ipBC8mitSP5vqod/5O2Mf1tSbAb8w7Dmcj4OZlCtpoUq07qYdbrSCa87TVwm/0/H
Jq8p/9GfBalHemutmjnRARLYsVEysaYcRZTZivy7Tbe6dceUduMtu34tvPfCCPkn
rfd8r9hgf4q9p1BEg0Eb7VCbko6/Ney2YETJvV6YpE1ebh1I7oSerfdGzP6CFgSg
jQN20HkGGEdw4mWtNDGNSwLRQgf1Mq+0xmXnwgLFg3YcjojiOJjBZikyAx4bG6f/
EBcXbAn6w4QxqPx9IFXXDIC9XK/9MZm++yWcHMrlefjlvm1unAP1wETnCzLXyC4K
+4vycdFalEnhjsh4PViO1UtHAOJaSlQAVUduLaZA/By+ZYdBY2yTa/b8cSXdnF5+
DiZv6j5JR1oKW5gN4aPs5d7klZhBkZNspyuQBsXTLH3tdeD657+bmH1T7tD2/E8a
RR6CIUyxQXWKDMJZlGdHmtbjRvLuKFrR2f8Zoi8oTB2LuuVk+tOK1wEldxDCJ1eB
pBU9YmQQ3jS17PKTxlpkhg5SUQBB+ofWFzjs9XycfR7Ndb/HbKUNvp2Cedrxa+9C
zXQF5sLVmgbpBb3AtVBWrbybKf0npA9iFlTDC3hhUes0dwBn8hd5Nelz6PpJ2OUV
K+qVTwiwILnKTZTnkUpRTzYi8NIWQ1RvizGh5CBTU/6VOYNKHoHBWZ4LuNRuCrc1
jDLb7NP2U5YgEbJrr/hP8+4hBUnsXiM/yGUhEaPwo4RnOEHpAIcFGZyOVYCxCJGG
C9hzZxXSXxupwbyaVajl0WeQCyHUdqSxQcxWX8clqiVZOdzkc6QfIFxA0/xhbGaP
2OCQqTA4VTi2R7LCEJfCDcgN98MK/w1Pp7XZnzif9Zf3Q9bvgIBkDILcWLkd/pFp
zcJgddYPgraZpH1gIfqnQxl0GPusiz1UYx/GwBDDgDTrQ0pDzZ+1E2YAvkjHdXic
0sV9Iso0ppQ8SQjjOtXsvGYwzEdcDIExJQpsC6eJTxAwy9cbmxBgJXsup/xkHVbQ
tVw9/VKKZLAQE3d7oikkIINqhanmQi/9XpviwebOMuYmFdQ3sMX/X1dzqijOHEtD
xe/lUaUnSrXoWrt+njjjxvnTysIJA1pCv9ofS7/xDkePUORKFyzZJseawsChwDlG
6RLpVIJ7FP21Uo5YbY9hHs0KoeNlw9gvMvguSxW6/1kr3a6hTkt2yVuuF+gh9weP
D6DDvn0GC5/270ruEL9Gfm8nGeDIggh9UgkQRDN3aVQMAUgqQxSebwsueNJSpcC3
UWScOIBbX3rPn3pW7DbZTuzmtVaqy30ukDyRVYUImZ+YmWKgGnJL4jWS6HpznRCZ
kSzIiKbNDi3XIFezgJW9l98bay4PDKbAGeFKhPAEkLGL9A/tVzoWzSwhv949r8d2
nBQnSBW6mWjWba6XFUtpu/ddS5EAmvOU8Zh58eDCs87eLN6dxQs7JmDn8ewknUu+
KzA+eKnCs/YeflSCXenm9tK04S3XNnfAP/OVu2mOu5IjxHyHvK8tu1F2YZJk+1ug
59kx6QGhX5SNWkblYgjYhXnSDuA13YpTpc2rfxqeV/Gj9e8HSHYFd9serMoJoHg/
QfhC5D96EU1FbSPwyeMyfgumde9SwPA8g4zgFFMdboU5C4cxkxeSRxEpXZmDAC0L
etgDkDa0E5tNQQlTP3E04ZACRT/WEIJmh+TjLtdL3bps8lPPuEOCUZJLvKBlNO9Z
upjhB6wacWONhR3Y+oXO8vj0v3sUZ/4a8h6xXZWaKKDeLQZ79qs+M5mrKOXpEGPK
jQgr97zypXgfIFEW8JdxwTxXiGzfR0q+8pc6S32lLShutVP0LZiYVNidzfjPBZlw
OQ3IxhsbjHwY2eyLG9bruub4uhhd4ezPbvm6+ipUrnN0DnKeWRaZxzJOl9AkRvIw
REx9yPHp6DpkF7Bw02u6RxWvEbXhCLaGZ+OTken8WbZnvtHh3v3FloMc/b5mrwlL
JfrXckh7EYtKPXXR8Up5dvkXK6BeD3QQo1mIF6U6DJQ3k3YPsUqTFqM2V1G5CE+2
EKdviHeLz9gS7Z9OJSgtCiBufSEvbPkygemh3PNbw32CuHh0T9qcwLo7v+z5SNV/
`protect END_PROTECTED
