`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EpTXZWUrinV2xzqQrzbD2WiqK9dYBYHLQOBTSKHd8cCx4D4SQd3TzweqTl61KwLZ
4FB14A/FFA8+kGsFr2dZCH99WwtI+YMj8oktmywutWc5Hi5hu5VDp0+iNDKVLWjS
ZfbAWsR1NXcw8gJg2Bqv7rK0i/7GCvbeIPd0GFGEnPnB0HD9Lpftax4HxkHQn+Pb
LOZ7tOm5V9BJci6if1Ug3Fdh2EbKXHtyfZ1NIR4VMsD3pmM+qYIb+Nsa6evvsdaT
hly48U8WoPvUkLTwUYHYzgg9DTaYZFGhODplCSKtCDQbF6f1qIPaMKk1n0i7bSIY
QrHKnpE/0ATpZTl6l4eT0Jczd9i8xDhFBbbXGI548rGkEUe+2m8rDEso+EQSkaiT
F1TMKaJLDJbrgBxelYnNOjo02ECC7vHkgCXEotmqP2QpKp6Xy/Hrf/eTZ4x1udHF
f+X9nSUxOVrlUwITfCuskvDCE4M9s3nWwJ/HrSW5wH/t3O+ClCNgtvw+q9LsXHzf
FQKTCLJtO/AJSnypWrBpwEZyoWDwxdRbaHlhYk0gMsNoYaUcGFLG37pCjZ0xp+hx
dAT6b6lOUsM78bfjaGOmn/t3/96M+r58tt3Z45pHIMKnN+/STMMT17poYHp4m4Cs
wvnvEWsuVSh0Y4MPKyiqi0KknFSwV7ssjHitpjE0xrRNQTJzuzdAf3YJ38W+sufA
BFT329v7WNVZOLSDi/CBoJiGMeKtOCmkHHcfJZINI8z88bcPwwZMtvx7KG5tsxh0
mFOd8s+giO63E8lejy42RgA0YSzMLg6q7/apqXIbi+Dut45a6NeTdOaXM0pfAHKZ
O1Aj7KUx1QrTCHr+oUAKMpyhdgcY65VLGs/rQ5qIranb+U2xSAEiL+VVFrjR0sa5
yUFZwhKtsgIe4I8rcxJ9qw==
`protect END_PROTECTED
