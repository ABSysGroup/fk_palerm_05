`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HphfvmUcjhcEJfpctKLNUNfsi2EKHnpZ74DloQ9vAPC/Pt0Qj0sc37uZbDdgglvK
qsf2JeoVSGGfS5V22Ag7q2cx2eMzHYBf7h5Z0UIuuI/GTywsM9BZCq73BCIMVxuv
rD4PFedjxRl05FY+2SVTVI73Q0pldFD5zm3ks1YQMmMWIWHwHygvqSGh6LrZETbK
ylRuNzRsFrg07gk/fDN1UsSHsWEYP5PFuejX/8IH8dERxxVPzfRWkBphA5R1nwgB
x7F+ntASdWxt33uQi5S5GvqXU1bWTS1SGT3h+FxuZmsUvqA2usXh0gFuBH89oOhY
G1gvQQIZX8O+/B3d1mpi4+zu96E2YbtqCQsmLnhTN+Knwhl5X+h2ii+qh1UBEvhh
btnETvxMDcODVYx2NPtIXMSpGiy3GST0xuXWUwxyvBvyBm+9/xbegaeeEg07OYXb
NOz/YYtC++vIdjrUmpPf/HVWrClkH2YxTsj8A0dTzr44+aZB+aPsOQxG4UMOp7d2
QcFd8AkOwu9CyJ/Z8FdJJ7vdKiQTNTGOUxWuI1RAQe2ZZqQAgewxEB4fYk7L8RVn
EGWnx1gFWgIN9Z5wE0If39jUhD4Hna1xcDYUXZG5bOf1tRmNz3yfVPg2HxdEaLlY
fj7oaS3kqxNttkj3HLrSpuiObOHR0PrTaULmr/aG1AP6WUeIeAKE79dsN1uDpidc
BhDCXhwm+MfoLHgCEjVDysKEBSprWuznAoOclwhjV4atqkjAvzcQzNJduV9XCuNM
/vcAKMz18PAesCh48LZlAOgnUugXDZENoL/+P2admJbSXkALN0Np/xUzWDF1UpZu
MDxzu/jrn2osNYWYsWnnE+ggPAj5hujZeRUB3ypqQtIiaLdr6FRc9yDkOdljy8xq
O+WdMyywZurioVpxGGZ3zz/JIURF2ytJchoV9Im9AXdc9Mj0MNEydCUBeib7YomD
iHkz57c6R0wPt+AxgwWLry7LtQ1PAfCyuqV9jtHLjF1w+wjDGzAQAltPdXtoRV6D
9p2NxNOjA2+8A9vyFRCS9W8Q+ZQCiuYRPFSn4m12UsZHvMfeIG3V9YOzkwWmssKA
hXKInQrvHmZUDaLfB/4sQoWmvwD3eChKfdCOwMOTxDKenKJFiE0OUZwz3vb1IL+6
ebFaJKkejWAyB99sJeT29kOZqFc1UqpPSzGHLwS1lTCELZtsFSRN5376jhHrRHgq
BejLpLDVaVzdMVB/PJBdLd945iYRDd7ueZuDUA5D92+/PewT7djSTzVIYhbzNFxp
92CuUm18AU1Nry7SdALGSk3UXyuitu8/FiHZfZIjKp/Fj0wrbladFfLIUcdGra5k
`protect END_PROTECTED
