`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
opE7z7ajImDsgwSAFK1oPo3FXiGI8ZUW+JRtWqvM6wFsA5BkzcNe//DuLYQz2NPR
Au1arTm4uJttXPHxPW0k1NEoWqJj6f21Vc0RNByYFiNz1s0eqOXsYQF+yUe2h2X7
fB2xUZyG4uSKEDxclTfGGEqTbcxfE3N27YzasZ8aKfGvZOvVEcg7NL1BOxyFNWnI
L3ZDKEjAdW6gE47/WWltpGJZxF6PdQ7mLvfk2ZAtPup7seDvCiAYhr1TwtTs35eK
Rd3Ttyu6bygNUMqnd89IT+DdNKx3N2ibQmCJbYGwMyZtHADxaYsPKIwtM427yb3f
QgdWEcB1FkV/fmJYmIMSkzYn5SkbmNUfcb6l1Qw1M0WG1yQeGnEIqKNai7XQWuhm
aB/JNWhEjJrC4NPW/yEnJMHGCmcCLPEWNH+9ENrsu96icgaWTFmlqfkfrxz/t2/2
N1bZp34vMVHszmIEN9HjWuySyD3ir+HjeZ0gJLOB0yokl4jDGWefEadIb4WdoKTS
0mSvi5yQ/Yd7iPfRlZMcwL/8updgVM6kz0TezwA3ow3nf/uaZJX6ge29IfdP11p0
c8eBfol/os6jkKNxIgxeokp9MgPxWAYdUx5DxioaPE6tGXv5d/fDlXxERg4LKl7a
y8C1SxmX8R1dn6IWEt3y+loFGE1MobgQv9PPDJtrUi1mPigcnnnxo2cCTF5F3CAb
P+0GAMRdxuaBHi3QlomXX43PQ1Ea2/wQHNNkppsQRDH6DVxi21roMpLbhIHqKgng
3V91UxQ+7SRaLWVZTr4LsRqq9zr64ljm0KgRw9GmgQEoI24umkxD9wywXSKAzDOM
R9x3Eh2VR9GBFvlhzfUJr+H5VBhL18eS0OK3TKsjYelpwKwf8avntBrtXQvfX4k0
mGrUO25jzzbdeZe4ZsVpKxmKS7L/5QC+bjg9e0MxHD3sIxcjorfS4/sdepU8q869
G/SAIL3Lj/wcE6yVI4i+/eZjzk5DcCIGtFSWFxem5SY=
`protect END_PROTECTED
