`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ln7mKvs4jeQ5qCM7S+CXUZnEA86AeAZEZSw7DaAOkZIGepnsGo+J74LUX4mQhcRn
wbxhtqRFhF8sHSiKQ6IQzf8k7IESdu9viDTmYtw4bg8ezOnVH0CoZejJ5kDYaoGM
acWvcbXwXV0pvNfGHfF12GICtM+zf9Tq2hiOuxqbP363OoRaqUSqvzmzKbCHRSIZ
LGdROWsI31OZ9Rv+M7h2W7by+yN9YnNKFIPRwekAjiMUkP2xOE6z6iUR4389tXoG
jXnNcVzbAqKUwpDotb2zDL7XUrmB0rSSuoIS45IcL4Ckt+Ocfoy6Fggs1DP1M9dp
P5tavW8982i2/lt036iEux2iWpa2B64vHS3/owNSFczvB3gyKYozTYQpdC8XexJj
e0rtj2KZYOq947DO5O6mnFlafQIk7I5Y3ooitxFC9XcpcIzbdKo0BhHUoyvImKfC
CIW6yGrYNU4z/8xstR9K9TWRqCuRxhdWhR0va60kITQ3Ue/+UvZfBJkDxoa9ps6G
e/yKrbteoCnCFffm8o/X9m5Lw6Mkhk7K2++rYP0d5uPxdfxkbIFFCGDP4rbTwSZe
ROkutWdyelxiElOkNc/92/cHY3p6i54mPzXSNvHGXE/0lDqls2sBvoniU6ycqaV5
kw2i9Z8nM0OofnGhKCJcA+7soXgv0wg/YL5bRLQ9Lfiknfm8FTXBUtwMDoQvwxrf
/BFkcsM9qM2L3UVv+Cjvx7OjEnymnnqG7dbC7ipOQ3m62YrwFSHKLW2PB3UFi+74
ughvIIXmbhldoZk+fiBrcYdg6hsju5bfJnlM6IGNXj3+DIIfKqfhuxPhKL+aX99x
5C0PYcK3kQdGFVH+WchS1oQSR//bggy/ltDCZJ0abrvMmZKq2iD+5l/Cv98Wq8Ie
741jGwQkDw22XHtp/HxVzrRPui6SPW9bHoqgAcIBJ3oT7LGsLYObzZT28IIZfPVL
nYZYkiiNcmk7OHGhvwLgi/MMJVyX9omfnhAEd+VIGFDMAhjuS0+f0gTDCsotNyJl
G/HsMBsCNcQcjNOQY9fZZtYBZjYbBmtg+Ig1qXt6dHbDrUg4dPsnsMEMLgMQZ33/
JVNXydZ7oWYmuk9+s7dpYZ1kkQ5AQ/rml+AEBLUc43WwQkm7qg1Nf7pgU+4KlpMt
MDt0KlOr4YsBZVvJjhARm268nvB8NtOxjdYlFefEpIDAh/JygDPmtz2Zz5BdBGnG
e7dTvvXKP+ihfFCqvj11FSLH4Vz0uUW2WFFcAFUsEl0p5gzAbIiw+HUBZPGv0Ppl
jRJS48mT7k2ZXAjcwUseC9JRo0pldpmLkqritFRc5vPjCB+grL8C2qRKbJ/NXMHP
GpSEaUPgNjn/SMp5DfcaUtXGGa7Laq/cC12gMZift5SowCqYKkOXiAlakcjJp54G
B9Jrq/284KtqKcYCHg3tw/nSm0pwpfN8NVtAfMt/1XQN+zBHRTECpQW0zgS02kpv
HW05PCqfQAgv+B/znpStfi9vD75obRvrY/vNYrEQtmocB+MUN4HOgvOu2VsT9XeX
s6HCf4JgFCYexTuVU3WeCimBIWb08D66kMu5AElBN8twtAOJYj6nazNHB3Z8NIjn
PtI6lJoQWIS4YJdOx7VGb0dB6+8ZZvWuAHO4IutFjzGbZes+JIbRtcRB29yka2GP
f+fGAmcBAIHKzCIHg2ib8Qn4dZAcBNSg5hxW/PVOx3HcH+WldM8l0QLQKfYCMCfR
Bem7jbf4xTQngk5uyXTm1yoApytT7MmU8CptLdfFC8cvGXlolHqXIULQv1R4DpAH
Ms93skL9Ab3NKvuyRyxcevdA+dw4QMWlCRjTD+w4af1kRcyFP6Qb+b9SfvFIX/wk
bCf+x2xaRfn4oA1CYxfqLPvF3EnlhVGpdl6Eihc99W5EpgLyagATvXt7puC66zDS
/mCR7MFbMoE5dgi9t/UXOGK/P9PJYTcEFfyywlttHRHg3W8qouXNYEoFxSeLOnLx
06lpn1PirDDDRxJhGIbXPBZCRuhJNtwcgOq6QSdsEmfTui4KBoBswsnIh/n6qzBx
A0xAhlZ5gCJcvShxfPbSpYS5vFJfrGnsJgDb0oVy7WGXyHi8mhkdZDurtPLkwry8
yOSRIYZ1MjWyuKyAqXvU/IrzjVkPloX+EYT+9h0RP3vIUPUdBMJpqrWKWw666fO/
6Tflhu7QOjvK+T/hYJthph7OSQZ8y3GDN0lCZiuF5nLLSLm8qdHjmPVqla/DDoDh
/CkgW1Z549V4JfZ5LoCCB8XPKkhDows/eIna6UCtdYR0oSFkqQmKLTskdz+7iprA
Vkwuh0BBipkJooGZgkZkfze5t/bPyFoXDKQrFBkiTlqMgZ5mURvTqSrw47HTxHQN
quRoMXECJq4XLAbJ2QIgFuheBMYM5aSOB0oDEgVC+ztaaMvqcS2hPtj9SlT31wWX
RJszEzuvqIbu+iNwmbPvjCvNsFPEzJcpYe69uc1TRlF4LReC6tSSQCMtHQ13fWpb
2B5nyzYHeaNRAFJIrEr20AOhTzXw04t1nza9UvZ5nHWUHRKpiNBneqd76ypw9KGN
a65DK35aTJHplolKhrTywPZda4JUP+T16TPbTSRvt2LpqK3TJPUniPkBUBFJXPFb
aFtyzRoCHeSaEI88oxlBjQY5vlrJQrS5L4roRqK2a74z6vHR3o4OaGARqVk+MaCr
vyGtp5388bQPzYVLqdaL5bv8mHxNYkgtxrmCPZleQrs+9l2CYVBgs8HSkWLc8Euz
vAdbL2+ERhUb3zgvEfTSFMwOmK8h0zMi+Bw11LijGV+AXUE5+ttgZLUFFaB4XCnR
IFBxjoQA+jf+dNYrM9DGVc8hqHragXZiWeR2s4oCvB0i+nVndT3AcbscZo+0O+DK
q+InR0kHsJYUA8BQhYDMd1UEdJJclrSsfzSMbf2X7LOfZe7nkn3lvzgGLZfo5Cjm
YynUVH2xd8MzhtbqFtS0+cbLVDsSpUR89DhB9yKzkKkn+es2fB20tL25qddAVJWx
/OCRmr4YR6PPRLim8yab0MSnMNAFhQdcD0MTmUCmV26lumVKj55lFqya7Fb8bu6L
VZCGGkRI1NWDYUjdiob2vt7BYwrEb9CUhsioynQf3iZ6aKvO80YzRUYHZimknWzY
vK8h6KmONsPwuougL9xlfVX0yIk2kDXj983bjmqj8c2R3lit8V8uXiFC7jigCXLf
04I6qvO31u7xHZK1RX0eOU0MiTvDfBWEEGkxD4y/Exyfa6GTLhinU1vmY2oak4qR
CdDfpT/U7b1g1V80Gc/JU+xL3z/pa6o62QqXZBOMhjPmAZAmmaGZVAGCgqTeMHfy
P3tGIC84lPmO42KyUXgFHBbg6FxM0Iwb+yoRoHvy6qO3KDmPPZCylMaZJLnsKCkm
mOaPJPj7GltYMiI5zR8+MPyDyD+sQLFoLHDRJpOqvx5xqagxzoMzDZcSEJ+IJBTO
gyVVT3seAABs9WJEcFgierlS5lLoAp2c7dVJ9uD3UT7auXm/ekCJy5g8sz8osAOa
b1ibDQF8IvgukTijf8fu+DyaSlG3O216j7e4Q6LGS+OXXi6lNVzPiFEFl+Xto7Fd
C7B5K416kix5emAuhmjRdYQsloPobJ0Uxjp6ovkwKFUsGH0HV/R/3vFa51WRT40n
wy2PkTskCfGAHf0KOHtxVhEz6dpyJR3hWPil2bmsT1m+ifCTAvMHXngUB8WRqt32
D1PKZ2GcEzNWjxggtN0IPxNt54bEERKnBkv3m0Vro+dKtfOpbZEAXMTksH7Pdqrk
bTpqrynJM2VBiRrxTFJ9nLSDcVXopoPJG3qKCIGisr2ePOyF4zJzzxbVU2SuifjZ
Bgtp/wGI4Qbi1x4ClO/bLK7kFJyeRL8USGtJknEQHhjFMwiFJB7l65bcD0KoZyZ1
baZs2vw3BAS6zWjyxAsZkx8Jd5vTGj3Ub3TYgOAtEmdokrdmUbGgHR+3qFkYoGP2
avzRvfmX5HSerJ60nT4BgnqZQT0oPVdgbuTdWQBq1x4cfGoGHo2R9jzuMLsEMzx/
0F5KUb6FfWJm7CD5yyDuDIJ2Liwh3xqyAU+hiP7ILlohxv9uXRLCTekmVw2cW40y
f+699QU3uHhqSM2RcN4tccNt2yGGmEDjYTzrArHrT7uky0li8hT8+FlzUDXYR7AY
9FHTMbDEyG08gU9qf8euif5UMH589Uwo0RvaoWJVl9QRJ1nGgCXHlmxb99j9Rd8G
+jAKBtBMG5joHNdNFk+5gbsSZqagR06k9kaaKOw1AtAZvN3tCMemI3Y7Qh3yvSPH
Azukdc6Ur8JB4DYL/jRn6sDA4lyZbTZ+GQuklCMZkMrnXAExqlJOxLXlBN1YS/zH
eh6afFv5RhPt9PtxjqOQTSSsrYjAq1+KSs3O74Yzw+GSzrQWpifA2Q/3YylyhiaI
yCtLCDpmCPSjVvBBvOH5kQ8qdee18fzzRSRDbNxggFz0KcwtDbLtGV5+BEgDH+Q5
m9Vbq5lfJHZP7LwfLfPMl/+9NWgP4i5CJq7YqsRBh/8BkTVR8WJ5jkKQitTeS3Ds
AibKRB32fk0KaZgJxhJxCKReiPVv2drqoqzgJdJGpuI/CJ3ZRMddkiA1DLQutaqL
09p4VVrS1fjdVLEOEUgCRIQOA6p0+Y+01oaSdjaS5LZxuaTVGHZRAzXm/zOgpJIg
o1Wgb1OeVFn+X24R1CTh5/JSam3q14en4zZFoBNvThqFC1G1ybjBvoCJCGGvXFoq
1C0JR+Lpu/g7HVnLljuSAc/etVb6nYTXsOQczh1pi7Vrk8xpbZHf+0BrU4898ytK
644lW42iRRd9bPJzA6DqJA4sn8xiK5uQDs7hMVR3okx6wTeEv6UklO4IY9W6I9DK
uoDVgnvmlyvPC1EdJEeR+gdEfspAIxQnvFeqqoDlXa7Oz9vlSn0eRjbeyoEsSPS8
bgWPYn77Pogs7TFAdIMXIfgnvDBk1PVINcBLdN/hC2nfecbOcTDhYVPDHvjuRH/V
NkFJ5tZzsTE42dI1yrRaFq3pULGc1zXpv/ju5kZJ5ep34jWKuRD3BhtHyhS/yh6O
JzF2qzwchDjHF01KItjqwdKZhULiFW5MJNb23PNEuAZ/4xXXGN8J90FEOkCZvvKJ
zdQCrHpUMw5vjIuIPY+0GRNFx5KRmTiKrWVx4ZJo2uoHrsyRvsemkhsT2lUxdXVO
6hGX4+zEyjCG96wP4bvNZvLZ/AjXLPgMgD/+05IRFX8G6SLHDLP3oJa8La8x2ZBj
KW1JWHkGWtiSsq41bhESjhwHGxep6+JJaQoGplWYwGCEfpfVe8HsKQpQ4bdIB2Pf
Xl4ixFe79pq68+VQzV54MCZgEdoDz1SnD+/m985oewgtoV1fTAFOEXKBnwBqFC+T
Jv896PfTPYd7kPpu2VGKA4RV+bHr9hzyd4OFZCmmmCc/GAdL/40REYYNJTWRCL87
RQ8UX/9CFbaHPLQNi2GrVqO5jJY4EmfyPGJ+BtdzC2TC4L1021dOmZdzcYx0EtPj
hAZ3mQ/7BuacPVxxL3a6vowcEse4ugumr6mOATeB7hftP8ei9RC+DK/IP9ZE8DJQ
FZdoxkiUwFU90JZUtdnqGkX2vzoZbWyH6WrcmOyIzGTHtfZaPdjlTQBXxbqW61FW
+ltDxg4soJ48csU8MqCEjPOyFLqYra9YqXeXz8FDcczgoCCZCTmoRM8xu397FqyE
3z2d1uoinrfvd7UNBzIjBVyqPozUOoZdxnIB+qxIx+PNEC0YX4XIi1FeuXD6Fp/K
43oBsAyI5/3qWcg3EVEFdDh1sXtEgFjVlV5B1Gs5cbyy5EYpQ2EzK22Ffucq70EG
UjJeALVq/LUyvRnfM6frT4hahN+J8v7otcQL2Chp/PW7Me8srdHzpyvPGWIBvtmz
jTmmK/rGRMFBLObgnEOXkB9KPA0UYjVXWUhgDUOylUspfeLb7oiXdF62C9gBOVpC
9OymSKobDxuLZVjmOkI6lOBZtKSw3a+e1Fi1E2OOmWJJiGMs5Fh7PyvhFVbgN8si
wOFjybQodUSOMJJw0IJGykZ8DOdOLrY8oqo+U6q4WNUaB7KYSM+kggAdPQv6kjwZ
3tS37aDGdXHLoSouLzi+tZaoLdZYvQRPP04tPKLGx4mr6cobAUKlV7cWLV4TKUB4
LWQzFo7SAh9UunaYaaCtuX1v8p5xDrZc1aN4R1+R/uhTyqk31mgCRgtPw65FF4uD
xEP0+Zibeb6XD30705T0HuTEMlL8OVbC5zJnKn4FaAZagXzydndtE6lseu80TA8G
KaatlOzqw1Y3OODbPXM1mQtBCMIm11MLpz3QwwxR4zDMaEs+MHOeRkSl6YO+L11d
jiFMPxcbWT+raTzxlhmHzuSBBS87vjKjB46pVasJS/IU0lNbG358nfZmjmoZgSy/
b9lC5J3keTVgtxjZ80tWgBzDRjJsYBJJJmcatygFI3k7N2TGDDNwFxWH7TU3b3rQ
oCfyqJOVMU+wDCjOZgj4dPawfT6SeCJiee2JVl8SBbR8bSbDvmck28xjLTA38ehB
h2xyfpJxegSrYXClFdsq9OFGTCdQjQI8E0GDlZF//SI+TrL4QJ9P5Ab6IqpqsDhp
rAa838STNwBV+AAWJgJ4kNpi29gLtTMC11j4Sb92JoYuzj6IF6QSuUCkIFfC4nT8
NbVL7+7pcoo3XfT6eM21kfHPBvvDuUJnMBZmCwnIchzfKYtf90+5R6pQdfYZDvml
eb+ko+l+Qqh9P6/a7dzRDg7lxS3OoSP9wHN0czcFDyWg8TMGWykZosUHZHhXFSqk
K1uXcrPQs9Fn+hpbyFVvyWWgDJhPPPqviV5Brtiaf71/SRHU3HLm3CcDqhWBBaz1
j9Jh33KseT/5MYpfFh0C+AnKrFGuUf/oRVqYahzaZ3Y+wvUZboQ7umKNnOBN2nMg
lXc4RINaRlREy0iZemI/Gc9VPcB9zJU56jCqjyNiuHf1E67KMPmjtbVrMAoV0geY
JOuq3Qf3AYKZIEkAW6zQH3FrLE6pcRAZm7vFLOxilSK5tn712PXcm/6Tmxx7MLb8
gnL0gEr7C0c5nbM0FOb09MdVTrDMoVBuHz3tiNS60VllSKEM7zKuTS7ZYZ8dwMPK
CW+wKdrcg/VZ1nHsUlK/PaL7ZwlhsSRf39QKfnewtYr/dZaVeBm2UBVM3WLaZple
fs33r1NGonEjPsg/tNriPQeBi95KZ4HrVXY1fA9lKeW/fwpTiF5pXhx5ZnqN/mAW
06U62Vz9Zu/mhKWekVRL0HWfuFbYsrvN98H1K0cFW70Vjmadq8VWhvW40umY0/52
M0B7SaF9Av6KlrSmkh7QH3Fcm0Gx99O9ceb6tMRx7TfbOBeFaBgDwsQmx7uYdS1d
ydUx/LnF24kN0+Jl517dOGwfekf/KZAf0V3br1ynN0Ke7BZ+9tXVBcdCBQAm5cAj
JDppSEOJ6BMVBh8QFu1/Yy9cKPnSY7ZYKdJUJKu3f0oW/wYKAAsp2bU7uS9XXYGd
/flp0Qt7mrnv2AIAxkuslnF0Xg113Sos+wIt22v+jS8vcm3nIljAlIjAt49UGQ1r
Qb7vzLcV4L+X6U61+Ie5g/aDiklgaqZi+J2+hvJ50pUWMUOjw26Tiaw3OZAVSUEj
c+awaFLnT+rdnD3EFz21JOxSLEXHFbNbPJMKKC/KUD2ZWtF98bGZbSy4G8sz1Vkx
s8bP62WXpAlUxi09WCRe/0hOK78lDp8vuI1Lrqfs9TAzpjNZhzjh/AxgGh3yT0jR
uFYqZPKHdXli1nCsRbEtkP0gbMoSHKIt9Z94SSK3wN1pNMcTVvUBAi4jnqpnwB8l
KP2aa7q73frOmc8lU7W2MltD41H1Rfq6IbcY6qDI5uerlWXtGXK2pKaqQ3Q9I+Tq
XYZvFtWYchzDco6I9N0OeHM5VwMvdu/Q2SBs2DWeb5KR6kU2S/d22BAXxzYPB5Sk
/sbhF0aCL5D5U1MPi1sg+N9GTe9c1UMH3L/o8z2fQiZp2xuqUUP9MSt5nI3EbhXL
tyFHGE3Fqbjh8aFsC9MRzvR0vRCFKLSIiLic4PBQEA0Jxxt8I2s0HbfT91c1dKl2
ebR9zAni1QoM9QaM6TfZdfd3I4/Uvu/u1i8314zk5QXNwIvkhWgq0OHBRhzt0+mV
mOD3F0+vGmPiu/ezjuD9AV69pPN0bXddmM1z19f6D7CimqUoeyY0D/NGFTsmnbvw
LPOgYnR8AD3EV1IZB1InoFgA6JaJzrpC6ZWmE+vaFJ/GKfeBWRvPN0poh/TvS74y
VOCwH5qOXdE16UgQ41EIU4YrcA0LnA+/gCAZvqRsa8XEi7DnctJYSbR6illVgKRd
4aMKyZYYGmkYSyts+r/PfmgWr0WVpZsJBCqI9tElU7TcoddWyHW8/yORlB2xdYRy
91SfQCSlOWT5zHaKOpAHdx3DIOjsUAMJiU+bzw44GOJhAF412g8izNh/n401eoe2
ejEpLofwc+B8SUNZL0uLh0u8bF++yezV4zM0pGb3VD0wrzqLv6xLf+EsovRFdDl+
oETjwLpduxGEXM0eLbPUw7WbbgFg/0D4oDcINBQuKnKKFowPnhbdyiQQH3qIGkhu
GJhh3HtluUaGn26baCmWFd0c3eKwCVMV+uJ7QxKhTF/Ea0W8gmO4tLm0oZyVjPby
JRr9AUhW4JHHo0qwoK7lYuhtGKKCI1fFw10GV3q0nAcnBT4e+TqYGg7LDSA59+zy
hjvE8MXTeimOD4dphnDP2AYQ17IDljjK3Wbw7Ab0xZmoTjglCwDDfm9Fzk7d+AX5
63uVe8uo4B1UV2Ma6/6Ixpz5mwQq+rpnfsPwZOezKdPLRr0qIzfHgsTy+u8hEJdP
kgXj2qpBRLaxTlMT4+JyJFwqIFrQSwtkVoYdCTbxNUpgTh2NdcSAE+S6pkSTDjho
+3jLDuB3uGhmwj8be14Y4WBC959oH0wLKBkkmt+oJMB3OVkJ9GS+9UFZCv8+AmO3
TSvQQC5R21pqsU8qfOmdziiEBRo1IUh0ZoKop3dRnopyogzQ+WaYk+7kQC3L/T/F
9bWdGXHSmNi+9lgBuGr559QzLKHgodPEk6I6Bp/WJwK4Ou2MQ2bQQT3QpXwpxvI0
kkEt/Qp4FGOlola/4T/4PLcIICb9NZzBdiKTr1GZueJsrGYGDGYg5wTZOuBQhLS5
v2IvWGL3Uh8C7D0Er1V3bTxvlkjwnZvxspXNfxgWOKDcrXDxxbHYJaRf/oIEhFdM
LMa3Jvxp+bu7hWgC2XQ3zLfw/4t9stNy3UD0A320GBDxCJpilfHaWAjJY7fuZmrP
hK2KnBC4/cOxfq+s6DfHR7KzARW8KIuNxnmq3b5/36eE67n7ziAH8uijdB+292YW
E3UIXKa7UHhLf5YHC2qRD9aCo5HZzLx2KD7v5yY7R2+KWH/ujVRYaHebIF4j+QIZ
1YyNOv/I7GtnTxgFEgZLRq5ENUs2co0EyVvepGJ4LKRp6Sapi4oBB0YfxJnKwXEe
Gg0Pnva3xPe+Pof54J2Aq9DpZcalRkBlvO1pVL10YZvm3P4rFoQ4RkJHuaWBO9xe
rpD6PA4SOPXvMrLka8374iZYE5hPKRzSaHAan1agqviXl7qSC4fTPWQcWAxdPr8T
UdN7P+SRLJLT4Nvl+CSJnWJUdF7J2nWAdtgTNoVZ13A2PTSiLMHgYSjN9wtXUQPq
y0s1kq/nxU/VtVFeStnkOw0u0WS/cLPWY10SUGlBsyNyPF3gstbx/m31Mov7krCH
9aBEVHVraa0JNEeOxIHUmZ8gnAGoRkmEqJZyXTyKDfQbYiSmCBxWFIVfw9409pGJ
3YF3SJYnDTWIjPDqKyoloEixivoS4p/ViJtI2HjBpXhZ+r+PzrX8GV2uHCvxhto5
NdPe3bPvLBEG+3BpIpivs7IJRFtNjm6H8EUhOfu94Zd4hsbVqVshOs4iHb5FGLi8
FyVwYQZuBP8MqNHA/fzbslGVtynRyeYcF5MIQKm3cQ9v1w60APdPe09o9aBoEU2Y
bq3tM8ED7u6UpNToMjxGu/zFy3UBzp1ullsxkr4vogaHz6WKqjjIiYMQRhjcKX5W
u2HwTrgagr5yChpdYMqbvTXgaE9S+bhpze+LNMv9E3EoNtw8crQWQuYPo6JvvRxB
nNKIDgJdpvk7nG8fjb3orf46a0x3HCr9Tvk4RXa49OvbEX4zrOqLsSOqgCYCa4VE
HzeoTZo3gxTTAMlVnMDC4gOSV4td6zlM7mnfr+6Vx+MlW/POXxLK3YfEzYyx9051
LOmy8zdmk1LtUqmRyJwOGOTIAzoRUcs04DKoRGkJj9WVhE+b2KaOpuTYABQiDIDk
Kxq+icpSFYZPdhhRjMWqPYz7pOWNa7ipmGK4Al8/FKiElsvb7gGQWdzIsV4+nOcO
uJ7Pqj0+xhXbuX5BuK0jayGuuvPBgfhslz4IKtAwHDLE4wKOMn9UhStWvdmzpa72
unkhzbdHPaJNXcTQnfwmILo6fxpcLFTBDVyN+pktMfjKwAGkOr9acR/3asCSOOJJ
Brx7u25qgQRNtUJLsCvNR9wdPmHrnelo82vTay4Vtk3d3/h9rDORUxxvmDRyK59f
zbZkV8NNnYaSPR9s8ibe51MqTGj+B4dxIePdAsGrY17rNGrWtVGuEZx9PqUjjbBW
PEE+vmig4JtLJaX5iQ/N5MtlnxiO+/PM7a3JH5EuTjO9EPDUGRSx3yLHAzKhkDh1
z/U5ugGciBA1Ki5n397c4K0FylLe3VEgbN+NdagPkCap/Yiakn7667mY1Oy0CFPK
+FVxgApWCCwYzFskMY1svuT4Up3UZeKcbwn+MtDNnAOvAG7IRBddYAQrxpPdygwa
kPVnSM1YMzg3WJKR1W9gkwiXmZB0J0x2tIiRIUuNmoQi6p+siUbhUhLqyEp1oNeM
Tx8BhMdZMaLbGi4IJEAGz71kyvEiouXBiiVAXd0IjyLB+Gq/f+w/5zURfYcOmxFO
0ycTN6Ano0bWrNuxuXDw1MmDvyLAplTVGEMGuthVrSyqOUcrQFoL5g1xkKMVkrJk
AV6HVZkJmE9CNl17ucN3xMZnkqU/69eX0zvEw2BVpbhD9HXQMM6YINCTBzhlzCmi
hy40lGsFfc5FWL+v3c/XbBC9qUwAa64UgVMyDqt91fxq08pVBIUo8BMbVtJeBaD4
bbD0N5rbaGfT8A+4SjZ4DdwMB8jZX25ZiVHkPgPHxYnO7AvV2QAAp+V2yrKdqLRI
FT0gKEvbdqyNBBC8xsMwfuMv3OnwQuNqrjMfIz0HrR3DmMqMKLCH3hvbSHH1aGv4
GQjsYHVYcMHTC/eTijV4mZY+PocNlKS4yxZkF//v00Yq9jlcLNuItiOc/d4Bd0qX
HBFcA8QLfm/dw2Sk7ruakY0RE9yQoojsrR9XL75s/8iHvYgLroj5vsHBNZTTp2kk
+1V5NkJkEbiDa0L/+QxFsycXRLUO/IhxZN5fgp5n28tLTjvFuf+NsQ7TL1yBjL2l
zSJq50Nm4gCba1eGtVk6jLKdPvAyDvapsZ+97hYnvd/2sJ3aylJOZIuB8m+ooG5a
GV+i2HjB3ftduD/ywn4xIbP1RiIjt8h0q+A5ZEas9OcHGfcABXvykelzwUUIuTYj
cPFMJGgt+/XRCpf3ZgIpHz9nYxYpZa+vIJkv1vir0g1UP0qsL2+Oepr+0ar0Buul
XBXozcFcwBpO/yQq9GFTdkud+YayHFKuBUHRq5Z/EliEhX2j2eVluKl3BOGtfMLF
ZyElvGZZARuv7zW4rL89nRZVkWmRSdzLQV4zxO6h3gBN/+jWBVbHKnW4RRUjM5ku
nPgPjr69mYcEwGyEszgn+KnziVD2GoSTJL1QQHpZbaUMYriXite/5McMSWfScUec
za6dD99YU5l71O8kUJ/qze5aYLGsigTL9TsNam52FqkEtWXDYHBYN37ELOGCw1Up
xIgA4Cj6NNEBRAx1xV0I/qA8IpKXo0YAwX+ozoTMRAnQcGObZRZKvSZDCFbFKFNf
dhHKE6+9QW9dbG64eSQpBaPUlMiY/CtEc3V+FwHZi9ISEOMMMSW8ZyewNSAlDdc6
Kf6/bYPRH4tZlcMSJs992DTDyLe6Kl7uE+zCYC6PeCuFFBktboOE9NH7lGsFqLN1
wmmVEVaDQ5VkGg14HGKHkJzdg7hfIHeBVAeD2r+RdEF+wjIQtlJkmnl1zM6/iqzA
YdvgckXIsQRV2J72iUhKYeCg22/LK4z6bLvqUUa/MMt9CQXKu1rmG7tepnxBkPJ8
q2v4UGLtNE3Up1pa7rIWmyYLV9Sk6euKp9NCCrukLPpHcL0dZQ0jLKkruPScNav4
cjbrYykUAtQbdCudk2KqnBLHFe5CsUaFPSGNOHBTD0sO7f/eNGfRby9GIXs784o5
QizHX9bUHEigYJg/GcVXE/wNy87E6y9ZHQ1krE0AKMzTaYt/WtYHhn6m3CUcZmtP
dXohpQbhLt8osmzRUw6Rp5pZsYhp+p1eafmJqRxlfqsiUeHvd4ipvxOykY70UCQ4
gbC+SOd+3AAOac2zQl+J8eCq+IcmjI5xAXD3nrkyKeJxejXIIiFj8mp3WNmwb0pE
/Tdu4Fi5es1kw22zG5A02xzO2P32bbfaIcYr91KpjMGisvPIRmYkAROG/jslRATf
M17PYDjLXKp50xliFx58I4NLtAjImP/N3qyFOdUJz5z1MgJ8lBgn+GLQA0N0NqQV
DG5KVv+wOUJDk8nqW3YSpL/TrdlYHF9hv+7kJIear8JxcoV+eysxgzR60Xsy+f4z
eWTvziDka6nGCJxKsjDHovWGGw3b6Q++6NQDWsKXiN0pepGOQqc7ag0bMH8pVZih
NwoQoOYF9oPz2PfvYhMB0lJgp5wYyeNzNCXoFJWWArUSObHzhfxACy6xm5iqeRq+
CvO9qjPLW9+ozFM8OdfgvG8uOOX97oGI8YU8wUOZYG3m84h4oCOvBa8YAob0MhXt
1kk/BihXOFnJmd/X+b9xW0OaVceRePeYvepyhwraDW9jloPrJjHq3kmLCegQ1eh0
WDSZDMPgnW4eMqpG41dU0YEIPuj7gLBn/QlIj/uqpBIebQUkzZCLkdiIBVMUQGEN
RIseIvf6Rayej+8WcCgGOhbXNVTkqZY7R1rofBb0tY1jtDXDBCrQG6tgKepVEBMS
VehFd3S1BVxssD8qU/R80Db3stGei+oml7GmxxzT6lNI5YqhExlHdYsGie7iGaj9
lEKR/DYgZOMwOSRKPSOk6yA6AEAn1MhdOf6zjM1l1lemR8d8yW7PAu2LS3oKn0Zu
Bgmplr7xSf9e+1forbVHrpj+QsGjrthXLRP/wvUht9wUV18MxJkjaGDOcgliOkGK
+L+bjmgVYGuSZFOhUyf9a0CJb5GhKLMOXJByNagYzmi1Nhl0gepiHfW4AC4GzrPd
nVqNPyKMzPvJZ1O0+x/ImqWnSX4muIR+/0Jxls7tOBTR12BfUxe5TV9dvYtqyh2t
2RhVV58BjgbFzFJ3ZFnAGXpXQF0eYnpC1jbY7GsSRwhJM9Y+Huv1NypDm5SiFFBg
5uOj4LH4a/5yxDlQB9MolkydtNWtFAP87UfOaLHdDnyDQGJT7oeGYVv0Fv1tasRy
eNHd9W9TErI27wevAUB229CdoYXkGsMZHNEWlRMtd8oWnRnQh1kr8wMZjSJI+W6a
f2mjYQEFDVixz1EtLNhvjtcPytkO/Z3np0or4v6eUZzOxwxQTRb4T1fHnfnSZUff
L+icDOVxK7z6NPNE64dR3KiknyVIRfB4ZGdefHeRfbgqKgO/G8v81jriUqQ74Kk7
5xnbgYED88nbV1M1GOIsaK0vdqPCYsPiCIqlMdw4S6zX1Do8EqP4lZVZATc5LzlL
TjSCc0vTGG9IPoFmsBNpkY9a3BBx4hvBu+Zl05tpuWpVTef1ptTTRmevDuaqx5rq
IZZ4Hn2ZxRfwXruz4BuBn7vL1bvIScCuLym1i1QfbvsLeFB7GvIXQ67NyHVdNKoj
yTf+TAFR/iyNVrZkjC2Ngmznhlup8R4yOlS7yBM5whJ/rXMrJx7r9K5/3K5I/22T
4MqIm3AezH+z9lD8oXpfs6n8+W9n/vXEIt7HAtbNneBFvkW46TbxCg1SqhIAl+aY
iWJB9YEgPRL7yF52oxC/kxZ+U/qU5V55KOOo8OHInQFgDj829N/viYqzQgooDUa6
YJTkECdEnTdS7cHlQhEsCyVD8s7IoBGVyIWcepisv6XXxal0dSip24oC3AHbtbga
SSGrFs2dWTWK8M74u8nFCF5aVFYbJIa+V9QHz2655pk6fO593UAM2duL6d83NN32
qCXHBB8zcabhRRLSsIscGlHKYdCY2zMRNOgvjUUmrdOxP1v932ePlyzMeXR4O41+
Ykhpz8C669J4ZHk0IMUg2vvdjLjg/CI390T2sbSjOb/P5at9YXINSffNkaDLUqsN
jBin5BeD8leeE2aQFUU32OYYSXf1jV0ft7JinYGuMf9BBqf2LqOA9DlrC7tR62z1
rPK6XndUQ5m51CHbCUgAjMaWAaCj3GwyJqsaq3fM3EJSaKeaE8D+IWySyW4c95+e
r0Otxb2G5H6r8n6JP0UyYJeYQwp2vY1UJmkVWHelvJU6CF1jqTn0OghR+nMbXHug
IjrOkYlbnke3JXc1EUFiKtk/NN/e8+cA2fg5nVeEqpv/dfYgb+MHKik8mSpoESTq
G8pjqhls8F2Bhow3eziwyr5JVw6J8fOUBQfU+mhNwq8adnTAOe/5LqmNmDw6w2JU
eQqgV7F8fVtH+iJFGBXWCriPquG8+W1xxxft/XWu24Z40u0ScyIBcRrCAQFvICRk
VyAWgKRulAeIPI5BcIuBK4Swcvo6JMPr6t1JZ+MUqJSUQF/gsE7yy/M8NFjk1HQ3
3fvu9shXxsVb2wgWfJXuxUeYUHyBkozlf9Ani2BCM3UVL0ri8i9pzS8JjL5/vyb3
dkUCj2q5w3xCksQs7ezcTuCOorMrt0l1hp9fNnfAHIs/gSjHCQx1mUglaCQ8Cgwh
lt8Jf4DSXT90DsBzMPvxL62Jvb5ACzGPtHoyGqUNuCuZeUUZeTCD3EKBixjCd/K6
4b0kTigHhCUo5ZTf27a4RWNUIVHl27orENg9Ycu8fFD1Soe0RaW/+5YIZZxa4Del
CVelQwqHDbzXvPdqXzCT4wg/+uxQ3I/bA/PvbK++LY33H1FeJkMw/IVeqKEWtRGj
IOcdfprD9AsofU33HdT6sbgsUBvULwecZC7YUX2ubzBKc316dE3P1jsBS4j0ykgC
ju7ReTJxqN0anUg5ZYdNkweXfBWt1UP58fWw9/Fvpn7TNwTRfvqNN2M29nXsqHRT
5qXQM9c6ALRtppEMJLND8xGB34wRIF3YgLZWTYXYNLRE8ViBANg/J2CZ8O8Io7vo
794noNMDN9MsZMsYo5DjdfuliWiqmwSPoc3CnmXHB0iwr1bRaPcQOWv8fxxyK1Xb
wLt49vzkSPKq6Do89ZJwdR7T5CG2grrkKfqlb7mOV9rzWA06snLACi8j6mhDnDyY
Pl7kSBTfbevvbtdvB3Y0Mesr5I+jLBDlLxJLTVbqSna6XssQActY9olxwY12FiSc
aPN2b4S9I+aFsRHOiotHlfmjosSoOe2k2XUlg+TRGeA5cIBV8iVK05FvIrgYXcQ5
7hL0L2Y+VL73EgyJ/LfjwlHK6IEbNxzp8aiZ5d5wpiY5l9AdzYHC0L0hbc/MXXWf
S7PBXIjXsoAs2FVL4XSfdyaj3cC15jqxfeIIgKpg2BvWc+Y71+ooj2MDLAPFW86Q
Tx/rRMLlTJs2jzNSnCzaP5vFb4qBHYPwuNHowBGzSDc03TydP2SOmzk6Ot4uU3Iu
C8SoiRHgyAJtd+OOpz5egtYNia8WPlXhk0Tv+Qnpqu4Z91rc1Ufb2VYUtmhgL76v
UhZgmeJZA5bcR4yl4YFRzev5Zh+gipBNftCcidHvdaioORkpQ3u/zhYsUrv2zBK8
suV4mmCQPOitIyusNjXOL7gcpsniCZQkQnRMEhk6yi3qvaP93VbWirDafgCvHytp
0FZAPKiSmNoun1sKj4YNLZxgBykQD+kwImQy94SieA10orJiMUou5at18Tsw1JEC
J4zJ0TzGJx33YbCk3/dPSqBG2cBZ2FKuPbSX6WWJZFiYbjYnDIc6SiDr2I8+hkSH
Ap5uZvPz3vOlRnfTs6OScGrqqtlrYLVTHDn28iC6uuL4QI2TAN0p6m4MFqufH2WS
1juFiL20rjBJw/jaYyGvfalqUuIAGCwAGUDwuGxogPbJ3pFFDInuXdOKKjlUBHd1
7oQJo16HSo2Tak9P1pF35qEHCt2AftjnK/G+GpDMpKmx7K2O5JEoRsOhgq54EhYM
jKQ1TzEotk8zQakx8cA8zOTdom0BCOyj++NZsbpmIy93F6LjFUcTlkxz+0K/EmGY
rpH0X/CSlQFrv24f+4i8G0JyVqB8L0JiahJlGrtGZWRTb4efxn5SfltLiVHJZ4Du
Ubes2w6Ip+XOfcQmFCIbyG4ohAmskaJ6yQLejrK6H3LaziFeNeLfwsaZakx+hABb
U2Gx4O+dUFN/At3LgxWUP4yNtsIcJDwUBzF6kp9I2Q6q2e6njdM09Zoo3cJOdfiY
JKDlNWWS9PKnP0BP3sPDhh9lbf6O7wNtm96wrbafHct2I4PvCCDEHkk+R8Ys5kdp
RkoeCBSOxbgZzxdbMmnHxnT8V+OuSkB8tLSQXSv5Tjw10Oq9PttbOfJ62vrh9hEV
8WZBL2yFwsC/LsFjD6N3My4vbcLonRNuYarAGLQhg788ihiCcTwYjbAH0hNmEP2O
f0lVZaHfTyQeEKwSUHnGc7OLFfNgHqJt73joeHNxY5n9z84f6PERqOWnbVrolY4Z
gQjztoMsRjNMOdVcX+prBaAzK25aX+mQH05AdtI6PWOJFEow7dfItZd++kg0osvy
pV9PsDjBDXiL9ai1P591CGXQSPLZ8ODN4RKrzAkbWAAeyA3fWLMZnhWD9osiTudM
tOrwNl60Pqk8ZA5nqxRMyDeHxgl0zafw1WyVSb1JCEvVP0pz3onMW2mMZS9LaWIB
9q3IN1BpTYSda5uFZwUfGJUVprUv4C3Ts3UmZSFyZtLbMBS1/itl9r0OZYTliJqH
pY/3UeyWlkeWYAduqL6JtxR5MlE7d8dnc9v3TV/SeBXF27KD878RUETLKGC1AvJC
RuxqQjEbM3ATDp/Hp6zcJ1XeWZsB22CHDpZOnDoaDfUdosKv1a3IB9ufxJKnjoQW
uRgoNpaZ+6nCp6s5kDeQOQoBY6eHnFrEvMWnfYcqsu3ysAGbbLVcidnZkbPhREMy
cZrPy7EjO/fo4ATgKUBR2Ouc+t5hHtfFanWA2CmAOGTNNUKRieZ0n4kwnc20Gl6E
fjvv/8YFqmGM4Ylx2vY1U96axa9ActboLY5ELNc0uLNPS7DAS9ul1MdxOJsLmlgK
nl5pqDtJjm+d3zB/t3zkJ8zvr05McoKqvrnABGh7mzKFfiCe/Hl8czxywJTiF/xQ
vppbsDebaus9hIrUBzwAQHSkI4miOq2Cwrli+B6+HSjTUBaOg1LlT2HhIq9QzKl3
PC3XPRydaXezrCqfkJIGkxSxYGTQ3BDzzOkF/syGKUOiohxz0F9UFdF1bSxLvG0X
XzA0HVeHKkp/InyBhGqZcWwQhv7qGCUM+SnJin2IjcyV+1PHCfXgauPDBAjcsK4Y
jZ/naYC63E2aqTv+VSblTw4nQ2+sOxjqFXm9bFkb7QdK6LxSefQZwmU/GgFL1Gr/
++Ertuu6XrAfRodySGcQ1ZrdwlmB02oq9Fe+BiVpqhKkrsOc/7p2EguhoGns8Y+a
A6EpM6Q/vvNRcwPIIaZJVTKLBR9gpH/WfGT/Q8J8w5PD085OQm8E3a6H6//UXe2l
zNywM2V0ZPG1nS5HqH7x7ET5vVwpy2QwUnLoOYIbiCCrsT0nt1pXtexIVn6PfG8Z
Z1FWdIF9lERvx0sbSSfNUc1YbI1uCiyNnRdxhv49Cn3jTYD+eNR2AM4fQz2KTO6q
5h0PjBGBaR7S/m6/J7beZ0iWC6xta8Y5cwC+JjXkglBFmgKy2tWFtsBrMvCwEzfT
OCjlT6uUGZs/xsxxG3Pu8WWUmIKDhQG857+Th/omnUAyU0C5bZPm1MSg9wSVhAgJ
40FdaW0kuU6fTxqhvdhJddA2rkwr3pjuhZD816t2juni9ONVkA4pVxy4QlkXmgJw
hRY9o2eAwc6oMYytdiY6sE8nFFnyIvlSOv9EUfjFeIcG1L2ZbbxQtpqumFUoDACz
1WORkzvT/HvUQSaxTjSUPW9riM/Wty0UliujcDrwg+9jvhEoZ2h8xNjEK/NNmjr/
3hFxraNLIHmEP7PhNjeoqw2sY1YnkpTCRUIiOHZ++GnhrGZTkwiQieg6HLRNUWvd
TBTsjjgS8D3MIST6FnxhOeAPTm4Epu7PYo5cL/up8qT5dmiwGr/I39WLW4z/B3bn
HnbAv/jURg6j5TeWvXdPC7/2aCR1nk7/fL7Zr0Rs7VZYp7Tcz+AM+BCoK0hX9CmI
m4XIEBhvd1jT0KVPABS72908iY1D2DyXh6jp642NO5zq4H43+vUxaehx3M7Xif/P
VnT+xG/9Vkhed/mnjxQ5QiT27tw+mBDw0RvT0KBNwy22pEyUycKeIPt2Ip9lXNND
9AO7Z2R4olEg80izZXdgjT+i9Wn+O913P3iogSb7ecFLKBoMEgp/impUZ89kjtcG
D4kE8MMybWJvcDM3qX/2gbUhPpc4i139RO4a8h69TuDhMQuG+q5XR5hHVl8KP03E
WRl1KxafMKh9XsrhFOzNNTQIzjRFWcmot6MX8Ymq8WZjeJR1gdgcLzFTWlKBihPV
TezI8uGlo+PQwf+SLbyN8uF97YZN470xtK3WplzAHZMwMaPQQmQSFiIhUbRCClHx
HkiTDwyR/bP9z1QmLpKK24JbDXetAbelIN7ZCxPzHUaV/y+QIvfjw/LKFpMDp0k2
9C2Kk9l9tmCCp3n2XP6Yd+BCmm0ob2S8cq8Rzle4ASpyH5y834ePA+icdCbDVofc
ZVO85DUv/wH/cJVrUDgeqWpCLWrSSu7BxY/1/9MqJJIqaDhtWC8e/PxoJrNQNCeM
0hWf6KqUi6IrBEFaKEco2kssY7IB+MdhXh/uhmgmkdcN+upAxwQZusf2c3Tmc6vG
Tjduy2giGKSI05jShRtyplpxuH4mqV9r+lp8nD0711/0papRiBOyBk3z5lbGdp4J
bEV6+Jje83c8jAAuCHj1AKMh1Oe104JsEBqhYl7Sa4PGzH+b1g44hoTi9v1HY0Vh
9LH4LYsvjKQZJj8DGYiY074UEsmZ7+/Ok4ROSgHNIkwuyaVTyK0s4M+JVDD5FnlU
K+ICV8Z1/fl69y+KxUHjU1+kZNA2uQSsKz6PSZcHckAdEgnGy90r2jAvgLxCo2o5
2rvaH8O7ewTN55q4pWAEOliwiEbmRDFnak7KuWIiKvf/p+eY6lG8UVdS5bQ/ed5Y
X9IsKx7XyRP/bPZYqgmZIWemh01CnV3TG1iVAdMsRHFXntvWcAdbzcIlBB+pT75s
xobGFFkrEfOf9kJPSlMB+YyV0vA4oqG6Ea1Wj8YcM25fSZRr35V1P0SKmP42n09t
xRWDdjwYpSxU/+ocWj7zBqto7Ee7kdiI9XH78nqH1NCdTNpRc0At31V/NRDebcB/
aJv2mLank3OzgpCc25A6plpxGC0VieBvFMJigXFwooEongnNgp8o1766bYDiMTVh
jEX9B8fSa/PGpiRy41KvWiz9AxzP+CartdSgX6YaUHc1WcNZGYkIUqNSb/JgfR+2
W9MbnGMXYT+kd1LFs8EcbZKPwfXyKY/bCJnxrFTR1CrAP2pMct9eusPzyiQqLyKf
0n3vupUu01yEat9Ni+wCHyKTup6DO9pDlAxOGaBR2tHdXeJ6w7U7uu4n9iNk1646
65Y4ZfYjs7BziDqnLBq9QjYqZ0A+Ae9Sjmh+02bg0Zi4DTdOof9iPfzyN27AF4cN
MrHZYsVbqRoUledNa5N6PHdacLXw0XBDmPRps8szAloAazhTrlpwUaGc2kLsL/eA
rN4Nr9y4IFRzEJ8JE/FDBXGoUDJBxpXsPklm7fcfAS+9PNi+8AIcdcLXxcZ7A+45
kmLLjNh9MHDjmrBi7kRQvXGvyGPf7ebLIRfSKVNI4LQsB7wzSjCgAE7YZBFFiG2Q
nmq+bBImtI3BSCFATufgRvS/A75ztE1YmSvXx68mzxlqfGKeoq7hAEPxwcWGA/XX
QGCyjYpLtvGp7i0a8SU9NDATIl9djCLLO6da30ADXRD3zzdQKZHzw1gwSK60Be/e
TbzRX0VY3sGMVYe3KO5jvKYYmwUMTY/DVpfiOZkGlD7ZXzjYGSM74NBOpGEjFGxZ
O9/uHOZnQUyJAn8jfiteBn221GN3cPqXJyUXQQP5ULZp0yD10klXMkCgPzYz319A
ZhhDOEZkz3TEx/R8XpnYUUNZ0OkK2wSKgSp//S81DtDveP1LBFO60ChXEqjDb+yc
Ei//2t91XMTkhU1bgRPK9IZ6qTNJxSz2pNvRIs1blb+vrnczSjb1YKwmNBmoDeC2
`protect END_PROTECTED
