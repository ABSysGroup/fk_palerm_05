`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aLUIGxH85YxnTQXer6/Qw1QH0vW1XH2VuwSlwk8x0w3I6LRgDEcjsd8EIp3J4aw+
E0bQ4DUXoquyYO6kO/KMhXsMZVgpWBeWTe2kEpj3MiezXT96tFD9E1bmIXKxVKaJ
4mwCqGdkiqSfNu7sDXQPjNaHpubZIkkwD7EDyjPpwmCcp+xSznoqHd2LdLtrDKsR
RoFkwBTOGsLKHOMz8Z3ro5ZC5/3iMvxP+gTSZJM9nrLRHcQql+Cpd6vcArxrNnma
8WRE3XxL50jrJuTpGCkNNxnpYv/zBo4dXvivp3dsWwTykNGbOqPcvX6z6BM/3QLN
wdIW6vBG7DtZ20GF0TF68KypoySoui5lth7BM42gSDxFHB3ie9s18VCcIrujc2nw
aG7iAYBz452zkv7rGL5SFigp83vPQgMiEXhAy/Uktrkwg3VNTFIxBOwTtiFN5ujS
AQ9ujVOZr44SE5HFrj+PD0OULl+5RrlIbI6INCqhq/+d95NJlGlz3R4oPHw5Osyt
iIhq97FDeHKVzDyNt6brB+txtRyhkoteQLsDZYnx6azdZEgTitR1P9Clc6lSTX3I
sZa1O765MskstkuDDXYgSdsgPocp55xGwuExuIKhz7l+EaPMgRxj3bLQleNXkcML
x7tRdgC6hmfwm9lsxTFh4nM3WNttggfoQD9Lb4o9X8VArLw2lQkDLDnFzp8r8SI/
/WtN9cbZl6O8lJNKZMV6Tbkqsr04HDg0l+QbcbbfJGl4AILkq7o42H+YjfB3dCmZ
3l3T34UuLXApB6qoXRcxlA1YyiEgZPLEiqJq2dLCtzaEzcAFaMaMBdX3Vbz3jpkK
Vb2ruqeX/8ZcEUZZVKoTurUflqcXLPrXWMF5x75fexb3NvnmWU+S85a4I2+K8+29
uRnQbZz2yko1RYOWYsx46xVHkb3sECnJ2+LKfwGLec7JolHKKtMNyGQuwyBGbll6
jyRe63cVdZP6YpfMagf3Xh0Mef03DnSxwio0NLuPFNHkwtQYzh4+6oyqBxCDugpl
zom6DjodgEN28V92EOTZbVqXVDq9EFg9r/bnTTYuG1ywwKtN2ldxL+2c49eyDWUb
yDqLICcnjJW9uoYO+snsVxByf6KVwk216bV31DxFOw3etdRHCChYlw/I60F+NUHS
e8BR575yDhwKfqTU2puII/e9NPyKJtg5EhzXLm+L42P53LyqORbbsChbk71dL861
FWDD4JTsy1WhxEkxhZFhOSpNAucr/svyYm2zaW9QD9+ddoc7nquukrm6vbTuNryb
apuWxhHQ4X/5QcEW2701JQ/arsPjYou1VVP9QVBl1/X4iYiDy8jrt/COVoNIxWIs
nxmC7tQZfZVr+P6nSB+z4y3wZcvZJV/1OJtayYqHC5HUDeC4bnqCvnHeEi+tP+Zg
hZ9e4b0Uy3uQ0SHFzhIMrozx6+7weLvQ/ic2Lw1tGAKloIOCNk0zKCKdJPiXxjgl
RUfsJ12yOZjkuWlJ1S8FzQg2p9ldXmt5SidD/2S7kQKX1mEIRLLQxjtAsYmlb7AN
DreCrBk6RKdzcWh0L1ItHGjvd4qFf0BcrmApsMvyri6x2smcLNktblJNTWDuBVLg
sq0PCjPXuc1/IUfruGPJWOuH6qvbzmvTKW4bQbUkEewX5Lj7Qd6DH+rwk6j0fmsD
ugPrR5/gqARtfWCEI2Rtvs51CAie8FbDwuOBefx0cWIIKxQahWaxQfzAOa22jXdi
Uw1mSzAm6/lqMSaceijRHRzj1Mm2o11DR0fguw1t3SGL8rc4TN7ICJlVhmBCDJz4
kPu4J+4M1gNFnswoSbT1adK74WE5Fohkd0VRZ81SCja8SyozpX7b3I5flud1fX8N
lhWxNRducgzkmYEjA1jUH+Ad7dffYXMV0mMy7aE4kEItCmq69PS4LF/xn34U910V
NRTRBT1846zi45HvFgVvu+GN5NyVKQ42aoSxPw1Xivqu6wI/q2Vf9t5G2nuaUkBO
HDXDZ71duJ9J5RFVExkH8RR8NM8qK4VSqfqibIR7+sWl6ecMdxVntFCCmI/mkeiY
q9c08a29Q+CqRLwO+a5lUvxBrdY5SF1Fa5ViAeex2EeiIpGtQNVnKFgZ6Xu/mn9G
QcXdapLY9Fi3rMOi0UJwYhAHdRpPRpLD/NTK8DJwXfazLkpzF7WILvPeFfARc1rt
O1shXQRaQ6dzoyTDLoVRPdr8doBQr7bN9/5UqHYrpdOUuueEz7EQIrEdnDKUSnx1
lbgfmZeLaAjRvWauxQGIIGo0hhVnciS49DNTjxDStTUFk8JslqSkIoA8hhl5N4+x
V8dSEDjr7cmjma1yeZsqDveJ3N/Q8F6lXXHMRJe2110FdkXOmgt/8fzPUtwjALcG
3bWiT6+0dXerGoc6HKwjgIIXA0ygZFqQIVfxFFBfUqVrVzjTJ3VaZQkwmQntgZUd
hnD1PlV1Ym6bqmUPinwnpZGsoj5EA9bt6ng6dyGOmT/t/WpfTNjS0QRKoLr5FVjd
0933ble9Hm2vnwKRiGH2jsCHRsFtlWclSMIqJFUnfb4=
`protect END_PROTECTED
