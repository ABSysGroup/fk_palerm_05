`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RdJSsib/8tmCghe2RFtLNe5dLbrq1d0q1+rmpqgXLjFlcbpKDnhBQqKbIh697wiD
yLbEmzNuAN3PZWnXSZtn9Yl6Hn3SeuuQf5xUDObsOsp1q/lP1p9uRe0eC9+XgmYO
xF1dhZQpx2fSDIEOIebKF4tJc8RK5NZC526JaYCYdZHsRm4ibMF35t1e4tvlht5g
lGAeafJTc+ELM93X6EJG6+kZZ2ebHSd+WktfHBIl6VxVnCYtvU3GFBd6N+CB+vSf
sSbJpTB8lYkIvYS7cjK7O0/Pe4QhrA9CPWy2rCT0cS4=
`protect END_PROTECTED
