`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
06E+ywoTc/dcbtie3CQHqqaZNoKaNtd0sSELDUUHfF48gSQCYyYJS5jxgxUs89Tv
u2l7+EIuSphPHwEj4KXF+Ai2Lss3Wem4SNo3zes2wWFEVEerhlMbGZpZNBB7YYvt
NpxMDRPiWbKdFYnk/4YUcvIc3KkWPWQEm35A/P0kHQhTpCP23sQaGFNB6LdERPtR
RvRiLNs/kEj7pWUdllmqPRaHC5PMnJ09U6LgrGVG21RR9+6JE3dteBfNlW6iCqo7
EZAreFFqIld5sGF4ipNDUF3Ip9FLikU2u7ZNFNgo0iaJwqpukFINDCjmgWFnb2uT
DuGL8yfKWasj/m1LCc1ODDQRdJXogn6YEBGpjeOStGaoumoUlwQbwrCL/yyCGGIx
1JQRMIy6Q57fZi0kCj7nlmPlYAAVvRhE7mwWaOzWCYDb5Xec9rpACuBfgYLeMbRh
yeuHzjAln1l1263je2ZaPqGkzNOdokSetllBZhCDHQI0MJu8j3bcd9X0GMIQwhNC
jTMne37ePQAj4BfdIiC/dYXE/FfFJKK0mvRE4sPSCSHNDWNsQrL6DdeepJXNrhjh
5jq74to8WExqGpQdnz0Xlrc5OjL68lCBDHSKnTAxqi6uNXj/W/3Gfjl8vjhm6vln
nPBwgsTqLIRa9WPSUqcj8lXeqVGCU0fyrrTc8dN3IccD2+0V2TtvvIynrScKn7M4
SUxhD2hiYcaKlJctcUKhWGGT6nz/QWTYn7vK6oBF2VxWNtjtInm27po/FujNzDQ3
8N0XOrZtY5DKHsnj/1ebb4k2+wHX7rrQaVq/DS7tLckxJHgq17hbV9D2s3jpdwhV
onhy098xoPxaMNgJZ/Y4/h24S22+McqBWVN3zwcUJfRexF38qOaPYOPKOlVLaOK3
IfwOFKFqNtFSlcd8/DbF5BqFV/rObWKWtKZowIMp2+2CIbgJNL2of01sWLs/N5+T
wofvRG5jV181IwT4x+jheOglUIcCbIdUXx7zdaKRz0D5FUM52+cOVQbiI2EhTPFA
57zWi/z7E8Sj+/mU4WwkEcfOX99oiJVanWTCBFVE6aL0piDVI8wCe/6aBkY/wn+e
3zL3o9MhSqlDt1qY+9IOo/qlIRY7l+V+9MKn6GG/qmhb4L+YfvuAsA+Ff7JfXSZv
PlCxi/tMO02cuh67jzRjGaKMYGzAY724p7bNuhngw4HZhMef+Bu30Aw+O508aYxU
ZXPb/GPPtEc9zoF3y2f0Sv1swoXE1MIXQIm+g02V2oq/k1xdBn4RBhOs25zqgLQn
IBiCbRmJdWgRlm7cRCdFbJXSV97bSsM5SUD1fBL4mxDC3g4MzQslYz9i/ognRvaH
eATs9aBZN5C4eEt1aGb9sCVR4rRRav/S4YcqiWU984EbfOcCGNXnzNwYD7Piax3d
e4UbzXqTz5hmrPTXJ7al2995mNymgiIIhd9b4GG360eXRSDvdIkgtkqCnZY6sf1u
apgwiN/JBFk26DV4Aaocz2FdnYtGIaBigDaP3tJU9z8ff8lab2hOm9z2HDDEvbCA
xm5fEqKVucmdpHpIfzHZBKEtKBsdAFNGwu1uSCNDsiqrJ8MLIHiaCCLEow8dpR8C
bnBSaHi+WF3mLyxXahe1fvCp0IBCjbSz5pMMnRaZ5ZgqVh0LccqE7r6YZ6+vauRy
k21i5saKJC8wKKqrMfDlP+NVgVy+/JY7TFZH9L0z/SRXcHDC+Qf0zWM2TUz8rV6i
/qAkPY9IX/v+2yQRvtpUTPlkz1Xc7gf2U4YbWAGk2MsV0ht3Xt3YY8p2B5RzJGk8
cJy+GkHW3RNriy69DGvNg5xZYpgNMz5P9zzQYa7fQ9DPbM82zGyQ6mU9zA9cAZD2
Z8fdT+LpMsw2KK+4tuKjMu7OzmPQ9eTGaGlAy9Nly7NicYdbIKk5W1ht+LDLO5Yc
X0wcMliKrfl9DBnyJdbQ9F/KNDtVQQ7ZBVi9EfIZ62MpSoJsWBcn37P7q0QrXR4A
EAuIJA73lmT3ja7R969KsHu1WK7DXWtAOe1nQRsLnMEVgdJBBGtxh1pQIIADbFSU
s0RV4MSIXS18xdy8tFRSAiB6JDBfA+saV6Je027paFvvTx44zWohCfd4VfC97I45
+JjB8ozcLFXBHr2qXXSae+fYN6QkOjAw/8pPnS16gPc=
`protect END_PROTECTED
