`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yIJvaEzgQaDHYUBFbzaqGO2rn8QWqxPsEWTHSvOcbCRR52rviQYxmnFrCX1Y5OJS
yWhUuhNu69QUFWdtVuugi8SFvDAD8CNgQmcSHbXJFU8mWLH0zyi5zUSmM42hKmAo
sUht5T8tirqo5nPcKo90LoJg1hpTjQthlzoOPc/Mr6V5IL/C8ggZNYJBH3UPHuSb
SBZ1AVqsU3mrE2pYRQwHX0XHHrRKI5B1YG8rGvRY36++joPjHIS9Hg6QVBqFPuGk
66pbtswvplvNqLntFgN07tAecWMJ12rGNDofsdt9E99cPjel3WAq0Mpd7/WkdprZ
9TGAZFXwHkOX+LGBZzcTpOxVuL12QgsrpDvYPLoWslEIlRT8BBdopscuzSzjJNMw
tm8iVVRCJceRBkoix4tTywg5GMM9s7XNrjTlasDQrkfXpC/jax6gS75WXbrjM+JQ
rJrV517dRe54xnplxOihq9ThzAx6fJwfooTPH1XOQHdBP4TUdDtrq5ke0aV+b2zw
4nlR+VumbJVsbN0NRzk6wd+M3x1gFJxfIPwTzqVamQ/VvGUw2vjr4OqpHpWEchJv
S2W9rrg/wyjruguuOzgZwjGje1/QmpOcjuCueGBiuq/Nu3/zjyRzGtrCsAc1/Pr3
pqk4RLO1JAQo8a17A9sYsx1pewnW5o64Xt2aJ3m4cYEjZXEsXNF7NYI+vM4bP+Gx
q8nZiJVFVLmSuv76CwCM4+66funoNIsNO4xiaVqsQppcAxUvRv03R43qeslCUMcN
xjdZCiuuOsR92Gyhue1lus4iSXKvuYRIBuRA4ofEkgtSLgABbqy8tlDicn7Vp4bt
S0Sccr6I/0BDAhaG7R/3DZiROgNB3ywx7PZAw4t99OMipELrHixR/rgon2Wmeo4J
DUDPtIscDfVw7iFOt794aVctdbeW6mlRy7CiC0Zw4Bd7VuaP1w0ioQ/10OLn+pZ9
TamR8JzEpqibql4ex16Kf6e2R3qfYrMpkVr89By4XSQdHcqshdgCMtUmQtFpZpR/
/RlSIYs7M+sjfy1uA5vTsYfgpBza56v9T974iNA2pR7B8EE56uzNu+HYD1biMaLS
HNvt3U24nFXmzMcZme/mvqsRA4bETZVPBNKBR5SpjQrIHJgt+xqwCWUWR71cG+bl
OMmqRG1e6Bo7Hr9cdJNMJk9uAreX3Lhz84blIMNbRYJNXrz6mn3bp2PRos0i1E3M
wbFvp3sGxbFs8TsqT/tM/frlV5H4eqmbUfmsy9FM6Dmgm2D9EuuE1MbjiKs9QFcf
RGB9guO/Rl/P5FUcXQw+dSO+5VaGAXHDcEKMZzp85DC2iV0BeupQFHYYaSJA/Nf4
QIiZrIuF7v0Skdwu/6sg90h69E4+BDfHcv6F2Gi76C7ZZ8F/CA21kM6HkxMSriNB
VQBW12IAxUsrldhiL7FX241lyn92cz9NwlV6SbLYlvUdhQsfWbM/8+DxhhpG5MRn
mpAeKNEDJRmIboAM5dFpUbblf8RhR0USeo1ZXs1p15nEvDkzDTRrnGUl/pgjwDV8
1HRvZaI3UGOeO3pbN7poOOuFcfGk7tZZWrNy4+PzH+oRpxA8TmhuA+Xr8k/vqtTx
NF8+DpJVllHrL8dCx3Srx2CvOuVR3OgSBG0OWh/2osWqX0FTfDmFjkMEvMXU3J85
KA1WPvjgXO0dYU2iIUVRe7vAIwPMJMjlCWK4XPTY3U5mictRDMW/TUIFmSXf/EC9
3XQZcvTYnnyMJaOa7b0DZov928KrQi6I4zUtPYWpnqILYE+VXsh2iFdHXmjbHMOG
+mBhGDZ40OZrxHIaz7xuV7VC8vsUycmM9SDZS7/jfZs4h8CdMBc3MmSqdHS6gbN/
uVkwIOmz2ghyz1cA105xWVQSUlQ4BBE5VXgqnPrvMJgya4JfifYilyJO07FXCjWG
i4+uryotMkdzIg1BnOOrZdrzmLFy2M17vhSU/SQcckb7rQWg5hKQ7A+DFrz6boe5
v36/i55jwnD8duubnq9ByctVmmpX/EtOd8YPmMdTMF2x8nczWTrOlg43qb4msGOo
cpmI4MMENpLeBm0as2oa2WL2O7mo2ar7M2g+A42RTwTi+XKOpYFySNRLYJzyGDs3
yDkdbHm8DsxFqjIW/u39v/cMyYa8qu7m/dn+aFzdwA/ozV74jgGUES1PBMjAL6v2
9do21F8Nxi1ck7XuIdut5XLmflDpjRUo/MsC3GgixSqFeY7ZxRk6LW5Ia4nxP+3R
VjCwNNl+klgpnlBHMlodATHped14LlbwXCU5mxK9pufbh12gPwo+ICB/sVyeBclt
MEvGGsYp/Tm6FTUcXc1zscKY/QlFBwVzGUi8cteVyp6ijV1lqSV19Puwac3Xgv0U
56/vKWm5fHs62BznMA11062LNcc/FKxYzVidMD8PapnIBTfvdga1kmOG491IIGjY
CwnJwbDbuAUxC0uFdYe4jd0VVD8THOVEbyWKJlJWtRX7kLJjvQrW+keYM7J5ZhX4
wbyKeks0+pjZ1c8px3nMhP1F7J4XO0XAjCT+AMZy/AcvKo2KAg27ieuU7or5ECez
RtrjIas3AG+WnXBrYQoOVgMmKFKwI023Cqd2YS2/Djhrd6x1zc/DSltmBbgkCD8d
Btr42isP5G5T7TWN0ouwhm15PKl7wZGo/8QOjaE7oa+uou7z3iLTqXi9zpn7F+wX
tq+Sd3bxtkoOsrEDiMHMdHI46av9DoCWO3q3cHF6yePwLR/k8Xd+9r+eCZZVLHFJ
DcDKsfj7Nw55pn7c8BJRJuRqpG9d5AXWsn7VMZQfZlMx/IW1VtZJQSPdp7+UGcrr
aC4qbrjoj3uXcHq4UBAy9ofIm1eEgdQ1FYTJX+sMZGI2vSbO6ZLxyXueeZSX48yQ
zO8GcOEdcxDR9Es/TgIzXJ87OeMVKg2H/JGXQhED9kqHag3DM2Wu2SHsig5yWjKy
Ey/WepH1vvEg4ph4on9GlVe0t1r3+QrKOlU1Iv3BKNarXQTsUc0Nje0Xg9Er+aUb
Vggi9u7kyj3RhnxqT3TAh7itYkeReouNL5873EMvob1y7Fk5d4t8gCrXDB0lbxnl
xJwprw8ygPcuugVqXwqiJbNpgIVFlIqrmVa1A4Sj3kFHZgVELREufU1U+5xG1l2d
x9QZNTV32LS3ZKF6qAmGaNXyCQ4xutjqjphRk2kokc4y2qR/zAsuGzR1Beqn5Qux
DmDNh5UXfGC6LV5Rlgc5UMTxiiZE7wT6Wt3Tm5TCZDbDGh9YBiTUfvI6aLiyXzK6
g8PfGUeBq67RJv78sirik9OY/T8pg+bd5BByopwcFv+7DWkwk1SV4/g3z4yFuI1g
E2jZxMrWKLfzmp6G1CuyHCXTspCJ3cRv80vEts9LwM1JX2ZlzPaVJosJ11BPrCOB
NlRsOpnqJi2fQuM53jUXUPFq8urvPjdA/ZAj/5ChJG4sXrFUNkkn/lBVNh0gOTSE
gfIKslYdFa1whaUoZLlh8xPQG5yl3ac1FrTlPNWedus2emRf/5hzRfZ/3OwRB6UF
0X/otb0EE01u073GG8W4NtmeMixf4nUZGlIpJJhlKe2kOXL+wN0K15rpgTfouOP2
4z15V632Rn13gYdGv6/ZTi3zeyxUJoN0etYcljs/EWCB/xN+9ZknOkedDPrPVqG4
K0NMcb787Bbe8C5SLboyZOW7OM3uA0QdBMoVoBK6oHz4XDTRnCn14PGykdqXs4sT
NPYUZJQbRErf/VuuneXY57DO+cRJL3dcNsx8O7snAWVGFVZOV8YSupHoM326troW
pdBKg98NAcb5+75hiGF6WeFVpHiiQQGsRwpogU+Ge4ZM+CJxuCZq2C0o2NVgtSKU
wycSR7iActEKsCADI3vgEoFS3PUnzR/XD1fYZn1zi2vGNbGqf1c8ue10j/Jxqy7q
kAulkXwNG41XGPqXwPVJkBwY7LYVn/23Y3KLkJuHKOe58Wi3OqHcBq5T1ZPK6qZz
ZXefVaWQryPTzEo58emdFEqzvSZy21M9CQzcKeUDwDOgh3RQpWlfL/OW/Mqpt9gF
6pgTL6pLnLz0tXsbmS0U0jilP4E6GcihTU+iUa7KCec6xXHj7uwGCBBif8Ihxx5T
zDN/p95NuIUWdfgfHU3LlC0CYBHVPz1ZWbL6EphObb+l60/VLUeNp8jHRHH8OwB1
FPJWjvxo19biqGchSnR5b7xQrLj3MwOgAJ+gEwIOWSRWBsPKKytjvTISwe1Eus+t
FZ294jEpg6a+hpT3NHl5eEqGR2nnXZKMfQ7BNA4T+xte/8W9TCF3yFaPVEWbQitK
2CSoPVTPgdSHfzmmclax64bjjJQ56gYipUcUdXvDqPLn9GlLGuCB3tKGeeifrpv2
WyMEcx1Bw5sctSyYGTAm+oQfuhCiri7CpYBoYPYzPM0H05bzqvGnXV//PbyFb4S8
faZdj45pecKK1iHEFRtxmDW6++fLEXgI4VOnmtX/+USBmUsT+3Ke35drr/8p0d1M
jOlcHpYySX4tmpCP2KCuIHIGqqk+u+hEHJ61ywEh5fU/Tys1CDsVhHTaXlaGVcs5
Xrb77YT8v7/NF34MRZzSOTa3ST+1aareOBQgboc+v9vjs6h0aIBUojGh5++AIEmS
TrZauo4WfOdLkS4MRjMHuHW1CfR9kPEdyMohTvuhVDstj48fzTtlxaUSUfZg+goS
Po8UAftmSKqCzRWokcbUnArPt/f4C3fRg6bAZoNa/Xis96mpJHXn94SxGV7ghCLe
LfZtjm2YXK84w5Z8JDBUPZVqeJwx9YsUjMyjBqJR45RwXH8OAHl4O7vuwlZm0GLp
SvQnQI+I1KJylVCQKL50a9icy0WMmDtHZZAIXQkP0w6nJpuyzzbB3krlkuRKkUel
S+s62SNYrgpnyVI4APfHnauh/K0qqfbD++YxpM+5Av0QLx66w+5GzNtRbgmXZdJ3
Ci5kChKJbSwCxMN56chEa3tYy/gUek4BhkZZmkvkZNk953vE1qnp3hUd/6RG6XN/
yE9Oc/BgW5AkRkf0Pdy+wX8m2FLJLEosxsCDi0ipKT70xIoNOtV96sCSMnx9qZTr
Ml+/x6F98kpsBhmGyMmCbt/D2gYdgY2DwBb7aF93eVcQUU5xjGB3kbHSphVFoYA9
dGNK5TByUBtAKezSp7giYMxzwD5MHMhYnooRqLrdL6x0nXan0AMk+pO2S7V2UZQo
tkNvqDIG32M7zSMpeGAg3A==
`protect END_PROTECTED
