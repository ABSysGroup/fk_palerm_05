`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h8r8w4sc4N0zEpQZvQ2zmie3CLNm8/bC3JKKOWmGnjwC+o6gWaOiKFuq7WlQrdcI
hL6O3Duqom2dyF1hLXUcovrMHvie4i6rp8RGlmcUI/8bgELPBq8ZZXYna8455rzU
Ax4KrTI23kM5CWTiGMP3Omhz17Wnfe4cu7tbGiawCWlPIMjbllaKPv3l5q20bau/
aMXSkncD0Q4hZQNXZXatc8sRv4pyNt9HoZBhbsILrISOKAAWFKtqo0jX5e8ln9Yu
+oDkOs8l3cXtUya6+jEINv1gkzDt0YUG+sLk/v7yUqHR0ku5pDwtUEg2j1NQ8wyF
NZtVEe5LCObg4SrqC1ygol/sJIMBI9CUHwUeQORqUtjrmiw9GVOZ/6dTphdeOwtG
BvuMJO9Akr4wY3F4ImMSTCxN1nH8134EB/xEoKjhsxJm5d+xEJs1YnWa87VG3+pW
lcy7dTDYM7cmZdaAC01fRYdZqtGlmT4qrwRTo+/cnu/j7YYyRxf4LkBY+gnY5tdM
r0Pji634e57uHdi3qC8JRWSSlekxSdUxc7OKoJ7vlFjpEIkXdsDijM5bWPT88VaL
vOrURbKJ7c2PVLry1ErDcvVE8IM9kC7MQGevR2Sp48OfMeAWZ4Efa3/hR6n8oE8t
ZC/MZDc+xMqA1S6MgUPlqf3rxwQL7wMPgrNhOpcze+Yl+M4QspfbvPYUXXheTM0i
AjGRnTM60VQ578ePniGzDERry0w6S+YI3IOMavyWYmwmf1hY5TFiAFtX30i/jC/3
BFPlLzfCWFXc8CUTmrRl8B0iHjEg+GhU1cdGbAmXmPWaLaaQ3dpDVU1hGWTsbTdk
ACErKVeRojucNBq4YmQ+BhoIsU+WoGzhj5TMFofHvVk5llqQo9i7TBcbCgNcrsIG
F8KyAWOIDb8VoNBD7mPUkhgRxv4rqB3cCSOmJo7l+BhtwudSt9y5dIHz80eyYYdf
4Pi35+qChllkHlJ++cPkxx2ZoHBy2aQNkRs6FusrSMJ4VdI/H+ED/LhDf21yNyD/
kNN7kTyagIwPi/rBgkNRzkaDZn/+yVUz8HxZIop7vo8Q3//upTaZkcJDgnbGzBqH
vnTPovdErS5BzEw1ztlRjSon5H1Nl6OYS6qwRb6pN7BZwaOENQv/Raqd7CRhlQ6x
OdilXAbTFOiQnPIgSj+znjiQ9F3lOKU4XjbfngslBNQyjbijqfzGNBthwYBHDZof
kwdnJtCRt35eqjsB3st1UagJOe5FtlNg3G7sMvLUWYe32pwis7GdzvEVxKZ6XsDh
Gi3JXVecRy718uXVtdqQYVD0I3q4eBEdbtjR1VQr81GuYDdrXxGOS2fykbq22DXp
0K5tBid3atv9A2lfof3htoCVd/U98xPaFMRmDt++YD8onDfSm9MkSUiTvMvOcD+d
HinIk23QhI7BZjhiM2ryhAvknx5Fl6x/ThMfkgNehWWXK+8FbS//fesbV5G00/ds
65lKiF1RSGfiDizNUmIL5L9slHPFrIxCsJmRysesg/3TXmUKSGaPL7NBZxfGGUlH
gAU9/BcMmmaNLIvLNjrk3dwkxG1Htw5AKSNU3V3kstTwkUZLj5gAnVXQDmQn72l9
3wiyREznznv8Ew7tFCxVMlOciOWP37cE+tftk+VuwlfoJH2JLuyI709z9Hxvk3CC
1ljZDOxujMLQBrQ2Wm8+/x+U+tZmkIBxF94yK8Su3ghzLOsLE9u2gmSg4eSLJe2g
XBoi4mgl5Al6dkNIswDCpDJcmca26K2hRSqnw0homueKXlfRCGRZn0eUH6/U6S2O
navha9AIOWFs2CVr/dmha2/VPazUkxV3goXcH5cZ1vhvtW3ivXSu8B+MroTjUJuD
bmJpIDmsaYwm8bEGFx4/hfY8u/LEpLyhyMCB7GxvX6MEZPdWQ2FCe6rB6N4ZN++N
J6Cidkvmd6yd1JeSC95m+5nioVAdkznmg74Janr4YXpLriJXpE63ZvAzdufRq1pg
Al+P9+vE3f+uAfkA2sF9Znka8iIANThfEN31M9Dwf/UuXXLp4N6Orq8x1KIY2wk4
RQkd7VBlApbAz6Z8UUEJ7nJnZyni6BVvsbML5NENAa+I9FdLkg5a+Qy1IbIbrPGL
kVdf9k1qq6TgkdYnaaJg/ArjnwRYhj6jZ9OxSXiNQHFzoBqG4dLxCuyvmrmcL89v
xxso1M+SrvfO9vSXZAb+jFpQe7Fny0SBF6e1UQIkrQNPGtFUJPrNhPFeDEW8BA8J
PM4rA+e/baJSgyagq6JGzNti3XUL3W4jD+kxKCaKglDZsJrJAW1mtS9x8zN3CiYu
TD6e1q+UNPZyBxqUIYEsg7EyXaCY2E4KIbrbMAB+W/IvphLAcAR/9o5Yd7XMFghA
VR7pBHbY/mFzn4pxnWkA8GsQm61TD1TVC3qJfV2WWAKxHhd50oMf58IfEn8vpPXD
4WlDepDLRgpHYgjPxxetLLyEwxiNtNl7G6exYoM5D9ue9qxhDzdQqWR/fjiJEvYa
JHV99UpSA5Dlou5ESUxUjBIoYYvKYNbGsxT7Nyvjqb2/erc4KTFFfZw4CzoXN5eK
bngsRUZRO6IQt2J3jGnkpoqhJRMZRV56Nn4fDIepQWhMSizLkMWCS5/IfXjPtsUa
NSZsazeSZWxwZm1pL8LXRl0/rwc4fqJ934NWamXIagHx3aqWwAc460ZlwRGweUNO
+8SxgsKzIbtQ2Bh0MZNTrMXsX9q6dEUBtBpAiEbwtItQy+w645OULi5GKrwGsEAV
R9VDpIF6psNsS0kNRPafFExsMxU3u89JYZGLuLOXnn2au+6fnWqHXuaoJ+GhQw9T
BNHfJm05p2jL/4wrbU462gI3ceHiMrxS6wfGqJUT+NxmnAaZBjf5jfERXMki9sFA
Xf/rwDj3j7dQp1MT8z8rSNQpauCh4LJHsMdeLQqKKLyvv5OuiHAwT2o0x3jlz1+h
qlDsIYQG9PSmSMSTHP+RPL54swmMiuR1NMYxpIeaW/mMshLrV0P3tchaz3BpFLjz
40Cgqs82mSLdSJyXkTJtKB2AQeNQPXIfeJ/mcWXtKCAxwSn/m4+vb4KpUQZEVehN
zQT5LTOkrbPF2muYLWCFb3nFAqxSUXCxSCbX8f6oWX2XOiqmZcaCdmYbp1YXcvCq
oXqBrglZVj7nI6Pf4f9gUpP9xC4mMVggcKYLx1l4i+Wsue0kAmUJALBkUTbppEtU
Cr1K0kVeEzA1MLNcfC5B5dcRfpfPxZvCADCfnsLXqCsnWSU8zPsgZy+v/FyF49+n
OYfznK0VG5MDRB/vZWZI3Hj2GC7e9t4zAixTx2cAhaeHNVFcL2QWEHr4CsAGvqyh
eye3Y1q2vMd4zifbwud1QupVANs37oYQjA76903eHZ1DUr8nB/vf0BoWnNmb96U5
`protect END_PROTECTED
