`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kZ/nDblz/3vmTy9SCbfq6M6CoY6+37OEd6cS4jbmda8hypIYW7dZh3SIRctxt7VC
sMrELOOUE0TYRxF5c6ElUxtNl6BSw89Vg22D2N+8J3Rf2qGMAw4joo0KD8CAuHFd
SuNLF0WkisCmcnP+SGldeRdkdC3qNytNedIICVQ2Gih505kO/i01ozH65ulc+hQs
VPJBsnrNPJJD/BKJrNfNaXrI4AE/zg2oKp7/tsHXuXF6zAyPJJw733KdszUqcayc
7Z+airF5bRpAqnxEdS9mbw==
`protect END_PROTECTED
