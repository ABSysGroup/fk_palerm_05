`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QcZfRDeIR9YU72Xh2HuaWy4AmSe/Q0bV4+F1irYN1M+5UVCmWCpa+OEXDUDhlJga
kiXyurERVPcjUIEoWXXZfp+Tsrx4QJ0ufvPfN7FAmGJAsIPopQcx6xFoYqWb83n7
HXGkdYNDB50W5kY1eQCkB1G1ypBIz5E5l/Zx2jl3b1wqvAzpXt4iRmOOL2R8OyOq
+V6hX0h0+3AZ5nGDD8wdIp1v1QtbkRSEX3dpojZiz7k5UiOFs6ghzDj9+D/QeWZt
KlpHpbHwBJYcnYmTFY/LSxgipWzEiDwtaNusi8NcxLb6bxSxMNfoOpUwZP1Yrlxp
H7Gb0eO7QaocnnRMYfQbVJnbbpmJT+ESdTSt3P6AUNsuNE2cy12QQiIHo69SR7EB
4m3S+Bx/CEO0hIZ7y+SBcgYtnE9HIBVTBCi5ARdW8sYuaqTljcSwmgRIza+QRJhM
r2Ct9SDV1bh5bO4MY0r8ElOfmIxm0oJ3aahQi8ymTre6CmSi6DBeTI83q0HW3TsT
neaojEiaUETiFIvWmbZVBdARJM4ScJF6+VaTxfmXqCPqYw+nFw18ET4njIQmM156
3pPc6mbMmIVgXs/rQ7NVsc2HbeYkHWSdcJp3+oJFqDPef1YWdxL1tfmq1jnAK0Qz
AJVlLj+rpgYjJRzl3uz8IGmubsGL1nS5NYOPQCRWvQYlyd9V25Ck1Vx2cOfv3AMI
+VlK7cEce8se/LbAJsi0TZKjpxnZEJgcflgVK66m0Bh0dTnKr69lSctUts5QjNzY
EMjXRsI1EuyYl8BPdyyswCFFYpFrBySlQ2EdLpKfvSG6Vfi8L1sz16/gVheNjahE
rj0+ejd6fe5150I9D/FbtFvandP7WdpTcSGRhjKhRwwVaHYqXiQhTRVKtlv+pxx8
nqjre+GSvNpB2lZxs4sKspDi8D6Tj8F3tc7w5r1Z51h1SN5ZX+IbJVapEsPxEuny
LCwTEDf0BR6B05tFMK6xPt5phUUEHDSsbQ8lFi+0qsh/982c4UsNvrx4ruq9MO3R
ysrFaWx+c+GkRbkYagC1qUYyOw1j8Ju7bPRIUh5q9oLvZO+6Bxv/OLVyDsgQDUXI
eThZjQ0pWl/tHQu4Yi3Ga6m2QQ9ccn4M0n7J6RH1SB0ruq+PtOJl2r8r94MghsyQ
klOz+mRwdpRXetcDNFkmL3QLW4VB3fZDLF5f5QUY3Ek8AGfCDJzYYD3jbwj4teDZ
gYNBNuPFyW71nNjty7YURVFCTBNcaT3SJo3Z4i+r1mJvPA0p2kmW9jQfZNWYbnQp
ezcL0ACeVUQeKc+Yy2we7omi08CTMQ5ORPPGUBMLV4xdJNcWMes2ZQMFmwkPsb4u
waEGb37WNdUovF3XW3i8cnKFOgTv+XOgbl28tk03DfedxpX0HnOGu8UGm5/O+KMx
Tg0eEabzwkkBE1Zv/n0qRS16dR/daSYsnvHrX/BkZT3tWe9g5S197KcperLCv/H8
06wH1zhpkD615IuPxb3KvcDN1D8jpiEcllvD+2YMZyewa8iroWm0eebIeRQMW/ac
VZoqiJM1rGmmuP4kLaqsEDwgqUnIUkSy0rPDPlh54c94tL28J45fMM0UMCkUkjLN
X7jJdMg/4qzvDececovDOiG2SU2SWTGa7WqtUIsBdtiafVKdn7YDlsNdJ+Xn6wMb
WMpKqGjDwOjoVdgbtqjHjq4KE/3+0bTJv7bhyHW/dFx8Up9V2JLA+AGpe3Rj40vb
JuKdM70YbUc9jizpWk2A41xYSjDjkXHUVIE6spnc+9olr0fapzEzoKYOJEmTXzuu
xn+v03ukNyXk1H7ibNhQOjatCs+wFwDa1DSIe21QNCqHkzdP+BcAeuBbFiSTzdk+
ufztckQ5tfYQxYaSBZmgcvgLVEx4vmh9uT9hooG67XsvMZ1lJUdJr/UCXJiD/vS0
pWdKXAV8DnxS+OOGYWDVlejTtbAFYo5D2wCkFeB2yNAtTIrquVOsvPIw205tat/l
gkzo+yWXMIIAzaDH+qNNTNiXgqVuxk6ZbB+n5f6F8+RmI7PJ5iO1t1fXkYT7tdTy
5h2e3Ih0052vpOgh0SnFkQl5vSHfS/17Io6Quk0dGRzeNgqlHeD+7y5ONonP4hJ9
sx3CH8dopAGxR9Jk4Y0S/cb8JTWpdIGVZVrk/oyQFXzaDKhwGiqya2Yd2hsc23qA
IJmY21arfPOPlLyOmy5bYiQTKRnwApQJAMuLk0IsajM6REA7HyzVal5QhoCd5JTB
+bQ7X5EVC1j7ZkrLmziSuMPBkHm8vUFG4fV3HBo2huAa+jLjw4jZtomD1l4cx6Gw
AiJo95jtw9DKN3FJHtgM8N3fZu3KDQ3q29oPkzCXKJbRRmtRj9Rm4mGVm2UJ4Qbt
bnrsQqUTwb3h5FN0w9egTyrjxim5QfUQLgf/WEFsGYeVqfIsLFJL/0ug7WFMFxd/
xvwxyHy0fuum4W2XdWnIPhLLE3ukkQYkmhiX6gegzk47CGpflv2fBrENvUIXcpKb
8hxlrKfymTecBHKfw4OgMNqHaD56HgFc+QrEgoilD6nOYGDnbVhXwQyHhSEnLf3u
EihJJm7SjtiVSmi50F2FDuOi7G9TkBkujCHLLUxp8Ot79Y17Z3uFgyo1Aq5hxq9D
Xitl3GA+1xpyGCdbhcsdJNkCff31MdP6VtMXI2yyPr98R+WmNldxFlvvp1BnVrls
EVc3vUVMWw3acmoNIbd0LVveArrZY4tnx0JNiwU1RkT4laGUuvqQmkv+it7QWP+A
6dlYMpkN2hexnqkwuxrwMv0LSoz0rsF+EKUUSsnwEr0x1e+zCK41SGjatB2aEugy
iMQ7EWTYy/JjQFwOWsWdpClytMmHlZmAXTGWxauLQtM5ZtC6ZZjDt4RBD7KMupUD
sX80EUm8qvtvGIaNNRoTDka7WdcBA/wvfVSiZhD9JJVFW9b/SNPlzfHpN6+WCHSb
btHnG/2+7NX+AXYVn5fRt4AUv1kWXAG4IQoFm4Cg+f+Ev+MX+vbiHiFL8/kEhbPr
0OAw1dWNEEif+K3UDt805FUEtInbIXO8o1iMPjmi+gYt1dUDrXkgTlwPKHWyucdq
vFWCiIKX1nIuOLNMavRSqnKSTqg3Q9OupuQNbasLRun95nnrnblISdCxUgJNbotA
gOPK9mlCNVmMCsDPAfhFfnY65itt+wijngA5Gn42cellU/C10HwzhN3y/wS+KrxU
HJ1EQZNt4/YdeDqd20LaYoC9Ig1WMsbHO0PUCaVlvPsmjkfZ2L79PkYMvpeFzQzb
k0qbjzi34315xS2SW20mB8zYYB/iKiiiRwefCqqBeiqe9IBYMXzydzcmqe0qDaSu
9lax4EyEPXi+M9x+3RrDIi8AsRnOM9sSnh013n1/qEYYyMo7kAIVf/EzTU8vvo0p
uH4VdBlmCOfnPz73KQkS4HNtx99RdXU6yK2CGVEWvTXzdt89jwf9OoyQfc+S7bFU
3d6wR5MyNlXogC2oKDbx8iuJ9/4893gDW8cQKtRA5QqPpnUVkBVu/L+V7okMaer1
IQeHYPn3GNp6Djv1V/vShrZmqHpgrV46rum1cdc7rqwjH2y6vnWe5MI6pGbucqK/
7zAOoTTLcyhVl42dvw++NVTcFFAkOw/f5V4tmWJmkNRl2dRbCLNzS1kxImxjD5+J
hJcKCDsEojuN9bwXTJ32lrzxDiChE6y54yP79q9SiSV6Eoc5pHbdmAe3H4E7/Ztf
TFnOcWIZD9AtJFzmh3wO1GkDNqFf6DY6dMosbnWTTnwwPK+pkvhe7qLN0naNOeMP
pCjIT/Gaz3Ghod+yQRYa92TPQRrYnkUmpUQCerU8T/KCZRXZ5z4nj8IIOGA1TdBr
wfr1s4JEE41WpSxu7+ptptw3bkBIvR04SQ8H3dxBJZWkRvHUSSktsGp0TnhoYZ33
z6ApSFFJD8+ItRsD3junvJyr+EoVA4JnaF4OoLA+vrkPIfPNXoZVQGL6ccIsQXri
OKL0yH4B3z5jlldlrVjafYH/ydPszYcJ3Cc1izwwrD4kPMQSnj12EMZ3mOkZM9uX
W5LOpsbsk+hkiCyChKJxu3NfAz64RDDXFwA6LQBEw7gVlTOawB0l6qw6SlTkF0mG
IWsgFjq2DyeNeSl4w3dm9H6h16jGoej5Hf1cWb8jABMTxbkTIGG7dhrMcKf+i/uD
KjButjcsgvnn+KnsdrdtV0AUd8N67/YOdmUxAorgVTm/yPlJ6n7y/6YS7edueP8B
fT51jSwCX95dOY/qYR+GzmgenUCC47NL45dR2sJXxrMWz+jWsFLhX0Y5DEmM0/q7
NHL+La5Ew3NhGPSrpBu5O5fNixQI5CEE/Wg73rSFeNNYWLlDXaucNXh8zCZD+E4W
4B6r8GS/fAHXbQCKugSEN9RBWSKTre7rAhGl1l/lPUNenZKTZzVy2mcMsToa8qGi
wFvSwjUSEOK4FLDUf6sdFeE8fkoikpIgY5+cPtR1tCdpVeCCmBHxmzce0Zo9Skw1
K8nAzhjlydfF/YhKCRnGeZdR0y9/63jTHKCPFk9icy67HZynnJeDRiZwYLSAf3KW
3oGSsQq/t5kE+v0izG+Vt3OfKTRBQ95BnXTc1Y7BWJ1Z09FPLGegwD6sJWj/5gV8
a3RcdcO1crLoM2QIEf1041AWX/tKz1e08YHd8aQY+zaE311Tzd/QiTQMfvSoUfJQ
VjFlIHerNEVZoE/pRcL2zA==
`protect END_PROTECTED
