`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z7W+f4WBSQp8anK9puQn/wOARzSM7fz7OO5jgWLK2FwCSWRwN0+HwFyVC0i615iM
bSy3epkU0H1kc+nO01WJeIEABJ94NrcrUleIdeag4dhz6394E889zbDrywqa3ujR
NAnbpwsfG3xD02go66YZdo2l6hgQq+zn+y7lnLK5YPGkPXYSBtk6VY2fLdodNXUU
S4mw64nzOall74A6mWx4ddjMCnCpmpGe1eEI0jQfnTWBeqhZioPbvkwbFjKfLp2s
a7kQLYGPqvxg5U8A1Mbyq+vV7TYvF2M1C9DATUFi1wkeUV4Jqabad0TVbTVJNgov
4zlWFM/jWmaukv0cWennMWbNV6gtDP6/batJQSN6ikHNLxHHGgB5MZTK5pps1xE4
CBN37xZYP9fgDhey5CmbL2W6ESo0pR0KJd4eztdifa3R/jd+Gv4MyxD5rMRSZuqP
Q0BD6qamtrQyzxGqpmPoNJFIdMyKLnWvxajpX7wvE6qd9BsumadIRtAULiXmqNtZ
f9ai8f8h95bz446eGwc/IWGxYF8eMTa8unuAHAX0kgRDRfJ3uCR0OlbZFA2Zd+zP
Vs7w2naSOHBIQ/PAhDU8HdRUrv9dTUN1CeV4vW2VI2cK2zFwzFnenRDoCoyV0IGR
TGxQ2ouZTnZaMAXyeWQQqf+g8qkrg2U00nsSpjfkKrzy+lVlPHLlfMH8QR8/p+OE
ZQ6P56G0gS/DTmRD6Ticc/jwJ41BqJidlPPnVKeSgcN//B3gTWeYL3jXEvmob1LV
MQQE+ldqDWGGYxqJSWBg7MsV6BQ7MIAvrfw46pUKKXs7HlmQB8HzZLvvdcfy274S
5MbNcU54uAfXGBeBGk0Rri0roxbcihnVx8gErO5eQFWYo+9yDS7SI+fT7I8sjC6X
lkrSD23+0tD3OmTuTPGXrdmFqzwvjH0I1hl2OPwyj57C4K2EONNGBEaK6/ftNNa0
`protect END_PROTECTED
