`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xtMowpjMRpj/lnqXhk43rzv0N48RonC452fZro874m2D/3QhyjJ4UrGXHjoxTrJZ
ETeQwLGpd47bCuQkXpCrydYCC9X4KNZYje/HeMaiqbsTk+VeFspVWfnmvOJNdB8F
LcNbp/2cq0og93tl9i3BDXhduyrS/XsXPQckU69NximS7ysaxD4Keiz1CiurECZX
97fuIZsae9TIRIIXZyaHKjj4PZ1ywDwTIbXap2PqXV2wrHgPuWXnzOK1MyfHBBDx
6l6DKJidhjACjhUvXPQhPANi82Wf53fykGHw+aEL+sX0dteubJw2OveZrHo1nr9Y
pqbo4ZqnbbM+igjU/YCimQ==
`protect END_PROTECTED
