`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
glDBVI2M1aeYPn0DL2nfdq3XEeeCItH/NkGp89cLZdYooZ/qOmgUponSdvmpBQRy
UE2sjGyfh43xb94jeObOHubrAI6UJCV2E8L8RWItgxQ/7szACw01C/8a9xFIHTnK
hg0TmsoECCTK5zIE8AkUyHX3ctUObxThAqFAM9wKfnVkpoxjt0Xm6nTXISgNQpOT
ufgZaZNhNL1J+tjY3r8vbt5CeaiigSsZRmLsIwm0waxIBDP6xwyxzv7iHga5pm7r
/wbmFnV9Q59zYu7s3tp86g==
`protect END_PROTECTED
