`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3d2d1ZasWg6IPhz7hrOoag0/EeIcvsmPx55xQTKET6S7RyivpnckxopjIu+to0vN
xqu6+cnydA4RxRRdTgkq6Gatja7KCKmp/y6nMzgmL85R/b2tp7eMrmLyjaS5dCm9
9QKRvBPtvRPQYZLQvngKhxXhDV0VZE0o0W6KTmBHbpqAGnOW69UAFUsv1UXv+1Fy
k/CEWtLUXgdalYGSnlql/hL/uFfCACON/lWCGOqoiGDr4ipmFaEdn61eol2Xqv6u
8udwu0/lHDclsluLrP+5+A4+NOONalz2ygO/hu/RHQiE4hT4IW5r8KxGrtCJFK2y
ePIMbWOsSXOYzj6DeAo5WtqgVLPdoh0oCQfVy6yME6l4xYf6NG13bHn4bBvt0TYy
UaSOISTdgDwzP6g5XxYt83tLu1fpkhrK8J9tWPmsiinKQtRIYOlYykRd/bk/Egfa
Pl8sgkta8WCHAAJbMaKi4FApesiGpuBf0b0GFoa7cqgvYKyqBgqkMNcsY5dNqlnK
Sr6c1jahNVyoEGojhybiDg+xSzYL8bjcXmSd7iBmFABeCQDJyBHJej+5XAqptU7S
NIZsC728zZXeeA2cXNrcBUWfwKk1r8+ylTgWel+nAUAo3h2yxl7wTarFwrlZgeld
8uRWaLNZrcZ5UMynZo+TImJuDVsvHKhft9hjEwGA6LFuhkC4Lk/+KlwsVaWkRjSH
fAUL4N+zCHqdwr8sTK+RmXE69+rbEsXVmroU93JdMJ67ef2HZnqtzmeCNaLAM60z
ncYtSVL20jSsJHhCp1GbDg==
`protect END_PROTECTED
