`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ncd56FfCEVX8Gcpjj8XHuV1iAS0/yrI2SMTqVMqtbpjH0ON84ybvd7gSU2lDXVic
yEjbc9qerdJ7plxcZ8GZ3PV7qN+muxAW7Bhf/wgD5IxVE/OPa0hqVVrv/zFRgtdG
sw2htn2EV3xouwarRYlT+rgsHs5KjCVWAdVwNtw+YGq3J4+E2SYqs/WZ7uiiPK97
wk2CWIliPuPMz0MNkcb0VjIVHNBCvWUwirSZvv/q+HaEcwN0+tMbGwExd1OwX2nV
V0G/Rf3sX9sU0iC+hjuUOQ==
`protect END_PROTECTED
