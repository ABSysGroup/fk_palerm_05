`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hOuL81uHEHXvgpF4d4Kih7fJo4o8Y/yXMQgVFUs0jPd1RXY/3ah03RBIOSR6iwka
NgmgXiYVyj3sVRrkD/AWTRMBIcYsFSiu+dPx7xf9H1Mg+z/E67C/pBy+sMTh3xRP
iqtegzlUgEaokoHDq/V6AM5ubwDphiX6H6MaKh8fkpX/iRV4Oswlv3Gf4z4QH2KO
yfeQ8Ms8hkrMFBbq872fBB2vie34WPQw8Drq3cBj1saUz1pigfvtLMpV6YHnB1D7
d5/tQwleAC/nZwmf1KzMOGaySFdoU+lEb26Qrx/0wp6nl3cbldgbI1CeXkrR/TZC
CijsIZo3aliBFlvcnYszNnlr30TmZfpJKF9wmgLYOWWnWM7b28Z2o9SYicVtqPIa
EmnxJoovY0fbdo+4xv3//CRe1CLSI3PtYqn9K9J4Wv/lvGIWMOSTGH1kYsm6uDfQ
Xf0uEU5qfxDB3+WQwW/EifzQAuy+W58WgYaMb3C4ryuvzOG7LvO9TF31cKk6jkri
IpExcaNtJ5NEJEa1Zy3pOMYAT9uCS2+yFN3oPs0dte2KFNUtKDDEKciQq71GNz22
SQc1df4HQnZLZcg+wN2faNu7eq0OMMpqfLbXy8mrlHuNlFdtmrs9Yl6R5oaH2b+J
XGZEZ0x5qd0nyp83Xen1Mg8/ieMe8Ll4pU4g7/RoBPZrCztojLEtwJT44wXY4vnq
0zyBzqZij3erEWD/Q6IaXq+9V2dA1b0agnvkaOSXjyHVS6w6XDxEyJ8pU7mtET71
GBcJn3zQ3vr5qLAmaAjrT0lacP3rfCLLgNKaztyMf6aOm5lrWn18b//olN56mF99
UnI+lb/+Z31rREwz6doqZYYvkvy653VMwt04WA1IqWsA7V7w+uTO4cyDG+tKLLTM
`protect END_PROTECTED
