`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NrRPRbMRtvtXtafplkwLIz/HbsuRJ3T8VKnDoNQKE0xCV3DCTp/wdf0aPxTLCXjI
/t2PP/xEKuZUJAumTnco9ldUTQPlTJwyM1jTfh0afITfCDygLpSppxr2X46KlSM9
0abwbRxAj7QnW2mbhN9o/ZsMk0Rk2mb40aM9m6JACR5Jvt4HvA2QkOy1GanTl0dk
s3oJTBY4Kr4D7/rJ+DTJXEDznNaabLzYhS0X972T6am3YbVlLbCgbpQ0aRRbFwT6
iaMQAG1Dr9YFs+47lfowrLJdWTymnhNNc3MtBIleUsCBvzRc75f2qsUO4TPfC6O5
AiV/0gx1QfgzApy9BwS1Ubyi4zCQ4lgIgcGA0TX1xdsOnhBZ6HmASfjMsmUhDads
ZLPfd5XuJ6tICJIrZn0fzYy/bub9ESJjCix8Zhciu80G7LOXO3mmBbkgTjKh7Zo8
0s6IjUl0SThr6JCihFkdjJxVox9CK5ZEAhVS3Rp1fQVpLcjoWF4Z3GEQuWQjNCs7
TrgDMN0VWLa6U/nYWg+a0X5DHcv+0070HWS2YxRSK26mbt0DDLKYAgd8soT/Kw0l
R7fV4e3rlxdMiRw8/3c2pfwTF1czrGxYoGvh06Ixdstjep8Wvw07ccjFsRfH1CoC
Es3iL040Uqn6cz+9CxNLtUVIrUAen0m0/oYjzA20YMMXrDFqHY5Yya0Qjc0Hbwua
Cj4cUTX4SYBIra00x42m4mu0gDt7/EPO0OmUL64iVo21m8ijdG5PTYKzN2qN5bsD
q/fe6SYew7KYiKDC0SbSGeVU26P+QBbmzXp1jg/6sANj6CkAMdBknDqFY2Vxr3EN
g5OPy6f3bgQ/B+kYkBN2Th2+13Pne5aG9jkw0FOrDszZITQ127Eh9R01MIkKpZ1r
yk8MDUMriJWIr4bavesdVWcLF5iiTC10Grj8vP/ga0xO7eR8YxMpp21I6BMjk/Eh
8YdC7Sopv764hR4TeQGGhoAz1bIPd9h7iH+6SNYclce+a9yVvR/KHrcXMoLNCiwn
KK5GgN1NZA29q36ml7c/71eCb+aSQ4lywZr/tdbKP0as+UWJkHsSY84GAMGjBEsQ
SLnn5HRUvoYUdj4T1pAXpx/Z93hO74wGDvs1643xSVhZyltLhbWmTkb5jYIB5hty
ZqrIJp3jzuKpS4K3kcInqsZtnRP1WJoghMtrBGofvJR6ezqoQxgBCHWCgQDWuOnu
kxoHB9GUCDZxZQCubVzVGn9gzj+n1utnN4zr3iAwDjoSowGSpvlJO2ED3Ov7dbBw
IylW6ufVQ/KGGWxDmPu4PMD4Lypw58ks6QAMk4zIdJtmmVJvK349S4TuFDsXiY5r
OUG7Kw30aipyMoFDER3RDas4R37EGFvhIpvgsUZGdrjgaBVF7wQphv1d9jPw8AIa
vfBZqolMSy/J7opaDaE8lA==
`protect END_PROTECTED
