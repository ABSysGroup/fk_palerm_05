`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VbFPzV3R+WrOh7o09wuSb1AttFSmwiro4kbMFl2NcesmTaIUZBVH1M8mbQD86lKH
ax4zFl8uoRfa23LTDtjLJa2iWs7e/W4LTARYYvJM2cQu32emUqZubnliA7WtD9rd
UkwOlWxYxrvfI4P053CFVoHgRmKFkW11LlRk3V6MTN5sBF+hYiUGAngYdc/M4i+n
qJ8kice27+uMNf/hFCbRSqIsDEer4WcUaSOkoLwbqsLGgW5xUROUW/PlPPGXfH2x
tpZXTQ1X7I80bwJMm/FCKNakEg+aTTm2M23BzK8l84X2/SVoinUh7sTglZBa3wt6
B09QKHTaDN7/VC3JrCLkqA==
`protect END_PROTECTED
