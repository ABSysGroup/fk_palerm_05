`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hdj9yU47JR08z3StJuMC0csC+sXxAHTVLpHhAlSqSfsLVahnJpif8Z1TNIU/HIh3
NL4RnU0liw2b9IIpE5L5xzKDbkD+Qx/6DdtGLAp7PhfGtvja6ipy0vq4ygTXW2sU
01FEzpn2trhA5CP6YftRjwGk3Te85I0F/Uo+55KfpfRBv4vdj3RTc4WF8SXIQD5/
4yVe/8J37NnMi/oqBfm1nOusPSOnr3+ltxFRiDW4XJIXs4rBvJDxvWhrgwT4BdU5
aPvpt8aBancTaP3r3OoyJIrFoEd/CADi/9R+fUzOf+yw6wvqSVLFXQdInp/QxLYS
Ma4oFHb8YYjnJsjIenft61G3W9aHjJmCPzVDiBdWuuqjtDJMeZnau6mIcj1wG8ao
k4T1HC17ekwl2lHS/S4rB6dja9pYXkKgK8ChkLuJKZhHwRNbFIBDTWON85uiumt4
MMst53ij0gSUhPVk7uc6NyezjcQLku1p6ZFUC0wT4MNpDRqI6LmYCvRkxa5NTO/H
dWYjcHj5BOPlvshxcmHm3xid0ehI003raC+sOh/16rm61oeyjK2I6kJ+qNAdYqZL
vwa30Njt5AEPiTq0q4fcYJLu+mGm77/X9OtA+4oeN1p96Yh7TNYvfPruHR9u/aRu
x1JKd7ywHP4n72KjADSUt4JkURGFerVAvUihPM9ttAAbPTzxhhNl4bDTYS77wfrh
w3RgE9p7ymPgpjM48x4VfQVt/Pg19tkcew+e5SUTdFQZoOu0/ZYEa0pZ3hMTXIs4
K0ke3+894Iog9B+x/y3F3S9nWurdFl6tN6u0ObVlDLn3ndH5p1G/yJARV9LjAZHL
9dzIldL3icJOenzNQA6TV/MzL2SbIA0eGvcQJZDPIQcqr3h4U0ulc6/hPbHM+kNk
bIr8fxpi7sshHurQf1QrjXVKwHbUCDAMdkNjfl/nki2NYMlU9Hl6bVtC723iCo4+
fTORCoDjP3tSiBuGe4Rb+aBlxa8tHlhwyqXRe7Njx+MGfONWonYid2dhTFT1bE/P
i2eEmEGHZ1IHk+WjAlbLzSAK0IXxoOvC32wkHVEDfOfYNwxeCsC/KkIvaeeKUI3J
4ECDUkPP/DNQ2acI84AzYaIoUsYp/8HM1cfHOOV5wJ8CsuFzqYXT5F4mDjW8kwfz
1eisB4o+AYjJwuRf4sUx33z5p40UKVBx2E3tj0IyD2xA+E8Jmb/3jayGVQtX/pCE
ld0qmKeVYFimJCcWNIIr//2C59+iDOlg/9So4orwfgfV0dEVJq1VCq7Kq3EnHzoF
mUu+kPqGVh4QHOQ1PEHE5/hui9C5wjBlGh/jZRBa8XKHV5t4Xesf95BPX0yvYRlw
P+9ByM5cB2zhKx6fFXYMjwMO0cwHe+S/ZSJIksb/3i6HJejGJ+D1oL5qeDWBIlBm
hDbH1n8s2t7nXj8EpZb2oldGhJD9U4FqRMGFdpv5F7yrymPqXDzORuQQtmW49KIC
t07JUMM9BTicHHCqKrtKXCIAXxrtoHmH1xd2GXFM95Bver78W9mg0MtpHQIsBPWA
r49AWEAvjXkCeYbNu9E8vHwOlR8TYUV2bqQ79f/SlOK2y42IObv6mT4xKQu00j7z
Ar7n8QCOcGzNBVO76D/miZkkMUxp5ILG462/Y41O5iyqI78MN8BgNwV8qqdPiGq9
7MxGRuUQ641sXG86mKGqkXFi0SZ4LQL6C2OJj44z1wFycd/ypI3fbdPWGwXlj1o3
wRDgiuVXhnUuyJN2D8q+JMh21EhaNZCNPkVgN3lyxoQnXUAQSF5qP07XlliQIJlI
UQl7vw61mikGmfUuJc+5p0CgTfnFfVDN12s82c2WvwS4n0tvH3YoSR5X4vC3VDQB
39ja2yLdCbdsNTQjI+/Mk7igVijCu0lHdgShOdjgSFhmhawHszUuRzadQ7nZBqNg
ppfEzOj6Gof9Jhn0BXca9fFYbehfjFr6aDPWxmsq5jPh7PLkKx6eeEonnJt+8z8e
mpcQxoNZ6hBKH5ibPThL+TKrvIAKmed94A5wTi1TWp0LFZbY3WgCIV1iaMsnJZA1
OXYKFRflNX+tdcIVyyWph7i5aeXU0H5+en+Y1W83VYhNDjAzoQb8ypy2LWnIPV2o
jz9CvMRDbXQbxVicFtgTAkYHcBTkzxkoEiCDbJUAIGFxy8SoAc18Vyz+v08NUmmh
J2d3U5wXG4LgMfhyCrORYPAX/lLJBRA067La4zjw/zhUd0mGPxm7SVNXcPsOPQx9
Srd+r7yMZjLdyy+wsxgemnonyMnD9aPf7UG1Im8vGrw0Utv1IYX9CCWfjKr/NovW
jSKQhWrVMR4DaIgVklIqrKYDXpl969gtiaLEqOBMecvm6hmI9OKdNbA4t/g+JEJ1
+6QvX1Y6Vcv8reWKkRSNY4cdvrAGhSIaVJTPyJNu17AfnN2g1aUxyS9pLH+WrEkg
6rjW3sQClcMIxjsqqX640v206koe9pH6sdUVJtntwlu5GaMjIeq3FEqCUO/NFF/z
HDDqc9NszzisCmIgcauSbY6b26eLPxej7GZ2okZv0h9JGPxWP4cYNTFwG/nxCpX5
YYux69ngddFeboMQPcOGWjI2VWoPh/4Pht1frW22SiNQ1V1Q5FdxM5otd19IkyJk
SRRKUpy0gF3gWbzO8i+Cj0LnO/Cw5k5yJ/54rAA/tvnYpxiYSWW2hmQz3LGsBNsH
K/OkDYc6BEUP18uxs2VHmkTs5ph6FxMtHC/V94THw7ZAZbz0RfXbR2+Tt++5QguB
HpbrzF61BVYa9LgrGL2C4XZ6SMnJkPTq3h670RSAbH856sj21wpgtZ4WN0y1VRSM
arQmsSt3uE2CUsu/6zEu6mzSkhOdnUdeO1ehB2wXxK889sOsS2dH8nXeHTjQf3vE
HRYyV+qbOGdk2/lqqm26YJCgauplT/riAqWM+IHEQuLIDIEJ4S/VQJ6rUJ6SAOau
1u8okZXxBk7l81qa0iXT+gc+CV56TTBBjxSf+x+W4r98ljAt86mFqMnOYcvcRNyx
mqzVhOxX8QrgfLw4u6L8OP1D9gmomWyGeCghsGl3mPRmYwHAnAekQ4i7acV+/yUu
Jcsa0crvf5ryOlDsqjOViY7E8T6h0ta35ejqaCPkZ+cqU2F0sr9We9HYNnxRYIfM
E9rW9rQi3Ps8XOXJVw5i9mF787lN6sz/rJRqAr2QqMEMefI7L68oDrL8EKylXb6+
1SgbVtftQYBTMOE2Qa5Iycd1TaLkcB0w0Aaiu13e5dGRTv6T1Eva1A5XdAUYhARj
5nO0IX9KtUCdRKpqSKuiGsyBadykUbSk3EeBJuoQUTT2m1g1veZpfWIWvXGJM05J
smZKiPb6IT+FcvsDFMJlxSVQww5YLr5ARQ19hf2AytjZXi9oUqXOH/Seu6LLN42/
HFq1U61TYjYBgOkuAR8IA6iHTn91iue4A1q5coDKZoDuUEuwtQDRUwVkfOchFUEQ
dR174P+7FqEaDmiZfvy5bXj17R+Pfne83hrKqgBoL0uix2Y1kcHALUkV6r0a4YQs
APVyZwZB9gI/S+jr8HECoCp8xTy8tVBLlic+pwJbC4KoDonZq6cEHsrv3Za2PNK+
KrNBXLQ9NrzFsayPPvRoGbThYUDEKn1GbVT2hTJTJnMpBfTMOI9RX1IFrSXTP4SE
fdSlZRrPRQiGdkQHFwA0nPxtSk/2o9wvc1zl69JkmEjnCm88AlyC38Y9R2tvpPdJ
f7Ygyfqj34yM//79CVz6sPBw3oTKVfGYzzlMNhJQ4o/spXraZlVpczSNv0csH628
Ennla5WvEpowIWmVU3IwJ9dgRxYq8VrKEvy5NUuxYmke70bkMhzragNZgY0tgSzq
Lcbm6E+fqB39enyGdEtMtAIuzdA0sUoP5jUI4gzhniCIbEh1whImnxwe5XlLXS4N
vaqg3SAXs3BOw6AJvt19xak4EcpFWYzZ1hcT33dhmvBJW7W/GbnPbHHmLrJwaBRf
cz8V1+IMX6//DA+e95kPkqfKS4DDdWyAClZaMzCYbaCU2M5e64Igz4ElDfT80RjJ
+3WPbXerAQFJN11tyD4a1v7936cLR0B0vEhX40CibNV/HdsP9WicXfBhnUhXtFt5
WxKeHeyxstbF7GdnG55ZVyt7E9Hjzd6G2VDwoHC88C12NNzDEL3gbfqCQLknhIO9
ZocoieBlNc9aXJwIQvovP4ftZYTsEFz80oMGFppW+5UZjLX0805Yoq+JiDVjCG2K
DKnKGnLdnfG0YyCmBRGc49VFmdW37V3Foisn5x7tj7MvqTewLQYj6PBhbpprk1MA
XoS4i2JxXjol8EaRhVKi2BNuEwKkm+TgpC5ddDL9k/uGeaMjYtKdkaYLzudaYszk
VXYC9j6T3k+IuOAvxYqTdU+XpZTJ7SNfoL7CJimsRxRNaYpIIRQkRJ7Nc4aBm9UR
nwMvWm7aZbnEqQOy+l05449nrb28gCVlm+3ZNKq9pd44RqMi/PWj6aJUNfx3IPIe
0H0zZOW6wmd1pow51Xzvxz4xRg72m4IOieKh4EVZN06pt8gNiq7weH8mT7c/2SgB
y8t0iB0ZAdNYV1sS9hO8fycoBmOIHIL/MkaD2mdbX4o2kEpxvVhXyG9mSA0ESLyT
s4s5r70MVMUn0MB0PjJvBT/pMue2Hzr22I23G6Xys7293WnEjuL2BZtuT5vO2HC0
nR/BualKsYrwyWmZOEnOCHnPCjIbMdm1OfO0yNYI04cti2XuHTfSZGwNSPl8znGa
ltp3LMFh+S7S8HVXWoA+N9g1gaX+fmpM0U5XalC79x46l5lguNlA+XL8YpwYbpNb
ZY1Oq/gUckM7AZWIxtK5VAb5Ij908zSsjHzqKtnp+BJTvnChRw38OViuDsEH5lJh
U52RIvPXQcCu9FIKNsJgYq8cpo6+ttrDMkPV/81D/FXtr781gFr5aD5JBpI57THq
Q0s+n2gbGHpLU6WF+oSlDwHQPz9Fvzd8gfx6VSUj2aATyH8PIRr0QaW+1XKwgb6u
OvTRO4pTe2PNF8CM27vXhXbm0Yq4vxzPRAJ8Yh4DRmtWDSdU+o4GA6/dkT0bxWIU
oj25znRBld5/WM3h0QihBiPyvE8NRj2KDaymY8Drpzji6n6TP8tSAM602WZ131Kj
rXqldQbHcsJx9Tp+Fi3goKndhvVi/JOd+YuOmQerAKI7ZPdgcDpCA5buAxlYEhhq
g0nQuz2Va+91g1ksvRP1t+FKiWLJcpc/vSnw+3BlL0mzH2tTB4Nh6hPjwdKg24PK
H1vrf573gLgTwvXTcgHmz1nkw2frU97JKB+Myp3EVMPsgcYNi00a63PDMPBiZRIp
ltOTpwrZd6fJ8+LQQPjtv7FEnx0g+2mn0pTuPSmUrghgVK1E6281vKOvH/LOiJQl
uoEab4vW0nJPCOFwj7xJX5aHsWJuwdSIqCFoPZHn0up79V06tDDpT1anIx1o3S23
oUNn7q8eYpUfeHEU3OZba8PqA0GSuyE0WlClA49WbUhcqOL7nlDHnJKFHl3oHJZb
cLLMfic9DobdXbsAQg9I7eKHoXaxDKOh8B2yZTdxXwObTrilDtsuYTQA39WFc612
Ip2Cn5oE5QllPWdTqt3NlTxnb5PRR0hQioR5ySdq4bRIm59LEYNUZyU7BZrwvEJF
bRTX8T6/+/YDD9bxG3qrCiAEYuBH47C4sNwGEBOz7lyYFf0vvWlivkdkF647VxeR
Px9pokVCKE0/kO7S41Y6M4GBYLEehN/EXHW1Mjk3eQfDJR2ynR4Ehu8A8b6bfmjT
/SAeAwm2TKuIsWuxD+Mm80CgDaynACk98oexkgHiQaFMH5ihWKIg1qT4nBxFI6D0
wiL+csTRxUhTsNR/w5gysiicNyjfh+VjVFTLh5HeNTBhwkLdX/X8nY/hn+qCQxtH
3QhyJ7m5i5hyv5w2Ci7t5JbbQKCyxRc8vTmay2SFvnjLcjMcjntf2j7dVwANBuic
xrBFS3QF2HgYU/te7z6gpWDDfAoJif8MgU8rUtYykRs2uUjLD3vjUq4C5pA974h8
371lcqTm42KSmHMCWMjiCiKmL+6Uos8a9CIZ6npLfEUSklJEjuAa48U7+it3iBcf
PfU2f9kzdQhFoUEnAFBsvUBUzYZgNtLLAe78Wvyn+FNatB8tX59G43spXC2py/2B
NWnFd/IywR4mmv5VGrGRpmObmQhcBqifau5GaHHTfxzF3g0gg8Wg6Sld4pn4gVgF
+5IXytl15ZreogGHd78ZKeSREVvc1T5etXWvTbQIbQdtqy0iAJj2BZLVmfUqgU8A
Z9OMcC1PwTCpjgXJ5L3B5h5fe+DnTqlmMwvlgxn/tu8VJeQM7MNKcJWog4xuy45/
Mn2PXarCGVYJNHueRVf5DQL8rU16miu13L/KJeguVIwuSMikBbKbgE9w5JUWHyJD
68fs2YAnE/ZFV/8sgSJQ9V2WqCGdaYSXtR4dGCwam0uf2JpyjgebX0/Lf8uGBD/D
qN+13hCT0a5JAZ7Aedr3JQ4CAXOBzw5q63aTZq3NbfAifkUjbcOsT6StguPNwccs
R9Wkjdr6Dij3mD6XXyEOcuDHo32cO34xA9V1nPEe4mkMUfg1u/sjI/3CastTFRY5
EplGjTa3QNqvidv0YdyTeFHBGwwF0/6V75j86Bjp7bE9jMrXzxSgND4hkyzg3D06
TAKEnoW9u3kUfEC+kUkceJFqwMiDx+WQEpxhSEMOm8Qe0PDoBCcFs2hWtvGvdpIy
MLtYdNcyWBdVxMoxQUDwZAfTio4UiE6BDCHK80IF+0oze8vP5ezHYhLgjjGECjsT
eNc8MONp20Fyhy5jeRcKBOWDDtJ39VjsPPeEIZX3V34yHADDtlD6nPLynPAWkYc/
iRxVd0/z0/EaTraTtdhhkEgrgW8Es2JrkDq4cpBTr8/PXfTiLhzoRMn/MGkGiTxO
xIOUjPimg7PziPFt9meH+8dcHq+8KdOIoibZGmAe91+Hb3QP5HwMU/JGosynPHpQ
j5N5fUcbb4bDyxTW44isE5g99PNa1owxd48rv8oW4v/ulzqCTKzwYs4Xaq3jYAJ1
OFceB7/F4w52vqOpWTHusAG+lLqBFK2qFJK/zMh/i27na+187LlQhvcfntgLjHN6
O2XjL5FgJJAp2+KTBO6znMUG73GVaxp2BYnV0x/Wtb0ik4kPWXlFmOXAugRNr7NK
6YwaOOqutDxOzDMEqLL20/xy/AyTOOcaSbESVf01X5ppQwu4gcMfNR/aacYwiViI
tEHVhaBi0KEsEX342PZ3/u+RjzAZrGl0WFBWyqmFkXXN/2ViuQJFm+U+oOevD4+6
qEYNLdp8fO3fqk/aYJM5EodLyrO2roeMG1ySKSu7eTXmg7U6XAZTXM7WZYkwyFUV
U/1oILMWord+IJ3y5tUR5Z9DYnos9DlFScpEASKFSIizTxFIPOC0Z8Gij+uham9i
IQRR7TDyNDRO5QhFn19jND/P2N6TcDzSRfdDcqPzHPjdLm5kVmV4ks8xrR4GzgyL
tFjQVj9xFkWxPeLEojS02eENYEBEjqBt47fS3jUPWgWfld8zQoczA1t2d+zW92+G
zVyEj0QqJs7BoB1vATlIIZyZ0nKFKarv+bqDrYeAl1TEMHZOHi2BaXvVO0oCzze5
+vmFg+F7N5q6Jp8C/3P5N5XXYwCAdhCZBTpz+0npoRLTvl/0nShBiRpjofukquR2
aH7etWlKxSAiYAoMvOkMKB8MuzYJzubfGN8l8OQdXnbX62Fi61ActgwGqHiG4kh0
R6rwX27vXT3JImXFStNwLboThpxOCcTkXJ9+dYOAc+c/bduroiS/3C4AJWfl5b0k
G+avKKCG3M/sitGMB92ibm1XB8dXRPQ/9L8eeNpfNHAWz+8vLA5D1DOYLcZkxZ4L
/Xyy5njX26+ozBfR7p0mYwDafq/pWqeo8+b61NsDrYIO6KWmNTSrXFKnYNKyhEPr
F5Pdwm2vJYv/yhDsTXU06q3Vo9lc9uny1pXZ7qwVznAntbxGIWRGa2zm9jrCQsBQ
vmOExp+J0kWMrzASmiZQ+FFotF1VQmHgFCprxGlo3EqEjqLfYk0qWVbHmyOUZ/kE
+SX0v9qOfeU7gBgYmuwdWUDxpkStelKrCE+epl2m6UkOJDMDxzwDMEanZ+e8vZvI
eNjmywwCpsQ/BhHmhRIFGPugEKrPaOqSFBZXI0/+N1a3j85mXzUGKXU0+NSDb69W
9u2N8mQwZ0niDFLdKrq4anJt4jkvqj7HBEVO+uEUUf1xxnNZMIS+q1DREr08xtDm
vqQfigApLxAE0fnonscFjpY4w+4YOgbVXqUC9I4CwqZ8oE3iBqueuwUQBDGvembO
P0ayoxajuZRTXfamuW9nJIKizFqbniRYy0UnEoRTpQVN2v1Vq3vLQjAQJTTB9hco
i4s6/0Jl1YEgdkAA0VSEAMghR6NWCiLfcFAq0+HuQeSWvvshldndO4qWMpXOXq5G
lhpq0nVa/LHTBinf7ht+5H21hrgIlT+SmYx2Iic11zOoE4qbRwbL8o0cAd255Slr
ZZX2fkLVROFPy2EKoluSXLoRyg1DWWw3BRYMZqfSeEP254K0eTn2ptcOXG4AnsRk
+ipmZ8S8VU9IGLUZFkxAClm0/gOLfFn2ChLsxMFQCRDXFlLzyHi5HrfGmO04V2QH
H+hQJwWs7jTV8E+hfeIUMrmv7+PhcjhDiiBgByea11E2X65Lq9SKt0yq72JioBOW
71r7mvgkSvrrgJCN1AuBb63XXZoGPt8rOQMqoyjdtlmETXqlnjN64pXuQpmac9Ud
dJFPT4rRTquPxSn6qY3ECixFKbJpNR7C3POkFz/NsKR510q6w0/zHaAivxl7EO+T
ZW4RX46rsvNc5VXsHBUnO3PvswFDZ7Vdi8KtlPZ3JCJaSg+CG/5+f/0owv6huQLQ
FCrbIWXV6Fs7DANwmAfxUj/H3dK7GKPlNTOIN11jYs8k93J4RcC2vLP9NvNw2POj
AKM+yH1rMZTkFEvQy5fYzhDzEeJ8kmM4xb/TsYnEsh8qOV5BW+B5u8TRwz6IWEgF
usYLDzoBcH1GumOSSFl0z9harhV9wmeEWxLi4aaRktrFnFPmcB3QaES6NjF2/1ny
59lVc0fLRkawQvUSxDf5ovI2+TxEdoRji3s1X9Fn07tPhcpT3/qUhSNrSAdUubiN
OivItlmf9H9OF5mtzlQpd+fWmYEcokYNZqJzq/gLV33xB/sxkMSu5J83pBLsMWcL
t5/rGYezgTH8HXg6rH9DZQprMkl5fbX7x6bOyV3PjK7rM2MfDj19BFT7YqE+2bGE
jagyrAut5msjtMVroKw37AH6CoTjmuMd+Ap7Ue+dXj8Ew5zqLlYJ4p0vvczvBm0v
6PhAfZuu0rP7Zeg+wfRlAOcBelxG0o5nVFM9jmaGhRwTiNX9TZwCeda8Il5DQmai
P71rczwOXjsTbkYnVVH8Nn5H9/UiiBGhWhHAfoiWxnQCK211vVg2P1KlWM0UPgcI
fUay1ao56hD3flump/F1DSYNMHgAeMU2CTjdPSJb/Pze/rN7YsTNJDnBR32va64E
5rcDrpBncr9r/+oXhKppveP7JFxu1iLjqMlawPA2X5/Udxs5TjyIY4MAlVmoqzbt
EiQcVfbQMh6WnmckaGeYmqw89QQV1a4+G+hdYqqAp1XEIdmb9veBEf1xvUX5EcMn
glNhT3aEmR9g8SknKm/R/CwQ+Y2cNEbCP+SO8W9q3O/SUlobTQyuDS7MT4L571wG
wllFiHFW0j+5s9es0nBnxawDnsvgAHInDXzLEm0L/18WHO7PkLW02wF3GO4U7ZeU
sTY9T5xkIst4ZoyMDcxnQQaPsd+auNfpXicQ1nfFWyObqRq2hor5x+SUL87XQhNI
UgnGFHd8G/IY3u9HbJK+xC9e9b1S/BEFiZo/S+oxN33VIx7eQzW7QBFP5mcD2kDg
WutLz+eH0wFX9B249vZPB2hTsFq128A3nafC6ApEDEdytiYi43XBwh7B/NRyWDv6
xw2vpMqTadf6YgYiS3GNEICnMxMBtB+2PRLBZe4qmKWoc+YR46aNn2cKNakveiK2
8Q8VTcy/7fmwll0eS1/V2Lz903YSdsvYyXkbst9BF3DFc5cenBrKz3rnA4d7HBZB
sGtcXWWyAbB9rxYZJ6YkYKtb7QhNSOILNHhVcNY+U/lg/RQRRwdtnErn6B+9EIVS
kJcfhnzGzzHfotPw763shB/rBb1oHwWrImMi+hAktDfSikimGQE3+BBRb6Ir7Uc2
G337MkEFGxSmIU88/I9wIMPmieua7Y1Zs1/rmcUPfIty5nrwG9UaFSRx6TJR5R2e
0ca7GOrujF6use6eIwIIGjrys3zCoHZnmyTK8twvOB141bHbx7H8OIQs5+nT2a91
wYkJ7lRjmPU1xq7WbLdULaPRf0rFzZqY+gR22vHZ1ypoKh13DAGfEFOwB5rGGS2Y
2fwO2SFi34BMxeLpJUhReF96wuV71PR4i7l0emuJrteYpscKvuQpKQVS1HeE83SF
OSw1PE6tt5RR3c+to7UyLRLkttfIEicVi6HYnSEJtoX0rhlJLN/MCwOY638B5ZWx
EF+6PJChDmM4xbQgosOKg3QHZsuJp9rIwkFRxHWWNuYFPJk/HMMrRgcLxKixoeqU
1iDkNGW0r6zYjyxkGvEGzzsLe8tYQyNanEnHbovX2qBypCDqpqOsISgnNFT4jPqV
mKFsEfmgUEbopBNURCguicPm7VuUaWOYHsj3Sp7gyTownsYhYyWKFaqfJYMdspVR
eXvALWlR+4EAW7p1ln8c3+/aGKK/lDpsXQLWlVWESNzIdzmUTf9erox15l5k/p4C
+6OqA74qYhqz/kEvrCsDMzYb1+z26keG9wEFjiw750XdKK0af2BDNmSCuajRh6OC
au3JzErd/PBnVydDf5XGkqK0tbBDjfKWnZ6pjUeIq2CA24c3gY1Yu9WidW70Xx47
XUnbFGyeQE+jtQNIKWfJXCwiXLgORSseNtzc7E2sFInOK4ozlHks2i8I2pKZ4086
N9LUJmf+qvHWPqU7qZQL7X1kXroJ065zeZdCdoGKYhNTQWvMTxkcLNokL5JSVfXU
+QcrVFSPLG2Da1YAEkQkxgttbN9FdsiaHyhrYN9wayO72ObVd6UC2o6RHIEAcMkD
C8xNFvOtaj8gr0+MR+w/xIVVqL6NjKSfbw/XwvshOL19QtAnCrUkEZBVQgArWVl6
/h9LgNilOt7VVVp+j0UUkSJrmT5GhlYejvFIoRGCiZTQr7elQtmTXoFKEcSqYT9c
lQzc1o2K6LLWImPrl33XSCkpxM3xkuWBHJvdqGHIxDgEcAfVteC3F9c+WGbS/lPJ
Mo7QQp0QGdNDJ8P9Y7Z8s6VOyMrrK/ooXx8dPGSRFqPgi+tQyTX5SS7Z/iQO7PC4
fO+8eVkgIQtKrYCMzdYW23OlL5+GxZH2mzIST1fRxd++zAZMIHnht5ZhU9H4PXBV
8jEBF2sxFMvNqidJrmpIRj0IYSHmO5xy2NPD//08JVlSjALBpp91lJ2y4Q7iKK1F
69WKooxWhkglwqEu4QKUJKnFE6lLd/NcJ9acQdIG6ttSW6cDi74dzJokaN8GByqP
j6SYXMxDVpcPE1vBEyRqC4vbmvclRNG/8eUbb1FGXYPLVHKkgljJNw+iGZ/iO1gD
aVbflnVuXJGvl//xVBzwkPUhIKn/da5cnhzDNKHM29PpGA/0oXbupqIBLuk8dV/J
l/Q9em1gE1rqI6ruUW87QWU7MhjOFO//irR5BhUJiAQYoaYAjJZn2PKGOiE4Kqas
BgaF3FBSuSMABUmT9LLZF5OXK2nqfhIOVAScvZFfvSZp5kQ5v4O9ZNDaW7fd8lE2
Q0MKZKoZ5Db9veICoAIC0ZZy9RBVEHUW4blM+vvq4XrJosxnzyA8uVTvZUapAg/B
P6ROaf6BBrNgMYxxlKFS0ZF5fU7ml0HGxtnwEblTcUX6U8FJVg0DwcQu17I/UzUa
ux9nIyl2dTKQ+1JO4PwFaQT0mEs2QafT7O07n+99T3uWBIBiLJHHodA+IHbCzMB+
LmrTanc8WfMz0kyxcskq2GoSagsq1uSjpzsxU8tP/6MRnBvnWdFfJX0qgX/M+ATc
9luhJnPZmUjkTE3BKzU+KOMv5gZVIXCDCK+axBn4QSq4LUH27BzHN/xDkrTyu7Z8
UPj1yo3Cc2n64mGiW1VOb5AiAi1H+DP6EAMP+sPYxtz+SfGXsM8p1aGAQN6MJHpD
ZuHwWptuPpGHmdo3Ks2LdLflkfEyxYpZwRXMiQZPH1wZ8HaMCv4vJ7rNnH59zDIw
qFiIaXD73pSP5Swv1nIutRzztc2k1g3PiAFNu65wx8PVyMLVdP0sm666MPjEYbL5
TqstEqfDfTuiHwZJFzYQT4z8xhT38/BbdNMqw7gfsaOtlHJk9hOsOuUHsaz4kBxl
PfLMhDlUXcMB7XUiWUsPuVGIdZe+AL920WqHB/VrDzHif8vfbQX1Whi6pecuI7be
juwNpQgrZa6pOaL2Yk6TXwQQ4oCgjx7XBEGPQGY7jdVOIcUuptzjOqRXxL2+JNog
YPpFX78l9y2nU/XQG9lVwEqI+4xHDfLkZ2sR3Scho1mtTpbylfA1D+zxJoyFfGnB
GNBcgTV1uoMCW1bQXbHApx2wo4eseib0YBPfJywWtWagekiao9JEC1woJE+nU6p1
2g0/Xgu35oMMEeMQJJ8Tw6WguVbxxC4RjI2WsrkIVgebiRY0q3HExL+XI1TDgq0D
usGLzDw6iPqgvhiiLH+7JP6ET5RvtGndkNQZQbB9Cbu9XsJCIPWJgbRTHo6u1rGZ
pRAcrCeaURUvj/1wkdRdlChnF2bWSFEUQe02fzqgOX9gODGPJSLZUMG0HJAdzACZ
uJYnofSEwOJV++wuV9C4ffxrOaJYm1TmHzfnVomxfZgO7YpsGkbguqaC6vDQaqg7
LI80ZYottbSYK1+HeXJAsFjikArwtu3hw+nBvDzdinbjDkFm2QSAoNhcoaidsn5+
ewc4TUhJ3hcY+3VMEpMA0GDb2P9wJrGcP5aqvaTQ5eXLO8eB5KCMOHjfuI4/FRl/
1mgsyRWr1iDpFNc7GUiRF09za0Bzq9VJvE7mcGa+AInS4r6bnfznKC5P1dDmGCNW
A6OGVwPdIJsKH/JnYoOUAsuAImqhIMwSsaQm1Zesv33qrwYCsLBlvo8BmdQZQFLS
ltsjYqDATcm/D6wjVfDW3OOH0JorYpmTLdXX3EoNFsnqWuNaMi0AJvCqihBecNTG
1XDrWdqcawLUNk8WMV7VcStPv3hI5pAwZpCF/nDCCFsMuTcx4/PkuAQcdv3gf7pO
UYpRHw/SwUTu8jFQ6m//6JDNpsOfhAZSVjwmrF3C6N4rINLqQiI54dI8qdJqyxHg
b0JamreJ/7FKqg+/QlvzuD3zodLvvF+11U/G9ZypBcHJSdLlU9fTemwf3UCQo+hX
C7f+40M/5hbByyLoin7AqGymkRBo/NOWEUbj9rRn8W4hulOkItF0j3qwnl1lb1dx
BFofq4rs1URPQTeuTZVOvdEhAePjjjZTjgrE6uBqbmrfMLPPIKivriUcxX424QS0
BBconwxtVhl7Yx3QexlplqWmbKPRqaWD1QbbE2tTSF5EvskHzZvG2lEInL0fZ3Z5
G/zvA+wy9K3hNApEQYfZl87JmeEAorYX8l5YEuwJ2NreWG3QCuUaOdb8vrEX+xqY
akkR+LWl2Edk5CTAD6gou2n+ielk2Fa7Vm41gtWgDcERcKibB3bJ9NBxufX7gcS1
3YfR/nLTUK2/tWheeC98hic0N/97s8HBjF9IehdziDtAuHv+5Oqs/+hpQ6j+o9h3
YaGVhOxxqagc9KN7H4Mc4XKHu9JuW4zyiX7cRJ+0Fe9ngtElk3iXTfJOqROgItMm
USRf9Tsp5pcHCbqAQ8zF/mPL8s9AI8TtdKH17qxXm/5dcwjEAMHrluJBnNc7xPNg
zNmTit9IyVMqDzjlDiHNX5LURhdnvGZivvsnp+13F+XOeIidxC68N3WeV6IVJBAN
64s7T/+TYZg89q10jUjfEI3v6reLShB5K/p06afB2Sx2SzFMqLn9+Q22xhWp4sBm
RMiiZ6t1o5qLWILhsDs5bSFJ3UF4G2GIlToaJs5YDngFRMixm+XhTNsBCBGuLfeL
wM36kujOhXsZ1DlxlYZH3voqLcTtVR2czgitOCi1DYVlyUdcNQBGQV4dDd4eFCF2
GR9DmI9KfGtoUKQwjeVTejOOgMOYI0jGwMNlXmVTrFZ8R0uuQCJK8cuXyIRoSXiE
FBWeFW7jd+cW7Vd8M2PKgYRkcRYhwi2o8P5WdBN7yWKmE5wqHNMZ/jVnC8JMmgiF
UijggNC2vsJBbtu5jJ2pW5DBxPD5FXBVApslt4JH9jsNC2C2G+YkVle9eGG6KiJR
FnJt3aTDfi8R306C+z4Z4FsVXZEF/lwV55VM1sWD2KhqN9AZdsclOTRiyIc5Qx/H
XGwvjF5RcL45y/je4fvVzNjUibgEt2SB6lolcRRFjabym3h/kaKJRap7X4fvIe/3
Igc+Rb6I7Tl+dfMMCvv71z7LSzF830Bt34PwKwK5PsGPw0kpPBpFE6LnuiIxltZh
MD5+pFWpfQFtXIBPTSxMxLEO9WJare2dzDmrnQcxGvlIWCadlqxcfJO5tDW17V/V
kJm1q2tL9Pv3kLx1Tv7+v6/cLjg2npeASD96ood+4K2xuZlBuTHAjbojTLDSRiGL
Wbv/qmDaTUfm3WBiqJH5HHDbtvh6CkdnLozw2UMmou/gVEXGPGAk9AG8IKshRt6J
E73XAXKarihLqzagF+0+lEOmKjbLcrPandK+J8iE958NkVUuZIAr1k/eQvqCwqUG
GiSXxRBhh6B/zhz7rbneXhbGmm1qy6emT03UbUIerxz8BAMrjQ3jLcjPMA8jikdM
9nFuXBxbdVA60jHuN1/PwtN+R8FQK/UtVq1DBfWn5IyG4hyQYOyS0yscEeh2Mg3C
bZd6BLWErxi0Lijx8iiliLFTUX9iNlcfOa4zQbjn2tar3GxPfw8u3hLfnvm71PRb
HS+jyL+o+DBwy1RaGYOIy9M/d49baKh1/UaB9z9zIvISUxJLD9i4vj7JSWAZBvBG
FpzmJUy2OgSNqJlQVSkQ8g7fCW55HcqJ7BjYdi2TRyZsMw2phDNLw0d/Fi2+rA0d
1EEt3ZCMKHqgF+RyabZOHBonQdEiMgRHuC26TlNPMqCoe/Y2+sdgJxmfdMEbislT
Fdg4Xtk6TSDfuK7/ZvkF6I/Z9FEQnpbTR447L1HoFFJgmIHaL95OyUAy+B8SXR+L
TB8VHPofoGfy3G6eEOwNZxdH1zP9nSxOcOBpir0abJLnFDXixi2v0Ve+kNtd1IFV
NlBZvDc72UNOSYiSWd2eRAF4lR7VrPWoj4BdlZxL/BTOk9jbCMJgXRPlzYjTKskW
lCoW0viCmbILee6m9AtMIvjqHd9VTRpsTdMsrzI+WuPlRhxXpxgVCy5VNNAbSbvs
WkiGAYgMQj/CnchB7xd2pJ88gshYolauP3BlU394nxr5+aNXdV6DUydQzuxerHG6
6pRFvdb3c1Cpf4fJpHirdO3XwGpdxgD+Ih1U9cA7soiDdg6NuUh3rUlWzl7mfnO7
x1sCHLAJtZ/Rd9tH0WVRbqeLrjlsABk/1Zc9s7Bt9FQ/QaH+FZYRgJInxG9znasl
waS9zZr/yNSU4EKdz4JZG0Fro1l9Q8DhJPT7GFxitGPtfwicbmKAI3/ZeAZ4H/po
EAyI+xnuIIy/SlN/kZFOz7n0zlC+U6jYvE2DUFxlqqiTWK0hi3u3xjC/kvnv4F0V
jpIF0ZIpD/0fKxGttpqp5HPbZLJXRA2BCRi72IkOqJcfQP/8eszgy7WWt4p8Isjn
eegI6KEjAGT09Ri5mE+J5zFLMe8asab6A0dot2m/gK1vwzB7hBYPFTEYOwvrj6GL
mXeT5nmkkLFQSF0DOz2t5XpkxFjsU5dWqBqBjDU6ALTZtjDqPe+SJRmLDD8P9acp
7ZM+27C2+OQxTnDWqkT/lYpw7kOtDBpihLbNSEACkXwWzNHH5redrbPJc3/7KUpG
fQ11glOkU7YIuWpPX7fHPlbo/tXawME2xdO+TL7r9fmQpKYCKr39mpt262YNJ6MA
u29PO1N7rZhV2NkFkd86eOfIQvl6IlDSyGdEPLJGYBhPWXe4I4rPBE1VCJPuZ/Zu
DwoU+1z4tLhPE4OzcdnvcP8x8otk8yH3KTCAYkfmWGS34mfSySJFTIDo2+OXffWU
sImOu9tyDCrmopP8Qa3fFg==
`protect END_PROTECTED
