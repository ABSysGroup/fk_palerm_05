`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v04B/KXJ9kfPICuVEJ40TF4FuzomE5hsDqV+A194Dw4p0FMDa70kxft21Hd34ygZ
cFPDOd+QPNScKv8A5hxhCFwFx9RO7oj+ST+XItuppBdmSraEvJYRVmdS5O0VoxPi
PwCFFG3gBuU8zCxxppWHzZHuZEej1xk7XXB1LdxnAw/+J/cnyb9WDAYm/LAvvr5v
Huuynt30mOxEK83u9rrO6T0gax2h7mf/Pp2GFtS9hq4rko+LJ9ynIWe2N45FLUsw
Z3X6DzeYqHaBfN8ZvR1zZOHBsaZMdNejRvvHKwqFRYBOvAOc5FsONVPlK8UMcrdh
er2U2oH83qUHXxXh7ADOFRRiijkAFfRah2+md7TCmRUKzvJ9z5NN29yIEcBqHTXC
1qy01p31lEBAykAbhLZ/pgEi2Whz/IOXFmudGLJvgz2iXjf+IxdOFA/2xlTqM5+O
1WTjVX6d9U/I7zUpjqXXXk893L+NrA1wY/SsFNtm5R4Cxy7GpkGMvEwJlIZMu9Ww
w5zMkZLutOzS0F9xVocQPY1FX5X5nmuVpRi0dDzTsRL43xrEHhzeNFLShUz1UpS2
vlhGID/hcKJ9eh5mLBdHBV7/vaQL111fy8Q1Admr01bDCpI1G/4v8Oj+2VPq+REh
QMmMbiJUTSMtUwO8eHOC/g==
`protect END_PROTECTED
