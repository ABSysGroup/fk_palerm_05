`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9wJ4WHYkyZSa4MoDym9poKurJ/FXh9CWJvRg2kyZo4rH/QZ9KMbg6du6nQLJzcGK
LB5hq8z/2GmQPW1YL8XWQ3R9uHCR6GbYTTVgwZi3HKNhQT464gqplnJ7KxthbgDV
fQLjLGLDCWoL0g39apg34wineuEk1ErIRZ9LKFAYW4KyVV6ptA+0o891sO78VpKh
X2cM6ZDf9c69NpfWzcSp+G3G6oROTm54TZ3m7oRFWXi890KALrNbrTMy3lSeVKZB
JoAAMNTCH8JomZCxsT9DKp48gcfrb4PhBAT5olJplt0FqGzvMxdECsMILZi3vzYu
zUdf8ILNQ5fgYGR+7KHX82Se6qijGTu0Vf0lfoL72lYAPuwAXY8d8m2FoFPcXATd
`protect END_PROTECTED
