`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D5LPSQSHohD1XSC0M05VRE03j/ePlRXkixtl8xeKRdvP9PKkBiTFe37Y3Dk76Ve4
1ano7+4K4BjMvsnDP2JuO+i8mRhZxlFOof/uxFRx/uUE9AhZ7L5VL+8dDer88wzW
gOeCZdfwRLhr5RwuxWRbKoI0a1WXmslZjB0HYJ4COZAO7G3tI/uIq7SizfTjXG1l
5g8+Lz3iJ6NAAMBLkso9WmVS/ZVnIveTqjKtWIMYcpVbs5J+ixwv5QLl5AajLJmA
Ur9TR8aJj6mhfxfnBYTwBvhb3V0Fn9owqNL8mwYOXSKTalngJPkdawzwAi8pPQ7n
wkBR5z5fYIVx3w9WaJeNHmqLLOaXcxgtT2Y+vCiQ4fNCKnMNnFv46WeWk3fwVOzt
fMNckE4tcg44qk6ppXYrxd5lQ/UBFtnSzywTcZMlkhJ25lbcGpyCXlOLsWB7BDRP
PsNoptozx3Mk3QgITmJZevj7Xpsj5dBsCvjnSYTB3hHv6fB6WRod6rQI1nHsYO7z
1xxgLd7Vmaet+B0QmiEwp8IOHy0T0b/0Cx576KibnT8=
`protect END_PROTECTED
