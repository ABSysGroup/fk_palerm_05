`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H2ue4nBzg4HOTNUBUem3a7+NxvA2zYbgz6IUIPNLNVWCUKcmVNCgK+V7TCzD0zA6
rNsVF+SFis8S3Hi6DKs0BrplgB9//lqx1fGyWZSSY/3MDEH4zT5vTNapZM1FA69e
8UCU7dglKSFtYuuEnzRp/KyXakwEGaAleiQb65pumhGDBPtJniU0Msf783qCMmki
RS7HEqJ696PQTSISdx9TXnMkZNNuJ8O3xdgYPFjDejAsU+CroQr0Akf7tC5TFBm/
HbJ90WryY0tiWuv1OYRUG0GF3Nd6oq6kPQMPkIGWllnFCBHj68USuZy8kCx1kdHk
l8e//bGhE6GfpgiCgxkkUBAr0cAZxrRaMnsLk7wMWjoWBbu0NjKt1FnH3c2VJQUr
fW9jG+2NZsHimeVUiSHWzmtuk7JcaX+aggjMtm8gs9S7cd5wddTef+cl8Q0Q5JYo
yfNOJN/UiO79T9EZCbCeBICoM4YpiKr6R80x7ZE2D50HlVtsNFugDj/H0+jTqhq7
sK7fMWOlNNnuSjff2Gj65vr/+5D5P3XyKBUbRDicIraSqBAN1PwhaPIgQUwCvak7
eX9NYWqAvQXGjJFKL8e65gA7xMJeHVcAAKowMOb5awhiUek8JGXWXIlg23dCangl
kggUm8n5cFBatwfRaejgwV3xl6bqBBSJ5SYr46cnsicrCqAeYSgGpQUvX0unwyrS
byFBMTb/INqf0S4kix5nBg==
`protect END_PROTECTED
