`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VBlgIOaP8h/xm41g+fBKpabiDrSx1DA6czZtT4eRqZ6BhchMae9qozzo8xyv/F8z
hhz1g39UxE6pajRZmAal/GmlvDWlE/IVv+tUSwjM5bMrCVr6uKlCk3QltGA9Tfz0
ncc7Dpjy7+me5fLvDWoKwdgQZyGftmHdPoQmKCvoFzv1Lf54erJ5zBy7XROFN4RJ
rfF8psPol9dwp+Q1i59zD0yjrLn8FfbObXxLSiCWytn9fquaL16OE+nkKUDSjSBk
H4buTwwiWu57S2BXrSTOzS8+mKTtFx/27j7jZh7vwmDqTjXrozc4B+dNA9onHrdW
mZO5j/yRaEtF8JVMuDR0G8D+X8PsSLRDVk8ttQl+Pk2co8oC7Sm5zDvFpXEVWwHf
feTzqKpseYIcz/JVwbgdVV8KI2Q5T5gkoMvmZaEBKnCDwr5OWv6Gn2wwHHqzab/o
qRwZBp40f7XU2/8cu+XFsf/+pGaX3+Fy4bYyjfUJpHklyTzrBxPR6W2qy90L4EZ7
`protect END_PROTECTED
