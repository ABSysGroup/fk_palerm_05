`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0DFjIREOCU6XoM3/e6DhuvtSxSjx88h/I3Ro+LYF5GEJVs/aReY2x5oPpUd6S2Nn
0YektMMU5nckJuGS/+5tOXLqabpAI7iivF86lhjmNrNQkMzi+A55MScBtyKEnkp3
IgScuwgQHk4DhS6IE+b9c6SATlCE25B81In/S/4jfhnv1kvk+9rqXIUS9rlOfDI8
6HUkVxJTdG6UvzYZnaS0Htc6kERMX9bxY/Wmf2zWr+DKTnT0+n/lfqWndawkGpcz
Pxp1S8fdDKbV5gmceqh+PVliZA60r2Q8H0NwJdI0U+tGpWOc4K2GhHnjPsHf8aAI
q2vbd1tIEguOxcJ2WbbMdfJma0rEZug/vnyYb2MKOY1ABe0iYn/WUJUBSCthvhpp
jwze+XY8Pw9DRufpNwI7VkgNssHoxO7XiLc8vO7LvWP/h23CxH2IGwdn5fx3lTB3
IrBtJHns4t7LB04/7txGLSMrPxIDKzO2I5bJ4S+IbqhsuE7WoQ2cqL9qoxEdZxj0
/dg3jwGhajeR04U0175nzw==
`protect END_PROTECTED
