`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R2Wx2Lh+AfaswJR2cvqTm/sH6jRwymVO/JbvsH7s00668I1GPASll7G7JOI+vegI
eM+am+KmgnqssFB6kKomvGfTRpYmjLx9H2FrlPCekDgh/KwiAmRlnoZUhF41oIH3
CTR+HIzu5kds1A9V27FMVtrKHx7aUjfT58UpsuMGMPxPu4eERHapGai9FQ3Y6dxs
rIUHqYODT3NJHZ93f+mxy8bm6S60iYNWUVb77pJ3v2uGmHI2rL+c+7lkaVNkJzzS
fCVpHw6Tcw0R78QP5v41/LbNHA8p7FdEnD7ifoYQcLKvbb8qjBzunlxZxUWGpRUd
dYrrBoHPMsXwb9A38viwEBPtRhBbjytjoRBi7L4qNhY96Rv3bC/nd3gJk5p/4IvA
x2MQ29JsyXyY218eX32BhkBfNjToOuhXpp0iujirFaXtQtdTrWZSMAZJWqRwCIFp
mLX0vCUygYaXRB9XPXKFHSQdPZ2wzOjip73Z3jj12EA/cUMgZkBW3fhkj7iLLbq9
VPV5DvH+alqeqNlefBzjM3PoKaPSF6MASFhM9FrV2/8zr22rSEBtOvE7eEfjM5GN
Cj8ONIYaan7LvciN3klOsrQ6HATdOhHgZeib1EbG0shvdjT+5i8gQQL3Go3PGBmq
+4kOQmPhsKV2zY3A5SAv1s+2DDQJIjMKREdB8Y53QLgBJCaRDMUwIwTgwIxkegY1
VIWErHX2eTHFz0ZZHHv/j0qHXTS5yUVuNg5vz8v0hDEXCJ4vJoTGRPv/MwoZYLSm
UxX47BIfOG/Y1bcTwfYhkCNGndZB5QjeT9PTfs7vpSPEAqPUnCyS/IbNNLy2KmK8
RCQoUFXuPRha7NHWDO1Ea6GxKYHHT0oqAq2Me9YindIhu7xpAVdAUcRFN3xaTByj
VkBeByQnIYwiVn95Wpw/oLIiOEulRRgDykM/Oe2f6//B71m2M82wfO3Jagr5idxJ
Ar0cBrNaOyva8HflyTySYruxkcbsuz5EG3Fr96PhpojUYcB34e2H4cJ/czDcfp7j
lH6SjxWNrgTRMSkOAg22I7+n5v4s/9cirDMiNS7h43h0PT1tB9w797ogzFE3oZwK
CB8+VbH5HlchITxBX0S4SX5RNQNBv+/euBoakD3eP0SXkM1YKIlpbgtlLAca1QhV
EUi063OZB83VRr8lGPjdceEUsiBOyOC5KHh2M+WEMF4LuV5TM2V16H+A0f+ahWNt
DjTdUiahhbtB/rq4Ox321LBQ+ipuUNeqdPZw2E1OSaljpWnTB67nXXlt4aOrg6vj
VLJgKjC8VgdzmMgB409xsiAJwWifqNKYNbxi1s6c0zJoQTyDBQKHv0pjLHXOsKF4
ojw1e0TUrwRovDjGoc9twVH/DjwWp4eNJxyxrazW67uKNL5YFFumKEvxBvabr0TN
HMQG8SwpkzPps/zPnIsWPdIFwRWlGTBhZGrcfA2PVAtBK/6iYTbpn535YNkCesuJ
DWwtwCApBw2Qq7Oh3oCNgFFnl6qqxkpQ0EhZ+YhWth19AbgFTBptkdDIvn4YSt9J
Nct0SUPpEB433ZVloJZXzBePGQDe8lba1cAJ3HuMZyySn+HMX+7TUkSTFU+NlMEq
VFsgVIsgg1yzUzwuTNdvFyfI+0tX4qATpLiuF/wUgOot9z10eu2PKL3xK3NDw51n
PNOWHIhqGIyRpfkwdyZAIjtpNBnjTM9UGip3XFfKWfkFVc8kIvBjQFOER02hAfpw
9zp3sumIyqmxcRt8G54iih7eRg0fhkLLJuQ4eWFzDpQMxGwZzWq9lqGeyNB4LI9c
SnqX10OoTlWeCXwUxuNlBkpIOQSuJwtc8/y/kC0HbTQAz1aMX8ZhzAn2t//WuiiZ
zES1IV2it0F/cdQRNiJs0tBfiFM9KCuS/KYYN8dnqtVbrFKiPzQoamcAe56MmkBH
/muBUDpsZOSoX7mquQyN+3cKzSamQJh+wDtGkpPAsVphxRgQn3YWEPYn2vN8ZJCN
vHV57exFAPTY3P3t85JQP57AHq4ZtItRQkQ/Ho3oyuuvY9YPAsJTj79zaT9CxUy6
rlz3ELPAVzzc+OE+DJ2uR77GXBFhGVCqACRkwGbGMCyDkcvQGalj3fRlE+rJIevS
Jre8Kn525Bd9YE23rjdvc5HEnVH1Tmo734L7oMY+elAzAYiiLstGzEVpH2rkKY95
r3g7TZefSxow6ZfTCnj7NaTGTY2xdjbuNAUNDWyz7YZLMl1NTAQXcCNE5FPPkqus
WS1DVYjsjZ7wZcL2gXYZZrzlEM1UWPOzYLAjnbzatrwWzLZiY260imU979rQv44W
iKSSJoItDjjeoNApE1nmlWOUyhVTwvD2BBcZ21hMOFYaDt4Ze3K/kzYV/T9Vqfcn
yCiGC4Ivhl57ZRpOIsW/9Cmv3ZGfoNsTs/1+oajBltYtyrEigy5yV7Yq+9t3PSxT
9UEx3EH5GSW6noQZZ/oOfbpGNVumy8zuG/73OOotSPYEztNWs87jMlI2e0tLQC4m
pH9A8xvm7uqV7wsu5Xp+AYG4yW1w4kg9BJGurmynnH/15+t8ZEcrsVMmTfaEFKbs
uK0uMM6CB3gj4N7QNAdU7dsLDNpbqOVaJ9kVcEtIdWdTi4Y1oh5ijpN7wFVXLOoE
N3gVmhXAJe7WSJvOgsYyJuhSz9NmqRePUBVb8V4LpRPRLgZF/v/Li8aho37lX8lW
SM3dRmRwRcKiKvu2LiwY/Eeaa51oPhVqkPue0PLDRyc74eVt905GGZMLW9ZIE5s2
f4dO9w4kFIV5hI7qHGcDMHAZYYestv9paQc6yQx0NW2AlHuV7dPPkM0m3v7jin13
0HbVD+hddO8GFUTAtwyL7dB7vqJ2fF5TVEy6hvNl/udcEpi3v5Z/Px9lQ/fXCLx3
5jeU+ci1hOzeVP2r0QlLl1aE3XcKc5CAYQnNRqyYahBwg2hmdRblfEKQYXpjvS0/
1tN84fB8QgzZiAIW0xlyJNyT+xacukct2JOXDgOwf2Va5DUL4eldErlRx3nLjAfD
zwiOOtP3FtPRoqXIIctjKW0m3+R6CA60UWxoPFULYik=
`protect END_PROTECTED
