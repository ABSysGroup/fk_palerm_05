`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o0ro1uodGKzrCRRHEFYgXO212kVl7CWb8r0s3QI88Wo1898XYWh6dX+dmq545It9
hgRHQBtPMcjfRAGTr3q2yVGOerwBi4bZD3vhKkceXk7kTJ37mtIm7fIwtKRE6Y6H
DqIpicwqJ6UbN785r3tFh3v3W29VXMwBe2q97lPAwBdSGyZdMdBYK9HqvAfIT4TS
MQY6/K7Qjdy3xjXuM6zh8MnI7O6DIkXAM7mbsR6mDdLr3jkOOQdiEzDnizX2O40I
QTDwVpB9QrHMBWJbRkMjzupIk/G+nY8AIMzSUvrpKn9K3UFjV0D2gsj6eiJF+yvT
jNpVn3nACNz1bI94Go10ShxrRj9PfoUP5PKHgcsP+wIjAYIrZV8QqEb/P0yrJ3V0
r58upGqNHX50vb8J09pohUD5bOhWjXd+wt1/Nxc0jWkUy6xQ1NMBMSqbs19aGIok
`protect END_PROTECTED
