`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qVZEyLRdHE3S/L7IBFwqe2+C7M9f3oeyBQXZLGVYB/furkpvnL8JuAWjFxNvS6gg
P3ZGef1kVhB+Sp7GikbqhrTMlwDGD26bu8wzrifkhX0cJHzP9Apfu1ZYwS/GX3IN
rfCglSaScEz6YFrOC7ZR3/bJypr7Rr4bsa0PPOPSmpvSuxWrjZdCaQro2On6Wb3g
35TObv+QdXgiitTswGXSU1LHtpFyDvd6y4YRjYBS1M48cOPWFmUHJfGt6pwe9hJ3
1WZxeuL4QzrVQHhF00A5lwLZSR7w+SR1tRS0E+aLDfrEvIJLnKH5emxcAfwjQwU3
7Zp0qucec4QI8KqknY23mPTW0Z9OUvMKkRqqghGo0D2AUuDYvgQJOROr2bOU8Dgq
hLbeKIf/bxzE+1m3fl0R0BXs1EgR95zjph71vQDvatGy1CG0Nshyzd0WzS3o16ua
G7EYfgI45wxeMNnFNnZgVqpObJGXYCYs9/1nPkirhGdiMsteG0WizVLfNhKqJzNe
HB0jeMo6u+8zAIRtQVfVvhN+U7WS6TtgdZRvUzThKT+IEZB3OaVNHewc4mlOgLPq
Xc2b89jyhhJV6vLYN1y6CoKagtNDFTxYfykvQDohlKoqO70SkyoRc2W4H/XORd6b
vpbQZm+qo3QnWNrjWrFc+w6MUCXjeKffatZfFzbqDIApJ2pNZTP7UawtNUTH6Buv
NXS0jRzlcThLhc2b7mcwmq9K0uGL0Cvva58HeW+tylJpoHXzatt2QUd4ejBOWE8+
NsBZU3/MTKlVWHJ+eUzcAYKiiHpgu+t0HIUQ1y/rX+eFwTe4wO5wBbYwKh5D9st3
QbsCtmOt21YRC70ThG2qHMhJVdADa0Ca7qsQz4Siyg8=
`protect END_PROTECTED
