`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gpSioxdl+MnUlqJa+SGckj8Pybm1mxCVKU8f67gYJTIGyaVOmi6DhSr/gZvqXt4z
b+Y3xgYUauXztWjbNSp+hRnxOhMRNuyHDBzKXcAiYhOKB/gQT4dDbZa0aWcJOx+y
zMg8g7wbW3YxkyGmq/+5D3RiwazgXM+Ow3+rTGS7sdQuTNqpjf318pFBOUdXHZuA
5oAH/8KIj8EZk9UbO4AUZsV9qTRYzlmrgnDwsg+SDDgh4PLeBKIJuo/17b51J2uO
CaxEsf2xLn0IgXXkLMvQWbxMLE7YdB87CuyiyYgJn+DAm8nU6Bs8eEtNqVn29ufo
aheq3CPYkMJcGaN/cUqYhAb6IjgGTi2CW36ycIrPDE95oApU6NKmQn4jCaP2jHXq
`protect END_PROTECTED
