`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PSCXD7hLXWAAfZwS5Hl3C0+sVEU0M29VScfJvzF38wRhVkPtFKaq/1+ZEvry7S23
E8H9km1jMPCIxnQzL6zwWCADCl5Tstlp1s1nxCTNuuEVqKTybUPgVIj2TPq1k36E
flhyhdJOpGFnUo++SU3WyZ62CqBnk72Jc76IFSwl6PUIOiN9249pQAvyOxSNPM9N
+JqYhAKgiZXo60hAnR7LYH94cnAiJdzUjMSNXh+EAJ5IT5NAfEPrYgGC+gGKh4FZ
f7T+jwlVFT27fht3u547qq+VRDawK6zGLbQRc42X4AR3Pt+jDnfjEYusd7ScusXe
/XwJPCDHQuZziqERVr9y+OE8nfmULRHRSCJHVCXG58Jai6iJ/GRHow/I8QvaO/nF
qjeQJvZi0zz9gM/Scb9GpHnhD0euLDLnnEVqE0JfbPwv++gGNujuifISEaep0UeZ
s4wz12+pWfuKz0OROx8/BoiyQy1DZM+TVnsB4gdsxvJDdGXYylTGBF+kXVTmJfIJ
mT0NmTYFAYIYwk5yIIyMlnLEwisqbIOAwyxTCnV2R9XdNmBZ0UBJ9oj+/xxLjAHJ
/JELB5bBI3ThOxouRX28rumbhFUxW0DB3uednyqJc4VvC3mZbp16XFCXUwsXUww0
UilbDvhG/CIV9ejr9IwHf11lfrEMNkT3Q6DVhFSAa5Zh1R3FIJ4AcP16lohWlJQS
3+WTAaWQHqqdPk8ANs5XTtO2CJ3cRX3FG/T7PV5RXuRW6qgEbdshy1M7dKooqPlB
bsUUIijJQ0BRoqJIjl9URhQF4qG6g6zjiw9qJjOAUhtHijVlCyyosD19N0OBfSNE
HXIMaH4PiQmKyLBTt/RcT6PdwAS037At6E+PNHIcUvJoqsEE3FxnaTmrD7KNo0Wo
gT/voqT5cVBU6v4SZFlIjBnneXatW5+Efd2DsskAh3TW2I/sOpxTSxbgnyh97ZUX
rYXNANcuuvTY+gRmkdhjF/zidWd9IKEq8UoR/sQr2SWCN1us0LgYzX4ozcAz95dp
8ExQMHi09YuvSg7Ya2l6MvNSC182a0/3SHqHq3UlIt6hquqR+G8CiqfxKW0/rnfu
xax3N6u2Yr2clNmrTLBGrTwXDFeexLAyZOuyicifetJ+tDxmYrt+sT3KO/i262Ba
w2G9GaTN8EQMtdSBerTMn+wJKcsXiwDw6yKzcrzyWxCMrfq18E8G7TH2TA9JUxzT
hmxs94HZmlUUIqeVPYBCcWcHUaHDWulKWE0H1XbT9fFp+NSO63qmkBlt0rbzGaDe
9EzDxWtuC8AZgHtPAh1NmeWRKihxH6WNOnXXFrBPmfH+Q/6VWcslpPHfIXiYkE5U
5kPHmar6sL3dxI98qeQRVlljWaWjIEcI738hm+2RlgTQYaNkGLqczfcDY01bmK5g
StEdL9DF8h+332O796k6bqEkJ3avcO1Gaj26ZmH99QxVhksa9hzUsBbPA3CwQDl4
pBTZnnunc6hCbj9KK61dZ3uEFb3hS8VqHcqY76FE8f9YRx75nitCYQczrvxKMoc8
aSyjS01Icf7JbTsbFK6dUNbzezllseNtuSgSFPqWix0XwfM20ay7IIOA+J5zmXEc
GE8kJ0p/O1GE0PYyYFUJpCUK1SKKOwYpIlVdbqA5nq9AsMVep4usr7TloJPhs2Z+
xipc2TkqWLumUKUXIkhP8M6TqlablbS5CJtBHYmsSIPkYkGu8jIEHoTqqKtko/Tu
MEHszDyZx092loWkf+bM7KjVWn/z+tsZl6mxFiRvJtX+zR9wiJYMoi0PZ3iMiQtY
LfZ/7fTIrdAFefuNA7Ia93IStWd8OtJ4H6RnLK+u5X2rDQYLOTY6k9uPboQZ1Z9t
tZk5uEF6s+vtdiRkwssELJW7uW/lPml07SdVasff2ZYNehkQcD/FIXwjjQ96L98L
vo++Q8xMm3NGh/4DkpcEnpMtVoner6JUteX1LaR/sXg+Yev8ZhfwagZP3bjYE3NG
EUuufoATQqpdJTH+k0KHCV06WDlE3ROsi8Zywdf7QQWrw1dh1AwZaDGZgGT0M2PF
TWj/GK+zxFxZlpt1HXTTpOwZVUhoodyGUUUHCj17/j/EUutEEDK1SUWUFO+Bv7ri
LDMeaHd0KMeYhJXerSj8vgOQAuqBYs+aC8wwc5ioY1PlyP3MBHO2WG4V9cS53qxi
mVidcZZpbCgt8yeVrtd1lD622BbmHiOwNYCrB5BLKwZPGMlk4O9uFRzlLKWpOGhI
XFrRglYitrAzGf543F838RTLQvxtuAWkzqygWLzxE/ruzlNWONLu99QV0CBtZFOk
K2Vy9QSWhFYcv2+50PpzL/UD/wU/LVeypv2+mYADiYZGLDmte8KzS9nQmOW8fmI6
6V5MJtr1qczEdv6skAMATdITV1TS/bCVTGN9F4b97O/rQHptqLl1NeTVEAktDTHd
YY9/M0Qd+c5cJVKRb8hrxBW+RH7jbRg+ymFqHse69rQjugZbWw3J2dvkl+nfB2FZ
/Dd1xs4ZsvxTTyEgNnRDZTESywesOStG+IDgL+IfQi8khR/hk/R9SOpaaOsqZslF
/MfBo4n7eAUhdxAxAGFsK70e6LwUcHHVkzF+cnibeMRcdYgeNCp0/vsa2ubOe5t/
49219jh/5/4tv9BhBd6AF261d07z8WHw4BJNuVYXhV8BiZcPccMd8JwhfJaoKYQ5
k5wKGOQa6HApPDBLR9UGZwVpK2SZdkQ/AanrPW0Bxn6CEAwnpsOpGCmHfYY20b2D
0A39oD1VIazs95JedzKdsIKHvPqtjivrjf6w9NqbEP74r55TN1OGkn71hwqre46o
txHvrAp2M1KSq3MVlfQTkAEDUIJyBiSU6e0TWjObOQlAisAQig30IzYKPbj0GstX
LOqVuda1LX8aLz56+qqo8bUSxr+PS36XJYeBulYudCBiFOn5Q5A41tWY/HNRNvZB
zeumyE0OTipnvwbXH9+PnkjYQc6fBL3CM5pV+vVQY10x5cZrnGKLeUeoWjjQtxLg
akqwybu5Ix+9xGPjbF3UxhAcowtOb29WZaSsXXCWX6bL1rV4/Gc+/3mGIW2QUAh7
gGlIG1KCZnhmxuG6GGW5xv5omsM4xG/RwvbsXtJi5j0sNU2owscHRwDUn8vpvfEN
O9OBDZ5K3hupAx4BWoqYCPzL+XyrT6pJKlu/wpnr2FLrjdZLnYzcqjZcXcz8Rz2n
0dBB3KZ45A2r1iMDOJU7Aa4GhhM6zxpsSC7saWJLQBnPvJaeXjedIjXwdzyDe+gW
LfXWw1aVD6UQkwHWgpMVpJsTli/GUthxOqxT4PycNYY=
`protect END_PROTECTED
