`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hmwZBWJedsnt2g04l0tiSGHsmFBoIA0hyRzkV0ygp/uuBRCigwvk5bIEJs7IbQBw
wv+q6+XrIyXVQGPbRLid85hFwm6axaIo2mnQnBIQRK3eM0GrnJd6UlfFMbb/xJsf
ioviYRt9LNYiHvEbrF/080iQ3CCZsoNEWxMTekfveLgEixMbs04IGSQ2g5ZfqAVY
UbKEoGWCAjR8uG3ZAEAG16GvPhYCH0dxHoHM+vQVPugPe6g4ed6K2dpwmoGQi57Y
ISYKVMaVT4vzAnf7ULl9NYmOJarfOM+5DbL/VFeYxLAA0K6zlNlmZ4KUlatYaJZJ
OD87thu+jgmDVEasGQXsjGJ+oGzj4m42I/UGjRsERiay75epYilUeJWpnngRxZQN
sKGSlSuU2IO5zkGltewynHpl/jmGgTENBOvG16++Cbwoslw+Jea/5pU7WbXjQ34R
`protect END_PROTECTED
