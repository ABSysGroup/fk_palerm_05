`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y8LRRilfHPFd/FG8j7nRmr2cyQj0+r8Jr0/fl6oyF8Cv1kgiUfWMadsb8tKeczLh
OQldkiAnLTTl3wsQi/T93D9SUqn22r7ZOhus4MRisWNk7x1p7etxrUodgceEKUz4
+YHbjcuLTNlAk48alAHNlfS67/TGlaBiRp/HXgmsO+LhZvkNWMLEZEhAnzyEwcc7
DU9uFRfCXh9jeK83H6f73wLDBm00VL+xiMtnyTyD4zJkoiEkvGMc4NMFVE4X6B1W
hgMLpOAQjKl0g23cgX0eD6LkLOOckRoKwUlk+OxMPiYxO3BC8eH9X/S+X2J4Q+h9
dqjdK+m2S/ratEE/kei1G2+mUtxgYS33dBuri1pndelF0m77mFXC6SiCyUDQW7Vj
qdbdNkbGCNJNJOy9WbniSH6unVYOSRJ0PodEe6PGVUWM0zEd98Oqs5pZcl0VtBwf
s3webiRcd4GGVjBXv2QPqV58E0a1GWGnHJvCQxusS4xXserS4S5UaY60Xmy9ZAHT
fp9RLAdMWJxTXpftFw4HNgLXqSoFnQWyzzY4b3ODrTti5FQ4loNL+iRxi3+/iSiy
mcnaoojIAQTjqZLvtQas0HtceNpiiQ6zfJzyBafrODYz1x1vJUdjvjU6YgGwvKNf
wabjq61XASAsZs6H+8H6xsKUKRDiUy6Kefpp7isAkP7A/gQ4hSLn0AF8XxbCfdbv
qevj/m9vxR13fXxWzKMhAjcAK7GioANVcXhZJ2DNIdg95acd/92P15Tg7+u1cDbj
dwBvjKiz8aoNgGws+YfGDF2SiD3wukdpZ1xa3JOtfpBONVoLzRiozw3aUgsPqGMc
fmF+OtKki0BzVK5DHCdd1JfaZKEfLw1fbXN3eStXa+Z7OTxyEVEygo7op1XiJxOe
lHfgC/LtC4QWBaEq5N//Ov+2QqGto5lgQLX2aBsRqWcskRpgIPv2PNfsgbugzq+O
PzPTB+AuNqDQ/JQ8/Ua2jS9zCFRQ/9HZ3EAuM+aXIQqIQiYqJ23NZhempFnPZNb7
LYQ+MHK0+mIfKZ3c0rw6GbP6FOqI3KBmxWhKGWMnPkPC9dOqxgSFWhD9bCCgJrls
yWeTd8uTz8PXFI9vEt2Ruq80fS18iJTtquKoMRpH75Xq6HxqaRkiNmBqUpMKXK+j
lwY37buhioErloDUfQZx8VunVjdhAIbozta1P/6Md1NEOANTnXkEecyJzktSGRik
+MvudVgJvQOT1mFBBfIhnVqvbzGMCwlNJEIfQ/3PdFwNUq+Qr5pfMk1SXewJEJSv
78+rPo6HCSj7qUcUc0+Wspg/rtRFo02svITonU2rbwRCtSNJ6/6wU/kqX74fEpMz
5LfURKq5XlmMStEjgSEnBauNFjaaeX3CuCIVUN9lcCn2tTYHo9DQct+DTAgRCzy8
WGJ5x3A7GOI3GsfrY/awhoJyloP8K7uhjSwCvaJEscdnhkKVITCfPNGbP7qv7Iny
M3dEaVIzaLyr6RhvTogouEOxil50UvveDGJiTSfjeU+2Da0bPehCQGNCeiHIpDAl
AC2dieieXi+z8spDszn+jlQokpQuGx0PcV0ohyebgTi2fO7L76d0I6o+oR7P494x
yjP3IujzuSXAfzP/QqVqaqEKWUqURi3yS/0zPN/gTMGc7ANKYRUbK4JkCo+5TG8u
lLbwRqIQR9vKeJPLyqJxhgVhPO0nveDP5Su9yFzoocc49+C03vf3r0em7EJiPf7L
wX0V5z13/rsWrDx07I68pWxV4OcGte0V9m6NlRdsN9UeyLe2IuNSW8nY7tGH4iv8
JUGEJxyVN6pxitIEMZvfoOL3/HGEw+GIoJTqrkXJ1w352Q++hgGv3K4NpBkUJGgB
ZYY4dgNVzFndrnA3QILAM17gOvhIyuqLcek+JWHx+iBx97i3HeVgktrFn7nnVcbz
Pa8oCTrFWDouN/7BfvuHGE/tm0SWXFx++AzALrI5ltfPsBhVcfWwWuLpEqYMVxvI
uwhVrlL7C/aJhyP2QR/eGVQlPplKYxHMg24zJ2sDZVvhEdHRv6Y7HSI/luQmnC5b
S9ycBKfeDGRWUP0UvT98iCN4AgowhrvB2CobVzzTAyGM8Ee0KGnrVfXiFi+SvUnt
vgvKAsyn3PRnvYaIUWtjCk3eFEjlTNODRJX7YCFHGt6E2RIRT8wJscMTae2M7j0g
7wNsD0oAPaFa4Fp9PYo7pvajjRa0LwjkaQVGfuMeW+kJ+ZmyrLD8YYaRVDjn0/Ue
qqfpyNeuCRl5u7KtBF98xkBhhKfjYiT+emqae5LBQUxzaC01IIacj2iItxg9ctFr
57tyZJuEQsnFkGchxIB6fyqc3k4cgP3XCfX7hjiQQdTy4/XhE5l+xg827M3T1TM7
RfohQhtNJ9YxxGKk6PM3wCshNSHkqczIP6ez9xUeXsLgt8M5Mle4ALEF4rZEXJcj
atZXHi+e22eLIOjPRl8cURkwxXpuXSesTGXSDckhRRxC66JT6JkZbawKelZSSdxw
jWsaPzYN01ca6/LyFn9/KRFalVxQEfWlILL74+UNp0gntm09+LrGaBv1nv45yOKv
dBxiOAISfk92i65U8YWYNLJ2GcTbF+s0nhjDxI5rBUtA4nfvqnRkvNgZQTy2vksJ
nqdydo5lFtzgpYY1h+rNWTE4dD7+6xKuLb4+f3Py8n7toCOkjlULCWQWQ0Dy3YUH
zXwWll2Mi+w+XD9E+pql73eGAXLDCA6X9An9i+J1CU9yk4IWy0pCGjOn5KXuPgID
mDH/uMp3Qv61XPNWK2xStVT6znNqMbjwO0LE+izGpjhRi2gyBMKyHI/UdXO4jbbS
XAV3KQyus++QtL+9apL+Xd8ZA450ptwEImh3q+NVk9evJkN+HmrY3SqBvLfF/bGI
mFNSae7E3JWI2z0JfzpcnL9hdOC9AThMTVAu0fAkbWJt1Ev2JOc4uosTFig2IMb0
CY6+fmB961Gl4Q1pUQgN5IoDC1cIFeoxF+qrYwxOhTyktLJYwxBBSuz70pSofohv
4OKWGm9yexRcSYePBlitTuFmTl4PzSWf2YJU+1/BKKD5zK8vVDufM7b/RzHMGyq0
/zlRoyrMdjskM+xUd+tEXNayydU/PQrLQds+2Bv7vp33RB0NODv/PyOXdiRpTTVB
cHlbFXRga/dRfkQuMeHOFnz+5kxre81sqtzKg4P/XGt8zK6Lt0E4gyDF9yHd7wh1
jfWvaV+js0U5Jua1UlA57pWKCqTY+ZsbTvBVfpKy5rGHqWlA9tuHcK9nwpxqnVkj
I+mqNe2cmy/DLKNi+YwP3pZCulmBltGkVEeXh/Ub+7ZHsv0virfiM56gUAIcDRHs
afs17Fh5QzFYrs6+slhexqgT3OT0dNHakGju6mpgl3EQWgCfTB3Q6GqJ6DFqS8JR
2Yc/217vGNj79ixHZQmtEcRFo3bLzmLa6TM+CLlo7W2cdw0fG0hykQA1SHs5nQU9
e7yj+iWqtUZ6pKoD1Hu9jPqHr1HT5br2//pGVD3Q9mBSMSoV0t4uEHiDL+M+HNwf
z7ChHd2zwZ7nKCQVlVhM333/GPl+i5PTCumVa5dkN+++JtYJLlMSrJRpjZmsKn0j
AkJstSkzRohkRKxZ7wxBr7wb6nCOUwqEnruSdpus3g40OYTRXWLD632VhvbjtTru
7KFFqN+qBpru//S/5RQuUpiTfdo6oac+1cN27vpPQnsLYr2OZ+AjoFeTb/Yl6gkf
BFr0hGRxs/W5uLlX3KO1onRIgoGAfJN0gAHa5zg06P5HDQ0ggMIElnW+7ktOmk9U
KI0Puf3VJP8zN3SRnp6BrxmD/I/dx31jXh+KUzhImhNUNZ1GgJusBc41CA7DlcSW
ZMS42hC8pnqLB/+Dfe4/o/RJgv1clN/1xgcc2hwy9rl0wJhWZGDAHqsfb6EXaPYY
tTcibGwMuLljAmzlB9dbD4hhUULZiN/dS9pyoYvxDmHNW9C0sC8G2WFmOi1y63ks
lZ29ym+U15XtJiCSKGI4wtVvY7tI+qK9FyU7Ytj7oiqTGWHZKBki4shehs3liIxf
cYqY9BUv5xfalJQat1f9gP/EQi8Yziysyj7KPr9S2m6V2HdjAP2ZmAY47xC6q4n1
kWjcqPHAY1MyGDRnc57hMy3VS1jPySmPMlwBEtN/Cu+e8Iusz/Fckd/46Y9RCUut
aRBlpUAS1QFxhBhblOzrtk/Q1Wox0vBilwJypp3ouU2cQbVudzo0RDdr47ZBxJyN
lJghgcbmbhsF+ZcbUnORaKVeQcPOGeEuo1y/WyO8qwy9VfzYaYazPNLX65FpoghN
+o2B5WzRA8/muIA0Wzkck8O5NWAna+LmlzyyN6F6uXj2X0Vr5zfX6qjd33JedUAJ
pYfDrEvL+cDyVsnVmYo1ICGVn7vRnCqixhPXjeInIHfbtl1Kndxr0nPwfmhG4t14
o4b5ZdZx86x0ulfgN0LDA8n7T/w3gu11ajdi9eRdtBjHXh+zZwTp/JG76sS7CRvi
xd3NygdFuDYyI23WKw7kHXZxS+iZudNm5ciZmTRMEsybJAKuNjFdmHFdtfpDywBk
nArD61km+5p0L6eIIX9e79EwQnNOYdAyMLQ2eyoUVjKGnNEYjuQQ2Bg3RlPExHE7
I2Vr8/kqN7Ecl8Nkpamvbuq7Hcw+nkmg0re48a1u5ExTx9BV6ueYlRMUst6WfuAE
faxXyFF9D/elYHz9gkx30IRG3EYGgltaxG/F035TbhedgGoOKcYmdZYFUIuiAHf9
DXyFtfkFjXT4eBU2u/35JhuLiMU25grrpdKtXuA0oqmRjH2kJI0gyzLBmoHzDjXg
UXbeRgOFi8y/hqRxKTEnMpNb+UekczzFR0V0r2c95/xrjJcKjKnfRRJixBAN6ecc
x1VkSaf7s7ilZBN9nVC48q6/kGAzV0k2Kos+5ZCuP10fhPyWmMmtAxDNpT4gcuHq
MjkkUp9v95eF4e/ow7fZNGYNX5PMkg05AN+XGSds1rlYjg8FOEvnb6nnwjKzMPUY
3dIk4Dar/TCAWtGsX6vbWxPDJnXh/dM0VV4JDoY7viSmooZ2BhDFwbfnVne2GDqf
ef1SoL7UTdkD5dUJ1XtEzgPdl6zE1Jj3QNP91aM7/O6V+OhieJjoLMIoK61UxDvO
`protect END_PROTECTED
