`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JNElaRfP6MIPhM/62CM/ZGTNOpBZM2MnGp/IOWRL0Sb/bUNfpCmliokF0f+aupXg
ueUneZWx0LhipAa6O3kDryDMOJMIf78pbhZ6Xe15Doo6/YNiw3UqZ63qQc08DJZj
cejwoWByHV32FcjTrZMiqJVjDFlpz5U82VNWTMm3K6FwlUhmHG4zmpsL/MPScz9J
gb3z03Z02DP9ZxEM7XtyAhMdvzO83rnVv9tQppM48WdhnHEeEZLLj9i3kHx6beXx
+2nE6QN9z5RRuqc6+sxWYB+eBtO6SVneZQR7rFVqB8ewdjTlvIFgV9FmSUU0UWCq
7G4SLshZpo9PO9u7DT6UcMwlLJqsatKOw/zXYoA2PHKafKAI7l/PzTN/TVjSNTaV
rxK2EOM5E6tZ75YnAjoGdeAMsDP0pE6dlrA0K+2XZuiXzQZIf2+wqu0V0TGLIiA8
QG2NQwX9jfTTgitOrWCeegt/7TodvgC0qFpr1hRK5HS0KACGuXuvzsbUhsIOvTuk
Ku9QqIzGocbkxe1bpvXMan5pXtdhv0gVkuCfQVgaQdsQQQav/jskKWvO2uiEk5HV
RSpJW6fSxxVCRlrH/fxg5m6T6tMyxAuhUuK+NlpxcfBWcU9/cTOL1SR75IFZ024k
lk/3fi2LLdzB2LA7L6zUfVnkjl3w9jT93cjQS3LxxvsSvJ+7ZJxf8nlAgks0mH6c
AqNvc+NIvIQo8mtq9gUKKkgdiyZFfVrqe9j2bg4yOWJgt2jw8UFL81JYtF+BYBeQ
jeb1qVJPt5T86bk2eRmSRMV9PsNRbBmt+dI9nGPi+33WY06vBQj/sfMriqrr/FxQ
alN8BV6WBnJrhuRSjOBsK9guGbdWASiLKfE/+OGQcqWXq2ujVPV6rFKf1K4/8yTA
nGiY/llnsVB/dA4bxxuqHtEHMRYnjJLsztrRFjdcKDnK8/iksUzqhhIq/qPDLKWG
ANFphbJXl4/DY1dsPcw10TZEdtYbCCYK8lthbpms67oOMHxPdHOK/GU1LKG27+cs
`protect END_PROTECTED
