`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m6eqhu8aIY6IkRJ7uhyGfT3IBHsUKH9VyTHPbi+vsFEPWaUWHI5h7TGHxqSuaBKI
TXa65dqNcWHfXPg9QTAujp2GAP0ocLBf2EXZdmcDOAZq8EaedkkVR6BAitl41H0V
p8n8oD1izFsQvrVcyUYQ//MEI3n7g4WbDlgwbNDhYWtipthE9jSYY9HkGCY5zKmA
436sb12m2AcIajpmIHSFH4jtMe7CoNx6PMcEVEueKq3azVkA24571+/M1ptIg2iy
GaMnZgIv/hJDy+tU6TIRFyIPpDaPFmPHTHpBRD9oz2bYVN6ejfsZ+Y6FUkckuyj5
YzMxlY0hsJeYd+n6aO8V9Ldb0xqqZD2XjMmfX0brTdo1JARqY1yms94uXZ3mV9dV
d8RdyENW4ANVNPsBGCRG66Xsk3CgEirlIW177F4NhazK53xTvE4poEQtoVZqEFs8
yUxftLKy4EuqeAYPH/Y7dVeH+0wagnCiJFLx4D2h5AmfoMnD/2+1SbwnPK3FLwDZ
f/NtzcGw9KmStEvoUQsrAZ7Df+45owyKdGSO5hEDf9ZBP62PizOWC7MXr/EuEaiO
5zOvmmDDQDkq9nLhTecIqFVqxY1uTUjUt/vlkr0rfxHAbeW7bjd52wz4Gtl/Oanr
1BRC9o4f5n789/EGl/dbhKM4imrTmV+FmkUIpqiH16yLiQ647T5UQNMvu0Oiif90
JWeMW7qjG8DzQeFChaZ3UDJZDzhCw9JdGpQ+b6dZ2idhaAO2h40a3m2v+G2T/GOB
UhbsTCYKx/D7pYO5ttEP2w==
`protect END_PROTECTED
