`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AzPOfYJfxf7zKjXVlrcNMX2aKkr5d0hafNO767LdtBIvYr72pT5ONgk/zxaQUq5z
Ls9TovmEFtTLZ2mkQKQk4mIVDpXQlPwNUKBDCOQNq2Zu9ompEvOi/b9ashMmIL+H
0Z0tX8IPstHtCtlua/X+Ymn6bGBhlldZJwSLK39Xrds3g4y4b3/AmvYa1mPGh3+u
ZEeZacAllYuCefBjavXjPE3f15WdBNCIEyGLN+7p9LDpKsqItc/Deg4mI4+OTfxL
2WzpnBh8VB89I4TulqU01qaIa2SpNMR2gxguElfojf0DUselbVFq+/j0VYbuzW6y
vIKUey4gbFzUG1GU09v+Ltm1xd33M+qFkeZlAMAz/A1UxUCZyUqIrvVTznv0W2+N
xWkBTcNoAc0rTAHsxlZdi6pSiYTecE1iZ+HOYsATgiqx1WJ0ZMPa5UAM/FSIS8OY
8atS2EtQl5oRyPsBEV51QKMH3TeFG5bKf74JSV1D4ElRpcEHbknfFk1fUi/a1DH+
PlcS01V0HtoUr6SMjFrewJAdcIc4biysjXRFOjZJh5Q8k/0I0B3t779wMmyui97o
RyFAX6NPHzCMN/tICRMOwzFNdhyehpDOzCCVY7gYU4jgrQM0f6vM0mxvYmonjo7G
hv1Gk2vskN5WlYx9LqPYVv/AaSqy6Cy6ZVFxJ8RRZmeVlK18YpORGiXlXjW1onGK
M8LJSJ8YP6skOrI1WYGolhdhYnjPo+rRG/LiK0p3ZrYscv2+Mg4wBf4J3uXqfysj
/TisRiCovaewzN5P6aS5LbRmDff8KGsdmiAXVcLZRSjcVe+/uifemNKg4kZcUduG
dCXYaNgfhO7hdvjFf6C8vZ3pYmIShvk60D5+3YRvijPy5Pra+EF7b8NDKYZbOAbu
GHgIU0exgxohBeD2rnLeohu3VsZYODHkZbXyyw4gzNGJYYWBRcVhQBTVS7bWX+Zo
`protect END_PROTECTED
