`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
se5Bq3d24XSgONvhkIrHO6C+pNrmta5J1FeiDjyFJeYn9Iit4deTk1+j+FH0N/Bc
lkolXAktOKdbxV2mdv2oR8F9LZL5qgO6w4GJRKo3nLkKAh6oNMSVdCQsupEjcuYz
Dpwq59dJNxDIo4SplqWcyouXzmcimWuJNnC+7VNEXDkg/2S/tzwTCIjh2F8QCM+Y
qLb00iQe5pxbDgfbiSRiM/3b7K689FQ8Xp7dWBqRrOCCcb7GWahPBd6+w/wvrhPA
OAyrzAKo0mxMWz2FQYb1JEgpx6wkc0cvZH3CeAsvpQwJoYELEolRbprCb4wdXNCM
vMpSEobrnIdMKkVLVa34sg==
`protect END_PROTECTED
