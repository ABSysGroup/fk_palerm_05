`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PXsIkNv9WM/ak/Vy7iUQNiFfR5ZGSaWVMZQB4M/COdep4r/QMUzYBwMC8elYFAVD
dlFb1K3Xzy/DQRQnIbbBnWKwEqQizuoz2UyvjqdBOk9tym3YvGlTjTxenf79+z5c
gzBB2cu0QCHNz4zmRPgR3Vw8ELx3F8hYrasrv1elJFWlkEIS/vVYzSjdkgIn+kh/
/NLexdbG2pTSgYkucds3EuZB44yXCd7yPfW5vDUQwfF1++Smm+OBHVi/xXevW57E
I/+kmAZu4AUubmVYNNy2NxGfMbXEcbeIA854ozwd6PtvmlK4o+mjUiLhq7JqTrgn
LPD+m9WoWNET3kbtWLLsb8XX0bXHCoDvE6qPyICzveIQwMmHlll89ZIPE5E4wL/H
R+qifkIcJpqgsEiR9c7fGjlmsCDiQPR6+0eZleYu99qPigvTPwwP6ve5uNlQlCsr
mcHOB6jqNYFFSqnKP7GxvFXk7aI0AY7tEY+RzZP4hF7mX0M36PHtEKnxQ6sqkO8n
`protect END_PROTECTED
