`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jueUWEq00mMHSuFMN0QwpO0dwyfjmhRULwvrjdrKs+DAQezd1Mp91L46ziZsNhBF
AfkEd/xBQtcJjjUaHd25tR0dWmdqocnnFMdMROWkDsd0qW3d/OpeLE1Jiot7HHxa
5vI1gPHkn7FVS4KPU2Am31WCnVKif/sfgK8NQj3QCwam8IxAc9e38urLvLVZw1wc
+QExqv6cmsuCGGS8k6mtjHlUNB46uCnm1KikWRnApYspVqPieS4I0swPe5Wp/Q8k
VkxgdNPmFPPumUtZcaSZ1SDEHsKRUP3hQA62jvREFViWvJRsgRw5/1Ys8D1ydBQl
1uRyM9rw0UfAe+Fn4WmYZxe+ksMHjteWHQ9lER7zs7ISHBQM/W9JSyg04IN65w3V
SUo2kDTEKKgMyGop6I2kT4eEbDUdfIEl7zD1Yn/9oxJyelenjCplHqSm94afTxL4
SUPj6WS0TdHwUTKwLfR3WgCIVP9AUWQYxamdI5RMR99BP2yQE4A1XfCZaoZ/CgMi
RQXbD9SYYTfxMU7dso/HrBxoIjh+NagKkNfZtVHNhWsRQHG4zTPvbTxA+qZHMd8R
1acAwX7z7SNmNItPUqqWiEeR+wFTLyWBqW9nQC/ttisabImQXW4W+BQtrYjcgZ+J
hAPv7Bup2kDKNXxHz8PNczv5A5wLjaYsJoIZlZUvOtkdjTtpPs18Mj5DJ1fuoh76
ZkjCAhOdFPMQZYxu2s91aZGWa9mKk3qScHP9dIzj+2oETuNj4Dv0EHdSot2yEuB1
BrNIjmRvgJyWNlOj+e+t2w==
`protect END_PROTECTED
