`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X1ZbCZubVeCiC8F+fmad4rC/JiJhY8SXKitWezcb5eMhJF/7Q/0UeLMrPc1yqyJO
gkuECeAztATiiIgRu+Gzc6UkehEup/5TUzz+CsoyY2y/F24l25iEB86XQecrWDk8
l6vA3b2n1RwXMJn/bISyj6VZ3BTHhbhy4taFEf4I9wn5/Gr6+K7584twt7u3DWuO
gJtcsZKEswKx/hkrhcGMbgMZkqcae9sqU0ZiBc4VWGcsWzab8kSduG5Ce1nXz8n/
eAxPTLNKPZggV7TZcSzG0w==
`protect END_PROTECTED
