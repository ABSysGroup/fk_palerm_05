`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
obLqsFB0ZgIaBvno2j3piWaf79kVHlR2DpNtvF8+DZbIo/tnq5R1k/AdbbqMCtvf
RFkdzu/jsTNZKflcjmY69LYk4iYA++cRsKXp+03SNgTQDmRrHt+FL4K/TZakslbS
aygvR+K/Y7Xa2GdoyAjzMj03NrulczFD3pPwOSSluPWTjzpK+LsnrQ8LPZpPrqeN
p476C4XnKYbryFN4zLQxG85LlBEJFQGqD/UQXeSk8UQ6aUpI/wQaO4V+0Bo1YbEs
FHVEOnPEz3RIyB7C8rQqPa8s+WO8VAVHnzM7EGiidDCCqgJA0BV7itfxihcz9BrY
nATETXvaduFfmU/C7k45BA==
`protect END_PROTECTED
