`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pcFjgwKyLehsM4cFlDCX861jH9SwiMu8Ctq4gtOghaOTNALr9MF6nJX5OZMt0gYv
WcZGm2TgqIMD1OTO7vLzQrylICwn41tMUUPQVVD0dFPbqMDFXjKb0lxqzPJYyvZy
pLGLju9mJnxgo/rwO4Baaz8GW3NIXCmwRopUN8RxsrOOmrVJH9sXWoHut6bdFTkE
9OAViH7Qmzwg46OI8lVX81hbhDghh+IiXSGGB0Gw43Hb6o514nr9Q9esdRaiIDtm
/QNuh7jEvr7KXQpnck+YbAQWuziQBD9OPIaqvgW7G8Z2RJJmJDseD/UNqNjFEdvu
A9qHZ9OFhkpsjBpL/a+Kn5UBCIIuaMCyDBAMqh1GWp3xDDDxi0aPUZAZoGoG5hTJ
BIAg2zNhAlkgpY8nuuKTHxfF0zOB0UCdoqyDmHuymfUg48eLSRLLFB3GNJsTWWWM
Gz5XcA5PE4b2vQBbxymJhTq+GXYtbZ0op8IU0EJbGRybzM0XvJ5wC81A9+TSrlwB
XZgUNo4GyxMW//A9e7GsN8e2Dit6XZ/ybHEKgwev53cT5XZR5VEmbm2yA7uUENbS
PTFIMSWo09o3e9cGOzS++p9GOBKAajD2ZMWeIUwqkBI=
`protect END_PROTECTED
