`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VB02VcVq8UQmXLT8aPBU6PmjdJeE4EaYOMvEdSEvqouFQrM1Vnz09pDna4u+auo9
0daKUcqNl6aQeK79aflGPhid8bMoAcd1LDzr000Cc+WEC8OJ+BWT/UuB3taverwU
AyB45hj8QVBT1PqtXJmixDDpvxi5aRBCH/ojQ93qVSb44+snJR+lE0pGxCSyV41k
Vx5VWgydd2N+Pg6Y8+iVijvVHD04SUzJ4nxB0l6IaxR/voP7zX+WMzbB5d2JrdHl
Zwgx3WKV8PT+9e6/J5i1q+mJ2vAuggjGI33RmGi9CFz+zZ7qTQ1WUiN9wKl3BEnv
xcXRVbNiy6v+bPoOZx2qT9chLR7pIy6NcJaz5CzvC9Fdpu3CLqEwvz6R89fp/dVQ
/K6DZaXD7lERzotRmL5C2XlZIGa1fAuCJ+dm9pSKgJOaGQTWJzNuGzkG/IlCuey9
rCTdJtV6rcNSiY+br/OTb94DVTu4uVMYDUof2Wn9T3XraY1MBhrmlUMd1N0js+ef
oJrLAZke5rgHUnQC+jce6K1T9g2CEY/kLCRfJ6254tUcDoLtu2r1guiGcYmp2hYe
rKlwCbwiyv9wETz/RX6zyahOQ03n/C72tT69KJi7G1IRsXBcvP3ywWb26Z5iVlfl
RzVq+cJ3Tz8Wyt3PVfL/277j+RMa5HUzu/yt33K0Rno=
`protect END_PROTECTED
