`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g/LBOLbuNVV8TS9SkHoSpxd5m5q+8CyfMNvvK3oexpV/kVUSlI0wLJHip5c2YYYP
mQlqEpAmqeKg+ONBDe/55fUwA4MQqCbclwrfN1i/plYFYaC8C5cma2C3Z4y4oqEx
tKOW1hugw5W4MezGJj3ozlFCcxvgEZFb0L0wcQRL5DZaApqnuS95tbk8R168pkY+
yIrdJiPi94fH2oH1bCbHYBkyzf6oxV588bn2oMUITu2VZsYpfG7yMW4WYSDFHZN8
9qg+E7+fGxU1TwPi0JCzCSpVaFtwDV/zuXkqXlEe+OvrrRuW59GWs1kmygKl0Jvj
1ie3Jej5NdAnT+9kx3U6+/MgJmcZoeIZiDY5SAASIlACVg7+DM0dJ2FlOGeczb6Q
GM/fmGiSZ3QZcM7VKWXeew==
`protect END_PROTECTED
