`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7h+7+MqFL6YdYC5LOOBhuAj3znTHNF8X8Vr48lW44Pzfi/OrGWCEmb6YKnhzC1Fk
iCCNd0E0ulk0A9XfMKDgyJoHYLi5sL0REYxhFYXfSGoGcjlH8ctSeL332ZSTFEUZ
bqJtKttu95g0ANrc9h9OBr6hiVkDGMI6tcn6ZtcX9WWf7MK2b95X15Fk9/+W7ZSG
OJh6RMjMW2wf9kMGyNL+9em7dYoX4vCVV2/uVzsb8i91wtW2NXuNdertkOy0phSd
A+L4eBIs/iCnBbwrAAv8EvcveBcyoz2O1A8mIyi09+NffEZcBk+i3Xu809P4bNZc
pCrcanWDdqHXpz7i43RgmGFnwh8foAUJEqnT7XttMDuykXkTYu+qo3BeYtqKfg1J
L84mOX1caoUNa4AB+0xlLfgOOJBDDikwR2DJ3MDEFteexdXtzzCUARBzC5EN8qjU
Jwo2ux4I5VpI2kLnFPKw0HuSEmyGNMZ7bQNcWDOFEi7JK6+LrEA+w/p0PZlYvPh5
LS60i65BAOzs2LSdcSjwjMEEu35882oqqihsUSDMqEArRWzP3bnAHUNhkEojSSpv
UA/8HuDIYN2nHXf8iXfEYHMRjd7tGecPOqXhfZZ7n6wtK8l8jXokaXjFlKSIEfDN
WxoiyMVgnTTRO0t8M9I3r6OVBOSUtGt6XKGV3z6kSQvfpEADTIIF7Y9vU5MgYU71
8e2xQYTXyG+ufhVq0hY3NE0wkuLOFpCNHF2IYl7Yv53QPvYhFqu6lkj8fdTfgHmy
TjTPlg/W1aZOUieNrh4bSTe2NxlMPNTv6B3bN9NKWdq/8yVTwGaesBow3plpSNwF
2tqA6SK8bWtxoSRPNgGyHnZwyGtcp8HusAilLZPHv7ZmJ6+EaZR6/HgXW6m67jlR
1vfRsothVIu8ne5g1ajYa5Rjnq6Xst03tUbeSjsAd4f52yQoD2ijsTKJLvLDnsUR
PirY3bm3eC5cEcy2FkMreGmmxmXp7NlpRu1z5+BEnQcL6eN+rD2/7M4KJ8Q2nn6F
Sph60nZHgzUqoThLTohGWDUGska9MPw45Dq0rMoqvP83wWZINH8gw5sbsdNHXMkg
J1f5mNC5UfCIowUlUlFMijOISJaN2IFR73DlTkeuRbaEaOSzm0SKaYsbqMBrG0T9
WbuKzJvxhXqup8SDjVpI9np8s7XDCoTw3jlKENpkkXqBxFeonEa4kk4rMDzykvs+
m/QQCN+boqqfEAVpTMlJks31eeZfihCCFP6vpCYiVKu12Sk4uWi9IPe66qyygVtJ
LI4r27dDkBHW3/LkhL4Iz0/Ql3NdIC2Ez2wBPEUC08aDoNltCuR7TE9PsJuweHur
+G4zUiu8v4ZD7x7cWWqEgiAIVDRUZXQ4ndRild7+MGpHO7PgAi7ZoYT9sTJ7bQyT
nMv+iPy1RF48gTR3XRkX/qWEIcLWXUT1PJJq4725qYxzOwpQ2zZmOK6hBsXqyY3t
H6Vc8qBnl3pgVcy2q7pxs3Kfgvv+hSXikeaMd6S7Wb5xI/YtPOvFb6HKj/9u3Lb1
VC660tQo+ScZeUyqa0TDglLXU1smM0zPdMBEHapj9WJr9x5KVKMHuVmZR+CPiIOO
Z8hHdFT375GVLlZF7byiGoLrx8Wxjr5x5mfieFM8axnWK36bvT5aMv8dYalOaIoC
rUnSntGTxUbMDzD0h6rNlciN/4pH/Vnnfqoq013cSbg8Aj6o7YQU0r2v7S2swXnR
XwOCjgtMd6BxjfaxNOSrLRQ9a7+Z8+uBooHpYZjRzTYr+5Md3i3t2enq1FmJzhTW
38TSw3GVgsmfBC2T8MuuPqo900Jz+dfSx0uxizvUE3SknRbUtgl1Gn4tXCfYFrBI
XnJpAe8f/4IuAy17Zl6V628SErt8XHsZCWsNWLT74Nf7LUeJ9PX7biY8ZklMyoYI
lt3FsL6aGJOa0/YgKnjM5cBHe9MASlrP8pDFJ1jN+0dhBILX1wg3Uq8871O32enk
YgGAoJGepMkAkjB0pX3NwbDpew1+urdFS7IjkeIFHGk+FmZLb0gPh/+tkj2cep3V
LSEHMYCzC0tGgp/pOpJTmIFrVjACucF3Rox5mKtdytD9u/HZQFaWKIPC93c+T1HO
X/L3WC2ZU1T8rmNji7HxcZCOFp+Ej1rSoeru0Qk2i1NIW5wCRc7O/Wm+QRmsp7Tu
6EmMyLdARy80YhLeIyAe2MGoI8N8zhZguHHubs5uBuyOwXs+1uNzfGialJmboY+v
2WjDpKs8PhAIhKTxgTolBOFWIr8yJe4+s4AFx6x8BhxDmL7SFOO0BjdDveIzMckq
GXLocZjSTI3oXh1loYkCsJqZUlQLL3uoWxz/IBkFRgE2WIZb1+69Tu9OhtKK9os4
YI93DrcrVYchlTvMZ/e40YQyn9UUlabMtBOVidn0DKjLDMYRJbvwyDH/SDE2rard
Rh4Nb5pNmbjgS8minTHKntFg8slpOZhztTorZjLJQsS/WjwGV/fVjs/RR3FXZXyd
BNrTM5EBdBVJx9BsPrDZFa6o1ykC/cEIpAjSNCiLFP0XGuOrxNLE5LXkYPfsV+pL
o9TNY+TIjM8JaCV1kPXtlWuiprSg+kSwUZMpu2jMxXRGoeCxf8ZifyBHHZb2/WYc
8lefAIfw//jT83FnyPSm7ZscYY+18zpDeYAcW4xkWDgnXOjR+9SXAyYFNaOriBKB
lTD8QiCvCxS/MZcgudU5bPbQqSrZfxtwGGbPvTRL7WCnm8gidh/GbnRq0jsNsZ8b
UKTLgwnjotdp6J+qrBTPZOeRwbFz4XwmluPV3t/qEDScowWNGV/Tg2cJtWOz1I4U
E7/t/cDA84rbQY/Jf0Ln+2adKySric4yR5tk//FxCRXgSKjMQlPBKPCDkboO8dk7
9uNx1CqpPn3QsxBGMj/ugXDlrSmpLGLkA1vMPXKeVWBiCU5LrPE2lGQSR1tqlSNX
Co/Ff6U6Ql3HafCef66x7NxymehTEwJUwQ6pjyNz6ot7ZDPHegKuZk4NY7AxpcEZ
0J6aobVSv0zR8Y3NBtR31g+zBtWUL0LXhHhy4OoXfTwl2Q+rKQq9P00gY4Rx/vRc
SA8gnujC9oOgt57AfRiaFxrAqZtvzqCXRcy9hKLENNVSnHFY0zBudUf0s0hGLWyc
Kz8/MvTXi5GEoFvmrt37fyaf5N6sSv3lWyOOMuXCC9Blx6cxrUmorRaNQmdPgusR
Q6RXB62bfnNUW1fW3H+r6RAP4lmlb7ZOVxbOFcFnuvFPTKxefb12qCLHFw2Q7kQu
IAcywaZKyMVP0Z6CHXzBrqVWeBBF/aRpN3UIcifN55B2dckefYNmyvqnmASEaYwS
X4rFhzvm+4QS/HKbkN82oDc8HpzPVOVPNMRkF0CwHM0j9kwSpcRVLtdyAS+hBkkO
GWV1G5JEnk25qWfpHtipV8xzgn6wYV3iePsD6+sYQs3nqjJREGbvQ4Dq4fuMFXgb
gn5xDKWlykgBN7yTk0ZsskpY8haLLkLOToVQhQmhXsTvMxxC9daAV7pUNyzClGPS
zFlIZ7dY6fjqLZhr6idGg0W32SXMRmdIZ55WyIeyi/ZeJXfuq5T0r76676DC2fWN
E2ef9CXqUdYhH+I2W4qi9OcoaBN6bi+fHAFsJOxDVjsBnHRIHwITZtNuOvEK5YEM
+Dp1UN0VqSzR8YKj38bKy6e8Pl4SU60PJN9AdR8hkY2oX/5t05LJXDd89Ko3jKfL
xAIwTNSqxGLXLcxARQC4Fl6vy8R0sptAuseFA41CyzR4dL3nBgpX2xf8EtQN00AD
Tr1LJNCVM1zXcG7dP/B6VmNKgiIB6blW9wtr2kgEg4wF0ljV/74WkGcRbiKmPDsM
UEJs/9CrGVUVEMcOV2DPZ9G/zoNzJ4fKFq7Nc/W0SYhMgjmczEhHWRxjrk7+Vk1S
+g/wB5YmRkyuXKYYQ7wHzuafaeOKm4H6rY0aabnWT2PfCZHndcOCKUYC72rinYZ1
jfXojhTIJFz8bgw9NZ4MEsNQtzprym/pdkUh5l3+oYPXnXLXyBIzFhLbL49Bc2iC
vWYiZiZzPiO5sEXbF57yqJ60CmFxqDEZ/9P046Wz6cb3aT5b+AG0AAwAioKOJKqW
hA5wzXWW8kF+ACmpJVfV5NaDSYu9z24dooOnerfiXPNDLMeAmCGpQsgO51rqe2tl
qOI26M4zxGnGP4cXUPVJE5vkJw5zYQg8VANLuy6+dGJnEQQtnGRecmNpebaOMaaH
dPtQH/tGzeXgdzeGEob192v8hYgkRJp0OhikmRAuNv1x7kaVQoU8hoTGFSCZ6nKt
`protect END_PROTECTED
