`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4dQyz3MVjpJiLZe2xF1zLZUWqElMIENdNFA0y0tIlZNuIxhkUI1x73DLGsX07er8
GOAbfo5g7J2XgrOBRw72oz5BWFUlfAEwOCxNbU+PdwCaI+J1bKboUXRLT/Q4IgZB
5Ws06Acm+Z3U0dxv/sxzgT6H4DQ2op1ygjLegsVWFRjAd0/jQzs65tzr425ftCph
2m4HMLtGry4aDBp3i/KNVPFI2tbzzlTeqF6OBVF1jA01o9+XvRH1kfw+YuRtx88c
S3S6hWnha09t7qE7r/9IvjW+9pjgSsWZ8xl77xB+HGmB3WwzamLgk9Y3+AvIBKf3
QTkx/f1GO6SVYY8BXCnPpLrTq5nbKeA0CHr9VTEaEzoYQwnOyWPSXXve5EnLiipD
1mk3d89CsDDQpzNUNlZbKLxY5rqREeDx0Ks5aT8xhS0kppZVXHcn/8G4h3FpsE1B
bTtMM4Vmnymmuyjx5BSpw0/q85vb3ICIVHTtGKYFiPw=
`protect END_PROTECTED
