`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vSMi6JNTXP8bYVPUNu3lAFj9j8+w7WPz9MlZEz0Nfndj+sRmYWCoc17+EUJ+wRQt
cuplWvzbU+V09BUWElBR9BtXxK2YnLvXa5joy0FKXR6gql4M88CXXN0UNApehjAB
bPZwaFAI/YLJoL0H0rPafwmv5IrOnBHO3uPms5Nis/BG8V+JjP/TtYPChdjj41qa
hPULWH49NXNSmN30i5GdY+hRkFS+u7ccCRhBeFf9tbg+2HjA7D/mSvZ70n3nVAlf
ZZ5LATE8lQCzqFLoLHVA0dgpP5V3RhCGvr6YaJ2W1mMgPu9t551G12bO7yFXmGZr
93zxttaywQ68QKlRimH6769CgOoj6shM/GAPdXohF1iSIZG/BbT2Ifiq0MEf4mHA
4nTmNBBAzxUmtHGuIRa9rm1hfAv/4MpK+xOrTBOFfDDQ7ooQqiJPkyRaZrCJOzwX
5L+RyGLgdxnnlu34LP+rLHXnMazEk72kB83VChgK8nOIthkt+tPzN02EE9UlrW21
Q2lEHx8TKRPm3xbWBBUT7ogGAdlz+91l5yQsIrxU2qh2Am+nZEzXJucj4we4bkbH
/Kfn/WYYwxZ7BBkvlqOiF04Otu3SHae6O+r9JPJwI6nqf9zcM+MWNu5vVTZcOva6
ngc5wBc8vdE2RDiGOw8haUjKpT7sZ5HsbvICUnQXW2j2KoFk9mIYo3YERGPhD5AG
00XDbNYtVegHRE8ljuxTd/yqbS9Xykqq+awUa/IPdU4ohI/x2JBNsKWfxn/sVxgr
cFjhXKP50+ODGBY/eCbG3KC7bAgZ9u9S8quVf7/qFvUw+xOTAXVl17QCt88tddtS
vyEXrfCvcuOlxPLO3wqzN919L/CXA3MfN3eexXB6uYivJrQ7VDVsTn9c5azh1xHH
HLf9n2SO2wjRfmVlMS5gIL2V9vZA1n1iKoNlNu4YRhlgNRCEGmDrDcwo29cfRnYX
+t3OSVzrOqJGvdLX3QYx5PbQK2GIhS92iGzoxBjnoTdJM9ELEYKYYljf7B2udgDY
G16bZMeaC/Zw+/GYnZT4/5UFKORQRQRg5N4GOFtCpZYRh0O61V4rnETaksIO7eul
I4Hc65Nky9q93rJq9TVeB2HVeaipVvn32OQjKRqPHMlJ2bkS7oSA0AYhck7liMpJ
CTNmIdytxOZMfBkbxtMJX+rtlB3rXxO6hwanwTvfYr3xzxV3dL12q5kJpb/ZgYqo
9knVjfmb3MvtockmlkGxyHqPN9yOkz5O3GQqtM+k7aRz1ZN/FRBVJeUneHMUxOp1
/zCcuYe6G2yOYJRwDEIyJktwXFLG3vYhJnXu6fZfFN7ddIvFJA37tb6ZGK4YEhfv
PpQlDcIG3Y2h6opd0C0hIK44u4Iec65N9DM5TJxo8rofq030VDhehMYekeXIOhih
wQksv0/UieWkdNRSv8D5HoZhj+k+EZTkpPHr72qfrASciNUqQK5KzzIdcYKH+NHP
FG9qDVADDlvpc/WxnVw5BpYHsf2gqMypOaWNwCLdq9oxaocnkn158m4Rqv1b3z3m
Rqxz3LTXhWvWa5bb4vdx6bpgXYaI1PXKh5fCVX1sQ7g0QRq3RQLwGmoS5EYgPX4E
EF1QwdTMYYYnCZyEbxJn5BiimKai/UiSKNOF1VF2x64+ImHWh3ZQ9G+Da3UC0cO9
+E5u/zQyFTZ6+AqgSMHQdhiuHPFw0lTuRMEwtxa82xlyEAL9SOqKn14P9RVyJlce
RNfo3TE0/JbAVpeNIjGDmWanl8wl07mA12ZgKCzcu36ACbKkiuWVKTObJkfG5zE6
7IDW16uYak5GXBirkiXe8flnwEoqU61h5gWEZetM+zkNo4sGFAukriLCQUF437zQ
oWdtdJwT5pm5FiuBZ6RWTayTS8y3wGItP+Zge6M3Ff6R2nJmMshjy8TG8jKTpteH
oWJDcEynpIoDlMPZ9sR4tQpO9wIfL/9qQZuycy/Pn9iKwJ1nctMpBoQMQfMHcrIN
hfBSOpHwpiYxhMnCUISv2kMcYX45rcNNKBuvNCJf05ba/FnpOhzTZh4m77sS/VVb
fObIhFeg7DHjfp/RbxUsILJjaVgAleZrHvi/QNTsWrkfi2mSeDUBku4iu1X7r+0s
bHMdAEN6AfCSsm/M6e1Rd5Jxdf9EjqJOLdofqyq9G9Ijjqlu4+ajmhSxpToLjWdQ
frBeBkuD6RW7s2V0XJOXL1Z034XRwuI166Mz7bqLuJHpL3UEPHWI5EWetwn8XAie
6AcSSsOobaZhSZHaEK3YcvpbaMwHPapNttzp+izl3XqQ88azns3KUPKpNu7PnmIa
ZsaGguvzrQHESwE75r6/k5p9nMJCS4nh4pI7KsisAMzPYCyMz9JG6mrVoasz04fM
kG4D5vUxhE0t4eawcRdR919vhH3CMVC+n4SpQhmws6MCNZWKT/ltyQ3bvSJ2Wq3a
APiEHOOyz7KI3ycKv0Yi84lKr2wHS7lWhEwnVkz70RH7r7YgFRz7M4vE0kPybeQh
KPmQJqH57rP+vb03Zu+4TSRyflCVci1kYMOeQVamBqlaHDcV9gMc4cpfZsnvwOCf
9HAhBgVXp9/jT19lkxgR3BoZFSs1Jt+4avTeVjr4W9L+wTg6NITnUkrRqS/2sx0C
pBXpK5t7ip7FvChi5B5okb7hrHKIcWEiHMFYX4X2aiZrrWATTgqHhr9/xtO8aKpc
qH7iF3qrovsnX1NAH9swHS2po1alGM2FKCp9FiKorRwovowCPUw4fNXTuQ+TFCFF
H4EFrbzaz1BYPPnvrlFpXJwYs4V/y031r1z96RTKaj6XIuye4qJYTm+KMd13JMl4
PDOmbRr1QhsysLlzKEyCuw==
`protect END_PROTECTED
