`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TX8moyVMYbZukYDizmlkOJpSuWsw4FRua5PMLQlYXY62cyHlpimhdoNNjvxPrG8u
e79QnHLym0fXx5dKTlSYzVYWjJ3B386P7cpZNpb6o8lM2jWip/Sw7PEZwX+yNjwC
/M154oPH26X26Ljg6tr4AX76x6vC5H1uEahLtlrF11Scf4bDBPmtJI56hf5by+BL
lZTvEs250Z0cxN1w2Ha5JZXvb/bQ2/KnskNgG3k9Apmup+KdKpu4E72KGHT249p6
QenFVJpqOvprAOIlPf9T0vt2Ehizqa3szkdxzltQlXtqU3uofIxASmDAzgGxm4cO
yk/Z3uv2MTRp3oniK4SAWkymivOHOi8VqQSnwvIwR0A9sQPULnZHpAq8W7rBFxb9
CrU36eCWd8YTSioxoteDSLWGOjz6Sqb3U2rHoiFnn52PF0ju69tf5ZVNXaKYaxuy
`protect END_PROTECTED
