`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8UAYxGxZTVj6S10xmI71KKbv5a2MkQhRMtlz5nbPbiM/h0C2h3uEcLMG3TlGLIZd
0xJa2Z4biJYLh19m+K242v4TAuXG7a/ubEG10M6QpOi56bjqhJGbeHBxxBhonqPy
UnavE34BIuwuTDJr/OYQ6lTxw86r+lS036p/XvvhY1krGsR4Pfe5R1QfqAyd+gI9
eZwYi0/x3PgZa97cSbczB+nwNg0CoG9YeQk0IT2cRdxw0OzU1UycInuE89reS2le
qdaNl+jhOHgh0yXCXGt79WOieTkKyJgXjv6WQSnysCuYWpjBDK/r5DejvjfA9bXG
jCgRs/iUYrDoUuC4XNMY23oFmNBYH92taFSCA7J0NqRGs6szWV7f0lQFpNC1vz7h
UFWy+Wzl7Xljwx/DQu8jQjL4AZWadbiuBLUa/iXBbRx5HFqj3xiR7kvyFclyI1YN
VaQaZDuSGGSl8MV2PQ1X38mPXvJe+EBKM1KE67snM4/Uj0pdeGDFdCQ4f5T4JqpJ
61JZvbRl8GfZoHq5HAdQkfm4N32T6X/9W7KFXgpuHMvyGKcU5c8ZN47p12vnVp+v
nHfiS32s2VsbbGjEC21G+wyArLwrrw7iAbst9RpKZd/JHxaqSGLELhtVrr+kvICS
u15Mmvl5xuX6Wbbs9zPsuxzSwsvNWrYp+d1sPJgBrarZnB+7BCuFwGxxKDeKHGOc
xNmD9cT+X1rwHECpx1SAZxOdZfXOmMulExxXwhPkcznrwkIPIpvn/tqyp0edcCuu
K+BuueBqsDFyMAyqK6FrGVrTZE592Xm6sDOWMKKQfyTiDVcQlWQPYfyqYIFSI0Qi
vvtNAtCfgAKhEe5/g+jPrIgwcwygLbOUsEguBrh30WXJvMKPVK7WcsmTjWYDahU3
iJjjDmeNPKPKJadkMZk1ajtAf1QH/Kxk3yS2BMydZFSu6UvoDJevBvScnzvxqxnW
vZJN27XlbS+VZuaLuGDU69TqJTxpoYdvtRPWp6Sg8FVGt9A5plLKEQfQ3xMUIRxj
WQaYpyO3i3G+ChnfcG0NUa+0F0n+ULjJsArJSkCHSGs86NzgNU8XM/VOnatT89Dn
p42b0hDhlcoDEG/QdJTKqF+aIurUv7Smzqu+OHWEBjI=
`protect END_PROTECTED
