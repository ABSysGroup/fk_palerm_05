`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
no5zKK4RdoScXYXcU+DizFybGiEFCgZKD1WZYqlo8NZ/KCXdVPymMSYiNl36nNI0
zONw5zBEjazNv1ys2fHv435nf9MuQ6ALvZ18Y+v1CgRmXhNjkzIfvAL4PLMdMqqg
YaUlJ9AOlk8qZvNChVVzUpgaAyt17tDlnEwZqOBHXoN5xM6+d4HpWvBDyK5WT+xk
gasZv1f/YIEUHEvaGgjqMuDTn4WWOwrbwTG9tySrHG0+u9LmKLacxfwpzgPHLYVE
iBIvTkGVi1oHoy7E97+qymeJNgML9wZNMSeQvwPPjBZd08VH3uvgwZXhv05ATi6Q
OeVwMmpht/1ZpMXsOIgIjg==
`protect END_PROTECTED
