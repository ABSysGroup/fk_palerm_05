`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y/0Zv5gP4gDe11U0bWpuupo1+WD9ytBxUCx77kA63BvwKtpPk+yZ2QmB1ntltd/v
uFBDbWC222zJ2F+p1wEc8OLsY0f9ZL4X3BHyrtsdvAIilHmh0j9Z5EVFdm88CQAQ
W+qVp37n7AJPMbUQ567LSJ9xPFe3Njpd9pf1zLHvWml9VcKeX+3E+b1PR8FVqBlX
nt16OVpspGQenIROHVpBUwl26Qb1yLwf9AbkiSaNOWe7arOXLqsWa2s1kDWQgCYW
1kaXzWrHPAPOMuXT3k6U86MQWUJHiT5grXu+sIbC0GsZMOqxJ467+QBvxsQviYoI
r2Z7RWOHXMoQ35vxzJU9em009opFXFqK+ldPVaz8B2I5HijYBsIZDcl2+KXsT9C4
SWbbZO18fMrtf0+Ur6qlnjSz6SkYfaKRA9ghc+XZ+yNNE4RrQITRIByunjHOi9cR
twUiqweLUvdLAesgyonWgA==
`protect END_PROTECTED
