`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g9XGLw445QiYL5INUQ7qL/D4JEWZEO3bCiMta0/2zyncMvU0zC2NvWfF7k7KSP7X
ENHarpXYMmiaBOcblg9OKKHbVa3DnhRGXvjNa4VFszymKrlaonj/ASz1o+1D1m/C
OFvZXbV3ff4M5zncTrP6PlPUIAOHC5+FsN1fx+B3sJZ75VrMof0rHhV3GvAXyITB
kYvnbJYXVf4TD6XNfFYRCw0iPgCKNdyDCNf9I6fK4IRgjNMif9oeogTTNSXUy4z3
AZtwj9QfENP8bugpox/zx3Twe6DJgMOIuyaa5YvxDp3coU4ojJyP+LeT9mZjNS6p
8CigbZ7b1rr7KPBHGR0oDwqSzPnOVapC397EGlCfhJ9RHkHh8f2MSYA15DdaHKQ+
kSDVxD+SV3wKXQ1kBZ0n1fm2PmtG9tfuY7XkmvlI9XN+llwbTJ6q6tQI05JSZEdM
fly0YrIl57ne9SSdm7YCI7FfSpkPA4smS7xk9ytHr6FyUPdjvhA4HKwQpAT/DvPN
f5PvFcqGwH9kPe2jKRds721ns/bwsdOMLAov5TT64JPnhmFyIX1b3jLeaKScY1o0
zP9wKkn9EcNNbpSQeNYz5iZKGNq8PhUR89pAgiOfdQWMsKW3gyPwT5NFwb/Bm9TF
aNFWL9csclNcF/RIenVuqlyxiqm9wn3daEQeKJNVW/kLRWRWr4CISxf1xx0ezygd
BPsLO8+kAXmKv67aQyoWfsmhA18hvRXSPM3Yt9+7VciuXPOq1hxfbwNzLFWcLBoA
9dF4xwb7Po1u6RezcDRXAVUHUlD5sHHpdJTmxjRHpy/wwut7CfV5WoOnsfzsmP84
+s+Y0Sv/IoX35rKgtUWa9ujyLJUdPD/ClDbOXXg2Q8e7JWnzUf8jkbzVdT16BkS0
SPCwQ1l4EW0nuKIsdFpinbGyQ9jscei09ld0wN61jPUEG/RMNsrU0A6SbV+ciHpC
1DAJpmp1iINZq2IOXLWIf12XgOOuEjCHtM08Jb0mmMHNHGDHrsEaLzgsdYlmAUwA
Pa+EOb0WfrRNe6JdELNpY5iRq5Nt093MKm8phUgCmtV0D3sSrbL8ilhVxl3HnuV/
I37CEgT/aFo48JOLQN0VbsGYdHm30L3HEpGTr/3DBi6fzRJUXhvCDzJl02iaSzFn
vNckRb13KyV+1ZAX74KDkc00aKLcrn6yJYPoQnkYkLNysRxkMRf0AQCxc+bdY5op
4zHqtkwM5kynmLzMoqz3t0hiz2tVC5GIcTplYbfXiffQmBAC1TN2E1BVtZF3L8F+
+PIVwZHFlriDyy4htGr/GJa7Smnog/mOERhSKmhFbwRkQ97GATrB7YCZb5XUqVEO
rZFZdpCxynKcODlOsTPbNI6ed+kFiAhkIaR6EKXXQTLhvdlMjTKAyVaq6n6eSl8d
sVizuX6moc83oy0v1X+2p+Td/VqSCa+dMR4T08M0VOVkDmKA4zcyc8bjiYokOBqs
Wo+nXUeeTNSgWnToBF9lzHYvt56baUfmJkDkMqs1e6qMHSlLciWgilMbYMP3EweV
aZYTfc4BfeeqSOuSvr9eCxMFEq0ZE/nxh6rMTlbvW7+O50KAzOWql5jFsfs106JB
D8JvnJZCILOZsHkcUCWAJoSKkNpMbrhW57mYexnNuYHOHXpXXR/sUpopnfZchGjN
HSKJq/yO0JPaVvs7shU3KKAHnKkU6FlHr+6g7ADIupfqdyWm8B1q3cbnKZZJtHNp
NaJ1oHXJlqxjy9A7XvC0JyiPY+lLGWwrZVsLcG8eUoda+yF+LpMHyZHWPN4wVKea
dgS3kUbwINhSazBa0Y9rnBNgShquwXKZKZxOJKJOy8x0pcC2N7oRBJTFRKyoUeLN
yuFzuT8hUGyRlm87YrXZSEM+puAtb6GDZwZqGqYfXxrAZDORi35EXZTEDpJ66Gwe
zk2M7+h+eRLlR8duWHF7JjSKNMyq7xiKrNesQR4CyfPudRIzr0sQj5PJnmU2D3Wg
D1W7gjJ4qHuT2ecUesTaXvfYsgxEydJsjJedHc3o1M9hS2falk7Faa815ZcuoudF
qSVwOwhvH3ULdQjnKCyVpbaskhRd6MG4cn8GKbuJOAWpNw5kfqkYklsrJgyAPEeV
9Yrz8b2+ZsofylbA/nl5dP8VBTTQigAofg4UhD+2AZy/nsZm0z263ewdHRpx+6n5
DYJR40pQClYMoZb9WbWfk3SPWJJ2ojJmhp9M4yUp9z4gcMFxeBCSw6X56o/4x6Tb
UybwGVD3qAQ4giBoht4omZf2hw5usBn1w1KovUzmaZkfChryBydnHWgNnD6Lk5HI
jJZ0ko/8eFOs7GBfpeTcMiojdpT/3Ix7wT1b3Zvt3+X5NYUQ6ds3FeN9QoVW1iZ3
QYne3B9q5ySqxqAmCPvgG6wtFbKISlYmHcLL63yV8urd7556SDL5FF31dX6N7S9F
LcV4KsBalt7HxkXpU9XOmMRJRV2OH7N2NXx4elu1U3T9Fo8TJgkSlCq71vWv0DXD
OnXfZ23pRKR2FOV0ruUerFCbQDrfU/d5TG++7dRv7oq437x8dYY6qnez2r5Vs4k+
3/h+q48cjGEWlHHk5IWw2i2/f/+AfO81b6CXD2Rkcjz6231X0S4EMDCieo3iqhE5
rtwAobS/wEwuJ5jyaKeBuSdHGajzEAtq6xXmgiHRanDKKwo5HGQXJJ0pGhTsXTT8
zaFT54saPv252E96Vs60KoNo9aO4VQHNCq4LeLjEaLNmVKSUXvDGfDIzOqn6hBKB
7sMTtwINOLfx6e4F4nwD1kcX/1Hc/XDivkGqRRMWPFZub5BLkVp6mINJgMvKSXxG
jwI1UAmP3jKUPj+rCVWdj669hLbSfxcvAWzJF2UPUKffMcewprRyR8EYLHDOwTwv
Sg7Tq/btgfWKXeATtxLEuBNaZ1xXXAt6frzNXJOkpGMFDVhL6ZSvrALSGEFFktAL
x8qOnQ3wQbJENqJ5aMMVjEpaZ4T82flnHqCtwHKN3s97Q1OJHaJa61FrNlC7YjtM
4uVZ8w4dEgRWhp7gQMLXjkQXWPdVXqT0QNLaHNwdHdR5mkEHra0rZubXww4phJXg
lCrhK38wxfwEzv3FRJgHp5TylL+S3VQKVGqdmOzKezO/bGFUr8cxylCZHTDttJCy
8c5tn4oNex8eAiWbvm5/1MwpSvlUy9Ww/Hi6AHk5Gc86h/qfzCTn5FMCly0CEcIX
HG7TQ1jG+HPSPaxp9kGAgI+sxh9+AU/ak9n9kTZFgb0y5hOG+XjEkzNvmyeFsWyN
OjUS9Z+YLMwAfj8HXW9O8yH4wNNlkjDF2N3nH9KqsW7xeSc53KbqW2+G96HJo+/3
tvoBm84LHp2VezvAszufTEMLsjQrKQ0EuvJ5t8NXPbdZpv7ZQpd/q3BDrM8bupou
ziC28eCeTSSgggJ7B3ePYIDDWzGJdRDb6yFwtklrV3Bjs0SBGOTqhL+6d5T79yDe
MTNb/tcbr8reRdnBYOX9dkWVyTFjZdbmYMM8bsRaKULC1Tx9Qy2AZrY+bvFUzmb4
nk6XUsTxFpGY9nVA1dsED1XEE5VMrXdEIKCOVBjxXfnCpgQQGCPyJ5qTdYAgZJPv
EZZA0lTlFDr5RR+tBz7tivGKewcx/pftNgLMB7GoEAP7Sh7GJqN1u5zg4yz6L/d4
/pSqvL7O31snYhpu1yVmxa/BwT3wabAuX5cDHQK/NgPpnxgW2vN9JEHDwQaDhpcr
hTv/J7xFknSJKt/L44TUIUH4pTJq1CQ/Za/Dfip+u26TCtUDBRYMNN/vvuxdtSiz
X7bZuAMCeQJ+AAmKQ8u7NNsGbU5fDVYHBhx98cfe1dCXTyttdhxp3b91y4rFv0oC
lXwPicv2lCzJOpib9NVRepyjLmWbD5pj8D0QuOzjsDX+WPjGHmMMPc31bwvXIy42
vc0TBTOFwUlMgjaHt5H23OGGB27RSWe2qmQ/2V0UnhbyRropx/bqexrhf59tcbYa
mh09U+HlHMuGxSBKO/MJpLy/ItzWZk0z2xC6rLvU05xH67Y19z9c2E5MqFiyh57k
c2UsDszHIuwYKkByOAQVyEHGS53lyU6bQbSSQpZcsFkbfOVLcizmz+l6qLfB6Nkg
Kv5I+MZCvL33y4OirLB2dniPCI2GDiwuuahCmsb936U+9S6+RUubJ0xShmNEopjG
izUJp2vSxEPm/U3mzYMm1nNzjdXNXfaLilzy5jSryboJdCIm4jFEDdmXVz/2DkCi
Od2ihX0u/D5xtHSM3bJI6GOVoH+eZb8T1I8uxcQWjUU+C9/rICR4l01NdcL4SUFF
oZQJYul6WAgPy6hNvA91IaKz6QR2is0xSrcUPLOHILXzSF86VR7amxVTbxH0KsaP
QnS6OMTp0KVd8e1TB3+ARjroB4OPevBqSYTIMO9XhaEe8pKhumlCWyDJzaagcaim
WrwllV3K7ufO11tqGFQ2JPn3PdzlQvkng5Ro+x7RdL0JIuERf04cwExKtsVkP+2o
aFV3I9eVvxA+uwpJqWNUS8j7SqaGmGhuqJrNnePSetq48tLXETJAGFvCSpiQt8SE
ycvVJM0JpmiFEvhi5skhLWBZODfqoYxOvx7xK4Px7JYoxg7cIOIzJrNZAH6ASI5Q
tWxuvro8+ny0RN0haCmJedgYDAaBX3YTR87NS/amwsrkewdT2lO1/xco/hJ1Xx8+
0FZvFL8OHOFOAyYSsZp/Uyj7zSZoNO8rAlHESUlq4aFl1heT10Hr8oBSim/EGzQu
Jxu3+zJjetNmHbK1qEt9hyKlz7fnppdpaG68XX+8wLepwJ/M+YjSUayzpuaybd+P
eIO25BJGMGmm+7tV81qXxv89nYRtb1D8Lh0NU7ZLS8ZvkuhD0dL8o/XHH6hZGVrY
zeeI1r9xvtZ9sIG5mnBed67rGXsKdLx7KstYVZs7is6eZXa7SRT4RfB1CTAt89yf
tyKB3C5mBIpGNSHJSB3joPj+ck1PpKYll5tv1V+Mo0D0OAy4ayEgZCy2nvg1ht0y
/plc4AHt6tfqfBduHJRwnQJHch/8rWP2hir1vyWln0C5S/ek/ml5puu9ni+nDQ/v
TGy36yAVl3jaBhw82heY5mM3j/wfUP2UFQlPZFJOfgbwayUvD+GVgpMz7xLwepds
Vf+dWTYc9bbekyfc4XRakg1cFIhcgEY7TjwYlKXLhET/tZJ6KkIRN2Ws2vPn31dP
dwr5d81tNKpgtT0suzw4kiW2gHXVE1K6DhczFwDfsGJEVzygx9DzzzA3ghGBWJV9
N1oQezsvwXltugfcuwPyez9bvQtsxLYK27WWHogMUcvy0krwyKgbXZmap+usXVOH
`protect END_PROTECTED
