`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
euzvT9n1Z6cZLT8eT3RyR2GEmqE7/rp8tZSdM1OoklkAQ0E28//+gXuF3/+0KmHS
Ma+xbop9AJQquxOPOABJkVT+W1npMHTZ0xeyxG8fp36blARz5grVOYv0Xg9D6rRr
3+daai3YftIQhEQb94O3oBPN9fE0n590yMRfUCJSrKeGamCSirbdZqvIOBgJrMgd
JRy18ECeiooLcB9phAcfYt4d9LW5U5dBxFM81rXHbKrIHFqe7AwgRgPVYRDH/cNy
EW4jdf57jUHDA8mIh3whAJBc6C7l+hKjZfW93J1IPlssqHe1KA3gtvJnTccJemfO
RfBFx9kj9u9qlqbNYQERt9bEo9pGrlyCwcX+qqzbX3sKwXjzUghi1fiQM0yhOP94
eQCSBEOkJkZu0kp9QEkjXnhBM815zIdDFU/BQVRhhIUdYhwPktRjmI6ZX5jMS20Q
pbG1Nkx/ZFj459FV4IBsKsSADEJL9RGOaSTJMqo2u8el3yKJuY8IywPiVFWtVzlw
Tgi0k4WcErZAY3qGOWKPA/I1ZmuvJRe3b5YHruT5EGf5Bm3BdhAdGOh54hczOE3y
S3H1PXrz5h0sWDnffZwuSOCGSaurIqlTtBbOKLttWqpTw7pB8BhsaaZs9slFIi8r
gIp/5HrpgI7CXhd1KBuOVY9lXxRBjWUWIJYigIl08355EWCG93gIJMWGdkVsn5Kx
iEjtHgeSd6ala2zw2J3Wteqgh7+IQrdGBGVneXEea9LOfA/g5EUcfitQ8haYicSL
QJLiscDNDfDBK6PQUxF5XzFWWfMSsS9fZ2ZMFUQBNaiDXk8+tez4SrLgJP4f17hM
A/cG32aJSG4lMOPayQ+PGM6WVWYwe9ZqZEL/vnSptMLUbJj0GsjtjGBR5xKQ1KiB
i4cAFpcuO0SDpi8Iqf1ewAJiYIq+SFj6cqiGp6GKHwCTfZtQJmn/Z3dDgFQQWGMg
n2fLCPODo6x0ENPBWe+JUWgN69xix0mvoS/gwYj9E76YNKQmsnFl5STIrD6dRNvZ
OpC4EVamVwggg/wrULIq/QsJgRuUp54qlit3ceHpyMRR+4foF35v9moOqQQc44Cp
63PHY0EwVMrzWrNRIGKUUViMO2uwb1vAovR9vWH6sbsJYq0LJpVujrOMc6o7MgRS
9hygJ+YCy0segVHeBri3owWJg9I2P4dm/yOJFXcmLNZzgThDr+AvHPALop86w9UV
kJV2HAXjCVpBD6zQ6FfyrqF+5BmAhsV1binFodgbwXeFCZvqpo1R28oH39zNAUfl
e9+Xg3JvXoY0AKZij1hoHBBmJNnCekuWsjcpQyZ9siOeb9wUsChc1H82SNCDyorx
UCoGqyQ8+2Nib+Um5INyB9jtPtLTmKb8A/yMdbBkbOLFjt0+3P1rk1Rv4v8RCrMY
G3RctiVtDkvR5On14dXt83A1tGjoUGrd1nJo7vBT0qN0kV3IzG7LfWLmBKBrIhW2
iVxsGYLjiISIspFi+9WrgjdJ9RSVMYuOG15Zt4/aBlN9lP+3rV2YR2qCdekFhPAg
PF4nW2cjQlu9Ru7uPmXvFtGX7eqUoCg8jmBA4P23MkVCjy50rSfKhAbwn3AmRKEV
QUpSrQBhp0xruLfril2g3rHinwXe0OkBDs6bUn0G2tzW+fWM9TTY3ByzzyeVAYlN
qSfb+RvoZUU5E6yp1T6BSWiLBGZnEXvaVnivHIawL45Z2pWsAARSjayur4K/Bifb
24t3ZhjaW3oDZqnrz54OftRgvlqTf1zPkBFPSJL5vHaLOhyAqgv+cy7IUi5FnqLg
UFIMt0ZGcpSkUmhv2y16C0MVV+3PRvmZrgPTb0MPSgEDwLufZ9FU9DJ47cTlxX9J
G3eCAWh/NyVvypbnZ6yAzNXaHjnt5eoXHyr6BZ6b8Dxo0i0mrpVfE7rX9nonSkoz
oZ6V/DHep4vp1EK3tYq/G0uqq/Svf+/Cf75U4KOfvrUIv4y1+sC/MlhUVc0Yl/w3
B+aJq8QD1ZZ86BaBFCtyDuccck4KeKZ0l0+gGll+jIAE23FyuISnxj2Mp6O2I8Pz
JnK7Meh7YKfOfR4VOQI34emtQ9vWzoa40BRaJWpqQJyqCQK8XsPP7+e9jfSHFLMB
v7FKCYylDq/yb5d7zKERoRx8JlRi6OOFJpsdEDQUsEDO5/dI5F0CTKCManWAqYT5
/l30g9B29LXxZbv/QWpwUVpJQ2mvGos5pa7w7+mAZmRp/gZ+3m6s+vds1/YbFAYl
8IXduR0YxTMmmzqC5n9CZdywhfIVxMUh8S1P4nub+Rlp1abqB9E3CY90FxANpgow
4BbdKTxwNMAsNoguj4j7j2lYDH1tWFqjdD72fiasP9XOrOJo6IA3yZg/FBFsioQs
9n71FPOJLxeDH+Me2roiINwPf/bfd0RtgM6t/OwQ7EAOu1gSfk0jGGvoAQsvbxHN
YXSzLn56JsQbL5rmQ7P/OeUxAmbXTD0QGVNtfdjfsE7qTbvntgB42ynE5sgCNkDC
eVpupEysMJ5PQJP6cROkjR8cxkMVagOOpcC+YZ9FYQO/1EKpqzGA6LNQnUyTha8z
zYKTmxvT3pUKbQ5sEZRUUoitsVepJPQGMDi7DtTFqXm/HIw2dep9gqHjmabbtXFT
HLH9DQ+Vfldj81yyLks+qWI9kRvh57lmGvQ8fLG2p4eM6p6Kp5kNqtSriDTJ6Xp1
nuIj5xK8ya9aWjaXJUDvzIjOdpFJzeXPzEHGBuTNF3wmn4KPEWyay02lIt++zL82
tDlPG8GGD68DuwOXtwNXv+bp5tVPwpdrooma71F3suVyvkD6oXYrZNbULJv7qaLJ
dgBK0QjyGj89JqESSdUgVXPnxptCHDk7YUYm1KFyd6diBZC/6CwZCtgHxJtDMkdK
YF72ZYM+Fpa2ygk2iVcuo0dLng6x0RZmtb74QYsG5QkDz0P0pVQn40mUqcPXtDBm
iGGcJMoNM5TLv1oY4KuDmoNbWSJCDPHx4P5L7N5xnocONBiPg7BHYaBJZIyJ1gOd
u5jNIB93dZYptqxAf3MdZa8tY2RIOzhnblC5O/dxOoPlTOGV1wdbNDNN23LO8qdq
e/8i0Elg4k2XsRtx+pGfVgewXSbFj8/HsdcbVLTofL9sIvmw2NyRPy+RoTltKBkn
EFDyvO96g38AOxS+0giyYJ+H60y/j/yK1U3eG0SwElHJopLz8AgTvNhW1FwjuhlC
HvHgBTgUiNHjrlzLhCfQEQcxfskHXvF6wMXW7w17PT2ZEoZIjMYbo+P3w+KpwmC7
GD557BvkLP21msJT84GuRxPeS52ukqJ2EsAG8tIYORWBA8pY5e8b1ZdmJiHOC8b3
NASs0+JEsUKfub4aCQCKo6Wp9EdqRGhG2gqVpi0fQKM9BHCXIHtYlMAPL614EUfR
F0tP8oT8eWD6Vu37sdkLRC88/q7Jrym1o9L84ApK2ICGItWa2hGQQzFkEP+CJt4P
QBcioEC+k5b5A6NGaiST8X2YyHl+tJo+pgG2+wwYbC92LJXGdYSZhRGGXlNYHrJu
J2a5QiilDQ5W8FQeJNBMhEfPKBz712RFDHNr65V9S+Dr9q1GYI5b46/EwZI2s4Nt
8zf09mp/UDKtKuDm/7DWALW+4/AsLsI9/rH1QCCbOkuoruhOx6VNI6gbSRxwmBiT
xcyNxppuNmOsFWdeJfszJxC/BNhP7b1+/jKIwV7EZmQwjLb8ygA04TPDJJbxNytk
9RDQmCDOUVeEyH01QJejXLWdmeXV9bC4lj03y9E3KdqdwdV+So4SWCXzkwpqTvMx
EseLKWjLKBTnnXy9Qj+XSgsUfeT3xADfRfY282UTmZEoihH+YGOOzlkFceYNzjiU
jlB4NRJMJE5HtE83TO8ICkzdSwVDZ2BbEkCNK3RD3GWST6yoxBGMMQ2heR2DwAM2
zcbjV73DpcoUAXcTu5n415iV9EcPKhfG/t+vHcvAwB4vb91zvfyuetfJJs/44qD5
zy0Dz7F102qXg9O5ZRP6ELgfTDZcFSwYWv/c9dIBCT+isH1vE5YWuKhIW1IG4hpO
mhfOq418qpG70JAzg+wgubZiO0hX7ghOikRVMruCCgJ6PwyLkMh5AifffPONpF7j
c7eXgPvC9huagMF5b4qrMOsDE9LbdpAoa61/djoupp4veR7giQVNSs1jirVffttm
ASsHrbBcWoqErW2xqvBKgMbvjXHMp1cYVFKuqGds/VeB8vRW0DJrG3fZzYoFtpJx
IXs1w9IY512vFjheQWXYBfCOltk8/Tn2CXViAon83r2C+lv3sVKUL7WyITXRi6td
TVUAEL8Z4YVb8mFwwW7DgV1HKAzZxrUtr+70Z5HXPw5ThyRBOzDzbq+BlEQkj5jw
qmHfgLYkFCfkiFVS73TomkUORE/rf9RWZTxdwXJ/uTERVER+LQVeJZJqMFf1vJZD
bMsGvuf5A0c0D0BsriRDHg5AYSQamSZiIRnwuqOG1+f6uCvJGIi+cSYH/aj0zU26
jl2GuDYHTqHOQ1rBNWZS7p3sQX/xr2HRuvnLA7zfRkLV3pBgpyZnNPOa2FSdieNp
d2iNZW7Pxx2xZc8IXonJE8duRWMIWZTVAY20ShHqLApEM81Oaq9WVusOn23YHGjE
JduKbXgS6jjucBTc9YltgizcpbDEJeZss0yaGHl+dAW5uzfuqCUh9VtPxlQeJTk9
8232nifMiZLnHSdOzd7UKclPr5WZIM2Fm113kqs2jVPqIJ1sjtj6dNEwi6F2Ngk2
d0DeH9VOnt58SuPAf4EoGhnPTlcUIQYOliIxVt6b10VTTX30HhHOSQCfL6HlEVp1
um7+VSfOeBFjaQcsSMG9zD8Lsxu67tLfe28EmuHtCe6d57MG/eTC5ZRpiRWcR/PR
LEovfV6+ywSTvOIH6hRz2dCUEV3A4Cyvgm7aykUxeqOLGUmgHkmzqE8gYihHSShi
Lo6Gf54sBu3WUTg4NGvPeUUo5YOJ7DnKWna5X8Bc/fQDnU+TuqwWMkUyXbhFhl0H
Pmne4nwAg88iWb0hrKM/UyH1iXKVvuPfze7yR3PQaKIdVTd4HXXxYbpJMAR6XPzv
twaGmKOZxaRVO35hM0gfMtUsnPisg+p+9+gaCz6K1L0DbfepjfTolZ6HrNCd96wV
/jRDAjThQRJEW9HcjyeB7vcWAu4a09nlh1ZsnVi3PsN9vK2vh/MrljPypO28/z2H
D6GL8Tws7B/08nIulkRGdwvkVtbpRW/YOWiBx9t7lEoi3Sj/gG1ZRzYzNifvH0bK
gHSJfn8ZMbdTd6orIEj3qgpeS1WYOVkQIxqeNKXsKuSGFqeBI/GWpHYwxW4qqOAK
mGfmfSNpjrFVke7BWigfYxTn9tK3rZlpvxmhIOVH1mS72+44EszhHsTzSqoipcAk
AiEEjDjN7sAAxiohO49JlxbTc8yXvlTPhPo6Y4SUQ3qUMCPiNa1MdZUC9q8jbCPc
+Vr/Hms8TAGrR6oh/giqnKsGPURG4wopdjehZhVm7w/xc1NAS34ILS0Fhk3r2/gU
giA+bmhEVwBw26WSegCeR9iuhRsxlY9h9zLBsSfNtDd8EnLV7eVqNzUHA8W1sevh
f5Y4oQ7Qhp/uV6UCY72pCTdPOyblmafnsxNBPKT7t6fEvqOTMj0JYYMn98PDqOIO
nfkmQLieaYHmbXPDAcZ0l9fo6nNRtDvhXT48Wx+yS89fZ8/9eYVXMokdrjHpgEFj
nZzef9+St6A3aKRcn6RVlA4DD2jQtjAqU63GGdgztRBTxtyWfiuMjdmStTnin+N7
yH6C7duJ0YYYhHcmSTafOyLpWVChURdl0dIy8cU69mNSasxo9vixzNf0HgpFXbwJ
gEfx5BSPrR3EYprbsd4RbMZ3i4cSK5Wtk/1xSlUkxATUIptOBvC3xM4BLtFSxohW
8bJ1FydP+G+ufHdpvnVWUOWQ7bjNtP9PwCDZtfOY4HNDRRQ1PC9U0lWnVhZnQY9X
ScyDa+24jvYG2iPfcRX9BDaaesMHBTJeWwwmmpbPx1A=
`protect END_PROTECTED
