`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PPsiu4wNIaVMYGOY5Oqx7vl8aVF/1xbqCs5juWyEaFYGF5w6ZtE0j7AW5Wz8Htlt
2rdMJHEKMws3dGgOkVnZKAa6DBju9DR73tHosvIJwr8AaEd9c24uuCurC4FToAdD
EDzneCy5CM1LPIh8IWhV9HJUCj3OmmDE8JUQ+lbmrtx5CCfvCrTptFug1/aAfOww
RZrr85Sj4INLiU16CjWqKnUBmCMWYNnv5AATzlLwonUhgAHSaVMjIK0D3HxVJDZ+
M8X5HbER/6MHjY24X9RH+D9gwGtnRnL3E34Wjw5dTr6WYk9OBTjZHSnaXHqIO50w
czO5w4QQSlLN2Xfwr/2OQm1B7vfRf4Ed/4PyawojK35mRi1Z/3Q0Bc9uOTmVGNXV
je8IC4k0xR3zsfRByJXuiZQ9A2Wux8KXpFUHD4kgxHG7iYF5KGAPEHQXYCNCGK5E
JXlU/kI8T7IU9vykpHFzEBjpTKUxa47XDNq49/A9eUFtoXEdTsmmfAUfw3/RblCa
2XZX8NgJXiZ2SrpB8cgZw6uBB8hW1w19119VdQPOzMmzOYSrf9Ph0+fRxe3czAty
DGJeV6Z+Sn2aL0wh0l50GCqLFIuvdNHkAstr1Oiw/+4=
`protect END_PROTECTED
