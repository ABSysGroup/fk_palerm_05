`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JZ1/jETW7sCuSVeRvokAh6A0R0WMs67TaLtIBQHHVkRM3aGY+mg109Rjpfcq9b3H
QEr9Fdc8T5wNDoMuocv5o5uaY1m/Hut28+OjoSxO/Q/tSUWkn8hLVfiIMujqyUmh
gy42BlsdRjguJM5WCaDNljWmlrYq2/fZpRiArHOR9kXZVNxS0o7AV+nQcNVkBWS+
d7LVFcNrJBW9ye/9uMU5kG6hckGpJ5ls+6oOlEoFuVb2BHmLnM91LVhqx0P0R+tr
m7eBvfLcksAwlv/uU8DgYdKqeXF55glxV7SRdAAbpSU=
`protect END_PROTECTED
