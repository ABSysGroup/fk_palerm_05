`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zq/FDO4XQDZjmJJgY3aWY2XNterv8J8QI/D8JL6Xnh0URG4EGKnyMeOhWp2jBcZB
wVPJsh1M+6Fyx24SIdfpxZivFolyubvZIsLXNABV6rHDsKuUY+v4nFAQrmoHQEwK
P6vpZc/xaB4IQdn0Uu5pp2PqaKNGGYBAOr0nqQ1VLnLOTBXsjQQi9ogmksWoo4Vg
TGubjZ+sjoSW8b4WD9NdrWAoqj0/a8NQeX/xtB7wZfRWZAoN7TP+NaQtB6qlduXh
PhDiyCMnkHmUJg84UwLqgCl4YwLqevByFSs9e2+lNl/bUVVGEoPk8SUhdjB4rkiJ
1BPSGcNSxRPObWVQy2Ob9GXpuYvc7AqvOdYbm4Bey1oQi7j5oL3Pg8PtQiwZbPJT
mudqw/93B7UugMuc+Ac+md97lxM0oBTH8Pu51sZeSUfHG+Dva9D6wPMvwsDVZYIs
x8fsP3awxGTFG+GDhtL5Elth6XihqViLBka25z/MOfW2id+bHcJkQ6qucFZhgvP5
fZkx10ex1gcXP/mRayVF7zWIfAJYqvCt9YFCFoAddxvuCaIVU6Ccj2gtnS8tyW39
3G6q4nFsyP5/7LiJjqz1nYoPFYH3rt2RgHJeELfdAlCsVIHYEkXYXkFMMEoSAWrO
rkN6JpUzVQl99AB+A1RJ3OsuDwol9BVp3E1xKrkFyDOcOo+BoK+Rw2ad229yleE6
KVUMZpIWqtBz6QOsUuJwzV+znbgEieB13XErsbbUnyUbk50SpswDoJCwoHcO+LGe
I7Os9dnfSL0n6RYslmll+ONI2qLZPqJjKqRoaEQ2/yGRPEzyYu80x8xNnOTGYaq4
KlDhN3I3AGoppt6QXieqNi18cxj7N8DqJc099nibEravNbCMUDlMjJhPesAa3Coh
LegfmH6zH7zSKeCfKIE5T+XadFuB0eHCXq49852NBYgUPb4qrv8+R1Y6xLE6SVJy
4zbzQYanbid4+RdqaaC/pZBGWOQAQ+AQGQMpskZP1KtpMgUvwuB3jDXy2VWs8/9v
r50LfALhHlJIEVysdoknfix7hU80Iut79KH6AgQW0bG5tSdip3QCzl5Jo+NJLgzY
DAEMZYYx1NFci531RR2xoXZmixEMNN2VHNjtQnlipS6p907FBXvrEpfwUKBDc+sI
jdIve/ni4Xh/3wlBhiw0hXd26bbBnO9hNktqdI/Pqpluj/lExui5Vzs6kq4sjuob
yhOKZIK0RQvugLKfQhGXA+7O1TIHIkf/F/+cusqC5wvKYSOxkwLcTqGV4jWEdcqs
IIEZHuakYkvQyQFAulzcu7x4OqA/V0HZqzgp2tBOnJCQnOPcrrGJoRmqXeWWfOQd
TLVN5oU+ySNKvDshABOCjsQfeichfV2LTH3g/yAqQk4aVKxgN8aVLd1DYHWXx8Sm
lHKlaa1pfHOfI0NZoZ4+101bkEf+9vvqYUCPO4FMgotprsqZp7+8EwcQ1zliZCEy
kF/rl6tAX63bxlFO0XeAxDOhs+Y1wdNXLke/eJeBwWc2vxZ5X3JnB08rj0uVHdcn
i5vlawrNQOdQ8J7FvtAVvpk5KtR2MD13txgTGdfkr/rM/cs9qZRgFh9sY2c080Pc
n1klnC/+YCFnG684FpPXn57pGswjhWJF6Q51mpmfmsFxCBJy7CX0xnTYfH6H1v10
wiMA79O+293Iai1NP14nPmUbcnkyJHqj/F5E50/c+IQPr/nkqW1AQTHrYuMar3AB
fFaUNr14sE31GcQ518JOnYIn+f1Mxo93IenKgm/vQqzNLXIbI/lu3frb0w45dlgQ
z7nhN6RE/mFDJWdg8254mtR8PlecYbDGmRiGegJG9CuhGVdToLnAnYAVZ09FQTML
i1f4Dd0C7LClgjoQx7etsidAYeoUtQBTkCHxua1Vn+ZoQLIjOaatOVRWUD6kk0xj
PXp7AfDQSaKzH46iUBj6rYtQMU/iDNsIyjBm+b9MXBWl3Y2TPmZG41mIBuweLHeM
jKVE6UeDY+7nGXqhlUts0sWS9VQ5wLX429T8Tsc2Pm8g+IDOZ96FFBld8LXHP5pf
PCyrxyeW24pFTg6LihJXptw1dFDK7lVd5A3fjf5U00/TSAqQ+aW2TY4SC67rYsVF
8VATB7qrV1vFGoenqU0tWiCw0Z/Cmye1ei6Wyrdmwr6a/3X4gMUyQKhVAie6vK8F
3wJgquS3kjm5L8kFZ4/l7e6stO0R+7RLqw+3/EzQcUf5rHh+AOjT/EVt+aEX5OdF
7KfDPvgcxiO8LO2WM5sQZDcZkZhsgbdshPjGSn4LgqhiiTOpGru5zq5Cfp2AHsRV
PVrF8/zXqC11ppHcgJaVBJ9s6UZPb8v9KVlHd3xib1KLFqHRQv9ID9+bPzAVtF3C
vOrLxSky/QqhYlOSozUo38Kmh+WRm9Ae6yNOLyAO8WyUGcrZKI1E3kTwPv9yxpnu
5YOiavTYbWU+e6ia1MR9wbOhYduU9td27nfkPzZVk01FDCu6jnHZnIR8PetnZCp4
u1c4/dhglvJMTA/VeW7ESgOIyXk/kxYWp2rHoc6g7V3sTRKEX/op1u378fSfs2Z4
syZy7H3P/icCJ8iB61iE6apw27yoraOj5p+n+W+doQYDu/jUx+Y2BTsPIcqXVrpW
HJvmkxN983IehAi4ztBSiin49dwwgQHyF58lHCs+Psz7ldeYBipq7rZSo5TMGeNs
PPB4bJyYezpgQ01kBFPJjKCmLGxacjgGtJPF7O7lHP525rxVrLq6ktvDa1dWvH3J
sv5sZgVOAfFfTfETp1lMGz85b8+BSdxQKG8C51v0b5K85v4u5+ScCuXgrphG9fZb
geRSHM1K4P6aD8SQcRP9J/Mb7V8BLP4HTAn2DNtgaAGlD0Js/dJ4nRjIGNY2/LsC
f30lHQbdIDCwseCQaXOcyKYle9xRKpdDi1YVPwWe3b12SRJ1xibDCd+11i7+0KEG
0sSnF1n0FhIXtZHOjrNHunYlxVs2oX7Is9URpYBqdOwzpSFbO5KXsGD6LKlVx35p
FDbm4WvcnrtZ4imVtE4kjLfT2pdcGdpbu/rZEvb0VrUelTp+py8sxuoBWnKuM31k
oWw56RStsRTwkiVOBnEqJphZrK+SQqulU/7jRTShWIU73ilN0Jaw9t6jzCJ59uOh
EkIH3+CSvhTRZmnbhtvflcYKmF00fIi64Mk2hVl5Cjhk2JJgjmGc5OQV3K2OmB6K
6p/lcoFp+IAczKiAzl6cTE+LRyOQ1kiZqswbFGBxHtXwd8SXr/NjJMSGorTdu9KI
L+It+7lfYD1sgu8lnGUqSoqhbEsvv+uhvh/D7xdRMDS8NpGy9VNj6Qv62ubsugjR
bn+0GRkhjgNKYY8mJXHOoGi31t8fv81HouTZ4Sjzfv10y35WOzs5t9YyEGqyjkSL
DXOrTGCWviDxFyc9t7w+t+JBF41PT024x34YM7cRn2wn8v638efd+/ZfEpNEKtqg
UCllwI3WzFvj6HgCLaTrQcJyvhlxKb+kLX9MUoyrHFA9uMGDln9PDW5rDLl4JyAQ
dlNqxKzzwxAhzVp+NpHzXLUDIDSXO2GMBR0S4zolX4Fm5bfAyaZbdavXo7uXtnR2
eozcXR+3tF9dSKIkVI41IaOXVWyKhXAR3e3gEeeIF+93k5vlKx9KhJ17iVL+73uH
6xpveyELMRHvi/2n6LnHvAF04jx3w/Tzhrt0Qcdsy1QeV32irI28kNBDP+kLrpu+
PkyGxn/ymY/LSTcHigMEnbqKKAd00zOMi+Ftb7IyHRo8Ni9Hg572S7FLKY2AeYq2
CriFCiNE8PzNhSNHwbBvr72muQ4jDVM/xvMqEmHOaPlc9ySVxv5QFkDSmS1pTqjX
fpE6L+pYEHbj4+Ay+stpKMB7oKVtnG3mxkJ/asAULlg=
`protect END_PROTECTED
