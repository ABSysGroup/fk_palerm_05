`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZkRgJGUXAhX6TuYqW7kDeCla5p3dXuL206v6yNUP/Al/FcD2nPHb9tAsMbaRjjvp
Al1BatIeaMtDCtsvL/iYs+eB7RG0uwcTO6GnCBVx4Z0fi4sz9wITByeq3aHiz3am
tul8cDApyVFM3h/VLIUNFyI5GMDF7fBnWKPyi9EJVKoKJ0upzMvDMSWtfItRYTjj
/S/GeJuBX3JM1paBwjQMt+0N36O9swISn2wpnbXWnLoY79tXDm2uftYicn9G7XWr
KTzgGhJbXk/bUILFa+wCIAas2lKEKtfLEotUGASU/oBeUUB3ncFgnDszKtDBSNlo
DzK3kQE3rvDR6VscKxRvXzYjMBQg1I5zCbYLVfAdkVspKL0r0fxCdBPErIpqglUh
IG6adKCJTZttthY6mX9r9nwctOSiIh1voMleR2Wo949pJEko53bsxjMXiyoBlvNW
x+n7Rnqt+R8T+h/gJSjVPq9QEGwMja3GwYknF+NaiZihXYfiyEbCApLdl17UYsun
+QYSjeOQd3DhJ2kVSEnQXsB/enHQi8TEoAD3RX4XFgBweRhK7rZXpEmRkQGdoMCT
1ZuhN67g477lnfvC6YMszRvRWTaUx4NthGtQ1K4SQ7eEroAyml6DkQSSc1N6u8AM
kcwKz8ayATQbAcvUMzIVhOPTcbwUhPxSvI8QXLGQsUABDv36g8hx4aisC0JKpXca
7AHJwVd20MIRqc7uHkgPer913jfElVovkLYLQNOecujJ+UPBTkHkoX3t0FVjOKS6
qz4n+lNIFeLreHOcqQduma88ouLMiR68u+y20nzk6Mime/QE6sUPVmCrcarzTq46
9IVemDHA41295eaTb8+TTGg5kzS1OnXSEdbYL5XQsuxVgQnDcSdFpKhMpv8ery1G
qKQ8C0Nc5AZyvf2S80vtPLtqTZKMb1r0ACUjWsW6MDiyzW1Ui5719mVY+3x8OOcO
PLFNpNoOBq1q8YmKyOUqqb3QQE0PYiAGcz/njYXS7a0k+s4unWBb2tvSPoy8whiB
1PZ1X8Zig39u98dfLU39A+mTt1vlqrrl2y6R6AsjNbk=
`protect END_PROTECTED
