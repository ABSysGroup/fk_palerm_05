`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QFGyce8pr2bSwDz8U4x2Max2+614Wh1a3hFUDchlgLA5w2zZ3aJT25FiM6Az2x0l
Jv61kGGcpFUdjsEwh+831RQPh2medkvjjmTHbD5yG0e9w+eknMh5ebHcRZg/Li65
AYesRQaupXLiFck2PqXANrAZkyOC4iezpn7jyBySYBJZF3b3Kcpp8K8VwO9vJoCU
wzF381HCOtpLxazR6TX6Q59jioCOcYSI/sdKz5mL+FvgfHCrg+0EpMitEbkOcX9G
OuSJ/yGZHI2AAMT6QfQIPf0T1S/icnXZThyKj55SSw0=
`protect END_PROTECTED
