`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R3CmXvyCx++gRhKE6KxS4LFPOCudTB5tYxJlNtsrKu9Kh+YfqLwP1oU3dna+z6yc
uGKLnIpW1M5mAb9w58ILIkmOwauGH0y+ECNX2444r+3d79RHhyGrTVQA9hBHzON0
mBc4z2ZmJSgFE597QFjjEGp+rdDXSbrOTjbbfCTCSgyEYt6CjYebBpe+E8yMlP5D
7c5bOyjR2NHqLDIJ+ceP7KtKcGherJ9WgXqRSeCjYOWpD8am0/cK/ZZi9mVKyA0L
sVvYjKcCkfLg+DiVl3PBxBojvIp93d0yJH3fziW44STVolDd5/4kneuMpngF6OEH
/1g/s3k7lyNWJjOy+Z6cbfEiy1GA89CgMXIi6kT91+t4hfw7Zi4ocNJFezXGNbjD
uNv6Q5fKK7IkBAPp3T3aFBgGlcT4F/qKGzAS7YAbrc8pokNzOgLz6rNfIij2w+o5
iDgvf1uTfZeQP/TP+CacxPDuk8R3C5vZBuEvfD6V6nrdGtgQeYDsNVFqNsSVakOT
94sSEcpOr1OvqVKCvBPzd/oqz8H5gcHNaLkejoptb/jln9125uTbYO81jGRJIAEg
Lsyn4NuvmbMppSBZM0RiFWrBgMeZpCpanT64Qd+WWhVzp+DUJl1+MtpTUbwqDkDs
9QKRrG8M579CbHfE707rQVV4IZ32uh6FToNSuawTqUgDyO1Xw54PC/IOAq9wa7T6
IGpXAuWdR6FyVosMqHnyxmRpfRfs/CYDAdHLDQKZTSkSDipAtsQD7YHi9oiedwc+
dcBQApNfIg0HgoPbQmeO5InllLiUz2Aakq6IxO2KSNStAVc4fKhfBgLyQZOi3ciO
aZoKgJcNCaSOE16n8AtMUbM20gHCaUyqnPUwsiV+H4wxFTMHqS3gUixK6gfat1Df
wx4xtrkBZ2/y8tWRpXZVoourJmlVYzh65GgA5QXnrPkOu4XsZMcZuj3JAxF8hInq
3L4nLQzcLB1fx476Z3ZKxV2++ZIzSVhKWGfbD9SfbcaFZ7qyzxh55LzRwmM+ZHa7
PoKRKxPPIAh5g7YXSwyZiRCtwrJRKz7C8V7fxa5lJdFy63gGyNVmhkBUMOgYu6bl
YT18oItssqbqSm/8YSEzSLZClX3JCdt+Ao945U1ShyAYHJdNlKscGuEkuS1O5fwo
tx+LXnD5nvbYhDsVXr6UOu6lRVfR0DJxfwz+r7/cmsXfIFoajV1yZdqkdMa9h2qO
rALpIb8UQ3bK+2nUCfQh3PCAGkbrng6SXyXwoGztD09QFKKWC/wbAarAzXG4Ztaq
TWMWWdW3ir9cj9JaCT0vZhJ5ll2hpyubfd5ZXdDNhnwDHEeRRgf/S0+YxaIu4U0+
3ozkG6MPSul7Mw+tfoEqnMlf6mKk/4HQVzxQxDAyyN+9jCgzQlY7bLkIiVKoJMYG
NBk7cQGVZgDNnv8jkucjhompjP7eNXBCJqmyLYgEPxOCod3BGkqz7ueTnk3O2cjO
/h/E0xEZ9iJl9RguWKeswxra6CAxsTfWJmchDm/yHZ8sUYaEUdI6WnMnRHBwp0d8
FhJAFHtebN7bLYkZxfvGo62y17RRK8V+0Y1PCETbyex3VUs/iQdtxGP12pWmWrQF
WSdJ3E/jsNDK3Z6FPUSHDBunBePNhsrfQEk9aUTkpKaZEo999TOQeAIsL82ZEswR
ZGXneSgNQHZFxNPfSOQGQw48LbTnorAx6lOjAKaGOGENEI3Q9SbnCKMnAAvqxUKp
XE1QXRbCLhXGozv0TvxvyArj1yJHu4sfzUftbqrx5cCQC3MsPSvfg1nRgtmhwKRO
HARDAN8QeVPwbPA8d/ZMwI8zKtHLc/o1aV+kc+GVXsQnW+8GyvMD2ZeiiRWxychH
XmD1ze3KiNM68epli52f3K8nvPGw7DAWJdEJgv5HQ2Rnb3xRYBaAyRfKb55ayrPG
Hh+vaC0P8NrwO50J32pViI9Lerq/L6bM2ShH2Ax70DMo0z1Wb37vETisWD74VWXI
47iooL/9HxXzUN7bVq1DFtsTgCQdF/j+goVaBPVgXdsONJ/Wr6BDaOIsOO7QYXoP
s++46lBndJ55vVqCiq06LFWmN4MqYRfMijs/RpBmo8Y9E+4Z2KelDQFSRE18e8Pe
aB4o3dAoujRY5/V/gJwmZSPfSN5jcfeK3f0Qh5i32ytvdgqkAuK64/xZsff+wv3I
oV0/T38Xp/kq/opPsE5IVhD8lDr1HzYduVUiBggCF3MfMaqFuXfvu8+EaNf9rriR
5iUtVKzawtvLmYQFXwMGGUAUbvTCU1mEuNAAfG9XtUllRumzbiLKrGLhke2qSX3b
Uo6IYg3a7VClwoCdc0kZe/0lNsA4pXfvoow+eMxvloFVyT8rq5F2X/B7tjWaYc9A
umbVtxCzKjU9yORFy6V6SOiKds6c+NwoCqqYFKYwcuB8ZgJpl5tr4K1uhxrmCAoQ
WGd20oLHlZsgv/6BfBGws9EiCf5+euAYfuK28KzfVCDoqdzG5NfZzYUNywmDWWl3
JQboXgb+TT4yDbLge6y5nSR3PZJ9pMxHJgV3ZUOl1SwHYTANYc+Qn+hUKZ0XybVW
BaPmQLJrnUloeYAFAw1Z4ldS08q1TVh7ewieLdwKmyiNMDYQBT+YPlaxWN1AZqZC
mRikkxIQCalwaiheSh1zHG+gnQlO/Gs9NGcucpYCcpNkh+yXeB7HvP2cJ/fko+cH
414eTDG2vNI1NsEGo/Q8lrJyhX5zPzxHErhitFolZS9K0g2nEQyLncXCTCj32fJC
KNkJaVN6sqyuQVZfgqQ1UD8wPdA76egKrP2fY2HBXji9K+HqXLjeTBxDb2Vk5aHH
yTKRsCp4aI1dm/hCGkuTM74uZ0/oRnab9tILghTlB5StImBL1tOXXt11z0Z/rqoK
bOr/76cp7gBFEAVZ1jSUM1ZLIXButFIu/mxHpyDor6IRmLfCBez4fff7Y2XhUxV+
aLIx5+zXa+IUItbCPyzyfLuSsQgwAnuhJW78yS4haD42IHZVyM35ShdqX2yFX6Jv
R2jwxu1C/OdXKmNErjCC36p/wug4el2H7Q5hKJscAa9rBbvJr0vvNbqFd/lh5QTB
ODAy4sL9Jom+P6UuXv4eGZ/YiahplDiCi/zZlqBoWfl2i4yApw3RmGbH1dlrAEEN
cW3d2oTY/iEhGy8FqTc2Isix2/CqHCwJQ18/W7GGyTG7xCqOsgqz6A8oLRdueaWz
oi+2CWMONdqA4B0ZewSbFIuq+if3veXp6VrZtLUqny8mWIp91Dl6QxdbuMypU/pG
1zhRiShpkgx5KP4EXuCaaDF0iovVSgZOS/tEdu+VxL9xYu1VYGd2RYU92LISiYC7
ahyBOUlkWJyvlxR6ElM7QcH8U7FjFoStRcOk0odUj9ZgGdpJCvcXlBrzDmid6m47
ATmyonpHbwNsfLw+rtf3Zmawz5FscL9Xt0QOI3v/0B8qg8uROItjZLr00rJw7CgX
20HBNRtY0ecqRfjYNriAIM27la4umQIBqP8ISV2RhgMJfH5r8vPj+tMxpLs88xws
DIB6fTAiDCHYPnLKRhFwgFQesaQ6v1fjaxdP2z9AoMxXAlr/YpPGDZYaPVyS21zy
xo1T91KO3fBGiYwb83nQAS016TimF6uwPqxTNu5DFuhTHHc4Hp2UksTMhvU4KE0Y
PrrCMogUirmDIRVtAy2ALUkAJXEVCeiMQdw7Kx931rA6xqy3BjhGkrJp8mYS75/f
0VmNtYiVCysq9geDgg5j2fGU1NTXp84Spsw1XEe9de04CuwvESCDAbOPs/+GW9VD
H2rR2JZFxNrYnuB7wDwshyuhTqqn0ZYcPX2TYwv77C4ZhimDkK5gx87R7M23qLQn
3qhifr9rQkflhwrotUjev5mSRs8G/PCfSxtbAYahMFlxmXoeR4YG1D/kyB7FylqB
ssfgzbDqE2KrwYGRQP4jbdNvByUr2sa1NOP32Ql+9W7TjZz4Wt6ype6OPk0SXnJW
YlSMkbdNosharGHB9pkX7VZHQPEqVFHLPNTbgWHNuWJhH6ewq1ymXxSCmwTkmz+t
SPvBae464NP8B0z9phkxVmFhBptBBEp3zmspj8O+tIIjiJDVe4W2FUbyTkgC/zUN
HiG44yPAAd4RbBwOVpOkkFGPdPoQX2X2DWG40CQ5f4DDgEtGEbHhdF/bYrQP1jhc
CesoUBf9MASsG+xNejn9wnGs0AugehxGeKChwwkK3nWalCC9pt+V/U5egcyu72FN
yB1QN7KBtQNxrMZG/pRsjgGVxJ9Yo5/HGU6JyvZcUaFW8OlPKw2jk/OFYMlmGTGp
m9Dw0zHkSO/PbezsWsD0iInxHYiTHpGaPBDuq9ITtYKVmPUzfWtY7s9vimhgzSPX
XigN2BA4e6J/FpBhf+8n8FwBgZQY3MfhPxbcCgECQkfa/sNR5+LjD7qCzcou/gJd
Y4mb9Je0quo31uw7hNJcazTpeTPjr76RVOYUUPnsX9W2RzZF0UZ5nItIXeC4SpcX
19e1nAbH5cYGrcn97b/fXYzxK6y9Is7UX4Nu4fZk6Zn0ESV1eN8sKP/o6FddlOBp
hxx//4uYIEQP8DkxMM/UyuXhkDmxv9QR6EV+MLKmy0hhrJ7umbxbad4mc+984j49
ICCZVGV5TOobIgy35osH3vrsG2WRsjz4AtHfYfWaWLCSlg5m77JrVt/c3H9OyN5T
mP6S7mSdjDazDD1kDRx8ghxCPIPurxEFlUmkL3nT24uv0FeysAzDUhBsox7sWEGv
fvDPqhZ8EFt965hbP7ZpbvxftF9syCLQv5cjG2O1Vdpd77srT5mzteABm4fBvUTF
2YA5k3Kkwr46KWPWAefQ9qgBZUBwBnpVWGK1MzZcW/VzYi2hj30Q5e8beH/C9pZt
EmZc32SDezcswNZokU/tsnIZ9glZtU60pzavSUT8credwtAM5ekmSZkMq3Ut0Rsq
Jbdfkw8dXABEndRaWWwKhdkElX+qXU20JNbGWD8qn68ljfEj6bCFGuzXqT62AhuC
a6wdZlQ7uyms0pPsr/RMawvIHUsuLIDzUce61UJZOSkKlgFz60LE9/a1SwkfoGAt
s1bIVp08j7/7BD2yprzc8nfbHdFeAMaDYmYRyHowDCmbeP+n+MiSrrl7i3p/QDM5
ykRqTv6H7gkrkMic4Bi2L3VJQ9xLD711rd6yJB8MYWf0SRNyGmHwBCtcA+mWo4tW
mWGcZaOrAIY9SAZQCAIonQw65lofKTLTAOpDIoW4mRuec+LqQgwyjUv2iXozkhMn
7v4/7xmvE8Bw1tXqZUWjrJx8MztWNIxlURmAxxZc8UY52vpojhNprvFKrNWS3W5I
I34coDqpxh6TeMi7kj8JihIFuX3F3QE3lt53sJ5IZFinlXy7FjSyDYFIy8DibCA6
O0muixciyzOuX893HBXTTV6F1hiu4v+eU/Cqp4AbPXmkCp1QZWeyYKZz17cxDah5
3ZlsELqrqtDc82KCq96HSLlw9Z9lFrGKk1gPrhMaZ+tXCCtZUwH7XLgdI06Bz60M
02nLcCAdWSL6jXRd4NHBlmzzcq7RBhHG+q7BJuDPIpN3SSiYj1JSbVnuPBQyPsTz
5ujgTBmCCa4f1Z3ZuuBYnj3xYg2fEorLTgFCQHpqXvyuvWvOe83qoHzvG+W3m3gB
XkgnNf9lzJcJwalkpzZJhPRQSNTfCYZDAkmRnBev/Gw=
`protect END_PROTECTED
