`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TXYyEjQ+AwqXAUtk1VZHmthOhXPz0lgwxyzVb0wlJ/7EneCJ/k8GdqXuBLOiyCB0
Drf2g0nzUSNtfA5xQNzibesfo4OSJKg0k15kk5EvlF7eSNfh8OyP3No6e992TAZ9
QQFpsNtCL+l8CcQije67nPLOB4lMaLScHe3ifbEIkMDU9MRtW9XcOsD5tCaGXDHi
OHChgRhZ9jJfA/Js1aWeSP5VoOANK2pJztBWE+TrcwKU1OZt9x7maBCJHxJ9zb86
d6PmWIrhjL17sTWgyy/B6J3xkNLrtQ7jNFH/1wn4MN1vh2M5843GW8lG/LimO9HW
eLTo1mzPGDA+XOkBnc5WEzk6gnphpk/a4bMlTwNUVGx1MlnK3qcXrHuMpUY85Gie
Kqf/D5xCDDJT8vQ5w5Md2bl5bam5dNYHxwuveGBFrNTlfWihatUUNFJCzOHlXfko
aG+fOVwSIOPpcgUh8hObLoZUOof+TpSv0sq9f2ogKFTfsJVJzHWCUFMiI2/8KZWM
8pgTghId+r5Cz1DDyIxEsxwqfnG+enrbiKo6aZ4oTQB0tpZ/TCzdehzMDAunt+N2
M+bOrLniow8WCaRU8dKGZvUFVQtNmW3sz8NVLLd3SiiwHVB4gDEGTNqr4eadXOei
c7apXmVUZSWm8enXU8qbgBgaPSwNSaq5vvXJ7NmDVmyLX3xBxYehyS9AWav/596f
uSai6yKVxXmY3TQML7RgIP3s3Zi+sLZ2lTn2LXKSv5IDQpuGDesFsLtXbvokQnHT
hLE4CMkSVmTQSq99Gptpx0buATDYiD7ZYGG5oVPJW7Qd3KTNx/L94g+caoh3hnDU
itlsVyQeZ7Q6L8ccQ6x6wWB0mxgyiiON/UC6nYG1x0mXtn9vKx+MbvdcwuCI3Gdj
Hh8zwaBL4BLREsrZVK9bXAczCitzfL2itibMeEe7HqtSiEXdLzhRCCsupu/LBpgr
yKuK+CT46HXJpfBpiCDWryZ/q2RroN+75iy4oXeFPz9U2o4XnIzvTKf6hxIycRXE
C1QhJoXfDdldwbk7Nr/X5ucgu3Spb8G50Tj41ATq4jyL/3vwlu9Y4l4fFEHPdhhp
LXi1qfS37Pq3mLP8Hnhs5OOMasxe3njVYWDpaZrmSP6/BVnsB6r+yKr3j8axv1dn
zTgyMb/o+oezPt/oeNRFEFqoYy5SufZLcLlkjF6fxXBF6j4f1gdMvZy6t3lFuRfN
mKJtRbIXkWfr8nGgs2Ami7eOhHgUmRYFQ/5TevsOPzA32BC9bhNowChJSEKgx2nq
EzRRf6cUq8Sat1wIytnbgjq+N93mNUxjyx1SNHFuP5Cqm2dTi3o7rqLByUOM40HM
yzWud27zjOYWEAa69d/QKqnfrotFMsHP6rQzVq9JK0BiEfBGetYIKFk5zVKk6opT
+2RF/NhAe0BQUEawjM6kdpqM26RHBTPI1eIfMCVENLc4JMLx36QQ+89FsvhVAVOS
OMEU1BhvAveVhnTG7uW7gsZ/Sc6rdVoQroE36V1001WeH2zZhF+7tr2U9m0f652w
0TjfuGdYk/AFbtJA4En4UyBt71gL1gdhHLLgcdzYuxutQ3Cz63ZInd0SJP8VArdI
/X+lGfRfmgIVgLC7ryncSvYgCzBiQLn9T16sLB/vu955HMkJSoVet/VDrAvJKHAw
y4/Oe2mKtVki11VkAOubhF8T6rmvHPHw/OPFQgqWq9I10GjokXHTwSt4phhuYAsV
BDhagD8LSp87rmq1XvWIVrGB5PvLAwroZIefeSiGG3IAr7Q4qQYETtRLGWrEpWQx
iIn7FchPU9Ae9BPq3kWKp0ryShy1uJkAVtaWCYrhUcJ8UdLLJKEoFZJ2YkFk2aEg
zcI65HVquwr9Lh2PJK//QJF78p4IbCUHXkM7A96oKHLpN+0L+UyOS4fsEnthTGc9
ELxuUT70XuJXP9wvcGycQQ3wie2+ryszLqPFR9hyySvQZyrAL0OEnKnrD0cSkbNM
8vevW4erIpDbKJ5mItDWiOoen14wmTc5IF4iPXAx2697ic+yGQ6EpPGrV7tWurWM
cxr7XCIi0E7b3/Q96KKUUS+uum/R93VbJSF8rj0IeqvJf+8bN5GDVuxaZU789ZAp
YkbTQUwP2KnSVSSru1mVdBxRrO9yuBV8T08g+5wLnnKJ/oc4EaLv/LpCGgYtDF7I
DMEhqkrpJOae/0quV+UNR8EtgacHJddAemHVfqQJLuPArDhmLP3TTtn/ENXV9+X7
I/EcT24bWGAlybqW22Cy7D2cADjYbckz+MAYB8lSa6MdECE2TSRhu7Qv2NN1omc4
PL1mjxp2ZwFSllEcOfyMzWyJt3LB0u09Zz2PtImVw7R+SO/PVNMcAhDyA8Qvv+Xj
9DuwXEDQyKd1/ShNhQlRxqo5J4R49pwK5Uw3TuxirfuanerANDRLQ396YB8HDKs3
lF7aVSrfgtT/ws7Q2+YNjy8nq4hz6tmLmqpl7QdDEMVwVHBcjzk6WD5QTPF6ZJ+M
teabAznHinyQeKnBzGcnXNF4ieMuaiowBC0c88xnTSlXM2YF3MboczKa3Hag6qQ7
9dOR98jqO/EWh8/g+3baOcYgIr/WoRHrRA/GJi0PQmZKPyV4tyXVlOY1+uiNWh8v
MQJe69aL+9//nN4WzG/emtUH0H+yKrAe7t5lU5Cvg0SPnsS8JE2ICv+3ZMWKnGwJ
1CNEmAzYtEOubT5uJAQQx5E11Axv8dAa5oAg7raWBSzoBZTlJ0pNNzfmhmJMVUFd
6tB+YSQTNkfuQyM/YN+8qYR8a8Va4D/IZXVkOVQWwsyklP4G0a7sg2uzRoj9npBy
AQqaioWAgRN2qqe3VqwSzYjrYTOTr1BCRrz/xbAQ3/HLuUaxXgQWaIh0+d/6BYgc
GkWEVAPE3PqSKpkafCd+CDFER9F3wZALDm49IW5EIgNpA6KvoGhgQFAygD3azzpy
V+5wjJiRWBbd3s75V1PMHb8g+8MtTK7m8CZKX6Tfl7dS/IncDADg0oYvZG2Ckhqp
B2gCcPrLd0gH4JysCVcewQ7Kivn83jk15JSjDk94TLWXJ+tr9LnJdrciFCQIk2p2
sKDnFTCCwvklg/glbRG0i6quycOa9hM8TZOZgOGIjakRurKvSiAYIPguZBpi4/UL
PaCq6O9rzDdguo9OdcuVWeZuGg8TNLEQRcFhR+NG+Bt3MAKaBG+0kpPVOmVJ3zPq
DnhnFmnb0gizIn5eu2lUr+6XDtRIbK/OgzwixjTf2w26DhK59W7bAHSQHi0lZSrI
PiqgmOCrsPWgWC/4CE6YXp4vqSoP3M/uZRVV+kM+woMIbKLguOfxkJ6CHqiUs5qA
yc0JnMMefvgr23g0Xb5LhpFDccXXOxg+8PsOCGLI519Mnx19gm7jiaoBalNeJEka
wuJ+yScaBMAiDH+LWBsKSm85tRQd98ElC76+hC3cqKo=
`protect END_PROTECTED
