`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mjUpiCnfFhWGTYATWTLeVuMNbYo8Rc3CIsUH0Lk0WTwkqnqHETs011eVExjjL91Q
Xk/NvvyhU/rNPNe6Oo5KngqdihldMlQcnnuR8W/ixeh+sVsWU2PnEQMOdHDWEGXY
Qp2Tg83dbZN+CXWYfsMirNGgPJOUaionmaTBI3rd+xoFOdf950SMBaUPpb+dZkyA
x9b8dehi+aYAU87pYwffcIOqhkIl157hv7VlnGLVV5XBjkYxA3xybyfZ+JV5AUz1
nlrKbFClbyhcyw/k+Md7yIrgvgxujqxNOn1S9djd0jiFQ8hm4VYQTaXM95JVip2R
o/bL94Ghjr1Ea3mc+G7Ka45X4+FZyqabQZ4Ovm61u/4UQXlcS10qj5NS3/WSsJYX
9iDv9OhWu+SBSymcm9Dj7CB+JfqB8e/7iR3NCdAl5XgoSrG2ETAgdFtAgxz4Lzhe
F1PfYhjOrG40d8kadon3YIOlkZqcidM/Rj1q9otSsYf9Y12ZOTsCEIFkBpYobYS5
KOeCN2GX1bbaePR/F6z4Zfvb5L01A6IGZy1gc+IbXl3QyN6mGqCIbN9oKjqsE0s3
8FPahOZMx2h2vMw9hxl34zudLbjNdgr/FOYFcO/WJ42r9wcR7IfJYkkMEl3oYDgN
UhrJ85nZLxdcFqCMHl6fjQUMwxYNA14Mi/RIHUgypTkn+hsvO+m8eD1L2aF9GpL7
i18o/ST/wlJSXVZEvlI+wA==
`protect END_PROTECTED
