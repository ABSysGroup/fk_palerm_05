`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+8t2yljVlD5r0v9sMGJYsmYu0yAato3AhBtS2jyAydH5ekIaxrbKWWRo+pDhnReV
V3WAlDVQ0W3XpBAMr6Y5H/KXBJ115pAiqxj9xMaMcyaB8yMPJ0z0dg+9mqxbMBO6
4LGm/zWYZVTC+L0qb9CajMHkmSVNiWK2hNyLdR94kxu9ilpkhu5UjKQP4KuVWSah
Ygzvpnq7gCP/kgZYXOjn9e8X6+aecmdIY0G9haxbxAPdjyb0NMRMuV/mQcg06Lqw
AB4/sSbDb7/k4/P7wxUufdypcPK4I0IJbfMPM+Gmh95W0VU2NcMFd8rifEzMFhUa
40m2WjyKos3fRdMg/9Tz1TJsn/ngI7va/piuEKFK0kqPCJinXhRtGElV3f5eLX9c
AxH/ZTWax3sJwK9c94TtXl6lmE2aEhDxzW9DrTSeXTDSJrF5ncZl1QfQQS6+yD8I
J2F6KXlhQ38o4KBSb8bNUw==
`protect END_PROTECTED
