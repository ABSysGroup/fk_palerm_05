`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0b2xLOOCfQrDgRZUfC1v1py6WEZNTyxy4n08eGkfUpjr+2xe69ErQpMc/F0Rw+J/
E6eXes09ZazJHsTjBIkxAfGNS4U21t7jscgbnZ2HWKYU9nbw2sT7blUFgEMPu5qO
G2pg+ngdDfGTBB7dOS3MRXIIOUFI1UH0O7lUTWGaJ8SHuy0Odeo5PLhoFmmA4eZj
1e158Lky5WT102DctT5XCmzzuWF0sT6XRY3nZHJvRNE78WmjkJ9QQe89q3zDHuyW
Udh/spBEFAHVGAGMK8zmoe8QAkkR+1PuPCB7G6NdXJXMf+DTLdwNEfUC4549K9AZ
XK0TSMcOU6D0s4O0o+hPJq+ayvbOzfhGDIl3SOLJdnsfpkbeNR0AFqCavru+/vLp
pqjvwiyof/hrei+CQUZ84i1tbGazliebefyDQ1tk2II2+YWphOUOrxgV8i0kHKFZ
1O1mSPNlfnwXrkJfkAqmV/rKjyxLwBRjhE6DM24MahIhvOtZy9eEHwQgh09AVCyF
F3ckglZ0Z+ue3ySJNVRuCDrr4Mzv5CJ7iVvBBhPYZ8SB6BB6QhtFhqPoK74/5+Vz
mhsr0JXE7hxlW55lz0mA8HxHR7n37CLTyusYHnCxjmGkw0nawIJrJOabuI33YoW+
qr/ij1wrMJo9htK4QwzwMyPm8DP+SB61r5F5IauFwWLYiVnNY9uwLXbhgfSjYgbs
`protect END_PROTECTED
