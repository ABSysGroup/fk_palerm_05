`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hsFw3WZrVibbVbWsA5xBmQTPaw39GPlCw1wU2+5srwieldygOZmMUe3hDXX66NcV
MWT4Jd4b86FYlyEszyXx4c8Af2Au3SVZQBUC7+Eo67e0wapAohKorPVfIt0aMA2N
9Q2e5woP4A6ZDVqRAwjUnyVgUIT/5FfwmqNoJen92QOFF+HjaPdaeCQkeJqU26Af
HtWScKSrWJCw2w7+fJ1S2B5WVgJvtVzoGz4f7Kj9mFLe0xd15Y46CTAFoIj4JpOB
jik7DAInc3IcN7oVVMcQnax6prwmHmLM1andCezstT0bg0CVuFIp27LPSsFcoYYd
uFETHH28TXaha126da7HnVoX2jkHmeFazPOaYllRLsRordQn5N9GcjyUTMK3+w3q
7mB845KrrpDgkV6tnCzOXf0DG6EK9TDn6/NRoiRqkLkf1IikQ43fVi6+30DkaDBw
vCoujxiNKQfOGOClDzOgSHNpybQ1ZIKfv2I7t9A5qSduduKudZG0Y+eq9iIJ5X/N
1lhFwITZmn33ChfVXcqeToF8QGwLBC/y/q19t6SRORABfoRlMVA2xAojcRag7l2E
vTUca47fBcaW2nJtwEz+F4uyuu4xqih1tkYnBQpsESifVgFY/ee/6Nk1RK5icrJU
GOErUKz87WSYfeDuIT6VbXKULWNZo3e3yGS0mfic1wzKilRW3vPtamGsBFVuogZ1
4HoyBs8U1hYNm5px9JRRBxUFz+YxPbKi//ClYbZoQn469/t7iwhpOkDckwrMG1x6
fM9GBrE5KkOY8AVWhiHI0FWCBRJCeX8VsUH4EYt9cen88hu7Mjx9zujLeK79ZkLF
7y0DmlWBTDQGdGY7HXEfvdYUJ+t0AJW3tDycrciUvBplBhhtsoOhhLiKdYNvd7Mk
gcQXePro7gbGLe86qDrnyOkryka27ayACPFFCPyFr4OJKn93Lad50EsCZaDDgYFK
vNjjlRdhYnaNDXq00hUzb8NKko1+NCfsMh3/eC7DyFFgabi07pFmO8ecBKb5zWhf
R49QM7zYyfAkaXI9QB2mkZhKJYaCyS/W/3Nx9iPXvhD968wJ0ubG0z56SVCPxP1G
uVrU3ze0TLGNjAdlPrHGFZ7E1lJ2eWXIO5b7Y4EKquoEDmsTVwO6SIIlCPpBpsD0
0SeJaHARS+az/RfJs2c3lxwtfdMQoBYlzqaA0xYo6Dj79eiRqAC7rSGa0PILkc26
BA1KFL5Onzli9aX3RT2nfsTjoEuGo9fg/m7+qCeke4XcD/q7TDpt7EDicnhrw+J8
re2UJJfXEcf8zSAWD5AOd7i4nJcxEtLNB3NNieCbgiNuSdmc9F7X06z10luTMqrB
36RPMJu7Jzjf/+PKcFrBxvr3u4gCn3HobB0FTQroLZcXee5LwK6CrtBx2Tm6Udnf
z8SS8yUtjLtVKXW7hMwjT3b8pfhLB3mGhKN7k5ZTE3Q=
`protect END_PROTECTED
