`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rVLmR6Q+1TISWYCRUzb1yjCVO2AIl9Nl3oW3T5wycLKHRhZFWm02QuEdcLx8dwN0
TGzNTz2vVlPiXMlNUtAGKm28gYvSrb0HxEvTyixcifTRmDeTBuE0zMIrRRQ/B2cp
k4Rsr0TxM0k2t9D54KclKUfA50v0We9tBCZmZlsMqb1q9r/i981o4l8WxHaMJ+YN
ZL1fRk5ES+fASO78smFu6Rm9jmgeZyqampCzSAveSKCQP8Iatf60eJcQnkNqVLxg
EywWdGCY/9NyRIHmMtvrbSyBHZSewou1HHjvWUCH867AjsCj5T27O9Jp4m1zO/+z
IhzV9Qwj24paZrz5ZZO9tw==
`protect END_PROTECTED
