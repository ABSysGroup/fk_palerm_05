`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ogpDZthbhwAaMxfMP2P1upW44wRl/9VAfXbEcp/e2W1j/w2oNMWiqJFh/3onIpZg
2k219GNqt8rUyfMhhU5D3UGzdvESrF18+NBn5Ekq3u8R1xRCYKgzduqah+qbYySV
+wKxy1MN5fiYpOafOAAbcl+e4eMEZzmO4ru1fYD9rvI2EB7qj/aBHf0SV0OqOvNt
DqtrgoDXAcOWcO7YjsL4cEBF9OpXw+iu9YhKS3JHRaK532wAf1sAeFfM3cSFRRlw
pzlezMIdnVS2+IzX6cDR2v2ZlsCCFc1hHPNn/wFBOJPitNtXiskyppGzGTDwJvHm
tTJkq+W1qCBgjg++ksfKh0R8onbKDWsPw4TFMyL/mqwEsW+JB+XBQM2CCTApXOVQ
YKa3BFO6orZbGgLUpn9yrokADKn2xhByH+Jv57f/2WkB1XFmOyNaSqge6P+fmkxR
rJiyVhRyra3qZBJsLQB4YWhe+WQIKH68cIzWBz2jko+B6poBNP49cRBBgYdUL6M4
sh0rkt8BopXehrRNEu+4dbwdVBzGSFyIXFKhRbRqlzGr/z9m+8GhiJ83NRHva2BP
j/gs2482XwZS9s8Ko4gNmPIwCrTpdBoyqtZBAB5FvM4zwv2ovBJIiyLD7fJ1FWsQ
lxkPLO3GkXepjth0e0ni81kLPwL4uED9PEBjUFLjwhSyg9f6ob0SVEsJ4PY/PrW1
n6Lg8M7i07GLzz/cmftG57adiV+amEgJeWYc9xvCcLgRJa4oDHFWoCxLaGq4WVwA
beLbqNpoJcqBdIRCsgTJnqlvyrrpTDwHnoGxi1PhuHItt+O8EznJaTrjPGhN2oLa
0IbuDUmfym5DItQEglGfRK6eyHB+zT6MC3KFYLS4temyPvKozztBYZG8K5/EE7JW
9eHu3nxfhjq6/k4qLYnqJ4shdvFwaJiiSnjo0pWntSQI1e5gleKCpFKuRRyJRIxJ
yRpzpDlHcbI9YicaFKD0DeVihvbWl5OSj99tdR/B/iPDEeIDJoxq8VW8xuqLCXMz
Cl4mG7QesfWaUEivb9pwQJH1gaWzFu7OD4leqLvNK6TzWjjdfMjLVoPQwL5CFdt0
mMVVPGru0zRevzcwWhmeH5pMzlD39eaJcbGuaZZ/PzE1nd1OPtwe5LdV2kZg8LiH
3f/Yylhl8T7BJa3QHWChPmYQ4cfVhI6WN0gkrwu4s636XvNOtKBqYoIvp1X4j+eq
qaAr2gxE6QYw725VYJf94Sphn0knESlA7crCc0deJ0NSLTpAJlz631ht0vph0SrM
tWt0oSEnoF0kd7W9KKJ9OngR5pRIf+Jtv8jwlLztTZQqxg7qyMhPi/ceh98s6JRV
jGgF4ad+KLmx185Ygf+PBg==
`protect END_PROTECTED
