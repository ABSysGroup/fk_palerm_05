`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HwfQEU641oZjgsu8lOg5VSxGMXfxBxAg/0/HEJI+YS+hMaZjSMzi4rcB59+qh65C
5+AKXV5oHi5k7AwwRj0FKtfzG3jd+WZrzJFc+Yo1h4KoN/3UFcDixR/HiFXHZIqR
uSFhcfrRvvOVAPHtvoWGXnMOxi5Yxevzx7zmcKDzkqUQQpqkXVA0UbhU4mnwJD++
9mdeqYhGDpWOoH3FEHD0OboGlGjDWnUwMV37Z6xEkSUWZdI6xehXPhfTm/mWC78i
r8ivGVfBT0StQsYpUxIWsaJ1MZ199aRI1v6x7tNfe2DOZKGwxuS3iX2JNWVzW1IE
6QhebPdI2AjtmyD2f9GBWe0g9iO8i5Bkn+zbXPY0kFXsAgpQyYTaURG4M4g84MiR
sL6cY4Mvud0N85Kr0MrZX2IK/FMHn3X/J2IR5awSWWSsYJJgI9pl7p8ej8t58lbo
YC1pkpUZ3ZyOdxLV9pp3oSDgZ5LCmPsg5UiM6424HMU8rnE5zqxeft/TTo6Lny6f
`protect END_PROTECTED
