`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hZCFoQEpoCS2+znlXs3Ztsusa9tHHJG9aLpfITw0LylPqalL7UKe70DsdtMH1+Z0
Sdp/90T69kg6XjdoT52HCqFOWIFL0F/pa3HoFtI08qbpI/X1y70InQXFtPpj8WQz
AHXEd+BPJMH0TwaPWC+DgZjf0bhs1zwItcaFFwhbLLLlshCAa1foNORj86KQW8zk
j7VTCKngCfTLykWmivwUxVel5H6L3i1bxhvAzncD/GoDA5gsstYftDpAUkwNjUa5
9QjspBbFtVsen/5fkgYgSTCI+xc7BltyO8RJmxx4QPJEx32jP2zqwV4whr+g/AoO
lvGyDQ7yddZzKG4+6pYi/cek9rgjLIMQTDX8ML3v22JJUk6Y5e+0R42iOEgINq/t
VLqwUJAM0Mj+GslK7GNDtkqDLcs01TrFNip/xN9MAJi71cJroZD4/jqDDprnZup1
38AW7+S3wrIvFoaCxZcZ0hLuCv5qT8TV3q6mLgVSApl/YlYkUNr1V9JSHNbjfs/e
wsdNWTnyrK48rA4zIOpapZ2YlxlZD7CM527RwLggdWz+CuRGXYiEEjaE0iQv1tdN
7IOw4gtKd4djDARrAY9+eNM3l5YUd2Njb+okHvXyZ7VCPljmV7b4MvenbS5tJnOn
hcVCYwJENHCqi9b+4Bz2Qk37v+YM/sZGW7OEdD7GtKfvKxX4A1LMN/xH+a1fq7Bz
LShCHyWxgccMFk/Gqhht7xG/6ynky+tUYDd893G2xc+TmzCjGPpq7YfBemGknZje
h8RTTGKUhucnulRNQ0gxxS2zcJPd4XZ3J/OO94SC/WgEEfnVgjrX1JBOc8bNzecz
piIooqJMMvU0lfBPs/ROEYYc/fpoqjjX6+D17+WpgKVF/weE1+0xKZ8DiXcf0mUn
s1V7F2m8KyDK/Qln++yC1EoOuquyy7TqI6XURs7P9EgSekxMpn2o9zy78gCdITEO
I+Jo2t/aQiidVLr3F1jV/EFdtJeq41sqdBH0854LPGpPjy+6QNntOjcGM/+g8Bey
hMCwzdCupn07IxZX4/GrL6a83glJNA3Gi2gv7SgchIwiqBatmuO/t5cjMH7+NPAa
ENf0nnmAL6ulqcEq0mBotnWBPPJhJampJXDkoa3DsS8/Ruo76QTrkzqbGKctIxAi
aMW+mQLt3+907kTMAJvifovgEBogVuf4kFj9SgLuDkK+bAiesbDszfK/w8GHkytc
W9iwSKXWUhtWXIORefsPqVH/jk0X7FePiP7QTwuoGunEcBR5QNYdBBNKpqGCQNn/
R7LNaXj8XihsYWyAaVQabDpVgYnU5/9Of7NRoIHvWIS9xaW/JJF2tF8/MYcrXAFD
GLZRQxEEXs+LlJ99mOs1kvOZmt0auyyBcE7oXNeWBG8L0ufRGl1dPCOjT8t0mxfX
sBeHdTY2tfpDpJ3Qb45ghEjXgEbrc73hTmXVwIijy16UyuSdPMsqrEgOfFrqu3Ao
t6HtjhTJSV5cNYoQH6saeuv3aHEU8S6Ms4LcDEgk2Oy3Wm/2wXdVOup4vPo+Z83N
pIIcwe7Cx3ct6WLjh9Y/86PdhlnqTisLAtih3sQsYysBf4Hp3jP9YgLw38sLHuwK
bwcB+OaZJidRRFBpFDIRiiiDmhUEnxx/UtL4Sueg514ooOzGEb3+CMfpQ7UKgWxx
QEQ1YnrbzM6nDxEB3Z+pHcgj+U6RCviq8GTUH+LBpQX8hvyCotAkFz2AttGo/Nnw
xZPEfiarPBmxO9Bf7tF1Vu8gGMYIla2uwGcjR0ixo3Yex5stI2AVRZRftVlvgujB
HPHizKsrIIbfnDfvB5mmB3OAs6kdM6QHBA9yHJcPk0M5BDa4QjvrbwjOK433Az6c
bi9wRW6tsVyRMQR2LxRv0Fm46FU78Wser4RKWL5Uwlllt99Uy6OH0/k+gXNoupXF
djWwMCRHPUUfEIOI3e0eRZ6SqQtUb+955U0dpftUmMkopJL9eCQmBcpvI9VSD2Fh
tjEisDQHyDxYwoPJQGiS8MiAsjyJkOYAY1aHyGYtvMX3cQqM/Xic+bWL/ofOAEyv
xJ8X8wNhDft9nuvao5mWW7slUrKn/fNbBpt8OLJXs5TNR4qi+I4vTThWjhis/yTr
lV1PhZ+9WDPf5SMVvQpkWSyG0OrQ51gAm1yHShafAGVfPrcLQSivkDv1JXOfgXLo
MQYdl2mYPdVzGVTRIVjtpjgHUO7Ow82Mnco+l9mX3NLA/MIQuF9EpQZnTI5wQe43
ORGkwYr0uHM6/8MN8ragR1Z1MIy3MhRhqQaKhYfA6G73GnglLDHkGiuD5TqTh4MO
PYcn+mdp7Hk2gmqj0rNukgf41X0B0T2+LS/aECS8mUe3WdRfgTYtnPUuqIkstUw6
ccIrjHeeVDJDowikSHsh/5ON89xF2+6s221a6hj1fEQRUud4R+hHsDx1Dnj4YrM5
zy7UIJJZYZxBzTsG7symON5RwHMxF/JfPUHQpBoNVv/h7keVP31LEXqTFiq/QPdY
qO9k5zcLJcPjj6RxOQK7wA+XWLRrijJaqrEF1UCdcPQoqaoJffW5wyptWZZhRxiC
bNE/pr9juZHUUHiQOiEi+ueqBE5sR+hGVxHixxi9mGixNryOlTwEHAcTZuloGmfS
XCXGt1zGNDRBsKyI//DRrzq4bfuIM1ea4pOdcxOetUcGVqrWVcxTSchXSNBwwkQR
8jiCP3h9NetM7BK7wrSwoliZmn3LRsV6ZBkV61zCaWINeHvRy4yVohdZ2c9lU/bU
sO0GoHvKLuYVGWhZSslTCmTAvCyCu3Rzv2V0jG8cUx450AZLymO3vw58lXYU7osL
s8iemRFjvWM2p36rmwch9+kCDTNd0R2ToeaKQLQpWx/PF6j5B+x+v0C+a7ZQD+ou
eEMSWSqBZevCgmHrqE0WSLtk1naqnKl3hSD/vTEbMeaGUt2rWC/MuURTHKTmdLyC
ESuYeJPPoWu0UXAs3JOKc74qOAG2bn0tEXhr1PUCPjBMLaitLujG1t64VWMuTHME
NqCTqY34LhM69C8a/g2CA9NhHbTgIohxeXEo8miWE8nS/uumuVIzPBxqVaKUqHRA
1FofY8xKq7FV4K056lq96clbkpuEasSCim7Jy5imdO8MZqK6IxCbNpZFO9RpjWMc
NpTGbkrvT9myFfmeSJz1QTd7NkVt0XgWxAA3Y1Gs8AEJAYTG69O3vVM9zQYzgzrm
+g8DyLRIiiMV4h/3Ln1rNSCmcFdHvtmj87E2NDGndj/QqBAMC6bljHhu3JiYgQhE
qnPEmolQiXx9qfWep+RDQpxNM8j3YAglnnK3d6Gbj7oYjd6bRg2IcZdD5g5jq6nB
MGLX0gIGqjMmPks49Tvz9RzEbEj4e2s2UwVAzZL8M8wIW/tSDQTOObJOpp5/Upa1
OOmci9jQ1f8gXivO9WQJObE20MmFAniRCo8ihz4jO6rahC4oqqdmTLZnzybVBHeO
LLtfxDPReTONMSVPpK26h8f+HyYMbrTDdTGEQm3OokdrWA+6cg9WpeioLwdXQVQ5
bbpq6jHcGxOorDpMO+hzPwoE7Ln/Q+hx32FWz37hZEXCmCNQguFoexCioClit7nK
r+tXRopdakBfqi+Xl56nZ6DknU/llXK5wcS/Mibg1PeMeXQ1bnEesnREN0sErU1U
3gv99Uskr56S7NWi9ilitvK772ijXB8QutuaD/wC25roS4mf5Ys47pzKygEf2E4c
77PONPrC/vsqFHQJKeyw4X+mqcZKbaWC6bRtXQm+UkdrEWpJBtzalVycE/y7fvQL
g2XwGHpy7HbHHsXa4gglcJ38tv3x5ZBR/N++kbZ5sdV8KLskeWxGDReVHd1LnFnV
AA/6RvHODpvTvsluUCoBKGLQ+r0OlVGIJfD+HNv5JY20A6iRXHvPb4y7hg9PA3Bd
YO2Ri5tPxSwpzVwKGbyhP9s9gEw738Vsvss3+cA2SZZFksE8XcG9NlJjj5XDhFzJ
a1Tm5Sxb0NWl1AZDAOBNN1fz/zaRDzux+Ac7fv16VNbFVz71V9M204QxTSuux9FD
IccaV137E5n7LcKDHgdjsrqW2RLkDdGBIL1OHZRnkBaEc3dNxzsFiuLrpIbcL+lN
mYM2g+f5zC7FeMOPOOXLVoSR4nUoJ/z2LuodErH/d3GxGHdtTTRxsLFxzHxQrLFS
SZUXYg/fF3E74LFuXSA8wDkz5MZwiM6g1jMDZKBsfZRNhGo9rhUjfqdOYLtkuDQr
iuyCYPhqZnZ/YF8skK2UREUv9Ti1T1C/mwICrmFZfhuLmNmGy5XPCtDNlgB+N0U+
cvVSqFVGevnFybeEHLVdZNVJkbpAfQCOIhyYy8abgB1gXpW+iiTJ/KLXbSY8F8Yr
dzFvi5ACuHg48oby6b2/Z63BTAfV7fMe7zJ6AHW+288Lb7RAqEBISB52+9boRWCj
sHvqBjLonL5Mlsj3Z3XA1YrK5dETAKjE2w/SPYW/kBZqTXiTM4afqkY0aiyW+IIf
/AuniMfGGaE5wDDUjKAhW39jdvPFh0K/8eTRb7KVPdR7Xa5NPT5+JvAh8I8hxwVC
M85SCVOHmttqydzgPlwgYeS8XxBTIQ8JAowbv6tBKSR7QEnTgV2kUkxGJFPZWMmv
0fgqWSQv+bRUO8gQKYoT5D+n7PeCMX0U+oP9+2Qb4MO03MNAhwUlAiBg7pG0cPEJ
iK3gSXsjZWy5nhe9Ao6Y/lkvmPzVp4Eqqwt3nYQh5Q2U2/KaRlmHtPlcPRQFeW0x
FOPOZUB2Y5FGYAHyovQHecm0prrwAihTGVvdBNMztB8xrfGh/QG6rOa3Z5g6moiO
IFKql4pAslCti5LhcOt+GLKCOmImOnoP3IPAO3EykyDBWmwto3XxSK5MayPPVHlm
n7c+ovATZmQOb6pOdXP1F7JqbAFLKCZBXE7V69RKxLd9+mkCEZjver6nNRQVyaPr
d5AKMtA4lVIQrdPRYHqkJ6VmKSlOCmQAZ12SLWd/1mhs2OkjNJJU592PoJg0bV/c
11/2/JGa7ZNjkanvGvlUpeL4Itw9OP4tfxwwTxIL7XNdIkgfovr2KcoMC/D4mIsS
DL5l0XEKX01PhQiK7jWM5zA2jahEOWeP6yTGmRvDvVg80cNawQmDkqkxOFohHy39
KKgEXIDsUmnO4EFTm7ItB/V8+klydwBG0Outd1DLzCJVrLXHQu3ScWmSusQxXnDr
+CnaO1ZMLRL358iwc5mXDxUGQxSxBXkuFSLT3Nx2Kwf1tRQFO51DelY07fi0tybr
/fefypNpsJqeh9/tmQJr4O7I4QKNDrhWdeVkwyg7Qzyvo3KsHoUQLux9rOlMwMIH
qKYYjwGblxuyDnPMO5QxbQt2kY6HePeWiJ3FwHn8U4sTwcppJY+8+zQapEiTb3L0
3e/rONEGVl8ou+hQr2VgQkh9B4LC/QNk2jk7YVgGgY8UaSnVatN/1Pn4vIUff9s0
9FxdTonoLt+Z80X113Eoc6N828LNVA4K9lr+GkpnDSDHrm47G4gGHPgx3mAgJDb0
QGGTY0oqFOJ6uh8IJBbC0rFvHg4nlLJ7hrOrsUHvF2nBx+9sdW6irTehW1eACXd+
U4iDoYQg5pcM8jxPehljUL6/oDrnr1MWl3CHLMS0ki1shU0AMVftFZPICC2Ny0bT
QQfQ2y/ivj2Tzt/PuCcO2lE3ImirwYUjG40WQqC30q+wG8mZxBJKQfti039TaK2I
f/e3DvA0klxpFd1m0Ln4yC0vuTGifD0FrO8nZK/TOraawpfyYYrCCQ43HN+OJ3A7
QFf9yzN7fMdNkwiSY36Mgs13OkUamH40As9X6sdWJMigOkhYMLzAUMJ6NUt1+fjN
QEpD5ZD8yyf+W/+7uqiCf0KDk7BKuQIv7FNROWUAXbkQ1hpN7LD4wwCP9BKPsL7f
O3es8SpJml94yiTkS3EOGORmuwaOzFrYsWX2uhjmv2mTf2Fdfq6a+y4gPlWLufgh
xyZ8PV5lmScU6yZFzogmdUWdNUppks9HRRdqQp44riCJ8Kg+I7aZmmGRRPnXsQ6C
X87Kwxs9b01uxze+N91urQu+u8GOzUZhMLrUtezhbGTUB0Gm/IIc6vcC2Ay2x0Ad
XpyNDctSE/Z1Gz9XqB7HFHUhDa+nsbtL+UYOo0pnEG3fQl9axl4I3BTpazEQOy4c
kH7dHhhNVqb6X0WgTgU0rfWwDVFOTRTUbgR57DWo/9rvoj92uphXEQ8snVr4o7Pu
IaSzNNn9p/EPl73Rzwl05uBriZp0XEe0eW0T5g0V8EmcZduDBxqhMMuYyvf8CjIM
ZA4PxZ07DOUh68MOg5Dc7O0r1xl4E7OhrtBe4v+htt9XsTU4MHM/dkCh4fGoDjDu
8KGXFg6nctcJAnyFgH2orc2DTp1EZ9qyc+8qeaXjUMioah1d1TqDaSt5DnvnUpQa
rY3V9Y+FZFXHcqo3pGfhhNpu+/ZfliM5VgLp/7dfDODGrG0UflPinduid/csgjq7
v6T8CFequLYELGikm89Blt6oS7CUZBsqQhno9u9SlbTc7+eSNqAwTKNfakJuht0y
kiXXNTFqXRrQyVHqLaNeQ6IruX3YATrhiJUR9HTUmLIrM+vQ3Tic67QRxB5uB0rf
bo9rL8Z/mep7n8J6JVjCy6tydfR5+Di3ksgYxSmYDRQaqGbecUQhT3MzfDl8O5lV
tBCZNY+TlOHi2d/rurFpqA==
`protect END_PROTECTED
