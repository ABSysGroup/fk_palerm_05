`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hJfcUdUjTlRd2lPnIGzmZpN0uP/60tNdMslXMg+Q4pjKjnQSxj+3azYDz0EF3PWc
F1HuAsEApdtTfpjWw7keRiDXNQ0Vlr+x8zn3Yl51luPjVm4woPxk6xnWlLc+cdj9
OyJEtt84BMMXC386qfcXV23FL5SSV8D4UvwUz4Cxjf0ytaco9tvPscQMbsDNnyYf
vLwsffXXBhFBvOa3u5A4IPI+oVGPtqRnNL5O7Xjs1JhOqAxR115JMIDb/nhI3cUN
UtVW51NEL8mV+g9bII2tfZFT3M5qgjLWsggR529VjUwiA3QyHPQbFOdfW5hw0lA7
b+huZ/EPPVFmshj/W4XUrvB0jajCS2fk9XWiYXQT3ahE6SswkZaNJgmFtIYHwur5
2gq2Z2SPPxadBD6wkSBGs1I3xNHqSbdDKF3u8cf2foAyCfn+7w9tkI4E5PNi+nPh
w1evfwCwYT9YSJ4c4kBiF3b7NHXmJ9YB+GisAl4wE4QHjBsOItm1ruvacCO9HpN2
jvpZB9DiOarDnZMqssBdyHf2B3Jx4uO0DnmLjdwjYbVRZeaMEccNQXA8cKUW+MoY
F2BIA5VoyiUNNf9BG4zYhA/NL/Su9Fv6jibqK2o5c/FAHABdVvPugNjerALvZn1Q
h0QLF6TDs5iszQXzW7nmGJvgOtW+mZAbg8cs8hIAzqwKApHSCgl4vjlcbqsf0nx6
XQ4Tp1gMu0fKS6YgPjbWzZvrbaM2K8HDuXPf4inypMnTVtjXBfyypZJ4+L9Ct9/o
Y+ohxxIsCSAwNvA2tXSWLToD/xB026v0QZ1dTcNoybifoWWqrRSfWW8VTwieWZ6p
0+SjIrjqqJEdrLhZCiVVBdhl/g2jdXqFlL4BFcymQJekS27cK2E+Q8bdL+bpAi1+
IiyGswbGO9OVQEVr647D8Q==
`protect END_PROTECTED
