`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IjVTX1Lx9aI46HIgKfv+UXP4DfqnjaKLVgffCDVHZMx2yyaSV/w8AgQoAPd+i1PE
WDQToXRDQGPh+KRQ4YjfXhpYW9Q0VapRuPlDp3y6GwCCo/Cx7WdxZ26SY1PSVVE6
/3wDvEtFJrO4iubzDG9uaWCx5jyWdX9XvwllnmIRy9QY0wR4Rkrt8BLq2SJT1UM4
G82pSUyIXaACIuSoJhR2S9hoi7a26ka9gfZO7DaNenpte3Xgdx1sqPoqSaNjWsqQ
MCqHXw0VR96g3ppDFAQwQSBfEFBFlhnM0425veQtREIB92/BkWsM42+QOmsOXud8
KBTjRs54s7Z3JJ784f5bskQ4VyA4Obzi9FifR51C8eQILTg9tQEom+NLjC6qeVPv
sC61vznLrQA9LHIbO1fL7oRq/kLu6mZgLv/CMo/7f6hMImkoGUkNc3cHA7e23j+m
y0X0yM2cMXiS2W+xqbGY8vv+7RUTCYdgKVIGH16sUQblUYI49zyz2bQAF5Yydux+
XYudDE5ozON7eXslRSXskBprLvb5rQxtlAGu3epHf9PPp90/rQU1mlrEjxW9QB0D
9A1SgRtxsAZHNEwc1t6WvrknaK0XOfAgyXIaprh0tLdrhMuutz14pgcGkRH0zGiI
IdRD+neY8iszG5rb3OxYpttpt0aJ2rr3ivyGo8Lgu/+MIJKjG0NBy/rACJRRG9fA
gZ6wCNqIvkqjtR0lRDXJNZ+xcTLQg/9d1NO4sAZCBb+2m4YLTEFSEiPXUihOJyVA
lB9tc0ewrP5NyUJqk2uVR5PzlDmmoSbu1kWhfabWwdcf3+8kONMR2AROkF192qNM
PaYt1n05A2HxJDHzCtU9D4cggl0sO7UweyGwlM/FPmv8mqoH2SULCgBUDIKmPV8/
aJTQvzLK47M4kAjaymOPExe5S7A+yM4yeKkJhQb0VVYl0Fhs90Ra1lxniJ+eKu9c
iGr4+wbFpuqX0fWPvvf4hOVrJKg6RIAQRyeWg3+IKruK6gWkATLCObv514sSrccW
pq/M1XmkOkQHgO4p7vgZuRJItgRaECRdLjYq9soXJ+bTk4xFXOJdhSnReGhxY7b/
uz1rlNCWZHD6UCczM33DxjVXQT8Yfr2ek7ax3Qk3GAqrTS5iMYaH44H0EPaHr9Hx
INE7NQNMl1FZqsFVBH/pwfryuJeEy+FZV2U+F0c7eXDGn2t0Y83v8ry0lA3tVI/j
+/g6ifH5Y+noRXfmA+k5YFyFADpqrUgTLkER+qN98Io0jfoIiAEPuaynlK9OLf2+
++jgGVgHXefJO9gAO8b14RzyDYdOMAhzHv4CMo6+l6irWey+ncA9vtSwePaobGV7
`protect END_PROTECTED
