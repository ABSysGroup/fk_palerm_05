`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mV2+ihdf93MegavjFI8SpW9YPevZ+RzhtlJo3TmS1LQc5WUb2XbEz3t5MvMnYBvs
qEVdolDgVgtzj2REM/TkzKjbAIY/bkL1AhMQNL0iskQyHMVekxqFIIA2Y5LjGE/u
iRlkSwlK1VkAgkaw3hYgw7JH2ps4zrgcyv0YhTxRgzax5uMrH6vauNhLOvuMdvVz
prdwphuWR2w+YT7B2KrcaK9sZrk7Obi8Zfog5HofPXrtNfj6M23nlvsnPrFaaSRF
QUEucpyD35t9Kg62OsJNvwtZWUCYDGPyQ/8sBvrjM/eAe+zVAYcg78+oTSgAhmOf
vbvTlkFUq+Nlo8znqJRmnIBjPhnVzgHTHcqGG+SiB1/zPxuwM4146ibLLt2x98xx
RRx45C2WSUSDKJ0KsKbZNE2Pk7AJsd3DSw6S1yAAVksdFqkZfn0QpefZntkLqlwC
Xdkw71/jjHOVcUkGy5YogPM0lemjNygHndtf3LJacb3U8+eF6bxqftL5gel08aGz
cF3sjU8qV7tL5UDZMPm+bDkKtFLznEhqoSP8GrgmqnNCAXpYXD51Rxp/9/YJP33k
u0bZKfyrvkbIT9k8eptk2dK/IwlK4jaeXh8FdaDP7KcS/7lPK4T6CTZWtosW9HUj
n10ufhbgB4hqIAxK4TbYy372pfWeB2TKNMUnuHFCfXtwRZkfghRCMi++BWmRW+S7
wZxRFOD1YjZyb6dFGE3gyX9VDihMKxMatLbUYxtG/gjE9j2oVswTowHKcJDgLnQH
7nd+rPJSfyjFQZIpLjTgog==
`protect END_PROTECTED
