`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rJfK7lO6dj/XGavC8bgQX2oheeJ+yGLWQu0cE02KTQ377lpkiB76BgIOZ4t6uQPO
IBxrsqll7iTBeOmy7p4jifORlaHbHLV6uSPkL4+TtoaCJiR2nDXappd0fEjuY6ds
NofeYTY8qAhDj+mSvcTdzkdbKt2zGlb6pGYM9Xdo70rk7MdE+9x8s7J22AqXsFtw
tyKS5LeLi++bf87sL2xg1wh5IIPMPSfBs7/4uVU23U02eICAA4+bkDIiS9EGzjWI
xnO+xjgruqg9y41JauxBwBGGB01pCfW1fq36NstC/mtThjkLXDmcAkxrPIpXv1KK
radTeC0BuDPU12QNEni/adjqcNpXhGXN3YFhKoqEYYYi81s0yspVF7wkWX3v3jT+
POWy6SwFYERkd9pelYgCt58ZJUewJ4wsild1yQb6qH7W8fBGvZbPLE+uJQf1BGpy
i3iuqZ1PKvfhz+p6Fn/fUg==
`protect END_PROTECTED
