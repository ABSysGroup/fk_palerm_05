`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n/nqBgn6IZeCLX1x/GtMXObLtTOUWISyuOgdrpJak0ljNwS6kGh6mIZouHkpuM1K
oAgXuoTb8aTDCJGhVddI3krE4lQxgr4nbDyAjR9+ReRbvjFuAGKJOg5o4TZ9aL+r
vnY1V3fK8rTMy8SsGfwOp9gI1wN2YDhGQmNkKh5JYhy9S2k4kRVypOSVHYrYCQ9x
ks7qqoMzK26CDUBUpjYYwq7KN4Wke+rYVNDGHnRvsrg+ekFiee1hZPLWhrVene+1
ZwFD0kC3RbWTW52EJTMSM7vZnCOkXFcJdoZkX8QMQhpUUXo1Ap6YbsBCj1io+oSR
Ybwp/0JTKrthJ+G3T6XPciuAzKxMCGqhlRxH8nPhjkFHEuP7DxQTr2KsgfFdL1lz
POCwRSecZaBHtCrCM0MyhgPl5+dRFoi57HPbJ/6+Mk3OzAmEl1k/lws7/s8Y4WtC
6tGdjYMs21n0EzBOV20m5g/bc2QHIY6Q0T5HG+NV6qexVkQVn8PyB/wdqN8ZZi3U
XN4FDqSL+gQYQ3xrvrWYw0FN96nHr7jvUyanubyICwwm2u7SV+zbJFH6CaFg/8vJ
Vfuy8o6CT0ZHhJe9qJRfyIa/FR6Q95NJhwKMNjxdZUrP8JTezFD1yIiO3pwinv0W
TdWbzphzTexhFQ+aMiRc3S5Z9C2PzqYg95ykSBRB5YIfOrc5QRIO0+C1oJkfrmvC
W7lI7CXAC4a2uTUBUj6yewplTRYRCCKt9CyMldmypaNG0zXNl6YpxIpa8gW6Jb7k
eKbLZ0jPwTcahT9Oy7Mw8wMolgMDG/IPmiF2VFsxr7AbhF7kQuLTVv6wVkQuKzz7
0+I/bxhxqnQLzK6hLXcn+xW9p+8bcLGVaJ0K36o+B9i/UfU9MgGfZnm2Jz2j3RRk
ALB+5hU6cla3DA955OAztM/TYe6poenBfVuRl1sfaHMB9bUZNJjddfz7v4j8UyNZ
I4cJLbpWEYrwEPqGkrDxwJHRyhJwZxPEf3ilBomhcgmSe0tCfxA3Hr0p7puqNNBT
UBt0Zu5ASofc+jPe0JnOHSUJtbHGOVnzTIIEc/j/0W08V5G42Eh1edUGkIWPDo0s
2NSdEpbS+ONdTxOw5/vYii1BelYEP/EQkgh9KTJg0HNFwSpMCJ3KQqGL9xfJfOce
fx36N0vZCpKLtwT9M2sOW8W2GTVk84WfAw5nbx5ysoTHB1OJaeb0kzm1en3waZ7O
SDyMQriRM80R13e28s5O/hqte47i31WpYt5aK5KoLjAvrXXAdcjVUJ97Mbn2moUX
MG6yqGmyCa++hKSovlIrNACGWbs9eImn0XDJPq/8H5V0v6GnT+lDHV4p6Wh+prs1
7OLYCDqz0qQaD+9KMmd+pfuU4wnBihFXZtq1JjzhplWD990ShQk7Ap7xnh1N0hxv
yvYGkoEQXSlGmvyeAdZMGjsyuhRQKm6Mz+MhBrLnLf/9EuyayCMat00gAnlZDHPk
fAqJwXqIhlhsxpjAV3JAP+t4ZfoAmfTkkUtl9AjSWIZs2KufU7fcwjDVYZKzZwpv
0PyOelLCKE8ezKeX1NfIhHsKDsuRDB1SYF0BhBozFhG8sgCKoDiO1j0iHgCBxVpQ
2MxC8i8hm+Gdb5D1EeM0ZTqCLiWXNZiPNo8g3UxMYN92OU9AQeQvOvhPG3gG2/G9
vyWSMOksGbwjef5K3Hn2RlRS7RSpmgNdqEX1eYSDZEAiETRwBCMlEDmSRXORtMmt
mY/skiMLlThu8BAsQvdf+xuHSF2rVt4JPB6GuWOjx/VAniCHs8efTkjujoZBWPsk
fp0fZV/ze3qhQ+MLsxeIf+5LDwMOH2fQaLJQY93bdS5mCa2HZrTYn5UDu6j+i/8l
x/s/HDidwiMiqoG52pnHA/59qQ5mePGw8jKothxa2YSu4soA7vk2SLje5B+OnLS5
nPb9pO5aSpT6Iv4DEvJyKOwf4idR9aiUoOFCesqf89tSnkS3Gy9SpcvadYAZaDKF
i7FFVScM1mHqe7FFLlglGOW6G9KYKrlFHTujU9eYiycQHEwiS7o/RIfOk54ln/N2
T/lvZjGJtfgkgvb89S4E9OWy/kbsTZkjUAY47pXjBacjQW3YH6NhDSehhBCfc2HC
PstUM0coLmL/ZsllsPvYr+731cFs/IF2nhcC/O4B3L9rAG8eiAZOvVTFMRsyUhZU
qj4rohZrTAx24cu9qufDT9VJX0dQvJZL9DMTIQjcS4mWjUxhsIMqAZGnQ/8FiCVv
hGFLBwoeK0L7+ErUuDle4AmbUxxGi8d7PtYdSAQiOtb92Qd4CDhr1QKr6FaRcG0S
azdYt6lSFycZI6GL1Xx1pIfGHm9EFUDU6ImBY8BOJ7j45VAQImLhIY5Jajx8eZ2H
rXgGcTltSygHjlRcRAT6pd4YJYC/jAf4TWbl8zfW9nRBfrzafFnteEhLTXe/tBB6
gt6s268hBRcEniRHMvhlFPGEELaKVvizTEwG7BHyJNML9SN1dwqYVWFeZZbsUU6E
8WkRyf8cjv5juFJ3ycORIPIG8uP9Qigz0dkVIq54l6s9xJ7qTCnalhh6k3Gm9oe6
2OhV+yuSnfmTSmlfElEt87iQPes73X4ZO2ZMPk4X9MUI3I3GNgi6d9FDFAHyzKe7
BYpncnyBsOnnFVpUXZOAfhs+ZXRVECdPZEfRuvR6jpM1j2sHQWUQwNBsFcEZypOD
Yfds+VeheZ4UjrhiINlkp7NroIQMhnt9fXeyhRnnq5eisXKuEH5ZISbzjyLnAns5
cg3gyVfsXg5pgMZoYXye0OJpKKA7jJ5cSRD5Z+Kp7eG+sQjJPNMmfa9LYl1u4FFa
r791GrWcbJfK65O2aj9KbymJN2rrxBXhnJVAd17jR4z+7TaKQfNcVyNB74f4bqhy
ud5HDPHTuyAvrlpYfQgoYBIkDCHlbsBt1wgtSb816rKCQ1g9BwC7ft0+TJGOhtuM
uuekxDfyMOig830MTB1rtmD5RwVebEsFtoF9xN63U0JypUcQEcTG2+spRHZ1CWrV
6mhJL5Pw3uwuyTBVUycrmok+bpO0X/B7fVB8WdiircgReaXtvOKzdaT3wVbJk2Mt
TJy/1NxpkcWEXHCu/2yUwAS6bYAUXptsd011UH8ZUUhWn/F1/182VT/h5SXz45za
9qPQpc7R3Og0sEA+WOlF069FtKIFVGnKMyV/GLm3ZWQA+QgmrrK13nsIDztHISbd
9y7C9rYOkdX3bVT47gspSekgl6dypsEnlmXsF5PeX4qnbbr2WGB7uBep/IMOQXfH
skqlncr1Q4UOD13OkEqrWSNLWxcgWfIS94AU+ujVvatBGmvtBrL3N+49iMWMip86
n2a1HEqAmTHYmAAyGi8CNed2aP4OpvZ+W1hiCI0a4xNnfvaVEs82FuoPvJZ805Xr
JDoJzLcctGpE70QTVUoliYMa+sCsvdCtILCSGmZUHmJFWOGZWTGw11dhldahB2O5
hOKhc3AgYk4dygUQBrhKkRz7VDxhqY4KPznVz05d/KdWHiBiE+N6T9Zy1+QLefjM
AqRfsXJXPeK7CBYDpYIzUVSoptXRTVvkmjN+3JN3PaUnIAxmK46/mkj1+jGWHI+7
TQyAVVEYwttcUURpTi5f1pfNONwSaGxSZsQatJOajcofkQc0s/VfKR+9mqdh/h9+
8eICgehCaMTx2ZW5+37r8OG77cVBm9CYbh5quRF+VA8X8iOdto84xW5hplxXSQVT
czSinV1Jt3Vfv3gkjJ2E36dA1t1kqC7+18PjHjXGYS66j7uNOhjFTg7PpR2s/ZHW
KoFy9zHl2bUQfCPpHTjTCxHTTFLteo4vZROXq/n6z848MAhynjnZWc47fO3EhcLD
KNjZjPaXSTCe0l0AvWnNiNvml7F77lFAtiWUBeQ8sfO22NlT7c3Mw5HoJBY+7wLN
HopqlCu5skvOlmS5Az4AfgemRGQeVVhEo+yxkix3TfEzHZCdoVioIE9d9vf6COnU
SAI+F5EDYCR0jR0Ou7D5v6PpRJYWKn6eOXLB+Xe17oxCaPJe//vULWvvPjcrCyXD
zVVXnbi4a2eLfkxYLmCXGxPD8aG+StSTwfG/1vNc4hyR5GSyhp4AUDQQ6+Vv46O8
ucnXobOqIvEdquvAtgbtM2AScH4zej4h/rh3FH9oQV/OvFBtCmoj3J2PFq2Cyf14
ure5AikxINbND7bnFU+DTpBQlOye2ti40eoKYpCCXbdyZ3uZlgJHu1am8ka1+aS9
ixXUVHMQJQDWgdlo7YkDcjiyf//fpjSr5grNrNmFKXc/c3YaV2FeGrXOAUE3pEnj
kJXxioQ3P3zYiKJpS1DHdEoYLSxxbZe8QX/B+o1Ge/6JYaaGOT77FK6l2sFcObTO
5Lab+CeuGQOMYuhZWjvgkScQWFDBWSzm5H/+gEMNfOwpJTYjIDu+eq45zX3U4wL0
gReW7104Hi0Psq+lq2ObmCjw5yak85lWZHIT7hxoErrGhJjWxsS4tTZxOIln1GPl
KeQh8w/J8ztzBhcfwDsF/NRR/blWG+6LVHa5WMZcFuzHNoZPcEd8eM9ZnOK4jIFy
613S+ORkl+7okkLOTtFQK0KcenOhNpEPhCpMat6n8fkHjIeMwt9kZdk4r1sByJGa
0Cv3NrSYIhdRNYGeC+kDU1qxGxAzNrOpIa1lP41ow8OlEw1L8CqVY6DUlGCKW5NN
`protect END_PROTECTED
