`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AxiwhEcSagQ9zsPLgLZ/oHsvXH5WwkCIhWOCTsGZt8pCW65LeSzr/CeN9JwZ4Bk1
96mpw670XYioMESDWwtM2xfZ0HBXzsXmH1Ug+ljQutIDb8865z9kfXvQGJmU2cTP
qtjq4BmiP0JLDHJaG51ugUjanBlyiVgXZkMgJM0klD5UGvCeu1L8ybdj1aifvqa0
Mqko9HSmPrLh1AuYtmg1bzmyXttVyaS8xQa/H6M/+FN8L6WV1Lz2sf9uJFD2mg81
UsnMoqYNFpRXPsK5Hx6dLqQL2X7Mdv/A7124tfj861aBPiqUW8hQimIRPOShOOAW
3TIqCBSIRvMtXI/8jrvJE7LMfx6DPU2SVY8sXJVjg7WfD1RVY9c5qfCqfhh58xL4
ZTeIySrVKdKniHzw7gBOAP+IuxnIsUxy/cdHN4wJnmEKP77lP5f45oMnuFe/ohSd
MPBk1BDKQYXGDczEpZbsftabpP2p03fC0aCaEO/N/boOFehpo0HYFTfpC/u/6HIA
TNZaGMW2txfkw7kNoC4CHefBRpcJAZC+mzzVokwJ2c6YHGX9Q0oR7V4V7uNEoMdV
`protect END_PROTECTED
