`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wyijTU7/69bYLdWMoWliKFnBHkAP2ZaHrctSBQugxnR4tw0T9FgvMI+741QoIsdu
9rMCsUF417EHjYuofplXs3oxAWcBy2qIRcN0fUVlA95k5mM6KMsbdq41MmMnc36a
hR4UHgbelIXpCE8OE7lOv1mzAGBqFiiCkf2uS+Yb/yXmQsYR+DaKhY4I/A1VWKEI
fI0eFIUSauf+3xY694K+iBo6Jjv4AvQDXMhxijSQJTLU9aVLeQFW4cxmPeewW9Mv
nSYvS4eKYiWQd4zlejx+T6LrWygWvGry5b0BpVmg24UDGIs6W2iCW4+/gyfmY7dE
saN+x54GCRtSOzMu5rKIFDTRgmCFQp9/cCa1+0MlkTQJr4WACG6YDigkwccE1Xs0
Us/4tmjAkkmCl1Zey65Ocx2yOhuychFKviIBy9BCE3RJs2LIfIIUogrFAS7jiENx
QJwa3LXDcE9kbGOCaIn16/MuCW9YHdPEiMRiHYN6aP1nW/OikzU03ZcZUwjWo0JR
1dwbfGOAfYckK/0d2hK3qW/0tnKIkOEecDxUucvHHqGpGP7I5vU3p8+28MzifOsx
qkv/sZfVUO7d501oPoz5xdv7GrY3Jgy2w8pfxzPRrLRZEYyV07l7WZw/otSQEzEn
jRec/BfLGjhXhSyrmP6Bc/XGjNcdfd5x2cLyrkN2z9tFkjbc1ci4skyDQ9OtHDH7
aIr2ogItklQEXTZKeCrgNgUcqky35v6s0M4ytse+JMfCb0GMLejuMfHeAxzk7HTp
BZARHrTg4WSLeBoKRNI0kTdLnNA7nE3d80OmbrUrjTf7Vh9F4iAMQStuUfwkHImJ
e8g3L4jvgrERXtFwb4S+avi2JSh8JIis0fqSwKuxbEApbPK1vNkjvyr+y5caOvIZ
Vjk1E8+rwTzwpTBs8SSv9B+mRXPRnT9Ns7ZYy6hj6rbTg7OBZ/zV2V8nV6IVs00v
`protect END_PROTECTED
