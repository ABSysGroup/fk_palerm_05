`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o1FaxBTNRD93APE5p3HaFhBEiikiwSqrUuYanRH10OVKvWUl/W05SoxSNz2qL3KY
MXL5iI7E5zXIzvPKqW88dtWUQGn9JfbqDBJ8e0ryrEO8kOC/UY+hdiUxwWWRlCng
0TNteLoHdLP/S4hJAgS3L8dtDALi1sxyz7xkAxVfWscNRVGprlII5cIlkMFJF12J
84vIEUQnc88jQjtrnrvKBqNM5pjvH1KNKrp+awXPA5XuMtJ6PumH39mbx5XS2NyQ
2nj0xhf9taFwxsok/5ZCaK5udvBO111+Ukj2yxwq7r2TadWuedB+oasouuXBJwwQ
mrA6t2Qxw0JrkErl+wJeTW+wj92KNVr6FJbWW19nDN8wknvrEoAVQEw9JSOQVr/6
boA7sAPNztNVfi+koXdy+wO2Tvdvvtz/BurH1POxjqSXmn7ELIkO6aDZwW59HbDf
gxMcSMkNTFSMXaSJwne6ro/O9ro6/AKOQYRUmWkPmv0y6Q7+G0dxoTKu9zPvV9RQ
xSeK8X63/Sj0LJKNvbN8IIz4KurgFCyBJeoTMry/AsLnR9X1wUouZkmmkzs+fo0N
PJJa8kvp8FcXMrx96SZ7hV1ox9BpwxE1Rwww7ksp+LRYxjtqMzYMleAKlReTrBoZ
sOs1v5ZJHxEh3G8730JXrpfP7p1M3w925wnqaCZvq1aiRDiizDfdzO+U3whi2+c7
L0MoLtTovhoSas1+uDXXnmrdKSBX3gRZuVz8tBpE5ZQZiuaEHUWU1zi4ZrVqoPPp
uSTUmA0xbwZrHJBTuVvj0ULO7ycZQRfevmOD79fr+OvferV0lgqD8/UPeJRJPzuF
Kcres2t/dxopfuhIv+FsMCtJwSiztHrjiLBiCaYUcKT3aIP+J2a2W46JTEJ3CKm9
pcAP8K+rtl3ueLTjUECSTHMZ55FzLL2zFefwPxdjgfHqkUnTfNpnb0Ljrwae+SzX
0RmDWS85/6DbANE8fvloTHP9wNVcAUtsy5bye9H54zc/zeGwYyQePcn7nFyMOUJi
dyaMnLOsx0o/49otDg1Z7rlEwByLwYqvlTn65+YUiIULhcAJ33xQVR3a77hSy9w3
Zl76/EY3cf6B5qY0fIq3Aw5EK6IL450bTaTLplychHbFUMbsMLZrs/xVSmSLOeQk
0YL48P1u/vQtJ37YdSN9IG0x43i55AiRpDG1aJuN05u9o6Ro4wRpNsNt+FRmedK6
BSl6K4soO1nqIjuRwpXug+LhSubgoWb4qr1N+Na7l1z2Hfnnaow1gSWkUhgnPOFz
DmoeGAKAo0GqfnBXV+hOCAjlN5m14fk80oyOyxvLOYMh/ytUkkCsy1YY/xkxVReB
lDPZpMD0BMq2vShOQK9Ea6rG/VtvxGQG9J9qFEm6Hfex6RAfsTCplb1MpntdHt2A
QLKxuWpe0Sr/6CeYmxr/4nRDPYsm3L3z313hyyyOikbx46FTJ99MTByEbWG1lEHR
pj7i2JfEpbraVWHsY5sm8eq7U1bgsSwQ67nHSeZ5rTn7l01VJzg2OsKKReTIzMGW
5nGZ1KPlbOFAD9VZ8APPs26r5igTnco88ZICfIwUHmTm+kfrlrqcamRBk9P24BvC
d3QsM09ixDhHzRC0Ely/dUSkUgwO7bT3r1Hp46EY4a9hQHw7tpAviOiARcdc1Dki
yhqyrR2A1l6J+1tldlUO8TLUUoEx/SHpgsGnVGRpE7ZEe6Lz/NacErRl+NfJK0JB
8A2sIy9pjvSi84e4oESmZuMrmpyMaJKvF9LdfNHCtpoKFgKQ0H5GCAIM9mnanXAi
lZPg7D7RP45ifG5BsWW9psN3oSvgysGsNe2VX00QSdtPozobV6mlbzKIjN7iqIXu
mql48CZ8hPTdjdueMTic2h2jsZyC4uoz3QxhCmKhT2N0PKEvQ5FoB0vJtQuZUVt0
WwtZA/VU/NQ7XJaKXbU3wlvbLqdSePF60XYlQNaTFAgliTSFPUlua4j5yy3VdoQB
7lt0aQUgvRkZG6LHci9UHsdEn28o/qiYKLkYsFhrLPSw22LmiS85b6l3QtofeAZa
ml+0lvcm0+o1QhRDz3XDje2aVNzv6TJY5h/4CiYtoN5IYN5H8+Wn5RK+8Cf/PqpT
uOpq630S+TWzDi1BX+TWAHScY7FWc70ZFA7RUzKeZGgY2+FSfCe7w5Qq4Br+CBLO
G5XtfN0LK3dMIFPFNAI1+j/v0DoF/FdTh7IYbYZy+hXwtCJL9qnmTIFpPpK3qB85
q1/yDJSAgt6uaZNtlzKEU3rTjdGSabzm9QohveqmWQ7GoKPRdO6Pmf/2lDF3gYzg
OuRbUFSMB/71xlkTHBK2bErhH1mJmUmOueABWAP/OiGlnDFK/nkYQrSmmygrPfug
6Gq3C7MN3zZhl5ThyzyF1Rzs0+qdSiGgj3HRVg2IsOJJyJOmT+JNgXk0cYuPKJNY
uiGAVQUxFb9ug5wHjqNV6vU9neyyw+8SU868Nu6uNRowgBZuUtAMoVBNtubEqpsf
b2IGnQlBEK0zag0QsK83k/t7ie8v5AvT+V4PuBML0liygvKd6gReVOa2Ur4ewG9x
MfUqU+azFjafGDeieOdorT9QZGxrPb1DjAwXjFtYfxaPU/jW5h+k/n0ny4kpAEva
s6AF+7VgfStyV79vaqWULT6c4v+JhIWGmE0FqRWiwN2FCCLovEDLhlC/zSDP67v+
lM7lSSEfznuGepHoc+6dCT4nyznvZOh/bRVDyPNNEjaSbxoHpWjNEMTTWuRyYbDv
msKUefVK9o5cnJB+OG5ND2kUfBBH+862fDwsLUUASwg3KSNY9gHvH4Nj07vzgb56
VwdUQZN13lDY4Y9l74uISoniy18JsEYFeC6UJAoQ58zprjzSx6S76bJflG4co357
NhfXgGsPtHdhIl1v5nO4Q5JjtsQBA51kFkYgHxbnoKDasK2SqJUa6Ya+ZaieDqLb
+1t71MQBkVT/cFsP8govowocFHbPNiGSs7RnX9fBpi0=
`protect END_PROTECTED
