`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mBxYMtcr8Rlfs6nkHoMsDGofC+mziIilUR8LPnQGzskGLUw4H4ryS0F/SA00lM5j
PfQCXU/50aR96j7uvD4RtwNPmk85ZLs8ng2ZCMuOLRVjaxIs17Z1Tkhx4rqrP5Sq
13GdG7ACZOcZIo0HAzj4n+3d8o+rlzFkPhry9z/4DsnuR9J63L4xpWZeNSP8/IRf
IF9IabqxHA7g33f2yQauLdaZPWoJVB81IqYavPzQ/B8l/AlVat7DLIowjFZfe9hO
OXRrQ6GFvkppSnbT5kU4P+zNYlIokTbgNgVMH6eq9CTBkoYfLpxQZgv5ajJQKYZL
qJHVDIVmPnAcCnRG230RH9upiRmalzmf3lm6LWM9ZI81Wtb4KsgojEs/o51nJVUK
qp1cUJCKc0XF8eFsgrMNtQ==
`protect END_PROTECTED
