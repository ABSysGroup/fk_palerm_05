`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3J896ZIEsSGwD9iJasNLy+8OLZFvaFJYXwmBAc+RGy20jK96apKxFY6NCuXrJ3PT
z+aDVXIdZA7fBecWCnnLrlL30G3wGhW5NQ/Tyfsj+oBNzyVFVIKsLDmVlqwy7I2t
+qyu0TziiL1ZOPBdAvDUnnEyIZz2TcihG8WmFan+/QKH7NfBcNKhxiFaUGAPIxIM
IRptEC22QayvY1kH9oLH4l/MMRL6dDXfdc9wShyNg7Qu5Kf5TMgyZqAzqKPcoz1K
RrGIAdrZ95TDA6wkSGR5AQp9EPtGc9M6gsvzdZnU6EsxwRwa6Qip6rAJofYCtf6I
kd0cKO2SaDrY2Tta7K40WuMuEeMwf6Kw0xE19iQfZAHlByPKXrFwF5xOpHVkfjs5
D+oMKr6reYoeLEPzSO6obitc1m/kPjhnpSPjSg9SOQARH72WsoEamDSZ2IbLIHYE
wHcMcT8VpXfSE9JuVonpSdIJ8pfQ0AZkyNyGQvYJqzOF58JpRSnj9ftx7OpVCyQz
QvmkG8ncly3R9fvw6CThhskTbIM0Fj1JhMqFXxztdCuWgWNHEmh0a8WNbPbxJ+pC
0phdpUWhvMGLktSlSwadI6xxF9GERqbT+E7kaQuxOooqHAgUHF+3ZCiTtjPakRnr
Giep6I8/duYMbQ+h3bShji+D6zQnI2kihOgEyVDAmn/cw7cxFY8eoaeHFUMeV1IU
GbEW5pfcKApBcrYr1+bhcpR2V4kyIGEsHJ5rPImurd3LGb4Gy2QS7NOr6ucGv/bQ
WCRy0OZwfzjVGHFk/PW9D8mIqSFY+dVKRIymZ60rjKIJnZSeuUynC8FaI7860x4j
ZLaxKPKmeOaP1cuP+O6GI+lMZnv66HPqoFuGidz4Erg=
`protect END_PROTECTED
