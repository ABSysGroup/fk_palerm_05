`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xbpnp5tXS9LuIW7KYJLiUUVikJt9y7l+tpPnAiAiA+tQaeqzM05N8Kh0TXYE0Xvu
5CdVPkMTrfoSxMBN1v9OObOCWyNymWxHAsxJounQB3Z9/KezuB4N7iyqFGOBlPHM
s9upPiZe9rDV4Gvvh447ZuKoNYzVGxa3oHKN+dPCBNAOySFc0/kdljdHuQz8qr1e
B0snpMqlwdOaDSFfhx4+79JyvpdIHuAfls0MugbQ6ePdvS1xmVfWOrQWsn70zVtD
OiiciX3nlIGEmf5R8bIcgjNtGP4vjN4ElEIIRd9MlWgbI+MHcEHtKZECGgAOcuoA
mLoT7Qwwl1oGVdIrDdDlTg==
`protect END_PROTECTED
