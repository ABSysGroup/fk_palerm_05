`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
00So5ypvSpzwWrbDy9C7dNXuRPcAGKazEdvCVoyh2CxZlNJi2QmzGKr2wHT8DvvY
gH2COky9cLMj9KD3uKI0oIQXdria3kF3dnQ0INWbF7kdYbD/iUSLM25D1hYR5jDM
faRqTR6O5/PhiN+adcLod0sy2vei3HMjW5fE0ywxguT7mXYybPut6ljSU9A0XtR8
0ZWqUrX2ue3DvjP1gkhzW7gxd4+5GhNrbUQCZqjkqqOLT7maoq48iW2JKUo9Idvq
tAlzdlO5mLsrkzHcsAD9mEdTrXcSNYdEWxvr9+w2m4hVsFahGG0zIzFDVVx2Fpjy
6PO/vnR1399kS+wms2wDPGWVIkcu51vxJ17FN1+QlGeqaB7YV6+nv4vxdpbKk+oa
MogSR1TUlFQ1/gclV323UUSEic23UoOk4i4WZhet21xTJjNUYrURL9+AQyMbkIpf
Bx7N8+MiORIqhBfAeW/lkZ1WCa8WqRK/prmHXWHUeB4kweaoIHpYbDaWLRKwUZJb
Uua2mNqLJk8fZdwpk+5e13kWNLzHx/Os59LgOyujWxJcP1wNAE5b4lCXg8vdoIDL
TxFRuKRrRINsHG8hKML8sinWBFxcgfeMoMPxfROUqsV8bR0K34ChPINCcf2Dn9CA
j50hUqNh3WIJRcK5zlsXFyDebD/efTqdqkpulfzHVtY=
`protect END_PROTECTED
