`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OoIyacjzS5HufJeEz8b6zgh5/br7qfEjPKw4nF6d7axoN8Qq/fqBM93Y/gLpjXSp
j45S5VipzP/mopk2WyuPbrHaoT3Y6KBnOxf2ndHmoiAner22GvrtcWs5N37klcuK
/j/k4p2o1aCBtS3A7KBWsNYGe7D799khCvgpCiD/uf3tV7hQkdgtFG+dMnkpqO1z
c5J/A9Lfo3/VKm9NSmn6jAWE9IcSpVgZpja+kicp6uCsfGOPNolprtWTUtNjXWfx
/sZXtr/3DJyrJYTujGiCmN1NbwZ3gRTCRrsFFYtihUpIpuBiYybAgdV8pn+76Ml0
27VpeGgQdFUT5Lxj6rrJKbPmSXZdRO0VN/4ap8VQ9UKLEuQllE3aWUWFLC7UsqvH
RwTv0i44tMXj+U176IegBA==
`protect END_PROTECTED
