`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uCH8dTTHsnD9hSJur1O8BWdLsJK8Wv+/jyvehuTwSEL0Yb20fKx2q0tMkIqGy+sB
RrLil1yzMYhcVhpOPeqRd7CiTibqzHDp9ABLtdx6o9flCIVB+kZyYt998le3B3Ux
MswY+FXJnip5ClYa9aXdedzvbJfWJkRVwFsiNGKC3gmHT58zRN4QizOrp6NSamZZ
cTrMi5pyaSbNVhafp88e0MMsCxVDg4I2OrNoKk+qcxWYiW0B65jcM3cD2SraxKQm
zX6lcmVoItCV7mv2RD8waKe1tG7/gbe+7TKcW5jYvOImoM1Bzg1STpeHM3Osh+aq
oWh7Ck3l8O9XjbttWdzDL8Qb9PL2cVIJp/qHVMtn45OvJMOIYwDCpTFFfc6EBhnp
o7wUX01ggvsp4TGOg+PQLwB8Cn+YbXWA0/np+MeNW1JI3H9ptRNxHwsnhuhCZVnQ
cdA59v4bgAc6ErzX8x/4NnFYqF1POqno+LzJwnVekr6/o4VJ+1HChSD75JjEg+f9
ZaT0O1E6TcQP1U6YJWMsOh53xhytMfYfPzmYY7hORu/hQEgLVvvkc9xX1algy6Bp
o4m+YPowNBuXn2FK2SEREIfIF1ZO+ncBe/CyAaHEZbtEaZHK4aXCCakhV4aQLAAf
N++niU6CDmyT74idapOUxNs3fabCVZlsGDPuWP/mVzjUKaNgWY63zP5jSXMurN77
FZ5RjMCaQ/Zx32Nyuny278iFbEs6gD6pJGQLZfn+39Nblb22yjCVAERLb5ApcOTw
9NDsYiJxiYM3CxQ0zVAnYmh95fWjzhULW/PIzInXsv5vr8M3SuE5TXuZu6UDG7Co
yJ9Bs7MvjyQvSdSLpUvYhYeyFYzPpV5sAKI5iBBZhbpJ0EJ0uoX6IgpLZtxr1KJs
QKboRJTmScaFCstqilR2noqMDBxjjc6+AplezaHDZv3l287LxYhiXyWmVt+l1q4N
4JhA4x2smj5BJLXFnEVdrjda5ywXqgxG8r1Les6fxRwaqpvuWuR2lJuUXVoxbhly
P6rNzaLeHmNJFNb4n3mbK2W7MgC1CI0BjqRCZ1I42UzsNQJ/v0f7P0mIu0b5IWmJ
cTCuKoWvYOXezrW/OXC/pbtFe1tR/YPWVqbV59eCPOoDxbBQsxOhlr+4vnF9tbcz
Z52ugy1tSzfJbVo1HotUiewOutIDp85KTXhv8DQzzgx2Sl7fOYFKEOJNlJBZAK/e
`protect END_PROTECTED
