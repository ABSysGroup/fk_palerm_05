`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bQMd2w3drZmqdiZtPQYlhGemJzSH8vve83KgshlUaiSI0j3voRwlu2KFlDOECAXa
W9q5mW58m/WHTRbI0xFEF0XXO5lN06SGeobWJ9k4h0ty9WuYEBrwBV6e1dQ9o+CW
8qfT9N1y/SPTM0Vpj5TTBppnDk1NJDf/+W4omTFjjPubak15R2ja5e+nbYvpNgGw
Ulaai1X/uIeNCDWDNVt2dnol2dU3r0V47Ql1M5pxGNWAJQ2XSeY77bPfCCyBmBfA
TmLn/TGvOeRc6sBuoxt3B7FxIte/5HGsYNOuODn74ticj9D9qNukbAjLxkCdRd0I
B63qH7uD6TKPst26U6tjHpUFrcVDG6/CE2qtXnixlWJqUFp/zo85nTOerTd+UwRb
KSHCu0OchjQm4hPHWefpf7Vzmgy16YY/jiV/KUD6yNe4f16FiwrptgxNyrXx06V0
IrYAOVSSZEBWRRhX3YOfb0SIQpVwN2/aT5hbmgbMjaCiz4sZIjVWLlT9nnsO0M0N
HQ3FObqooi3STgJJpl/Vb5qq2jNA55581ijAckstZdmV2zyjkJxFZPbm0PTVdtLB
KAOo2e2dNB07XGg/TRVac952z8i5IdkxrCMBFikkBNcpA3NY/TsU7JkAxeefzlmL
tVZBxQl61w6gzeUDv0iPAJ60iDsTqQ5uzaAOUwI3ZkbIBeKwe/5FgBQMhny8FGXN
SZbGQ2SKfuO8V0YKIdcQ9ck3fokjXBb4CL2e7/hySucZXljT2ldQONekT6HhTXva
e7hofv1OEfqkHDE6bsVrCYKGBA4OLKLP636X69RK1yqdWDHdw0hGk5eozeUXQsf+
zXgAAnuD4KOw7W/PiJZtauEKvskgGSAUZAaNTUMbwDOgolL3Mf0lNqdSoX9oBvp0
vpOvNpLm4cX07llrbLnwcZClyS8dReMF+Jz+nbtmjIh5jzKDbUlNIINovoySYhQ3
ebjTCZpA1/Ddv4Wapb/YmG+5rE900PBfmr8J4c+jB5tqZxHkB2cqAR0XVm523ySb
HisCJwl/fxaZcOVGCJ83/D9uO6TYvLzEkm/wC+NX/sUo5Tvj+EYs0YGccHGN5XAR
lhFbWUIThyy0vtYZlbCzrd37bMlt4asC8YPulWa9IsCsQqSt33murtE/mR2wC4RP
e8Szs8idRgR1qJLv7SS3FvBuxhZNOO27YPcq3wiE9baDUDWwYTQiQNW4shj4rlBw
11lSuFgRM4Q57GIxrVFIklOwpWl2TSVbegeJDxbRmfXluzKTKiUbbTDwb63A5/hv
tAv9qHEGrpUiWMJHNvebXiENCp4dJJKm2ElMQQgR8u7yp/Otkd3HDA5YrsLlMtv5
+VVVHpN3iwlWwJCg/bgiJzWuMQiu+Cn4LW06GCuNRclnZTAPCOrSQQgrAX5/gLs3
FMeLmFwozBMRDRIeFs1peYP38oYXsRTUMb2j+qnseFXneJTYifVI1fCQHQvgbYlz
ZcLT3p1hkaGbjwSDwTfLfdJHc98y9/aAVNu/6SCrzClhlSTMcPxxqAT1R8D5K0qy
qzkzBVoP1bl56U2cEV9LFGyQPPtqN4ybJYGOS3M+mUeTTS1tbUdH8W2YxJ4KD2uO
LSe8tj88HYbxARrYBn4z7mEjmB93CdPYSNJvdqGb3eDZ0wY8jMIe94qecLQuboal
SPz73hfFWH+6qq9nBa0slRovMtobhd22EP+eKD+YosmkvfFwor5AVPdH3f1vLKOm
US5S3avfTTIBb9h8dPWpZIZ06ORs9ABSpCjrNAU85ZI2dQJFZhE+POLHhMP3wM2+
8HjsfXWWy0APfs0a0iJjYk87cV3hN4TNL91PtQccD8bu+aT31nIVYtXCwZKJyXH6
9LLj9JW7qNQYkD+eipOMTGWHlT1g+MulYa/9+OsV9pl4rgNV/4mtRKiDLz+b9DqF
DPqMoLnXXoMfbdjNf/LzcmigziRC9Wqt1NxEncGs95pqrFgP2nEs8+qVl7w8LA/V
4HaxpY8h8lfowUaM3NNbcPOInpMUHWc3ongXH5wmhukGlFe8ywbBz+BJZ634m1cb
vPG/V6epyIuMn8plnGOOhvE+jLlWqtufZ2UhB8/TQXf5DXb+miIZKOD+R7edDTeq
yY68luAh18NZ2YD67ptWBuuaPXP8wJRaZ1uZeHR9IK5t8W/WNHuJ6WyxNRJ7DS1/
Z4I5aIhdWRP8QqYF8aZ4YwgM0kMdsz14GSFq4wx98f1hFOBXsZm7XgA5Vv3Pe58b
pNddiGJeCpeSSCYH4G26KaL9i0BlSgmRn9P7xpvBCzO7+i2NzSufDq5hdyJJjuoS
ykVLGk5rWMKihA7wXwKa121stx8w6LwjQH6Ag5+im3k90NKCkld7oM7epSfcfQcy
J+UYnce8kpXHp0bwKMv2NbmFD3ohtvW5tBmrx1uym8vJFsnAMg4LP0rPAec5MG2U
6/2wsIJx/G2NDkwpbKXWJE98NcMHkt60Ne9mkfmCeNuUCKU5D1C0hTsTjHxo/U0S
nwyeOL9SVPQ3C06Jc9Fc9iy3UjxUOzuBMisy2s6ppVeKNgU7RYPPy7TFkTvoRWsx
GQIPvZl3pJ4DWD29BPMFpCsumJH9GtM/GxE+VD8HC2z+3N5KN0DBgPV8KOStJ8dw
fk7KKW+vuIWw997ux3uTN4KghY9/3yWR2Iffktzu79I9AayCP5hLOwi5UIWr/Ah/
FGboUAn94qwWSPlUI3NnQcG5iYVMyHcKKlv7BNXVgaVPU29aPDbcggSkYjnwUDPe
Y7WqbIfJ9Cpv7o7/EVA6iUHVnBmJRCyv5WPbiOtlTQmqdtfMJ74xVjWJ11I0jkkA
UyVzbgCzdWOFQSU0fRgU4Lq57vs1JR17f1FYIUrfPGPoeU71JfXzTH9QbWmKr+O2
Zx4FBdxUObezNbXRMCLUbV7GcpgR6sNQjSVs2AwjKBBbvCpBGdwITlf0DCRVozGc
polY7lx6OV4FmOIOKosLdjogq8o08/G3QfnqDYYk/w/BPda66G9YZQ+u3k7tAkh4
sSMkCoQNZw4L6uODAVnVIWUyCqTBW/azJjPRDcz5CriPeh28iE6Wu0luXVzbbKZK
g28VolV0MqV8w8l3LAkrkCCxbfZgEWvSvkuODERioKo3G6V2rsCkUhGeod1hKmZE
g8ppGjnt+xuK+oOB64juMOQVrneEyFx2Z7vka8PMutitZu5926jgkdkJqpcA3UIE
Co7+CNPdtD8G+E+pAHfQeMsNTfcjSZrzf5PL4iIe5ACjk8HHbnjgM1GmH5Li+dQ0
EcxB3SYLYDRb0AAuZSIboEvfMd4x4v8tM26oucW8zCmuE7GnS7J2vJpIc59GzfNy
X9Xwv5XRGHnfdEybE5ddEahi18F8UDlt05XHpIJDEgAHk99Qs5IJHXOOgibuWsEp
VJxaV15f004ZBMU9KK7FQqLB3OHm7N8VUL8m8GWaCp5DcJMdbpwoXHnqJeiqPQUM
Gbc44N5SUZjy0O3BfPJkViM+Jd5LA9AdJwK/TTR19d/Vg4l9Lkqsr6meQHqE1l1f
jSw3Qnup5EDZe4D6tyPDAXqLKEsJxSMTzErQxmfYZgJC85mk5Wpb3mbmXBY/lPI0
znczI+au+kTR8jT37skTkUoyxvb76h6gryZ+P22Vc/zW7ntUhu/Zq616D6UP980c
1plqDzAM8czmDxpN+1HAFUBO3gf8NYrauPNAnMcsOHihLL1zV79PjAL519E2j8k/
Irhsw7VOwdFha2L7CviZZRAygfYWWKP+xi5Gz6ERRwsQuYkKA7HMyBN3pATKMixp
F2nrgU0oVYrPmmYSoQqp54HLAUaznvIUyCsfsnmTW6xgouTpURV+O3zF2SReccuz
sEU3uyNDjBJ7n8aGNw7GJvdnf9FnAdP12AR0ptMq5/LMhgiWInDowoY31IPFLC8y
CF9yR+8CDTjjPZWDOAoXKYOzXUQ7vDz32HgUe2pFNR1rU28uv9VqiHOQfSr58roq
PJY+F+GkZuGoA27UC/tjuZMXzqGbr8hmBETasXCEvH5rUoC+lwNFEx7PeT24m+Ez
IvS01g6VtmkwQ8TKt3TqAXyvbIUAK+K8Z5HCtJr24dFshZoS1uHLunuFNyZ5i8E1
3tWGn6aIuwKAVTd7e7s5xwWboX5mYNyqnPdNxARYZ7eKO0GFZ+XMTFotjMn/sQlK
o577dXaGSY30qUS3FII7Bnd2RpUPZTRYgSBkctsO8L0RCH4H0UCPSpDMCVvFJsT3
M9mkepS32L0J8rtYLG1iOxce/pGIcc/zQ0ENdCDbzB9R1GYJG3DWXipvJVWQSt7Q
D9LWKgwcFy3MG53+7o3qeuI9kE40wf0xGHhnIZ9vX50/5zAW3PqnsYln0FR4OiG9
tDg3q+74H7Nga0ybLvwi5HWZpK8viGDNmLuTbqaXlf53FnDg5VvpLhrV0iC/49VD
48uTJq8tfJ1DUwpErYEez3u0bijFyufVG+bIvFzgcIQnBfFeDAmWchYN7o4joex7
3NMwT8qoYCDmbxBcrezuQw9bwKjjxmJrMWyYsbuODUSDsejDg0Ek1DFK66Jw9g3Y
k6ru33kYzsD6XQIbeUA7RJN37Bn43cbmjiOHIl6Oj//iAy16F7NTPEuO277bwogv
SfZRIUrIck7lAwUEdHka5DdxKOQKzjJrLUQNa4zAu6Lm1laFS+w/qzS0P9FMcOvM
C5ItrzgPwTcw4hflw9vsWvt4LtpZcRa+HH+dhi3Zsirz8ZPXC8Pc2H1G6GXdzuKu
Qp2SxQS4MbOdzpUCnv2luD8NJeqQlZW9oqysTSoQ586WLcxWqSXVbqhcYmM1nuHn
7NXdn10R99VoYGZN09wgHb5G+ipCIlnug7GeoNBXmPuvBRtpQri1Ud+fn1aZo9wu
z5KgA0NAhGvQgt4u2nk/PIOj2CGDogb+TcP/n07l+c7cgi7JEFTmOe5HW4LTqy41
AVAkV6CD0o6aFrd7R7IkBMRRIOffTJGAAtyadohyX2ESOZcTarEUBEkt12kNAAlc
RurDwNmos1xI0xEkVOy3KWgrdyKKtF9pHx44x5TSk1tp3egcV0WvC6Cve498dsv9
uz6OLrCl0tGjDzdAadpO8cEYaAYhIQmJW99p4i4R8qvHEvz408Af7mOgLfehpU+S
660Au+icSvpehKaclMw98zUHs8q0H/yD4WBzh4Mt9ddVIGMpR5/65uJ+d0ybJeG4
tXW9qfFAVnUznobfxcOenKAFbNBF/rRRXYqnx3/ZqE8NiHN/ByPvVutJElaJpvJb
CXRopcSuUMXWRFaQWFF9mOTpFWFgqzOhrZ4bf9Bc8SU1ITa41Yi5glIHke8cHJsi
sOgDwOINzHHyPLZ8w3kpPX+hoqwO8ZIJtF8bkeRw8hHSdVwlCgouXG+y1n5QbCDN
t3yhjxHDi+QZNYx3YzOxhTZshqYVgmQm1KljGgSbsKOTCdkbmSlslKGhIx3d+61r
B9mzs6H6N6N5XYa/Xnd9lxtUYeop5z6cvvz1MCN8DeCdkHoqMf3wTYeVjc7bx/9W
U3AQ2HjFAUe4jhQshGkit0+WEcE+3nfOi1I7SYfGMxSpWR4arUyxImiY8lBd0vu8
rl/9k+Zz7rXGcuC5tWwaKIAtWTgeQ3xkTfqvv7TZ5rZxGmVwx05sq0C8/2POM3Ur
2rjQnn3zF6q1LcervG9Tf1QYqN7LtXnoGD3N7jqclljHxoMtjpbNgIJ0Q9IJzksm
/PZTvF8KYOwy5g9Bs/XN95TpTEEDvcHpVaROVconKsk57oc8ck+YZk7pqguGxfKS
A0A04LD0d1ZKra1yX5pOE1r8Ou6ZfT3MjdrFF8k3rTyG8t/CsZ8R7YadlHllDOgQ
xael0I8bsm0ijZxPelCeVrZNCWSLveklK8u+zm0heYZLDDGz7sn4icXnmwJF2Z4l
E7CYIPgDqNfcY/xDVAGwy4nKB15HN3PR8mcwp/1cpFDkKDxOeNO5VjQcdAqytjUo
v9giHcBICLWu6tS6x2PtzDIwsune3IaRwtluk63GfQXyaxFUkQ7iR1HbO19kQJ1r
sC6r3tPRsrhnFXnAjsKJi+MU7BJWDlSXYWOTI/aKCwWfZdJdshFnd9i3doIBbOrI
vYyFTJnx3M0fyrdV08WHXVVrNZ64Tox71Hr1vE5S6vzttz75oSo0MQnDO1GihpK+
CljgHRVB3D8fxZPXSbTz5kCNz/q/Zh9AMBZD8V1Wq5OL/M1nHDsPSxxaGt7WVm40
FOc6zdto6wEnx6Ti+SSFb+EdSfgUfkWBmpeIn6SnE8KJvxfwbpK2Cpf//CEWXZ2Y
7LZYjqnWx45NJbFYUMiFim+WDsu4ag3Z+JVIJ1WBTY364nPKaiTv2Zn1NcOeOiEB
0Kg0UsEGxYLTlePFgvpLWrowTilT2pW51PTN7q/tILbOU5HIlwIWvf/pwOsBXo1F
Z82WEwUKdW9TEtE6Te+WTSp9DUotMJJgFgadRqgoavJ4Os2RfZ8clXm0eGb344Yf
Vdlk87pXCs78IKCDsiDXKW2UVCPlEqJ2pXGi2rzP2Et5LQvgNp75XLA+2zTfWhTs
K7hzp8k6Nygpl2aAac/N9hlvX8g/1Q6lfEHS1W5CoDdd/AEtE/vQuWJAvydRRGXs
nfDNXLPj0ejM10ixBW5jE3b3M/bGVVh/SRffV5uB/KsAv8GHwW9+99azqxAbh1uv
4aDle24OqNNVIo4bWXIrM4QU5/+bECk25UqmEZfikyLavp+Ifte0Cjb4LuTCFJxa
8K28j46q6VAbkfR4G272vcMUjO9PsVxsUgSMjUgL1sNMi0RcxZHg7KoUlXJaWHWI
Gd449L6ejJwb25cjhEnwBjVjOm8IILZ/i45X5D8VMoVbDmxLW+S+MOa0vXK5kbJJ
5UCPWojKkbDSAGcpuFRVAeuB7kO+frh3R7TNstxktt2qMEeF8lr3SVAN3mdNf5uq
rOEhiL9pyE1NvKmUs1FkPdeR2jiVbEgj9TOszbcoOurjqICIGCAjAeltrhnoqg+Y
86JMCO675LnbiR/Rc/aWF7J7q9QHnHHVwyM6suP5VQ+1VZn1oXGIhQPExA1b8Kqg
ABdTkyMDElM/PvfzG76RQjby0Pa1UWMRLsMovAZDxC2TV03+QJUG11KW1eFccr97
hD2dkd3dc0UI7Dr0iEcok0dKvJbbKTiN/OCJoII9pI4Lz0Klc9cBVvr59Jnh736o
/M8xLZH5nCYmYD2QLcWKiH1s01M73zy/rja7lfegR8d3V8Ug1vwc+uc9JAtHbAQz
sArjjuJp4twhSsGQbKr6J9AXFEFmIWn/h/LbmnmxtTwC2//Uo6v0GGJEN4g6txYQ
AQsab6PSxsoUe43JZOAaj2r+7rILuYE4GNh9rBlMAWLquPJg1TO29UEtgadw9v30
NHbT6u46+Kj1hIDu2R+ly27z5gZTjDfLfTQLjgjW8qyNNYPn/ggGjqDdq/CCBEpz
fYs3DO5KhKuyO8aInfj42Dbp4XQ39miUIXRc2cyONCmk42C3jRzpVhwSDXyROKx6
TCEAda/iv/cExeW5Ie8EwKRjuc//mVuS8R/uJUKXP0yMB1AIhCmpz6MOie2szWQF
a4RSBFMTNthYFmx8FiyH6MdPXbFIC8JMd910NKDHG6jzQS0mhMKq3vcsZjJtH0Wy
2n6j4d23M4v0qiDJHEzY7bvswXpeI88vP29TYIJiI4W3IZhRs8IeHbNxoxCHxDb+
fwT8Qc7ZUmfw2a8uJ0NQCE2y5otVzowMryjhkjWOt0gMcdMlusWXmN/hBS41WfCR
0XavvlX6jZVQoMoTyja/lXrQsqbMJUwxdM8AIW/wTtSX3E8tp/Vk36qaIFI0d2+m
+xLm8uGrvPXHSILDkXJkgP92gTzhx9nKWZBigcWIhzgAob16ckbIlkkCBZGvZ1J/
E+gB1M8+kZwI2kgeFhFzZqFDbr7DEYA3xv4ecO3BskDU4y8IJM/yFY3qnB1Tsrn3
fDu9DBNbOHtln0ZHjSijRshpPCXe12BOj6Vsm/BO+NP41rEd0L8syTP/4/MK3WCb
M+rf0M3X2DZIaVx4mci9JqixllAHnpURvUNmYl375Z22XWTJE5IMYFwKgbXB5Xg4
q2BwAUjMFsVMaDQYGE6ThlrPAXwmPOE91M7ns32DYia7YFX8MBAo1L/OdZr+jgbf
Tcj55PkBnuYd7jUTJ2+30rClcxYmt9pADhsfxhDUre3i4mI2sVpTRNqcfGm4m7t7
AWye0AAqHYNycxlUwo+/pLoD0JCbgdf640hfWE2JV+60Cz19D3+dnVHbaVS5iqST
VeQyeuZuQV7DS8sJbbkq2hBf6EXkN4eQtR3NI3/cSpQvHP9i2PcgMCv81G8HDdeK
GhNjBuJPyBfvVdvQZtV+eHMTOvq6+g83ihxU0sF1y3FD7+VetaAir+e/ErlS36Du
q2BuDl9wIYnJQNh7oAIcMcNYhVLnLNz5pChmKKTPL+1GKRf6EnknLQ8Ei8eSCYVB
u56fRcuB4sfVyFjDRXKKt56KtEPNvIFXx/HebZJk1mq8rfMaU7Ujap53qy6n3/ZT
DqBBrSxqhnK2UE4ietXMCpSOb7QkeNIPhN9D09Ky1xKuYe5xyHg9rnwgJgc4gy1u
3HepESsTESypqdu801cRor+jvx8Uys87wB4/fWw1oKw2XtreAqkwbxmVOnTYP9Ka
Pp8tJWXKULPZy1XGE8bzJtIzCFm0emeS64lEJIa/UAlLSWPtNIDFqnjOFOmPtPMi
eKxpJjvCZSanlLNoAmj+yTWMjUB8mBokMKlv56FV/xhGJ9Q+wnqChMlcH8YYHcyv
6fnCFfJoO8wjdxN+EL9jOYvrqOY0MR8HDplAYquHoLi+HJeJfOwuv/9nouao6cHQ
m+43b/EmrS9LbbnDxzoVgIgJPNWEpi64gCVgmNWOcbJpN9IaHdwa3mGwdcd+J9xp
asR3eLYaTvpgGe3AjGin+e+eUkpWJPCwCHQwi8rUcUG/hkdpFisb5/G1B0GU4gUx
b5ixPYlraiN1FMAXNmEg1EdrC2ef6xNbdUBOfdWGtM4hdVWD1Gn1s9C/v85wrtLr
R2a+TeDlDsImzn7MT/moLY2lui3U5YS4lnT42Q74yWlCLzd7esWrot7v9D6zQw6u
GNZFlnuOKOQEjqF1ZK5avz/Aos2Tx9c7vTeHoplDKnnbgskWii2BXatW1szIYGQt
6DvZFZsoRYwNtknfjh6oGfvXM5ujociOIG/PxpKITPeQJuUOncJbJSCF2UnODYuE
IZTCGKD63zzwBUgsCVeDeW5v5HmRPDJHcNselH6W0JWa/ueBNYOzWg+3CCI8BnZE
SrB8SAk1mxsbeNp/y73HLvfMILJ/jVIZG4RhvCTK4t/sKXBJyev9F/Qoysye1KBZ
6A+/oPc4t44SOrl1NP8EWK6xeW9MHOGkIRZHOpm6UejqI0RhSmLHz3PYT2dBC8/8
kQ6/jBzyAaUXcHYs8h26duXTUpqdrC+XjXJV+VUY5hpotrWAdL37bhT29xzfMKmm
VgQYkoGFVvHLoWJiJV0eF9Z1HyU0n/Vcnwo/fNuQVt9J3LLsQPz7ydsoDaxHWMIs
JRiTqS97F3zCdRfx4WKLJQanJ7YbfYlkaJe+tu/7O8dI3gc1cXREicfD8oCMIdZy
ks6QdU8KQGRFo76+Agg4pNWw28PjYuc0aNoUxPPdP9KFt+EyqxIPWQYi1Xef6Fom
cpfYUyENAAnfbTXOsJ15YMVaEhV50U+d5qHt/7PLdobOx14fIPVyrcecRaTPzPhc
gAi8neUxg2jsjWoQy5jUkv+tNUjS1N9BFJbmc6xi/x6W6JRPckGhDiX0xWdhLKD2
6vf84p3sbgYsPbftgk3xjO3rUhp5oNSt13wAZ3LO8H9ek7fJZKPlfa5bhV2vU7hk
CtklP8gob1FVYf49fkPtInIzVxOpw2zdPHhrrrRdlz1CVRccJBCx+rZINGLJLPH1
BzUYOYQdoITRX2MCWlPS2bjyWY/c/qv2F3OPJ1tx7vqseYyCMbfrvdkdfCFPdcp0
wrkYyPKUtyH4JwZkbOlE6HngfFThBUtbL+0F4+mFffAy1ZM7Z0aq8i7RrIySQxJf
gxVO/ZwiaOn6gFmaPPLyWg/0RshrjaCNp22+5HK0/WWAZqnQqjDdcZFSAOguzVGK
XzWwtG5ZbLsSETkRAQzLGNaAQZG+Vho39Zbgt9AbK8X8GpFb1E/gbs/BTAgNL6Ir
KG92l8zbV/3IfwFrrhiA8a2fS6P1ah9hKdl+Xkdc6Z22Ffw3tvdjMlU0CuE8+H9l
JuW3OA7mHrhZAY1CglB374zysE7ecOwXxrafclwiTyph8rB2ojQDs1Yu/sPZO5xq
htPRmMzIJBOvzwmcUp5Lfg8JzT5tIVBL7Ga5mfzsAlSc+rIKdTG6Nz8CEibjPKH7
sUqrcsrJFmJnF0oMNMk9G1PNxt/kpuizBnUBL5FxqwKxaw+q9GW8yEDn3zEmP4yi
rJFjVF7JJeORRUAQqidjaeS4S79WVIKfH/UkL2yXb2Rw9wRMta2f8mdM9G/EPbCZ
t5jFojq2v7K5cK5WURKenG7678I5TeenT+0Hbd9e0Iv0NzRtfIfl8kZl72hWzotF
If4+kKlDb9SgM4SD00h2SvrpNUkxtlnLFmFgmc42N7Qes5lZSV2YQStdQYaUg1+Y
4PFW4f0K6HBksduyp+LubvPovJv1gYUeyYmsdZJBgKLL6bL9QSH2B9zjQ7yl9dml
3dY7MTu1nfcT2XnIbSaYrWihUavy5YHbZYKKRVV9nrPnxT9jhbnTffwsROYXkTj9
63a9lD5l9OYgArX8/pE482fX7n4jw9rDKY2S5It9MERbPli/e96ivhYSPbp+Un8J
KGCYYpInaeP7FNVIIyCFRBEwGPskRZxkNbhqM0YkLZJjwflJxQHEm5LeOkTHIQB6
ywR+H2zCVenpBsiiS8YmyoBUmLo1jwOYWtuFptd9m1crZZ6pmIt8yYljpRgy1or6
flDzbdFLolD5GuDbAEDw8FDou+FIpMPAtjM9LpWDPWOJFPj070XHEBwiOan+8Wss
l6I6MmA30qmR3QwBXNLu9f3jo6vOi1mXWXaj8nV66klNYbvvabgUfvzqNE27wvgF
hksuiqVI8/udwJB2XIXF1zAquduTQSIdOYwiNLG7S8ZsYJhzFghgSsz0COV8Oagr
84mR2Q7fYmBn+jdGMfjx2M0S63tx1ZJE5gRmdNR7hrR7lrfa+LtYL8Xh9kXiXsY1
OP+Uor3GWaH/bdRIA3iImqY7qsIrjKXtWKQVwQxURgPnDzoTYFOuhKCNCFehz2qM
QGeObU9FLobMYNBxULfPUp/43lY+U5HAe/l7amjG/bVt7/6iXLFLs6ZHdb42Nlt2
ECEaY8avzvxP9t31wXvr6csuVOMI7DKhwpQk1Gwa7Kb37nCuuvQItfdF1L05teQF
o/t5n4DYrXWf/PBwrFahPZCwy1+FaIGhzz2U8xUd4sDlRurPJkAlo6c55MZFD7Xy
+13S+UfHHBHiL0Sp++prOgQ+42Yjwl+ulo645WlTaOMr44XQq5ltfLhtAC6kqSPp
d8wvrjk185oQtdi2+hmbw4n0CRbNPcWsIh3U/xK419QoMoN+bLB8AJ588cYDtrX/
rSlMvUzL88eHFMusHeoGmRbBkXhumD7Tfwn1GhXYSjdG1gXPuoFRq0pWggkFRpK4
+/xh9ugWB1MtFLS7oI2X4eBEBMbSzZDoBZiAsK9Je6geXf1+iepytRizxXmFYAWg
6pBhuAeGrPiHF7eD0gVKA479BizhTRZ+Nv7YnlqwHdh+enEI4TLHe9uEHj9t49IH
iMWluMrf6xtDtL/uxI1c+thj3wwNVyn8CC5L2Vq2vibOGYozlA4ymXhVUVuKoRRP
/CcaZ24FC0XGFI8QSvfH6+v2g0BXbffij85kbKkLC57YgduJB/Sgc7u7KeAmPitY
Q/tfokCrAJ7HxLP60aiYPFwfiu5HGGklIhc3fY2qp8iyD4W6R7jD6wl699JYsiRN
SDJ8972OpVa/Qye730I7752BdahYrQ4oH/FAEZb4vQ5RnYXnfCNphDKNagadoClo
nIHnhHc4LV29YOKKxnlikxT5HJSW6hHCn9Mlg3qLI3WOPmusykKtSlsjiY22ZWKC
RCAGJOpaZJ+ZEPdVAyNT+36hf+3kBQySzNu01du2NLLe4AZJLti/FrXAQVH8rfQ3
ZLdVpwUThQKPfrRRac86/+zryQwXwbibJUfJJdl0Ad2dFcOGZ8Zr3YACpUZKG435
jIcu8SPpBOhJwT/Vv+r4ZyGeeg+w7Hy8GwL+O2lYWSvBQV3oRhAbYA7YaMokl+Sb
nkBIXdkVHELrgnUbf1of2YAtOJE6qjSQXMEA9l94oC9PgXzF6mfhCFTl3u69GKs3
z+wLD8PIKn0inld+489NSV7TBVTbyKHGbNM7iqguurQdFSav1A76XM6LowBDMK35
yFrJwibxtpPWB2bCUA4I4UnKekUKu4WR7dyFOfkK+p/34n1qooHas3rNXFOXZhSG
lOxEWS0GmKbftWKbu3u+ihGCcjvBIWeq+rAKwRk3U87xRxpsFxTlu38z8xmsiIYX
3zcAHRLyDthW+/7ZcUjH1RyaW8R4gMpS4EdgmXpcOc3ptrRCijmjxGuFMjEpO2Pb
2GS/eeMdf0bWqI50r2tV1dgEjS6SaWYl4RBb4NEyNSAjQFIKoaPLab8C+l9caO1B
1/7nvH13qvtmoXMEVNXx2ktl2G8vqEDFKLstIYM8w/reSXB3IO/5gjTb+m3QwQXQ
i1qhJJfd3h6oiboSfdDuaUoRVy0Rl3pG/QJkb4dBjTwtwDHsi5vRfIXaomcJXLaV
qoNrWqsTslgXVxwHA2SrZcmUtbPc2mEMmH5hkxv52kPSlGrQavL3l8p/AMTCufW1
p+5l6V+TwYN/ksrBY2OGZTNULIX1HZCOwhAdHl/QQlbsfHOJoRdod4x7fTajnjiL
IomrV/sSkL13vFH1oYz/ep7zfjhBZiD/Oc3O6TM0/OmiTQd6AfopM5+9I8Bvj1iQ
DczIZdRV478j7cZtQghtZ055HJsHvgW6SMPJsY/LYgzVYG5eDET/oyw+6rDKkhYt
zEOh7RDmXXQOBJYl3LzZfAdu7nVFcRXV/A5ZRcmoSge/67XMZIhW40o3kanotA7e
v7aoFs5b2/7RwZ6A+GX6VxlYTYEkNQqlp/3TUynUpJs0SOVG7k4hPQXSwHbYyatM
KWQlrQbgk9y5a923Akx0NKbD/oSrtdnxWGgNJpFeLia3AukYqCoYkmBz6b0KnI4t
bCQ9hMesXSZUDdfOxzVmdnF2TPGe6xcJ/XbKLQGl7tk+tMvh6wVDC5G3M1lo7M8B
pLzXugZB/3n+qvAHSDYfRg/6ZWnFecq1WMRm2uCRBTTHsfTBBZjGB0UxyVs8weCb
bxRW7CZyd6EA7Cl+3bXnht+y3VWbQUBXWK9sdME6z1ZXvyQl6XlMmXfb8Z9RpxUr
EGYCwBZkiGrPtua8BE4ln29dvgx1oPxOpq3Nxh2ScIGEXFLQh2yWKKvQveC0zrUz
7L1gq3GO6HX8wjrcHUlGnz9oNmfozihHCmqr6tI6zlhXmTA97XlTcBmj4wNinYU8
uAbem65ON0x7Y+PIsvlW0VOpOUQquOLmgNIssqVCuM1Me/3H3VleslrUZ+YYVQEG
xu5vCv+xcxpdu69EJvr1pDeDQanrsrU0AVMVgw+Pu8ABzkdzHzPbKyiZp7odptvg
a85paJ9Rkeckx+IkdcCCgkkON/G4CB5TKm0fuWTmh6ZSJGIgHq6Ka0scY72qv0bA
/oVgUNxSL6p0vay1m0vES/HY2nJCu08L5DevRTUzz1KpZm8gVVpSiwNt0TnXyE/4
otecMPMi4c7WCqZdPGOj3rnvjams9uKlrQQH71hN9DOrRbmmHtqF6LrTR77b2F0f
aiJoVEvsalz1TGzr9o5En+VNjZep1r4c1R0ygLBQ9vhRABnoAYDVnifXHzcqfNez
ZjXC7oZl9Hwg28wqD4FcMjM3WLb4+TZaE/ZTrEDRvlJjvIv6iH8X478e4Wde+nm+
0Ys/Z05BGky1iez0w78tA7W+oED95cK28UsKCTGekp2L4HqHjEvgnm3+WCX9QHuB
hCH8lqlc3E6Vh5JxX+pqziuhOnqHNOuhOQYwxeIhHV2HwyCVmUe2PP6rUTfG64mt
ucN6L7qz3uFkVJvEQwdIlwE4B2RISzHHUfQ1qLNH5Zv+ZQakkWSDbJX3P1fBuvZl
0f6VtJnbqXjkn59Tcg4riS06qEFsiu0lirrTU66s292Nyc847mNNtdjBwVdg8ZvH
CnyJT5GBNojZaOG8O2D8lJZZf1FHr3YBRyZ55XHUGkRNyqGB05bsQHRL5ELwed8M
oxIavbpjOQyr+zZg31dy9Q3B4tbK1JeJkm0nu7HerSTm3PaKtHSLgmX6owuckzqr
NgDLj60nYQR0FbiSXOjnKcXvQeOKF3VGHUwr6yu1r8uxeqkRGkYYBdXI8iskgMcf
wY+RV/f+wfGz8ElfmxDr4avhbk7qrIigG0r/QVZMdSQDqQiwMr4KmHq8qaz93g6i
L6vfMifzI9m/BXsc05Kk0aqvG/U1EqKyVMxr5u8YBx2ujWGDgYneNSVQpwjSvo4z
9pSIetuKEnPQofxJ/y33CQKBh6kIkWbyJMWW41Uz4cpQqjaAFnd4VCx/OgTXttVt
s5FTPiBlWd4pcKG2FtkrbnsNUlEwVEgqYeNrdyEc10288HHp55qnIM3nExhVjARF
E9Ft6cVLJIrhPsnRXZPoMumbplw2VFClcEhx+1baupF3TyvM8cVHlnI7sCa1XcQV
QTp8Tj5o1EnEgnhYO733izetZhZfaRrCwPx/2Ce3fUvCCyoNL6mcHQVQOip1axdY
sFVG0rD5PN9QisRXrlF6ZA1II42ImPffH6pFEejSyIiwt/HFI/sum0OpXSzoU4Xp
l0FCnxKjIJojEMmu56rSxdqiB1LYa5ub1vZJ9VCmkurVjrRNtJf64+2pCh/C915Q
xHltqnlC2CGhGtz5hZR44FAdzu4MT74+EfpmUmp3nltHKVVpHVzLtdd+YX8Mj+ek
K6j3Iooc833Cv2cNHlGSSnsdDNVd3l+zMqtoFu6gOZhUSevmSjojSeYMIPHQ3FND
YP2tAnhpkTI3rcrEA8ktQ5jWklCCuJJ7Ovh83mBXIBlznX+ct5aAcmcNyxPZyQ3K
ikufR9dF21riK7k1PJzHT3IdnR21enQCMxkJJWOBXRH9Bbp2aBDXBGknB5CP6Sst
TTNzzGuZaoytKKj9X4SbxpPWgy2bybok1qVLF+5DArEp7KEwxdu4MYtJHyuOppBg
i55o+vkgGvc4GnWPgJxhpkZwnuGfHi5cVp4pYKThLfJ0l5aquFiPGCQiA+qiBC0R
dKV6RIdctIksknScPPNqvdvifIELvLMb45yP6Yv4az4v2AJa0OeXqc8T6G28KRJP
YU1VjrM+evvLDsrO2Jh5v0l4em4ORZazfC3lcWQH0E4QW7mKt+klgrN2Y0lQG783
BUmwmT9WpwHFGcreJWlPJ9L7j3352rHruvfLCEk//wOgAP8FIKHNZ9zDZIBfXeFB
mMZCB+7Ab5vzuz114DKjrNKTw4u9gI8uynU8I/tfVEGNxQ7XyubYhAoD4vgbkinb
G9xk/ipBxjCbNH/SuTFgOYVCjP45tJqNi63qEu8rxxz0wPNEctoZ2P8T9rP7B7+j
IeFPAFal5ojB4La5JbaoGcRRGUvqjVnGVoF0343pY4945TYj3KjqRYICw5fm1A12
8bIXB614tZQ1Fn+g8VrhIXCHVce7yy9V3IKPA552b8qIYl47tvCY9q61caOUXjnT
fH5+0fcQsLpWyJa1HcjZvOQ1y0ySQtYmKYDDKEYZsa6fOI1ZtW/WkwhFqnlgoooY
d7KHFgcrAS9eWKbhGv1bsFKAFgs55vkXdR17l8m2RKry0whwU464RJAmPhURbG89
SeqTKHWYVApLjx/479fR9o3lyZzIsfg5+qh862XNF8xESRCRzcaF0I3yOqh0gfQq
fH9VXKeMdskiY6Fd9C8VT7IDVAUkr/C7xyiuIj4B+/+bycc4RcxXEoVM3t2AtO3k
0NHNTN/QPBZfQoHUB1s2WFmBXdLAC5G20oVB4H6vkPPILBjxs34PKczS1ixvQevm
ZYYZcdeq2vLIIhCx1sxBS/OmCphHFNMNTJszeiz+sRRUkdLMVFEHNZfGFIAw52bw
kpqW++JOZMdySu0bAT805D3wt6yWKsasNp28mhuMf8bzzR8BrpJkjFuYAB3KpP/9
9arI+Sj4Uf4tBrnSsdxZXgBlJDa/GkbTvl+fejB7XUj+5BsTBAKPgmjvhH0y8m56
w0AsxXuYTdvFZKUA5wIFAicvt6h2ml1WDg0u+I6hBXzyK4Mox1sBjBgh2rmhVnhe
+CGh2nS6xMgBDrdCu3x1JP0pDbHF5MlQ8dz6PsAk4dipCJYDrqJnOPgvtSXXDYkD
Jhy/ppK9RnXVoyqvmyTwP4TfJz+j+uL4PkhQlD0N9wLHUlTjutoL+qaO2UhhHJHC
4zUnNNDM+jGkUvANFPjS/HOPM6uiyaL9Ps8LfAPj1xsm1OGv+tvypn9TS2THI5jm
bYOsitcnm/RVQPaFS4iRUuBa8OTZWLij97zoY9KZjKn8C5vTPpDC/1eg5zwqQ3Fb
UYABiLuDSV58fI1hftikI7ip6b9JnCDiUONSV0GDgRS4/JvUgvm3wUKm7fqcGgMN
Y+7QYR9h9jb5mj8x2i6fD0heWusCgy/uEZzehE87mOlznpEB/PHtwUoKOwlLOAd8
zcnXu8fdOyn2HtbxUdMVsTgGy8sqZ3UCTSol0ZxnD36V6Z6Z0ro+WeAYIStnsW0+
M5KI+XOQVEd2tGoYDr5N8eDOqHWM+AZ09gBfRgW0vOQX27Et/0+OZQg1qR9RCbgU
aa0+wnZ6hPZyVrNG4j0HD2J2sypVqFgySCWbb/hovOz00K2jomgnQa/u4QOV6N6g
+oCYTkXpnCNzAw//DIdPY5i5ztABBEBnaaLP4mMpq8Q0c3mprRcRbnj/Oajf1zxY
jdrbtGVtuq7O+jkmOp/PbsdhdWcB6pQLZpJjQSK/rUKvz4uew+h+l55Q5mLSDMA6
ER0Weesm8rK5fQg5OUrA72QFdOJ5UtH8Nl1uOG3NAy0/SW4volOKQyPtH+ZiekCu
ipH4o1xCIwgcSjKJbgnxoEw8WNybrq9RdWIccqBVLdkYklivBoP52iiZVHqbem0G
8n+/qibwDUF8L96tbZUJ8nv99QbiymNLzC1uD5kH6TuewlAF8G/wbPIeJf/ZEerw
CLQvZcN9QLMnm0lv1LcJyrW3frKFkl/rDUKVOFg9QH1X4/W6U0idogJa4hmRKzlU
cI2gQ6Rd7aFvd0DI45mx8O3nWJVddPYxujBfP+ooj3M86nSYuOhJ41CUFy0n2SlQ
4ATeKIqnnOYECDMuHwdrFFlsgbXDouHW68uXhStEC0/4d7i4QwJR8w/odNcN72g3
oaOAk4V7lh/NKs0Td2LtirtbwNUtj8/CIdMM7yKPjAH8FLSWeA79YLAt7BPLiuhD
lzRVDqFiHiTv7kN58u6kxKTs8+IPpkLmPUw7YscLQESeggbfSbUnE2iHaCMoj2M8
/59+DlFe1/4uAmQT0LIMUEpAOOB3oiarW/PPUaSZORsjFJBHyDqs+6BrxShdyMA2
W9Wkdukuzw+LhDV8iEuehOR65ZqkYtpQLe0GS9/UWxC0/jVWPvWpEs2x0eQ3rUDz
VQJiTUQ4xwvaPfrT94XTDOAGub42oyu+T4bra+fD33ukGSxfTw4fljAZygeAtTfa
Njl0Ut37M8jafuDUaJmo2IA7suTY/LgVmdanOrHhDADFBQScPjpiFCWybxnA+oGY
YjAPmEo6DtlVb9MYocilYfAmXoTNV7MspcAGEKyVf1GLBP+/h+l5AfBljks7+9bs
8ZIoOjsaQmAhc+/hi/0e6MylcC6X7gfiQ5HTPSe+0fmFiCW9YR3GSEV42NTbR+Li
jRffhgbg3yKrBiEQKr/j6CQHIShNFP690ZlLEIBpgMms15HaGTCyGFAUBGEd9m+f
hxLXoinauum/Xfj/sO45uLps2HP8wZ0dT15VhbRDYwbZaiOEWm1rIPqO7/cEzehl
LtyhhaySDwtbklpXoi8kNCY77rrpf1y81LIVFS7P0IIazTaYqWNmVFJemIMceEhQ
2CoV2JO20NL2hc9UnIl6J3ftwXokPW30saYPK6peKO4EzNm0xBSD2ycJcWNKva/n
y/NC4DjXL4a5b4pQOOD5/yjjJru41EPtCtyK4wOSIkXuKPqJmaDvSgM0loZVvK3G
hHNHvNHh+oYDhKs6AMgYogxF08KPz3DxtenYjkPgklQL3PJqUC9FtWZ5GAXRoEO7
Xq/JRImkpTSOqGmnlhjuC2dNPIOLmkv5qd2bVovKyRbkzEz8pVyLBbSLkETUcqHa
djJ5TzSHcsNgIu88ho7ifM/PhhichsZ47g0Sel3BIi86yXnaiPPhRuHynWBSFH5S
rq8CEpDT7scTkPIlRxn1Z4oxBq+5hl3Kmp7nTLUTNDhrUiySZnkfPZfFdVylR6w/
k3VHiEzCAUqNNghCLb37qj4n/KfB4zgl15HPdbbf/p9YXC/nGFCMl2wsRI7srfrF
DQz55KNrdmrUxibqXpAnv89vicpuiCMpwRQTHVDAqd8X/5X01UvzVn/lBHe6u5QM
09++YJB1MCTJzEWSNrPlxQb0/o9dAfIv6wilwPSyoNSi6rocghuRbIOnn8odkAoS
8gUlK9FgGU9OPwXqebRes81Vqg7zuJogXlY8SJDqHbYxliBMevRkJr/uUeTL6iVX
YsYR5yZcuGUNK6KE7tdt8mdkkg4j0ZacVggfHzOlzsJFLKMXySwZT0+x2ZPlIdIK
i+1Hcs8Z/5BM3EIJqFA6jtmk2N4+Qb2ZrgYa8n0DI0gAwRz3prh8DtZb5kRJxYij
0XU/mHJPQtaMoNKKCuWfEHJqUbifH9Z/2WG89AcFv1dMo7MMVlr95e7X53D2JJmY
lrFaORu1t7+RxGMR/ACclzx+aBiNZtFbRsoikXphyvdLXfx8KJcEVSt0BtveDlap
mnFzHFxXSkCnBmbMD0WTPWwMHY+qsLNP64VDV7gfnlPqVP9IID4ljkTzEl85TLXp
y2ccdB7cmoqBwyyi/sMlv1clCVWQBbRhLIt0k4cwcnQU5YyX5Fip+j66SH4TfoJF
0PwxNbsxi53Q6u8x6nLphaz/wGlnxccBidv6T+csFhQeYCAwnpqygvTvgWnGZZrI
E2BFQ0I2WTkgO9EeplT/NA3BlduQJtYVbfeX80FHCgeng2sIBuwAF1NC8MvFYmmi
e2jMOcRQTV4PoSiZk60Py7T/pP0f7+ns+XgFdtv5dZ9X4yZtt0osZ9HCm76EYWw7
aG8gGc9gmZGooMUoU7W4iFGxaWNEfD9g0XS5IoEr5MLTaSBo5YOnWpoYWhzvorq6
rlMfvtaS8TlaoDwH/tUKA0n/vldzlsmvEnW8zKajmI57Zzul9I9fj+Onwk7GEvFn
X1Tazl4amf1n/f0vHpY9m93lShxtE35e0+h8cyEVBJyFtQu1w4qtPQ4iUw3W6LiY
m7zi4kojV8vRd8X1ueZ1yG+I1SR/ab5d8HBSABnMgD25ZfKzcSQ4dmdQd2oVu/7K
HwoWy0UjKhM3MGhW9mjePDo9PXNoEwGC6Q1va4qlBUG9TcU+iEaK8sdATexnsdud
X2t45poyhRz/G9pM6/bZWNwnv/ldfgz4s37a5VBlGAJJZ293S+si+TrVfQYXMvon
KiXObqlMxVQGPqUa3J5/bWbgAoUK8hKtMHBUGTrYtUIog76yuT3Sl+lJZKRCPL+J
X6RBlVDqfRUx6ciFKPAW6Puo3pMHhewAxbgRrC4R4jBzIWRHkXL0qwoMeBzzsn/E
MFj/ehOocxJj9A544OWvO9MMdJZPtJ8LasIny4PDvpVoZVD3z1qXUhHM8WggRTiV
0tjqNYbHSQdq/Ffuov6VZHHE4kBXaRbj7491hhEHO9yjaOL5Kb4BVzMfBBrTW2sH
/bjrk0/CprcMLYdg+SDSDjg6+GUPmVQVtNJkqXvkhyLMxy7bY85Pb2jFNV5dAVuu
UQo1y/kp4wNFFhyLNLxeFM6Hi/GARh3McVQ633ro07eLu8HcppenY14SX9uZLHO8
d5RAjLdozDjV6vZJLVnXhOen6YEAFQUASHZ90pXmhpt9/S6LH/B8m9+Ph/pgXBT8
dgiXei6EiMGKC+ch8yzggrAkZ1dc572qAS+mxlBpScrr5jFbAi8PftCUo2uMR7fg
BesK+BlDoLSOdQO7lfIf6PeJZVKpTbTg4EgxgCFCU5ol5xshv3jSEhMJCw5NHBCF
9f5VwCXUD/MBAAQQLTNct6DYSqFns0rURmql45WWr4W6au4R5V/AX4rKLjEHyYIo
odw1bYuy4HLj6tsRLgkRI259GIvp+jSPtpJrTD/EYavks3jjlg8VFqSAxPrfTJq3
qEBW+Nzdtqul1p5xKg0f9qKzr5efDrQ0YwUY+x4xU3Ezx8mrEyQG7ypKZU8QsLdB
NoyyRn1ON1xZl5Ge4sG5wTeqZZpeVYgUor87Kjct9+syT9wCj1oRNBxAhfPBMZom
LJutUVwKHKQnmRHoZNDPGE/H2FJfdn8T2vKc2r6afg42CRq/P23sxGXBu7AFBLBk
W49a8gWnATtlbTanXtM1QYuQ/nnXaDQVn3oP5cYkh4D+hugXmeeHq0b0jmpRwvqf
i8TUEg1yK5sNSVcMRflq4kRHbOOM/R/2DBYf7+3Xlsy4wQNIjvKfxl8uJJXWjSSg
9cfBvUuYBQmtzJfm0X4puJ9t4jG319xQWQe+HaWBruwCs88Ldz+KF5iMND5zRbl4
oAmSAo4ljiwmTqdHYw2sxJtvnu4JDHqT80dQ3r7tj55W5rkZ8D0742DWjKuMKmRi
Up6ICAjUHb0+WWTq7Xxx2RjPZWIJfA5DGf+pOtax8/bp0Hk2Z/jXNCWsD9QgtqKs
p8CSPR0Wwruv4Xi9f/sZkpOBJRE5iAg5/lZ/YaH+FDbT8AUxng3xzEf4hcdzWesb
Yejuph8dfEDH5ArNzzO+2LVmvqNvYjyNjYcsSCLLpPc6R5+Sb3GfU+25dbOb1dC0
gBiL8akY4GHEYIcGmoWycckQJhjeBCmpTGgUDeH1hH0L3TQ+Twqzyi0ZMP5ZACDW
9MkzUoILR0BIjNRySl+xJI5cBJ//dMnsqHT/LhCBPrSFllI2QBZ6AN/r2Cct/uWY
BPmBj+abwSCdKIK5EqkHgzvpWqErfbOczev+jyvoF0rUix8b54M+9zKYNiJpqTX6
ehHaehxZHLMDohfjgb94xL9YRcjNNeBW9wL7Ly0LkRpLOSWTndvHlkUe+t32c0/B
SoG4uSf62KtTqsk/0oSqD1wDuvjfUcXcdYUhxpwUw7JMYK3qKd2F/tVCqKTRTCKN
C1jGbp2mTQ+z6HusIFieU109MzDPa9jsJ0y4VD8+m+Olnc+7rwOXZARRtp2m8IzP
M8EHefi38vQPmWCkgOdfBHfknA7o4psR0N3hhTA5VapYDS+EmtcIG2j6EY/0JF8R
filLQCCAH3gp19bcJ42BsSi4nDMvr0Rz4h7y4QyvkvtoFBXBA6H/46/AllK71NPW
pL5Awd3xNCl8qlu+kWHp/kRusAaGxnxu1NHO+p5R/q6M+vnDb4/164d0wunmcIgN
qo/vILFxM6xhcEuU3ofZStHyEuNzVEJBDCHvtvgyu4nJ4ztCrIV8frok7Kftj3f3
ZxISRNkCC1EEXEDJtbjBRR+E3zfJnHoj2S6E2eoxmyvu7MYN78O4qfH2dzMsMoEG
LrlqvSVDCavH3CUxTa9nE8RZI+a5JlqHi6szjeeYVm9LJNW0qo9LmEXQwsQhywdv
Jxn49tGvXs/ROojVcXMKWrWevGmflHt7iKnq+YYXmVb2ooeYwJIzFWSmBHECGlqC
gKkhyMDgEOm5YL23tch2SUsmP0VrtlLOIzM64LfNv4DRm1ntmZGR4dqSRVVAhtAJ
jK3ljgPa16Z6RYR5B6m0QRibrDjPpWOFxfSBodei+ZRLjKlzdXxmpEwU2EnceT8w
4jLVveQCSu0s2glX9+76XXnpBT6A83vRyBkhRG+4g6EVcq9sDdJuUskIjsUQMhfw
7d3+daufjQ/h9sn5oIN61caOW44jeXFJenkOP9EJ0SQRSzOPVdBQJTWFexWvgYps
zvsBnl57LQCNRWV3dvlUtlOfRcxc6TYs/GrXI9J36/1fi44mz2rn+0gdayJwib0t
FygBasq5jGrrpNqWESmZVhjsGQ3/4v8VUsSmURyb/dYuXkW2pbuEQ7YG+t/MydwN
qSOD4ko8s91Cdx8+uL1Yu/X/hrLjXhLHirSCIJwXV7bLhIx694nRydyVKnopQ2uj
OVjnmLqqjRtyHsw83dw4ENvo1ncGFEGEBSewFDYfc+Aco1qbXUKgoH3c7gaGtSAe
plIdZ+qLjGLjuP+3Mkt2FDRHOpV1M87k5vFrb1xnQ316+dLxPSB4Tw51xdaEgKA6
L93jRGYM+ct45Yn/87VTO10xcUdZ8fgsuP8ksQbCH0kOEh1z65Yjgb8AoHN69bOs
QYH5OBooj38zxH32x6T1lOU6fFEGfLM0vZCMah5hCYp5nPmHNF63cCvyYSHRds12
ztfq3gncEATi7X9RE3WDh25FfPywMczISrXvwgqz8EemZm5WuNh4mlXKIGy1IO9q
sOlNgPr3oXHnQTPAbp5YQGV4V1ubcKEKPpSv2u05R4i+R0MZcgnUrubGEUsb3lTc
hIKFtBUID+564/OF6iHc6fOsHOQ2IdIcrAYSRXTx5EQ404kxL/LiShLSjUVcBP2y
/KmB7GLPBtc4RRitYv3DEuxpivx7Mzw9xlfNMmHKVrUcYt0wY5g4eFnu8jaUPa4X
FuMoDfOtRmKM+rFpX/3H6dNu3ed+wzvW+uHfh2+hPpd4+DhqYm4XFzQhV9ffhR++
ZabnYigX+8BQPauH79SznCYrkEdxDSt6lGKjrWdYlcSA0cvTlkk1sBFZYRtjPrAz
pjk8OildWcdGo8Jh6nOVo6EfVCnlqPVfR7xf25DrLlOmhQjSmPUAaSJmjD6s4RT8
t3DCOopwBz6yYkLAhr53K9nVwAhEFFPGyK8e0LeD5aFiQw0uh/yp9I9qMRrslM19
0bK+1MPSvlOY4hxHC00Gx6OnGKaM24oXNW0fdKBpIu6jOokdkopSzYV5YvH1WaQl
T65UOTG1O+x5csWW1uxTJhYb8oH44tf1Lo5F+sM+rKuULxuLK7uC4RQ7vl3GmK72
LCYplPbOa9394lx/7fdWg+QR9g6kIcyURbQuZgjv8W9Mwbv/QJA5JEKM+xNzFH/u
XvqgFqGTtanO7V+CmSO89qvZycqjPSUHVMX84Ue0KVvZEBkmqdLX8j7N59zuXEgD
mcC7njx2Cn/U2Vz20afBa+zezgluVTik0Duj2a65xKU6aa+AN4xvZzzAZO63/tpE
wpcUq3EdyTB+g1jRuz5q+kdpsnVnL+1EI43PttIy2lAOpfuHQ20hR+Cg4z3uzitr
o+cUj4NDhDM04DaPTQmWKFJhCP2KB5b1YueTEdXfZKZBckAQAZYrVRLdVqV/woN9
/rAqz4PVb6IlCkIRwSZhMS8Ir2dzQABTSrbLUVl9hcJMtXVCpRxdQgVwkKdfWxaV
wE6NfFnnIt/tgT5DEn4f9WBh/mY7iPh2eyLt5a9PkOznwjZDG7saZ92DEhqTQqiu
bBOFl+ZmiWeOC/Xe7or4InHSNO9Alee9w6PdeyJ7KwfGt0eglfet0ztfTZpubGXW
2PR6oL7XshwFU0jJVrn9zbYj2l9MOc/rXuSvGRnW4K0GX3Csf6UJmCG6ILL3sDFy
g0k7Qe8lZD8v1IV5rRkBwKCuuKSZ00rWNAZMsDMmMun1592fhCapcN9MRy6tqeQm
7x1KxFVwsyLgn0T7XAv0d/EPNijxEXfcvS5x8vrhXWo5leKqZq1mYSIYdZ7rnFKX
76N12bofkYYUnpdqkt5BETPnjMP9eDYqAcfxqmJaqcamnOBNU7S/il8S4KlNriOP
j9KqtQnDIYdTWygQGF3HdDzqRSkEDGJD5hpPHw2VzuC9geNFgdx8GeN5U45QyhVT
U454RDFNNEvKZ/Yl4vv+zrHJmGXMsxmlBHqc/aDBBFHqHKsYpwPWnGkpfpGRMaSb
SL2Z9Dx5FXndINZLya96Nmxb4OUf5EI2PNcOeOdZ/XDSlq8m9LRtwPojxls23OVQ
KQqM7/Gk9X5UTCAHIhaUXeW5mQm43Z+H80XOpXIlHp4AGlWgJyxu7DSNY1qRtAAf
9mDdjMWi5vkaf3QWPXkPbtmiDZtzhDYd5mkrpwNLoNhU2ham4B+LQb++NTZXKFOk
eb2EZnu9/yVY51kFU6lC0NabZ+xqNEHb08XuOmYKeNMf7Wi6aiVcrlXCFlt2Ql/R
RqO327c1VC3FKYUtZhqw/pGwRrlVLZSRswuEhfQzCuo5xTuS5kaWfg6X51CdxMjo
8G6M80TC/f6g0p2qqSCtogWjuX4pVDO593Gw1GLi4nWMrxZfiztaFd3vFE24DCqK
vIiMbj+ipUIccrL+TClShLavx6HtRQIrTn/MpHuVqf37/qJjjbklP4fketaNzNK6
rY4Cb5GGhTWXDPKaB8tzOiy2n7zeedkwBXrDwrRlw3ecFTmvJ4mCPEgi9ePyn1uf
BL4EeJgvJ3NZeCtqHQOElQI5TsHBBgpTPHUrWmVwrGuaByaMM6m1PqpBCzM6tobx
yQsdkJmF0wI93zoeihu83BcCHccA768C90GYqZ287xJOEZwAZ3nDVQBDGvTyDpMt
KcMNoLRVaZeufr3fwieDGclGckwpLzaE3jcwMJ66+sBkvWrSOi/7rTSusJqUmX6s
ieYQRj0qaRdnHDDSC8bGJ7yYoNfC2GQ4qMzvtRDjl5qKV6Bye/RDI5n4eA6te4Af
6UWaxBU2bIyBmGFgZMYJXftlJ/hwXe8vggg+IhQb0zD0+F4GO72w8d5EKY9mEIeb
4tWlsauiif5jKN73SzXOLQTLzjpmWM0LPPVl2TpDoWSNIMQGfiXpmKPACdWT8hGr
asVu9xAk9JnpAHcoa0HHLSi7bpLwJjh/l275cpFi3wOWcBse79SSx0fHwOz9jEfK
kSqk/nWD5kFBUvuZrXAAEsyq3W/A9b708xBh425obVylxdEB3VdFeR6okbtIAHbo
Dq+96Z7Rr0jjQVCId9zkE34r2vExLvUuW0xFWoX8FiJE7XBgKGs8VrzReI4uFHrw
qum9vd1YiMsWaFSkGsEfgzWjeRUDmHxJlwDdpQJ+BYk3DNzCVpbyj2rHKiRKGoOk
GK9vIfMQFI1M6SvpmUin071Jo2rT9Nkkz2iC/Fowxcvg5RNEKhYjzHLR8S5sUYYF
zqQSJmubHzEI4Nss87QYcXmjEoF+Vga80jExILDVUF6rrwAR0EIyMz1BeiESpa0L
NWVI32tUffucWdlT2IycTeBaK83nRZvbQFF43otIG++mJKRLoOFEIw7nJGhfeptY
ah6+LQha+HrzBAl0GMWKnhF/4typmSWHt2AK2WJJhwbWfJMMzSOXoHkgZFMViJiP
nIC8if0QYcnQ31uf3JCoALtci+Lap1pJ7LqS/vSK9vWWrW7+yIZk3MY7woXJsJ7z
DpxqYMAAQZa5gnl6+/QlNlBmlVRfbpd9fconxAjUsIBGJ4L5Y86iXAVs7Ee5fT6X
qXQ16B4j7EM4nfvYZ2eI3GY5xUO9RF79FDKRuAjDURZydcUcgo2POvTGlrstajkW
VfulrEQc/09nsBjoiAWybymWgrkVJwXadloR/SYylHnuI1BOgCcgQcVKs1Mq2/E8
uv7GXaP3lWWdRQ2VLC4/S3pLpxxvH5jEgnBhb/WPZSp418jcZnvmVkVIfHtxqOMe
I6803Op+UGKJVaokZtnlBAdjzYmyhG1eO1LP4Ch546doGfibyvtIlUJzWWsbcqpV
I0zekh6JpfQhg0erjuL3oLBZS4KU3SL6kfZSLsOdktEgnTWnAxjE2iQjqjmovmyu
XqetVo0YPMN/tQfBol89O0cu2jyWXxttKwmeeAgUNsncDvBGSC/tVInmDROdN0xU
8tYfcUi0E4tPxEmkaWwsEZXxZbnX2aBz65RO4UbckrrEhDiK6SqS3eup4TMhPRjB
nVDiQ0jIJK8zf+G6Hgw6gdWJlneSehowfkzzNnlZVGRZFUYfT3pl86+zW4Zv+iGk
k0iOl+yLQw2mmo1bXZCplRfMxolVmF/oyOiMTmXSoGLpMvyBUKrHmJQxBQTXUZxr
IKEBIia7fwv8DZUwFi6Wcumzyypctkn3pELMB5o6ZyBmTKiYeVKkyC0uaz/Lgctr
7EF0x/xfkuRoPK3wv2hN/QITPPELCNzOi5MVL7CqhToXUOlDa/xbdaWKb7e24YDR
RZhO7sFFrwHnkj37AKqSYC3seqjt8WjZxQhnszV63X7/mJ7qV6D6ZOci9eCEZRqJ
7Z/F+qH6y4UZydIHC8Hsgy5rRIhvbWkLhiB7xxVZGI6YYN+4ZjwecZo++pAx09Fb
yQOPdfTt/agezTcRavw6SaYh3yeajFPqVmc3RtiQSEXdLFmLGg1JZ51IXMSrKovG
x8D2x2E6Zk1UsJteJoUHEiHJhvhPMsVrj/+kyVHd+wKjgXK3+BsPo5uyOEAD5vTO
SQ9Io6wYSZww/+TQaxGvMN3dOyJ/15NEWow44hF1o51Fr01yWJwbgbKyOjsvXQMA
bN9hjeYH2KDYtPPXfPcl9n/9Ln0CJbPpeitUPWGKHMmC+XjkTvfbQ6xrrJU0hsXv
trx+A2Yv4ucM1fkbDyOO2oxiHyvWxYTueeQHkQp/JPb8iyTCqts4Ws1cmSfHZerf
8LBWeD1pRi7VXsgP7zodyPVTgdTo7xulJR4WvS6K9Z3zgoDhWnxVRhVitl1IVKJJ
eUZ08Es9aVGmgF7YxLVmRGWyyJmxSjF3394deneTNkU6c2eUv0M5Amm4zNrZzS+P
2fC67zUYFawFrrkye2ilqQVO/u5N+vaAwGeoO1SjEs7ku6sFkhIEFI43sIMWxKfk
Wvq14+cStA1yWm4LRdQASR84CDG1EVkwakDgimYNv09RxeTCGrALtFb3ivTy/Q7N
rYPGYSvrxrb+23mY/jPiiFrxWgnM2pVgR+hiDivtKpgoPts6F2mG4KtF4WrJXUYg
2KSuQNLyA1896+wH2wNG2Hb8YnUUiVRYCWOMWA+W0srytQH4ZdtMZc4e+QcCo4xI
2ScMQbO+475qIvEimYSSA35LfgI51dyb71fgyeiMguuLIe3vxhevr8oGmXR3Fl+E
BVN520e6wm2kwqrU9bPq+bpaU6XXyWE/9LgjY8Ta6RqfHZQuJz55SDBSZRvqq3hE
U93w5KaeD6yAwQH3RQyG0jec/Wt3tKmJfXrgv4TxoTj5Lj6M5X9jY36I/sevvNcN
NDIYuUwMH7EGtwilY4flUZuGOBfypWgXuUb6bHVeFXszCQwQPzfZE4rDZrLsSSaR
ArOrpclyN6mHtJCfrwWO+NAeL4IlGbmMWMWrtQDF9MUG9e88O75qB6JF2GCr+Pdr
9s3Uc/rP62QZVwNaFrKHztUyNFX2YULj6F1MUBMIC9OfX7kPlWawlTjXgKNVO1Ba
OGxXYCao48rtBbLgoEWoguOcIdaoX+DF47u2dIGOz81qr8wMsblg0WCUpKaw5Q98
IGrsSNgF04qfuVVj2JWvgZTg6MqvUVlJQNHuoxFjc9ui9MpogfWXnWDbcKP6HvHc
Duokl8x/UKiE757ywKq49ZAO5EQrYV2SQrpmLFPHxdiclcLZUUpO4lT23RISgKvk
n137vWi+zoH+buKclF9K3cKvadZ9apPXysmB75Ob7JYAIOG/M3CqVoRNmTzbQIMA
3sysaOQRnH+GiHeiWKI3sYOEOO+XAQbKa7Ll2QbKr3c0/+N1994mrpD2YLmdO08X
t/md0FAH69KSYTVLjeaE/0JlcSvYx0cirRGmzz/LBQPzxoLsjKm1VzDq25iZ0bYm
Xoixe2u4hX/t/HwHa1ZS1c4HEYr6SR6Ba8yd1SMdowzQ249y+oB8BzfLO/0z6pa1
5bwQn/PlXhJkm4hgOe5EYPpinI+Wo0bUpIMcrWYJw/jxkhpIWcQiqV0TDyQYAPMW
8rHPhjMZUPCwxdqks3hTbc5gIyrG7lO+8U6ltykvWBRjlo04oAqMLZj20au84GAr
RLLwOp50f0f5ug6VKCaqFIDO4RkkpNDdhvkDJi+TSzvkxPW5lyUtDNqXQhtWwLs9
4Rizf02WMGAT0WtO/m2ZjlrkkBQmEPl48ROdPxTZP+ZGvwjzj92UDWTnPofWZefJ
FQAPcdDriYay40QVqLBFa6jUnJeXkNaGlmLQy8eq/SYGubqRvRM7GTZQHB0Shf8q
YhAwGbonfOkMsURI6eu/GEb2O4aVsrJ1H1CSIq+Y75V/kFa+nN57zT6Sbzsw4FJV
E3iQFeLXpYvKYSMOF1t+CtgInkfhN/IeGOhmENgrAp0AMCdJn4Nj5uwAWmk/+/6v
FBGasAQ1D9x5urtpMf/T26gxrFQpZwZBqKa0iCMU79pKAgIbAQmvsI0gpEHnMX6u
HEDFM0KFrZFMciJP4ndjANAriEUPPweQBU2IvFBrCl/v6nSfUv3JqgIpO2wD9ldj
NUNJXJVWqqpgk8mnkJLOnB0P+cWyXVLrj1vnAK0nU8Xk9BEMQQnC2E0p+4VtfCfN
jVyhthD+QxTW6gcx6AWo8jmYGHG8i03Q6ZueFscL56mINfclCHw3GInBKJUmGvJM
H3yjLJZLC53T8kAqzU0egOF7mHfOEhW1VyKNo/xlS1KCdcPJuHFcI2XUwiIjCTJp
irYwdYJ0U5uKaKjIUUFISQWsnuRhFD/btH0nXDJtBbJbuBm+/TpMvpHhuHrns0hN
LtnAbiWj3IlA1pYFOuLED6w5jFNo7+gv+KM2OQUWcdh9n2ysoWvO03TzZoekGHoP
BkXT3PBvVndHrtKaO9h9D0FcLdCiw1cKTUzzGU1ZgeH/MmFe31w5NTwzWAA7x3VJ
CICjej/C19ezCSBYNdzjFW3mxrL2pzKR/gcutfxnz3nfXZw2xXS8l3Dv4HCLwHFe
ph2ICGirJxYBfEPDmgO/TuVkkRDUSbwoc6UbohKyQTxxCwimYqALLsHD1GJFhaqG
oAndSfLdtB13ueU4qaD0XkNCkpXLMDCGRzBzbkXj6q4X7CnWY3SptWoBMOpRIxDC
FmVr8DSdStoEzxNfTTOxT8CqV4Y6/YGySyehlPBSoQP3mAc3blcX6HjNqNyNohbe
YRRIPAPqyA/Y/b5xQvEy0slWIUaeT93sZKC3sCl2AwFBIjPWAeT1wpfMY9JQDmeZ
o+uQpF23JzhEfm/3+q6Hm5whbX4KwFQiNWA18hSH2YsNSxeSjF4csga+q5eGk1QM
rKbApKL9S1tFESygiCpQwXFdfCltCYGWGa95xCnfFEEfOpmJIkMVt90kz9bDXPJz
+WqBlE70ObcW8iS/WFzbHWMvZfOIucIcZUPdlLdatfe5D2D/Z9dS2L5JS4KKtO3O
NUn1QfXfBtcQvrBdShrpVg/lna8z8vadqjlyp8AbTvIN3cxM3OYiIYRgXNOLGI/6
Nev9d1zUeg0SMf5WMgmF/DyJYin+7z10sgP7MR1UYy6RRMmye0qJ1H5VoUt0aHrm
wlLeRA7tHJzEItrNIDNO4m1V819dsa5L5ZhS/pH0ucpBDw9hZn4sFT3c3LV6s51Q
Dp7t82zImGe0TMBsOLdAAIvq/ETR9vZKvBizP2G5ewT4VVku0pSvmO2C+GODM4AS
eavER6vqGxXDRa/PtdGSOzQAH34pJ7vvYyZtEJBBOgx2HncsgI5RAsCQY7ebhkTA
KQGRby9Ql7x9ekVX6zCDaHHLvr6sUtGeJEwx8vvuD3zrXqKj/ELPookKUcafbwUS
0uI78SjdMcxUg1Z3kFFLnWdaZ7HnDBmdOU6zTeESlNiQi2MeRdR00n4H62dTGqSU
HLVFqqbhI/NcGUU/5qC1a7wSQt5Rpv7CyDO9XO/RfmELpD0Go0bV5LvJfNq44lAp
OyqnzhEkFLjnHLLzcW6FAh45ywByZrMRiK8xEn5TT5ejHuoEW9gPH/Fu7ObfA/8+
8NeiBpVbq3+qeCErJCYOXRSuTPelFweTkgSxrtTt8Jr9h6ydNtenTBZOi94taxRD
L/WvoDT2feQ4wxFawvuiwOhWwDsgRIpy/ehIVO1H7QLxJmCTirKt9NBZqS71/3ew
/1k8e2meUF90qx5xMy0cloZQagYU96fjfz9ehkL8RhUFOeN4atg2vzltEdwvdQAj
nywm2GRMYOCm1/BObzIS/WFUyPHSDDGPMW1niWJAzQRWR9dTIkt8/viC10Zpky0l
9gHx1sTM4w4tzkq3Yze5EyLUmld4CRsT2jyrmza0XTc0ZR3qjQbdq8Pz5DNF6fJo
EFk81lOsiwFHk6huELKjrxMMl2TV4fYZleBMuuLHHzELh+4uLzJN9mPv9ixmqcoO
PX55yuesvl1bN0iKmJbMNfKX07vYhnvRhGDwmi2PSEf5xONfHfL+Fcjwt/AaOoQi
bwTvF4+7FKNno+/6+zKCELWvZXo2XCxReNvbRP1+74AmeM+z8qeOohm8UMqjsEt4
wTCz5oJM8STycNUJsHSYSlm4koJ8DaJ8eYBvae0kNPpBd0KgpF24NhhDFpta9MB7
jJDg7wRi/7eK3cgwZJ7ayCCV5AhaJ7X3YV7Qbi+Sj+H1i6N5/UUj+UL2caogPg9+
M9MKekUoqEoHMGGQhz7bEk75sOjeRxburUeHiya4lxgaQtVW+cZPWzQ5do1zv9A/
ROyU9gTW0UcMubV7wMWy072c/T/w2h2sq6LO8Qr0TGuyyJNGz4cAfAhLlbWWNPuI
gkXpYvLDvuz4f9nZiDH/8iBlQhCoSFdUz0YdjbqxTVyZMXySzlAjKXm3o9SVb8Lj
RJO6vm89mwjPuOtzCwFoMBAVp0reH9C+yqPRSBBBjLTr1x0TFsJACDlhPsZ6ah//
q7OO+dHrZysmF1JtKFfVngq/WaFrFAZ/X7hoqFrvuTtXUp6pjK4ZLwwdyjCmlIUx
2sFu65MJTp79X/UsPPQ/WEDhdRG9RZp8QXe6xf3sy4qO+CVe+ZVPrgk8ciJh7uXR
Jt0L6Z/pYT2UcyTyNArlGjUDR5J7lfBM1ztcdNg/GbWTDmgDCF5R76XPXyNJwMaq
JtMEjPT3ZB4EtG0ko2B2c+ps77H4WTkFCGxZovOXBB4R8Hmh69tYMfUi6l7XG+CY
0co3C79J7EvM+IOQOK+z/XPzg3GhjwQXHAj1xgbiCOxeIcAN2zY7JVFDwq/WZGUO
mOU1fZqxZpffjak5S8FQKjbC40SPED+h1+XVhoPDG474DwaVARin1aIyvSwRiWvy
+YIv9JWiPAXo5tOiddnVQgeK+T8smpfQVfuT5vOHVfHB+C6HpebOyNSavDM39nOH
kSvNgnWuzF6xm5KCfgBiimEHCadGKn3eavIFx3xppLlZu2N9cLRKRi54fZx5voiO
DKA9dKd9L9ODojkJ0tveRYPAeUnjtLmuzGMsuMGkJoC9Qj2uKLGHvQnlQhT2WlWk
n4/MOrCniIy0w/6sTJKTL88Xk24fhvglUF23zGVNxeMjdz+ADGRzTRN3wYRNxtwj
BsUSmR/kycQIRXyCbpQbGzFcVJKSFU7Ny7BGacdV8fRufgLispMnl2A71UdBYnWe
efYYjhpi/ZAdmOGkcMpZiFNPey8ocJtcIge33RZn/gMTDU9djD0EQfab2bHt8VYE
TdxPFyH2/3MkYhe5qzA053ZYFnDFFc2z9t3hOThr/YGj+72rdNN+JuBSRphqTw+s
UoCdoPpxeJEXxVwNwKtfG3Ez3UI2Hudj+EtuRFQ8Fjux1+tDOzfJ8TrQc16guCDe
QqDPa0mvfnoI4MumjGu6iig3D6ovXZtYBYmq2rF9J3Cj68pBKmlGxEhTAlwL/ZmF
ikI8xMcLZN+/FpgFrnfTZFL1JSut9EttV1PL8PSvVj5x63Z4gN/34XqdUI0KJ6y7
kOUBZ3ekpOpQFHs91lIMFmMGK3/esNaoz7ijK+QeGtrBk8V0GRcuhpIDS5hO+ApT
MlgXLZrdmyxn4AeK9dz3zZ4WIEaVnI8iFW4Oz6Z86FCAAwq+LI7sr9pcxMQFWtU0
fJJRL5fn8d/1q1vuZ4Yb84BaRsO9KWvmcwErG4TeqN5f+XZWH75BPJsLw23uAV8j
AUirYGhKuCN3YJELNbcRpfQozac4Z3R3c5bpHIwnRS+3xZOwjIRiGDer7IWyByxV
UvrNjAYWdDYkq4IkckBFZwSqlCMm9dD8sKE0HbY506mWQPz6SuHUuWTMA95FRRLk
dHeXAFeqB5q95f0ROydbQiHJRHqN0OolIb3aEGSY/OrqYgwRaY2kd3+7XsLVzwfK
IWvRdpfQ+yxYLriv1rwg1097xywbpNq58GZTY8501NE0Ft2W9d3ObirdYUq1t6TM
95ZiUHGDU7cMQRwkXEuM2re/2us+rSwJ+I3RZXk/yCsiBkGKM0NdaJIrLGCSeYOk
g/GNtzj/KZAd0UCy9fM5KIaOoH9K5Fo9zVBuW/uEgqaTxSCKcnJPvIIPI4gPgImV
IxlLGL/xs1G2sLU/nT930JqoTUh0IW4n4AGPtBD+vvccVuMrmGYVG7vzxaE/oS8G
ZLf/7L9SWBO8sqist0n+eQ05ssnMTESMWxhKax1ulB8ksaIqto5nj/iFT3fhL96k
SbMEIilggjICU1GN5g/AeLeHuqhyJ+TMiEuQJ/+PndHBZSewGFq/VcjLyt1TZQo7
O34h6GbIlCOG5EvIqVOuzfT3E8OfM88CLw90ID9ZB/1/i31RuoTEk+Is/z7901o1
FleClRkLLVJmvKk0eQYrD27b6/VtPd+2VvdyJzS+q3uPJ+mrUnTQzxvtpR/bHN26
VRCU3vgGtDlOVOlh4sqm5OZvkj4+C7w2zMsLBVtnDZMSX4EfbmivRcfJWdiPtKBB
Lg7BNkNgNpY+5r6vP281dPw+12C/s0uuBM2P2brk638AUFGC8tcvuxHpi2dEWO4C
TBTupXuMgNKPpqMqU1fC8JAPuWRRx0Jolh9HMBL7X4Vxb6+ywVwpEUb6k+ORh5Iv
HeILHeuNT7VOrn9RinkcEBEUI+UL3HUXo8XkFlGt4gyhacqQBHJdWIIXuj/a7z4t
3q4+4UP9Gols4W0gIa1otzPkWKtAzzwd8h5yBZgLapVWumE3091ZBMam/PEIpgo/
r8JUO22IqF5UujzrHkmFgln7EAhXo6MIsymRVrxfehqTamRaPTt0VDxDTOYMiwMg
qpTgwSeOlJVtLtDbDha2+k2a1q9OINGP43k4YGuTeOlIY/7KRrmbq3HRwll94hrK
X/GHJxOTncgSG6uDx814wFbvuDWRses5DE+FUSX9kv2THdLB+iCmqgTLeMLCqol2
6zd34AGelAD0E/aNWEDKvVQhCCuP13iTBouDZs9X5zfYpdETnsgo174t7pPBjNr+
dMk9UPEbCpR0zv2tNXYRet7hm25AByJKU7PzZ+5O8er0dJ5etvgkXMTcjHY59nNr
y/Bb2YifZTUusQ8t/AC432bJAm/WWdeKjEI96lUSDE0tlXeo/nE9dya0phf03Eo9
AxmC7pLwJc8Py7v/H3/LbFK6xYCgEUpk6NoQ/Tg64Ic748Tihzj4uhqlSfKSa++n
Qy3u++78tAOGvgteMRtYPCmYmvQYroDbfE0zwpZ1yQ5RKCrPcMHNVixI7nansHh6
Z9EZjtXVMB3TZGkRmxq6CNcgoNSb/o1Si/yg7knoHk1eqbPB8b/MIuXsFy4YJdFd
oyY7ZbCmYI1df1SavD8XpFlXuQe/a4+FLwhNUZId8tb/Zg+cMQvPDi4VHMi6P3Hs
ooJzE+D8YkWJ6B7KGt4pFeFk3iCifDmhwRTvM0QdufuVXqKzocLBOm3MaSU4xMks
k3yq/ax6ti0ozXWgDjumLEM+Ul5eDp+jb8ZAOrobHlo9h3ZIvqYrA8oN0I/wiPZG
ZV2/KCs9XbYrqJbxWCP2M4lp+Mw12fmO8R7C0JKzQ1xk3v64bX2pqwtSM59lvhep
hObqB+hQ2UUEatY6cB/EynXTe+eFI0+fIgABR2/3OVZc/gjIU6eVNL45cnfyANsL
LAWxcOE6TKJr2g69Euv6X1LEnKoZsHKOTvVqgPz/5u7OpD47PEJpqjeRmpm9vXBq
5ADVcRKTrhq50lFaiXTQKpUNeqwD9quZo9eVOcUwCpNe7+Zi1YXUw9FFR8zhUFcr
QTtt9F1KzYkjmlkm/h6shpGMvwZY/sgwwD/I2EhnRuIy8+sIXKR7EBm7FE8juHUd
8CtWCCrl65cYL9HKBGnsbH2ogKtRhr/Elz43g+BcQ3pr/prbxF63qx2F5pHX0zK9
WPc6CNlwEwG2/S/YOuOket4nhJRt9O7L3mXK4le4Sn3irVlp/598PBXX9Lqx7XSl
OREAMwnAhdh/PDyUWHcUOrt1BCPzvPWfd1vEMSOPems6UMVF0mKsWAArq1a8Had8
eG1naoS7sT/2VS5uhbWbUNBE7eC9InivES/PH4h/XA7QFRvpISNr9GsDUWbjPTB4
FXIYAA+CJzwFDmEHYMckprRmAxA5YIBwxpiKG9kZISAlwjQXsvS2xE57FjdWqbVx
lIT+CQHu/UcwSOBEcwOxl2ga42xgidxl6uXcTNIwmlK9PRZCd1xq62AhiS6zSZ9C
aKnNlw9/+ecVNmCej8Yfe3OKJIOWkVAlqvu2Cv7e5g21HfNGLqtUUDrOJWMYeyxb
L4oKGK5nBVHveMJJpfOZq0kN9gvGSD0izSRFh3j+PWJ3hyaaWByKmK0FFq56CwUq
STXhbC7Zti4fCjWdKqY8u95IkKfmOPFsn4KiMMUS2GLj0Ie11gVK24E6Y4N7K3HL
WguB2VcbFQhfG3NSyN3uLp2PWQxYztbQ1aIyt11Oa/kEkCNVo1QGFEmRhtRdwRNa
a1uG+IEgzyY6QRS5MhO6nT2b/HAnbN7tEHnbdWSR4cSj4GClnQrc+oEO4Qd5HYjo
MjGpw/dweLdPBVcBHNOyK1MVOgPSK6MWt6gXYFk/LOfznAvfw6lq014iYldGe/h6
WKlMlKAT6sqV1mCfI542QRDpHBdgSaTGMlDJHMkccytZoZSfkf2k2IU5mdGR2olW
BeyHG9uv2a7XIBYyPf0v3N+xkQueAV/97Ik4gwr/aH9XhJchcN+9k+tljgiEkBL3
iAUX2QCApH99EVXelHwv1ZO4pkbmP4JQzrYyhvPmW46Fe0Xu1G0kIaTKH0igbKLG
lB+o077D/lQ8/rdycgvWWL5OVJk7lgkWNvuQevknouAvbwYBlAlEFVw5OPYsAYF6
aqld5qC6mppaSzVI9O+G5FccTx9dGrXAp7jI+0Hd0DzawQ421TJk+MFQ30kAFOB8
ty6uISNtRJ1OnuzRE7/gXCezD0f8pyfg3jIgIDT8K1NoiQ0rOHSGXO1E+QeETwUy
UNaubmrEjCRv5j6MIDrX8IgHXMlwkK5JmzPs8FVJG25o2cYuBZujfg96y6Hw3AS8
WueXPuNTz8MDC5kb3XKCr8c8HqevVHuloVp4VZ2qeoElrC8uwV4cLQKzPKmlK0AI
kxOMLiRaLuxx2gtE9vnrBCmR/GzztB8iSd0nwMR8XW2xqY+pwm7zZaYJJRxyAtuS
puzXH2iH1MTemAK6eUbLFeh+kJt41fg9z22POCsYZfjdlm/ZGh9ug36PgUrwW6kD
c8TmDOVx55pnjoqWP16qZCU/l1X79CuU3We/7Vm9R/9+2beSuW7cLe0nlTX/xkhN
A9yqkdyb+XCeAPj6U3XNkMvL944DDaPlMURFTkBzlPbkWRZejEOuFR7Q8ZC0REEg
eqhhFsM+VfQcZZu6GtELf45l8k8Mt08SmFEk+cdgnz5KkDt3pxvmBxLGNX6hzOal
B+5sgP3CSCQkf4qdHfKnYHLKFUg9KfmAfxReZbS35r4xUS3rYG42MRtJnWoCHoh6
uhhrktO3FgShHdNlE4yAf/YXDwflFdomE5Ic8BeJ4GcWKnP6jL3GAIMJdepOTEEb
4wVPXsR5e8dT6yh1zzapon8KdTrscoqtJrxMinZNvq5ZW9meplTdhPgfIQOfuDm3
q/71Kla6NaMpcQkNVkwsNVmZ+tThNowWkT99NIqfgooYaEIZpVSLDFNIxKTt24y8
yEGzmw2cKflm2jY+LgL26Ga2dmC9ckjUFbL+XpUCpZ3Oh0PPojAlfE/jn8z53+BZ
p3q9cH9YteYI635LlY0wJ3Z7+Jj58wJllm4NBgkAQju3myiNiTpPhJGLwwhNEBo6
ZEDvlyNzHjgxBB5UwwmQ5dj9idij4rEhRERDk/146XAaWE7UclcAmm5RrdXKEiLW
zi9+9ddmjQ9FNNID/iFvp2cFj2lDDopQeP490DlfB1VENAzDcxEEqYsSQ6Koomvp
ZW4I2ie/XKFL1onqDHgJeMUILMVsKR6UhLvBwPrrAe6gSFSR39bwzpD8TsNnNpzz
XtgWpzvOYgr5t0lCIrZ8hJRxDdzWhezwVjkQ7lS5mqEOZTUBPq80Vrp8MZCHplbT
eq3w+0JcQ1nepsP2aWUvaB4R9cQVlSxcgu6zT+0rl5r1avkbdkOx8l2ux3Nwo/xL
TDt3UsnhCPe6hz7mjJ1HCedZj3VErFG+3CZfUaWYc3DFsiSI+ywjFGz854K/21wE
53f2logitKO6RNzDfTEEpyl+Ytx7DKsX3xWyS7X0zLtPb1ygO7UTfroPYsQ5Ygdd
vmOxlhZCRd2ITlwQ+bvAmj9QMvnIwTIhMTfnRPekK7NVw0qMcc+Gj0SsXw+RN5KO
iG2igvNCT/OHYMqlwjvyDrX0CoEhq6S6Yh0LnZ4xzUq6rifOEZ5lEzDgT83opNjX
OVBRTcD3ql1ookfRLw4zLq1vTKwqYI3Jo3K09Xt/2W7OcxJcZ5U6ITXdY4lGZStv
vpClCCZxfiSJCUYwgAZB1doOCDOhDsynrvJQVERKfCMKTOGlpjkT68CE0zzOP/si
l6ozoM/K4bYifJHHpexPRB51aDkdVynxEbFDwIGAZ4PuV7sU2+jMzcjwYYJK21AG
jxsY4/PINRR4Vbb8I2maSjJGkwF8UtRAMZTBHDM6DpuuCz4Et+wvo9dJVt2MpAl3
foVBEegLKS/+DNudTucSdVNDG3ERWGkaVmxtaV+Zh4M97IEoyMqNTfrJiR2d1Rto
mpSrrlTV2vEXlyIAyD5hT1gXVTAsTGVXkjqrRuCPPz71sAeMcAl7CB2TGIl3xVEG
gBbM1py4ZRWmuvhVmvYjWiEi6kDao6dwQyx+lFfZ1SId5TRkus2lkf60Khv41pUF
ShMpVDYT1CwSuGr+GR3Q6fpfiFPSGg0GQ90UTeoETx7xy/S3uRGIHZ9aiMTmSx4S
M2sVYE6e6QJ3ueU/NyDx0Ze5x2IkfpcKM65y2Y2wASH24ia5xdCzLxr2tr+OWE0C
uUB5qP/eQXBrkxyUYdZ11pcu/wswH7uWzDNlS0A4/Oe77a+ouQ9xlkT1ZxTwDoKl
aCjv5g1ug2TKIaEvfB6Dw26VlaALB8JT6fA7VDENXbLXD4tZQSxNaiuzKEr25hwy
LTtjsltC3gEKhZwjFTWcCYUiwhY24iBlE7nQjjoUdojIoVqXvS1AKCZcGWSFdk9K
yu9gy1fUnz3HKsTxsT9Ee8G9i7uQ3iymD2zueL6SAIZmqVskGqOvYU0SZy5CMDM4
ZEvq4PSatolMojVDHJfl7acz1m0FQxolWk5kiZTnF68i6GV7kkmvtLQUdDa8wANM
b2Fz2KxJ33ltF54ry+AU+teMDIdk55EtKvICl/9JoShrVSKEABbdngCNuQpozyRv
SCNZ0YrSBUB78iwPWhbwpV6sx657a/uXKXwY1UrNKSVRor05Y3wvKq7wyR6q6Iwg
R0ao+P+f5Nfeh0ydjEg3Tab6pMQBtHTo5bfGk5iukrUZMa3JtUaqxBwx8Ptqe0Af
7n9Vd0lv/T6RK8uUSc6TEGtG55ct0KOWIuqItpHwdamLd19mddrhb+ezXlELVyHq
L3zhWuTnHA6xNTRkYJXUUaK4KlABBmqKLsyoMS1eEEavugICiCjTLXCF6mVd8Auw
vuCzV3vwYn+zZmUV32CS6jVpaT//wFU2Cebvi18G7v7gNgOgoWZN99qNSSdJP0/C
Ttaty2vXuDvHfd9yEPUu5M8F5H4LZZOOTcoGpvSqjQ3Uq32dYKXQ9QQYMs22D0uz
gnf628RYMZlhamVj1HXEaPGy4gSb4h3ClsEVhioTtvtp2Ks3DkQS/EUKtB/gMn/m
oL2t9ujorL8JW9NRy0PZjLZM5l/2bxGI+poyScSc2liOzoXRBwzcoLchITB1qOPx
ac5AEJkqHayDAiGLCUCKpEXNaYPeEHc6xEG2NaXvBKwayDQT2J9hCoKa4Ga4hG0t
yLURngKEOIwgRa+jsO+jf+oDl8P9KOYdop+eYWOio8U1huENRx5Ref9WihxRirpO
f4qB6s3QUkQcWGoX6gpVz79jCkPzqeJb82i9U9BnFl0DyLK66ufZmHGhVl+Kkb/s
/xf1XSuCEI8Uan6HV5kvAwPUew/X0Dyw8ZN6sJwbKlZzOFN5p2f1UjbYP3PVEixv
Jph54VtGFCy7fQZASGp8iBAxfXjsPzr93VIWbCvwrUuV91raIribnc9JKQdKTT4P
DaMZBhNnPClrJS3W1b5dIOnK/vcaPBz+zEDPYMoaaYgZeLzecY4wfH6Cb74jxiw2
IUXBPw92GMpwTHM9CPdPs54UIP60i5pcnyQKz3+JHMB+bOnoJYgiOWrPl9dySznh
4u1C/H5WUZWl52eNNvxeCr4Ie1v/98dUYPhdJXoulW9LSfyLaOFKze+TpLY+gh41
KWjzkjmycF1jXB6gv1tWTWBIUoP0Vng/MOMni2ABGc3QkjS9SKp/sHXF0ruahp5l
NwXurZIzFdzj6BNFhj4riPm84SEb6A9JED1PWM0u0+LeNJLEYXrhF0Yg/ZBw/mms
m1vcUof7ELy+kMcvwT8/h4QQ5+34qluLquTJ1mqWKZk2nQBtp8Z/0ba98a6Eu3vF
36e0qTSGEjxaAt6gc8MaEbPN0d+fS+lJcpOAbDPZ6ozfVG78DrPtB0NcVi6wv+B+
f/QKdKs6p/Eb/3rxZ35n493JUJT0ARkDZt5HWpwKOmCVdXjiMZYmLMI7hbNgrgmo
E4u0zzCfns3Qqae61yF/rNl4NNYmh++5p3XOK2E+J2uGoYnR1DoYMI5mryxnerUB
42XjVo5ksRlQLl4M6uADTk1j5D6PS1sZmL2sCbjuaahNrVabQvEKdTK6NJ91bIS2
+BZcN3Dev0xZgmto0Xm9tRJP5fv1bNKKA7QIpi/MgpmIuJBMZHHyezQfwFD0fvgN
N8+EAdJmGq6wHdH1L1dh8p+CNR7GDSl2BUA79I8ZGYacpG0UMYGKWcH6hYycxgx/
j2/wX23/cAMwqBMhr7RX5JFDvWS0LwVrxBW9Y83fLiBe4dblqIXfd47f8uhBelpS
UdTBeVxi/8COBaTCGK4YSohBnbUKfwF3MODuo0W3KNVSxVJhObzGtZDp98h6mbc8
uo9Afykz/3CRtdmgXwQ9qyRV5viK7NDuSfNd62ki2YCEb+RwBO33d5G83m/MG0Ho
2WJ089ndkD4iCowh+Rj5aAwlhMMrdnr3xTa0N9Vs9mI3SPiuy3kaxAXnOarS+O7k
Kw9fZPyYTqgrDenWmJa6wELvpxr8hSv8L9DaYDgiEemxpAZMcrSjhnsFQFyNc9DB
rNVpaq9G2+ARPdlaRhq0xnkp3IwqSmqCmEBAF07nlUQGuEX71uwAxfj6L5qvoBwY
5fBfAzN/m9kv2G5mFO4RsFRV+9Wmau/ZIz3r2hutVEwEmr9rypd4khk2TjgKOfvO
GbqQI+ENeYqF+WHwi6Qoa7UorpP48o/KM5ct1g9Lxe/Zlz7Y0n0xe0n8V2Oc3meZ
tpZcoitY5YJKkICD71sk/FTiwsIYwQT0y5Nnh0aoHjH2+6GrsbvdMbOkMTRGWp/p
tRKLP/iQ9NJ8yrGrw8DPOhgieUCNOXoDvLX7azMuaT7BAVQeJeNxPRBCCTG+iHHi
Ax8Ai0bcJNqKyfWfux/1lfXxJ2+HAulIDX2MJ8WOXx85KMROnsbxZrZgsB60xHfs
3J4XSBWCDmBxNS2XZ6u67w7WJwW8kd87UDWMEFHfQGGRmvcUHUXSDnqZJyZXl3CX
WZB1UmwWcM8Fii4WnwEW/MRp5pUTqBFQvgOdma2sLNoV+3ScyvQBEcRZmPQb0cKy
N13xGX/pceOcxm6pK6St68rOOf+WCQrNdIZc6zVcmy6WNZ6e5pwl1fZNLKFJbVpX
7UZJcPe1zXmPZy4R/fKbZU1vZ1FpQRd3/Wh+jI7ixNA3lOav8/4yuN3nP5LOfpD+
7NPIs8ASJUUulGJTBrVYke5c5F9g7AGuyr54OhQfnygoQDwqPDMXuWhecc15arrf
CrQq9qh1LBMW2bK6ZFKUn5gaq6w3LMpX4GF22GkGmqVg61HcdqhFf+r/cpevNJlp
ksQrKtxkWRFnfaYZUzOz427a2IF4oWR7/lZUAuUhPDONUyqE9MGCw3u/jdWM/GfA
3FtPDNyczM3ndGhlFk3cL2noNRB128egyOFx5Vyfdm43UeKmWhT/B4fWHaWMRlNV
UPdLDVC+IzpAIFff4vbtu+MuYJ4/o8edWyVwMw0OzrktW1+QlzgxkNcv1s6tMBfp
/RvM7D20Dc0oLgBD1rIYdrzs00i18TH6gA4uprQw97YCHw6wTvv/gu+9L2IPik9M
gV/EIuqDL1fQwfukovpO4ORhhFwADWxwoyEaEEMfJVIx/bIO5oBjBp7QjXwWLg31
uqtdc1rnRqINgeRP/3qENlJQL3/MTwCAwdabl7I59y0zHkMIz+bZ77oW6IB/i7qG
F/ezgWcLuMxw1KKhBZnJdVgiYUKhMu1lsXUd8+/JbkUwys60hR03ogoWHOBC7wdX
gVLvIlIxr/x2x3xK/cmybL8Ehq4nGJBZaPi8CtNmsp3m+aj/Yf13dCIZqHnQc6OX
BAIdfDGCW5VqksjtfR6VOOyAE/UgL9zjO/DlC5ugDOdFU38lI/SZuy07Z/it7/Y/
opicEDNXYHedwbAXNLY02nha8WmYxVAfjEmwYO9xKANadGUo9wKSS6MKrOV0irBK
fSNo+d0GZqTrIXdog287fqO/l/AJCUbR5w7bkkVvCRrzMUXOJ4DI7fLKpkY5R9aN
U4hbFquQv6EuJRcgOHVLWoScqJeKA2W5HTGy1esx4e86QMu48WulUQn12jyghvQ2
FBCWb2gkIHqyH/SPNU0tFQqp+Me3c3vwokHqZAc1rWQSCkcEydvfglcYsY34EYlb
6V5/ETWgFqH2fKa6ilQvR/nIiDXscXxJlUr438WZsfhgJxq44x4OugWcNSu/SWji
RCsBYtU7RHjg0K9XNNEYYGl/6FGBsPO5xGYPZwNb7iqX1YpInomdxkXu5ypPVpuu
WJFC7cp6mFTJPbCmg7ZU3wXvtMGZazZFDhGLrpqDzf1OJSdYTOV4OZMb6e/oJSgI
Eaj+65DQhwOZRbtJqwL5sr7X2uoN1yDa26AFpJkL1RFoEYgohRxgYRiu7ZB28Rjn
QKysv1MpBusG3TcngyTpQYP6O3o+d1stkiTgaAep/o+fUEyOJMqDSDTwUY5CjuH3
Pww3DuRPZo/00JO++FElFWiS14XNfKcJZEsyNQ17b3kKoJ+vLT75yzOZwqe3lbQY
CM6ER0gglp0MSqwTlWlRLmaufhk7VDsSvvwpV7Z6P2BRwkp2FqKBgQsBTB2i0euJ
nOj9r6/JewoTnfE3PR0vvYX/iL+D2D1+cvPPtqrywyd85QbWR4vtXwAr+sV9+upG
kInZBF78y5GEnaxofaJGYlw4pTVXeKHgM/7MTkx7mxqoPB60qEAvCdmzPePH2o+t
hmvXF1r4KuM//AgX4KihXG6fU0t9LBi7i8MJzbDBEOHsQ/fgLihjgWYKTpMoTMvW
dNGjAJbA5SegRmurLm6mS0ESZr96uxoB2XuCiNzWxugN/JAWxK3RTwe2f5DYe5NU
ZEI3RNtfz3yhTL85IYYWa9wV89RJJx5oOCuzms3R1G/DAEZR2La9DgESsdBox5Z2
QznPkTD+0NZepWmsJ9eMY5XXX26lVtipU+qH+gN1rMjsPYD9GiE16J7U6Fik24QC
uRZeVmdnDmRU2uaVr/Yl+aCFrQaKctUrEGOBXX7hbtkteTVhroEzvZ2895r4rhm9
qtG5LTe+BsphcndWPel0aTnzYpU1MQh8kxFgeMfSxZxkcU6PL3UEEKBpV54eAeZg
aycdyA/pimQCXfdMwLwVVQSUEQIfEJnP8oUCTYYl7vr2dOtbRHbgq4xm9l+wsHND
qfAZHxRBtvKSTH7x0/SnNHPFTQENcaQEuAW4Zeffj5yEOvwj1xmzlwaV4s9mvZx4
ESygWZzTBHX/5Fu4sJixC4kT9XIcOmWZcTQC5mLnXCAaUxpVIOu8lGpNBG48Q6gs
xAu4rulGjSFDhbKHpGJvhqIrsBclJ3R5i+vK1Gtirk5xiycZl8KlVr4zWskfCYAf
nRqEZ/Vg8MHtX70xyG8Dyim+exWeHYIEs8CuFUiEZ6NHyg21/dg6XPG0n1jxL7v1
+9JseOr7P4/XkgZRJyasWKOYOZWcdBMmwnqk0upQMslYwSv/KxdImv8xwg83hw3Q
vNcU31lc444TVAC2OlsYuu43Lg5ue0bfZXvvvPr/8q25K1rj9P5voCr8/TBNxXGy
SaSu2MMaxbQqF0mGe/TrOaBIlrjwBXOXnc3hSqq6rJyDE1fk6llZDcOm5neOOtQA
8ZInk9YV+mQeH85FrIiDNC2CBYNXkyr55XOd2TCssQHcpTpZQcPNdmQS8YRGiDGr
1nzeclsuMstJI7uMg7Gb0/rYTAu9HtOhKU2+TwCSQE/q60o3TmORpBTNpsBpG605
WGwIsV9wZXLfW5pcUrf7/ADDHQF+bH7JeVx7M6V0+PNv/z9yyBLpUYr+eqrr+pX9
7e3+ni7v/xd8pG6Ckp2XHEzkevypr8UouXTn/pbnAgJ43XNh0vHVefzmPjiO76Is
eUrKGfd1zYAotZ3oLpYJj7knSJxriBy1gUFIYLKKoQGjJL4nl7tfNvMQ54fzkHmk
xUu2AgeaM3ESNh8doNl1Qtf2qO7MTt5hOdvfTXyanznDbKyTzJ4P/6z5HUoH2Xfy
s/JrEv65sZ4t5HYoQrZb17LK7E1Gz421IbnOaRU0BpIhKhNLZ1oeD/dy3uru8VvC
Eo9FWLXcKfd4bqPAXA5FyA6TEjyoCCUMkKLFuPiPsj25k5Lf7Af4wSp3RUuOD3b6
pS7nPZqiTiIckDobBC0IBBrLPgiBZI6eBmjrGpCpGXUsJv+TJgDibL1anuOg6nkw
8PKC/C+zB0EXdBGnEy4uns13AP8p0KfsP8Is+lPxPNX+XHfWt83WcFLi4Vy2BWkq
3poCs/Bu/+1xM+f5NOpq/U6V7nKBnX9jnoc+cbvU54EPy6l0Wscf6W1+Xw6TKV2s
wua1t/H4wcy9qptbgFtx+HleqVQ6nLPLTb+/LTQHL5vEASS+PShQe5DbUl5bEWNW
+1Aw9NyfbceUTJ+1YKpMwO01Qem0kTO0Bu0f8pts4eKjsyq49WpDx0iePwrTCwYx
YpT6HUdyatLYag9hVZMtt04KTKZRVtF6V0cx9WrHD0bhRJHRGbSzicnnh+hiCsxb
oituHWl2svcJNVslxZM7ssPfSRiA1RbTT4znBw9VBATX40QKOaYUhzm/XvH5+kf/
EsiT40vsedjKtYEhhRmSIRvCTKgtsSqvqAu3KTyShmshpoFiBaQBuCadRcvLnXTn
qDeDn1ifYqAZ96evH1i73uBnUrf2DTJvE4mWJf8jtZMYdsUaiyHukBI/QhWWQhs2
MHOBa6jre8BmPLqpDY57W6HEuUMiXkkJcE/yauk1EqdKWLsuqIG4Zpj4B+ktGikk
+pZ8Dt/QdmBKy+shYqGyzWCNYK/rP0MOxp3rwDvCMNbHA5kg8VmrNIC4+s9Gd+dJ
7Xz7VOoXnKg8GSftQLNolswqX1Lo0jcfUoexumL/3+i94w6y2po4PCktOZBB9Emn
CPpAH6LsgL3l+8XaXy6IgWXnxpWp6PNScnKbyLy5wAQW4HKYCedXuhZW/mz7/q8U
fOZk38K7Iq3jkgDAnss0OQFiN5SCZAXyR8Lxm7PLya5ENGDD3yduAdmc0t1On3hF
h/yF/m8vt6kzEEN6+UzPZLxkdpSietifujO+rdZjNgwzI0OBrsneaRq2b0eOlLzS
V0ZuLu8i5M8hM7fuSSRAgiN4/L8BmpUV5U+Ez20W06yRIH3SaGkudTKs6kZ8HDMc
sAebQdUdLvomqxxSyCVJDY5Vqfuyyg3R+pwZeJvzGwO9kv2vU4pOgohoQxxiBo6I
ZatHyw6FyDKAK6upkKTi7ZL1zdE9yvxHUw9L+5OvM9G28uFQz73hq3UTd5WKT4cz
jIv2mPLS6akSd1EzGyzU8RU0Tq+CoiLEfIBDL7JsTQpcUSDt9hjFOdBiVhvmVtAx
qbZveWTLu+2wJfSUG4mTrTEg/uPa7IOoJNtkO/Or1ykSza6VNh3bmSzvyTxYU4Vw
AFF30IdxRPD5xZWak2xYJo5ZVHVoK1U71crd2Hz2THMopG7bvnqc/JWiHamhM/s5
U+vXVffnYShhzK89LFDtXijtPAi/56OExg4UAMLUnYFgqHNhZDmAddBMrkyAl6io
LSF6P4HQRSnms0j0J5tB6UmxqhAnkK43pNvrntnLQqjQUeEX3BwFr2w8XRoDKeVr
kShxwx279G8fSEwgwfaplZc3RUAlEcDq7EXIGwB/5F6Aq62e25AoBfsCZLXFMF0s
Q8o6In7GKet3rNDCNELb0PpCbBX6g4KMHTYnFNtWv07V5MsNKMbgDHZxvEm+hcWX
Nspdknm6IEmL0Uy9zgg8BNS/2HAk6DsaLY0ytoxMb+gTfldts7wXozDonz0CwOLo
5m9EQG7KY+3iV6GliMV+8DLx8ADi5DcZvWd0hCt/mwKuUYuhzFN+VJtTFNlB348H
gcrpOphLKl7a2ZvEkc93j2ry53Q2ZT9sLQS3kOgM3JmR5qyICpW5gUawz9UQKsWh
JJ3zaeI+slTXEQo8JBomMLghgWfo0hbJkTVn/6Ac/fg/9YzECAAHd6IiqdOoHkgm
VRXXmpFzB14zCpQjtUJUBwmsYh4KkKk7cjEJvABtXOpnMKiudO5IdYCrx3LwAVoy
5bveyIr23xsPQfC1z4ZVVisEI1OvlKOow9Obf1RyE8pKeac0DSDDDCl9jHHbf7x6
yu/HXCq4SCtFRF/J6gcCEfPxgJkCC0RpPa+fC9uLxjS6QRMAddu77howaKDoj3DA
1WuAXDehdWzkJZLmLDlTrSkpaTgfIVA6ttC1Sv3eP5VWOUZHRpc1BSFZx3O9idct
KiIBT2vK9JZC7CbR5z5t2Fm+pFMoahEd6Q0zrn/3kUEwiVHgsD960zmmJrjL61sQ
idMCWu3FLb9X0z9qb2WKuwfoL7At0YWut7U+XWMNFNgVKmps6U4loSVB7gE8/Mww
hYw0J9IW+gIY//16BbWPQx8h/9HVBRolss/5mNAeARL4lxkHtBiGcd5ZkL0HBIWR
GMIunyoAjA8qjdKk+TNl8xsKyP7FJKX6TOkPnBGaAG+FkBrpZATb4De/rgTUSo/j
VW6iFWxVaZdLWAtTBNGq9BHh6Ggr3gsHQf0ZjhtXio0chWWU5EDYVo2X1VWABDFU
/WepL+HTS4noyRDr9bo/gMv+VT7QNWkEusg+13gJ6dhPCZ1tHAmx/xRUkDNcwSeC
loKlttcsrOM6RVMIOIGcR9Ay8CGVbhPwAm/VAGXiRCkMFqyG1jv4+QiYgDVroemB
1k5EIyzc9GNxZEDphKurIjYzKOJGgB7WCc/VpnV+WKPNgZJitlijxFeO0pGqcEXp
+yweQ0Qit0Nhfb1N4xC7lpNCd/9YxARuR5iQ+EUq0qz2tHe8wj87fxibhgdAXxTT
246Or1+aDFr5jsF2EKT3Bg9EKcP/UaZ2iYtpjEyFInaGJqvvgousRedZS1F3f/8f
tmXvbj2fitQ+khrqEYbW6SNM0t/OIUwc0TM9s5Cb96xPQ3Zmq6mqD2NGSubFRGU9
5ehEMBG6MHYev10FT2jKU6q1ZSWP4BjP7Eh4xkXzDaU8DbeZx39xaEvDte3qxxCK
CY5gxM17X5OLEilwmbHAMu5Wl30AOftnw4swubatsJXcdBPVGYOyrSe+mKPI9BZZ
sOJwLF0pdGoJzhszlaEn5AemR6o62w/D/gFpQNjz3D5qGu+262LKisoREXyJnw68
CmeWnBhvQdUTuETM5CBazfrfJTG8ACmHlEyrlHpUXYjeyBZMd1mWaCJQMUoDwU8H
dNAJmjE2maLNF9JxRgVl0HVr5jdP6uPsN5ka1g1Sq9yeIbbihAkbJ6s+8BKRPWc4
1r5gqZYl1psu/PRQA1TvkFe8tR7PuVUeSS6/pIzXLStUO+xg/FeYybQOb1XnkLCX
znXZHD4ePwWSVbqCeQAI46SnxCA8Hc4ULawlFo7heTpcwdQnC1Ltrx+gldtSSmn6
zyKQDMxY1QGKCQn/1ulOT2oalbH01uSmWa1HpFK6rebPrQIOZa4b6Re629UKZ5vT
ni2w9QGKtCemw+4HZhF4GT8ustj00GkNj2H7/lZJJtVXwcFWr0G4NygF4d9JBOyY
dpvzdulfIiqdLzZgC0yzbyrNB212VduGDIN7NfBgWVNXdrgXwRSZTnZtZnSTrVzC
0G2pTUk24TJmZRMFy21ufFPkvs4AKchOwZuB3q8/Hrlj6U8sB5Qfva6MlGEy/SOY
XjC2tiWMA6Q7j+qREww7IH9wC8csmKleR09IpfEGyWwpHCuGIY0/4uD7Axs5a0wX
fC7Kj/djQClmXwKd0qaGZxa6+615gNVB+dpsyyA4kqjzPHOn3al6DKiuayftsjJt
FscI0J72Tf9cSBXDs+0AjYPJUA8IRsuTp3uxpWnmobffqTB56gQmwwdZpWVqEe0Z
aFblNNIoFLH1IMLGhmm1KW2CyOoVaaeYVC1llPet/7sU84Xczer6YV+/cI2eSre5
hWxbVsOVNYm4GSGDkQ6MWfspFtDdN6yaPxDc5vhKqQpjuyGftJf+AeG4cufNoswo
hqv0HF63i2YyEQGWOxMLpi19tH3CxRKdtv//H8502B2jWlptDhj65YJjzqlPlymR
XZWnoMtpOBagEjw2xkBylTc5SQux8tOqOrpCrrYhB4w4cecRf6GXWDY/tQpECDaf
ozQC+7PWMWEdtkV/Ficv+02nFY3ipROzfrvra8aXOw9Xkbl4GuyfGcEcJXrvZomM
o//5L+TVpBkhrDzY+V78/TjIY1jKpAqcTfF7+qMvxtkDc4WOC2wB5K/qB6ZYl33n
4JMb5GfPLKRKa2tnkQ5VB+sSwvziyOEUXxi8zalAm1kL70OeQBpBl9Bo5+i2hfjE
ibcWJCNj5QJY0Ak836hpBb70VLzEFjZSC+g6JGDjie81jmukT9Q5ktRflQGrLyIO
nw7hVVH0Jl1xJC5HrdcSDtnP1d0k+8clcPTjktdUCpNR8igDQdhRNEKP6dRzZuMt
sZ8yHyRCWP02B+cW+W1HCi6EmdQt27OBT+KRod9LE07NYJim0d4AOQZ4GCIo3h9e
8xuSwL2lN1I4rBJrP6GBr267jewQ5Dy3/gpEsyGePmjWL9XW7zY8b+R+R+SuYD+A
/tGRl+LP+z29hDx7fb0FKTIMEi/NLDdhdxFGqkpzpIMCW5qq6kt1ub+53Zea29OM
4Av4IUOwucm0vBe/nfvMZqLZ5DqXab46O5l1vvvmUeoDL7n0yKFQU6aISQhbd9eO
lyLb0WxxWO98wD5Xtu6Sg6j3WKlkhAqZgoRt2PIfVO5IOh8vjWtNFxHzIngD3Rme
PHYcLn36OEi6dOaHLvtDn1RWT+6tO7oHX3AbzLzKFjr2UNErx2rqCFDqP/n5bO7X
EtyidM26DpfPzU6iBOpx6n3C/+8WoaXPvmoXEyeWwnQb9/WGxR0J2nL6T7JR5K9B
O30FzYXuUTG30BFQE4B+JSeDDnEjQ9XGqUwLVLMwG0Z7ui1uNJfpo2b9l9JHrdB1
FIOOeEcga2nNPmONVhBK35pRvNt9QN0cZlroPVjugsOUh3aq/jzI3nrj0OgTc/wx
+aW+sNjY0P7WpuXDFoWVzNFKN/9On90N4wQSx46dBKNBSfgnOthw+/n7sCNCHAB7
JnnxZxph1IOdqc+l9MOg8ZJ0z3DgwZ7tHNALqHtcKhx4xiwfFGGYfC9srCSqhJ4f
s9y/mHqckrHfXu1+OBAZmxSZP8L2sgEJnG3CVo2b/PyUD9Cr/ZssKR9hqfcL0jY0
XN4dUEC4CnE4eSL/kNtjzE97DIBoXlqF0sLbb/vS+s9W8weblWhEb9vSXoR4rewK
Cy0k9uquOC7C7wOFn+fpSYfp0SUO77W7cgFSiOiGVjj6/9igBJHYC8HiL1bKP7Wn
py0Rn52YLHvmokYqXbYkmSa4EY7pq/8w4cglgyywR7Dey4jq1dd3xZ5qvwMARlzN
3Odvb0QBA+9bMyl9B0q2XfO0pzZPpEI/xUhlXu/qxTAqkucalTZflmX+vET9DuiU
8LdYUmijYf49jGWeS1vMvmUp6FqCJJ+C1xypm1BigN76QBX4IdU6gfSLtWChTx8z
COPfvZ6XWqwbfd8kqayHhcQJyo68GBMXMwhC5Z5Mc/ibUcS6eld9h+7uz1rl+1Qm
9ENL5qTVxJoYz+5kApZNQyNNN9m4QNj+sMWnUlBCWNI0Zueva3glYFTa1LnGsKEo
2Nue8tLrxdahCo9Ia2DjNikl012zK5qXJXM6As4NYCPbiedrygJAXy04vEiRMGLZ
Rhf9J9r0PcPaTPV1Lz8BNUbNsk9vzeyqmuSFxtFO9uQLdtzVQsl0F0Bhlcxgug4s
Ky+UaXnjXf6Fx87GpjFs7jMvVqdWpxsww8M3jH2UHjwq6wJUdXXttjydsGXJma9b
EXTJJmJisOixgA355LjFSKs9k8168SsEKJgHfvHfOKn8mZJpVKa8Wu4XW0YIVGCF
vxwFrOcmJDMEvxh7fT/KAaJDZZp1n3MGHniKmSt5ezH2tczZgftrlx7BXPYEzKJo
0T/iqw1p4LMargWHcVmTuDYbSsShoPK8HwcvJCClGHvyBLBeEkYQivpJT9FH5C3v
QjoilVpvtHMN8L9grH+PkglkaugRWjO5HsuqQf+VRfa9U4nJGwVO32ech7NKWU0w
GwjUUWRUX0ukyvMt3kmG3L3Bk5zBypR5FmM2XLGEyicjFxuwONEsb6Wzdr6Q/y85
voLRP411579EGTd/qvwUyC0Dxic71jJm4tgNsBbp5cWWcQvDoKaH8EeNMJpny8y7
3IefTK0VM1LMszns3MtWpDAPJHjyzTammwHVE906FWaWcNRm8TY3kZns/HPDi0ma
/HdDaatRQB9EikQvpXUrb2BH64DX/6TeEJ0+GJlU1KQI1qzOOd3YsQLiL6D5I0N9
VlMfqbdx5YuWAOYpWnc1XeX6t47XYZkYasX0F7om9zqWoDU6Utf8V+UTZDT6eWOM
L6QX/stoVhG1iwqnfxOuuYUoen7LTTAb4jCG+V48WKHg+KJ217Uz6GhQBGz0WEhK
91AqQm+NuYDGiE8KBpVPFMNK6mKO8ENzAgI2whYLke2LD9HEZaH0URPjXkd1/8BI
as5lFzSgGnFc8lRg16z6eIhneT1B/JZMcudzXetzJT5DpKpYaO7VcnIeyJ9by/T/
y2JyNZJHMSLvnjksoI4tgXhD8S6YI6TOxkfZixp1hqq0QzlP2nJQdJl1AJv7aM/l
iOb0DRxD1VUsA7vybc0GtSMbZoIo1pfh6KWMv2c4UCThUi8qCtyefAZ/DKPJIAyU
o+ebtVliFR6dU7yJgLrMtO8a1pmwi9BR64vAwntqHjVeGeBsmqRRCeQZRaevO4WK
TkHeCE2X0mOaNx6oUGYpeMD3Qr3Fa7OJLW4EAbGZLCWvMPNm75v/exXI/r0Uu51M
rDERMn1NF6xHHiOnbDrtuMfCjIZQZO0/ApdLj7OMX+1luGETdZN5ZQUfH7sUFo7G
2TZ/1ehhqXgNIeSk0ncPyVhlEHWjHFLdxWIaSP9HFoE1Avll+TLsLN6Un/IR//CB
vrxdXwn1peXcd6pZ10M40vMgG/fgZxwI9xKFamCe4GHlbsuQYIpZCo4EL/t28NrC
HJu+CqHXICogfmpSLg04MEG+VjNTeACD+FrHJqRb8vBMcmY+yQxa+/AR3H3yY0DK
tr3xMXczOgK+iwDCUcF1TP5CNGAa8vem1VNJF9AkX4gBKw/qtL7NCdNJfltVCqDZ
02ALLReeFrLRuiobjVu6Xo6CSsmUHyCCbx3dX7dGvqgxyLXGayZ0P3pXXk0Y3lgp
c+Mauon5pArNlU6HukYXaKj3tX9rhIQ3EWHGjbFe6daqJ3VUbANa82ykX2x9ipEM
J58lTFZnhCi1HXCkngeI7OCPikrBr9wkVbiFFr6XJh5xU7Ell0OIEibtXx6v+YNQ
bwGMm3hJTqRZCo72hMTQj9dev3ACRy5dLYOxgo9g3uWtqPQvudSWk1Zc+laFzZvY
bUK+IObG63kDzD4h9e0LJ163WfW2CnGYy7U9IVtX56tnODZx2nXSeOPehn+f3mOE
4tFzOGd6yexmt1QaqzmdhaL5FjFAsc1kK8Z6xsUA0mCnLmIHXsn2WFgXyYPfdISA
lrru7NJcL9rZepzUGbX32h881bv1aYVontIUfRM2dCI+TBMPmUrnMw+1bvu5/fgc
7hYeowRMiAKxGr4YfOU+jbsy+d/xiG8/irrJhPqIdhmYZbgYLZjuColhTwVxaFsH
D/t/jfQp1viZ4IZrfEeczNaI9T+3RNvOmuSinX8t5tHT5XcaFM5Zk3tp1L04nsar
PbNiE+6X9TID3mX90XarhtJ6Md7BjMXq+IK95sjOCK53WnOoyhj9Mzr7SlUee667
w6omEinySb0SRX3XhX51+Z9rx7I8XCmhtWZytVrf2YOJztjCwUkFEqPt51Ehqa0Y
x/5GzFCL46bdaTEyiJQ5MzSZVg0RpmQIAx4pF018ccEZg/eMuNV/0pZTjCXaIY9+
1Tz10bFo9xOubRc0XXd6fj+QJxmKgoMqTwVSm+PT1iUL3YWCciw4OEMJlSQOYe/S
1EIx3TANFPQmv0JVYrTuOGZDgkx4lJjqQJlonuZB/86sEWNGcQ1ey03Aat82oBMs
svp0NMJo87hHM64pBp6jLRq8lULNK3scT0zuWBnB2FLsbAG8+iKgr8xsr4HZ68oN
x+vdtjKleWwZzAKRxWEggFJ0cmVc9fi7BvLMjWA7fu5PbVmqey36EiKyrzkQQ0gb
/OwvT1Jw8vhGR9c8YDnNbZTo5Q0aaCdvBmKB1DuP+d1Xs0euS2mN/5P0iaY+p9CV
Uhjz78tPjVLDg+vVUR8vtW/h7/M4Z56LRxnzaiTVQG0A1PsTWdY1b6zhk2g5fIPQ
OG8w2fmcxmQD0A9FRkAxBAAL99iMQiZQ4nU+nallBL7Baa6up3Dgh5ZqtvmIzBD3
kYFkO7kn9qE2a4Z4DRUcMF6IbGWREK+MF/WEwarrIjt8Yoi6djO2i59Rs/yR4Dc4
MzCHloEvqsq4lpl4zsosXr0MeA0LneKd+r4tLtzlJxQMCul/Pl01iLcc4J/2e0Uy
S3wDS6KRDkvM8t7YHtEd3P6rBXIhKIDl4M7RMxOmtE6wUns2ph0Jq7eKKMSm5SFF
DIUSovOVv1XeOPuUnAx5ADclgaPG9h+iqrcLUiMX8JZuSFFabQ5DZDjxe0mY0ERx
M+FbysSIT3cf4huBC9qABHQwqyQ9RHKcexn0VpMWEiNjug1zmZwemMmyyv4zVLI+
48+4rcVbmKoeBFDlt8+6cm1est9XblzUdcmySZOEpJErj9bdHG2Dt2r0FjRyl6zF
ktdzyME19AzXmedVsOIDfDJuXR9VCYmXu/CzXJG3wO24OvWkeMbDvtmCKZ+xcxso
glJyqKnq498xi2Jf/D5ZQ4PjIytNETzFcr5H7BOcj2HcSUqf9NznWZggxaEwStdS
44GCKous0i1GVSQLNQfDMbbMK+iJGbYInHPCWaLdQsvNa2SUYxMNsdm8phaXbqtL
TEEQycIclFiTeAVwI/Qs6ntfVQVlD8KSDvBNYBztzFK40na7E9ZvhmudIXfYjEiR
9EGXQA7r1cmNrPtcs6PIkSGdsi2S/Q5NqSQUuNt89yBJBA4/TpfzSSMpx3h3pG58
EUF8X5UTzEXaAua6MPW38vntWO5jj9406o9UBrreNz3jma45ZYOr4AjDuXR7HVPv
NQQVzUhA4vGjlPQ9feALmMhWKMcdltKsYwVOqaPPoY1honfK64/91MY3yB9PHIRB
lUI6suj/P40PRwPvvnA/8LA46ndhdhYCUApNScd5hhuJL0LEj8aY9LxlgCzM1bt4
5MAdta8DWQzYuCB9T4QVwWBrEkTTdNtiK7s+qW3JK90gXXMTYucjqjEXdScR78nJ
F0CNzGA/KeDm2ma4pfqGN7yIRHBT0GNY1vlQvsGt+uBxqiKzq5Zp35tJ6IwUBy9o
KjdYPvrr843lYIRsL49nuusoIqo33Rsz7vi3Fa5l/GTvxxR5FJBHU+1g4MdfP6Dz
UNwdjaOklMsMPIUGEg9IANbh8WXECAFqILpyQPU4zKKKSHqyOdcOQmQkH+FXUsuk
wvyJOTNlsFh7IqlbtFaOhNcPlXS6xl3aD6vmFd9N9/dJCRiFX60BDMRQBpUsdcWW
vi9mvNIwR8BF+QHtFxtQbEIW8niU1G+1dG4B/S/JPMmj2GrwRDB2TMExqw0R7+h5
0s6WeL0/8tDoYBhAsxmagMbO8xN1pISDDLjUvVBZU43wq/s9G5C+fSRl+eCuSpoJ
a9CLNv6cA5pukbU7N1DeyAs4bZlQz7bys/VPAI/guAuGvbSoqgYnW3mAf1CbBdU/
IlIwB7MVUKDhN4Y7mVlCav++IW0QOt9HE1UZ2I8TY9PoreY6jF8zqEXSL13hs9Y/
1/NEFxxSYmtwR3foktuP7zuvRo0No3v6+B62Y7rxzIrVhFx364v1lzU6Nu5XFj6z
JSVWMRaA2USD+8QcPHKYHYu/wYIsxLInrGZ5KLkl/UkytCv8KxP65lpynhIaFEeX
QIGZ8iBovJSr4d9UdeuCPrj2sWBfvnN2zKkbe7aTn0D6bix5firZ2WoO9OoV+dbd
lvxZq6RhpNY+D97zu4/yN31TQj2rU8IOqlD+Pxn4Gtaq34oGXf4GBDroq5EpFRd0
ZorS+0dOtMoprdj4JE/io+590EKN2mY4X8pNr+07oiOU1Z98+anAULz7b5c+AsDN
faqaQnnieauHWljd/WWU9ssTJMN3FQU72sUzi7E7q5UB0jTdEOAS63SZ9VmdxEzN
zET1CjS2R4AaXJRKVVZS4Pz5rxNnIpdginJmbs5kjTQYSiBrZzcqbr+lEd98+KFw
YhLwAL+sCdVpG5UMimlGjvYI5RV7q+elWo+Zyg5W7BPixJTnt0lT2sl14obGUUPl
u831b3JCYgWJsBA3F0AW0M7L1QjvgSQVJ5jxkBBXGT4fTi4bYvjH1mHGMubCqNza
5RBCWXF3IZmoAdeOPbdxfPppq990mpeIENpiCWNLsYCIT+Xp/6zsLB719lh1hg8S
Uv8uWJ+WecgbgQFnI1CK2B8ZZmG9Gcj91raSiwhXbX4RTmYWiK99qW1gf9IsZY0M
XxF8paElAf9aeqpLHCFVoYM2fM1HERrBQbJSTRN3+8RaiL3D9vSxOIpqwlMzwmc4
dwRJ2+3xbOT8Fx2Ce64KA6k2HUMbnOC4Gthw1z+CzJP0LErf+qVS8kzhajJG0GjY
TAAmMsU2ools2bZWb97IxoTKs8kvPAlgiwKs2bihtbi24VYFwgG93ewu9D7lmTJn
csZIM1RGGjHBHjL86kSpmTkWwN6YuScxr19uUBHQpW0X/vQN+7GWxqlZUjMGhVwM
bx9kVMfnIE17M/B1zl8tvHLtgzgvHAGmCWtyNsOgYCinlCUxQoPUzsCu6S/aYb7r
1Vlw1aCwrTwayH0nhzSdkvmgUcjGA3er1EsopaMTUD21IAq/P4Em4ddyFTPcCSbR
HgRPGQA35DR/89ImI1DrbQObqX5N1o9edS5nqZBWRzrphHXk4coAg7ODVBkaJ3XV
6h504wwcsnLrnDCi0nqNQpKQ6jefO0BFLqBdLr11BspbGraYGxqvNrEdCOqPe/MK
XMcmrT1qHbhujQzJRSqb7vWyz5hzghJ4Bk2qPedHYKagvUy1xcvAIW4l2OT8skEW
E1CNDkdggWIIUZ718fXO8Clz1WnZ1AK7VIdUA60Miqj0srIOYzfRegPwZBuEC2rz
Y0PYSHzthflMgIv2Y1eiaR/pjyx7y7X9YpcyaALRn4LzNHzuur35STcNwcxZpTuo
YZ6itPYSpR/KJqtBxG9BRaCV9ehi8o3bjEgKfyUIU5lBqSjVpDSE5I81SBdCqVFr
05djspOXT/TMQ6cW4cwlt3tY8CHIW0x+pTlVCPgNN2p6PsuNSkz/sEUZeCS0zUAM
M5JWE4FGcV8/XuRvHok1lQIuQpHBTb28fgwa4Gpm7zs5XN08rzUVrWln5W2et+8M
9Edqq81iqZ42EcMGP14uzM6Zj2y4nl5a2ZgRSOiB8zcietnsMMqRoYQ+RA/kOzcD
AjuGuffNFEv/0u/9Iu3Z+tCfR2e3Hl7I0fX13dy+TJrx1Xi4/tFhejj6BDaoeh/T
zc/A+ZnE7xqyFNyDVisGxbzjNID3efGq8TewyzLllr4LWcVMsh7HTPlkuTjZLL+f
FDh9NjZrx3sy/4ayiYG9NYraK1xIgywX9OOpNjf0fHrgk1oo4ZkmKJm6zDQu0Q+n
0eZ36CKcecJmMRUmOk8Tjzyua2lK7l9E3jzgR8oczCZEsFdTE/zI91hOa8BQVy/3
QSiaqEE96o2lqT0Ov+4ailU+sSAxLQ0CstQbujI3pmLPNuSHGJ5pmrk58w5ApCMo
x91HJ5odERRO7iXlhrRZtfug9m5TBGBkCGB/Uchb/LV0VsKKJhNLR7NwUnPsXBSb
b+6xnTvwDPsIt+MqpLO7U3p2zUD/dRmCLcEww4JkTSLNayXB6dTRk/KtN29GTXMT
bQv+yibliVv7YRsl97OuNxVXid70Y/1K4jk3h4Dq5z0aAfGvsqdJufSAChVT+yU7
DQCnEpgTDEpoyFGomyraDXNDkxPk123sPo/32xvueH7QR6eSrDlsozqkpITw53oP
4G8gR2xUXIeJt1hLDx3ksjmf7ZS0tc6Zcn4LRpNqE1tuuwcLoB5VMVL1cEGChZPa
D/7+7SMHBVqL4vb/SwXJj0z9ruuUl7hixinBWZsYkApH6lHZca9CRrqi6uXJm7xq
sYwbmpBNMyDsXf+/ExCyk8wsKn8CkUXd4ggJGoiQKxWIwSX/sWjfPCBhqbv+uhll
3nm+mDBZCMWSr2s4kDIpIHPYebLqIS2WF8Zsrd5kHBjdwhVFlR6nd3wyJR98oZNS
rUZIRssQTPjE6CIOzYucnOhXpRgmmANR9kATiloxw6GnhFqzwvBu9+wiQ4hdIwq+
bG4kG5rQprVZ8WEtL8h6s6efqasX/zVUjpdz1MjgNwBnnz1N+gvQmaEr64vl09IK
xwbPV/XGVuwNtkvFrZquyY/UxWYlJanvujHemOKIKZj22BrE1SERLh30apEd6OEK
a1rhK25Ok5ZD9H4McKtEElQolb1AeZLZZLCg7g5nm/v4+nqO5kvY7re6fi7pZf8p
Ls++/PJgO5q0dB0o/9s4rujkr6yKg6koXRNDckttq5GLq8KplvkoAMiMxsDxZioY
d/Uq3wjuH3YPC1edBKKgIxVKzYjvV/S4D+GV6zhyIubB8thU6WiA93lA0Vo/ZA5Z
GwjV1GzW5/q4FLddHkyj/jCFrvNHQicERaaLXQTxThOlff1ea4bf4bm1/tDZSB2A
q+ovYzCOsaXHq6WYCQ7puS+HL0lTkVcamLrOauGZQM3O/JjQVpeuB7UhZjD+p+nB
rS7VbqTJ/9LkGT7PZLabUdMCtmblP+jE+lb2zJ20eWjYsPvi255KX/eM32Mj9Bot
GqTo2YcnrYkNSVmcWlmjcXSAJRnwz94LssMM9kQLYK6hsixCGeg8VTbtN0rPoeIX
dy9zwo+5cExsCvGLstq57F/lv04EG0j0jF5SW/64IZKVZ3eB8ukFDVztbr71yWHo
9QBeFwMSaFb4TRAndQ7MFmMgd+AXRuSA4uJ17XO4+dXk5Nfq3WP/gcw4n76J06o+
36+Y+PIRDbq2yF6vXjOO6wdj64rnDy5Mng8TEMw9TFQkxetB15GJNjgs2u0HMDIZ
SWeZUZwrFpQCGgtRm1a51oCOtECZpLp7y/gZILfMIoLo6MuZoAy3cwcGaxO9abAQ
asl/g6Ee2i7t4fEVaDQrGFueHVuM21f887N1OaEJbvBf3jlqptVmN3PSyMOqSjjZ
G3pmjwUre70UJ372zDv1MKE/eGht9WWnVbISkvVW2QSyI3nsTTRc/EjurwehfslO
eLg/z2T1KKmrw2hjvuxsa102rcZZj/I4nLdvNKsRXF3fRMVOIAtNHPg8toiruFwi
/JqddboyM1uHaoRQfbNUOTROG6IRUGkx09XVAiD9cm0a+Xm8ssGTiPOTVVsmPNa6
bVAPFUpLSj1mzc+54dGWymZw2Kko6n3eo+dM+TRh/zgZ8SpAyoWkXRJhj6jomO+n
gxjOatkcKbaJccwFNMYe/8Qa7RfRkUXWJBu72oIEjRHw/SoCOmyELWZoYtyGBHRG
lrVyF2BYlQ/KOLUV998VIHfLEL++HJvmXCL4hq3SwFmFr1ARC+WjQqgRacnMIjGn
b48Tj5/5uup6jVqKGUEk1NqRET214itMytSBD30CPDA0yRK5AgKSkLTbJrp6yXq9
aiDSngYa5gFYeMi9Gn199W4PZwRBkrkk+H4EfibFVbhJtxqgv1bLDqgeOVpPNhfy
2Fnn6C8mCbUwJ1hStLKMZ9DCo4rCJAd3uYFYHt6VySCzDzMHl02NhP1cuevhQy1h
yN8FzxqGV9OUeLn+/343uCvSQfyYy9ps1jdBcw5OdFF+fPiHenJ6DVIluPnkV5b9
qStvOrMSHQcgAo3Wh5ECcTBjHvuThwOAcu2GSWZxv5IrObHIAkcjUWeTt70xfdCy
GMubUOpLD3KDGs0k4Z9HH5glcC90bIliwUyqb8E0dGoCis5MAY72Ie60Jh+aIh/n
LsqAwYmkVDO5fdsNxkfJx+hTA+r1vL/zy5ha1FnYQ+WejCwbO0sKCzwX0MrqdrOi
7cd2705oGbB0s/nZ9rplOWJ8SlcOtJHjfduIlPYjE6GvYfksbTxtk93YfDTcD/KF
HQIm7X6MNXPyjFWwgCw2Dmqpo1iz95hPOB0fhl/8tpGT6RQ2ahIfBZYIIRPhXJq8
vDgYAFxqn+B8gcmfUZMAvasiE+lGnLmKktbXXa1UstFat39S0+OdE4gc0JpHeVBd
wQuukuULpqG5TZKELmQXo/qssJpEPZawx5ezNIWqBoO/a/Ls9vi+l0KCTI8FY3Ai
WVBPJv6WA1AiMBEFTA255lTHCgRSSIevtLhgEmd1QAWe3FP72AeKYR+vrA1j0OXO
I+1S9mShplb67/pFb/sOUwdsw8WTPwpvgCYNSb52I7OxX6qZDQz46jTITUqITLE0
aQ500cCujMxAEo8QJO/5W/3Aor9Wzlm9+TKaiudIXjO0ctK3HWosJmVBiD20Bo74
XjvLCiCrHkdcP39ag4kEDzLlov58XueSSHvb0AkU3IGry6Exn9sgI6mo/mjwTPQR
n/6Xcz+4ahC/+YvKOyDaX3GAhAOktoLQhkENdvktppIdKaJVT3xJTWvpvI/buQgR
D2DrbiGi2/eaKVM6JI+1mHchsjIZDXZpoecxIOQW6ukt+U8pScFRRebaLU3hUMVz
YGWj82yolfzZv7XIRueuc12dWTZozI3dmldtmCI78ZO1bb1RlslsYF3fBNwMlaHr
k81hrs4t4Hrx+UgN5oVNQaIRwuKWCzhwbYhHoEHvGlkuz82cZMKtXDCyB21VpIRq
6F8hE86CSA/iLaW6AODHt0h9hoV3YOlvcIO7k/+TTtFCc/aIMnH3OYLZeqhS1jry
0SzErFUGXSJfxEKZYM6Gvj4EQC7rfpU2UU8jKYpQsgnYG0Q4o7sbwumoaObSTvmE
HdsuN5nFsr1gjyO2e9z9GMVXK7DMFO2uYV9AV9qV7m+YJospEvUyDxEml8vkJu2V
5Nj47cqfrrUvOtGgS0KNo4uB9+/H9dhpbZ8U2x1BVG2sb8plQQhzNoG4l0ZhLHqM
LBGSRVX2KEhCPaTBG00wMclJXol5eqG8dn+xCCfCn/0YUO43LD2YnkvXC6OQXA8+
EiXhB72HoMCr8+gRUdpZiSyVQ+bnc4ZpoxYm10LUvA2v8dhm9zC2zgVmtv0hCId7
gmKZl24sNXbn+jR5/XZ+LKi4W1LPCIae3dnMx0g6+GbX/9NgEESyela3NfDKXKsa
m1oL4y6YddxCiIvJdOvLbNvWjTQao0IqaUXNhIoFnO8MK8qDm5aGtcZJNrZwga6E
PD7Yrw6CpluHMIiHiQSq+jjhs3khP7FXpDC5Hsl0MfuW4HaHt0UsuV51HdtsmzAK
ttg0VyHpCnWGKefbuKUdkCdFZURkbv3x2BmUXBnhguceErlGAgupKjCJ8hFuLr0h
++Q9SUUkSFNZxbmoh6eNePpVonvFI9Kjatj7wqDDWVQ4IwAKnGpXIRLjpICBKrYr
kWbIL+qPgHoW5D9qBEBSrw62kcfj0ZyW1tFYHYXaXkZMzGVO1MA4rzS5rTsbSYd6
MF7jJ+F6010meosHYDTQKMWtojvu4eEGHDl3DJOzJFHkJTFA/vHx8v8hj2FA8Czg
n/KIZ9/UldEZUB9p0prWz4omoxOh0dYgMmLLWMlbEsF2ckUGheV99EfioYcUPQJp
XCaoJXsthUpl7ifcsxv2AdknzA1G8TBuprrAmeHjqdfUDeJJqcDAfExCKOauJsxG
JJ+cecV3zlUtbRX+psG7flLmNjGZidBxo6eB6kmDuIevZoySGIafHppxcdwDVzQm
jmPVqumt3uMqxhjBZVOKsQ2TXCGeSWjBNR83HfBNaH1EijlLJ32VkniqZxSPDinK
Qvk1Fjt8aj0Hq8ktoKX4RHlk/Xe3jFRA3DzOrmwHGtUq64G84vgGzyIeJ8eYnY1O
SGMujCWXZdjMRcQ1CAquCUhQo3qfoR4BRaUT34a+FZDlNRrBf31AHf/Kxs9YRV4V
BwxgnRSpoHhY6JVRZfE5FFDaEzRuAMoDmoWxOg2D2BL7mja9WU0yg+82yo2GLnRL
FZJq9JC7DZuOuoUrTR+9X3TIm92P/3TJo8+kKcKQKCoqAfy//E8KBLMjlDjtEryD
RsPm+duWNj16L1SYbTbMlthIO/l5LBfcwOWm773xEaRvQpC1xNu1r62/VNjxz5W4
Lf/VObK7ii5nNgH83hfhJw4zQg4foJTvyAFb024H3G/1Ukks6+AvOK/CJwbjDiqT
2716GMw9DsNUjJOJrixLgZz7Wqtff0bDKNEJRG7qnKb0BuCRZpB3AX7GO2sxXjNW
S5C0q74grI9D2y9vfaswDfK3WYirRWPcQCuLYqQFfJKhUwe65LPoN8axxQgEM5MU
yIaiIUhzEtBp434htyU8Tq5lPh82dOp/ZNTZe872z1o6kEHG7uIFiViltnBFiZzc
qu0TEx2zJq1pA+1tlP7OAc4FbdfyBfLibS2Ad40zHEasslaXz0lMSUQrd9pxg/2k
jGvWSiBDBLZlLXsGxufHswqzwren1lf4MnQT2beYncKbVv4Gpaeik9IfoFoKfdJb
xTxV4rUKXzDrHMfAusLhiUcYjmpr0/8U5iR3W1g0vOhemDsIiv3Jb/lb6TqzfgaY
RoquDqm1gPM9A84ajxRt6FrQA/Il/qTMa3TgWlYxlDEJRl8pqlOmljFv+kfUU9Rn
wpwUKnQvCZqiYL8Hw9EvjjP9O50HdMAKwbS9AJHxs2aZkDYKqv3EwH6fb9AvyuRI
fn18WCLavbqcQCsVbWexcNR5O8T3Tq4xpiw6trTwq2WcPAV9rE8pd0wZJJ/4btaL
zA9Z1uMzn5URMsh8P5zXH1Pz1mNH4MdxISvYc9ZV+2EJfm1mG3jaXUOd3g8oVWtr
Zpmn0XGjh2ZF5aHoFWec0fwIKTZ6I5iuBn2wTa843icXL0u3FelorjtQor49FHPW
8dsh5URGQq0MbhI4OtUvV9dmW7COjW6N7XCLp7bR8tBvV6mx5aHzIVNFjhkYIgof
FvJ+dsjyxupiS4TlvFhF7BNbNAQTviSv6u84Pvc/u31gTfjJYZqQ4k+T65Tp1ltR
MX4y9U9GL51oC1PpNfGdejkKchr4mIKiYAJ3inGH+gq6kcU52ItS0zMrY2GccG/G
iYdOyH8GFaRyTHIvDgIn5x2QJV/bzHvdQbOt28zL+j2+xgOm3QDoXF9j7nRkBKqd
JHDXzfpsrw97SsALb/+UE52y7kZnenb7G/3xtQdxAwdDMLQ+q/SVHR9+tI/wlLr8
g5OJYmMs/L9AYQDlzM1gDNj/2K/4zIirPgsRQSlUZ7jFC5q8MJHXZN/Omm2n9Oky
o7Q+1HpwbyMt37/yuumKNFiSuMwls14kSwnntcnQXk2e3T475MHd64Vc4THHVg6n
Q6iaxZ9E3qGp9Fidc6Yln1dfqeUW8ahLl6ZWJA6VMib3io47ZGdvFPAUdSjxPokm
62hkyVnksOHmSs+3j3RP/QSRaF1H5iBivn9dT3woket6dWmRvVfg5qwjTnLp5JZZ
WncrBmVz0YTRkZlJEaiJgDjMj4K5HXpEHAcrQJN3MgbXsvneAvuFJHn4AGi/yf66
S7cPlksskcgnjtcOMA4mMybTxvU9mCiNUEOACqrqfK9/wHq+ieX6UtsIGrW8lBwT
cYUMULYvRkW3xn+I5nuIZaS2IMkWIFagPzfJ0wEkStGfbHmczVv5ZVUDIQNX9Awl
FJswXVq3EqjHQuIRwQ2IBDcBgJJZhTMbg97vuPRG4cq2rkeLV7HgHc+aNvjvJDqG
07HoY+2Bc8pI5zybkru69svuNFlrXullXAO5hWR0uXPYcQodlihbK0kXr8jtgdU9
LC5NbRXxjwJD9SGMkqE3/+V1vmENm/9hprszu2UJyO/3xTIKAEJYRroVIpsw/07L
ZVtNwcQ44UFs2Ma0JRQP8q57p2W8cU8BUw5wStjXOEO79WNtQHmiRMZOAArSWDgg
nPPsufNsNJEC684wIx2kXnTtfCfaC2P6rW4kU2K5WIrEAjeUx4yrPQueXdaIyvyJ
wPSxUhkGie9Rj6ac89iNKlj2JKvbq8fZFXMIHg6xDMn5fOZAisDyFUmNV2lHQHHv
XSl4G51/+bTtkwIb2VdcC548jQcy95vy3mxpvnDUrRixxVFD3Tp7sz1rYv2jPcUS
gKxU9g2jiV6/CYGFZbfdEFkjC1L5xNCarkvdEJOxidF+sH3QFwGtoCWLEWYvqYX3
KzdFFXcQev6xHEf3+KWcifmSvPbwFddgIq3XdH3gPJc6i/tfoU/gdlPis8SwVpfM
wGw5tcjjg5WqnB4OqicIK6C07vdHaoHOe8gsX4rPMr4upc/OoTYuo7AxpgGCVGkr
SYScziZRBbMjHudDalu8ZkFlNIlTZxrfwXJrA4Ye2GPJ/FhuGL7XP5YLdv+UkMTy
usRlhEjih/eabxiHvOQgn8WkVR2ZblPWrhA+7bTqpsFOjA614yNcEdomE0e3CxbK
tPLH8Vgzpa3Dd/8NZvQ09jp/D5+n3sk7kWkXl/aqBCA0lTEYk3jFqf7CAdeTQnVV
VGqyKuZa8wF0MBPYBlJXYhQpOwfPcGE5WAh+nz6UsXCZagePn9gUBdD7N8rSmVJ/
L4Knj7upf5++wiRg4q89YPPAdTPggQvYGxYPQFxLRsB8AvTUEZxVR4dp4mrckNyF
Foxay6kBqlSGBtuvTIMepsGX8FOIGOqmOKEImfw0tbDpwzZZBi01hDm63z0mTH9M
0QAGGUKm7SGvVKK1kEn1dgFoXeZbGFdH6Ek2vPxvXZskmmOV44mWgERjP2iMcNg7
5gNZszih+WlIbKfk5jwRmcdDZKmnt41+YAEzBbN4Lq/qOmNJdfDtRpdpGWAP07B3
ay9L22jVxSV1QqaH+u5GygRRIIiMz2Hkb89QPZixVmr6XcfWXzM2KbPnzN93atB9
EefwbApVnr+8TdL+av7uglmKLaGNdh9D0d+KaVFeP2JFJneX7shasxWQ6+GsqUFK
XIv6EP1vvuJd5M68MNe5JLtIQUuVFvM0Naj84CkOc8vPQpPHGqZsKy8ZTxRPMhsh
3Q7WRBtZcbBkImwxLVlA//XWdGOEzU1WHIxRfG1VYyrPNpFyeXwHT3L8sOEBSl9W
jDUUMzm86sqwC8FL4DEX9vH1lJuP6QXiu4gIfX1mkdobI0eTjJtrdepAXh4E9QrC
6GvsGsSj4m2pUTQ24WEyaSYxWPNK9hwrNyLp0Bboax4FwSSObsPc39g9z11l922P
5zMO9Y+u6HJVUh44v9cV29UnbAsA8vXOvDPvvSjFl8kY94INKCxcVddzH0eE+xtB
mwAkRHAb5SFZyA5e2EhSoz6SQ4/PdUfC4RMVULX9JA1K6hBGkghc8KwmiQSd2el/
8BU1kFTI1kHDvdWr0Bmeetanc/2AZMSmwDItf00k48hEWIss5H63ha6KhyMuP+MB
YQETlXdEIGVpEFZA5ZZ8sovQHgqlNywOWg34FI2jtMgc57bEIEvCU7ZWNH4Z3ZH/
/AAtvvYVngc3LnjcBFz+CsWjVXBItv+yQdfr0c6GywFLmAErfGVjaCc9w8rmpOE1
tw1dg9HdGODxlEcXLDW9WiXLLPz2ioaQDa9Fw6cHD1tY1lHTkjXO8uhgVU7JxRnc
0q+gz+F89bxoUv5d8+GFS7V6MwuHVE7jfXvXcwdAzYSQ7NDVIe6XTA5QDk/FejFU
QypdG3VTP2s3kgAzqluvNibSOQQsox/quZ/umKx+v50WwnBLZeSEQdnjH4/IPHzE
NBJE4QH/zqj/AHwnmo9X3etjdHPmLyQx+cOvWJkLaDKrXNuFvRBA35QD4YMOIi63
5IHWwyXKdVqqpqfUoZfyE4Brdiq21UDOwo3V6Lkm4fz+QDUfeVjcjnZWVBBVpn8p
FDDVC+kmQzZUT+xtxEUhss5OU0IQkzldGk/rzyQHPrBv9E5wSW5UILrVfSi4nVYw
vcNb4ObjOpOGbse3wB+QsRMWIf+q6k8eTLrq9wAKlcdiQtq1e3+E0RdKMZDg8NmO
E/dhubju6qnOzfqvfTFiz3R7UQt/WyIT/DKm1s+r7DCcOgSEjEXlNp1NZ8k/AgSP
Js+kT9qYVGIiSrvDRBc4SjtNTnXl8ELxEUvAfF91wD4BI9EatGcDkJDwEad0Pr8S
B6zk3WSTKiYT4DwKahyAYLflONKnU/a/mcB8Wtj3eIte7PnP3l06buzlIuneCOjI
jE9QnlaKxD3dcdlvPP3a8nnA9kAdB9IBkS4VNoco8XNeL33slonGkSZ9lAEiGeb2
ChwPncJ6jQeC78sfQypcIpONV5nDM3QyqBsGJ9SiPRsqZaLY6nxswVKouaqLDf/r
Y/M1MeZanHHdK1TWx0wAmcyvTGeGgSV9cjjfxwnlCBYDHTh3EYmKgY7Tj5kEGcyX
hnVod+gOPPW6neZlInZFQQfVBfHclNmgLyYh1OsGf9rgPR4Y7pi1NxhfQ368clO4
QYB93AcjiuwS2K3useyDPPJUbQTGer8mJG0+U6cznsIKBIH3kqSTnBJFFHs94qJt
oaTtnqiNwCgCtt2KJ04z8nThFVoqk13EcBtBfQdxB4Td8U8Xpwcka5rnyzZAM92E
ZNY0MXQSAHqOQlq4GTWEhXMuKlU/rVubNBAOSIFnoE9aY2b01Qzl2pUlzWRx+8+A
NtskiSLrLcPTNC9WyzG01VYZPOTMolClo9obHMTr3HM3XhrTa9/dte/S/sqhvp4r
5VoDtDIneBjvFB9npTGuMsNm83dze7hmqTTxh0r0eKi/xGfXDwFpyybNWtvygyrq
3xFK3YBRGw09mpdMOpj05jXS1Xa1Dh6Bki89cw9IxtZ3Co/OFnNAyXrOd8Ed18MV
zX3u9OGfnUI2C7XQ/e6IsaqDDi79yGT7zHYg8Yk+uguXWR1XS2F40nPk7R3IsEdl
BmfY1zqe3dFgG/Ruv48MsNRiMrICgNOjSFWWEOkm+wwgbLJmGSwZeg4WUe8/dbZe
KgbSLFMrjgyknkpk2bMjymrU4SQDi5NJsEfqCM3vk6G3GDehVvP2EKuI+hF2j1N3
MMC5lF5BJ6DGyceAgfdLJ0BGXKMixvFvwqcNttg2TtRHcV+EMb/MObh2ydPXcwkA
pBV95JXgg88pek0jnLdc93ymL+dvHSl0UWoNh9V3zYjk1zDJxUooOgPsacySVmj9
dfMTCxRYDZakn07Rs3GPUyoBlJWGaIEYnu6+qnrtU5CFQ4mubSdkpYkVpSm1nbi5
o4RbnRp8amsLj69KNC/uy+0XAmNLHnP7W/D8x7GDxAsexngR/w9mOTQzKhBWMBru
aQVwehtDge+gHwVTDMG2QY3ysoXU29Q/9R+W2rDHuqMtJHzUsUg3QLro5hJ6abLG
IAsNIbWzZQv1cB3OnTLYf7sa7S7n2TOOh9mlzQMeuGbfNFgTzhTI7udN3xsG0Jje
F5IE/HtIOHrNADGAo602LMgtsomXQflOJKKHrUrlTI3n5kvxLC4thSZFf1mdkby7
I75FRjDnzLhxVjr8dm6TYzUrRVizE5SHXYJq0da607SE7hCzUnwkK8bHeITk5/EE
Vyu0n+CsUCb/mPGfs1jUqrjVVdK1SdwFRRHWyv+/WnF5D/iJ7dAwtreAWHMpWjUU
DQUxsXL37dmvUqid/QDhaGQnnBoWeWy+WV/LYGAm+ehMgSdyQKXDhUaEniA4SvcY
SV9lS7QkOQiw0FQYK1Aqvj/jpqrulbG93apfwhs2fJ1QCrbQtAoEX6IoWAPaHvEi
3DMTyhuuQSwtpPmLcZFevu81nwKjpLRSGTEaIzZXF7fR0bPtzde/WwDp7fH8I64m
qxlpFUXN36Ye62HULbo5uNXStU9atXAOB+ZlZgMkRRTQDIuFhA3e0uOCPvyd2PZL
4MhTGCE0nFAPli8Wy5JKqBPuzv2454C0cCaWSzEsUcX1lDYINSJdxLOUtY3uQsRU
Jzie7Um60VNnxeiU/Uid9xKjYZFx4hhIhOeig+9l3UCkjuiOhYQ13PPLvjYeLXCQ
nxKh3+DyZ5qwwIPsO1Vuli1gMa9TaTFdRbW7fz0sJg/lLTwsQN3x/7OnRc5K8V6b
v1tjR7aPX30dRT9s9rm1+3DgCkqOi00NCUpfRrNpoVk6yeQyQ28RBhVMQy4aiE3Q
MtTLc0PtN/pPzshtHjPUhQ83yT7yhmPcOBDgs9o6ePqUNKeKw+zvUzlR9KPyd0OA
nfKovkkFZkkNd3dj6fCo6ERXr/zdhg3GK5mDqFuMkg4xByG6hMqKdkHywckOU366
9QrVV/oqm4eVEXXZq0PniMfTugBSLBCbc4YYIug+yI7Ef2WwwyWUlfB11qZU1+vK
wYKd8RR1xq2laaHrcmww5ijcSouKrJRpjHQGrJLMitY0YGzbWg+ch6eOaJzZ8T1h
IOkS+XK6hrJ/NN+kIYAJUK0n45vH/3y6k7uS0MFIXHaRstbIjpTcCOC/wKLjyztV
Y2FYHgG5u6dg+Lz3JPqO3sl9D6/hj/170u7vQgxYpparCgh6p28FZJZAMAiIkywH
0FxWUv8dmv0W3W14at6OjAph8TkzhIkDEBRtiCJwIHtQJAiofWTwX806z7zaSjKd
POf5L/Sr4MYGSpyyG8C6ggzAnayz+k+nqOqHX0nPp/tzuFcQWxNR9kx/SuC4iTyO
vTHWSjBq07slOEtJxrfLVsf3OJfiCmOhYPlKLIEfqnxPd36VAQVGhYA0rFNJSoe/
onJzZfVAYX/8b43v9iHg3pORji6umC5zHF6gNkJGUpdK3sMH4NskCBIpHa1AhPIR
HK8sDt3axqAkaj/kwKvwbK3yEJ53lLZ7w1IsXyTLHljfDoQCA0P93Sakr4jqDTou
uNNTiNSuqmDdUt4tjQKaFUDmR2z4NwOsFDLrEjc9N41Ny7xZpTql3qbdDVL0X9yn
ew6ggx3xMIIhZ5GSD2tGQyVrFQVPIhx7SjUBAHmDSKr9117jmlNfbbSnbin6ZEbc
C8a2su7PPCGBiBs1BBcfYQaFNF4JtiiNvcDbsLm2q0LomLAfESLjRNMF8+0aGGIs
sM53ZcdTBO9CCLCWSNrfpPkP5yWnTopiJdT9koQ88WTsxz8P1vKr2aanQB8MXka9
XkV68BUeD7W4oSScMIUh64BYc+91nmZZe8nuuCW04tSojKUk3k1313aRAIqv26iL
G5Pa1eHbDcOT+J3z4Tr4I4QxVkjLSoWKdMYcpFso3pYjw0oa1Ncty43icIGpxYGi
iXNqsadmii9kDjVibJP8aJw1xZmLTRv1wQ5gY02qo1OiTLk4035cC1ZBcb89Tovr
ioF56zSBzQGpwGv/jNSZflhXsrfbVLzjYrPm3z/8SurqRsSlAofaKcAQ5+hKKvIE
SSV/3ktfquQnucp46pzf6lW591znBHxGIV3ZR/d5JBcbDM8/lrMROFB/CqJZlrxO
oa+Rbv5QNm3jZFIwNXrrNlUy1s2lKRjVxXCKE1LWwnLIzB4NkWYuBHKdpeVFP5wu
EFEfCAimkJ1Ifp4pYpzKmq4O7oCqafz1BfyZonvB5CDivC5y48ntvqZylNJ/GuMo
09NzYWB1e2TFuoh0tU0mYl4C249uctctXH+B4pWzsi0QW5gBBYdx2BsTYW8RR1Sc
66ekM94bX72OK5fMgpTWecnCXYzQEMKdZicRN5OKn6ygA/eC8nHz/Yfi/AwHDNVR
xEk2tQd3xUX/n5EV8svwTF04WDutFXTLvJjCr6daCCsbVl2i4AIKB6iWL1/re7P0
s5KkVZdXbmJ2Kzbqibx3YUVn79BVNBd46dCFSiFSd5aAlq17YOwRnsozkMSHMcy2
8VgR3vk7IvgJvTtGdN7ti5znTRisal5nTfLLHzZHlZkuTag+/Xz+PHygaDfeMAWQ
E7J4cpaOlZncw0pGPMCFXW7ud99QydLMWEJDxPcM0UtSvpEjPpramJHp5xTqqpGM
Yn3+zN/9n2LbhbdZuoY2lSbJinZvwX9CungWxAfRv+0GtBA6r+l2PWmFBA+PzOmq
UViqwZqB8y/QuYYc003is7qx93v3EYOEghQT2hegqzvGQaw/YQ+sXx8LjlYJR2RZ
c2FqHlfDFyFlFKAjSHn0RxptCFlyIQHifXjLgz540DtxlvjhftYZILJcog84uvMd
9q0DA2NSI8IUbfeuT6AKfhDtJXZPUM1jDrctp7fCvDgBmUZ1O9sbIR00hrnQ7x45
OyvI9+nrtgN+KfjjEI80fOp0Sb8v6eiBPa6ughBxfT7DDAPerlpsElTGGKxlWLpd
ETrDtv5sNRCQk4QXAqZGaI55wdF7mzQ2xQD2Ikt48ngpynziZaaipow+3tkfgbSN
Pp4WYQwRpO1OmCdITUbNfECgIpAI4wDB94Wyh7ob1dYPuFl5e1lisMDptu4BaAoH
CGTWTnVEcJWQGdbT3tpVG7LQqrJ/hGoIZ9Gx8UWXXbOrzlQY8zY7iKWt6t72uIrP
i15hQOPt1Ns3+4fnEI/m46vddvCPxmtNJ2HJuwmzNUQmfgQolh54br4RtplQN9Ro
VePJZAMQjyqDBI+LTrijrZ//QQiWWr8bZMYO6Dyw8bZ+4aguAt8FBn8KaOSG7Efc
rIILAwaTl/dshkizQTVApUaRCaKK7k0L6LaVOLselM4NfU9VDuuxz7UcEx1REl+o
jAEY8z5ugPl+bPvzfWXP4SgJnS3uj+EemTTunk2zqRrHwvZtNSGdivpdW6kQdKeK
bmhXhyeoH6W5nGlRUvYpc9GadIhw2splOrlEd7PBPb0UyOt+B/gIa+HHP15oG2Ea
bKpDelVwYXpDZSyz+hs6k2gwrzx9GiFlP0BYzyCUsgr3/PS2zwhtdn1SJu+dcZT3
fr4OD4qzVYBzOGT/VPdExfcbObck91zj7US7+lbYRqZAfYi0I7Q+uUFRPkC/yhyy
1h8+d+/Coq8Zr5Ndo/emC2c50OjSYpd2WaU7e9JJPAhST/CpatHux7utoBu5uvpN
bO5+6v86pemuvL22XJhOQm60FhpsEaSjrkTHVrgp3+MzvxKoAjNr52XtRXGHG9lb
lhCsFwozoyxe1kOKaOBGY7RFxmMiKyMqDkk5s4wLaQSwT36/uHIkl6aMoJhD+MPU
VspEQGOwy53QwXNH0TLaSIatIiKh0BSMn6qgygwsGK0qv45+Ifxomx3ck5eC9+jP
4Rar3rZZWHZrxYQUwRqRBHtbU3QL/Pzuo7CSGxZzWbIDy50kQZLl3OAiAopTMuJO
F6yCQ/0A8yjz9v6HnwbsrHQUGb/XrBamt3wQGw/5P28ysNBZhFbk64rITwbaTv/G
69msImSTq/xxa7K34G9eB1FTz0msiT9zB2cx3k+FHIeTX015eZEw+BG+ZlFyHSyo
i8/QuBH/+lCx2AlX8gZzaIaLDkXlCWvLzJ4IxmewEm6gop6Mb6hFXVC5t+hFvvwG
aBbrqGKv+YC9xFrLkK1dqQLEwQ1SWsoH40ml+jBZIkcuDwEbUAJUoSpSqgMRAqyb
MI37AKO4lzWh4TwTFTD+j8GU08GgtAlsQsCuNSltZJRidPHf/BySMOvshFj1XVbM
ClY4Ck43I943zxNEOYimWXiA5es7oVuxi0kuontLzuRrk2R0AH9S0PX+2ESiCFdj
mCqJQtdCZJt4xI5BZmFePa7D9lJQxPeX4MQhFsP5Q8mhZijUDauuyk9pfB51uveE
XZcEeydAcq+gWsMUKMr4XCNQEiV357dqMZFIBqR7RW548Yd/PRLgBeS+ApcvMYmC
sxmOFFiMBBdFWAaUySjqtMLuR+c9+KNv8Q4bSb4rSkNKTPJQGwOTIPEnIOkBLKW5
lCo2++Jrtt4+dOnC6WRL/qk5z7PwbwEirpBuXqjGiIcSyRNiKPfqSuSChSTG042R
rquNhCpYWtZeYqxBFvFLiqmPnHmc0B3M/QP3jObaKy/ZYGHv9IdX/6jeHW8lhrgB
60Z43ZfjwW+ViBTu59vCJueuN6LkDWGkRuKSetlH365XdykpgrLUVvhu+WA9OWgc
2CUlLB0za73drniowUIc1+gMF21F4yNNP0jVKJmtdd0ciQZCmcSfim60rFmh4gL9
NlccOi+8YDEakJUfcwIoVZnvxiH11Z5RvFROm8MN6FDDt6KvtDeBVyki/wCajKL+
YenV1c7QcpZrcFerAJnnJzxn/OxOR8WUI1ROliyShJhokr+TpPW+K0t+EF2w0l/d
D9k7pOHcMHHtBPEUAwVe0o4oS5y48AhJXrayJA1bKwUuyzgq/o4ziwNd8n1BKcy1
5pHmWsjzNojAkM5E3DkYKmUJEewK4sFHl9+rhhhY0PS6uTOjnVinBlhT/ksiNvEh
YBGbjAv0btdRsqHJFUt8gss8Rpse9N3zoPl/ZrxsXj6e8EyDxxT9tiUOGkK1zb+1
abDMYc59FSx5QYMS6zPFxPYZRgKPrcywhggiSusOTA0hDnKcjm6Tx42GBGqlMhZC
7JRCHosFWeHQVqDrPhdp2yQGqnjf1z9nEpsJX9jIOt7zkaUSjTX8eo69No8fgU75
J4rRE9izxOsc1yOVwHdvVGTHMdfQeuCydoSXAqqvDC6Yv71l+cVsU4EIYFAg2Ykr
810R9COQtTAB7UkPggP791HuG+KXUpVRCQ6PKSd35988J43oJnDMb6XfGvfHYhJB
wpbq7yrgBBckgKZBR+6uDeCqLjeDwC5wwb/+wbKQuvvMBxc9qT/C/jAq5OMmch6E
9G8nwpQGsdTPqzUiUG75GPNbwZcYX5QnjFnvCgPPCxAPNDNqYwVNbCF5qYOGLz4r
1GteXEzlB6F1gRzad+U45B/tFLmK5Z1njzmTTvKZPx6nHdsNSOp5+bo2Avw9iigp
QkpY2dW2zXsE7V1MTMwIvyTMEdZlXUS947dtUuFUEWGYOzFYS8FDaXkp7c17l+Cn
BgEMY9z7O47J3i+ZK8Ff/O1jKjAL4ifycigJ4A4Hy7ZqBYiRfoJ/nQkepL4WKy5c
6vo3ZPtYMQstiTrVNlAnJK9Rk3VqZnOkXy81IDIFDalhqT/jKa3NUuN9Bc+doOMv
tkBoDx54+uMVKCu2KrsNxB9Kb4j2DWlvksvAnIiwfu2qd95K3lqNb3fPSe7uPrhB
mZWK8Dn4+c7N85QxW7eUqjCU4XpuFjpQgQD4j8y9eXvC1Ir9kzHy8n+s28OjFSIV
apu3THshXxQllpZhPjCS+e2BRJn/AR27bXMxqNsK5MWZC+6t2r9NS7xdvu0urJNs
dxbcugJKGmbOiEVW3PGHLxunctQO8h3xjgsNOrA7WLfeA6J4Hb/myDsT2q8lY4iE
te2Ep/2RtasOpv2vrXJUNXTaUlyiCeMTY1czuERrBcbPp3NGmoHZ2S+FQHQMAkoP
oy+eyKQoqE7a3cAogtB4d7Ax+pQG3vlhDpCB+GKutTxeEXsCTTRpmRRFtHNQre/3
dDBQQROnJ/47gjpLqyknJ0sgC2VAMNwo68KzCZmZL6x1OGfjCSBmJKE0PY8VF14u
BXU3Sb/3qM3m1WjvUowtZ8fmRm7VBiyPcCAD5/bLy52wGRF9sKMXx0RraTHcTv0Y
A16eKLgMwC57HhT6cM9QFulcWsf17kwAzyM/4it95yLb64EMPf50w/Ece9ID9QPg
r4YWgun9damhdosGYw/l71hCMzwEzYru2xm+rQfOOq/3ItC2XsMAJdab05FGCQsn
iQBTQ1E1jdAH5ABtdyHVP4yy1rAf+XHD57o5+XKXBfzems1d7jDutrQdsleF+P2l
gdpsO9VIcFTWyzywu/fggqdtmQHvx+FCcyQsy0XfN9wIPlh2RqAojE74KPlHf+tG
WFXX4b38bDb0Go3RfMv8cFMT0mrCPi8AhuKZZViD1Fqkppl+rA5uWdt/7FdtPYRz
D3IUtgDyCXJYqMXRDmbw2OUEgL9+aFl2GIwg0f6w4UzOc9j0fG1atuUTpuH2nNZF
WM7ehFTgHC+FsagjIc45MQZ8s+j5RYuPYoCnGdUOmGGekTVZgca5/yqGij0vlVI5
ng4273UJbQH91OHQWAeHw78/b2tVPPs+GMJpnVrAsAJf4O/OZnMcQiIUdgQcU0VO
FBGPykqCgkRYOAuD+2vlmC15q7zNnXHKUOVbfzyAQVkxwSttUYdQZNc9TiuJAnEk
97/YBCGTo60j5dTwkqbGBb3iyhvgwtNqGRzMTW8AAxuLJyrIJvCR18GsVosmEdT2
a7gDEnALwy2wVwagSCQrjhE6qHSYnpZMUEI5FTBegajtNi3WpaDbYB0fAFS1n3UJ
3WqrkWFJ/+BXRhzwQVsAfQreyB/krCkoCT5VBLN0WxaTDsd0R4e3n0IQ+fvmCsYl
ATB2ygMZ4ZRlliltdLh6yQrSaJkxviN23pU3DQN+PDsEwPAQ0vs54NTjXrurY0Xk
9VsunsC0ny03nz9xTYaTr3oWM/ndYSvHhURbAcWOegcKZ3Xt1Itwghg2UCtEIAPz
/OEAHLyR8lwdvNNbpcE3MHuj3TCd/JkOgcOw+2gfEqS86XWPVwubSdxp9ZWFA1/x
Jec5U3BkMMGPLfhpvybR7L1uxcOif6V0uiZq4aIyk2tYIfr7FCwhBOH42l3Wz/uF
BTywtA6HDLY1mV5WupJgiRS1VVbWajyz19P17eACwyzaw4DTuTiakgCzQfAa+Qfp
9Iw5zzZlXnMRpQ7NXPyy/mPIRkj78+z4mjCJFsmYNYo0n5VyaIxjqfpM9juqMMk9
WzmrieXEW6BJ+eK6qADmuXnBH1sRY/DzbkLCODmdYUWrIYTjGs1Zmfddxm8hKkHl
+7kG2Qy0CatbEvyZwwphMzJXoZ4q7U+XUWerczQY6MKjCBl8t/mlqtI8bAi6GXv9
gRGf16fUdmqpUW+z6A4B4dwNNNuzBRWGrkCYs91VjY/EZgp+lFBkJnnIDyEE3M1R
I0KDxDfT16FMG2fi5s2UtFE2LAsgrKZXZAHw8IsZICjORekOk+XNbIzZX0mk//th
rRHIaPPQOvWDdXjprc0UVkHZYXM5ypfYECSLpvgw3jYKxt/7Nt7qVp2b6IxetZPy
Zncf9YqLmC3Fwxk372wJLw9+0ZWtOk/UnS6B9oEwcxrFnnBUTqtoXLV8kjqciDeT
bM/T/Sf1YcMEU00siSPzvXFS3i2US4FA3l15lBuukFYx+McdFGO2GbBZ+fYGuP3q
7MXv7wZRsfl3rnIFrVDuY/bJ6xVgNd2nh+Cw+dNg7L0RayZmqFFjehTpwmt1x/Jp
1Aqzw6FxECcBY+MAemkksnd+iqGjWgVuK8jSS0eqdMELcurOy4uU6X+62gmyIniX
GvfkZPxgvZtKCN0FxfKw+1LSdMSUEfJIb+q5cGo6RLp3XuDFLzx4An/82P5uLQTf
wYBwYXf4rx8MUa9vOjCMB7ZkzC/8Q7tVmTqwr/u6fje5KVrJ1RmMjJAiyVmOH5e3
DJMBXQTzEoEgA4g4ghjqlCE6VXDQyeyr5pypQwcUKisbDPLpuvisjiiA0qDIat/d
MQnvxZVzRXAoblzjVY/g7PRUqkfQ1hqf1K0z1SoJTL2ZI082s2c/HQPBAZM5JszV
twwlK0v2/potCiUooaThQKVj09j/GrAII1pJYzAeADD7shm97Pc4df312NGF40MN
+2kbewce6w7y1j6cvSL3wtVze2B/31IBjc0PSbgVzkw3OkgxWvigiqEsiK8YzxXb
ylAkcBtzWqtJMRZEYnXOPUKkbd31w4PsnZ//gGCfoDRxEkUSPF65LikB1athMXmt
kTcyicos/mm+abLYpQBV8n3v+lrJpxuXCtE+qzGK6Adf9WFLd6PsbR1OLgCFj5Tz
T0mnVipAXtiuMbQtVGRG8zv/gHpJsG+pLUuixrxncfvybX596JlwzREOl74TqsGV
a0wXeL31402pxRYYg1K2ud4/XMHoSyYoqbi042mseRmt1IFJ00gGDvP4TaR22hZj
tq7y+cX8WNfdRVM6tde0pMUFE8SAjdWXFbx8Z3ZMI5+bTZKr5h+jzqrezH8yMnvj
zQuPLugTWaXaJnIHYy+zQ7eGr0vx6xWtw8Yh/mUBaXAsh9hElGfrJIOjK0c1eReV
6ru35AHNd8jrh2RwXOcudjdYulVDySbQTdKVm/x2Zfn9EDaCiGLZoG8Jz0SVV7tK
xHRjDxPeLecI6KQHyiYHXlZltIqeeiNKLFqN3osvBrZLuqmTyjQh8wyi3nNfvwLK
4AUAJDcALDqX9R6sXYMybVWhmzPKe4vft0wqe1Twyrjbu4FWxkDThZgzUwvUBMQf
86ddnkP8SKQHwGXSNyzJWpTkMliWugGhvodoact2RBTIgCpAjkc0ZAQ2nKHKxwV4
h7YzWItu8kvpBvrI0gucXEdATuKm0ZkX1E8jK0ukKQ+Amkh2HooCGl8RCoOK720O
BF3eMjFaZkiZ8X4KyKlFp6IxBxp+JSg4tyvxbxYfh+iqN2iSBXgS7ejwL91bXK+p
wd70kuJPvn4Fd5wCo+ZNV1p7Z1riwdnVCwiP1ilTz2tW4pjMP/9Y+GXnhlSTd59D
Nj0oXOGjZxlFWwSDWkuSDcSL4jRgueprtH2RpkYVMpxmCP49w+vrb+7yFXiL0jEz
NMMtm7a6wgVLqzD7/zlICZyHqVrLNwhhrfmO6BPuvq3ycDtc+G9Qy+9IuCG9V3Ah
/in0T1TLVkikhnX/mOpeTszrzTpUh+YNTnlWNaaabNu8v34dwwVyDb8c64S1T4Qc
4qT1MeuZcUZ2lDFqRX47UwIn4Q34XrIlMhaa81cG3wrDTD8emjOHMK0gXr1dikRQ
u8oBQqz7ToNku1+Yc6rSTLWLv8SvKHabjSAaVAHJxZAl9VKtrwp+gbcZ/b7S7G2d
PRCaxl4TGgOa71hlx8fYfJBVj7T+0ErdU6XRrXgE6axnUpXYt6rlI9oXiTgBMu7B
4LiKWtF8mmxlNl/iYMc6lIrETuEbK9gRIkzYLTFy4CHc4on0BeSl6c5kcuXO5+Fq
tOfbAJf1Qh/SVA6KRGS7XIlhW3HuBNP+qpXWZetgKardwxjrDSqtPSeZ5GhyukbT
inr0m8cHiguJTMf/Wmun7MtvcY8fcjcEI9beh0lFgTxrH08jhQkVCEsXsQEkx14e
64w4r3e4RnZf2aHdnZZPyVzhrQgS9DKb+fgUhdL+DlMym4cfqRm+1E3TCEpOg3E/
RocO2UIt9c2G+5laFrZcWrd+8W8NVySW5L2aIhBC5koG+DCgD7ygOXuDTIg3VjxE
x9FSYVgPW2aWvaoeo3taCjrYPIBNIbkXqpelHIqwItOuig/ywTJuauDf4UY4rj5b
lNyXJtlii9I8bo1E1N4PpShFH/tY6urQsVAwV6VSocGW/1U+8l6nWKancQ9LxRCs
HY8w+SCS+ROFQeqsar3hf72+NIz0uWicV0Rj6NZRaYaTsfo0zu23eP/lKEJbRCNh
B7kck+j5+oUVgyBuTASY0e42y0VhYggEgzYJJAagomrpZDUaq4DBFSl1lWj28cUL
9WcAPi3MWBV0RKJ/zruLw++BF6AL48a6jV+CMGxPAFTMUByQWuG+bDcjAy6cVNXB
+GcOH9ylOiUOD6RiZyeZVWL+GS0bK3/88nYRfAbGb5MWeqdG3jiIx8W58H3QQkvy
9HmSqtMW4Ja9uq0l+DM9Snw1QyxrLYAXD74ELb3SNDcKV1oy+P97U/38bfTGni7T
wuQQDJXZ06jqQBCR/3Yl6iY7fxQgwVtzvcubJITTDlWTopWEEVMePmkKxFJ46v39
znGXROHXFp7723TOWj9/bSd3aO7V+IY/9nopKDP1/+A5DpI71GUe5VTPRyGW8xel
QkuT0myavy4i0hrATBq/ngUAY6N8s2Xh8SJ/QZZEaPTQ8XwEysgjp65YANRAi1k9
hFaZkcrcJonLSYGX0kMMqEKMvtwk9Gq1zCrBzBkCGzpDbMmTbUgWMss2ZCzTmsWC
WK2ImsehSpMgM+Q4Ky/P1yWOEDuaHwz+yzXfz6xHELAi0nGbvqXwVKpZIaIbeijA
NLL6/o/GGQIMoNcT1Y0bCsihx6pWINAWfDvB/4VyEEQYHqmoqMmI88R9B7rqPWTy
zlPyu7bqKCs+0OyXHYa+idFw0HvQny7NcnT83Ve/QyCoXb0ferckejPH2f2+9sL5
UXgJ0ZSgpZaAnJxasIADPF+j6V1h/oWKLpJ5akWdlCPgtIp1R4x5fptz9VZ4Zkih
e8QfWQvWHmptvOz8QQx5Cg6MeiSeWEoHoDD/GzGnBWNg45TYPuacCpvY2pTv4wd3
nBgXWmnTw4WxGXCHDvLu0mFOoP2lUYznZ+4QLUzxCnZkKWX3LWjnoAJaOopykIDD
YGywBgrqw/aZ5xpf1LuDWP8MddNG+HvFnpK8bNL/pSXn3z4m8Lis5IyqPEe5RTso
hEVnxxYme0RuvgRQqN7M+D5fZFbo/QPXc6CyC5X+RdO5DCWqB0v600a/CYgImvIR
geTAmiMgp1r1uIj6b9Fzomnh006XpTNP4IrfQe3c6WqMpnhK0gb8YSga9qhGvn/N
uohAu+Us0aFlKwUN5DOTW641gB2r/tamdH5ebYaumnYAoWAbfb1YLyN7qzrp3ucj
DSwd1zjSrtWMncmaYnKbiOoXDzW9QAV/gCWG/A6DBAexxC6i54u/I3QNJGxqWfQZ
Qx4QpNOMMZbZz8Y3XgOs3dKaayCtTh+H9kGmLj6GOcR2iGuoYn6zzw7qn+lpiwnI
jvNhHm1CdDBYi621x3mO750ji+yOz5/HwPuK0qhnfmg1libNJrqo3beDUMMWZnHA
TVcDCMxDqaB6Q/cE8akR1uw0DlYx+BgRIxxQanhaNN6HxOOTl5ehUglgsON7wH4q
Smqjl1OD5/ZbZyskSyu+NiWO/3+id7cR0E3GHRmQUXiMbfmWcsB+zAliVWoUdkPO
nu5rtlVo5S9HN1oVQaWwSokCJvsKZskOVxTyM0JaNm4txYCO+Z0vWTMhPN4zyr3l
rheAlnJQhw8VeZawW1gO74OUVRwxmcjGJL+m6Lea+eSpMPsuaUIHv/1c+wDcRoUk
up2JI66BQ1CxOh4I7Kc8QvC4L9ZJBcGZ1wo03cWk6TffHRH4gUW9935NUUyRw4IC
+FI/vaeammdXnh+ogBWXavIImFKTBGDoiAnOFjwQ7dpUOWaeXIt1yuOZ+id/d1fm
6CU9CkwR7Q3JZwlWpGdtgOr9pX1gaFrQoNZxvyb4a2wLCxVz3VsHoEacrFo3xnQO
EM/qlhtrQaLwZH+wPagvye16OHDPGiq+aLx6xFjyOU2TfGgoYT9JN/a7n9TFGd/C
FTLGcudyrjDit/VK/8ExSbCaBSXkBdGFFm0qKVoiklsgDuyo7KEb3SlrjUbh2uoS
Qnh/yMr2oTvku53kjftXNy8Rkq4sgcmPPme2C3jq6Hx7TLoD9ozz8zreew++cC64
ouy0kgaFE8D85RjvGvwa2dL8vdJ/ZEXJc76Ofv9Ak40B/2ES2sbX1Hbd15zNFZUn
VzWVlGnz1nDWRVDIulJr8RKxFStU1DpyeNLzzHUFIpmcNvw+MzT+Bp97zZkjvq1S
5MPOCTko7uf/yKvox37oTtT6R37ayVvazMWV+k/0dXU+MQRLAZuoVNN23Rxo6aBo
3VESfyZI4EnfgDn6SUYEwZUyzbQLlV8LuAKru0JnQn8J3D5vRC8nyC/d1I8mUJ44
ZXdlptH6iXZVtkWtt1ZOnnIuDoWw0/ihdfMYhOpw8FpAq313+EsPS6yyqCqiMyY1
vCOq52PwpVpsATJ55RZrb4DbEXGjtm18ylwCQxb/2+Iz+4I/ZoDSSVo5m/KOV5wg
y3kwIDlh2N8eqbUq4x/rtG1UPyNd9urtNkpAltXdxuyHmCgAr0KMCwwyYIRhHN9d
QvtUdaqv25z7LZNiNEV0/bGuBsWthadt4RiqlyE42fHk4GBSl881LShBcXYLokYl
wZeolV1VLBh1yzP27JoRekxCBCBgAsGyhulx8bJIHJZcS2O2euVFGNk/NiS6lnvi
FMa1PSbA7dx8m8bnLifttALq9J4Ee1Z17p54BRUGBIdCNch8PFbuFogfIM+/mtCe
V2W/x6cvB57tvjxSnO0/TGvSmDaOJyCY3jF+KYBW5k5HOxFGqn4/ZiAVMT2nlpcO
+75AOhBoGbzx9Se1sO6NDW0+OmgcrzjVaoNnKUBzDO4W39LxFoZqvm3y3uxIeHKR
33did5fuElN1rdQN6gE4j3X7i/nTsNCaplvT2T2d0qX279dypT5ZzDywetdyof1Y
OwDV+MQi/wgVAFI6VhG9lyEBBgLqb8vg26L+u/oijUByH7FCw4k/JkmN4Tizs1Ww
xY0wIXctwCCKF4J5VJVZSN1pynGFhY9BvkBfnToDi65Org+eDpfe9k3mNuZzhlQc
vnV1699FCGFf31AZiWdO/ZHO8o3p//S23b90fTu5tFGwANYgHvfLNXAVBPb+vAe0
KJTAUdAn5fjm1XQYnySiry0PzExdCxSkGGYFo7on4IALv+vgLwY2RrY7+jqg8wo6
cEeUWN589ansedg0LlrUTYJ38Y5iPyZJGIpwdGyawgLz658THOzsW0YBKBopYFbJ
bj2kID7fwXKZPE3UxPoTxjKBKCOcvRYsO8EUkFinrpX303j2SqRtMJeWFkIqAQVT
EVUuCgl2YovpVz9zNoRHviEpPe08+QFnTo96nW9Mb5f7bPVI3R8T0qOnkC5ovD7V
7BAPc2gwSZlwJkeHLQhVv2Fg807ebFQ8iRt8mWhqRr+RleXzg3ryTK/GLZLWcObq
GcJsvM+nRq4n0k3eJFkmmhj30sXv1ltHtlKC0xR8Ieham9CQlgcna42dcWqY6KzI
0eOe3OHAHpU/mXj+UJROIRWt9AkedMPPLGrhJz2r09VU2e6qNeMu7dit31P8CC4g
2pGB6AziVLxSDxYGbxIEOEsoM3Y0WNTgNSt5mtG8nGv8vlr7vTBGV6moSjKmVBCn
pvoc6b072qMmlvSVt/s260nmz+r6jp4zPTFhd5+/Cqn8l7d5nvg8KS+VwDbUcQV9
/kSDGW02k28vVHAyoqo5IIysDslpQygkeZhWb1OL1cQ72ivjW00gaYcyCrCkzx+a
s6A+0raApHpgvOceCLCaAX4QBpOxz3wukhmT4LDivL14TqT9aMq5EeEPCaMnRloD
i6gB0IYrgjvAJBUjr4OEkLNN9jDhkY1VGi3uGxo8G56r0+bVOqDJCR69w002bdnD
Ac5aDMtj3a4dyAKyjiXI8uvAg5n1WN1pWaJTcgVLntiamq40g8Y6mogZi5YGIMy7
d1gLLllhYHFGu6swpY7nLNAQ31pKEjRFzq2M91Altco1BoWZV0wIe088H+wQaqBj
t6dhNsCLrsOUd6SZ1u4wXrk7y2Z5q1YOruhvbtHKEKKwWrQuO9LSeXxxT6U4HU33
sruovgZPloLFNO6y3DesgP41LctsqPNuwJEE49fUJmpgwTTVPCWwiuOyZysEPkIN
k8vv21gPPNeO78ZdKMdJL3NJqqP4akrO4uW5uVaD5vZGyAeGoLPdXilx4+invuZe
xjD9mhpBsuqi6KGDvQtUbVWsuFAZToaDEprfmvq6hj99kU67U7Tw7fVTuTZHIsRV
0bdq7oePpwrG50XKoVQnzPFsi6ASuM3NS00HTu5Oa0gldyo/ZdEN65+5HoCsl33e
rmzsfL00zg3p8CWqh41cqc284aSJn/cWrF/1t85H1cCOTF8319ort1Jqw1AUmDZ8
uowR48a38lWT7XJJsdLA03w2Xne2bm0j0eQcj2ZeGCIGbgGApEXcTYi1iSlKmLWf
z9SQhv4C8j2AvAW0VcnsLzS2TKh9yWEAKHp4p08Ec3z5pQj2Lw0FRb9ldc2g0PFd
KQNVTY4Q5lPFtRpkqTSOEbFHMwGOJpjDqHzHi5pvoThuXyyPloLSqrHY5sOB9miO
ID3PVQfWayJVFq8fxrs5YLHIjyOXB2beLcq4iubKnvNBPkQy8Z+73vFlGpxGkLy4
2C41t91V0n6yTQ4s46GtjT5YfHqzHQiwLf5LFQ4NZ3qUjtmvWz+MniBELv88i7l8
IBeE/bZH+jWWsGG+EmbCtutuctflMADxmNRnYQcytu1jYs81J+sOewAo6EsdPVr9
VsRqgNgLDjCR2IF4dsICQYECC9xjzGhYxFjhNEQHtdPrwp11nxO+5JDk9UpN26rG
qv9eQwlJHMV/TlsJiLQt7Iie1Sy7yunJBCndzCwI2khFTelREgjlPS5/Rbmf3yDc
RQGi4Gg1ua+eHMdbhXdpKUvs4Rwn7Ne+Z250EEQJq9wc22nSRfjdFa9jByVa8OPw
L5OlmWvZdqh/sibtQC4fESexNFSnL2IdSo3MwWaK/3VG/bUVPSc6CHSy8mWqU3Rl
eZTsvpCnWhk2E4Q9Wr4bDxyjibLTobYj36q8kxA2iabsPwoWK2KvXXqrNxk1mqP/
Qf+qVc5agIfKO77AAlnbmF1ciV5Ip/gWbLrZ+GOem2k2FcMlG5QjMRryGjG/NykH
4RHV9rbfMgmZoZ9DttPRtRAloSK2HO4aQu9Q2E0etXAr45p06d1rtMCXRiXm8puT
WxifLkt87KkNelyGK3qJczpxeNIMJHR5pwiegs5mfSXyfQni3I8lfN5HTflLGeKs
TrIMSiYi1UvONZktNkA3cJqpyesHyab8DzzlFxhOxHy7xTiTsHl1TjYJyskyiivI
6qhNIyNkex7FwlzYVx8+qyFDq1Pc8g3KkcPvuWDfPjWkGOGJLqFiYCXc3p8Ll15D
KrRilXsjRRPQecrTFIqOjG02isH2tGyW1dKVozq/ap+DHr1kY1vczcuJLt05sVdt
ALAcb2GFQwOy6THsFwd+Vr7abMS9Yv2EnbgWcJSkjWiwffZJocU7hL7hPKJDcM9+
gHA5RLf1qesz8bDblN/+psHoAOw++0zIb4yZMU19dY8Rfdggmakh4NnDSsB4ClPw
ps+D5X/67ZrGsyNiNz+jtSlO83lAQysNpCitOdziDSEtDPBIczIVNGedKml/GBfx
1FQtD8/cd2y1XTOHUaPTepICM3np/P13MkdgRVvg3S3NQ+JJhftTex7SNJNADqDZ
0Ej8RnxX8Ed5f+s4EQtN6/LKEC1K02xnfA1XT2dI5RYoGAowzqKgjuhMm5GKmci7
awe5SPjsZ2uXzZ/cLQdCR7RjSb5kjBXbhiwCs2Txf48+dDQCu9BlOJ1/bp+D/5TO
YhBf13OmrP2fXmkM/3jcOQY+LvbMvWM1dNLHowmI36MgUqdRF5TJO9/u+QKAYRzY
qepm7u+7ABx0dG0hhnillFpbVpRwa9RFbG9OHMWIhGmu7ZwkAWH/B4d/9cPBUgvu
PuLEdbfboEPWvN+3vOUZTcsYUNpNGYfiS8aKSS9fd2VAUc4P0Z2KoDKc5RSlpsFi
9Az4Nxrc8XeAkI9fzKi1vAA8l3UNsPi6PmC3DpaQcO+RZdMNbsm545x+6AyIk+y9
cRNhadzmfsVnVFfCZR41BTfpsZrv9hf5WSRd541A47zF+dEhDXl0OpDQZSbEM9YR
uIOi9FhjoiPxTxIyGpxLfy1IhxzFE4yz5Zs2A6YPwXiQXjHb9BUKIgaDiKgyxWr1
PwZX59utrdxn6mR7Ot887+vHprfiGhYZN2SMSy+v7Ln73+0IemKlwaiz5Zi+b9gK
y0h9Xz1oSgKyWeTWmjlcw1qOHydmAHX+9fTtbtj+QhSBps/CpaV4B7BysILia6Ks
0dcFrUCSzEEYG89ALkp3j1Pz7GqDUm/uoMaYBuCjL3n6ETGyTIpgDeIj23cFgiiq
xM4pX/d+xELtRTAD5PlBZIY70mWJ7vJ54JZc5H0uRcMhYQcWF4yMng4+MPMKhNIx
wzszQzLttodaqrz+L4OHhxZ5wrOXq2sQpZLZaogwQfGoOpGNzBrCdkN8rOLsv8xm
P7qpEiQgV7Pttt6NY3p3/rhxkbfM3yRjAMMBKlS/Sc0xPYkgP9jf2K8Qf2et89Jt
paOPMf6WlUnk4SF5GpC3Gwf5RGLr7ACNN14J4HSvmrRlopz6FuJrck90dGSFtsBo
i63oLOgEzd80fpL9Qiqp5CCzaasgboereN5dkgvaiVdzDeqTdyoOqo7FMKE9xFu1
JBXr/wEhYXfkFXc72afhdxMdiqSpI6BWexS94ePXQSzAYZsNz2a5QtTAW5kq+FJg
dvF05FxEESclMcZGGQ3x66Ym3ITTznZYIXuIKvBPEM96rMYfxfT6WH1ve2lDdqDP
QYE/ePK4avPSbokv2VEaTDJHbKY1NSHqKWJq2U78Lt+pI5sNe6QlZUBdzbHsyqaD
Az9dbJe5w0Z8t3VIPO5/HRaCYWV8na1yPRvKkzYu1NG+jcpoMWXIUCv6jLySmxh4
eKKLttIPZwAx7Lf7spls1fo7jlpV6cBiV7mka93gXZ+S0iQCXmw0XrJ+AZUoQMqS
go7Tb521rcjbz0S/oniii3cD44zXN4n++RJnfMTzQzcZX20iNau8wanKLbMHzr52
FMqDyfNyAaCjRD+fqr/KMW0l4U1J3LKy3Ieffky/CMUCrlLy78Nk5Z4Mkrd3gevG
OxKY58XZwlVfq2LWBWQgRPHsl8u3Bs+SYvSC26pbQjMzNj+PZKE69F+MUjkS7bCD
1nNKVV2y/3Lj43LnYNlDKe1jcBmLDd0eQxMLD7mtUrx8+O//ycbyfx2ZmCsp4ztd
kWa3ZEngdatIqgqnHp9/AqT8XtrvhKsTyCVWDnXEAQT8LpWBvzGEpcCGXzPI8yQj
sxuaFBIYzQ2OzgIjDtYullUqZB72GZ9wKCligjjxTtz0vHV1BSRs+rL9cXeB4Z8F
Ls8B9v4uyBPFX0LeIF9vLNJ7RiCYYXWxnaHyAITGABv7ViL811z8yJ4BHXxyr/ZE
dHOvwapJnfEYqU8zDELOn53f4C3Vt2lkvVqRq+rtkfxrypaXWiD58JBUPmrrzLBn
qexgQ23rQmNsf+ojA6u9xl6S5jsMTqj1BzJJWqfLKEcM6iAv4IGM8tykrpq/hWK6
sIb/CV6I3l23/Ybx7E+O6pGCNy/UqjtAO8CuVdGFIHz56ZC5LlLDd+miZBx7X7b1
EUEL04x6yBvJZVzbe8AKx0zdxGyvARTJynKSQAQNnCizDp/kVTUGxClO9u+wC1Wc
BbhsuHDGOENNm+KChj+67qkglFkLt07G3pbImdmkn+SkGVxI17ZA/qJ4MFMUOso3
TGkVR0OIZVIFGGej6GgHwDGVqj65rnmDQSOgpPfKnKzVOGMSnUNbM6BjikTHiNSR
4nUW9Z6NHkQsfGT1ONlZFMscSV0nCRLl0OzW5wMXY4UDRlO3bl8q0RFP4X8Me71X
G108vFRCX/AYA7gjxvWri2enjfE2gr58AUIVhhgjS3i/JK21HvzHeU+Y+qqIc1td
f5bAiere9QTnmyyy2UilygUWBHXocWL3rVhHvSnS7GuKOn9SJzAOsNAE5tMg0h8F
UvbNDrb4pC7dbtbpvDrrmRI7RnmPbaSy1rNyer7z2EcrPscPIo/nw6tqTw8Xe0gZ
jjPSAtJ9mjsspVy9dYk2VBwNU3Y4ZkfY+7kmWk32xFWib44Q9dNe0hI9tFvbJt29
YRQltLXC+5hG7ygs58LBRBHZPY1Boz04S1M3ntOmAvcF/Ql7aMwAPVTwzIrSwd1A
Oa2SATFEWuo4DH7oLt5GF3U9kE5Jb55qGK/3G674xrsYA7C33F1xdGS+RP/lj43p
P97JHfs/rtIsd/SGfsXjzq7xarEuKC850d3VEhnBouarohyUUXtox4Z042Cnt09q
hy4YougUamb7u3YCiGbwehFI48bmIDusQaPVcW837Xv4W1aR233yQ/vmeAc9H7SH
aiZnOp4L0tELNqXWlJDb+Z5F/LNv29jAJkLOHVTlQnw+jPWzkHEayfurVXRymhRV
Sz2AE0FxrxI0YLIAoDKt69s1mt3NV1CnccNUvUJqpXN3Mg4v23VCQMtfEaQ/6SSl
pJzuprY3U0URO3rFiUAYGsQcYY8o7ksIJYU+FINPAKQ1FJHP3ds/Ed+L7R6sz4dQ
OGTAHN9UzbRrd5/wAk0kqjmi3csr1r2+pYCjsPio+rpuKt+wgREq1UbkhkNaBJkY
zjHhwg/Q/yIs3sBRJG/A9x+dcE3Q3NjJkaYITiprPCiS+ECqhayenxo1z/l916JR
nQrA0BcIX4wkx+vvkhwO4z5o4gFWfZQuCGGxOo7/8EmDpyF0X5HsQ7w73eDqySWi
chbwg7q1zWNv9gK3DlJfcu3iLjZvsPJuxRmOdbjCu4DKsP1yFiS2HH9sSk+AQCtH
uBb/uaxEuWRAogHpyVayWzp6Yr5AZp3CWPg8FPOUENs61OLvpizcMWd6xeZu22mT
lzkLwwQEIbDkUy7lkaSFAvMqH374hs+USaHz/+d4QvWDRa7aJW2vlOVgB4Liuejx
FV0bBQ3IY0+Mkkecb94tMG6vtsGWw+ReVw/oHYqyVMo7IvmNlzkkaPk9ogaozGtI
si6F8G6YH0jaiijmZQcBeqsn+dZTv4tmOM2CHAoiiczxmlu8t58K8RUvIjsTZfup
s5JbYKBAmnnw3UQKvWb0VGBqNNEXsXN7rbjV4BDxj2cJKTC9Llvfs/ooeNpG7+RF
7shKUFN0UT1j39hnKXQfd/QQmFtaVXKsjB311V2DXzSJq/HoOgLnhx6hdB/ExbyX
mvEzp8euFgh6/mb9z101P3EC7YwwOFNKVNqGox7LYNrCuGuLWc+DRalUyV5uHxDi
6bS16HunX2BL0vsBeG1+rXRZFURiF6ji9cEkRcNUE27zZ8oQLvvlCD5PNxj2tK4f
JnuRcu0If/CYVMTyYLQFg/RRJ89Sg6qfFjl6OuL8fN9MPIYQlwzPV2+JPLMx58s4
DkjzMAx1vChDGYP5Z45FCIXBFBPtXB8/0lc0LQpdCNR85IcZKRfQMsZcWO0YhxaB
5f6Y1+D3OEjUrlw24xBysknVw69lh7C99joyKafgTo64lT1WiX09GSt3xX0/FlJg
9gIkot8nX0LFytDPyXaZbghNWLCqdKPo7a2Nm4pslCV8m40lcrp5ZwaDR3MEtnu0
5Q7TAoCK79XFQOrWDbJ/ZL5sc6WrknsYWNth7kVHHOLYdh6njfGZPTcVHvg0UWWe
ijkkVzAxS4CgWWN08GOiAYSVMJFIwOatuCJ9aoFlH9u9+qXQ5cx85X6pmAqknvvm
MtcFlLL4MUrfsZarKCbYb5tfEnkAO7K1BH4qsQ33IWfVQ4s0rRMTNrqfOyyqvuHe
lF2ZhleaYvZQZ0CbsCGVMneXyqKwubwmngp0nKFLp5ToRwODLMa+66qtJmtfjVX3
uR/SsrjPki9Ij/GVxswG9FJaNIKZ0kXxLRiWG/fEUrf+4LsIHUDrc0mmcToUpC3F
HrbafNA6BE9Hme3SBtLqFIyXGsfNcfsNWWhlzpcIAlqfJtI6599Xy8pw+uk81bn2
IJsCoO6g9FH39fxAucWC0sPc4lEp1GsDfV0MAgIQcm7IITmwtknY+5bjEc160wYz
MHgQuoSpWUSE66lkg2tVGyRGxNk3nzLuJ3gtB7sm9WbVCTdkXOVlatVIhepjO8z7
zfipyR2JG25a4HxZ19r91e/JXxWTZujjSrorBNxCPxorNPpx8nZYCohn0cqimR40
obNMa4DAr4ZcJEUytcRoyLp5Iu7iNu6xFIFxgoDsXmDCUrJiBqcnOG/R82snqC8V
E2+l36ri3YtKM8LxGyzK19LYwyWSH/9ntDY0/RqoDfw6uMg9H4x9oDVq60cILH4M
LfxpSQ1ydeZOPE/V2s9k5DAPydwIkJP+/N6X0qua2wBNJJCKOuWs4DQ/NT+mDOp8
ehAlwa3C+CjEcWsMYWLMlm7rxXaIKdBOjnBLyXM3UnPFxiXZk1L93b6dmKOz34+a
wA1Lg7UlzlVVsZ9M9EBNB7fnLDkEq1UfM7UOHenbNh1MOn5l57LhCkGXOo93aw/4
Yrj4+EXnKbOlr7flQvH/p9ZbgunQ/hbe0uxeI4YLELXj1cIxyuUP3zt11OsxxtLj
kCrxyplL60QHOowUi2i9YLIMy/x65W2tCSAyr3+sOXCYVFnPfrJER5tZ4yuP6lDl
J27ynlGn35iD3T7eamxLdSCCm6geQDsBpmi9qplMZ69JEZwyIex8v8DqNDZiZ6a2
TCPq+DrVlgkK6bs922BElDv1phkm6PjeFXN2W+CBnAzSnHBA4Akepw/DgDdqaRmg
W3UXwnTvDL/c3AzJqGkzYsFFGyh7KMrIirg6lyeiSYq5DOeFk/uhHiImlw4T5oHC
cXtWH33tGLGuon3w27zY/rwzM7w+9xXwDMiQ7d1BhwnnupbyFxMlv3HOIxet36Vp
J7cwu0UF1o9Fn6smWu54NOWu20Qo9sTSoAHcHaYtDYfu2aaVc2cJNo9cIQCcxPjw
dV3TXIMdhnU/KbKgE6EHxkkdp1/q2TBOxZ1oPPv9s08bfKlKy8p3o61cerZlsWCs
Z2cmjboUHkOX3fve2kmFrDwY3Xiw/CcNN8jfgZ4XALfsLGtCyN11+mrL7Ji26cE+
rYZfY+hYAlV1eAeGH377Al8dkyfzXtPi5xFdGcnMeGdjj89+nFU/EeHKoGg/iety
e5FEryM04WYa5YvgeBHUH1ipYIw230n0TgWdw6HeVZZl3u3tP/xXdqWEb+81CteK
Mu78HqDn1Qtjv324Yz5E07zM5BELR8Q9P7atx6ullCQvTWXcBnkb570FQcB/1QlJ
WBUXa19wUk04XzYP0vmzkA5gNuZ6SwNlFf0aOy5gPk+v6VTzQUuM8o3N91iHLE4w
chmzdVq+nkVz9jON3i5arpyrN0TQ2n2wCSNskxReLn1tp2jSJuwoA6Kv17gtTCSw
T65m6DsJXTqtcj7DmfjpxZUjzZgUus/wXBp4DNyt8RJI0swI028GFaqjYl5h3Cgk
6Wj3cP0MDrMiaFX+wg+2GPDeCmRoX/V30jA2MtCMnJhiUIT04NbyHW6eJJfppNzt
/lpVv/5IJ4sN9+/RR3fYoyK0BTHltiJIe9tEfbDh9QoxEeiBuRdT27A/8HaYaa29
MBEGE+2BffwA32PLuTyz/u/8QIcnSWGDcbJi4l76GV2jyTSbhMz7qiGTsY/4Ovu/
g8OUzzsohNaQXlAZ9L754lbSb6xki9yXwTdzJpGKDNCPK8zrImTWdEBTgFwPwQ8G
jrKjFxoWusRD4cfItoF6PFgpXR9uPtX7Zu4DYPktMrqX9RJzxUPzKhgmiTdD42q4
unoVH1MgYtbo0Ysm1rRlunjRVjwwQy7EswxAyWWMpamTQor6RYgQh44SRXIsAxju
dqdPN19YsHyeJMwknH6DIRu4rPV0pXciIFfCGjXlSkJPCl7CbEZ3YZuUT1ywo5oF
YrRZxgxaY3PLQllMZNXataYuZFZ7Hen4bMvLOHxhD2GTmlySh+jt0vPfuEHPAg1U
ktuLaB16yzAYp4m7lDZasIoTMoNyRYCKlP43/7DnDjnHYPGmYH2Ki9jT8aoTQ54u
Xd8lVEbCynU1aKzozEPz69/D4xrY9t5HCMglg9IwJ/RwGLNjkxUo6THFLO/zkOg2
BFkahw5RnIwc/Fp83PwinBEyph1J9oObMp8LGinNLhWp4L2sPnCPq+qZlPGrEkkg
mvZC8tI06dH/LJ8G/Gt8R2mZOuLZ6SmFQhNEEvONn6eeu5N134lEc3mHUGguQxMm
Wb+jkQI8nRZth9Q06ZlG5zEvpjCQ3KHSZw3OOGmZ9F3+PPzh5HwkvOsyy8y/gJyY
ShqgPFYNaaUENAU7j7ukTdFPDCW595X8x9din7CVlPBNHDl0trMx3hC2g3Qzggji
ji4Ec1rpO4l/iOSR4K2fCMZoUbkUE7S9Ht1o2KaqFDM0xRnHOPUA0cHbY9xJe9BC
G1yDuzZHQLEFxIuXH6aqoP0vs6GV8/J/jkiFTlgRNHoHOLotqTgGqC2thyU9a4Z/
jzsw3wtbZAYRTrntLO5WTEjCxvj3APdcimHFNiXudszmGssx4WWwbSz+RI/t7GkE
he6/p6Ff152hkGKslnKaIjqoljAQF/VO3uquWeyn04uUOkCBg086yQXSzoaQnN5a
2+qdMKje/xd3ShE+oIVA9tHOidTLheVIgSFytdrBtIe3oPlg+w8bdgfe322jkfWB
SN5lNCs0NZEf8QCwSDIFbGBoxM8TfDLaRzKQ5rcWqxU6/ut7PmlCYCJKpsN7vJCS
0TYI/optBkqbc+UkSmQXnGKax+e86ukuXuDuDgXrlCcp6IoxAAgcYUu+rMyUrnVC
x4Q+ZUwcCJwKXdgySxrWw8vRJ46R5l8JvSKQS7rGRTUTzxaJMhq4h5Y7CvVZozfN
XVSdX3RQy/KlaVXg8zDn65ErlVDOdVhFQmFkhnvFPjpw4+haK7G5PVOyFAC5uOAW
UT3kJ/90ermdywUQGjn7lKTtGLORsKmKY+Iepq+tE6p/h240WaM4hjXPbZDqnPfG
p0J1Si/SHcXd9D29lRefp154Y5Nzqiz9fow6xbsNivOHLhTRURWvMFAYD+92067j
QbGCTZRnyRhvU0sUD7f2Xp8s6pL9Z7Scw58q4iC/FacKdT0ao8u+50rzvRrvCW+7
ElSQKaP7rhffoXNSQYCDxKflWZXq5Vhi7GysX1d/XutQrhZyDChYx1szgMLrZto0
YdAVNyUq4vIDjwPAFNZKP/uNuGYxvUtg5rufuYQNkBIOZ+eIv+3eYiEDdRS1uXdi
WKxGXrl5hBNWGCl4djkSL1WNgP+26iRLvctWoCwhva0d3FiBeOHR6mKwVNm7BL3o
YVC7nDsoGdS84x8qVCJJzW6d9FQzElo+X53nsMSFBR8XjY65Ii94Ie2oszI8UC4b
6K2LAlcRmevTbu2uLG39B0HAxYREEw8ic1ufk0Zek7ZIZ/8nIhGX8PtOYuFy6O8n
mySL8XtToor8qCLPWuPEiTEM8xhd+eYE6pvpzp4vQkQBHAtIXWQcu4CYRWgKSHnM
Ef7kJO6BuqQhbf8f//Mhwfj7tq4qWbfpFLF2aa5fITlI2b3Loc2i8DPWTbLnjoYq
29FlRf5cXhf5t4qG8wmmkvcWkCPWi+8cCy9uvGSsCZOXFoCC52XQ+Dydk2shSWge
GDWeeKJ+UqkTJhzUT5x9dIQ/cU2OEXHLOMvnR8wB+NLoLQrk6QDH3eD+NrvUzqh9
SjZrO0cTOiNDl2hNi77NtcqdN7IfivN1mB+N9JRMCOEkg4M0GaazetA81YC4I8PP
ZcVSMmX7woA18dUcrvM82TH5uvws5iXH++9H1mvnoZDcbSzWydhJiXB75FjQ9PQ1
lQQLt0kwq9pB31OKxLh9ETNuxreJRVYS7T8RQNt79gFLpMwasY/ZbzE8nyYekJrj
sblOvXqaBw+SLyojuZ6Bm1D+OrVkGrP7ii9Y+UqPWSKnleV4lbdRwKjxJhHAJbo1
unP2QtnMUlMp/wl53e3x3FjRtsrlujenNQPYlv+lJQagutUoOYasdpU3jGUWFZKa
WHmEStTHujPp5D0pf0bMnWoFuCOxjTdPkpfcBrCcNNAcO0852aOOfHro1fdJbmur
NFcE8pDOxCV5+mm/6D/6LsfsSKDSEFLMXI5OuS0VH+9TQc3TcNI5yqq6RB+bZ8fz
v82sPdmEU6ixKpPdhIObDdJisxXFp6WFQnGtebYmRay8FOaL9AF98eNIFsskvIa8
PpbgWQE+o15AdBSdA7MoaCS3LeBfLUXrQL+lrXZcaTualYwjZUGB67IZAJQ7ax3O
WQMg6aKN6Vu8InHOrEiUDE4Foi0UVCiOVVvuSNbhI5a+i92VsgX2MTwUouEdtxet
B8XMYr4klga92V+YJ0V0EF7DWR6HT9+thRq7Qvwi+8pPljUDG+aBPFHoD8JnN0cv
t76yNwcjm7eZdaHp0gQaNgekqGrsajkkjY1pBGtOcIvWR7n6JinN9Ug6cbIekXFp
kyDJBAF4qmJjaliYUBerhsDG3GyKep40G0HrjY/XcDMH0WfLsIeTLfX6xIxPofJd
UnkuuuTlMR+fq/nEQQFUFfoRilqswfL+v54m3p8MSAyXise5uXuatSwbusesmvSn
9m+ySOoEdQ5HYmyIiXLs5WH93onPij83P571rQWG26603qKHHFf5CP92i0NaN3qx
v9mLwaNVF47kpZgcCUSmcOKXpps19CRxpMcYr0Ac6Ur1ymEcogAA7ikjdK355Y8K
1ogaJo/nGN639PwNmdJBzqS8YikMaIhcNXM7/ezxV8d/Ff2JP6R1WLH4RgRcg4s0
FfK22LrQAsh37H3Pd5tve9vy2Xbd2FY/hwoVnlGUW5V44DWwpu1aZw5IVgfOJcoU
RDFG32KOlyvpqs+5MZ2mFarWJoHs4M+MM5u1/wzxeJEjhkRoVPNyhinKXG4rqr5r
jehUJ5zmLwgAf6YghzzyOKMmzZdHN2JVEAO/ay3SQNk4MACXGRPCjlGmlR4/1OVK
AT7eAp0OJsnfPk0lLJriHYmMx1hEUOPSW7O3BsZqFOrx18Uxzkm/BdyPgHRLurGC
Woxwf7av6vbtigaP2V7c9qR9PJsMuRupjrxASQd2eL0ZzqTSINpuM1dN/PWXtz9/
YAOEZFxgxtb15FS2/1PWMFPPPDQ4YaIPj83ebUhn9vaggfNvGwz/6/e2Ku0nn0Tt
vY0VnhgZE2fPm9UO9NlSPU9J04+79DSpzyLJVRdpsBJb361NlpYXhx6hMEjlzQPX
xiMgGA9/n0LNezA6TjGFJjCEKCXZTkZ3AH+867sE41zXsdg09VTbfvNpU7OycHAe
BFKH4z/Nl5aYZcYmvQR9MYiaE2BOQseFRIQN7FEiIsWOg1jLuuBqHbDj1lH8Zrn2
8+c1uYs+8IXSyZhic0JVPCRpkjTLGqVpempLB6LuIZonAgZDQ0qiy8z+20ZusgHm
xLFI29FMxPPBwt7nyWT8xo7hJtsp4+x1M2fXoaKBUn6L0eXete3YDjKBNdNTK8Y4
okkQdV/5EKnUIYr9Mknbxn0SQyfLx7z7NT6Oupnmd2iPZJp6dvt1P0jk0mnp7dhM
U17mDaPA1cLo/gAKozRIA+O28T9OGYc8RWfZlt3qr8tqoGsZSHS8gupP6/0cgiKR
97r1BuGj+KEiTqMjpU35FrG/mWvFLNJAQ7zF8T76hYkK96MiPzfj46rENyTOMEKl
u4v40wpnl3qkZ/Nkb/4gYURRIia7tWT/FWKyeUQNW/FdTad8dc5UM80afp3X6NBr
cvadtJk1vyzmA9bKNHI0rNgcuTiZCKcpP5AAOWwYkleFmF3yIV08sHROpMzaWhN2
We8jMP5kdw1in+iD9uovHhELodIZ/yJ+9PC41CM1HYoopaX8P6L8+FxpfzUPzsNH
K03Z/oXQJUyYmTgB0i35VSZuacTDo6b+Z4oCE/I93C0XexFrcoQQZCsqj0LTxrGu
dFpKUYkU+kSipzZbykiSf8N9RgI0lwCBTsey9UJ0EZo7ab+wJrNSwwgNjgD4yObw
d8Cr0xzT8psYTz4dgChU+zfD6HyGleGBUaKJl3okkanCASxtnDTBwYF0IlUk9YKY
T1i3y1kCZW7kZ6COaRVmYhCkgmPizbxggVUJvQm9peTn9lN988NIp5Lae5QZCvbE
LXWpZeip/dB2FWAVrQvNUQutQo4hy4lRSnoeFnWvMwavI5uhSQZYdbXyAHRaiofN
khTYbDIiZRNygzY3meNomwWDH7EweI0GgQvscSb4Sv6y6ISeYE7Muas+iisKxoja
atdyf6mdDyMV8z9CBkozNc4f/LRQFuEuD0eivw4r//u/fGH6fRdgboxU1udbYymt
g6c2KmyWuAEOItql/TX6r/ERfLhi6CPwv3gp+CoQFj1JVKKkQQA34cJiBfMrD1md
2TsYeBOsaLLd3/mRk4c/7DZMnSYf3ohHaUmDdN2Z050nOlh+ZTvkvfDyaEzr67gG
xx7vcoNPFwwedgJed0Wgw/JpxAhPC8S37MZ1hpv+gQW7IHC8hbNxoaoJCzppp8ml
dSkoqH9oHgO9clcmkhNCaBUuW6mp7npspmmVOVkDhKlGvrEx3Hm8SnjF7m0+Zfbq
ITexOgbj1Dcv+WxDxrS6ahjjwd8946fV9BjkERDi6b91C7Y2teE00xEH7+JxJiiy
cYno59BLvWQS1AOnG8UwGdj2YBHhM1Z3AaG/Kykgc6x6cwKXYFPkbNaf0Xn7UkHL
b0KEQhSKjz+UDc3tEZcgxgQKeeHldLUQLx//f61F+I/U3aEN94efYiPb8nIyyuZ5
jC6YIn5kqhXm3sM63JvJ7IUfztj++OaXiPhAMkMOJEEqSr8TtNQSRfz+os3cusCQ
ql1RKcTUZqX/OS/sYItbRZSzshAyu+1robZiD8r+pQbiz+ydgCxZLyAzbcgBn96P
0glZNcgKhKdVPGfr8AzalsHUveJgsRz0yygmiDNyZukJA3VJWziACpKeFEd5qpkK
wvW4r99Kd/7jQP/dY4mxc3bdfnu/MjBwnBKhBEpHWIsLgWX7M69UvbqaPeuY0yNc
7MNDJA4S7O6QURMrAQMF4uXomzM1RHgLmVXzeJ2FBwTAX8whz+ASKMsmu2XU4TD/
5TFccQqlSLe1PEeASkpynyslQmcO2id8svRx4HqxwXQCCOQDVwe+JeOeFuHFjPI/
Ov1p+DVD4iBXdGsl8CDljDPrEJo4hEJrrjEGeeVWu6lml3eREee27YpNb1+68yV6
1tNqOD/5rnx1VQHImCb8q/ajDxoNM8bBRoVn5lYBRMt22LP2XcrTLiYiyHwTZVkW
wRhaP6xEK050tBcQUeA5gEAousqbrij/E72GI6Dt6I4E2/p9dWWJn80lDRWeB6NG
dJQwUBsuAYkUAnS4cJ7LZeTcnkf4GlZjHgxqR7a1sLp8ZsDazN6OetjNT2b7UHzl
AkV1ZSqv4twyy45W+yIkt5nV/q/5hMQRxzEiTkCgTqDmHGff89ZxAIp4TlxSvsbX
BB3h+phqO5cipCqXdTiIzR+haWVCVg4rSeW+HeOCd0sFB+vpWTTfGxu9VVMnZ6eK
LfwMz3gghwURwM9DktqXZsMVEI137GTqDGSiwGUJBLmVCeSwZB2dApqWv5o0CeJV
T87zhY2NsBQ4HxHudZo1A9kSHIk6ERRE8j7N076vW/VCw4XIhTod7MI5FVgDD4pe
tLM2GlgUJc+Ey/l8K3OuVtDSJ24tGGDOpfx7c615S05OI+hOGQaF+ufhwy1izIlr
v33Vagge2Bi+Znta2bMhEG7srlfRta1KloFz35rbTq9I45sheXdbmtUeRbmetD4I
d/+0i0FJcYEDQR713q4ASULdriwywYk9SDf01Ujhuw/tbfO9A7o3RX8ivCGpeR5A
xpLwfZts+/zqQEJxLlM/hPCQ9YRruv4S9VAG7qdArzPxTzD0/clEUoJyRCVIQqux
aPoCunGDpCGs0aLKBAvsbR4KzJu/WPsGvAr0BURqURzNZEezkjdx9Rw0IF6gxSqy
D7ps1IouwqHFxvUnyczIVGcyxNAy5c6y9Qz0TIr5wBKhX4ZwxKjnTePryGZoIo0m
50vLOq6O0WopKMtyOU4HjesFIo/iZNcWuKfCmeZhQwDDLPznxbusCfCy0Sn0fudR
x8cnArFyPbRgeygZAlksckwR6kJu9ccBd+vsBfOhbsrqmeQqP8YotubUid31aNBR
5kyeBXJYNJCg32FNe7kCQu55JcKkpYfvKQTVuOezGOj7fNZ3hcVCOE8iuSE2RXTz
PKvBShBCjA5WH/D3dWQxD6TwWfPBMFRRf924Btyf1YaO2Z1i07dui7Pnt7Yfm9en
upUYeGw+qQ95rkG8ObPXzrYhzo4M6IG6TYyePzIRl4GAijQUHSCHjq8bJtHZlECQ
+zMxgRusc1WB+WIGspNTIh86/mKa4yxkeTahTiu1NLmQw02D/uZMdg7a8OnQP8jY
y4EU7kaYMIA7dPDXI0FubIY0y2oUWJxxVAQEp1c0AdJVkvzL+9f7cyGZFVWqpvWW
i3/ZvZJ3WQXGvahjPYJwn/skahFCBDzE0vrjSKVpV17T3aRn1NHA1hwIc0IBvw8u
Z/FgGeyM7VMePlyaSvw7eUOpfWFbBT4+pTO7WwnEe6mwyccXxW6x39xWrzVs0qSn
pS0HErr7n8iEeaeMFb+oWjXpl4XA1Tgi5VWyylt4k+EcHnAho8aWhG8cj1pUlfRB
z6x7C6JMiZxy/dWlVVYVYdq2NYmRmPOFnRcrzDq2gOPQHsMUaOTzdZ685AkC9Qz0
pLlY6NOl7NcyRn00wZPCXTJd46hIFzV6dYrYZy1FSoAzjP59GJf3fo/p7OJfN3kB
y6W1uQrSm21kXQ+V5Dk6HMHiW60p5RKfGnbJZZdMzvazLg55Yl8ltZ9gZdw8sgwo
gIb14a4cJjX+kBEJHoAPIgvgxMCePIo2JhDURemxluJM2jAojhVKqSQFOe0Q8E46
ddntBpnYY6JA1P01tvGcd0eXJQxttGAonDtx0Zm8ljC8vlf7SQtoJP9SNK5+/GE/
/OKsM44p4Obc934NWOYHVavuSGszXTHQpIGoeSs/ZE3nBUAHUBYDwFTK6Eg6IwM4
lriN4h1/n0aZ0kjPBBVDjreWNGIrhi+JcTt3bwcYcEPs5DynLwzieDiZxXBSmfTZ
wFctWwvRMQF66o89+Tf3RqQkKcLTQcKqntERf2wPxUZrrSo7dJe007JUrTx8d+Lt
5KzIWdzW+NJklAZGgm79f/UfHPDvubjKftbXnjLMlG0SANzZ75vj5LHvgAEHzo1g
m9HtShDeS/A7OtRpQqNMkzsGCGxSad0JYfw5mAhVAbGwrk4QUEdBvoZV1mi0sHHW
0LlczlC4KZcg0785kF7OvJa15o8QTWR8838AI3WhtTkNLyyTzVJy3TQ+zhVg3+T8
LAiX0UJaIpcClAI6SZXclTD6GjxlQEQZII3zbSj3rypNXYT+ifutJcY2KqgbGYA5
RUt5Nj3mEMlh5viK6Z095dj0f+2yUpaCEa3oe1PuED1wBumC4/3SIKHzLEpAzW3Y
ZDl1Z/3Su1bKAP3H1ocC0v3W1aK3+oJCUc3D/MGcq7jZ7u/h3wWmUXzZWxgYaak0
B+jQyA6BjL0PNg59k56hGV4CtF2i5Rs2AU55DGEaP4Cwpe1Hrmi2Xm9sZOLVeolq
mileOWJrlCwghw3RqrNPtrnh3O1GJoMn8X+Wf1+Db9mIapDjULkBKUOKdgkSbEeh
KhojkcvMWFiCwU/RGkWVtGnIMaZHhgx9oM8Qe6Ygvzjv3ITP5ND3zpvun0h0qb4o
bJfUNEcxHWFsWDPxqvxb3Fxri+k4Y+fF6yY0pJB+PE283V6EItVnoaflwjLUnLRp
x6ZYyMBYB2quGZw+vPrETGinU2MLbHOmu1MAzMr4ijG1/HxTBYDnuvgr7uu/7kCJ
I0lB9LGGGpwbT3/Jn6R57lrTu8sotoYnsrunZMgqnwAgSWUUhweW8GGDgdms4Wfm
Pzl/RRybbuAyzMaoueP1ya46lOuC4NYwB5mDARicsk+ujLweZAJ7aB1oOUcdI0wP
1LLqNDXlrq1x9OclF4L90w679tvdiaGyGhCK+4r6Ctqt/GjBzysYxwCkzr9Rpvjy
j7P2arUXoXRJXtAxmBFaSXH6weIjHs2BhDp981OsDeZDjCh4DxXKUDpDu7DR3Rh8
QyD1e6FqDkAyfq0zzv2QlTR7y5yCYYMrTgynrqaqxuMlemq/H3pY83B7pnHgXrKs
durSPxWzYmFSFONTfot4l9MIxbumNdAqr1gEJUqf4L5Fmm3N/CE7/gwdKhNyaeL1
+g8xLbUjN5SReKrcpFuKQiYU8AJ7yRmI31q8xScjZl5ITE0XK5rmDDItrxyXrQR1
TGUI0QYICdaqZFgi99F2NVS3Y6wpOE75MZd+Xo+aulXyaZbRj8Fe65D+tyRbRt8q
huGHZ/HDU5+7I7Ie/DnQg2KuKdzSIRKBzZh1WtOBQUuQc25yBuNmOu9wXUe9m16J
kwHLLDSDFyUqUjwXsvVr6AQHLOCJzpH8qS3wxM7OlIGdLgUEdl8KoZXro8XPWXhO
mmjoU2L7WszvZa1A6YXZrxIEJw7t6mqto6psx9c9nH/uKyI6MATPumQG4KSfCGMp
rJerxnmwpNMGKjtFpm8QZQpnlJAAJ/1RWS5Q70Mm33OC92VfYCT1c24Gl+zIpaAq
G0G5ZtkFNmPfIAKZD0pedGKu8zJwXjQGEFX505SejHKiaNJmPJZaob518cQWsaYW
mwr7nK+yJp5qdVlb9AyTo/XXNahzNoYnDqoosTAoyeyfFOAQuV/CSOouc6RZlWdr
7L1dGwmAGzE3Oty1PBMhgQ4ot1oGqREekYlSyWnIQifN4yWzW5xi/IswQo7OiC7c
vfTnZh6wjiaXEdeFADVuRhF5lZHTKuG0d5u4oWvrJksLOTlvBPsSUbN5XV0mZhQi
tRo6SvYPN/j44Ui9LpeCNdZIHJbVlfy3/Pson+LZzjj6FLib29APSDdk70vvcikl
mfIjbXKG3FfqPZkOwywv9DCsrArRZtDGq+p2Gwj8f8AXkpYPjP9UmQu+A9NChlzz
YG+4Zlx9hDXAhfgRVJzNV56E3X4xgpIeR9AceNowb4sqIY+YGraqVmMqdGW0fQUV
5j7jIOpTk/fKwjK2zeaEMLnP8PUoWfnmxXdEW7+BTP1NvKGbYBUWDJ8JWuMGrTBW
tMJ5o5IuYQufPqIisDEcBHfjqaa5X3DLtZuclTJs/31daQ0vrdPAq0sSToQiEso0
EwSSLFmPkGgYPEM2AeeBlUKAkyADG7pNVyLCcvZ9ylvtW8hrASk238h5brGLet1f
g/O6ZaMfmULF8AXtNSE5ZO2rBoEOBORgDIJimWTfdJpv+Aka/4Xx5qBqIQAYqWsi
EpUaiLcesY4AMGDiijpaIVtYCTR2p6mWeZXU5vnd7TBAgRFC5+OsWZXFDDqOTZGp
eV5n1Gs2JOc2PmIdyNv9JQuOpWNPbkR+vXxqtiCYFWAKFqSuX1YyBnpgV2PZDOND
EHlLI5uUwY6FzRee78e5wWV2RBeGhrUY9zq9LgYZLT/lMbSGf1+i/n5bjl33Bj0f
O8dpWffC6O7PRXlki0eDrrGQvglkjlNlWzcdpT8w9jO7QUXIB0Dda1X+x42rl5MQ
2V+Wzma1yasz38HbIuLcUGh2T1wdUej3LWHmSnkh9vvkmSeGdtbZcgsPVkQ7TSfH
+vDJEMhe2MHAhnpdIaDm9f3/WVSGGt0VcLnmz3ewQ0vi6v4nUUSaNxNjAb/VmpBg
ijMRqHTijwEwP/z/uIwPs9WNu62j62KL1kV17M6J0A2h0xiiNd07/8ZFwzuuqpvm
tK8uTyuTMPe/JSEe7X/MQGJYXwZZAsRYc+AlE+yNGk6TvjN9Qk7JnwxUAfEE2+LS
PacT6JgTdia3k8wmgp6sa60SU/q5+N4+BJmhLtlmz5jIt7BV8pwxAqCl/T0uhJLw
9triY0cijjGNqZTOHDueL1K5iqwVD9pZVASDJfggvTo9XwsGxblblQwgVpslroBM
s6K8X+iDtl8pXh9uciyEr6iYIfzDS1uRR5sI/3JYm6BkjSaoyLwp9JPzuH8i+lDn
0rCM4GAS3e3hQPVtBf2nIT6+YNtiZk81XcoU/ErV+MPFXu90rhqOiFl+epAN56Tk
SU1NUykBtHojq/IWNXQWzRbT6T7rHnaJRSheY3IKty9ZlPHxzriFSx3RTTa59jYK
YcemM27D8vCIzOOmv4lXNyQ7cOCoPXlK3udaMJRNmQVGJ0VqkxUWXMUfT7eMcoBT
19c7G9pOp4q/p8HJabo7rj1FB6dtRpGAFPE4W5aIkH5DJUCT7ixctu/EA+0t9yvS
B/aUYIIQdwvIGvjieRq2NyImcknhKHBosNtvFE17sMjxOkPF7+bhcDkK9lEl/Zo2
yTSvkeJGAn0Bt6Th3ixDJdkPgojNAjzBmHbgUaAVye7enHg6MzQI/Lvx6CLA+mED
OOGMhAyHYv0uyDQBoI97m2nva52z1hscsVGvDX9lA5jBDFebK4+dvUnBBHJ/5GRs
178pKhXB5aVgBPKYnHEpcr5MlI3i97fxXOxIVJcDiEd1OoF9aLwZ8lXfUVbbnTaC
CRTDxbGeTvvGPdbude8XC6jHYxyPCe1UZ1LJSXPYmbvwwrn65zSoim6HHzTPiKY7
yIubFRg0U4FH1aB1zh9PxJGvf+S+HgKWtdF+7+ldpmtzjBI+OR8GrEvnF31arSOt
y0fhhPAGqoCnx6NEn+cQTVcBo2SU0ATICdV0tXoDvAW4SAy0160CDLGhNRrnHiOO
nOLxH5MguAKPrB6OqfOUWTQDiPJAjxBu5sDEjEH3XQQZZisly9/2UtlRjYk2wyOh
xQtqABPMjzS0zg9ndqryiDsD2yaitSKj4aqNnMtqlUZPgHcAEsO+CpbclWirmCu3
LXcyb/RS1hd7lWWxuNiVIsKjiioXYWxQpLmEIeN7KFQ9p4MbhVZTlkAsnfE/c+Lu
wVp2m2oMofo6hFetLN5al18S/NZp5Uo9AJFv6ajtEs5PpKxEo5Gc6cgceRCFfz8U
flJLouKEHCci9uy1vnWVt0pkHsVBUgdSkBMHwaAvhsjnueWfaoBlrfx8WoEbAwry
5d3+3R0ne82jDB6r5yGU/7Lb7ileYVo2HT9U7HceYY9tIvpRwjWsz47/qeJICuBe
zGC5uyMvMyNlpculEfFf0GaNcBkXVKdyFaAwwYAJnV7nAi0u5AdmdohvPyE3T5Of
YbTkUIAYlypQYq96+BgWeI1dd1Bpvgn11R0ZggDE3KYqzTYVhUf8t583u3/lCe3k
pa3t2kgcyIm6ZFKi3iDmRUfStVOTMxHU0h+676mz5MFv4iTUxEsXcuV3YUjlkrHC
4CSixJ0J5/xjh8vVIc+Ct6hu34DaLf0ZV/vrdKYyr1teFFXOfmDnuNHT8HOXyTev
yPdJQuSS/4KXezqqga9ZesEsZVDpdirzhO1LL4cyBjn3qkvTvnyOBe/uj4+78oHD
iEDtOLEugDFqL9HU2N6XS8drkzjFAbjTvheX6/+abvZ8rPLtMWc9bjW1nUfYvph5
17or/AwrmWO1pSy/1WkvUdEJJvlvu18SdHSBSl1KHWH7tREGZbVtVgl9N9ftWMQt
85acoF7GqSw8GwyFuC85hg3eT6E7IQL+htyb5KgDKXzhAKTzJxqAiyg3UDv97Crw
2v1k0kQpEsYFfCXQO+Oyq8tT1KcitEn4oDFO2R3mfVBkZHYqesViBueCUXoX+Pus
eG68pyZNUtrC9Owe529ozpMi9VPy+iUKLdwh8ZOqKd3N6lOCn3A5l6yKXDA2VVOV
4n3cYAui1hqUmzTiDo3n1cT09TDMVvWJ6dCUQsutaPhMES5+fACjco0rUfmX5fHz
ngxKbq258cy0Bbs21QwpXkejNgfHWBgq5RiBCv0hPeBYUaLVdsf/+jchuAPztWu1
5oWL2jmsR0whWxYW57PKBUJ7idVoG7wE9Jt/+XR31Di4VIj1td8WNz7fTN3IEA7K
YMW79275ANU2jiPgr0MyQGzTnm65Z4irq5nl1IcPWRiSQOmU8o0dS2B6u5vSbFBT
pqbB/rOI7wMs+jOW5FpnKpsP3NgR1xBAprdoBaQ+CqpYr408bmBY/3ZcdtD91yF5
WzeLr2sR7emXKhsX/1bcFvRJMCMsPxZMm8LRH5LVFybGmfvhU5rPZdddIlWknjm7
g/OVauvPaTZaxuUF7fefa6AsLHGvaLYsvmOKlJKjLfx+s7Xf3VbrlR76FsEBeTPU
4dq9M+ZL2Jv07qK4UQtgIxgi8nNC+ir2oEWzss5LCbD/Gbf2mrczjU7MaiZrjs6i
XyK65aN9vXC5EaiVgk2SQHGbPB0I5j3fg4HYY5MgBw5evtmGuuyjTOVPnd5GfgLa
MXD2uo/CjAzPzH4/NfcOwz9pJ3bLt6CP84eGboqbArNj55QIDRa2EVVx4wr4hkSI
HGAhII69CRSmO/giHJjxOWXRU2a++8xrlFOZ9PJx0vK7p+XMlBRA8vVZKOXgrLvj
MyWrYxhsZJXv3PDI6Aqz0kv50Hl9MsxbtviVug3U1vpMi5Sfyp/KiH+lsMxp6sMC
7GmWMULY9X7hghS6Po5Xq3k1dzBKyW00bjodQPjrl2PPJUSBBMkzZDz4rEKHOMIv
95WPpBSAOEmERENTH0Acr6EYBy86INQ6MBIDPwFw7gQVYf9av05ZS6wBnCKfp+dT
XM9PucSR9baPAZ6R+SuCL1BqwCzCJ1/STrnIAQ+z5xewo3bb83kLzQxRDFa9KIn4
W8A17egSDPrsUc0QeR7wF91rpq4IsVyMVlY4z2HPKD0bBMs6WiaOX10AcB99tGDl
I61DNfGXxzZZpMJYF5i+hdxArivDKXyCReOyhNbwCHeMqQD/z/V5KdPJrSVQpxqi
vgy7t8b/odACf2Cg3c9IFPnNZ0eqDbFQyXlQBT3J/wXTHN72Os+XsrJ0SIy7Vc+B
mCXbnNSCCWQDSGxJYozMHJ4NbcW+52m32jmVtaMCarVHCnNCKMWvh7p8Ao9ZaEI6
q05qig4mA9s2VpROCXVZ7l26k+QqMhvt+kMfVCRiVe64QR7wztThZkRrND9GKlG8
/MdWx/JJoxKR4WqmoPlDuPq0gl7bthDNlHAJKfvGTfov/qvfvtBGXkVURXk/aSKD
M0pL77RG9FoO2OxBZjEe8K595PTevmnUdCxvwm8nwETtIgtp4kgBXPeaOOoLAx4R
eXa8wrBujU2EoQvSZlD13u+/HinJ0Z/sQhIhOt/gqewkDAbK0XdNRi0OvvEopdw6
kL/Pdlc5qzSZbbqhfEX1KJcq9QB3sln2geCg+Z0NkiG8Fk8xvoDKrxQ8mma/yC78
UIo2agkoIQHpStLycFv+kKrcCt5NjxL2OILBDaxLaJ623P/jmb9WgDdm5C6gn4x6
lokYydwT7sv/wywMrhX021kIIVcHmbotuMI/cOwBXen74huYnM99qQcGu+EgU61d
EhS8P/wIvgz4I10OUj5yM3nvJiY+nUT3Mre4rSz4fEaBaKBQ5+z0kebqeVYu5v8T
P2Um4CDj6BRACksjJUo4OFNQSdf4oCVbJ+HuL0SIXZZdLjesFPTL8U2iPwEdcVqK
KBDSQAoXDP5D48hgn4cdf8DacfexN8bHX/MFunhbGGYtMJHioDe4GLQop85Mg9Li
/mrURQroLkGDuIWB6THyCAUtlzShKLYrk6Q9pQ0utRDAsrROcWWlOKDzReSGM5WU
zzLCTE0AAe01XrTDrMby4dbvfweR6IS+O99q0wXk9npe45zTjg6HMSBTIwEVSmhX
IjL9yu0GxcssjZvPYqI0SXGYbs0N+Nqw7mXBZtvYW8Gh5Xd5NQstFHjzjhznWbrj
mVo3xppElhQYn9yEel2ui6N+V16G/cPLQ1vPpazmy3uCxW5u1kDjjA2Ol9Z400gd
UD8dkkd8c3Yj5E8nVdbgQ/xCsnEyzcWSWVx+Zfxw3jZVSj7GJCcDV/NFqFtBofVs
qi7oxzwv5JjZq4bU+djMsZwxHjsA7mZHa5JKfPKcj46/tyJDdf/fGyObOG5Nx1eN
g4zoOtLAyrRkRo8R81E1zLCKK1zi8bo2KhZdK8EnX1zarZU1MB2RHR++mphA9cr4
FNymfh0QgVT3oDve2N2h56+1eAaCb5lltHPmnQ2gemqx8xqTtooy70Uj6oRWLQoI
6Mrsug1loOJZAvwzsN6VOR4VmXTHxYqxWJV0mWs2vjVu0w43HqMAU0aQ0iCV6JW4
NH5e0rqDRfFEsCXOw6hy+QF08HuyG5EsEXTv5hjMYXoWmaJIIjhQlLaRKTMdRO6a
eWnfdoPMKDLId5MvefEYJUSBbqmZ/sOtHfuqi+iAKk+RJnq0vvwjs/ySDWYuG1aN
EPrwCG2yJl0mvJlKF4PgTDUOZHTwDhe3UvjVTX4ohmz5gWA+g6N34ii+JuR5I5xl
iRYstAMlALRb9hc5shPt2E3A4lw6Af+jdl6OWob4iyi9VRW5IWJPKlI6dPEhbWo5
CtUCYY1iKX6DDN5dlABltWYOCA0GMzwGSv8fwtGDKESMoQU29eezWcbXskqQD/aK
PcRU1VaMy5moNN6Lo3g5qPIy0Rq0fY/xCItXPT4jI99OkK9jvyrooUFLJ8nbqGeb
g4INDtjWauTXrdFVVH2oRtJ1CwbuuSUzZlb2RvHx+Aix2lNr77YTUlS6Fzb00Zw9
rcqf980+UcBe8i5hEBQpz0yZthwmRPxhLFZchdGwXhL7wjq3m4+H/Ntg9RbiAH9X
nOOCkZX2PA0Xs/FF0sNEhHkWIjZP/PO+KsVV5wJxlBPz3YrSGpU3LiS10P8N9Vz0
wATvZ7fSITGgbqpzFBDg4dt50opLru6aeuGXJ+8HWULpILpEbLPyIXqdUAaMdWk+
VmELkVRF3vUVA3sFS8xDf++5rmn7ycZ1B9iG/TGoGGINO+kk1NiwJdHJHAZetiDC
iSyKJ5Ettt3ViNOlnPfSYIG35zuK4ob6AVuTjXE85/c47OkGtSRABOKkWHe2lC/G
QvY+VRFKM5b9TOOlX/ZzAzRSJqaDG+2e5nJu+WusSmKNykqSPPGtmP5VmwHOgIoA
B9w/pI14V57QCIxqB5Yq2Q0bMATFtPRw+Pu527iegIoZyb4ZQoF+fLITs50aKHv3
gFEvA4s9op60EYFSKLjqaV8PFavNPwRv/ynD2c6+DbmEK7KxC7H1TB7wuaoy/gUP
z6xr80hyBJI7L5Yy3qejfPN0KxYJLJ46pM/y7WJhRo8NJYJ24EGo90g2np3CiE06
HwZaDIyTgW/iVRANpO3XXxotogieUjLeF84qI1CHc2Mr7zyNSGXkut8HYNK1a905
ZOQW1pzRjoT06cIgaoqxki0Gmm7XE0RYlEBcz6W9FyZMCbV5hppekGf5b4PA0adG
lEzUYAgcK4HsLgtS9ne/M3NvnvvXDoi1f4Mf39lj3irVLO7PLIkDCdk9UMW+QXGW
lJvnVX4c9fz6oXTEXfHWAvo+Z3frrZC0Ap+aJQxAzrWMQOPZ9JmfZ1Z9fn6bdNL8
0esc056pY1ZGTA0xLnzmYSFaEAAY5uIxcO+/m5y4C/pB0vbIee9cbDDYsRwIvHEc
Oym68tn7iOKvT09wV62rF+65HlnqP2pvPasq07GTuVTEKb/CKoaO/CDSuyxcgrgL
LqzZPX0pEHMYSaJcErt78E4nho0BvS5t5csfhqRou45ClpXEys+Aa1dlqN74SPi4
zNNa9QX6QlGHjJ7qSCSAZcG/iSVlxi1WXHnt09X1AYYRVFqREEb8ok592tOJsuZY
j7UmmRswCwZ2aVB8j5uOqB6a08zOxFRtUNx0fJcp7gGytTxkxEtXNSVU3NF79ZBQ
3WhOOUmCFyDU/HCWOaYeerqAm2PcFvp+yKiJj7hJSqsF+gcXk0xgVo8ioArt58dU
VhX7zCqJCbjC8PRpF2grQZiICN+jw3PPIGKulz46zQMXFKRIfVqRkuPdIc9ZRUoL
CWGAfDAwg0j4LQMBrXXFhRjbKCt5GUotmbmSIQFZGUviQ+XKEQ+1TsSB6n7+59Zq
3BeHPttAJMWQ2qVBcp2BxmWCp/i7m5lYcqFmE6BIGVi7Xvq8+HA5CXUuD9txNtXN
h5iUJ2rrTSUyw3zLhull0I2gPwf7mL90B7KaGxcPWAkLAl+vis5SrBbxGOeVWxd5
p9bZmkGPXAB4Q2ev7k3dGgv5Gxb1dJSzQeURkYavqXOmodZfvWLXlZxFop7uJOiS
IlxxNswqH022W1hW5Bek4ev+6aTugRR65QqBMnYGnkbHNauBvt6zMMvrfQUXLoYX
ksKw09Yyaz5LkaVASBp3QQLB9ARntZqM6YBdrsIohk0bNtG7+bvKHXNGDdypRDur
Zqox1UMGK0zzKmTtTBoPBhpv06PmRHUgM/0dT9AdSo+4qb5J1oM185SuVlGHnGYY
JNIWeLK0tWfmiuIXBa0P3AKRCnTjT13M1t0/Vb/jyTapsPqZ+06sfWYJZMHP6LBI
tsfFO95bRM2d3YD34025vsjCJMfrS2nYQuuPIBoviro4MUo+jPPov59qGFLjQtO1
almUMx8c0FyMZFocJSiCZAnCHJWPFVX3G+66nqOwQ1Hpcm3S642MmuG++v/1FpQm
0zGr3VRt5i3k36/7Vjp1A8kOOjl+meIeVn1pUo6fT6u4QBk+IOZ4+1j2f0JPxolH
FYpAkMtmI6FkTeGrNFW5EElJKaoIrL1Qxj0POmiDJbvGNcTqjkzieVJgtgxpYJ24
3GjKrRFdpgdwmQhQKPrWm6qgSb7OBEroHqsmI0YNus21wEjnlvAK99D4dzYdfe8+
owG3FKiqAUK8zGOnSOhAY5ruOa6tykMeolyBp2OH5U4tiIbF54Ao1HAhTmHTqo8c
p9S5RA41GvT/rwldu71CMm9EHol8hAZvSyjO+8Wp07n6Xms2FIqylj7MgTY8wUj8
l8uoZ/bOtIumBaLDFD5gjem3nLQYNNDCDi3cn2s3FQuII4cYtxwsK8u+Bz02Xhd1
wQ+zY4LgjaNeCadahkJCv7QZDdocgyyA0fbbfkilWZCe0j5FrONwfGrJh8xW2FGD
GJHCvhdpnU25np6xtfWZ4dc3YWwAyBNS2G1K65i8SZUCXcEOsh5egEUJJUBvNdVj
pBQbUjkTPjwNd1JZw7YdzldzZHwcZudETndnCOf7LDqJCeujHIvFxIbbJbbV3iRQ
Cf3yR8fg68LXv5SxKZ0oKOCacAa4o5yGZHPFbQrG8knJHDRbIpmU0NmkeZc06MHA
HYSvRLnOlHHnDND4PrEZ6ar1IirZ99OaGfBkkAm0vWTp47KJSBCESABknuME78Mi
nFjKX3naMfWA4uAERrox2bk/jXCE+DwZ2aTnfvNMG2FfqJ0tf0/Pio9bAVNnYiBB
D4BF2tJUyK9Q6QyhCVF6NAUo69xFWQGU9b7xXqs7pOup8I1dzKrWrHFss2dwoJJT
KBatN12dIsc4N333oKhl2f4mT6by/2nRY3N0aGLkDw2GyC4cUv4yFgRcl0jVVnjy
j3+2NPEHLsZGdcpFLLV92nOZeDCEQTpuV3jloQ55r40GFys3uxyW3B1AlBPLCngW
NEhEeAHNOvSgHDu41Gg4L3URb0UtzZw/B+DA/oAk8yLBZEdx45DquoOjNTXzhxJs
n7KOhaPkyg7WM62zpzzYiokXX27Qt3IL12R2OMWCpp37RSfy0a2gG+YRGyxvahB4
saGwZtlZj8roDkd7H8oIFPooWwHkjOlY/Hi5jp35UzgqWuAHyLdBFwyE3TQH8AmS
AfAw5cN6MbIxHInPAULE2KXTNBjnNG4mtH+XOo9vOnW6rLDAnUatnWJZbiwc6yGB
KqVdeoztzcQl/Mx/qh2S0TqoIMzehbOllsxPrvc4njBYrFkeyj45CpK4hMA9aRH5
MZSi4WyPkDjbj0XxKyK/wcwk8wHrHjtcAp2wuLzGs5HkzCj/bZ7OJCnT5FImz6w2
9JkZiAPCWL8mh1CYwpwzESDJ5KanQe8hEJPs3JGriwMTYlLfwTUAT/XgGLMDsPTE
4ju13G0e8G2IxhDeW+bmYUKvXZNaSQeAS/VRPXIOgkyeQNpQsHUhHIqDKwan1Xts
aO+wS/Misg//ynC4wnZw4g16ucuNvGx+9MHUkgCYRT4MnvdP5qqTFGQrUBD/czAW
vsbunbVl4u5Oy/MP62zL3dPSxG10YBnjwM0wF5PWi6EF4xTPZSom0BHCwfGT8oYT
wfLwOn7y+1t6GV7vuoXB2J0PyOVRMo0NgAlzuxIDTSfikggfHYoK+q06erxcb1UA
Xlkc+giDSCOt2XKjufAgkEOQWDVwKFlAACBI7ihah0WLW3xp6bQGhSwNbP4ylIPA
rgbEM1zN0M4rPxCLkFdAMT672OXOFr7iakFb8TGofiINs4egclJ1qy4w2uMFLQeF
1s3hHNeve9DGywq5kR7ya44DGHTuglh7JgU054W+hvspEYUlpqmYSA861xWN53uK
C1ak6Ef8YMsU3FrxEZfq6cV9DPI0GfXFw2H4MpzRqpQ/JYKdGMooNiqWr4d0t0Kk
TWSVpjquRn9E1K0jK2Ml3dl8SYqUNAahNUPbZBNgE3qMDDCHjHSu02gP0Ku4bNEK
bPFEmNT4u1gCbOnN41IdTJudgkbPUgd6N4XRBZpBPQEzIruqLrAxLiSwXClsdYkq
1X4jVXbEoTlWX9mrzNY73ZO+prt9GsG6Bt+tvE743thWeY7sjY0d5De2PONx/N2d
/7C2Xr8DoJiZmECktKIujddy1mtVBKjLYgNhdOxYfh3OmN7uGwXsqdH2HI4zNndZ
Ieboj27GdXwgRbOgzDCBX4UE5YCMQ12FoeJtga4yBDHKKlmEUqJ2jcBoGnXf6/cN
J3UNzlN+uH0JNj7GRxqKeYmun5l2grlRjfR3UbCHtr8G/KvR0G3gucy+h6AOszLF
SG9j5IOWh326qY/akQsiiJ8On1VVFRmk+qiH18xi4R1fo1VS1R/D3iyoli+CwRrR
4tLeo9gVFhzERz8+N/x75THaiT+/lGB3RjQ1Uhx6jOueX7F0G5YkvMoq9uGN0ZlO
lIFOzWjAF+8KQO7SbpMxnKgEtic5rINp3i4i6Byz6urqUj+d3O+dhSTTImUep/3Q
SppYQnSjgmUtW0dqrlxWIInusENOMGkEgG8gbXlTQVCKYBtujPNbBK4cvBKJK3vo
ZqG52XJYsa54Tp31AAdrkQy60VyUT3WiBe0vqQATAujtvX0F0B2Bvw/W5EKjM5Oz
MoeL9TN/y/GbIizHxOz0IKwoLxpWticDDJ+bg8YFoV9vPAA+ZkRk6sEktKDKpC8Y
NAKb16bNFQSx4E8m1kDYipJ+Ps6LxJshpd3WVEJUqlovCaKafql5/Z6mfPQI82ap
gqH3QIk2QJYQL/h4kHMlXFJ1N6pEIrxvj2BWfL5pkX6s5kqGJnCbOELW5HcVKV0b
lN+SkMSXz9q91j7tb3bi069DOX4U3O6VxOb77qFCwitCzvRwFoqLU4nkXy1ocsaG
NlM4dpUg0TIsmwdRjhf1hTeU8mfiTFb+ClReXWwkQQooXFMYUc9HkQyJJA4Oo9hC
cUi3fGP2KCuC+x1QQLj6ygIDKwH5nD+tpc0f8muHRhjVnP/zinv13czWKsKwS/C1
KPksny1YkUzJf9cq/gXajlXZjDGLm6wMFVnnp4o4U3FWpsawOpA1OeZ6ZN3P6cVv
/GMCjmGigVRsvTycnZsIqqk0uckccUiphQ1xb88PdBCOAdK3BUqnZwPj9uJcDgPV
6ikhvIV785HrYb8koiZBnaiSDU3xta0tXqHvBW/6TmnToRwzhPHco4UMHv6iIiIX
+k4odbmZ/wB9aMmcPUGcCw5gMrV6bhJSZ5PnmNut5l9Iy16ZcNrj5eda4wwkiJQ3
aJ8i25YGa0tpsGJTfFEBYqWYlnZth0ehmAH0DMNzq/BBivR83kbC2Q9AKYEnFCqr
cuuzXOufve/htQfQ7K5Z4C+lv3X/aIcgCaBq2MnY4c55n3fmYBH1EGWLjQLsUDLS
5P4k0oyGq3EXJIiORiyYhC6mO/VPi0TC5OHKMu1cZG0YQZ2wVlMiBvgYfIuEQ4tl
JkUjhM2GZ6tUJrPBn1QZQVLIeWxjnb5sHouD5HDoumuVzSzBGX98Qvn0cTLFNKE5
H8eKFfBejwWt++OueXcCgC61uo4H0p8jCemOlUZA1/xOe5rj7my338Bio57pI3Vi
yO/10BLbT31Nf8WD+cJj2/lnamz/nhEDFirYa7zwfuRRx9jE47b1UQ1Oy7HQzVs1
JUy7sd24DowuuWnK57QAO9FPt0gnLsQHbPxa2lJsK2aeFfN9iUlMI0Tce5Dv85o7
lWet0zZzAZSszuMmKeOoWsaW6KBa5wIGDZI1nx+YO6OLIzxVoVWpTYOq+DYS0QYn
0Yyf9uMwigtdeDBZKwdy06Q9vYfXXaR72Hsc517ENMAbZgOxjLj0BGwNaHRX6KyC
DfE7vN/CbnCBNDu1+bJDbOESZqhSPzr2tyXyifpfTMUKbpQpXQNINvTTrcHdTbmV
I2oUARztrDDqWywsuolzJoOKiCPjjbhtT05svhY1joV1XjDqPALlwmTd0vnEY3SO
sm1SbzIuoRu3k6LzhZWdUbg3jyXMynIKegDpNocS1g9xXHLOa7lzxOdFLY5CeDTa
OTSjbRYf8bOxTRSRq7/rFy17GF0mKWvUPTTkHa58XYoP/MMMtk38jNG+popC8FPf
lL3Qy3/OWvxIoO4yRo7lAv9iYPp3DdRsdqHzh8T3DV41JSr0edQvgf0dJ8nIc+/k
a3dL7/UsEOGNCSKNVmWtiTeA1m1j38nqtKYqIEyPb6Kz78Po0raC1/RU9VyGWniD
v9+GTE854aHYATnZnleMjZlSR3vOXu8pVhaqBzF6xCG/g0iPk3gsjLU3vDwf7wBY
be4GnUnGfnb/wXAVSHrLjsesf4tHiw9duAK5D4ctsPqxXm1Vwt+i3jTTJxFUxASL
HJV2Bykzn2d6xFUK59H32sN7LA6zbbJAfIU5EJ+WXUaz+TQ1geoWyUpauSiuhp60
oHxxXfqhNRuvqdmb9xpXu0NRMlCnjSrLagsHvj7eTGRi7JKYLtdSMrFekjzIiZ4B
oEJDzA2n5Ab8FeMURnWYaOWavh7p1RuPY69K54czZMC4VVnECS4PwzYweC5rjvB+
05WgG90rBqsKwfvJs+QJdND0bINVta0lSp65cj0BAS0T1svTtyqUaxefnUyOjsm6
6ut/Co791Xca/oLg4MqkkvhRF4NPC5flBNreVuDiSKw61UcS+EHkzKcrpvYGgKTh
DL7ujDi1Xe41S7vQFy+2jCFLTV2+aI4Q2TnM4/qjxhxz78I4rP52sSK7oizpyzxx
fxr74lMdF1pv0sLcgaVSUraB1BP9aoDiV8vRUKE8l4LJzUMzjuCrF5MfPbZ8Eq2v
6wytkIaQE1Yuv0CAXHG9IpCE/gD7fG74O7+i4Jq/gs+smmJmuP2lgBmcbzETBs+R
2NES5Y8G4GhUBUo8Q9CBxGoy6YNv9vuQbXASxjvVHeTs+od1C/Y4wku+2lzexBZY
e9jwxp/gh1jOSOtK8egOh5CHe6yCLfQXs9x6zBwoONVa7DI5clSK/Fmy/cQQ0lap
31OCtwAjOkL5H6X1VLPv/EM1CMkQZb50DNE8p1eg11cY4oyVj1x9rPDpK+fIPBHr
LLS+GKICCBEN4lQFuJN8wQ103t1gMxwPTC7QwgnJqyBLrZJM/buW3iSc1bf7Au4d
Lv0D4uYX4iixjAFbKIQRHrTm0dJNnN35sMkIXn+pAINBCKdqYIBEKYUpKJ8N5oxp
9Kdoqtw2NCtsI+y6GeRNyf84mGJ2EsLLXWl7fgH2UBpXnk835SUU6cGN5liuk/A/
AeDm+wRX8QDTRGH1G25jLI6b/RQPSAFinRoSyADeL+f2npbOHBMwQSaX5zn1Sinf
oo6tLrTuXrq1TVMb6WaAhgNGlLbdmMZTt4dXs1nAUVZmU4FeQjP/1qI+mKDWWt0K
XXEgVA5iw32lbSacqPq5HfHUizMsKYcoEq/M/3eL9WfALh5QMDBEFGlBeWh88Yes
xOeOksSvZl/zeNvx1oa29BbaVHCUi6s8hzJFF1VGhusCkJO8BbsVBK5q4lOFSg24
ISMZj7qfvZbPfoW1EVVo68Y2t1V21G7rQhQcEuIQWbyRokiTe8lAhxuJ1Nmg1hKB
30jKAPv6M/d54LpqfKSPWi2FJFdMCf0XVYjYS3NthUkK2u+Cjj5EZsgJpHDqM6Lc
RMeqmgc0+S/qd0MN3bzksL2REI8uXqFPqeXAXN+oBHrQk9gI/lKjrDEXhRn5TYhM
52I8gdarPkNjkZYWya6dGTpeIzY1L1miPAJVGFPaxN/lquOYl3BaFQchu/uSRQ3F
1ZD0yfkMlkwhPoJPGSq8gTwL6PYTNfgTAoR/JtWawgacGw3AnM7z5AahEGdFlrTd
/RKnm2lmiR6JqEpw6Otk7VdK8xG0S0Ip2KP0dv5kW8/wH9DSRhUZazt6UpgP1zPm
UC5zOlEcKwRGn9h1QtnnAjW+LkTB+hnaMH8vuL9tiE+sFQaoUHEcRwOW8qNzjSfa
UtTNWPcG04OlsM2q8zkOg5uvaJ0qYD5MdN+F90fGh/Zqxmyop83WfHkpzDg5bTI2
/RoTX2QSiWjLbg11r8eXR1eLk51UNlDCivciMhpDYHIBh3I+Jj4BRoRzSnc3fEKu
WwX51rlEaojKp1ariyyaFJysv22vSLcULbtpGy4b0I7nbC5DcATnVRUFoCK48TFb
+hbhNC/HIT+DNkqJ7rHsBvnMWw8rlPcbZaLTOjWWjWqkITZCc83nnaa4IHuH0sR1
0nDmH4ATDmnFQEw7GNVRMS7N9ZpnHFm4+Ll6ISCyVjCkCGnOotCFDUIYfPqGMtTp
J8eTJORYlFlhPrgx+HkAWp0wDEbJxB0waVYRrAlhfc9leBKWyvIaXCDX/kcAyLkn
HTxaa6hMQ7jlChuIwL2aFFSCR/B+t3iyReuRfPl//rDz0ufV3O5wftFRYkLdtZc0
4XmiEOHOW/voJXhsWzByXIPmr/eGRobh9oPJVp7Xpw7wA6SltIanrk3mc7Xk2j6Y
lu+O9Xmv5nW7MfCJoKDjqUQwkEB3cUp4qA6anr42fcTVKC4YHKO+2OJXvw6yoCgc
gVtq62ovvhL4zqggqv+9Wsg+q1UWFuTfdr8dogd4LBCPPED/8l2U1LMYYQR/BqT3
BW/q5etH5wBHV5lnnsZASzdZBjbg+F6qLoKSp62TV6WDFCpZyFv/HqXXtaCx2ZUS
KlUeSvv+Gh2jqb2oaik+OhqhwoNQgNaHpDVgz4gip5sREza6rm3sgNHw1iLdX0cS
LB8BUOvVJDhD8xms2d1byIekfp4W4Kc0Kb8c7uthdOEkw+ssy1M6zaD8seLL2Q9e
RN+t15JL/cscP9+oktkQX+d8XmMSEId1g7B2pIYoA0x6STMm3L6IAyD1d2twLKhn
R1k+wXKhlfnlRlkHvdWVBGrrMyMPoZFy7Aw0zOV71GjTaCmMS6M8bedK6qLcQGPT
TbUc0PIVtEvtuFy4Zezq/M+m2rjDef/4tSJ5fdM09FYo19QCxKgCps5NWeu7VhMV
xmgjLeDC9Fh0bQ5iDHIlXuSP9ny3NH1cTUwZYudcCpXJbYKLtthBsPlNAlxL2fHj
YB8+oOCJTdVRvB1btT8QS/Plt8V7hCCmx/wzR0hnKzuRLzkz+sDr0MNX+TX10JSO
Xbdimt8y4EbsbL3Beh7EBsNcggaTfQoIHjflkirV56PNLx7nTdnwNsc7kyDrVPVh
1l03nUNPCYyokGBr26E8ncliOfidwWsCBbFcrujkJ3h1hZeypVddnAHdMjjA1tTU
mAvJPIbwN03wxwmtr6/hG4S2tDnwDYCaxm+Hiq0TYL72iQyM9lvJfkCiQYwFWsYv
/6P9XyegiVP2TIFzjXGQsZaiU7Lr4mi5stHs6i5xLEKK1592hKVdSgD9L81/cIOC
bZbsYiApa9cJ5mFa8PGlnMtnx0sgt0n5k8ia2KCG/r7Dm49+yfJ57HkAKacHgL0Y
W2WEFspp3rxO8ZUOnd8M9EIOlWsTjWfcFQseOgyoRV7zmggGBoMNG4lsozq2bm/z
o2OWTud+K8PaUFBpi8KGzc07lDsulaFdamWnEOrH6Yo6AoowPSBRjIlswx3F3Fqq
GX8N7keyITeJoSP6PCGboisaeLMFbfPI4ZHYB6MM8AlQgKXnsaz9l+ECtcbwT5M5
vJdVzU9TXdqCg8Bf6gpTjRB+WEKXLSHbTDjtHdYtG2cxTsbqySQNgEjWD4G/pScV
WOj/DLISrUw/GfVQIXOJ9PZhbG0Tq3gIlY+vPIM0tgx3YJDgCwN1AU1hTxjjedo5
G/gHO+y7sIOCnyvkckRyy83TM7qNxdxkjp4weGD4jV4XdOO1Luw1+UwMRx3zWD1D
VoL7ViY5vRPa4+tPdi29zUJ0J9R0VFUpFwW+qSQZgBKoiM+ayNBsot056Y7iDWJY
JscFWtIItvp5vUAF8XOesQr4hQkuBKd63vOOARYBD1QGVtAbcq9Ra8ERDMSKkGHk
qsNc/U/APSP2sDn4f4VeYv/3tTDC9iwj/nPyeaeI/3FrJ2yHrzMZR9EiO7dJ/pBZ
jqS8N6hfi7LP0tH1eNvJcKNhowywKhYskAerhumVW35I1Z5FSobd9PhtHWMeN1ai
acAuFH7PCBLwLlXHAkBy8N+imWPIPyIfIfSw34hbMHzDPCpH497icWxretogwoQb
OyB/V6gCRwe8EXviD2Ja8gW6JNLrroaRMC1ZvOWqGDadimlvFP2EYLy5lEwJCY/a
lkBH1w4RirKpFbOe3kv4KosW8iZ15+CcN6MUTAh/MyyuHHZt0gvhmpvI/TA2lZ5b
sf6TNQLt/Bq4iZ4gVWI6GLQCOnl69uvgn4vW1gDosbBJcAblzgeSFAOLeK0ucESd
Yi+M0dwW8n63u6gO6uyjU6moEMPS03gGRHiAkK6p81xAIJXlfwsU3JbOrg3RBMBI
RMcjsb+3EWb21ppqyn3M3YTo6yxCQxXrK4HokxVK0K07A7mpI9XvGBeVa9VXAf7u
qNPHuVtH08bHKWsXjEKIEmyL3FmqYNJB/3f+19HaOXCMyDmAkKjx4FJ7Sisl2DdO
mAyofp/z5bOMpl7baoT70VL0lrocyCbYiwTyQJgkZi/MW3s497fAu2+GhKTBM6vk
YUjjXhIzSanw2flRbfKhLYz3hsJ0a8XfK5yKpS1ohIwLfwgL0goiJRwDA2r+7TzP
bcD5IG6rkDe8eI1yt3T1w/CcqAlNI5TYw6ZJUDUf2qWsc/CUBBmfn1qUA7UZ5sJu
pB1goop6Axx37xMT4wDpkLnL15g9r1dttQMeinVRJB4p7+TMlisunlcoeTLq05OQ
93jB750PoBa0ZuxZOjtFufBSCB0JWgZqU+jyF3bHAL5dgn7u3HrKjX7ApwuxIHKP
pp74lbEOex/uuOi2GnJMiIYs8N5yjXBcTid1+1ir41eHfvdkHrmIdldsTe8IlFfm
8pZtl/SmFKSbKT2Kg3r9CIwesJSZx8iK4rL0vH6SM34QX2DCCSlkscnqR84YENT6
4io3BOLFVV0hOopIcE7J94t1pg51tejUZul3kwa0csHjfCtl7KnHJvyVYpNcRSDU
bXxVg/JzbeQJM8fnVWlq6zZlkFrmKtwoZw2QVsMeiQO87lTf83i/Kxxu12JuSsse
AAZDg7laFWVTI833G7Jydeo2WZgNhal4mgzoNpEWFQeQ4zoWtX9xLSYuPcD9g1B3
fyPPDgGOfeHTCvrQeQw7qlDYdU0OsEcf2CogfH8H/oPfod2aNIc3NheFd3mRok+j
VhhFyIGbCwJNs0aIujsGzEl9EnAL7oObu9YuhekNz+pslXxbKVzm7KyupQWjlotX
zC4LnRMQS4KIaqCCokMuO3b+Ko7V86uaoT5itUXA+8thkbVefyOajUKpQ8bkSZMS
PPBsKKSHIbviYn8t9BdQWDuyTrhrLn8KWvqZrYaz4dvylRF8PNqP9epVOBqcwVcU
Eo3+ZB1XEW2xw5oQt7AIPn+AZWqheihm3qqIg/3QpMqTp4Wffp5Hjav5Cy+Etwgp
4dKuKyLi+f9u9IsWEltP66qr4P76R20H+dP/wzNv4pTBglCNrtJHOcEWDCg3UP++
QmqdmNtt9RgalAIs4P3gK62+uj3GQ67nvGsQnLDPqc/8hZ2hJsIZzcKH47qs3Zq4
HkaeVDLZay/2O0m+L1wP4mW9tUF850fxhcnSz9VwJTAMQSnfwVzHI5q+c5hhXRAr
aXCf7hCiQQ2AVQonUTYz+CcYDHyHpafn+gdXLnnjCi6FP5qPd2vOfsgUsC4GOniD
n9ag3MQCFagf5YpUIaVVjevllmWOGXX/zR6hDlL7Zz+lcZOSw0sZNATZnMCUchIU
tQroLJ5Y3d1CUeFDBGxLBidx9UlVD2ObN8vbZ+7aX6U6PWQdKykNHZMp24Ihj4QB
8nyyrVYy3B26VLe1Xs2OVmQLX6xPBBrYj8sG7bosTdLPcBiS4ShhDYdiMwJf1EV7
D99Tx2p0FTnOLRzY0dIkhPAnaInLfqaGF9FIam1mLlV7e5VHRgj+on6yXudd6OeV
IVXfr5uYuq2ThV+DqsZzw8ZxHCIH8N/+TYgu4WnPnQ+3M8YjB+8n6mu7x8UUZQNu
fJoQrQDbBzARmrQpUEX80GCW5DouM8lvy21rbC5mTa9YqqJCdVZF9RUjyOT+Bjq9
JrFQOVD2kDDH1MMsNn+0+cm5ndj6ghxv9sBwlLJBR7wJxLfF36Ez3UFT4P1IoNwg
pRGf4D1HgWT2Z/JLYyjbVVtoSfWTuT6041HTR11dCr96e3lHeqL5pvI4bqZunpuO
CdRz6JQOWM6F6kr5GLlfS9O4qkapCTrshuubUTBSilCANkvAPWlcAyqSAhjUkuMX
x2zNG95NCd5Z2u7gDAx0O5RcNbT5NPSkuOjChje2wS8svBWUVU8yyIdcG7bNL1Ls
QIplxRJGb1J6Cjpuc6UsW5F7YLwZqExU+hgwG8TKj7nVOrEHeADTW+rgb0WgjMe8
T40BD+VF1IDqbSQ4Z1GY9KS6qGwM6Tuyy5PRcIrdUNY7Ex/dOnnv0KUcAu9mtEQ3
NHBr1zM6VN2LedmN6lVcR6+yTCo1JHTtUpyGv6bg2+3MmlJzslJ0wlRfUrlt8ynG
sIw9opZ+bZCiAt9gDmd1RD3WJK3maeLaqRjWrEdUcVUj5ImRtFkjGZl7lo6yvfSg
ROPQXthM5oM103a0i5f2ZLngVitvtQIYgPvBxqvzDZ6mXuqyV/VSdLZp1kjA48tM
XCYwttDIKQAnFtPHBClpvlQGUpCXWVWE+xr9b5ERcTLH6GM/NoxuxOeI2pm56tE8
1qWZHYc3IPQFrgJ8gUP0kJPKi9Eqw/3HPtxYTTOY6WR7faaN3JOhBoQt1apoEvhr
U6n8HwPQOXjtbo68ncgVLqM4SHhSsZUawljPhVdWFQp8kHli59ZyEik9sw2At8G4
QazpgIyv5lT7ksv9beEH6C/H51gh+5O6o+6Took9NNUFt+pZcwafTBOS7stwKB6O
OKbo++j2VwqI8GlV6wHbIdbCTSmzHJ+bKIMF0BRntjWhQNo4bkM8Ks3+IMNC9isg
u5/XKRDGHmP3yCsXBTR/k+Uup1CLBPhFe4qd+stErYlbpG/CDkrvI0R6Nf4utAKo
wCzvSl8ddZTbeHoW/FLHVlmSiV+c2H6W5ef/37FwaoXErhLKSlaZBLRP4jECmMIJ
OFz7zv253Ki70hhNMTtsMKB/H9ibuv3zVIKH/OGMeUpNdar8jvJUOn3IZZy1fpvL
gnJ+r9yOjd46POPwDHzzoLwbOpu102+aUoULluBHVVYPDLRgb0U3CUKqsIfaOXdd
cJFtjXj4BV6TEVVvKHE78jXcFSFbXhHc0/4LuY3wYB5v9Cwd2egsvXkKHRV+D3Wn
h2c1maU+fWRs1uEc1o1Ct690+pB7oGVPeQL4Xbv9pVzksk4RnO9EtlB7+CMpvm+Y
tlZ3ujaCYOOz8isg4h9ilOaNAA4LSUCOMjUQBuCxxMVQ1dWYvxetx1LTbKWmswPi
eyB2fQ4ZDs92I5klBw3S8iZc6uEsSRdBGe57iC6jZPwEmZOwTFR4du3dIWKqy0pV
HLf0B6TuMu9SJxPy7v1Gyw1QNC/kWF+GNYfi2G95m9ynEAS/rExXNpt+jNfWXvMI
8kuX/ix/2wyalx9ZahM/fyRvgMrjYBTA7rSazYLwpdyR687TwUcdA+QBW2FdATVC
GnrAbNadEcNdb/nb6PDley5hs5nbPlo6NF584xMuEkZqphL60RHYQF9l3+0BFTkl
+uYfi0eQ4EMX4O1VVhbCV/S7i9d+MBinMhWJ/L7gujKZ8goqi15wtc53t60x1pyb
orWJFt1Xjf8qNFKhYQ27hswqG046RhyiyzpWDjYK9A0bJO/eu5R6Ie1nnYD/MUfS
nLrzl/guI1izoHK28+LfM1k0eW1aJlt5iOZiYweMQ7LnPNRIah0f7BlEaL9wPgw+
VNI6IuE6kExITERRSiHNilT4jPmlQl6Y31bduUe68t6v55IUO0lU8iSJSQLeDOOs
fqHNBk+0pJQD5Kc14J5RhFH3YAhbI/1wHflP9rfKkLiyLYvW72t/czeLkCkub8gp
dYWqa7Q+ngIlBLzMiH2aB1NMBMuApOPiGvUM9hYkFRF+X9PI3AAAo6qa1Kz8vgnq
Zvw/qkH5KrTv48j0Kg7iJeyfaO+LdyLevoJOLZiGT66RBObs+Yrof/EPH7iznxW/
2ODLvaSu3HJD8KUnrvgdGFqQY+NuNnuNI+onhnOdhSspYtNtnXiVU0TluFLLz4Me
6VvqKEfdy07BwBoXNQ5huVzWJGvvs9zWG3KjI9rmTxA2LZ0c0DSk/D3ovOOBWCky
drEkbyeukjxMGJBH9b+HBryr1s+Q3fXkewbBv/C0MHiTYLUsR5Kogc9zeedA+pTE
RY4imt+uUx5iMagNO72ShrtVPn7v3pH3oUwyzXGI4SVpnZ+YZjQn5wcJu2QBXjEH
oNBypigTnSgRFCoKYa+3XZYnatIJdUVufE1rcnpXmic4YyMPJsNbD/W/l798gaAt
F6sIX1AJ3OiMa1aihE0+u9M1HQHo5rN2rGqN62QJqFVdik2BpBq87Ruo202Th7rP
vqS1wWqeu5Uao+4+qN3DXh+JGEF8jJfbHDBzcamu0bGKamlGIYQaBnCasijUlSkC
aNsVzS3uO1iJDGioKHqGylW/b9CbscJQYuCF4ZuQYsNGtiC8kJedvzbhwrJWUPHc
3KKECGNmT1ZEya6LHhvE3J3kn4HpMHlbcKR1B14rG+XjmlYYrsWNs5AHoiA4EjVG
7mWfDxDukJgMCIKVC9NwlXqD28i+8d66pK/XmhOtPqyau/gOH8+MjUt44JMpft33
+zUeqq0pQkQeuQ0VraM9jq31hAOjxDYUQ1nFm/5BgWM9vI8/FAq0YtcV5pp/r9ZW
pGDIVpwV00MaflhK5wGXcke1qVDIgeKTLtt0jwzalGsoeUiq0XVQCA51KGXuNSSb
IYeu8xXSoDqPNTmntOlFVBmectckgc9OFqbx/MXVTx97Pm0DRjWjJb5Ne32Ls8q2
Xm0X2R6yNC2cRt1nwHgT3xm4Ke3uQuI04Ofmt+KH7sz58cmqdR1WlK30lzGxvC6c
k5zmokXX87xIiFAtj9CUEjQoBIb3QwtifRwzjef1bUfcClB9sgIL4mGoe3IvU6z5
rEYoAg8e5xMxr6BQ6wHaE40RcaAFdvedaJD2Km3PHLr5D3n1weyFDYvIt62nwTNr
YGXddJ/DN8HAN6RA3xbMvARL9vXiqu+pNaB56Ew60ufDLYr1ghf43UCtK7lMeW7+
8P0QN4s2bFyG8WdSTGdkpIlGcRR60VX0RzNs4NDhMajgSCKbDzFSNoMOoEx7olh1
w0FSXdCs5QpewojksKMaLUcbWs0Z6UKNzvuq8aT7L0zw5SNinxoj/zYxBQyI/e1F
bNOGL6Y2bib/EiFNEp7D2Jn5N0uKt+AFnla3SypdAznJLNb3G/pP9xKe+0dfdQbQ
7SFxIuMWvcTgZ9xOPFTwEGj7zctTCdFvRK0m72ZZXg0s9H1bNYU1vA3/pOLqoYU6
8U3VGw40Vd2bZKeyZacE9fc4/1UJPCKpQuZs3jVSGgH+3yrxtHjmBGILTjutjoPp
aF/xvlNxLkfnhZEJ7L3m4Dp28MoWy2mC8KpwdqDdjervCDvH8lv5OxEdeaXqaGu+
rYTAdc+cw41viO9vmXukbRunWmCR1YuwUOD3lvLs+gQ16SvNymf36ro6VTA8rfc4
KE1uDJWUtyY8K/cnFiu0CBwUBrgYvegvJgqh580PtD8LoMoUc2u9vBohL/pdhkg2
b8bK/1DOoVve3J/p/0yb+jilZdAwfnBgOiM3HzUp4u6vZrXQCaihVjx5c/iVZRph
SuRHpXaUxxbb7Niu1On/60FxfscenAIaV3mUrINLtHxdv9S6aXv7k6fDKQrXlrFn
loTeg6GpITWQq+n6K7Ij2Z4Fz3X+2z3EOI82n5eGZUPSyPJrazRjhO2zq1Z+svv0
E5Rs4js2nOd0oJBh+3s5g+UYXS0SZIe1UktyHFXBNWZQnLswzUoZPsKWHE0MAfyT
QrSO1wgxhMgc5MNBsz7/m35bhJYuQJ8cm7MKiehprkdso/vmLo6zs7na/3gl+20F
+oMIm9YijRT1PnywqHkDEPfz5+eH6FTrPW4SxDSxKJrsKGUKWuxTl7DO0wbDbN6m
ym9ngG1K4bWzwWirx9FuxFFKwT5IQCaa9lixuX6QDQZE2WYNdTh+HBuQaIsYmLg7
YUwf+n+KKsTexs6pXnAXWsvVi1m3pDBeY8budj8ScQ3x1JsZ0TFRw2AFXoN06Srx
q7bBKb9+GoJw3THg6FEComDT6ar1ELHqCVFDXWYaxq/LVbRBlJmOGfhtVD6oT8XJ
PlxN8Zfc/q3fRBj76rwRtQNe5ORHrEu2/n9mneqXyS5iE+I2JFRwr7Dw4bHsRr4T
ZNLWnx0c1kfCI/bXPRpzBYAo0OMKhcCmHgYqcUpAXwyxHi+47hcFM3Z78oJ66vkD
bvWN8JcNiyv/VcnwWWGMTqK4bPB1RRYWI124eCnR3SUddNrDON75sEpSamQxVk4M
4jgAHfZ6miPr9LlZp4FsNYRT+tCb+A7SWHHveyNS8GA3DZ7w9MovWFuZ6ANh8Iu/
qfTrxQRs0VwmSr1NQ7ozKCchSwYzAPiBULCE+E7MLpEKigJgUYG5Xp1vqEvjTfpK
rt9lnKSr/vFssVurWzs5a/9r2t8AHhw0sCGWRKnxnEZpg5FgS0Eb2x29h9EIkJ3v
VQ0rOV2fe3DZyt9ShLrDH12s+2lXl36Y/+ybdp9lJLV5ybsUZCvydlYKalOcsvpK
c8gH8y1pYCsAeGfYdQSQ15uG+2w6DTSyE0SkPnZAsv+kfkd2Bdh83K28kZplb0Ja
8gIb9u7kFoRVhHHoNYkrPTk1wLteZFiVdxY3ceuB+/VdC4+uFVLnRDiakomXWmXA
GsicioFozfy6wnqTar+EjMs1PulhlcviSPk4xx6oQkfm618n0iIMgJUBv9B01kF6
Wr08Vh2ngV6xhfTAkCm5LipuJtKYQizb3KcjR5GY8uHaTHYFofa+6wcktVYBM2OG
9UOf+KtBFn2jMvDwzU/kyjowAJrPbhaCd14QcMj93gLz05wZ+53iv/MtZoySbtP+
ggcih5MqgZoENAkSbG6PwOpFeVXyZYEkHq5u9KptRU8si2mMqvyC97bJmmVU78Ds
P9XdTPM6yz1dX/6f7Wmx7zR6EbjW73Fw8oMqUTPUEW5e2yCKOt3XlJzs8D87lpfj
/HfaLSULl66ciB6efN8WGUPkxKWiftC0tTQ4FKQkQBMj8/fgWE7c8ycIyhVZh4Bb
1WUsXhg/M7SnZouZllszg2rbVg5EWjNyv38xe4MnJ7kM00czi1oKJyv/I5o8pWiT
QrikxWQnpiu+TmSVBsbbw0G3LYyw12ohXl3RB75QFvpE31rTpCxYEpW5hcqAIxQn
Rf31nyZHP1HTv2GGn6zyOQeUUhfFNium5iwmUWANIKJTGbvPu5ezyxdtINZ8BWw6
UY58DJHgB63p1JVZ7XWDRyt+mASrO3cwGg/RXnFXFviiPo0EerwfWM9rrTpchPa8
aB8UQaBaMPhTz+iNeAUr/5xuw3nivBFjE5TELryUSUq6rCkxifOc8U8lTGR6qxlG
kRFic71Z3d6M/T7wooIDXYWVDL4yw6ZwHRM/OCwVJHWoibCTU4pRh2vGuMZC5wNs
Xhy3l2/MWWnAx86nS3hYkDa4dn9UvpsfWXtxGpNB31UPD7ieDPXnTlCclYoBNXrH
Fujye6lbkAMYUIofOWEabDjIYQaLIk2HXQkTunJF7hVXyhNguW0IEdhtE04Ss6uf
gwaUiv3hOUA0iwQXB/BNcFzqUjDi8cZ2L+gDrcDhoXJh7nRaRY5kUCuStrJZNGWT
NH3fkVmYUFcQg09eCsS8RFnQDFbyhMuoEKfd1pIxb20TFJYCUweWrfyoPqSpUHgp
JLu/quwYozjRUNUpp7PnrPDhiqcw3hMfpy9kxMXiaL6ExjAwF3aAYcm1aDfnkByf
YD0iBlP0EWgP4puV8Pvm4UU3hHclzggzc1b/WYVHDuEkrWVNaPcdaSOUFYgMhVzt
xmTQVNY7cOb2K6hi1eXEp+ek6XHS7ZZ5q77vQkKM+8QnDxLPPhvcVBLVdGU4EeY0
0Vtk6LXZJfRrUQ9VwUINVjOgSVSNfJ4y1fG2aHbJ0uwO/AC3x5uE1skCMV6yPMOH
RQwITbaEPGlGIfizEGMqBrEGe6kJQhpeKRmf9WOEj8iF25BsUN8U5k7zpMlxxpGK
TTf0D5dfPV6jxFJucU6CTdhpPExo9lKJq8jIBHQXjtwJbdydphG8wO4zTCIVIWCu
4iuzWOS9NMgFT0jQKnjFXNTr79ZAIkB8ukCbJEqgssnsPndrImbBZnIrslznd0/w
X/pR6GQmgbxs/4swOiNU3Jfoo1Qr7qBAG94cFA5yNdIN5SadxuL6lTlbfk5GgnHc
eynKCNB6wJovacffUi2ZwrezLI/jpXQw/ahG3JbZ9z45JsWizdP5KJFfYufzEagg
LBgUgpgtpI4McIQUzb6mUJzepVYsEltga7iKEwT+s9FQBn/5Uem2h5m0wBkBL8l3
P4S5C5uCj3IWhELEcUPD74UuULUknrrEH/r5Fd5m1V0j3vQaZdslt6n5WSuVIIY9
an0RdJylTrxJ8y2dr0UaMfyQrSwiGNuI5sV0rryyiI92ixEujqbrOm/LRm3DBxF2
2OWnwzNdg3UCH6ZBNzgVA2djKunic/jaA/mOl6ptRKqPNpUjDd5tGTHuQE/z0cuT
QCG+3Buu492lM3j7w6N8j4Boh3hmcSaRsYiJehGtvuG9y5OM0TND0NTKlM5UqvWv
Ew4gWGyc2meWhcEW3pDWiANr3/sTtswgULFv7cu70jBceWAZrLqYcOIYdS38gZ7+
Og47t5Yb8CfFdU2AWl56u9633h5rgGUPg5GibLHvTeFyLgM0Fw/1R/zZMM1KK6wX
v0VRtYhiMWb5phKPCLK8te3kFDjAKT6cAncxhj5m3kYN44cpiYvPq4prbjd/I2EY
HFX15jjvjjolkUDD8K67KKn1aKiXjSWyeswvQvTPTdKmIvJIe121uMuXTf/QH45V
gzQWSGPW6HjnUzRcdcu68WE60AfuJcVp4r+9Y4SGLAF5arFiBLSUTeOpCN28mbo3
cIyyan/sHx/ksVeaTjNLM6uT1PT8xZLy1BKyCZ1zZGiIPfIFkQD9V0T1CUFPJ04k
7T4+u3/r3htau7wr8x/g6xk0ym47a4ido3VDFPLb5gNjqG3x8nJxmsoARAgEuUCF
gUlvA+PdFFwx36WH6xN4H2LLdxWQs6SD465KgdzHnTbKNfEaAoyzDHoaLklve/Ki
gF2CYR46c2tEg2mLyZ/iswb8ySrw7+JX5BVw8txC5Iw=
`protect END_PROTECTED
