`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v7X7+GoFso8CAFNxjmkER8S0MqctKZeYAEc6qq61n9/x2aNVImBpG2EwjPILfFuJ
6RVgpsP0DNEX5o/Kqg+7QEKs+8510wbgj69aIU2Hp5tHdIFmd82pYdC5SAPpvDR7
aa4PFsZG21WEJ0jxmQn4jtGO6D8Pn2/t8MhbQ19UsGtKsJBOyDVYxYH1YvXL2rGh
8H1My/M4NizrZKqrPHoMTMBfm3fYUVcmtrJRoj7K8k6eC+Qju6zseS88smD/R6IT
iAOmg0cxTqEUpzpfixw+Yd296vHOrkSwm76OnH4F90NUwOUvEIddkA4XMMaotwwO
onDzwqZ3Pq222j8xoPba/A==
`protect END_PROTECTED
