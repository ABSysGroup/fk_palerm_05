`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uxe1QXlvlY351cXO0vp+iJCXxIbuI1vCXiJJq3jhsICOZDO3UI5iINBN6ddsOjV5
iY+ZA0LlMqR7kFAAuHHQUYfUPZWIgiRMzk3JlWaw9RoOcxB59cFm/HrrcNGSarAe
jvaRP8YAEiCXh2FJYJDYdjyf107VnxR+ivw6vlPyn/Cqgxv3HjLFL90V5R0UJzhR
oQzY0m/iY9WppJv0ZohJicpVwav7S46dDoc+v9SNJETaL3sLeFdmwUWDlO6WHibN
KGYJcNzMVrs+p2GKblQwol/BzMBK21pXl0fLIafM6R/zlN+clUN8GKvwzHznoOT3
Q/ZlR4x2eVLV4tN8JX4lE0lbRy9Cl3oWnzveqqIEgvjK5TJPVTK08cjgkrngvxTJ
/6o088j4GFqjouFOfjTWDC4lkqteGj4BMQEg62pYl2b7AsZDOERiIRF13fyAst8A
A4ETqsfD5cBrtaREJLTP9ME8w8McTTe8/FKXvdrK5LPxSQwrxUEfqg+HEHSLOw3A
v9ouXrkDB4Bs1phwPHOm8SpcvTJsz0UiUCccB2eZeJBms5KPEy0fd7P8xqP1r3BQ
pcRG/FUQmMJjVK57FUoHWLKTnEBHOreBMS4UmL1ktXfz+mw4LmIGAYIHuZvFYtXn
bxdheWcCHytbTJMa72lEae6jXTOSKGEK5CC4TsluId7kCucK0GkC/ZvfPF/1hk85
jasR1joyaKUjomhQSFyAEAMX4n04iUYVAvj4jpB1zEM=
`protect END_PROTECTED
