`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4YNN5PAKH9FlNwHTIdhgO2nH20oka84/0cl5LWig2i9QUI59bmScb6z7ixBsTY9d
uJPbEbTRbuzI8ZA59TgAKQDEbABu4j4hvCs7dxiP4By/as+B2Nq5/tjW3r6WJTa3
E1hsH7uxiNkwRorov5TTKtqgTpHcGShoD4QIM/JhreP6nW1WurjSQY7whS7A2miB
BuAwjjDjpnve3jmYfHdbOjTxKg1KXXq+JiT28qvPiyFg8KHO3XJldrxnNcSLysHs
LRO4VlGVC/xvqsjOK4nlDByXz5qH5COmgidYGckRbmeNB2pdXv3XQqJOxfXt6rzC
DtOmEEFnkpqrO0nKybR724zYU77JX6K5DAT+/4MxUN9qWOtI8tb2+77YeJuAiGO3
qbUB4fV88/BuB+NP/BzKWmPrSD64aUcdnNK3okYKfimYhKgq+7SaHG4X0/hUk1MS
JEVqlMntkBvwGE+xCYp8JfJGWC5Ii58Kdsh31rJQD6A7zWH4/aJsdgYi0X8pLtd/
hwQDLULa3KAIqQcUalqD1Rrzj+cSgohIzizjuZZAAW+KFtNX0sFc5eeDCB1TBavZ
4dwYfS0lJnzzrYXo4lJqIg4YbJAXfguFiy+pTQ9GrMY=
`protect END_PROTECTED
