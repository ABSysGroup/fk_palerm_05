`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pGm7OZl3HtpyCGpphAgm0RPk5iAIkAYyCTkiP3fdiz8Sdu5HlPokGa8/6+mBJvPr
feHmkgH+NwEOWzEIAdVxJdnV4hZpqQQuOujBVdJeaLm0KWMCKYXC5V4sflDhra9r
ld6EzW7zSavV1VMq+8le33i7jlK0iUchwt8xW3RJYDBYDlt5w9gD3jhzK+OM44Z9
3aNElyPBdGv7/Y8vULU+hNZ3O/E6e09Ftf9xRT/9Lz3BLybww2xKAcLmcW8zXhnD
ZSaAL9xZt0VZ8rdk3JR0nFJSabDUw4Foq7bT+lEqeEESFphifAp0hKTRZLNeMqXQ
GF8PH9tpxKQ9OzkExnmB5iLOoO9H3kIAh1CTyyzTaI54ZXHG1epfHS8uhKaNEJAU
AKd6JS24hf+n7S64OMnboF1UhRP+1h88M72ZCPfkMhu1CpCgIn15pa9vMphsd35z
ZnqOg8kgfJqfD1V3ex7vKWDAlqs1azy4UeKSOjHc/Ah6XBbuWQRG2Wht7Hon6TbL
KAVybpx7OQZANBBSUDiDOrp22vDsQvLdtmfOk4BshD4XSKUVUNbFKXHMaPr6QFD3
l3vQgWcQDO3yoNPLQjZjtx48N63YzitVrcuKUa/WtoiGXk2ZGye93zgdHAmUCGQu
HjBVf3k1mJH3f8yzfHa6pPUlNh+IAbkjXXH61Eh6LEeiEAUz3skCAjjPSzCbNvml
4c1zYeOWwa+hScR4svoRbMS9+qbnsimIBZVPn+QE49KIzOsrQLprlVJ1SyRw0lCX
2Y7803lRQmeTODuZpDHIWoKrXKy8U2IrL7TZ44a8VU8FKuZJUTleIEDB8PA1yQjR
eJnrYdO8n4du2xFwtvB/NiDp2RaCr+Uokdywz0k69TB62Zk4ZCXln/rPHMP6OKMl
xy1rkl6sqJ92gw2F31EYwOLL7Vcfqp0JyEM+VRU1cTiluai4R8tghVOPhFpYUvyO
9Hp1dWMEbS82afWMbrcjpN3xa7HsgHeLLNMr58G10EyD5VtHqYxOhemgNWdDvcye
E3O342rHR2Yp7EjdL0/RvOFhv5v95TqWKUe2/Y3ebgeYg6XaAbG3xDia6i3+Zixp
AtnaStq259rECvi/dgS/H69DGb8obBE4Z7VtWbBifl0=
`protect END_PROTECTED
