`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EqIBqRTl/wrgOnTK+STH2rTjYQE1yQfFioHQrw77eclLDevAWNyZMWWiwNq/6CTm
UoUQcs8xYZ/N2HvYLop2rSCTG/W08gR96gyXdmdlpjUZnEbZfKfkzOSGv+AHgcNN
URRPSGgGApPKC3c9m/jC+k5rcGZCAmTaYiERt5c93LnqVTaVE8wXiGF867E/taA9
lHFR8JSY7UeC72ujrPwMPnawPvQu/zFR08nuy2S1WsAYAKxlLHv1r3iuGhJ9fGpG
aWPbg5PWRwHvoU8n5/pMwA5kZmkK5hxXCbn1kQC/fh8efnw/rZ7MHuskuq/GOxm3
TZ4zvCZhIQN1AljbuNzhylStCLa4yoSzr4UASvVi1I6BVoqAiMIE/9kJkkDOM7Ti
skH52mXtUCuZDG3R3fPELAGn8r6Nt+MNmySGyjdogRoJET4Tl83nHrq4DYXLzzzh
dDPAhLI1OKUNId120lkCe1bgCXdcOtyICHqQRrlzLwU/hSxEUqwjLTRoNfTIxX+q
3RYVYVNp7A2S/tJk01jVOK8kGIrsUoTt6pf4JMPi4OWblQWvrl8QRAOG7y+DLLvR
+7qzEaiAhWa3Nsum3Zxi2qUv8PhdED4+9y1PAiBaSbKTJsd/tqvHe6vCfMQPBjio
WJ578o1jSCDl1rMz3ho+olMoU4OH+cXXK3k7GLdnQAYWzDlsHWyYUo63ycZfVLXI
wtSuH2UEiu2V+lamgOggpw==
`protect END_PROTECTED
