`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tihzj8o990rEOLUpKf2WngxmQPgZ/pCOVZnsaWcISIxEPAxFKS/pQdHGHKPjeYpE
AlQtGC9LSk2tGtbCZ4BQ/IE3ZEG7AHAgRrnAH148dQ6hKGErCxSSTvlxCXB3QtWZ
4qYmxQ/1HlvUEAfGFSgkga5rYAZ735lR9T9qla3U6NKViV9SgpXZo3gJ/yv1RElq
TVPBs9PDY10Dw9cRprPGQkAwthidkmYyQtI7k9RKxoa4Wg4eA5CLol3xkKuhWWlY
`protect END_PROTECTED
