`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dHYGP6scAQP8VxRB66QKDu3qjdjljODm9ixk+F8ase/zR5zK37lVtcam8bCo7m7S
X6i+CGXMz7m2i8VEA9dMT1UlHyS+WJ4de/AXVNruMUpzkIYmoAqOGnYk80SAS1dz
ZwFQuUuMRSSQMT+dF3J6bAzTBFavg6CapN18OWwodk4iB8wbUrSwDoPXDrqcnVGL
O0AgVoMk2ngW3zAGa/jGLpVrk/rZwIQb61ERM+//q+HGGBkvS3EBcVmLEJkpkLa0
v6MTFFdjrsfB1uzRumlxsJK34r7sTIJrk3ilE5VXs7k=
`protect END_PROTECTED
