`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bGwZ5bDuD+avUUlARSbQ9d0/eQMGR6ZMO4Kstw9mJdhDz+CL4/HraAfpeSCGVdcR
2SP7/e551ksJzuHUYkDPib4ouDpMPfb4G3uW5hoB4AArElrP9qj3s5CvFy2MCJ3Z
MEnSmnnHs2YgTD4XHBFOXTJuk9nPLVIaKsjNqfZQKB30RU2RQCDp+1vb3tEJZkU0
p6475gRNs8cLs95o6WzUboY+P3kcTuyMWSnA9EmOjdKWj++JRf/ynLz4Vd3pho8S
E/0JQ5z3QzOFftOwrFP7iu8X7niUHT8Frmh+eQ7zKWhzAzfV7t8gtKV5ICE3ld1B
QCyJbMe4cqdvxtYd7ykXMIxxvaVEtYy4YvFtT1ue0bY=
`protect END_PROTECTED
