`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pXF/wOvrihWbCBPDUkduzzDcSdS+GWqm1tvMpMJdj7GHsIGuub31Lo1iLtniUhN1
Gq6wEraH5j2KpQ5B5wttq+tG9F7MESg5F7l3JGE+raoH0LKUwP9+NumtEbspOTAR
JcpVNSPCsfXx6Ls3wUL0saxGYG6la6Vzzkrlf4DJ4ZctZHUNmYR0VcrcoILpfQx3
VtUdssrncimfmUsjQAidFwNBrYErxfACwb/aurBFZRxnKOBewq5gqzIbKYxsQtcb
JcjaOpI/AaL/DkqLEcJ7FhtV5i/rcWsviUxLs5rEDNx22aj9Vzmh+d18e9ThWbfF
FGwakaUDCXL3jTd9veP6/J0GmsiTUSn/s1ywcRMpOGVjuzC6rKwZ69AMPohk4CSd
V0FQntYOmK6L2+YVZmwfQ4pv7GvgOhzSfjSLlY4Vwda4ysmV0oo8ThEWNdI3SpOm
9lu/1sd6qGFneLQKevaDU0GIhi5FoZ3pDej4WhPeLd4aFgfntDTbG+e7z16D6jX5
5AHU3kUAWAgjz/x9TFo0I2kAsdEMmnWYau+BOPKTvNkIuVZ8YqP1/29k8GoP5fnf
hQWwMgFh1CbVasUoY9QTvb82rjMixfjNhMYPcCl/t8EIGwSKSRaR+ovE4P/WYebA
VJ2dTjmTxCkwJrus1SzblzrEpWTt8ho+gPbfdql8LvCUmgtTyxlZQqO2EAQL/faA
ZpIia27LLVM9kwnAQjn/r4m783Mjid+pXU4HIqtt+pJydOv1BU4TJLeNWYCpqjTy
Hh4AZG2gmWkAX/xf5viruEXxB7x9p3fFuTVmNSo2fQZljvdzuDfPmUPHBuK7qcYh
hlJy4OOXdnovLMe3f8Xm7+TH2RY84sih0C4SO6e0reYxFchP2i3aqv8n2dl0lQPJ
0MhFICdwO1If22GcFyLifuzj2yhNFKFxSoc3T+gd7dprmV4Fw6HfGlhAlOom8x3E
9fyWXbWHsXQf3knshoyRJdt2VtvL0ypXDSCLnau1eG7APrxpF7HpNPosoxZdaxRw
toAX1ezYMaUt1AUXB204hwGtZaFKSbrSPcafCe0TvyvINBTxSKO7/Lzc8rZsQHol
VaP6LI9iqbqqoEfrpGqGD/t/Q7/lg1d9ZpEyNpd7TZEPAAaX1MDfpoLgDSr+KsiJ
Yt4N++SmNN+e4qqXRdQBEBvDCxIHT0T97zzU4pQs1ZXVhc03Ul0b2bfqB/aIGV2J
g2kfhfiTNsRmGHbHbXrfJL3HI4OEEpE/hbgRC8hrIZKshQOfFomhSyHgahwA+ocX
nlOj7WenO4iv4dYQIX9x9syABUPwdhzJyVd1wZ+kb1j5EE/3poV4jZ82YfeTMvV2
EPN5D36X6o+haALuG9+gVm/bZeZDWCxE/e434A6x7RvCouaosgNU/y/PAUwy3bbj
MLfzQ8ZOhC9/aNTdsvkRHdkCcMerDQd/ROrd+6qKp8bdzXnyBYne+IJj1WzXcYBo
kOueqO2jzdUt/Du/GD5xd6twPtGOTINWg0uyAgiDIQFtlI8BPrQBCTgqhY+zbsw9
BT67ed6dxsrw8wfoC1pNUHX/tNrMuFO8+VoEurtIl3w4l6B8eaGrqh3wm3v2JEjq
iAJkOU2Q2HVBnzEPRrGw3zFFO6LwHIxIqwbnr8dchMPevexOP28ojzFmFeN36Blk
j7jMqcM3V0lrsxN27mk7ouDNS9rIb2JcU/Ep7XBSzmOXCG9OZRuN6rPVOLumuDLF
in0oQpbmOY/D9tUZXn/N4oSrWYvD+vWgs1oFemiBwaBNnVPuMYvrpBDAoijhJr/1
4+QmYHaZC1HHxxpLfCsMd4lHC/xzhvXV9VPRypJ75eo=
`protect END_PROTECTED
