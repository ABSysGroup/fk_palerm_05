`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LpJv5IHflXBp2oizjQVE5zX+8qnwJBplQTnyUGJ9D/Xo2GjBJ1GHEWPtAHl4JDZW
Kps4GuCKXVXj403GUbWBxJWjCH/ztehTev9mCqjPy1lQOpb5Gqzi2dXl3YJUZ0x1
DLv9Kns/hwqOJfHZVW/0cnf2tEMNyVDPNcZAnNASfFbIsqzk7/3NqXwHqdt56agS
aFXYlFzgC5rKeWSz7Gvs7z4DTkkQP2yS3irmnstRUbORYHwxn1+7deV/jAAGOrlI
WUHdFaMRTlfJ0uBA4WGo8lTjmflVikD3adYwEbs0X4XC1IKRWgBAVJLyffTrRm2b
XvpDqlYYEZzizkYRMJtGhe7r05NmiTYlstN069rD5zt+/Zgl9W9eZxc2313VQMOs
15Dy880G/DbAsrpXPi8V/6lzugFS/at52pRaBx7HuN9ti3OP3GMG2TTeyNSOaT2W
w2bBOynLfT6VCeL4B7ZtH6YdBMuGvA0QaWhwTmLnjCxKL/9JwVWGu4VtuIXgdkfh
PN6iU8s1ZP5V1A+Ttjl9KU/BJT3+WnOKMsTan8A0eRY+8yYynxeLEY2Qfa3yY64u
l345rdpCJVSDpuTAMO58bZaY9Ic27MpSD9+/b6Z/WImeA7f+ZPR1YXuuxVsBsqZG
dj9ZmcSaDmU3DgMFIj+e3MXzonK6P8ZYbEsvqI/TqRsmkyoqELad2GiLttq8Guxe
BTcAj6WNpsIjwpkwOvJhL4IgZ8VRBTxu8wmbtT2dM+SVoGmtJAZNd/YW4kpRZOOK
LyApPXM3UaCSVYSYaZu9LPsUCtO7xb5H0PHZZc9VBYAETh+p9v7aXtkL7xVn56MP
prkGCLWyVmOghM6zx+x/qg==
`protect END_PROTECTED
