`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DoB+yaKeUNNrsP/j0qeaKPZgRj8D7Ewv9HZ7Xy5cCjWSySuJQRZSrI+9vUd2KE8D
V2ERHQp5vetMLjZFFIVqNsh/MtSKuL1eFW90jihsJdy+KRagPT1Wp9r/vXUa6UQZ
/iNrASnoHp2jVCjc7pxlN2U590Arfp5SrAnNjOqc/E1UfrC0UYSv0xJ5jsEV5Xud
ZFtgOhFWr7rjJ3KHmvx8SgKxd/a9lOYncvFDWdUrtHQkUZo0Fr20JkrcJFXWiwuN
Tugv/s+MbY4Z2emX85ViMTSanRGCbbY0mtIqQZxev9TK677FJwsExg1jKsIlG0e2
H0xcGnbkPju5HPQxDByoccbwBHoFA/VnOlWACiC6ir3cKqGJDf2NE7OeAU3MyhGS
HZh2Q9jwSP6/OqPj21+oykbPFnKukFkMxuQJ1ntxQPi7g3uQELgpxR5u7uw4TrP7
6JlwjOXMamL1eUVG83ikmYvlql+Un7Us7Z86o5wCSJB1uGTvqpOyXI6JxL7b/KFs
hMdPYK9xC9JiHW9QS8S70gYQoQh6/0W++sfS6fBXf5mgZf9lZxvelcKTHJSV7SHA
fDqrbSdRPOLN3StjD2FspOcpo0ZC2C9V1oXDziMsRVOiZkA93CFaJWVnr/uCVen8
VQnEokhCFuvvVKOUF5EW4oe9JCPw3jpMg0meMKlzJvKbHSDoEjBg6Q1osn7OmEsh
NEtsoZRtM7Jg41SWMR+YFAAGwKMEf6TMai+/odWReHtsgh+ULj9tBihbnVL1XZGZ
RLceLw4rG1U3ZZm3V0lUg6SnKtmjmtoXzWcJd/iTmO954LYLCdCi4UQNFCzh16N0
NFtVcYLi39UJlnFs8xZ4DONvnCgN3I4pHwO6gvvMPzZxf35RQToa6kEr2Rf0Z726
TfFYWgRrCrUqu1RZjqBx4fIRxk/N5ZCXaWZ/0lFKb9o3M5/YlNnaBfJivs2+NmOW
HXJXX3rrKowCm+WaH22NhUpHKJWAt/nv997jrnUCe1fadnqgtuIEHl6FUxL/DScK
oRdN8X/B7LXqu3eZBXOB2g9NFw1+BgvP2NWoLhVIhhRkrjcfOZNmUjvM1JI3J2bA
YSjbzzmQZkkvA4vbpNYYcQOomKzp2Sf6fMT/5r0ak7N+8W9+93Mqn5pc/aAK/G2y
FpHinoSqUd0woc6WZYNSiSLw7ujFoOOlVNDRLnsYHocn+p6DDcfOI7kbTy8u/b72
eXJQWE8FYBeqUE+GByeaAFUUjHIJUYs2XxT+E80e75ZjEruGZp1D8xJTOb4/32eM
`protect END_PROTECTED
