`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
98QoYCJj0AZNix+fpdhni18WF6ukTkS5YdxmbFh+xlB5rLIr/z3DwulU+qRwOXEW
/UNwrH2nqah8/C/BmBuot95UZB/FnIZZqLNDn6Dej2C+6MaL5QFKX+xKDGouQN8n
+I/cujBSPh7Kh8CaOeKCWGzuexFJQM3xw6caKqyCCMQL6DapQePgKOjZM6BvXvw8
Ukt6nD8vWauivqhnE7fqflVND0chkkCRF0vTSycWoGRykbcAZJsr96GKRB9xvJSY
EMIzsxmMihmgSArFcuFsDZWaycmGCDZkiqyC9oo3nIK80f+tRle/OMHTHIHW4jKd
/fJkhEQa1sGUQEuXi5eiEJUkN//iz2O8o5rzmOyCXPmoQQNn/5J3WYX4Z1aQXiMz
of+IjAMPVXYMCXaK5AdlpzLSR3FS3s1aL9Bu0Lt64ApiqxPwp4qtHPKnwnW58e41
Fqc9j4zl+j336myjbJculWRK/dL4GiUz5WANTuHQVTgclmhL8XQ4uGqvHXlyKhYV
lFgNRTL3ynqjSr7eO6+YhQ==
`protect END_PROTECTED
