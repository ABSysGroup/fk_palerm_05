`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VwIx+m1wlfvuju/jFnqqMRqHFbfd49ggbyj7sqWs5o3ktVTO8zg6VHoMCcSeU2PR
mjQAewNNIkEc4i1FQjM6nDJXb7iu+iyZ5cvZ3r9r5MUZXk7OGvbXqe1vRXNTv9+/
ZuNtwy8bW15Djlvw8jPAQPoSkQsAr4DsUzmwzrxquMMXx7Pl+3hdIQ/rTT521FwZ
IYrwayt8vblUegyuHJF+1CzVqI1uu5I8t6fKPHDINg4hXFA8mh1sFNMCapZcq8Pw
JhFXmM20BYnCpCDEdKgVbDShvYFGK94flIhwC7zxCAASB3p/103cYmPbR+wrcarp
TbHqbUgtsYMtQ1k0H7cW1ndSeL6mxFI5lBlWe2pGfdwAJPRmr1IWljsVNTF1EZdv
ypKj29dmraisLMS4lYJcT/Mvve7AUVkU3DjHeYB+OXcH82wNI5ErT0VhCUUJ/6ye
VskXwvmwhP9tJivs8qNLjXKhCtJQ3EXVYWW0/t6TX9lshGi1T6NYwzojKRvWTM8a
g0KU1sgMUPJppANmQmNifHYt5LC65TgW9ip3iveNStSWaEThRupIvycenzJ53l7Q
ZxLcAJXeGqANnBQSKGI0e1j6R/oGd+TtFTNqdFdTAMQma0dJuKVi3ydyTRv3fcJh
sLT9e+YrsnP0Gz/CwkM7GKQeF6imvV1TZGAKq3a2xBKPfred5GcRwePrd3zbG3uz
A/cUNq6NVoOzWW6XBRCc6g==
`protect END_PROTECTED
