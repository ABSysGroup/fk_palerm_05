`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I/MimWJxGFjKJVlf9BGOPZmqEANwY1JdDj1ecUj48cCWv2bdjfF1ceCGt3RpPhSF
GhzViXlZZ00lboJuFaE3pQY94oHzgaFKWX7pqOXnhKflZxrwRJjQ2tWoSGzLhHQ7
ZKiVRuZnasQrvCGQ5XoN5RBSE4dn1Jdo4VJ9k/tgYG3SWR22Yxk1JnBlgtr13GwX
aQkKd4v7XTxWj4OC+3dW/jLhQUieJE8DvMQPK6sXQgnC73Ub54d4URTzdU3g5/ML
E58RXytpPw42GfrmdzUmpQ==
`protect END_PROTECTED
