`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j4o7lfbiH03gU4haUiAfiASn7a2RtboOimHRXz9eKNyUFEUgn2Bh++Ig82VHOF0Y
3F9doZF0cYWztT/+slEyoIUgim5xmc55cLw9Qbgt81S4xDLNEossyBzEKzBvqgvi
Lu8uKERoMYhGpSUbdJitDvScYeXdacgDmgzzK+azOLuoFyn6dXNweBcbTGZEh/Qc
aBQ2RrxJlWiO1q3WHD6dE3yHm2g3lXpvjYeRnFGVIZaQTrWTjWwH8SiiIgyAlI6J
AtA3DHEYOGKi2+eHH9uQCJ7QqdLAcpazW/B9rY1rNkKwPqC4gPya4kVgacSr0dCS
bJZuKpcQCapBInnX56AurrxSyf9V9nlMg5tW0dqbokxQzrapypx6Lm1JWa98ISu7
5pLLKdizEesrZlKp2yMfSls/zoM4pJcrD1lg2uHgcpp7oMax3jDaE00MGHnCAgYX
VDuM0ajDoeJ+6z/MUdgI9/lw+KTImYUiOnmfz5PJGPBozFHSmT9HE0Cl0de6gIRI
Q1/pKalmSQAKlOZgLaO5CHkbX8ulqEI+BX2OLfE45fNEl7aqfAAqVwDiw+AWh8J4
gzt0eS6ge5hyW7qJmYmryWNrbpMMgYRHTbOzMncTg7r1sxrveYfs+ykxDT+XrKa1
`protect END_PROTECTED
