`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kWKerOAMy7+Q36zuO1mBNnj1b5AXemoEbfEyT5C650wkBDXZduVd/B8YoOPsauel
bN+T76m/kPAzJElrLqZk30MyAuMOr+2OqAb7qxd22aR5+A7q7NQN1Jl6vPVn++zw
7ARzdVi9yPF5H1GX6h5zMo06ba+wTy99L/nV6R5Fs99fllPHhVJJYG2mg1JeNptI
XYs4EtR5q2EzfZJ/ruBtvCtI9MlPLfA/Salvyt/eqDjr9cGlu0ZXLR7uhX6yjBhp
W6S/Ve/YX2lbJvylp48nTl6BbNMPdmqOwEP/H1SpZ25t/uNJTo1SJ+FotX4Qlz1E
XX2F9zQ7kbrsib1sZazrAy9YuJ6KdsqyLegX3wRbdFRDQdpzTZt/uv9zbXKbkKXo
SAxkPsgONm4usYpn1YYE8nVoLOPPtouUqqxC1zJW+F+vLQLlHuThMFQ9o1ZV+q++
ojXU5jmQmMOKqrYTiaIX5JTFf5e8r7P5rBw2r1mn5fBzA8D+iQMZqtKJxMVysFrw
UjFQu1JpX0DSVhRTncfjPgUuc7kCFvtPkDE44ibZEyG9MxB/ujvokl7A63egm7qh
D09NTWvtybnx15fORWHKbrBmD5A0/3NnGkOg8IUDlQYXAVZt3KDVEHwLuj3oViRa
Hoy6q70BLXNpPd5vi1u1IDQQdfalWS0DYk9dOOKWU6/+3HYv+GaR6u/pv5YqGA0N
syPORkLHIGkBfea1dq4/zAtP0UbFohQeqC0/VopHnlTDlSUnpE5DfbF0NuPm8Hbr
wGET23s3FJZZYnKFNnDTRR5F4UTGesTVGsAspnD5Qw20JtGW3JsDzW/0Fy4StzZr
tE9VvHizDpyjarlRPonak25YTp4UB2p+nPfczQJgc0asEIyYbAKszocO8gA+JbJW
XdQHSl3pzwBCenk2FHl03kbTGC2zYAa3lC35/cpUAjfF50x8adyZQQqRNtYErEou
GgTjs1NPNtAALrhmgVdM1Zf/7RyvKXsHz0BdniLbmLOSUyTYxJL0IW31I2vJy0uo
Yp6iXiRYgPVu8TEvGi9upQ==
`protect END_PROTECTED
