`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qbc5wgJU0GDZLwpULKSZa6T703NctJM7PKQUU1hbbwT3fi3ug7Rg/YOM5MZeGSdJ
RM2Ka+lclZ3SJSkxUYtWe2FSop4izwFFzDpnBJZvYfjWeKBTc0MCAL+PtRbYMURm
TJbuVW7qpMNKaBwMf0fQVx/+spCRaDtBn/xdIJuQO6REHjqoYOiRM8lFwAXFue5u
c3tCPVHONvbRizM/y/gRIHh+BPtqlHDVne1VbNz1ZQZh0C6u7VgldxraIWk1a5BB
d5j3Df9C9e0h7svqF4GgnIjAvPvKpDPAyrsGauCOz5qfRhynybXdKYe9iBgGlcwc
oigUd5MjTPfIT3mLg087NUYBBgIMKuD45UrSsja82b8DE4ElsfHT7p93ksh5e739
thIRi5VUiBL5j2kMmZIk/z5Huo23NHqz8VgmCgn3/s+ewD706TyVGK9utxCk3ksa
uYtVfgiMoA8wwrJSwNDYWUqPa3JdePEFBPN2CH1c5YReMuSDqqR8tVMc9uIUQNmU
OYj6UO/HIKWhh4DLYfoe+A60NLujc8kkINljC2nzy8SFMK1TR1M6qi9jcbYlNJJg
`protect END_PROTECTED
