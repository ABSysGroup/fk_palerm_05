`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bV5yp6VCgHRUC81riBN4easRCiGouR5r4edjfboLo6k/ARWBlFif33l3y5MkF+Uq
zLjKwrNgsXy6+wk340YTdaZmNZuRHaFuN+3CKbH25pSS0gvad2vvhgB/gG45hzst
Ea1pmS8/N8RoTjOoEBTeZ3eCwkKImwJ1WzLcVkoNOj63IY5CLqeUOI5gvU5Cye2N
ztu3DzYdSA3hJxxDMCdbbe0I00skn/Vw87c/yZZCXkuaxlrjrrfrLoQ1U05Z0zfo
dYi64ThEfoX83PNFHenY4d/hqx+uPAoGyb5pve6Cw/zH2lsMXYtb9PCQR89EMqZw
NQyaGY5sd1+ZJb7sfLsYFmVAg/uagPc6Jfctl68zw1mwCz/Th0Dt1cNoGze2M25f
3QQNWvtTd6xfuTfG3yCHSN4s580jh/QkzVoXT1lPr7mMBvCa//h4kXNDc5EPp//G
QRMQUiovnnLft0+j1yC4VqCKyrHPSH4y1w7XM2UyquziTNpnTWCPolNozFfKyU3j
ldU0s+iuFMQoLvOAfOFLjZFzALk8n27iRBhh2HN5SHHdsi6B/z0makDnCxRRiSV1
oTDiReAK7Tf45jhEB0e2qgxyh+Wrg9GVxbowT68WghaVDlN07HE8TQhLrzXJedK/
0XLsXRRP4IbXOe+iLgX4Qg==
`protect END_PROTECTED
