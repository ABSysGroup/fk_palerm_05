`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oi9UgLBQqkjbyVEmQKnkfGxwl5bkorR8Qzl8yK2nt+Pjhq6ZJ1Hz4AY2sT4mQNCG
i6H/bXWKDlDlY1BrB2lEcP9QExdfTUy2iV6N1N1aGd80q17ofUwm6hPH8kzJmdfr
5u/7mBFlEeTiDoxrxQawXhYAKsSG9OVC4lqSICeNnCldk8EXaQ25PA6m8fd894Ga
3jZ7qyWQ3dFoIHuc5H5zpiYqtmtBhqVTEQRz1Gz6UMo09pWgKu/sflwTkxCQt2xv
SITOUeLHSOp+tMgZ06rfFyLg0jBaRSiPKW3eM8ewzrnnnQIcQ4W+ewUW9HHtqbut
wKFolL6FWudrDVk/iSqpJnGXwElYaCeyj562G33sQ3Ax+LZGrNPna2FmAxvxmrD8
VNeOI9dm96sYQfKjJ67omN43UOazbNZifTSBQDqT9A5lCdJkmrF3Gmy1Jeh0hbbZ
kFkS5mknPo+t1MtZWySs7f/RhjesLe7jX7U25Ebn7Ae1hJS0KhD1Fi0SN1nsRPpi
rT1vDZy5L6mlZt02kC9lMniREr70cUJcBqWJWmHxCnN5yb289DuK/VQFLdnU/aN1
SyI2XaODNHzWzFqIRFOTvxqDOG3W+M8s7weZaCSBRfoD+9p3Y62LwRm2lviBLVu2
X4ra27A/c4EMtSZiZkPLga9kzpLoEVze+nTwFfIlOANqsFTXXRUIPi8YmuhEYdYA
9IuWPbX1tK3vK6oW72wgeVnFCvlPa6zeLS7kPRxLqgexM5rZrTKJHFHUmW6gNY8n
KQvdc7by/MjEgCcw7vxwew==
`protect END_PROTECTED
