`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B54EEP99kg2mMbVov3wHQZn9dYP38YJ4dJyREJSxGfnk1mJAPtyt/XSanad+dRwV
BLlQLiW9YykNjGXgf28caoxZJm23XMpAlqarRiVpLZ6qgPDIqGvfcnmp9SUIyBxr
b32kd1M/tcG0V7+VpfNf6X8TWlFy7Dgc+PLP0dNZzNKJpDKhNHoMTHqmdVznmnkA
NP9JYnwjm5mdnmvObguWxz1MMFjcQ7lu+lvbnKQyFNh9OyiQDILj83kKQLVpiHrF
0TmYK4PKxmSV+gwYeeCxqSVS0Ej+aTl0Q39I04Hy7hl3MDqnhsaK0xxIKYcoovKh
ATDwIkV2wn2yeTm2Z/XtpCjhPqSN6+nvi+WPi7N7jZotoHVRcFzniHXCwiG+/nt4
5dT6ul+3VbOLP7Fcr6X8VC4eZ+jfV6hr5Z/yyrPy0jnn56qdJ5daoTj22J/N0ynZ
`protect END_PROTECTED
