`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C8rN0qJPOBE3qJyZQK4NyDpauc3Yrqg5/o+RqSxaTgv7OsoVFIT6FolOu8+hukHu
/vyBF3ntQX9QN+769j6Hu9rXv7kARbXnTx4q14+I6wF0sekpbFR2jB41ARFI9Pp8
t6fg6zjsgdstCNNgf6xqwK1BLq3CFHHsu47nxi4ZEZyMZcJAzHRoyEz5mKbxWqaA
UeBQqIvLJiDzAu7yQCqrqH32Xmux3TdAN7A4cnwXgNRhvtYTWRx8Il+RK0uxR5k7
zIev+eyM18OFHQgE1HGDogNPyDq4PxwdFMhCecVU2nxYTyqnZP+keuY9ZGQgW7GO
r/egjE1wCXMa4BJ8pz+uRfnNjxVjIto8BUigzPqnmm9jtF777K6yzpwa6wzVGNMB
0u8gL1Gc46KYoQHfi6XNJv7P4AfFgHUdNVoL7xlKAlNlHCrpArcDAYO3kMs0rv4H
nyFTkoPEOEdiTxSxXR+CL6EgWYZFvTR9wvWu/YvD9Q1hKh/GZHMcBH9lTrutpJC5
5634N3S1iGqpkJ2LTAhfaNFc71vo2NVwGtvDK4BlXyZ+kqvIa5JE2+3RMvvu7K/1
mwsk4/9aXAluUt1ISLOgdTUG7fnugAmlOe0wGvnRDlhlXBMw/8ghZ4NiBc5yqfQ8
fwxgotiQpNJ8xxpTL6mJlcp9WJ/UYeGT09k+s1etfcKcMu50cwulnVlpza4dZPAP
f+RjtAOrZax6ufpOjpqwevlGpc3wmrHFLVfqT/J1b1RkqLKBRHbldLzx3OD9pUN+
//GTm1xnTxd1obbVx07L85VXBznLeUBTO/Uh5ZNHuonfFwsQyh128CLzwGlcZtQl
5Go+uHRxBy8vDA/oY2VSsUQGrNItw3tB8C2hHo3+9PQmPdnOozVrht2ZaF0fAwsF
sTuyXTIYsb5VhHU6T86Z0voL+b2eqMh2Gh/mHlOzSO081KrsnHZK6U9PCXUgtJqv
rt9ziOBCq2d5BTHYnDzSAwZY0lFRHydfFo5K07acC+Wz/J5uo+HpOUl8v6MDlock
Bly/+ssNrPql7pmReiKAT63T5UG167Sv4Uh8FOE6YIqWaWl8Z6/nA6oc9xQpojh/
YdnMemAKAJ6oug9QIBXgksgh34zSSIwrDICnhrogt6mFj1PyB+7g8eJ0cOdilJsV
OC8JNSax2HljX1i/MSLKgCVpJlPOyVcsgM0LhTfl4BNcBZBLOzbw+xfpJRZVfOAZ
j6Vp9KXZ0Kj/SJQdvFvqC1wKXijsFRkLuTs5vD7bNhgLGwkbQC0uz2/wterw7qFF
5GaYGtXqZc1ybzyg8T6ttUipQjkNtKjsxuNSpGxwZIfjLSN3E5AilIKsXlYPazEx
/g9WvFXFYRpQQQc1pE5QQYJ1FZ6H6AMKzdWitL9C/qWUw63LTRVdB87MAFPkSySE
7tixKdQ8+g4GYwwYXQVydYHXfCoyeIAhxG4+5iqih/uZTK0KAqR94wyvzq3OPv1z
FnAmdpdgB9njOYYQB3sCp6XqLgVwEkY/N5iRjY7JIw+vFqfeSeD156XtZfdqhLcv
fkZI8PxdyGwDFDcAH6n8vw0JrOOdjqyMc3J+0W1Dpt7GkJBpHNa0aLrjAoR+HlWw
lt+QJHzUuiJ9LoJnaRi9MTCc68nagF2/qUP/4VNwqRlDOwah+Ip5c6n6Ii/xiVwl
IQEQ4flBTIZomz90JtrS3zT78lhWcrBYGK8jk21+mFf22IOsN6F97f5fqMO/AWtE
/VGOG9d5flp01NRfUAedjZk+emCxkfaBb09XCUaxC27/nAiMudMXO79qQVdYy8MX
gp1PhuWihacdnO76OGlQMLi1wDdr1NA3pjpjLxulOjBRC3wKPJYc+Ka21UlHirM1
OiUx2mQ4vYDHfuSbRuxqdJy8rhzzO3C14cPmD73Hba2thnJq2nHlEbLtW4pfINCY
7d+3o0vb1/Gkynz1a6gdr9ej4qb3ESGCFjeUyBLlkQ915OgRxDzNx5weZLDgSv3S
0oM26b1xH6/nrSf8wUvqPsdbLd8aJWc4m3m94NuWoMKOPnePzPeqF9+RZC4Lgl34
EL5pyp2xTOubp+bOLEWIGSwXU7JVgOPTnH55LSrUFY2ERv0+P53NQNG2wufArvuG
c8w/TBo1xrNMXRY5JXJlGPdbA+saEc5Wfzi7vdtKZABG4ggJXwEmdZAtRRIHWkDu
oSvGaizEmCl4C7Du455DRxebQvDLreoZ8CFGx/7PWUKwSc3T0hyX7dnXiXPXq1ia
cGchSRB/up0hf/0BIV9Zq46oWIorILEYptABqD42dhi9GrRx+ND034QtHvUdPXlC
CFhFJczJXccpaw4GwpRb4pVybNSsujSUIQM7FvXTZf+apjCrh5sVJN92KEQP8YpK
pXcINPxk6DzlfaVObgGauLgkiiRQ2MdPE4X0SX4KnO1FD+Ye1EMuYQHeWZl8bPN9
Gglfx9s3aNP0+eX47GSIJCLeOZSPrNDPaQWFIKQQlmOHZPYIUtVS5PW9xyhfdAK8
1MS2Kqw/+kQcsiHvgmXspl5VOxaN+jkzaiC6fWfZAGvrFW+vIbtYnJnpDK1AZwEF
WqNkyHs25af/B9TSRaoAR8PnauStA/0wYP7HVl8PFdbqCr2HA4MpM1wXD1YJ5fH+
URvJh9SnkLBgTMU/QvKC732ifLQiiWCuTaIf0RZvXWQy3d5mksx84MBWwYWl4t+l
jccTnHGjbhfy/bXgT8jw/YOR63JCORqLcEPgoArHO4DnXIWsPCHcKmC2w/AVW4Dd
qG/RoqEVmuQ6EwYG5o9c33adve0Er1Mly/gI9ObjSA+nWHHOB7LUp3xbZQQ5Sj+P
n7lYVP7mgBZYP19u/UM+gfMc+z1mTPlo16cP3MAR1i8tBIaaCW7j7v9u2eIVtp2l
jTVg7/GajCwGkJI+2Kv5ZbnplObBb5psBkFrNPN+iUB6PtF2QdqbGToUfvN26phO
53HDg4cVUNbNP6fQ/B7C2+93StcqdJpNyen9Ches3/kiHW2xMfRc3nJT6HzlXQRx
QCzodZGK94gCBwxnNSUEt2rxgJXWVAv4AxboMIfwEqjU5gMzgeUlcy0Djsw4bCVA
sOk4t+KKig6Tn114YH6AhS2VZEp4aXaFZoqb/KfxvDeIfS5365+l0bx3ql+pkw+D
PFVdjk0uWSXfoau6Ztn7Xzh6YyqXRDVjF0y9/2EUvJuI5ONwy+fT1SaUw9qptHu5
+CJX7I64S5iU/yEH9egIN7J7ZbNE+nD1L4uBJhFdIwmRM9Ytm77x01YXQYnxzA6l
02CBMJVFlGRBXgeu/wd0J2QT/jALzAhP4lm4WP2e0Ob+4PdFcl+AJbdKrqr7yE73
ebZV3jByCuYc8316dbAF1YxFdN8x4q2aThbsqSJrtyP6KxOwuJ05T00ewg1a2Ws4
gj9EmIReC9V+rl/3SO+I4cKIOkkyLH9FFaQQqWTXtyWrSM4LWDMRKh5f/DCgo041
RYK3RmkIHFyd8U5HPrL31Rt5mmZvElkdbvgHoCaGCSvpMyTL3pfPK9SCjm1yjV3D
S78EzcEb+m3ODPVEZzpfZcbZPbjDbL44MhiEMEZbAPoL1prklxblirfZ8QXKKx3W
Fg0Bjznd+uj6gzTswUsw92M1hWdUWsBs6WdFrO7AhM4FILWxCy973OUYxeTjLZil
swkPw0G8vLqCKxCZHhnCN3CLK1mTHIj/+q3UkJJIHezHJUlmiFxXLga7hFPBXzWx
qNGu51I5SpKqlHtlbdDICd/S/2uo8bjOn2pKVEEmagCO9dD3AztXK2JQDp09Q5sz
RPWuv44uD7qQtbU5RqBqYhFYmA42xquyf7ognvs20D5e+UaIGe8H5EZvfHAWDGQ1
0YIocMtLnRmtNi1BycO3dDctf58WhS6IksqT2bhvwfy5Vs7oxDX2LxjqXPRNOcAm
sVJqoTPBjr/t188OJrCkWRtQVjulQheZrG4aEY2sQ8SaptuMVtvR4PaJh0EG7dhX
gU8jbUdVnGHiziKjQOr+mj8h2uR1zRK6BWHLE34lqLmJPiP+OslPj68PNDen3gMJ
UhWOOjiIQvwvMK0CBc+9xr7eC1G4dpGcrFrMNrEUI6TMQcm/39iTpBTEmrdPNIJ1
VRVYSB7eTJpRuA+OoxxjQBdgnnHiNiyKtqhzQozoWeWxnIHMEsJ3TZ3jhlyOuq3I
h9KVF14xB7TEZ83DhxXFbrQQGDX4NmngQxgAlhlikZbJgi8gpsFv+Kmen2ZZ6o+O
hbjsjPokMDhvk9bCE6dTvZvz4yppLGe8Je3VITr8ByWke5qHsIKjHni4yUmQtlM8
GkuZ0XKsq91SPROWgjGcs57pfZNwtMUxLm45wOiHGb7lEPCnr+3zeuB0UDjGq7o1
ZzvicynY4ljSJPwBvrCHHLqfHKEBhbNVWWrcuqatTcksjd3iMEArHS3wI4YU3fxn
IljZbEXnCzi4tCHvwqbGc+7sSkIz471E2dpsV+nZvzJzWNnVsSDGeK7+5q6Rb7sW
lKRkSnsM18ZBD9t3K/fEJOt5Cz3f3U2CevW2g7XHQmhNQ030WN/xNOAE+zne3Hxi
NskoBy8DTEwWg8Kz+QNgqpe6emvbsnK0neaCjbJlIrYjXlEO5/iHVCKetgjMdr28
W6SN+6iUXyHXe0+juW8Zj1volVLNGH/9wa9puWnhrxj0Je/rO8N0Or9mISBv8POM
R0n+rVahve3Bwu+SZIU3k8QzpDXNWcf1O0S+IE24nyFr/uZWy+KVCO5lfLFt78Fj
Hq08u/gc9+/d9cJ+s4X9nm0pDZC1zjY/6PvzPbhVwC/OVzbvKslzjBkRPPSdAhdL
9i1rUSI+jbfVhRQBtVPZIVwJetEYaWxiEDUGB/0mosjXcDk9s4asxvtf0IHd8oDr
9WCiJDXAx5YemF2tTPm8/zcmi0J/T0B62fFWhIds2Eo3Rs70cOyqEnoBlE+EV6bW
OKY+4/myF+z8sz6ag/wrH116IwjmkrH2jjMh/7DUQxfqCXxqbPp4oBHYsxwIjC5E
59HIErdXk6G3HsKyoJhWzZYwHXyn1ELT2WgE63PwT+r7evv0RNCcST8MesTsPbsE
88fAEGvqbPtMVLeT6T4o19ZMrQ1g41wrumGgQgrDtmfOQTDAnTAokpnU6CFulBEK
ZdPRITQ0Z9zQ9m/y2wCzqsvqkz84rKj1688V+G78/Ohhuos/q6Y6g35qLTe0/fRM
/yqQbbnbv1LR2JWkr0E+dYBZaBUkLP5qDTRlllpV/wgB2+7sBoXxKEn3c5UYJfbM
/rqeycl9PO+As6pFG8/GHtDfmk1+Y14r6TRNMbKtPtvi490cqKfn4gI1HZmsstIN
ujuhCaRvT6QWNtUd+urFPqnNAuCKf1anJrR/gTrvh8nWAFdP/BxY2iLIc/51VvBk
yfLpofTCWI1oklkW4qEr+llRQWZwltEeVp7qbs72bsfo5sUmGsH3RxGfuoluKmss
ZXYUK8EVSkROE09EtQ9nSBdTkaViRnNi2mIPbTrnL/v/F1ZIIG0fR4g9ilnu0hpi
/VKIcICA3w2oLUkdGnOJtWP6GV/ZzwYy56wZa7j7omN9+YDPb/34YGB5S9s7Dd9V
DTwPdBmoqAsJm6puZJFEmOKzY2qd4/P3pCcfjIdlbVYa5b4PKslnoev2IDuyXQbO
hGB+4Nrj8bpL4Wzw125L+UmH7cVuadkR9Hpj0V8G+/0cwQavTVyNW3uk5aBxkyOP
M6cZQ9DraNosZn43PrhVaguTW0Xb+7uRWQk2QKjFMSMDSca8iS9SpL1zuklJhajN
yhUt/zCTA8I485qr5h7v1yqRH0gbwsEL+fY5JrjW/xMahQlMSMCaUuO2RFy0qqTO
l+bBLzbf0C5evGPPjVaQqagV1SkJ0g2D0T9SvqV84HWl1/I2Z1URnGJgBD8L6s5Z
JYMCgnZ0/FR+gBlMB9fMg04l5jAfwsNfDRwzKEq+dJ61qrlcFQL3qdkE8zqxsz9u
VJHNkcFi/5lwC9XKDsFFdaBYdFusbDxD+2ojQ+KAS8U7OmuGlmk7ExuCWxP8ujz8
KqPgst1/aogooFNvY3Yv/5SlwDWMuBdwzzHcsjcVLAWfaNHn+bCXPuQDMZ5DjkcM
5/XZV5hW7Uxr9bm8UUe36OQ6kj4gtF0y4vb2xz/83/t0xr5EvHtUHMp5Srr7UtoI
eUZRkihrXoQfX3IXOL3ffZIHFt1jBfhxMQZfvdXW2d2jPWdHXR6HqsitKlIqML55
vQLoSZQH/dIt46jhQsRw8VDp+taq+nibHEfnOO8CyZKEkQq0V5tWSnZ7XUGL/YAG
KB04vQqq8e32mf/IpnXwYHTZZD0QrNbkQCprKeoLyk88f5oDfZ4UCQtMkSfqE2Rh
/5cwypTQQPfZh0v2TGvoqJyofoCSqVBhielgmvn5Ak7c6jQpp6UELE+dU+2L2bFT
C5Wq2MfhYFeUFe2pHiJFoio1ps7fHIJb/SVD+99mdlXHy1Gw/8jI2Aj25UGiiFSK
Z91+dhlRIEoFxgR1MWOtP8hg92PoURIU7NOChZNGIEMP40l59YpGGol/vbeGGkgs
IW5i+qoIUx0o1HRCd4K5fku3e4bYvRkjTC/O/StK1GITC4ikRcyWbHOxWR2ZHXla
lqH+UX4NvmZWhrVFxmdVonAGXbP3UBFBfRHWOZlIiAWEIb5B4TU8uU6Q3IB0R3TW
xFoWdLnk19Z9YIF0EVNsjpIboR6eb0RbncP4cLml2RNDn6aQqOT6Z7dU5pha3EBW
LbeCCIdxlvHKV7AeTxYlX3r9o1UqpgKEf4t6u+yzIBFfXNpLaGu+bIzQLKc95DAF
/OJQgzw4GeautOiovYxneXN27te2f8yTKjblifG4uhVY0PaE31MM972c3Oo4CI/G
LJ20Q/oKw1nlahDg3A4wau82VbTUq/JEBP4Go6Wvji3g5G9ySqdWGIgMJ8M4BWVS
je/8B8wcfm2klWauJXd5CJHGLLBgaGH9iZD7OaPv5dBRBbCdTKM8VGbZt9og6WFU
vBvGtT05c4irYma1t0nRwsFdBfawWkWYwN4ze5RWv1qlJ0iB1UJvR1pztt/5AxUt
St4yZBEUt7NiV4MXDWhC0sMfLaTnPHVaL+z0MZHPrc8WTxZuGLEq2wlH4nrgMm2G
vCorD/EvjCtdXWK/xUVrfdau/gHP8W+meCJeZ+iyITKH44IkmC42CSUZJyW6r40H
rBtt50JgVZF1gIOtes3dtQCLhlIwKfdmEIT3E2gWgMRNV9s5uKzpRBjsIxRVbRZ9
FFN491K51DM6Y/X8q0V3ODVteh4kVI4gD+TwwqEsM0NybsZgfD3pg84jkX03mrTs
1//CiZhMGd18lo0JeYPlBmltJzRDR3JEe8WN9/sZMthZcGoYPR+Mzf/o8qWgwLmn
tnibRNWIVPo2AeaTJk2KeunO/5cMH6HmORJLHGtEoADlQsMyekQ034YB4EAjim/Y
serZtAgSn1mhWgSVN9GL/EdGbvzj3zzUQ5lwtzCjaaqFwPEzhVOYxR2Mk25sGPTS
GrhcPoGg4YlCg4YD2hfE29V4tuRj2Oky3XL93ZlOaEDe6ma03WX0Il7Gs7050OqB
ruuQp+oXSk0O+povzFDzHu3Za9COKqAC8pazZ5ZY7iQXtEVPz82t/PfvLHr8llcw
R+Veho/I9xcKftCYg2T/pqwq1DhM4J0oCvLpDF8qWbXdB125AQX5jEXtqmGxe/r8
7pQg3UZ58OM+/veZZWngl/9dlRGKc6SUbj/1/0TkOrLlsYxclHjVogVHeUls+XZh
GgtABwlH7XvgBGMHQJ83oA==
`protect END_PROTECTED
