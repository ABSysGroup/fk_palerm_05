`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nls2GZknRiTx+25/KXBUABW8ZMJDIPix6DSBxJCS7I3K9iip1kHXxkbE/BJZQfdJ
EQwX6zZNnCipmpBYSaSCBp2KA4lI/MGV1uN96JVuV56PzIcPpFlZN+7kurdnT457
N5avuF0udV6pe/tMwlDTRaHXzFS39cZvrsLClBiL3nTnK9AQ9h7i3aEVfvF7IDI8
DUr1bY7spuGvxzvAPem6T29fmKzTUDI6hK9Pmn7/vQXyNjwTIb/Wf7wa82IW4Jeo
Et4NNF49Iqlz4GMWSZWsrpN1/u4c8SBWYHRJOg6tpN/g8s4DGwkD7fZ9JM0ovTYH
EqUG6tio8ctyjPGl/2Ope6/ltkHkFLO87lSvRQVsOi6RKQnVggxKExDikDEieksC
wz2W3mmTmJSzM9tgQljOX4PKgybEExZNU/W75e2csIb4jZjg1sCsaRw1fTMt4Rfv
Dn6tShiL883Ff3vunKDY4WC1RalFIEBKicRiOv4KbNFTQ0sA8uejOdmJJeqZMVhV
WiLz0WoHN2LeUEAQAZf+cZF88sUgU5WQaSw977MzMe6Zb7XixrOjtdK56FdlaGcL
+WrVCkZJNeY3L4pXvpEqjeJNP26dOQBtNJArDN9WNe9pg5U3JnyKs+BgKC0DIK+P
zjIVtA3KsrYVvcLtfsyYV3HWL5A/eU2s9vspWuFgO/ZsunQqygWdqinEIT4LKqzV
0Ex6uJkl4OUDMFrPKSi/bAl8N3klfg2xGqemt3XNqe5fkcMYQwC1vXmnXe+rIH8+
`protect END_PROTECTED
