`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ztu89jF1HLsKBuGJx2K17FF6qybG6/g8D/J1fa4RdEexILY7gO4IOHfsdZdg1qM
y6I+IKN+PlYQL9ChUAuJn4Acekf4i/b89HMXAw3WlQmHQtkYo+DFxETvVT8tfrYV
UNTIUK2Gpi0EJ19Hm+PaaUXlyVyIxT9Y/2ciGtwO4U+ptlbtOOyYkrXTLPlJVwg1
eNI5HyzAJoQ3m4GEa5GyUm/r6eAFRX93cEVexdX2A8iCMEE8xSdAF5LSZSTQ1fON
NRdXInNxyCH0EplzjUp96FLUNn96r9hvwO1IECfdV1+svxETpdjg18AvA/+IwWxS
H9UAF07ECRMtB6ATxeprbNuKYtZM9UyAb9A/+QZuxBSGVR5cxt1ou3Io5vaAhBra
tdl77ugohfLHd0djtNIetHIvTzBcHxwYuJtOFk5NOC7fIMhUWhEZm7P2Q0Cvn+j3
FiO3K/2Wf8bs6hnksrnUmMqYES0sPcNXnzr0zkHrYJrdxAQIs2P9eIy+lQ02cU+O
JA8oiYG+NIBsThplr0CvVDn1TUKpUy/4F9Be3TvSjWjaNWKCIKLjZLLpIG5TU0zD
IWx+UBg1IGLnjmLrmzntemvwT+kuvVwyPdSwsROJloJ6IMxK+LcaBDtrDuuVxtnM
V9mLiE8SPVkBYIf2bTalEcycWhOzjtAs/0V34p1pBoIsDIYhnXdfiJbsBWi7XHff
AcO19yOJUK92ZEQkiJjkpp2Jzu6heGldcKLfH2IyxvJP6mDXqzTkUZKX5IK0Lbld
`protect END_PROTECTED
