`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZhCZ5h199q386TxpDbQuW8eEn8d8fLWPfFppCt58YVW5mkh8Pp5dNFa1Sa5Zif8Z
+siQmZPXCGkmgZD4y3oyZxiMSRZ9r74CYZib+bHLPwZ159ls5L9vtjtSQLZU0cDw
8DRYfF/8UnYO6P+lOBIzJgrixbF0qPHKGz2tBjaDmmg3C6A7CNL50rDRa7wByN/L
aJkPb/HzkaVoKSy9QcAleaetmrW0RwRN+4kfbJY2/sDySWDzji+XUltyBHzhnnzb
p43ICQhzKvmdc9KsMRxAAd3pc+1l2l/6KWvwgvVuoU82YnBzc7zYfTPlwh6aG8sd
ylr6cUGpXbLTMnwqR5u0B9KjTwZijphuF6Z78FL+p74g5pt7yYjJwqDECCE12Bb9
A0KWH8gPjdwfOViBeIbKnmtTdOczsBCyYVs/Vd2HIT9o9dZyxBxTmdHswUE2y8Fu
xpO0MpAJ/Cgbc+isxjaWvvw8TNAykq8zM+mAg2miC/O9eOhZmwBveIILpJOiWuNK
k6J6tdAcVsCvavkYnvuE4jx196JVnT5sB2yxpqcnkSIjkj+3/GQxIxUfQdlSBs8W
6KpsuLpVw8suauz/2ypJSbRdeiHdaGHBLeV0ovRtTqIjTKmFt1rKl8zuD120s9hz
i83pj94YIxHwmx17+hb4xw==
`protect END_PROTECTED
