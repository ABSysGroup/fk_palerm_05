`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WnxN/SaG7KBBRDRPsxoL9DC6vOoaa4l2xg6IYyNbsMz3DDPEPzYwc2koM8w6toPc
jvoqe25IML3q4mtrw22Fq5CVp4Ynn638bunpqx1H4ev79cvGpkkobclgH3hthHF4
Fi4s/E/0tbKBb5U5KKnBwfWAp3oub7C0ZD+MjT60oZZrbItYz0UQxFNqHeuQeudc
0+iPO5rMWjAJOzrRLjjwnqAsOEeSuueMVMEhSM5HEmjQa/16uNStDaQEXBIJ+Gue
v54P+XRQeBY6jzpc5HOqujaGojl4ZTMpW3Tb+mV2gn4=
`protect END_PROTECTED
