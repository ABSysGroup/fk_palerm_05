`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5MQ5987ZP9sKf1TgL2o5RNDYh/04yQOjFBcm2UYa1y+wN+x7r1WUUcCsAb5nW9y6
IHlIvZ7o2sgtSSFpmLIz5oSoRkKvWT/59iXExIZvR1qM53VVMBs35Mrf+C39KWEc
l3QjN/wMGic4WDh+zp7a6xFgfvcLDFZLKz8JkyjSvi3w37NURY7Iya4iHrGWuS9k
pkdN0Bf2EfFpgsCeK9Tr8Mjl6y8Ojaj4byQZ9YA2YFz/q6eetcOTS/L0dNjrznoB
lz3v3y0MD5qPxxFX3wpAfQ9pQDO+X9w0xuomU6qF/t+Fup7j7VINRbpbfP+o8Hf4
seN8nK2+ElUDEmjkQ29478EANJCZA5Tg/XI9cY+lPx4qYFxSFXl0zXnA9eLOPkKt
lBRVFsDbluF1gb9ap7/qryqwtmjsa7szZwJY1IG7bAoDJIfc+3NMDbbk7v5p/q5V
LmQouCvj9vBpHHXNBxtldk2boSaTERanymM40S73z0HYYebqWfic2yUzE1nOrmna
N8MfIO6eWUKjXoMF8nZbY0eoNKPZuNwdIwdaBkO5iH4u70I+vIb5Puc39R0Z4yfR
mWuyQh6tzfYdF9Naafg4biIgD25FgYC0+pdAbKLdAfeZ2tuS8ZII4RZblcMN/Sct
19ifDfd/AWBb15OY1jCZjd+2fSny85i1MBR05LFqbWi6iEITQTbIR6iXT4bRkzS7
a0aj8HAxGRqw7e79llDwzIfXE2zbZCOw+w3Wv04+Z4cRaCZjqKo6cx5vbLlLBdoK
FFWMt3YX/9bUlzLQ+si5b/y/IcgHYutShn8pAQ3H5SJp1HRTIBzSomFn0dCeaDZS
5D6kDJYBTRzlpP9/tBoox5m0ATAE8LI3SZ6kttbtgbER1eU14l/PQhywIzvfvsoa
YmWBG7BgofPEbMM2aPVWz4QM88F48ImSNb6mOzovvgGCBb3cHlP4M2SJNhYnAqO7
O0FFQCtqCgCCJWlgKqKNbjBCDr1D8JNtRZ2w/hFf4qGy5sLbFJJ3oqd/TNM0uZeq
`protect END_PROTECTED
