`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pLlZFgu8SgTrHiE8x2mdC2VviR5O9N03fGf9yay1/YnjAhgEXt82FxGHNpJAeOkZ
MzoSqbQGTetMmAUX47Fah3rG2UZEAtSYTRdpJEkGNkLn1jaRsQ81wLvLYfHy6HVJ
36EdWlKjzEg/G8XmyVyZO4gQU8Ap+a+gAtFHLxLL2os6f57ByK0xgZY/4aV6OkEC
zgvFfA+enETDTRVj2MYrA9wbPpyTUymoQTTbXuPKFNZjWA45XPyZtmrdPsclVLmI
kxM5znU3fivSe55zYNHgs85+Jx7D22jGcgLyjCJmg8YkNfxJ4vfq5rApDnX6ZZbA
AmcSqySHVIA26TkME3kAjsirf2+haahtY4tzfJQKt0Idf7IU/eqzelQ0CVNCbWDJ
kRUMRhIic/H6XBCiJtMGZ2e4Z8SWi9sv+ihEvdpjIbxLK/V/xCUEMD+emWlNVB7Z
kFOBj7OoTKFFxf05nPbU8uNF8Bo3+hcADcIXrnrcIaY+gYaivnrgGLIrizxB/3gd
QjTGmO+Kby0iMx5wWkQ0GZ8Lvv8arldOmplsP5ZIpmrgmuCtlPGah2c+ba5/4CgR
AAjBRrqktvi60LZ1y5spUpWMlQ/+sJPe0MKlnfNqWA0lR+ZEghx6KcRo0gHT/09c
UaF+HX4YLLSl7PvAjQPUNg==
`protect END_PROTECTED
