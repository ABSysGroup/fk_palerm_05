`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zX5KG9qUDhjnn/KSLuyccsZDbHzUfJ2KGz40yTHhqk5MWPxHQwuxBmbfYEsanP2K
feBTxkrk5sy5UUFcdHsxkhTPLz+NvhcmMgI7I2hCYDnc+BgtErsDDbITw1TtmDWt
pMtuK14TukzboWTunGnnzOJ6dGp3ERDTGF1Gqff0Gjvdytqu3xa8wvMWes7dBc+b
0XcU3x/Al/RaaX4oszOoGtVukJKHWoV6GjMOsxdO6kyRSvp9F+CKzLRKPIbqsqhW
T/tLaO8nCJH1kgOREVBppj0jJd+9A3q5/5/Nl2xYN7uTdGs3Cv0oflqQExVoyf06
3ohM2figN3u9tmX4zCbsS/KrONeRW2kXfsBic7zzTDZZTL3IL2tthUUrAZR+bNbd
hk20GSr/PqJ6KHq4WiqGSdRZYVWdRXDJDUy8qEwT2+hpnhIsvVSeh0LET5uUHGaz
dySxIU3IR1HwZ9b2d/6HLZsCDikuPEAilPtI6sw/KYvVDweBdEa3ceBTrVOxAOj1
my8f/mFnljFqbB96Lg6lHc6Jkyh+HRP4RLmG9IPwkNVV5N+DBGjePZr+OaxTWASn
HQXz9fzLGcsSp20iJh7FkB/TFsCXzygVl+7dInt3W0WIwgotfow8vvzxYOA32iOJ
Uapxoa1eeZhHXIWpdKRYlM/6e4/RHR+B4WhKDJvrbsyd5qOfwBfdMDZsXHqk67wm
rEYYHdaDdWv06a1IFbRWi1+uta+Z2FDyZXZEm1T9YuRBwFefo1gNxwzZbMrK6pNK
h7wMabzS24ZzR8kmVsVWVkligz2W9KK7YVTaDAyGfOXJ3dvC++ruAXGin1KbJkUM
pqDTF2c8lVxQKO4Krm3CCTzfyEVBJ1V2XqGVT8eVtlJ0U+8vYEAGjZ6UaDcDmDKb
81CfCRYlnuyoJrYkvsHfXoR/kBaAHNCB4ytw+AkYXhQ5QLzGRDvBIuat9fVWiIjy
srwvw9/uOb8Np9fe6P/CVXkyzZG1bG7Q+P0r6iegIZRfdidQk40RsBJGw8hssMTF
1stHAYn2S4qBGKaWJDDubMXZ9tnIn+lgep5sXUmXCctzGkoodWBissqPGekwpDXd
4eys0nhCXG0VMTd0QDeXjwEwU9tVpyJVXlF3iBKTOWMb6eyQN8aHNlW4aIVqPyQL
3NJ26uxkPvcYFLeCsBv3cBxGrDvA5YNJEltc649ByhoIdQMN9iPLLMujNI8j2Dsj
8Qn1iab1IAARgM5lYf0sk79xmQnYQPVE0mbzibu0fB9LfmNUHlXGH4MQklSPAZQF
mCtGZKNEC1wm2KQp7kTG8ofbRhM3M/oD0I/1p+J4nyXXfW8BojxaFtxy3wq9l+/X
EhP4CKttIJSXKiCOoTPgA9r83sZMfGAR+VP6BtHUuDQnBv9bn10iofUqJmeq2EoG
5Q4p4u8gqpezRBaqLMzl9xArF7jNvastKnu05fj8W+NTnVbyorpIvtQn63x+gj24
vOBHvP2JCNKIkuyifHcI9zRH+umusZPdPj7Q27uhCBBiQWCCOxZC1S1WRM5N+oOX
DRsOpwW2NV5J67Dt1/Y9DPQpglS5+rKrvicz/Ybb5wXTL5UJRDMTUD1YvDhQfEPI
BDnEtjgLiSshLwXD0N6Qh7hmhNdrmnXnoVwCbpuolaz/kJn1KpR9QuOc3carcpCp
gqJGp1HgY9LMRAC05ieaTCjDSufng45dVwREhcWyR7iJooeeQtH8FyiRHO81VC9S
KAuuBYB5yBqwKN7ojHh62+BCzpLozct0gF0YAcvw73y6KiM+dWDKms7hrpdgwnrj
o/Mz1YLuvr8zjqED4y8KF9D+PglgCoxlV9968ZaC+AxJTrPSfDf2cNWwnwMl1I26
lHyUMddG9DgOqlV2ZD2IycV8HrUEq2IX6Qb4EHeCJp9w2gTPwoFAUnCIYFFuJshH
QfCkpP/DONmuHiWblAV3dHB1vbC9AGa0+aMfVJV0YOoeyRBraq6c99+CH0gOuHxl
8cn/ugDnFw7BzQm7jc7JPqAnjmzjYd5QjJVplYH29Z74OQJbOIS21s9n4q8NJb5u
ySBDlKq22tcGftqSRho7tBvMlFUg5HPonP79QwGA8XhpXZ/V0pMTdGRYaf+4xLqV
YGYaqab9lu0wYvo56SCu9STaDbF9ZeLqTtiZlZ4drgBCpybbgv98jrnLlrCGKNaK
u6jJBRAOTBqLVzHbPAJGGStIIFT6FOT3fay46mAOHAQFqdz25v3cXvafs9/PDC03
ueA0hTHgvEqOwZU5qgnk5VN8X8zwm6Q/jyTcrQ5zdGssMyedpRdVfSuZw0lrtTjG
gllCduWWCpuMa5e3H5DFp5lvUrmWk+6IJyfpYoOwc3cgeHyw1EOh8d1WegmYCEk7
VvvqvYuRHmqO1GKq9gtyNeo1JM4BZP9BDz+u+xMZVaF3pSzyOEMh5waZTg9/+32/
H9LDeBUGR4paih30kSnIZqlALUuajR09y+j64piRCZWPwOuPwogjg6iJ00/rffMg
Z5y7K3OErzmkedd1J8wxJjiojMVEJ/CwdMxXtCMWOZO+gbv5oYNDadcdGV8X3pOe
aqE0A2UhAqI63uzoVSU1YRnuTTnQO5SJdGwkzGjOtBqthjBnAMSC4Sy5OSJW8SGv
WfyrxQK6Vml17fBj26B93kmBGZbC89fkj7H79B69yluzuThKc8tpa1GyqpfF0WTD
IujWhaqzi/sfB9Yk9PaPCpJKqMWoEB5odeNfuMz03QL/evIPDN9ypt7M6+FCrkX+
yjfOJ9pSWABEtxhJ3/EWTvSXzq+Chn3nNhWY8AyJkEYBhIKn3SlSBgngipbzUnDw
GMQ/1W0SZ7gWZMUzRyDaalkcu0HzFkKx413LdQgFUJyZpwlaw61IrAGylPx5iGTa
wC9iKcQXkPXkkhO0F75Lp8wm1I5h9FuoCmW4LFnDml7Nsx54NFmMCB3LHP3Stkm9
j22sXRyX+x/F4mqyo5dcTpWwNBZ6b9Ur3ZktvGw/xKcIFL/iJUa/2rl6BgU7Tnyh
84CfOQU8ZPNMjmxc7pXGxglfswtecewtqtQpLzvKpivC9pIdNXlBrvW/v1Ynmi16
Q1mkeiAtWrmYF8dDSF+PxeZGVZXhY8Y9gInXtN8rIKAkhhksXgSTrr6fNPjznwr7
aG2SyKlcwAbz39y/tt827H5D0JxzPG3Zq71AkFOWcih/djWRuvbWnPh6qQ/sDRYm
0wIJNluwfzYGmlRmiQEmTI4KtKGje0pGWzcWKvLoRlnTww6z47EomrjD0ar9hypU
DHs0vTlowtS9n4eKuVCJEtyR2VGu1iZSqPFh+SE7Uorc9DDlDZ8PABdqhy8EmiaK
p+LzxrIuI4/+XAk3ut09SK810tw8DoJEEzlgQqZ1pTr+F7sEZ361DhZ/Nnhrx09f
mLU8jUSAHjNTNwHOLFXq68G6gM/IFEQ4qMuPlOBl8DtfH/+ueLjrLHsHpLISLNys
Cv+avIhFmvvV1Y/puxNpfAB4w8R1JFW3BvEEKos1TaXI9xR11m/oSEoC9YZa/MEg
Xwk/mTGeVHeM3FZwdJYCNwqk5aPMqV1IsU+U0R0gIl6r8NHPdXGoL6ZUxKJGEZgQ
1Sag06poS3/5u2Lv+f2IgA==
`protect END_PROTECTED
