`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wcb67BHAXwNR459zu8GhySp68RLh1PmVBZE13I5naO/Zaiqn1Odpie/wRL9tUOjh
VLJ+7X8QlV3//5e3j/Uzj0P3WLtAF3ICYCGeT8gGi4Eaf4S4JZdU6xz2yoTybV+r
zZE5rq4ZPIY4tN4rDdVsOF4/Tf3w2hG1fhC8CaRtV2PZTRvnagQX5HH3fvKuPcR6
NNcTo5fXjPaw9Hn/kW04/u+qokMUxM0dN+yQdQkZ1VwoMWXu4n/tpnU+zpWy/7pf
BiU9R6BnSKDi5582+B443CFwe4YCugMS7jR2qaqzHLBGHM06gh3e9tegTm4mn7X7
NliSIzkZjP4RM+UVoZhCL7Sy66nyGfHVt9XlQzzXs2v4qABpnEOq8Pd5r9ulKL/Q
mq1WDn4m0F2vQArDV1PdagBn+3yYWlVr60N/lTYomeQBokb0eO85HcASECHznPic
7EjQ7ctooHtGDYNdR9H28T8MjNx/GKZ+qX47JcCNqIFHI/Ep+IkAS5hhubXGJJ3D
FaGqehLiTIHACnj+80gyDquBq2iyRxq7NqfJCYSwH1oBnkVIS5X2SusoAUywTaOQ
Uk5rbaAZ/M70dMv1nQYQ4/UwYQbamKrF4fQ5jnwa4gm5BRKIng7qsEGEnKulIFDt
6cvNqR++ff0CmAnvWryfHaMOxZn8pNhfNfFp1IeoaoyM9l7wWyyniNeN46RIuM7C
WKY0MrzuPo4t6LAnFg9aV04IYiOmTLb33KdJJLRG5uYP+Y63iCFdEy25yGo/CtCv
bOEwVENH2TNiZtF4OnS7OA==
`protect END_PROTECTED
