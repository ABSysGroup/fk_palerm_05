`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VZR2VWUAOwcwnTYrUcLkWzQKveRFnAojeFrKp5qN/fJPMZJ6kzTdrRMLSr5XScpF
A3B6UO+dSEDkOYoT4qcgjp9ISY8qHrWSDsugfF76lNh+ireDESQMYqppIW9f0PAz
6gfMopyW7qvKTMX94ZRvpFCAVJ5HljyN7LCsgb/MpT5Jopp749tmcs3PvoG1Ru/5
YbFnPukF7Lox5DKgSdknfODowKSSWAMkk3a8n1sZVJa1PPruB7bHpszKx441hr5e
LYlf4tTOy1FqWBjE/IchBPRbUx7ZLPmpVtx4j/pAlSMxisoC9eKk1sTQpin2cA/7
dpsWLESBu8pELyhDtxiLVt0YH7Gn6mfR0nIBrhrdDAhVZHFuH6fZ4mpFlAoPV9mx
sHYLxV8xeFT9W+I1doPNceEenZUQwHD9hHYjgeAxTLGJSVxhfgHfWW7PhcwL60Sk
ZgjL3KHLlefiJy4BNAIYHUHzfBbaXR4jyRZ/8sEk2XpBPn6lEmANLUIIur71fQT7
p4y5gH8DtxkXMInOvQsnVKYBIZGp2QP4yBive2V75io4Wnd0zOINslAbgY9jHLsj
1z84PcAyPeuJb7DDyi+cIrK7ItRlsENhqTc3b5rz4ViIm+wD7YfyUpYG7MhqwNcl
PCjoT34ohv1wCz7awMtLvSg7zVgr2mQ82xNICesAnxoAFnYRsDAKpvt8ua9T3G38
q79rwRfVKbp++6ZbPPLtFraM7EyCOS90vAbWwdVeXxUV9kHeGMumNWrQ0Jvsk90o
X46CxYv5brCq/bHHWctJzM+R5pbO5mTWSQ+EZbKWmUOWtrsMfCO+DI9kF0ftTd9S
h53AHwqnzk5sHHQGaC0I3ZDO0ZqV8l2odZFk7dXjOzCSQa464p61D4gxblfO6hkm
bTOLeWxJgCR2+pKHvJJVfvGANUuOFqQMwiAJ9W6cAIu5rNpqT8/KSCPXLay2AvEZ
OAfH1Eya2pZQZFM0MFrAvT3W9wWXIoIcYygX6CC+J3WIL8RN+Z+Y0U14gdmcgZp5
mANlsdnz9D3byIrqcbVXsHHhDFw+1sSUMa+ZhJGtb+ViQp1MEILrps9lebuHPI/i
mXe0yjVoGDWrd5vZFFKjSg26xSdMPUMGiTqzqHm0j5qUjuyx13WFnj1ronOuoReQ
Kjhc3QKYIxL9QjwdtVvKSPMQG9g4BDdsB8GJ4r6hPBB66HAPJmbAEMDuxbZAUk5D
PGV5+u51NAH9iT6YABRA9MhWbBZ0SY1fQ3+1S2LbLLVmmLLWwCKaZIuLUVH5bhKa
yQSA3Dqiu613auDw+l70QmOl4+6rMkWlX8mJNMoGz7BO1txPIDwH7xNm4HJTM2G9
jzKuGY2KpbaE0bN7a1ljugVhSFq0kKIKCY9R10nljvDMZQ105Umv6c3PRwRyvYGJ
EcDiyru9u80MCLNFT2Txc7zwVxKonH7bI54L+6wde3+WRyj+GI2AyOb3Hb5bsROk
n4KIoz8vg7R+KNTRU1OpUqPLr6G9SXGF1vsw2WRjExof8fkJ0Kc03R8zr/D/1tx4
`protect END_PROTECTED
