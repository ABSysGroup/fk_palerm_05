`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WqTAZ3t8HRi2wsvxuwpFAceqSjuU2sFkrLEXfWtuOmLNOTG4sT9DmYFXJPqVwPuV
j1A5U7a6cYoe0GcTLqWKl6fEWzRcDJeOUGgBicqnrPO3i98mCXnFzFoUXQMarXEa
XihvewhTdLeNA65mroVuOo0H8QR6wlNiseI2WUBWmH5SuFxbjOwNBvP7zWFURfJc
ZPS+WY/FuB4owaUE04iXCsAs5vulcvLwN/qcNPfV8vkEbDBCpOktGlgyZB7qOmN6
z6dm1WtLDmE7PF8Q9T/9xajb+RpYrfIChQqBR594w9VVg9Idt1cEm+ZuBpIo6wud
34Xfrf/IMCsmykW5pc/omRLhJKtdphYWafT5ktoMdrxo20njyakn7XioAYR48z4K
aR3X0aPH4wJF76pydtsqURBf1GQulbUUvw7MbmuonqtIj/j4xHNiwFzo798licdr
zxIYXYzJu/kwygMmg0KEDaK4JRYtRbsDvlPfJWrxFLp5XkSH/Tc499GdcNMnFSoW
`protect END_PROTECTED
