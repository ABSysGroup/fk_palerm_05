`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2PGKnpPtgwO7kdHKtZO5jMEy4cwkgUl43mKcaLXza2I8Qx65xwqbZGWTut9frikc
sm3ustj+GgM7cqXUgMdObtPmMCaMEXerRvq+FrmZVpt5m4mzVQwSRabt9b8cjEns
4q5WeBTXJUlRCO+doHZTk4KvGjHvC254EqcUoYloxUuJRDxFQ6SVFD1ydXoBuWL+
e9T2pZquwG1QhMd+wdVaWwLJCJm2hy5kIevTWImXpoqGLPC7Pol+OTdzktFu1RLl
IJ/uoVfbdiH4lgMEcodew1y3ZL5bmUa2J7Fppgb4TSCJqEbO2z9oD3DgUMtx3nTY
5SQryFaPlFcpa8knzSx64U9vmUckH/OV1KYeMLZuhNDnznt3a35b000ctiODNnYE
a44uaXEiqvhlULBA6tU2aBkEV/rYLlVu6YbiID9CXDbUU0eeF7hZplfVlh7P9TL+
vwxLgRULHMT3fEWsfG/BhJp33mCdWHS+y/uxyJ2NetLmzqlu52xwcUlvxfjT/FSW
mzudbz2i3dE7RnHLwiFXwSoRywAQhZPq+V2drT30E2TN+FExgq+B11EPKLIYnYf+
u6qc9rNP+jyTNeEVWhjqF7hGIu4nskBQ3bP0C77yXGWhuRy/WhxZWwJSsm2j8Mhf
Ed9y4OK74F3WNGYBKOo0R72oFsMlB4KUZl/4mKZ0rl74p91RbYdeP/q7G5V2aTrl
sCZwo0auSNMpfjxAVEG0UA==
`protect END_PROTECTED
