`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rLIPiV6lRgna98c3yb9gc5Xr6Xy2HqEz8ajLj8BSpY/Z1QOEWjKNZPfIeA8DLm1D
Xf8yQUZUtOU4Dp09Eu+Cx6PHJODbMCtYE339ty28zAzG6fNjXvkanfc+QkIaDKao
IJewvODQxqi+OpxJ9aGKiDA7kaaCpPJoO+Wz2lzbmVqCvomk7PNp049FoN8HuUnU
YIzpGFe7MUgndzkR3HCniixApvuUBiTE8fQs9rmlpUBo/d99/IxZkwlgHJoEKpsY
KeQzOIWJKn/rvjj2+7QeDRYyH9+gE0iICpV1Q0Fogj0snOs8Vnb/OkPNMZqWzWF8
bgCTSw6ld/yuv9LaAxdHgw==
`protect END_PROTECTED
