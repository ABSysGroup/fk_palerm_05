`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ffwnDAFWQ2qQg9ncVDlA4S/GjazSjA5TyLKUrxcpA/xiTPhksRAt2LI9Hxbbh7Zb
A5KI1Zc3jHxQ1ze+22HOGs2tIDw1ZOVO1Da+n1kF5UUNPlqBXl0zWZt8wGUb77gS
ohP/b1w6D6/tPfjC+umeDTg2n6h9RVLEFqvoR+wJSsPnvLH3jSVTXBMxQ+PvyJKm
MXwVilt/nvhvDbBoMy8AySsQFAKlgxStUrzvAPErXrdT5ZDNygPm1G859yciL7VT
LH3lXMerhe5PrhYytQElgLc/ddZuXYXegHQYohKLL6S/yNdm4JdYG0k6CeZle8Ef
jgHk/q/SbjO1773wJAMxxC4UZwElGfp7kClmyUfdEZHo+JG1Q0W0iDN2k/LyTmgE
E+jyZIX4oOFOjNNexrvDOVymTeuEZyOrX8D3n/UNt7bk+vi598O1YeY7Dp+lJ2vo
`protect END_PROTECTED
