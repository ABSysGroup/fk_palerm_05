`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
irFDCsoaVnFChoc8qZ12Ycva0/MUFUlP5tA7VZ6iIsoXOzzOCvpyOHihokOaTEes
A2n484EJBiFR4TfSRLsMTNIy7cW/3GfHVlwyUslCcZej3KqMlkHFLlCiggBdHUNC
eLxamGnW9prV9NsVC7LgOLCEnd3etTAxRo+SmkAZsWeN6VE4GB2obHkdUDLTmCgY
y+1z9njTZy4sIaN/6P1/mOapTTVQqSX5pHylBYXMBQcxkXG7djNNV0zdTP+DEYpu
7jAyN4dIwp3EjT9aCwls0htpIAYAiSUGcsVnUEEjlro03W6nZkSC+0mT92SWQSdd
pKVmuucG16398pHYNja5WCPZzGlgGDz3S0XOWfA+uYuO/j9iZNHah3fLbp6zY3t/
xV3JmmO9/3HjYD734v/joTLRb6KILFZvGQCTXpnod+OuLzqKx3YKtdmqpSaa6GPL
7DkZF+YoCbREF9oo2SGh8sILfl39F9kbQdZYDTDSNHpk0QQhCg5PmDQGixLhyaki
z9OveL5rYRjz9g4Hy6hrduN//HF8iBAStVRa8cw5V5lPrjYvtEuUuHDeiqo+CsIM
LJPnKu74tSqPniuugkiodqAvw55rFN2bYgoQYbcPYNoYJKrdRs/KRFsPElPOAlTE
P3OrzdZMERvZ10QmyOWcCA==
`protect END_PROTECTED
