`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aMGzzKWOmbC2v2GOmX5oryoYb2UkCVYQ550Sh1SSciuKBOpHXWJfszn/6fF9HVeB
H6aVROen7j5oxAjfBhG/T3DBjnxZ7y536eSv9M1YKAqsd5lvoWDMGMQbyVPxI82J
YfqxH7zFf3OnH2a8wrhV4Jsbb9EdBGtwSrYA6BXaaMashnF8WfqUOAatK+S09HW0
4D9ZYYlW1cenUdZMmvV+1AFxW1agHKcRO/ebjXPvyiYGuantbBbBvyAdBPnNqzlw
D5Q6E/e90BOFJY6Gxh2tLUmh1vwmPgpIDDHPlwEQ3QuhBuG6af4XI00lQqaWW6pW
ikr2/iWMJUY3dSvMGeD23afiMzVVziR67tJDanrMb3AQCeHtEjtJwBUzD439I00d
AyTAgonbNvDQyQ0zFVP5+yuc+IpSOY3gckkIG9fQVlNHJTZlUogwDsnyWW10VN21
6hgSdCdGDaET/BpxbtZjCScY3iwzKJeTyfhV8bz01FDHhczgRSKKModJck73VxJE
im210dC82Pb3Gu4JWHRj8spcvRi4S8yQS7Q2rl3fw9HLaa08qmPMNl8me0RcopQq
5Uusk52fForWcVWY1mYc6hJDE1ElGaL6KfHopzlpJ+Y=
`protect END_PROTECTED
