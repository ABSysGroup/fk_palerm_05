`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T5LXsukj+IqxppZM+gknoFclI1ewy50DSPAlrGAI9cCOoPLRDvjRayZxyi2f7WOw
dj7X698Y6vq1Vjq5O4TrQWOxsZ6uTGJSbiZYRAWzetMbX7WSl2RJACFWnIOR5ib6
xIiMSnyUWKJJb6gW9w1yufFJchu8uUGnBur/VQqIGBdKZbClCbH2TZ7TYqe5/hfT
TBobwRntcM8iLJs4tyF0tYnUOOz6RJsDExwlIQ9GfeOsgGLI/644UOsQVfyd2Sdq
`protect END_PROTECTED
