`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8rnWGH6/6sNzHsD9siAn+GRFG8VPSELTdBwwqTf28BT2lClk+NU1N1hdqUK0NG2Z
Y40BpmAjoYNwT4aH02Yd+Bgn2faHI8adXHu3z8q0QUph7XIhOsjORw6ivNx5mhoB
jgt1sQ0sCO1xJ53vUJh/fPDJ4zP1b8Ih9rzf6Jb19RUHQndraLd5neBQAn0ZaHmE
GrKvrSTJcL5jIrr8pHt5Gp1Lyki0W2srvYzOulj78fLiHoEeJykONP5aO5f3tPGV
1Ptjx/ryCfOnf0TvBuppOPoRGbRACs9OMAAidYdpM8LSfx9LpqZObVv1rDc1P7SH
7a74PCV+F9QhwtYGuXwVB/1GQWP0YYBwtUyhuEY4lVBQz9sroDKjAL+J9Pzxiv6/
rN1z4yMAfTE5dcV0yL3WLKM20kq+52wRySda8ciX/iDILdM6JUpDECr5kwZ+P+tX
5yqpte98lnoUq26K8CZZVGoKy714sniwawdepH517hb5ZxVgWzWDsuaag/rO0WVh
`protect END_PROTECTED
