`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ggHcwIiNVm7NVy57BYORfKOs+nv74SHWjUXQ0a0dQg8dtU6u2FSWIvP7ke9uWRs1
Ic0aSzylrJ/jM5bbb3icE0D7uXeb2DxyGV0k27jD3zEMijafFB1xtUgANZMx4zYu
34Aoxjp/wLybXtpAjTnBezgF7CdbjzNhPEH5h3mAyhkVKeVJYbt0Fh2FwBS0A+/B
Y7qWNebnlwd9Z1xhsap7iYZVUTJ5A7VgV8MwMXauKyE8WwjzDy5pjnNpwBe8yH9F
0+Rl2FCQUOtcu7kFhxdCVw==
`protect END_PROTECTED
