`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Amuahh65gua7y4QPqWQhs7G8SaaMOYQTJ2kjOcC9+3VtHk6eTW1klaQBI0bZ/DA8
njGWC0aRtih6RJ2MyzNKE7pHHO9lZRTG9Aj6CrSOKWjb+7RJ4V5KCrWZw8+SUoQi
X+d41jutgVIbwG+ZrznkXVtDVKnh9+84f0+FtGM2/CyfHAdF0VGoCLreGDCnOXLG
D4QLdzAQj/D+yMBCrRfePYYuE1ltpWJibFAzVdDQcst0cZW84wwivbFix7IQCh5m
wmmAgdLxdnDL8x4u0fe4F9ocdvxuLkNpgegRQArWdvdfgZOHN8sCDETSJA6WsfB9
m/klfdGor4eFDXgJYOr6+pyHkumMlTc1xYY0rVJ+v0lopVcqRf2Ax3aDbs4/tNN7
Gc0oL0+aTef/XAg5cZLOClyuy79N8oponu3tHfu1L0RzG59/q5NOy1Z/qlSqSmJ6
utFT77DtfTlt85c2Tsm31WShPE9N31Mga2JVAhs5gPbktlIQrIBTrx5Tdimlc3a+
pCJYH3UfjEhwcNz0yD0YHiu5QkohXfAkbQNYHh9lY+Fz46TYdCvel/phzh5QRV8K
vuvYZaBrF6cB8roJ5/XSLwZXxU2wW7wAe9sNZuIahICrWqLEvj79FTb4IKmPiUta
SVSuJ9rmaAUO405XaY/rjYbUhqlFZDgfMT/bCPkylux3sE412aWBvWOokfseW3tp
ZuT0/nVdm3DiASXOzumI88BFDVoRUVbmgecKaAjZkh+qKrveIXk3LnszMEKln01M
r8JLwRhHlmd6vbRaFVRfaRvVtIPL0Oq4y+BkDOCZiEe6NPkDjiZ7nXLbzvJ1vIjl
yDrBI74kYgSS0fyyJKm0qF+pzL2hPnYjZYnnzt9EQdpn4WDSfdv7qfXR4BYdL4Ul
TiujrXTv85+goiAxIi+Ggv84VeLkh9GRtsftzRSloQ8YC5TCzTMuxQpb6MtExsDo
jrBsd9AG8Nu/qj6lNJgjSv9r/0tVLvSeY1ZDpaEZqfBJdHNFsIQSuiP1a1H9nvl7
aR0L9tim9zR/4gYHxBdOsnNTWfUX3ucpcQ0guZAxESbBOmue6Mb0b0Q3WsUibzE1
ouxAUhLxEqPk6UeXCtE1xMIC2GddQMMBTzkkVNvYJWoomxjm4w9DbOG0yrdv1Iex
OwwIm0zI9BdC4lwAzWwGU1X9gUR3DNUvawbElaiZe30upqcpkZCiEaYPFW/Ca/TA
lRb1odtAi7cMEvW13QEaJixc41q856tij6c/2s/WPlH52gU9Av3Dbpyd6+Gpojuj
ZjFG7mR/ty18i75m1RdQ/Qg25T2uAk36kTQcUOmScYd95zzTlJ5IgX25rMMgQQLV
93ZLX5El/q7PJh4/Ng7wb5IXAxjs9d1d2qU3uLRob8Ujp5mXiwumueh91RJetogd
P+LkRxZ9vbXUzFaVUQ9RAjFbJyHi5iV4wTk2I1NzQKXwi8DfiuRy7HPtdRJGYaOy
YzkDMQMGXYvzMCWiT22f2T+Q6gkG5RSMtphR1inff5JCNw6MQM3KNcpv8pWnbhfC
lJssU9JT0qMxnW46yM/HV0mY5Ys0vI31yqIClt4nMod4vgukR3+y9C25jKww/DFb
vaa6VX4ILvW8kBi0FFHeR1DXTxe+s3vhnyUl52UnRFho1lFbweFC0nhHCxl+gzb7
uznsaJRKrfIgtOjk/7d+TCl9eL6eGPpFkfD06GbSHWoT7M78MxoRq1u6cu6H6I3q
ghKUyO5ODO+Dv+e446zEYLV9cHbuBQ30tsQsUlfM9aEuGiJkF/eGl1sgijD9+79+
FXfJFqwKzpjHhK5pNoriqCsdMLGtv5pXey6ceAx9Yd/89R3HMgethJabwxPYZ5OD
FS3kAWJC4Ax81fagLZnO2Yz9VTXlR2V4Juc5PG+spB75aBrU4UnECLgkpEgKSKgl
WRQ/n+g6RuTHLvqGAFSt9XxiaLVux+bw8s3PAJRekIS2M5mMVdafyorEaQhIGTTe
iQB4Jict91bZuzAi92edcnviQkewQOoiOto7UnjnfUZLSBfZAlua1VuCsoIO4tLt
a04LstbOPEzqijG87zZ9gWPdxGtcXhVFXvOkfxiiQTrCfUJ8yREsLGxyzaETyPZH
NJs7n198FrnQr/fEsHQVeA8TtJWgu+z5oAnJuv9K2Rx6QM5MBI8g4z/oYMo6j6GX
EyxemmaBCkqwCiSBXtl+qPpR9hbifkaZDXClXW0m9ahE5hHGV2oPXWmjeMBajOoE
9QjAX+MIS5uhANCsev6aXYmDvYSavly5pj86wC03hGJxBVY5V5x+hjrlBZw2Ah8E
MCw3FI7tLwptkgcSyD25H4U1W9wjzp3sRtzTlHU4RNtC/wXd9wRHu3ctEtc96k6x
5LZ+EsA5SmReKA0p89ylCNvKGG/8zuk5cOhCo/rlho8FyldNPrQsy53mD73pbMOT
2sT1xSZkLtrPNVjb9e8BghJ36nmLi7Z0tSY6VBL78SIbdhynPzFnsYB3S6/louHE
v1T9GvjXlnml6a8GvCgrURW27G/X3cu/0vxuG7h8Sjx61dhK18eADBrZLFusbnyN
Bt/zolTXzOdTRNWXcNSoryV96BW2IbZ0bEzBoPkuBChSINU7rA3RTXPnS7Mo+YKU
xlxDkd/ACFrbBcv4UADoNWchnUDufIPl7jeG4QPIhl29bna2DEWe4yd+6HFv+646
tHnCazvFoaRk3jBr+tgjKZVuT0xkg7k+60ovhwrP4zWb2a4lF4VHgNIYpi4Sn0z/
mpzgzJ26TMCPe7pAhgk5wag1vjhY+WS9pJQusxMAzRODOm9/NHMqJ/Ezvj3rQSNX
yq+AE7p7wolGTk1K1ffz5B6aAgXyGndqM7JlNWwYiX4jlnistgAw4h8NeO2xaRd7
Q9/0FGhLmIK+3kJrbTwLVVn/8SO1CW5vrNuWgpPrbxz6eXjmQXU5VS+ArZ4VhPAS
tRBH4gaRdniKyduKCfK35FJ+do2NooKBMoXa80MhgI5O3NCHtn+dBxLbIAsfOboo
3RmGFQwneE9wCdeKyO8cmEAz1RLK/sTR0+utF4EUcpFYHLEvvI4iozqIRpN56bhd
sHZH1heDaTydtrXaa67nVV66+SjpfYt4yhqfaR+VZBJMFU+4Opw4FqBdXiHluzQV
6I4ohqnOfd6gEfCzfj+xmw5meHPbCr74ZUAJVR/+mxbCp99WIUYfK+NKieiwGbMd
8PaVXC1YJiPa21/AZJwWwXZXOs6QtQrJHC4mQsGLaom7td41ttF0EKMeYiDiMIi8
QzEqT/Bwn+Nk/d4upo++7lJR4gcUYqNPpfdx0d+g/p7reGs3S4g6ofZwY6SGROAq
MlvamPR/QJ8uXDqRRl4+PRGkGxh5LUQCrCW3jr/Vfsd5GgCgOwmdRmEnjd6h6OFV
yp4DoTa8+hwMpSugPn7nZ4iNChn3PhQ6qX+pORdQBCY1txqhVRVtNiunrewsdVIK
fpfxAhTsg9w1I/v3IGpO6p6FtQIzD8mQbmCAp/hxAdkkGqC3oTImFrdELSNFUbAB
kABxuo8Zj+pnp0KhQXJNanzcGqisXdPfTBclSmG6HBcj533V732BpkUTB3ktzy8x
tdcfrVCEdZMqBzg37x9IXarpSFGNB5IKxYSLzg3J0sDd9y5qtSO0cgRTu0FWzzfy
S90FXB3qHRzCi3v8MzWVzDvrD3dFMqYUBJV8p/jD5sug8woWN8j98VS4oj0+5KX7
uDkRM1MxzgRyFzULYPVuqb0HSX6g5Guoh0iuLEwf2SXCG7pz82aCQAiMbG0fdztU
iysJAyvtwCjWRDIFmtWXmM4H9Za3fgrZinnt7Cx61+YC/wpkm16yLI3QVWneeukz
0xYn0JJcRH4XZ8gAeMJTTphlevDq0Brb99LY9DnC7rOzRF1UqCbdfnLKAmF34lWl
ZcBDWpIj4oWHp7DPTnsMCNEQPj2CwNqakMz5ujdVuEBj4ATCG+JjX7XufZdXlPGv
f2xPm3LiFEfYWhRXKpNCscZNMUeRwUyG/9pw+mVluz7BzFZSrLn8kAzwMwpP0MPk
urHeYSUAu86Ua0kLzHf4MbFMtopD031THYvYb9x/91sDD9SS6nurCqWE+NR+bwy/
oEN9jprhUQdIGHINQTF3mDE03gzh0ebJ5EnaiVviovVUQx8jzOcFV1Y2QfmqKBQj
QBfzQMn/SDho/wRZGFx2znFewNxTWDvoGzRL2qTx7Z1UbiNaL30tJqw9zSQMe+lo
+sn+OgI8XnBKtMpygvzs4167la9UeEbQ8GlbAAuo5CnqCh/5X2Si5KfxOhqYFaq9
/AlsR+XMt+RY3gx+Rq5wZdaL+jDhDpf9O0XrSCaW0PZ02quNT24RLLAjrbkOokDU
ctmWuQIOfA8P7pni7u0NieJbS0YpKZu18er/ZtsyrWwNSbObb7IsJHJSKo+E56Nf
v7omoURVjn3zMskG8D8OSWWM6h59mrWQ2a2nXj/p3fiuqPPTMuZcc6CK3r21yGUT
fk0vST6u/PJ22NlClXUePwpFQ0M+xVZ48ldjiT09iNuTW41HW2MxUp9BmQL0skii
+inrkpruapPtdw9NytaInA==
`protect END_PROTECTED
