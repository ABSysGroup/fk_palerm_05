`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aYrWy6mGDlGDDqsPSjmAxXJsmc3XCM3fP6YA1V46kIox2eNaJ0gDy6IDG+r7AWV/
OlmBhcuUBjT9gIO4c3WhgreH4Ahw23WlAINeZ5IFGMNFRLj+xfIGcNA4RUu6buuE
JXBRDr7D4Z4xBVmH6DTwW+NW5o6+4PJDP0vyd07X9K+XBnTWJ7SAV3GByYp0RSdW
fKRD0quV49G7P4rl21LAtU2PNZYRonT0ABATMZESVFVuYbQOt8z7E9xFttF7hnNN
lA3WNKnLFzhULAW9JKC/HhE3Y5+ePNWG0PwJ/qDJCBAd3wRsOQwGJ9vZPXYmQ024
mX5m7R+ns0dajMU+Wm8tKjC3mMRvU3ck3AhktKxfZ57iunA/bA8B1NT6d/r/2CFy
K5JBhqHaDg80rNNj3HTtShwan8tKYd/VXoeLlc3jNo8SAcC0Bucmf0/wiFp0H2a+
pijhy04AzVcuzQT/Mb0oPgI1HxisRZfKDv8pNtnyEE667yTlUvdA9f5P6Jp1MeKK
887ZJLJCotrEb7x6oBj2UOYxwgDD/VjLbS0efwG4dUN9xHR6ZUdHfct9AD5yy0mN
o5wJniRzWTCMeStTnIZ6+zuR+CppFnJI2I4A021XeAU1KZVZLenc7L5mS9bPznf1
J+KZSuhgwGAOFaf3eeVnrcwnwmkoiMKr9Nn/48bf0sGSq3iRiE4zYidQh7ztRcWJ
H9IEWosKNMeTRCC5QlevLigE08e7l31UuEvuPwBATkBsBMfo3BwH52bDVxhgZkVQ
ukGOeSowxjNm/pdvUw6uhVYxZbNzUQ2vgpyTC6IDdRPtq5cPxY6QVMbhefdCj9v6
5gLt/QjoQ2updK3rDOZFg7UA2ge2ipRTUcSTEqjFqB/J1q5RGsKbRfdemeFFVNBp
pA/pCb7pvOPkYz8/xDjH0ghgUi9bD5chORdmreJcFa5WpI/TaVrVT1WmZg8vFlkz
dbhMV86aU5nr233kBT8AMuk4tA5tuww9vQ4J9rk4NfdG2rRSqUHHdyGepKKXTbr1
Iu9/Oiq/IqHZeiRjfU3sgQpNkQWGMEwcYvy3WiXqcuiDD1A4it3FcPF/blAPu4FR
EypYWjI4eUAaXkEiH7hZJdfnXIVNnH4RjK8941oV77aBdvgmsPXRcRknqTsXewjz
W9oomTeo8eYqJdl6jxjuYMEjD7ti2Nb5yQ0vIpvEi4qnTIqsG8nF+3DT8MXpkmJr
b38Li+5uAPWCQzjj/D6MyqKjTUP7QHsPyRsAhKrPNag10TkE2BJ7SL6wgcK7PPSM
1Du5d4ipX4sIz73QBFkcuLR8gg6SureXHcpUoBHWevT3y4bWeorfbUuAyR+xWSSp
q4NGAfGqMKWdNj819zjOTw==
`protect END_PROTECTED
