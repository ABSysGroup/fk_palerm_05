`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vHIk6nLwddm8wP4bbYouAks8yfkJW1hHI2kD+MZPjE8grNSDebwHWTqnIbf4Pcy4
qFCFCEkJN8yQtiPyc6/+O7z2aSSgHjcrvfqZ5yX9pJESmGyVUdJqg65+6bwcEx2k
cjHUuCnaZNmLrzAr/UFliUhgkyPRGT/++Apld2pD770ZhCrYWSrJX5+kJW8Xuq6M
8xaoG3s6ssXEizL0oqPuzkUGSTr91vwQlD7Gh+PiYeLKWBgJcsZMIB1nNmTWcf3r
UYELBTqph11Pg/Aj1VRmARra44iTEcZuKQTd7NN6WvWiweZq9noGQJ4eR7oaL6Ym
EG2hbZVXtXcvah28m1yorxPbDI0ZgOW8I7+Oi3EIpmojIj763GWgiLC07RYED2al
N0Ckl760cE6O4zrY3XxYtx5QY5M5GlDiEmRe22onGGnLgTVp0vUB2qbBUq14mLOM
ereSAV8DDsgCL9EOPlKk9qgotDfl03EXTZlJoyRx4F2Rfffv6q4hEmf8jBSLZMvG
xZHGP+z7pR+oqahlhWyDxX8usYBPKaZ1xJZlbCRg7uXAeCMHGEJo5SADGOck5tM8
GM21ZinN7R04J5JPF+2nRTZN5PJUpOSe4QAu+8kXfloT8SoGfOXlFRaZiPjvF+Si
mOdEObFh8MVGtNdPglFAVOGszFZU2X/JBlTsWJ6jNIyVw+6crzgv66/DFp7ndiyX
fp+NF3HOV650XvEPLjF58j6m9qQiYxWZnUESYUXK7d+xZ+6vXQvcqrVAhyK/6TNP
UyBXN1PNgY7U4LuqQZ3tdg==
`protect END_PROTECTED
