`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ue3jR2+5g8vr5ONgT0fbkICqwvkG4kY/cD7l52FmNuzn2qIF/9bD7iWlKZfDI0EV
qgz6s8uAjMSeNfF0cEyhBo6f1N1Ys2S68Cw+KQSutJT1jceobVOKnRTeOJEgmEXm
5kkDU2U0VyjmiocsVMNVaWx6DoJZ/HMkD312ydJPLR1LKmmXgv51DzZky7gEwhAE
sEwb43Uhkucm13K10fqMem4lAVIUjiiy4JLxSo1PcJQHAwAZ/DEGUC1LTcMgTUaI
9wlUxqed4G16BsWYrLtsBXQLQb28D4WTb5TfcIe5vtC/bx5OJfjFA/c+0cJj7cF2
Nwh7n7D+5NYyOtK0eT7stuJ808vrmVzBrCJzYyvciFuuORLU+5a7/q3W/NQnbwq1
bk7nUgjakWUB4NZYmU6HNrGybzlKJZQK3oXm1HRMVicTdqTW6SV5ym1zSaJgTSN9
IxOhEJ1N61NL1p/d1TBGMfkTxZPJ4Iof7taBCRA9OTuorALIw0xBIMjLE9Nf7VpL
T/84pW3hY44KIlfv/LsXegu2DWcYPvDTzv5Uf2AEfH+XzjxCrpaq0HioMwjLcb44
8kCaHULt6671aAUlCw3oJ09nFJ0r16JqwmwniG7wcaEJD0A18r/y02hAQH4vLaTN
v9s18ckb4ybrIIT5sJHdKq3EwLimZefVMZ4cGUFaF8wRzAIRL79ULb/uonVaR77y
VdriqABoXf6YXF009LQS5zAsV+qnFWKgmJjKsav3OiAQLnxicyyawomLPGploAA/
HBruDrNvE3EgfiU0Z8wnUK/pd7dHt0MUzCQxI7vIRxpzXnisK/oJuyV0FyihARw6
XSyYuR2qz7uHyhZDVJtN3RCqp02ik7zm4Q+RR+S6/7Tc1tujYe9mBEnESldc8kY+
5pqn9eZZ0hTrYXx4dEREgfIc66QdD/YRBrErOPXaZ4rA7PGaTHL3P2R/eU2Y/guj
Mljzjwg+09Uk10lXnCbaZfCTxdwX6PECovgHTc7RjuI/BPpJVZ3nnGtM/HeKpj6x
uHtqlpWUPSvkiDedtomLq0YuoNrmCEIGhVfzWfU1bjuOLkHKSyjW3QhZ0+SJ3yGu
Nx9COYbTm3nTYAO763PG2MXK4o4z+ZSgvenkynceR5ZYaEFJEL82pX++xvI9qVef
FKMdjNtKM4F2nvfQiCrZe54PsN9YTYdFu18V4Vfhi+Zwm9RzB8CW0TmDcXY8Calj
k8f/LIqQSMvrHdDXpb2y0BCQEtX7hJXFJoQMelLU+BPAq5d+18RjPhp+bEISbcfM
hhXlS80WlQuyRgf+HWlR/FNw50SWn7fo5bEYDZNHz2+du+QZyWJNXTWBPRQgYwqN
0OW0hQ4c9BTsFUUhx0jbflr3aGLFwZNDiayBA0pLC1rq+u8SZDnls3qMTmS4sewq
8u8xO5bwQCjonvjzZeYSv5tmMvQQkPLAoM73OwDklw0NGqTnStgCiLGcMWGGeEaI
wCgs91Wb0VvcCQ5+IOznSFrmJMvQLGCWZmui+ZBREnJGbGeASss4ujcvVW7iFMZC
4e/BnZqht7LJm3uQq/Wu4uI8MAyHxLv7o2+uCK+P2ECf7K3TY3LmDZ9g6SHoN54s
7EdbZ8G0WCiaAEcVC7W+Zemz4Ouy5oXkGgLU7/AE9W5VsCmvAArFUdt5BvXf81Ae
+am4q3n7yYwumb63NiyAPq78qeJh2lVjRDZKxCROhs0hXV/s7GvWUzYNwpbAfgSB
fy3K/m3T6ooyWfHRzukHTmrPZ0TXtNphERkOfTxN0qtEcEpAnKEfbUbA+/vu/3Bf
lgGZODVkiFrtAxQqhJzzklJSnwvLksPyBsDGWnCbnQ1uFB3+IT6nEO+amdzmnMC8
OJYxBYK1IozlWzRmOQifBRXX24Mc2IUUIui+PTahZ1HGmAWZAZhtHw7LWVnOo7iV
qG5Di0tJ5X7AXSvCewGbQBQeD7OzW8hx1T6rzncX+cMrp0MPUqmz7fM+lea8ObT1
1AxJ4JNZRtY5CvmuyMxZCnxq53cY5uh4HOKsLSPXwhYPsMS+m08eJ9M/zUBLtZSe
vfG8Ycj53sxM1sPh0tQ9fJ/rnHKH+pArIsABL1Rop5HNgq2xoFmspwumf8YpYviR
pDDp3MTZGz6wYZrXCCH5hETajS3i3bK0mhW5xjtEaligFvvLIQV+K8FUBJzbu5YZ
MYdHSl8xGjtRxR+q+rX0J9kIRiz7jG+wBFUuW6jHDxJl3lqu3+FIV3uzzWc4RzTu
gr/SKMFdnT/oiPmw9kcuue+ZGRRsx6J8hh87oV04McxyIvBcAqpaxQZeMOBlsCX+
PXsFnJn2Z8dmZjWKToQBaUA672mrdTQic1/xQKAEFqvEHeehM5UXsRN1Jx9alJFx
kXd6m4tI60M5rB1qXz//XSSAlPwSwAm9PGV5PuRQ7bCWsG6uZJuOpexTR90OFx2P
uqZktcE7+4HGtrVepjJWfZaAJlkoXefjJG+XGQmrogiVRUHzDCCbyJXW1FUrwbCl
Ksfns/8snEED4sPtz0eLEbd6JmvuX6blaIeTavt++52VsE+mDh4aOMqAQbXLjqLm
EP3gf73Fx2l0+IJFafIAGMHyj7BgvQs+HqVM5fxd0D0RET+Da4hp/CJ9j4hV+ZUQ
P+LKjwv/KT6U20ggFL8YoGvGsXwsHMSpwx5GgIuKIt06+NBhIGKicy151TH90CD7
GyC9hOYLM7TY0Kl47m1Hhnj2L05unK5AjJEHApqNl3LgMXU9R9U3wNdXskYQJBWt
6kPamacQCQO30sZZslrjk/RpLoFPC2biu/c5if4MHo9sTOWcPuQHyTuFCuG4DjlS
30D5NS/5ghJ3NPQUuNJACS4r3WWRb9/QPxqzmNUFK08XvaV1Ttqdl3xkeGuEjZBQ
mlL2/G4iuahwuI09mU6vt7qoPctQ8IbDRhxKmfJvRjc8dZPLdH5GqJS0jx+2GQpW
FrC4eRQp3D55PYbIw0V57LlKALXHcELfxHTX3OFSi4v0gJS3TQ/D7MNHbfVaMfox
8dzxrVYe5A85mEHuxGkcrWXVuOb1Tj65X3/WKdv9WMM8ElWVDhmytNI2TsWqNVTO
sPOkNA0OCC1EZ1sw4l71G/ujLdQk0WW63HAekAHxSNZb0ByzDOvV6ReQvLLyduOM
Mpp2teykrRE6dT6CcMCtMCF6oz6GXfwj0p1cf1ud7vacLj1fTJgn75PqXlYdiRCE
DUDuOn0LNU4lJgYssn+nHoAn73mb/dWMW9HCVWz9/RF20g38nChrFAMYBHUxXoeE
fVZdEg0V+XSw6n/6hrt2kLoUd2/iEPWoYURF7MbtokWKEQyKTWSE5pT9qDuVmi0M
cVy9h2D6dXgv8H4rA2On7vq90vcLKnBIP0GonTN2wXCpHS8FucxqU5XwoiNBjICQ
jbg696WfbcE2C4Qw4bxRYD1IiEaa2+UXU/6OA6V8blSN8C3fP0dhdrNitKBA1Fxu
Fh8jnqGM10OtR/+m00jlG4AsL+0S1O6cV7pPpGjkIMgbjZfVsNEJByvE69gf9v8j
reLBkfbD0bWlD3XPOR0QdKhWyM9tH5QMX+OV/mYl3KCym6x7+111UTzh1Or5/7Uz
nfUFbHGwnRDp1LYATewQNKh7m6YrFnVQOWIpBi2moQCeRBV+J9ZzUvQ6Oy6yRFHB
lcY4YO29nyqMBiNypWRWQrOfi0DSMvkxb8vAHcEzdf1UcmnUC1kyXSl7tPRBENOQ
FcURE7/Zva8CW+rBl4bt+WpWcpGyhtmjjAcE1Thq2IE90kA13f61XUZxVhES/f9y
N8wSd8jSiQsEh6xD7vw0wsImSrVg5rflf2EkMkVo3RUFt3SDpQMABGJYAOfJmgDs
DF0zYyh54guQI6UExrxIBbIbBxKiug3BcJ8lClm18l7rgFDmieARSufyT+bHnCuC
jw6yMCk+1bFaza227LTowjszvTWS7AI+CZriH0KIxzmD+1Y/2SNjdLQIoEHwex/L
PwLgFzWoz1ft2Cgtw9zrKe8H7fp4oPoU31aMuy9t5MCn55FuV785E8SupC8vkrwj
S0dcbptzzWJs6QUzce6aFYlGdywUkC+MNP/HVw8nyneBLu0WfsCeVwM0YfqvEKmG
g0CXNS0es5k7Y/HvbwX7m9d3JagfTBcwffavit6MCXq37Is039Ax0V1mWBGj95zb
Ol0tWRSwZAOQ3x9QRdgZ0qZWJop9X9EcI8yDVTCnp3vV3Sq0IivB26aedh4rqvFW
4hWab3a4fpwnMjBz5mKr0tBhhKXdzBHlMlMUy89N2zoxwE2BRXA02Lh57kcjtVN8
nH8GzVicwv27fP6R99fRwrCrY5NmOdghMFdLdnf6pDx6duea8kU6YBP/N6diqdB+
hlscnXxWEwbamhG6ytwT2StFAdlU71DZTMzaHVWyc/EBzsrefNtvSMwo2Azbi+XL
b5AOwHz+GlE7OgrT3EIah214aLPtN3TUX3WFq1MtE5ILvTRaJV1nDeg+3FsnBseY
LAJI5iTa5MD/PzhxKoQ9E0LrQ+VSZnwtrxf4LIciSoDnpfKF1uFWex0C/mRFxvoe
eJ7XTYkNsdaGZqhI9RnxLcZes7loMgTfYP1t5Jfwe/oZuQp1vWRBhUoUmsGvj6np
BrKEqgPfFBkju04wXtkufRqvw20BVprtdst1bJaymlXYGF0KkujS8GqmV15d0IxB
9xLL34T60iiKEbJSrq7WWKl/U7vKhLfxq9V74sioEBASDNmHHvUD8kpmRBCW+t19
vKN2Msc4UGJd4fNY/LjtBNLVMRfHQhpWt6EPcmK3+K7bRQ7+/x/IzoPhT2KcKnYd
BNXExGnOSAR/3xgcViaQ/cox3Wp44ALYbiBXJ181vjk+V+/WWw5JfC4vKEwh3ZZ6
yIPsm7aiE9HbpOzKlF8SmekgCOOCuPhs0Qa2S/TF2CjBV+pLQYL48hyIlKwWU9sO
KXMXL9QsLi9newmKfZtJWEXVWgzCCcUBU5Tmhe9KIRN/yFDdZ7u67TTdzz+yWAp9
gDUZg4aLN3Cy4VieVBF3e/nErXb24xBs62yHsOq34fP86i077RRcsa4FVjHiXVz5
ZN3jbMO/KYZfrSkbwbP+uZYiBewtvg13IUf/c4ti0szciAtnnONt6ZueA0VeoF/M
LYDCaGVD91Sd+SW0C/kZYfiXTmuMs5wty7ztwvIvjp08hvLNHzHvctSldkmcoOH2
F56l0RbGSd5pP0057NAaZGfcFNqsOVhr8ONC9QPEVnS33QWwZnGgoYJxcYOJgRb7
sUsI3jJFh82BYRr9vVNTnLQg8ZlC3BXDN2Fi0dg86MkOWo69/pJFFFOu2S/W1GWO
uatu+fXsJiwqW9EZu+xBoXv5ogtteLrRuEvYPUT77AdFhTzHEkbbzJAHFWSnLsPC
kG31GTAdVBM5nRn36nRfcVdVdIi71K12SX/BkKyOOsYk+HL5Feuitr+/6TpiSBto
O9AA8IFeaO37DDP4X4Yvv9Gx15doCWWjRNtyzS17a2spPXZBf8te/xEkqK8hccan
udvVUX9RKd5vQpRwqJNZynKI+fFS8BzwLPM9x+Hfw3MQYN3L7sXD0tif5FLi7Tln
0LRYpxq5Hs6tRgSeFjpUwn4SSxsa/bDGzWOpKEj3IMJlQFlXHR5ILv3jzNWMA8Ah
STQdCjljksmu/jCH5VviYeAEOglOgTod0oAdbveCfvISvHHX7L4DeO5ahN7F1sxQ
glOOs0cAmp5jFo2iiW9pzbIAjYczOfkUMSXg9W65JyTF9qwR+Qk11xxBEPzWQB3f
i+4NEA1uhqHy1UwSwG5Cyji0iHJJWn4sMBWvVdetFi4z8GvqAngen1n7eRLq6ms6
9aC078Bon+fBwxqTS2jljSApdzn8TZBZ2ZlUmqh47PCdNnXpPj4xiq9g96hBWUgK
B/MriiAG7hMvj30ehAFIw39ckugPV21GSNVzc1h9vOEMlyVxHvVPrljNpmLx9w2F
Vu2AGAU8oCP0m8iLD77exWhm0CoTxJ8AnpVcBdMpknH5c+XTY4aNSY2cZQOgITyO
dCWbbykz/YlQfqeue9p5O56CqGKFhdz5/dQiaWjf6pybIkJnPioNBpdjt6ttBuMu
uutCSQHmh35OV77d2M33T+F1Y2J3u809rIktTKN6LZsSUoDv6rd+ceowgQ/bPiMW
ngmTTy2VRkvG0F7YfExvqwq0sWBNadLaOm7kBW0aMW/fFa4T+0RqeByPts95dDmu
+cNLXt5qPG+qBiuZQQbpDMatpaf0TpUODeu4e3ChQ6EGc88Ohl9XkjEj74FbXF9E
iuB5hqbLYrnKCCLxIj7ITBjnjVXoqcEsj1QztK35NBcl+0v8Dt8GHD1QbQslCG57
lAdpTVhmxVNnA7K/BTwz6X8+3b/C8MFu4tTlptFf9Z3wZVVT/sM9HBMzaLzYaYrs
elqjDTUDk+LWRNDCBRJErRhkej/skk69MbQmRf192dGhdOW7zoFsnVfQYy6Bnj7f
mqwOeVMC16kFWi5fL9Mp/tYyQxgxnTiIKXSGT1SABqAoLgxq4Tx6DlVaerss/Ygq
JQbRrLc1/0qgj033jaaScjvfjH+/FiAibhc+ZA91Nb1hS/DywRRGzb/+XWUGlJT1
0DmgBD0Yw58bAvOm3R/XMi2a/68zWl1ciCG6EhugnXNt+RaTgy0GYOL+8joZoo5h
Eix1ceWYuASYNtxPwRytRJAS3zhoY3AbGoQu1xHN5V8r79YGz9lrYTDcgkxD2n5L
qcNYwboIl2t8Y+H5IyolR5j3LXFJFbN2xOvdjhzDQY6jRCTmwGafi1168rBhiRlG
VemnEu9sNCGwQ5QUHkAzlrKg2ULPm5R1Mhl6sJcw9NDMPSvLnF/IqOaoFbAsJ5EF
xVkcIBatCL4ADTixNh3XwHviuCTgh08j0ykYCkn/rFpfwV94CaPJdhCNajrxVts0
k1mAcRWxio024/ZjLmPcEa/R1ir6eYaWtzJD3g5TGOiBWl3lVmzXbzCscaq9o+MI
iYHRe4ghSm8zktKYRkvWmVXchOQr1B0N1ok0d6N+/kuxMJakuBUgm79N7QZ7O85g
X9ex/WUDmlZAnkEk7l+O/l7br1f0COdkn4ky6xuHHrE3QLtmkXn4wTi0agkez2nU
UXnV20D9LcrvML1oRF6O1nkfQBte+FwVyhLlqYYb1N40FPpJ/tPMt0r7oasyWgFh
w+J2A2tF7iOKA/2GaQURKh8t+/WEORaRvLc6qk0C+60i610fFU06GDIP+3yfcFv3
x5OGiWecVsrTkSecpka0D9QzKaBXk6yoHz5wlY6sGlDkH/sI07jKpQQt8guyy14x
pAnsBD2mUNbeAdVN7sn66Ld0x5abqrL4jSswgy66rbnko19BWn2byPLvw3otNu/I
yyfSeGQeiN7rs/osP+E0WLa1niPa735hFoEgOGxOIRST/Z0oBYRBLqJf0LYSyzuH
LybO38l9hPpUkvQ8pBLsQdvRLsP69Aqe70mZUWhSS4ZP8uSLcoSgLgi4j853YXNc
+ZlW9jKnkjYP+Q2ZloSkWhPNksBXKjbDnAzQ9ub+HCpjU5OWu0m3FL2XYj1KNQhi
Daz+Mxcyy78WKjeUaA5cLQR/vaPOn4Wssn6/1xrTQd+yP4u9EXB67HmT57AY90z7
9mIfd7tqvUyjGDbJWVFGXa1OwGxCAj7H1dANt/ZDXhIXiWNkJTC/svblHtTbWUvT
MKwMNWpzj1TKy7seRzQKtut/G7p7lEMgUnSRcSCq3+q+CTVX5Q+Es9JkdDhdokpS
UVgjP2zchLZ0b+ok6n7kz79rx5CpBoVXQ9QJ/Isi1giqEBvP8BPUVYB3t9g35X96
t8dEsHchixuWL50kkYHGfQ==
`protect END_PROTECTED
