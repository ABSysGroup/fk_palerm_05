`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5k+tj+qNJfZGAQIUg5PCLl0bFw/n73EesIaOZqmEzCf3TDfZJeFKwUcxuvztDhnr
MQudnt7nm4rYgWF45b9KphxnwPCx07q5flj53kl3Iqffo/ruU0Qpy8FF1OE4hkn3
4UaQ/t4FGyovvs948j023c4jb+3I2GLYgS7+cE8j3koP3ZkSTT/8t5JwoVqfbRZ6
PD611r3sjNoEbN47vyzandfUaQfgfOywDVJPG1dlluLsjgVYoV/CV2F3CxDnYA+j
vCohUDlSW4P9esx3/UaP2VGbVMXg5G/HyaV2Fh+dqArd8bmKubezeTcI72fEGXoA
g0xxyVuBiubUK28FwGhX/dkhxVS726FZ7ZsO4lbNtFM41zSnTCUCUiKRtUPm5ZJk
5WQtv5Mz98sCH+6T4yxszwmZt7lGIa+S3rtjbqMOdrH43eN0PP4jDCMPy3/cMjUy
OIgdIH5WgYgt/ePtFFnopaQk+X1vG0CGHDl7kuoth1/pMuaAjPSxwaU9m/cvi9/B
9RGxjPbhCUIws6ybaay53UCv3IFm/LAD+qmu/pAWTm0J3MhUlcHIlYLYe7eNApBv
HPpgkIq6Q2PPPGT+fCyRjx6MU/azdAvGauReWgfpG6G8owIS41zo+JK9xU23/B5B
zk9zCESGkjz0/vEwCZkehYy9GKb4oeaMZZb4iIENeIUd52GCJJ7jWzAFI3kApRMc
3Mpo9pwR6w1BqQ1vvr99u4iaM0e3IATdeRvYAAIJS9iW8muqOkvwxJZa6rzfWimR
8CTOzSA2znyj7+UGq1x9Vlf9FUcXuqMQIaUJpPS6iYMBQHdvihkA+EVYmmlBWA13
VbT1JtgESNVW7z/4g/n0yRUGL3kUEOZOVzHEgPcNNzeYFCm1ugIQt5w20kHT5MnN
0Ttc/LUjoaYQNyQrF597OzMytbE7KCGN9NjK4jakbmGqaA+/2NlFtto1gSPFA6Ta
LfElED/fOn2tXNChVIi9si7TihR8o8z1yzcXVjcEy7fbx06/u16j9cvZNz9xLec2
zIx4qxJfKuZkKDJBA0ONHgWWyN8Nl6Xq+WeuYQS32t7erOr1zy8CQgKFiDeJSEaD
09pBkfUX2OyLlGSQ8s0c+omPg4sJ/8yNGLwMr2MsbaMsnq16YU1b5aTxbXtUzglr
WqRaJaA1Ru4qLM2e7Vf5DTEiHjoskaIQXO51PhxMz4pObFIMysQb0Xmg7IDr4joX
JeFA+OpPJNUN8PgdWPE2f6A4/2fryk43Df1BN/aYPwJ1YOLkw5Qes9t0oIZu//S9
VD7eleSHxlO/j6EjPG5kIIG8gmPs4Wp2qDHk8vAgu0mbZ8kLwHxH316JNZBt4H5E
53RND6USAbSzU5IcbUEPHF/7sHX4/gDquFnOQowi07mKHJaT6BqUp1YIGYRX8MMs
`protect END_PROTECTED
