`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YFhKx6vjwlOzcfSuysdeoOl45B9yf/aljx+7/l/riOvf49Oer4U20VpLmssbffgq
83ChtyHqsw2KkexoqybtFcV5wansgR8PoPyLSnqsIxb4W5pE3uzH7eI401LRdlEz
TMbTWkSc23+MfWoFmMLZ6mBC07IfefX47NcNKykakZVQsroEqhCl+/tx3LW4HMZn
3MXimx3N6Ig3SG6ABVUEIITow7ACu/Dh5u9nnwlCy319a2O04z6/xjiSuGJWYMz5
Q6DZkcYuMWKhMkydS9MrCw==
`protect END_PROTECTED
