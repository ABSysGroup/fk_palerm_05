`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LyuKdb0qWO3qV/FMyEc+v86xKIZz7V3aaCKxz7A6oJHtXCOgAIqtPrzQo5ptOS0e
vgSSNVsf9wNY/6Gc61W+O7DaPyrjD7BupNtmNOykrmvfPfCe6gO430fjv2nQzxYz
wzew+ihrvbUj2S9dE4+mFppJpskXonaFQuAABZFYzZCo/IfiPvOCFgagThQZGFPQ
Oxs1Slo0WbEMBCW1uIq82KUdJfQnkozxWNDfW1Tt0YM0cuTfiYdxA9d/BDVqf5pf
YYp/q3Mq7ZjAOFG55aJP9OcljaMEMh+vhjzYnSz3BsPG+69vZ9hdQcBQyABqgfhH
8BmmKc8N8rAyf4IM/AuO5N1Kwd9qyczA9n8d1DvKSqfskm8XqDMACxhP09P7RTto
Yb7izTiPMX588dpjCwAIhO4MjQmWRQ/+Y/A+C/y1wpF1b06OqqZ3YDSnlkLUsDpa
GHSqdTMBRQBhXYAHqJNJtEhtZ3eygyCL80G6hB/8OVhOcbWlMo9nf3aA3Bfm77rV
WlcpWshwNVvoHCmQAlb+F+XIAPAJgslh5qJgH14Gi1QpPw+9EsIFgQZAiaO3OJox
SYTLqB6UkMYwooBpt2KfOeLp3+RaAizrtH6DDEWtOo+3EqgRVRn+LJq9+W6RrLOh
H4kGCIhMFocosgtY8pUu55HiOrAaim1fP+jxOXJFXgBX3kZPypHLHh3XB34jftaX
HPqlFU+IvsLi1QkvtmLUyvNnqo2uKmQ+v+b43uQjdak=
`protect END_PROTECTED
