`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5YL0GcZCdH0SDidVJxzCTRpf+4DyRwxbVvrtoEAMWLJFUZ7p3RXoh2/yZzSuWYmM
FS6N33RFTrOLjC/+yFE14m4bNS2F4vxJPM4Zy4K6GJhL3c4Wkc0w2OoADHx0EKVq
phYjoNxUZwkZ/P2zRqnmOQ==
`protect END_PROTECTED
