`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AH/gjc/OrEFO2C1ZbX9wLc5CvAyu12LiOe6jZUgJ9qdwp/BQ+qkf1jP2LWOMuMNu
bUhVIFWwfhddAXZbesofTcFVrvQbtY6tW8kihUziBgEfKuA/VPorbiCFlx9coLvV
qHax/0cFFMwssJMZoTAe0EF1BSP//KXVhpzo4Lnlj2audJzJbM4PH9cCShp+Wryr
fQ/a59Tf2dZPH0qfSz27OhbJXOSIbP91DqBIedx3BFikxRxz0C7e+fmKMadZ8XWq
55EOiSzV9AYCO8/pkmIQwUbw+lSbJrFUU8aa612BSRwidDvi5GC4YmnbOV2xItHH
elbEr9DGMGE9ySUS2obkv35Hwhnk2onXgd6OZwxcZ83+6yjFgve4axrdb1avuYnl
BHlx6DQZv5TU8fqH3yX0ym15oaB72sWLd4M6EHD6EEsyvTChavFdQ0AtfJiBo7BF
h91OOKi5ZESuWaDqXg1H9Q5do+VTCk0/6IxOVxqjj8dTml7tfjm4si9OUrcR3ABo
G2B3lwCo4dtOLFXKaQENgJZxB9KJBjrRchUdUm65RyRF5jK3XSNNVY055RdcMXmW
heEzfu5a8asSlIrhs9KNA6aMcfg2MvYRP8QoldSvjiXUsTQzJWmtZTz8885G50QS
L2pW/ue6fb1FByeSK/sWuGWX9EyZTsUoLO2N4N/IE//vdfkWPj9ThqA3E/td1Hjk
ML4T7ZVM6CHJ7nv4wHepWGX1h9h4AlbYb5JSmmAz1KLFNGu9WpFDCx+Jt9xUbtoI
fEj1zPvLXF9VPAUcwN5gsg==
`protect END_PROTECTED
