`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e8pOi9LgVPt4YJrhVQIozmv6UQf2NpTkfDqZiu3at4n1zPrAGClvmPqKfUZZX2Jl
Mj3Hl3iLNOQvGf0YzUOVDM4WwTpyeMIJubrDUD6hloLOziIn5FKk6Z5zRfI2MwUm
9KqhMhJXEfGp+b3/Q0LdvZv7NeugS3zkav6yK19PNS5B02iI7iiwFNqan6TpcayO
6wyDPGZ/maOBmDl05aBhTgRxC7KTFKF/4gGO5JLVKMAWlCUoDpMY4KmoKKcp28cr
G/ANYXuHLPGjTBzBKmOtB4+A0EyEAjSGyPDv9TVtUShD6E3hyCg+sG7wvT8xMXOA
4y6gfmvZ3rcRZmlJCtI6yYUOZbh/YBQu1wIBEBsuQxvHAIk5uRUeKwMPoRNKocD7
w1Lsi80kIeK6K4muA+l4r/m5QaXrCgw2YtBbRM+OUPDON7I35/bYUImOb3/zj960
R7Ag+JLWFD+4RC6k3qgDAs3SQq4BeYEIlW7yiUj3fIp4JqXRcXonYVsKOzo30GOW
6Qxkr/tDLdqjvmCVq21jH+PHZepW/mIgSYV42E3HVg20gOb6K95J73CeC4mGx+4c
qPK0f2Ln4VI99uNjrsnjOiQ5spTGwtM1UTyhCBQz6BwHjrfkR7vxeQIDTIeRp/A0
ZDyTmJ8TIA+Je1KFehNU2Nkf4x1ZXiak/q7Cov5TBH2V8s8r8zNkHqDak1FJHqW3
Iv45CGTPPsGrnsAXMdlfhJcceSCdT3RDyw4X0bnTQawP0MqpUpR5p9n8ao7Xg9ft
pQGrwBOln/9UmNL+ER96/n/sF68j107hPjSKSYdlKpWBEBI2HuXuaPmiauP6Obas
qmhuhn9rGtWrAumo7pVCA7qZa0C0Kyc3I71LcYFcpzovq659A22WdIUi22/Pumso
ZZfC5lX9JEADBObjwkS4J1dDqWUY8jadHS9xGGkr7egPN6hO6xXhljfDYp+cxgVj
`protect END_PROTECTED
