`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V3rbZL3lDU2V7YTRHQC5VEKVJ10xRACku6P/MEXfqIb7UG/Hx7mWHvKNuARJXjQe
Z9ma79JSH0TAK0Jt2f4hlRDdK2+TGlydcwSFgVk10LefKyIkdUjtkz2M6FmYu6XG
D4uqBgR3PegudZfpFtzcTHqmCgiYfq8Jx2CiNQrLKZaww+jHBS/99ALqZFI5ical
daZtMhSHfp8M/weM2WBeHwmVn40TpqGODeNTAH/iIweuEM21Fr0Y2YCvMe5cn/Wz
Z4dwUBchKtqogNYGdrOAKFYN6rC/2DX/wYwH/AuV4L/vRIrG8BitEQyoBEzCoIxm
GwULLk7z78JL4gjWLQ1VFdDRORof42P60kvmKNEBrto8ndv10upyGdkmiIAdfOtp
ZSDsRyygL6w4vsN2WiFKpqoT++ruCE3qtzSOLRcLw8/HCIcg18/QTibvQTaW8JVe
dvW8a2HpjyfzNFlQW9mtTbX67aRgj42ayP/7aN5HQHRW3Gel5SaR5I307ydhZS5o
g0i79XjUNBsv0EnGFdleio2XCG78Qltr6smSkuCYqSqOKeYoXkdIBmW/Z78r+6fv
oFaFl71LBKrtoN3d0Aw52VjkZnYERciY0i6ie0u4nuE0Qrg1R7NRXteco0FfUnbV
X3SznsLeKvjeT8qy82rqqaZXsgcftqp5RJUGR6Su0qTcjMEN9t0lbRFH5dbTgzn9
ae4tET8pT070aBXkdtdvR2PXifDJbmc7u5Kns3opjvIGeEtRxODN6iQCK3a4WM0+
PYLcQVr7MaYZ/Y6BEeoh/YhUrwUxVPbtfZ4QRu5S+G01I/hPiTvji04F9+/lMxMp
QVwToB5fbRUsZcdGhXFvEQ==
`protect END_PROTECTED
