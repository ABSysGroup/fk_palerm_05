`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Z2H8z6OdEy0UlkQJF+WQ6AT3zjY50tNDlUT8YIMWHUdKi60UeUmu4Hv5bPZsrG/
Z+v9KXjuKJqzGZUvODTsdY1WJ7CKsy4o8sfw+9MVu+eaUSumzAy+0Osl7yc14wEF
8e9pBE22Bn22BZF9pmgOoMsYuOf6Z+eQ4G6kEsPLJAA+zwz3Y6lbylnGkYzj2uAZ
j9cf0wxLgxmV4P3v+dzIFA+5ye8BWy6PfXK7wP75RRYZp6xLGaO+aaVAVLWp/JML
0VWD0FFc+fqMxMvUtOWLy8qKxkvCIZj/PJZuKymBgjAokCxwGFRnX3uhK4wirZmn
uwIAIYcqcKLtqTjzBPvIdGbqBGO/G0LvvWhklrgyGeQJMD6EYCV0zr1GLHc29Q3J
50wyyZjNUk1n3KCo1Uahs75cG+WA5uiyAfhXrJ/cPmzQfGdF39tXQDr6n0hk0aDG
tQluaI+Xoyt3AoXbarIaZk1syymqPyUBTatW3UBIjKyo7df+zIy1wluzUrCC6ztw
0s6Q/16cY8NdRau9UwDf8Yjl89lGSSVCXmUqC08Tr6UzneTej62mtwHbE346enGE
Gfs0qxqNVdcAbNjsz+p1ApuBofY5AtQxFOOhH4hMxb0gIhsbWxhWQRsdHI7LfJv2
FJBZXVwt7LVGQ9p9XbDnzwxhzYIpO0FyDTY9YKJuyBsPuD9+SIlh3Uj/V/25z5+D
FWOGZztPvYcDt08XsljAFPOmWZGjud4HaB3aonRjDXSd7FAJTvPqWKIAnm+4Xyqd
dkhzzWyDOnAd+0U1+gf0/tB3oAwViGhYs5znB12eMdB/jBQ+dANO80I9qUw6oYqq
6I7NoVKYlNWKG6ITmtWCXXnEZyqvdQ48ji9/iFogMe1MQc0RTNP2uWp1sh5KeGgg
GoN9uRrKz10sHeAQU9QhzGmSjQjg/C2cP5CMDHAVVYlArHn7S16iSJiU4dAxAXoQ
VlVCi1sORJ/TByhZYj5g4A==
`protect END_PROTECTED
