`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0a8a5yrxZUdyeh2sHyW4t5L4uyacLAvR+xNO60fItBTlLmu1ltsbqQV07C0p6KnF
4q3qdeQzEJyYmOcUQ2XA/+fSPfao3WO+FYgyAHCEZbAyqYU6ZZeH4wy3Z5C7wy6p
OLSsC1QIezj3XRNcD7rXK1xfrdWZqP+A4L1V6KiUVlWixYlbrzCw8HzH/ZetF5gn
pVy+dwg2oiYKYITKgwM+sG4q0sGzTsjelViRy58tiq3HsHzv3sHiSX9spAr+nPNs
OfY+M5i1JuKkJcNVwkqA1f2gNraQcWmy9jz6qtslgSMuMS8icPhzdMJrCXQoEcrM
QJcQ7zyqG3v/ERuuXQkjvC2vrqk0MGcVsfkywuEAkROVAv9elA/DyBqVV+UIH2jl
uzdHDxShtuqvaI6RaL6O45Oc8Drt8gzOiYUfwpvaE3bdaTJVINGE/F29w2Bj/E9w
7/juy6KpK9KmWZeZjDp6MX1QdWICgDjiH9YOTlniSIP/4qVBCNUQ2mB2DOPAM1db
tPBGR/SX0h6YK2tJ8GpEqTgJIddkOfPWcuGb7XkBkTBLA+DCRXKvuxpdLFaWTQBn
Hsms6LFb8U6IS5AOhN2K5FA1HYDXecAaD4jUXzU6QT88bUYsOoffYI+kaEini2/2
`protect END_PROTECTED
