`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vVZpQM9DNQ/U0YqdDsaC10OSxmpwhNxwtmjmWDCZJ6KzL5s4DOiAiSJkb5qlN1g3
wGkj+ZfEmR803AEWw8nIN8OfQDgZkFUp54AKc3MvJuyMt7lwEL4v2uB4UPwYfVKJ
8Ahmt4oqv9+Dg4szcfBZi3CA+67GmiDWhoR6jrJwnJcdRUr8vtJ5RVVlEPI2Wc+o
wx2jXtf4r+dWRZpq4PTaUCefbIbVP+H5oWaC6PRA1X0ZVs7f7aeGgYiM8q3YGVje
KRbRvsWMP1gWUFnZGBUcPYmZN3P7TYPLOj0EwTAB2t+4F9BynS5LRhF2QYLbbRMr
mDFtUmM3kT1F+cYwxX6REy9fdQChvdQBBMo1LQQwaXui8k/xVVBQzUbACZpfuGWU
vImivEO5XEHIThwUmPwhLpa7L3vLYHoKKugLOgk5wdnGAoPZPZkjv9CqQf1Fjvw3
5UP+YRpc0M0cyFdAd5rakOLxqmqxUWWBqWTEYM4f7wSlKquqrkgFK+MYP3/97ffY
JH764fwyAV0cFJomoNMpBhDEkP41eUFXwYbWJtkG6Zpkbor1UaxiGvyYbtq4yEsr
XGYsP1O2kOnKjn0aQ2YL01Qlg55VHEEvzn22lBDn0FZKQeOZvfmO8HqhrqN+qpg3
nmU9kNPavWGszgeBmJ/xWA==
`protect END_PROTECTED
