`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xFhxGtgewZRtCgaEVVKBDRUg7zD/DelRhOmEUKF9+mTIMcikgDPK93IEiA8nnCvk
e0VbMrc6OBQ2AjXPJKXFBsRQX1qL6y7VcufMWb/M75Fm0ccrH0HNHt4UjHoB7edN
Ab3e5vOF2YNrxJK25TYY0K073GBGbwTSMdPMzY1DHICNOU9BRCeRBRe79XHCy1m4
5AE/Xe1uqpq1vNr6CvcpTB9WdRSsDXgGDyh/44opRtjxTp5+NWAyxXxTrlFnNVg2
9G7JkRVm6F7f7dbbfrLHPq8Eem0vCI3qthNnVSffBtTiqTNVUMKdUTF5kwR7rLbf
3Fnq8EL7Qck696jVcYp95Dl7KwFbJn7cJPvmP6KJyWNl+tB3d5z8cBJ733GFGx5G
N5tpAogCO98gYFZA9Az5WAbjolLZWm80sLMe9V/t5dqBtZBHETdXHhzaKXi1LPPW
2semV/e0jGjYrurZ3hhBa8jcdDauoC9/npgWP2ikJS21SKYWbZcytlwBnv24Jqda
F2Omj4M/OaVc7viAKt0Wpgcujy8TFmldA10O3/nhWzgC/TOsT1AxTUc8MRj3YT/G
mnrV8pHYJ8grfIthemgRO1deJuahurDmPuc4hkZ3fkgMRlybWV5oznjDAfV2+FxY
c+LmcquIIW+tMtEpAAF5QKyAAxZQVyhrKx2bTM4QA1lKyvjIH3Cf+K5BBXtHLn7s
8zWnQyV4IgiFnheq/xQVICVFiiYfPvTF8uJ013Bp/9Srr9hEvLpoMIne4Kg4hmoc
pYW1h5Ey8OiCvdAqx9rwB+NZXcYt7PIqx1QiJOOJp82gW331nddxVA3OmnRBSJ3i
1wXYPd/Z9BVIkjbvIWRLrRn/wxxAKoW2kevY0E7NoJDtxnxijDwVCOtbGBm/vKc1
9e0UW5b6iy3x4hpVPPvdOcKat0UFVxq/jVnhZe/bzDWWycROgw9fJN86//6D/nWr
/WPh8MpLVL/kBYcBJYLw2/KC+uiHZfOv4l7OoNaLTMS3+6RslebBGr+Is311Tr30
7AWhjZnliVtrmQfvWhf6cwiW8uG7CGEyN3Jau1mELdVT4/AdtZoL1gWMHPpX7fKU
uAz5T67w64zYJuD2Tr10t7bRAtSD703Lnjij9ZhFd1RJUybWorRsSJ8WMPn+pv/k
5UaJJxgK68hhWhEVms8ND6oQFW0HJFvuqCu90gkKXfEG7NyRs1UDDw4z5X/jaMPy
8y8g9OFaWHvwDVDDzrNoYmXtepYoByE8MmmZzRfnIQIS1fQ0hDBCO+MiwmnOeYBg
7bpN4eNPlCLafuZxi4JQH7dCdS15YwzykOJCo5ZQzw1TF1BQrNfhituud8rbGW2L
TseyDgFBiIvZGJrdi0U/nnMRyxmhl26hUEMOdSf2RdCEYDLC6jJHRkr/QjRDX2Re
p0VisQKPKC7aD/aDYwCBraxK9MS8xgYk/zdep5OOY0e1x8znRNuRk3QUg6mMIo3k
XBjTsxwjZP9HrMvhDTozVZQoyCyY4KFlRqNkpyILY08uUm8XU77KQEldydp8qzm5
sUMJ55llciS6OPXtNd4t3DjYtgudfQO2QNeUQ5f7Z0nhXXqLxCRvbEzSGRuj5E2B
JKIZOVl6R2rP/phRf1NEJgLxWF2mjDFaZPxv/EPbJYQFgHO3IgT8Pm2CWNlcLpKl
pxQgVGkOrcRY4EWSSRG/2Orv5AnKXpvPG34BDTOQ+uRi59/WRgmRYeZhEz4eHwFq
tenHELWQwngGITsgGtfMldpMT6ziTfyGxxqKwBcfTV7kdqB6KlgcqfHqVogEJdmT
WhfL5I78/iXQHdO+3aviU/OhgjZ5pdDnZQrtnzJq72cHB9U2COaIEVWzwrW326mJ
ykVeiXsWVak7dn8Zp2RLUtQgWd2duAwJJz0YdRplp7LN68VopCaCJgEVIYX6IArz
cbcidHFptfpQS/Bfm0f4w6xBYht5FvAMsHMUrp9oJqriJo4Fw4Cm6YlAL6r/dnlN
JVMTSVxeT01H9bpSSudWPArsCuw7LXsMx2xh1B+3C9kgF/qQwDXGdxCFsChJAclw
7nSsKa93Bscw+XcmXVVJNdOJJJscIOYYtQYTEdQFwx1OrcPJ780XOOb5Dd3VFVqI
4oDl6u/yd6mGn0PLy/mXd3fovGucgxcshZmwAalKJlJfsCYGJYvQGyrTBRFt2uL9
Vc7PPZktDPoDUTK+lVSMPUmZRRc1Zx4PZ+MdblY4vEQr6p4tkYzl5ALdgdrAc2cr
IQ5i4uOa1uvz1fxJRU8jo5FiwfvBJ8RDo2cdFuMAh8rzUaB7wLRK9wVdV3wlAHqX
AdpSQKUnlISEiMOai+su9RAunICkPsGL3QQgBA37C8mqwE9QVWJ+jmAzCzMBVhHY
5scedkQ0db/+59nT+BtGcQmM8uamaUsp17/2a6Vk41VrItQ83rm/EbefF2coGPcS
e74Z2U30sq2eo0IU30ULqf1sOPo+ZhVK8R1j2HoShxbP54vrt0G9376b8AHBzCQN
Rv5TRUzgQPTzO8YcFdWropVfFQB83jiaksesW+b4QcZd2HqGnTJVwMejKXwoSS0m
eikyP3EBfrCfRm1B0LlGqbYahYDoGRPC2La5iHddo9lBq9GqYOXqnRmBjM3Z8oqS
PABZzhzcuIHPlGMk6iI4cQky714wDIwSsdX8ZXSaX092iHk8zA62qHA6asafnl6I
guzgNQIUv2ffRlBOQKHTsBs9/orxyFCSMb0DRmje+zcFAg/BTSpqkfB/Ay9m9xmj
owyrseRcGOO3CgKsMzH1C4pYoCxqF8Pa/Olv7FN2XpFJSbPrbzFYF4vfJjRS059X
SkqqZjhHo3Y2Sp4QFiBAt1O2R5OUQXG1KR1wVOX5Dd5MKTE5928TJmfHJ5d8CbYl
QFvLpd7Ouo5dOByHxh3bYNf9oFZ3dy6XocKE1TPigWuKZDvHte78Qc9ITvt+kGvS
HnS7AV20QItEnptDLrrlq4qQd1/6Y6RfAHSxqgO10+RHeighT6UgM8p9I0ooBlgU
IuujFeIhejT63iG6JPqUehUh5k/elVjm429XCisrB+G8CZhTMHb29WJkZ/mVIOnK
5CGmbxKv4y0B9zs+A8CztQj8oHZYctNbbVBUpiEUNCMrdye6NFRHHwhKU6WfAKt3
KJow3XYsy3dZegSodf2IdcBQHXANeVSxZ94ME38JDVhmgdRPU1i22PB2U8OXg2KV
r4myOhrEhFRzI/0fY/HVqyGEIRLw5sZv4E3PmvljV2DscMbEMW8l3KkJKv0MbmW8
nRNLUcIspwgcJ1I6ZWoeoTeqH8qgY9FHvg0DGgGF7w2qOu1DyJDbRk8v57+07/vu
O6nY5BKTen4tw9XiNkzZ6AhGCqqSNfT26H82Je28WWDiLsbcgDk3qPUpcqX91nti
73jVdFuikGxl35feNF+FpPo74FXpAJpc2LmN83bX3hPd7uvvcyrS2RN7Mrwew1Qp
PBidh3n4ek12TdTYmNUyrw3E3Z7E3aDHf4U86KwQRBYhSWDjt0G1cmRHaNAV5TMF
LxWdUGe1HR+TLhNGkumKfo5xcnDqLExVV1ImuAYuz+QCL9+sTz+I4M+eD4+1Xxh8
+3c92HB8STu2CKO1pFxzVDuj2T76oY0KBI5sBV/Kq/F1XnUTi6+rOoqcjDpfg1RT
aTIHFmPOTy6D84lPSoxJmBYsa8XR0qhcq5dbepf1A2EG/vhoZKOkhHuv7e8UXClE
oAh513CGdhDQp93LFWlCjmgnc8BABtCG5o1rcdRFheFKDrtbFFuW/qUvaB8pSQu1
+zft6h9Q7NGhWhkolCk5ezPtqSgp2NqiPwfQrP3+xcBGfS+zIOq2e+zH9lBoB5Ey
UXNv2ZKTD6koaWK73vSIfXGqaOSICBSdiSWbL7HoCkdDLDW6dVDDY+Ofe30ZWIwA
6PFvEhnYRNZxYr/RHkk2trX8/BiWNW4bxvNe3ESGRVkU3MvaF9YcIcD6hvndSzET
4bf7zOzpIcUrxwzDBiveKs9pidXzMKkFvtndMOrinexz9q/ddoXO/tSvmZcuGAde
fkqsSo5/HUPPGmSEui3vPnqe26mVF5JFuik5vCGc8KPWATQU5TFhLE4WyVoDih97
ZmWYgy0ZynRropCnz5dt9m2t/W3lEp4/b6qdkuLDhpk6DhuiLdfaOlWt77+rbTtp
uLk7Ne/swhkyDAaga4pze8Nrqyoz+eHguyvkJuj+DStLRB+eW13X6dc/3i4143Vt
L1koVI7CYP8dWb7CfmeNrrKv8bFWKydObVHfu7DsJpnZgygtN0fFBbjQJo1ojLv7
Nng1p+oy0gVOE+VZGWzdSJJLAPmwmxeXo8klz6c1uEt73b/+HtWMn6lyWcDMergy
21BgLdAMmFpVZsneHGfAnLioFLu0KdIcBz4kcTHfvlfw6hDv/JdyfMMc2xfNlBzT
6MM4bc279RpRJdwIt7Oq+G7hvHU+0rV7OUT+FNqq5NJIj1Isw3X7Xm34KgMz1lAi
CQEohGflnkmW4fV5CQBO77ZUEpHzHw7SQWtuu5HrwbLZKMhKWXyuvjK6VB/w+s+R
yVE8LvAoqnas94hnNluTl1cBA0lQ9YnxHAKLi3vuSER1am80+U5RSgy4g9WbIO/P
7S7/efT0XxBS4P8XN0wkOLOorcaipsMuT9Cc0DxMW4LF8Yq4jy2Pu+vl2MxeNCwH
XYXi521JVaICt5VHbxXs1sp6etKG0Mdv6VvtGU4OTl6gMSuM819lTnCac6+UgQp0
rmwEG/gxFzGJaARS9rYOG0FDxbLMVNobFItSBwGkufQWoj2CaUbSDMpZGjJQTluM
TtwCdrqYAOX1rfH3Isr4X32NRGgM7oH2nlPmi+wfUfgUm+tim9X/zEV1MvqzomgT
oIWhoTSCEf8ZsKjS2DHRIdBNt59ofK+JyxooIjhodb6ItnC1kKQpEwYSSN8NBVxE
ck89jqoxUg9i33sm+u+JZiwsZJoezN9ni/jNzl76pJrWjsC9MiM+7HUr7JrPaPJr
J3QVaJA2hY9JbvEM/S0fBQMu8UoOnIjM0LXW5yNvTm/6nBf4QL8p2k/CYYj5Nt22
s9UyLPvpfJOD5piI6P2ET3x+sWfcgVKF2T/Qj/Js4P+KqFAUPNTX2RFy/VKdkTty
YHhdZnGzEsuH7iga6mEGPjbsnufWDlqgf5rZ7umIztl3plbMK5RGNRSErcZYkfDd
z302J8IYJWTVGrljV3qSKywTTZogeKr24PXBKQQJQB/ISINwPsR6bTZiPfWcqoV2
7q4EyEWH/TSWavQGGQr6PiHeRIxeRqgrsL6T5FWVY+LX/HkXM7FBtGJluWeX/izZ
hJLD2vbNCPDitsc6ZPV2yarv2nrxX49ZQQxLaRzqJynDbIYEB2wNT0QG7fsoKiit
V/iimw3jJcmghur2xBbWxKEBEafIaY/vtvrcWRFiZ9D0F/sJmfxYif0jUBXen1G7
vcZF3BBwoKkbWH46/IFBBKhuUVswJNimXjZ++TC3C5FT/QGFZGMB1MWnbK43O/nF
qKeJ7OuU1tZp13+AL3WrAWqnZLPrfBeYaEKFG8jFakZvGq8O7g+Jf37+3DpBfI7p
nRWrD4pS+FRAiBpsmM8MccjAiRI+YG9lyiJKNkZGzI1nUrtG3RYNspx3kMIE6SLW
oCiqFo8RFVnK520ndbtWvBEGm6P+Hgi5ZTCbIuNgkg/ZTk2RhJOQdL1lks6CGQNM
XSIkhHZV/fMukec99A0t+vQ78My9yoej6G3IuFPVzHE64c5yvj9zsTPyMiNwrmEL
Dm/NfXI6HAyjLAQ/1RFRt5df79401mIic3hkjhTO5+YqT4QRbllARKiJAw7NXFNV
vYQiY/CXXsgXmH0lELd0PzA73fJIZv0ZgvSOAXIK1E9CS5pUhDnSsQQxCkPeD6rI
Djg+603DvIMrkuEro4qUhJSqkg/pAZMu2Dto63ozxYOrDGh+DEmzGQRSvPB2S0TV
ouP0m/3xtMK2K9eRf+v7rgiu9akYVdagqh/5JMiyJsMleFwpu+mBIAnmrLTbsYtP
3rk5nszKcwJvl9OsepdWOancvIBlMQCb8ArNI63RnOHDXcoeatwypcciwmXhxEH5
MlHZe4sjInWJnt1bjnpMAsHkdZzo3q87LSSXYOkNIZxaihp4k6GvYxO0FbIXR4pH
MNOfjOH5RfaYOcY1Ziy/44TgoG2AgqWPbQPTQjILz3uF/d7LBJThNOnUr51EChns
0fYAM4dj5M5v7LG7B5pJVISs37H8HoBaGUQh8tKmDq/I4qcGd8cjQzQtAKl8+/P3
jNPU9DJlenkgvOTPigpg1yK9NpRcTtjD/OlQf4mBLONdBH8Mlfe/XynLKCQPuuD1
9D3W+3HGSSV4kFhNRtqPT0mT4L2ikg+PRX1zI6lohh92ARHxLKO4/EP8UaiLQu73
La1Pf4/7xy4mIcr/ptts5i64D8pbtOI3RAsdW/dSlIGcRnLtdnz+0n+f3hyDCwT3
Ba2WxMTLEaOdHV3Eq1Uu8YidBSA4TDHUw0rkdIoi4e6csnDkzmeCkuWMrFyP6BiG
s0/y5F3raARkfXdh7GzPQ9wIZ3hwla7G7J2SSxjewv5w3YSv2J2Zfi/skzRg6G8s
Nn2Ycb4kqL0qfXYSSD6VPh36IyWixKs79oX9OQZZsGjVlWWoV7tNb64+broSArq6
ADVR8ziFLapObiT8NmW3so3u4I2eAZvQqPs4OmGRyv1fpOxZCuwG4gmwMxO2VMU0
tJsQJHg6FZJYVO2CNu0QXMm+8XM5NStD67ST+1pG7nVsyB19fQoX7MpUC+uCKUzt
zPdl4o6AoGnneVZlIPPOaGJ8HfG3jpr6t2fHgcfLNUq/fhZQV5+M80/uOwza8ZcM
qwYNgCGM5wS9yuaPWBdOiHhGDVLrvzuEcRDKSsU4ymDXgXjunolHzsxFV/UXyKsL
rBv2UgTkJ7rxFwnriINJVB80VPcVWqzKEKhKJ6KKAcGIwoPtsEdajGKn9tNdt83z
q368f3iJmJQi7CLlMDWU3MV0HNhGbVrT99uFsqQPqnTTo964WTWsZEyIEEkJOxDc
IwXj1aPaBZQIjZpAccQns4EnEaVi+qhT4XQCYtURfKchsNo2yYlDc9vNI7u968zz
CFnlTRZMrI6pe8PqbYETjFO7KEc7m1XHzmYrocN9Y41D8ydGFkbEaSFERe8X31IU
FVJkbAiOXzdFEz5yCiMOY2VPB0CiEi8MiXVtbiIa7jwIduogFrSp3ipL85nhkQuF
h3JzydbsHQKPXdYKs5hMZ2PEUCQxIhifCEPgaX7cvgBhVRJRMXBdFqUtyGSEtlev
GLRmDbHo1NykvazJz3yt+98DddePqtkBU89o8UcsxGxeXnPN4RAly3ogNQtcHmP9
kHtGqydVRo0ko07sv5EJW4nasPHe03MMwlEMoxvkuJ8EWlUVfI2T5ynVh0BitFvS
1V1f3W9dstUpHbT+j5GlgC3sNBeFn9hqJIVv7VfgrLf/ivfQZC4kvoft6Lfy4tch
+bfdEDASROmfDZFuCiUG8vNfsA2BiOds0467dZU/Zvut9T7rFHWgEsrSmORzNAT0
s7J4sq0LM0aY5Qpoqy7AnUxmsI9OqfUWrxevkxUXGpXAJUWi0QgFnjSX5fJNp5Pv
N8YSvm9vZlwmCkh4JgpNZKKqKtdqtZ+IWBvTOS4VrK/uR4nQ2QYtE6UYlb/KUr72
C6e1z8rC18jLqwjyMMXUjoiY3RWHxIxfPHfy15GIFK0pF+duUr1Kyo9GZE6uj5JS
sEjxc/aNinVjoEPUxbACxthC0hf1/IAbeu5rILkoxwBC92aNJ70Qhv0ieIeza27l
F2vwVaZZWQmrcSUDh2Fj8lEvFpokI5OMhY5QVWufO0VzolcjVF/zwNpK4VwiK9Fd
r4g/79cRX7M8jvq/o/kJAd+uTd4067WNkZaPnYXDrSO8WKIzwG+nfLO3yg2/ZQTc
tq2Jgk350fw53+Pf23yEcBv6yhXTraCWYt2EOZJa+xgX9jV/Hvg5hokYkBoo2YKM
e7rs5wo3f0cYYEpMr4lQW1MyibKPh2mMNQ5K9HTdEXsj7a+1jTX8CvxWpaVTzHNj
6tlL9mQiSV31FJTVDRmnvKWU8jHnHQ8xrReGT9gjeNWWtASKiItvntCqIQNvB0wh
VLiybftzc3pIU02vTHojv24ryc1Toja8G0tA9kiMtlmDv7Du5cqboF+TCCNInqwz
+yb/K+IIWx9XLXOS+ADfqRl16baG3DAcwF96SwOtRBK8rDxfS04nDUlM8WfDz2ex
DtDnPdjb7Dr1elTJwzm7bZE2pIDt7xz5wzd7EY206frntpWGlkluFQg16/nUniEB
g1Pg/HfSDX9DCuPd8nFxZGc1Ylekk7x7KsflQ1VAQkvFU0yAHmtu8N3BD0wYFJ1O
oBIizymkADVYMy+mMuI0dq3cwcz3Vn7itdJ/5cs9QDBirbjKgoHcyxBmFy20HeCi
9wLOHJJe6GZSUorcXy/T6q6JmZNNmTQjhgTYeDZ1R6DHaQXhc+4GlmL6bYomn+0f
8YbKaiikstUtQJ5xKWugkXeFh6nx9CG1We7SHuq463l2i4jkw71dd54MBcAN2VvM
4jSpQdVct70YiqJe7BN0FrzM26lE4F/N4MmPr/0UcSOlHA753qDYF5A0DJVyTT1N
7EbbnTy5iWd+Vi9Dny7nLa6OWudyj7Md+rOL1YLclJW6hFBc8KSdkHvgx/vaB0wk
mNwdo3fCJUn10h34GUtGk2u0TUeEIRLPieuM9siTXp6AjOq/6GIkEVl1XBkCgiT6
P3npgnAvg9fX9CkvYmP3Ju61uXJRICZjsQISdE06FQtT0IZtVy9buqRDIb8mOWFt
JKTDggLZ4NtcA7NAQ5gbuFGquOcqxsKCbYTxD1yz6oaOQJbPyqKO3VdcgHe6epjv
flGBR4DavBXqCvugylGrpkfdVRw6RQzaw7nqKu3VCf4V2he/HY9ilNe9zJE/KMfo
bOojtnVhnpPywYs/gmbWIaUbl6TJkgruHSRicQ9WulatZOKl8hoJloti78m6U4X8
zEV6/8ip9nNuylKjpuHoJpq1bF7v9kJvdHjMYtxUN6Uc4PYOSi1fvwB7lX5JxWyF
6NPTpXAFgGtfzHeUmoBMak/RkC4/l2A20Vji21fkFuoRz4ug3Q0JWsPz+tzZdkmp
dy5cvHqQpzUabxHMX3r1Re1oWl3booMPNZ17l9ois9wmFltmO3QfAMs8iKZWwPYX
0m/Mwwfl44cbuecX3VaR+VANT0gm//anznAM+bhK7NhdS2832FW9jT5fB4T71lpM
rGsxgtX2bHH9wP47HkQpm5I9PEyl/PFp9Tp2y+gJgLqozUvNKz9YkorPMsvBb2/F
aniyEXSOaradlgbIevyDIHTufo0RU/bffMP5g2601isTpZQhsc4dr6JREN0nQC1x
HT6dDx35HFW6xDleoImPVPFfyusA/F7Wm6tqq5ZAdtKywaXc9z7/j+cF9BkJH0uc
sdsRogbnp34StrxGVDYXeyQ3ZPikGgCtt9A0rSto/C1ixrRBfClZ8d083iRQRSUj
EtTvmPcBipumOzxxf4Xgott6CWvpPR0KdgilQD7LpxyZMje091YDgwCFJerS315i
gMfztBWSnHj2DjiDlinhDFxaPvoYIuT87oH1KPISBeeYq4/9FTxWmTKLpN0fvEFo
2TMp//hzF/yun2vI0tArP83YDAD5+Dpj+kmZN3iPhb8rO9Hqaxz7JAxjYwKn9bg1
5zz9RSMMpbuzVjZU0HW0xsnv10mg7xwpXCrQkP59fBFtZihJaGT2KxfgDgOSYU/i
J0BUuyA1m2kFT0jxsUJl59GxykW/TyA5/Uzd+oTrzOFq2jgiS+oKF93z5hQ7n5Mb
ozK76d/AGjWMlu9oEraRG1S/CH0zUlh06PqlUY4ETzFnD5I5hAdHgqJ6/0w6LYA0
CxkM4FxdcKfFQtTGDdYHD7dHhQusev3SbeIp2JpgTA2GRXAVeHBTadhiCNWJP3I9
OL3aaFrdByLeCqhU9J/G+TnRQLobSWzSPQRCvCDVjq06pCx6TtW7xX29vBQr9aMk
YK9rPHDMn+jz+GE2+MB+4DgNZjBMaFuuT1GnMlbBCuamvG1oU8KEd1pmX/wGV3Pl
AOF3jRdlm6POLyFCewUiQaSJefiMh651Y+4JEGL/et1aM1VQ71S4IRVCjCPVaQk2
UHKuTOGxjF24QxAg036DGDpas+AqY4VQ6sm/zJr6jLhrXJsubVR89qA5XkFQaQug
3zBDivjIGqi77nukJjixBf82QE1Idl7cBrz220RxTrjQEHnRkBcimrDxKPfyRvtY
ReokDLJz7Ad8sQtYjwkC3iCCnNr4I6+D5zG9OKluMelKPGnNwHfnjJkPWztGBJye
w7aSdGi6QDVL7ExYgeHalUKbuSbZfENT788qmQxzpzU1qfJ2Z96ieEJERYXpaxHF
mIa6sslQmPf+GnlJmrTkPQbUtuxNYK9nLbWtVibONYHI+tWTZT2OBdLJd0Tqtz7l
g1or2D+ygul7ReGgtxBPDzhc4cFeB4krNYybSS7GWShdXg6A5vsE9uENT5/WdRRp
GLC/Bc3IsaO+rcJwDxrQL2/DhSs47RbinJ17GSLzHPn0AT6aK7Yy1R0JPMMOuNdg
O9mBp4mmZzOblIX+BncwMpBk1730xjLq1LvJp6IWrcm0fmce+w5CBnW+dYPaUTZI
YwRbGJUY2ZxSIroTFvwA3teoqsIiiW+fFGQZacLFTXrXqDqMmscg3kbtvmTfB6OL
qy4ZyEHm9T89j/gz1KtXbEHJ8d91/WdtNCMmh6qCMzW7z9vb2rXNnr/T5N+Xmw1J
VKjyVDH98OO2kwMP+QS4DSuJb4wk0qj6RkitirECm+m1wOfwT+V1MyP3BPtHHcwu
dl4PlqQMEpzyPvG2D0uaXDrz+tp89gcsVnaDMy7OPipvIYVA4lT+xGY0bRiAkdbl
SlaxlkkhFxdUkeZgEGDlvbAFQ+d2tromsQN6nkVDkSJ11oIH6BDGsuS6HGs8SxE/
rcir7CLvd4QqVfjOlijqVIeh/pO6MjleTMOXPVq0OwEY8XlgXHW6VjfjGlhvjp2e
VmQyb/DItKEaapqITqHfZgB3jpPo/u2WTzLIm9Ffp4GrspK6D6cz7NVZx7LJrEJk
+sBQT+t8PsibRsC9sxUe8fcrd+q4VnbC87OCitVHlcOioIT8sn9Ox3COlrKhiGww
IxB1Mfk6kMurqleaiqXqijK8eYpJUnhYGy2IltJuDAb9mSQ/E/hpHd2xzzPdlz+e
/j7xa312fBQ+hy3aPz33/dmKjw9b6sVQ17lP+UMyQ7+UzR1u0J5XKPisRV0Ne0TU
9tpoh/FpNMRNhPDY7HSWs9PubYblPruooQ8SBKQxK50S7sjM1bWLgEEBpG6oYbEC
U6AadaqalWXvJWCmjEfHyv5QfP7og/oEqXJf9TrdYJzhtT28R2GFlE1Rl1P96/Vd
Pxv5yjc4tfsR2YCTHzNdzJmPlkB/6dQGOi7Bhsiw3eokWhtJ9uJmaIe/FiKcXVjU
gG0aguEos7LxE2dKVuxO8RFlDo1N5KQNIoGksyW8cqR3dWD2MBZ/zs/DEBvZ8U+f
VP/ca0m7RZwKscKea7BDj9lJsJGm/RhaBX2eBfLteJ3HFvFJQ+XyAXQ7UtQcf9m6
EDqQ3qyH+MuCv/h6q/vUdNyU0GcsKbdKm62q774y61jBPLxx3Tszo70eGWga40v+
QWiIpdwQU1sDbsyyDrnrWNh1yfmllp4BktxfqRRBEfLX/wbSAh8kA/S5Ja3f0tDI
EO49v1ubNB/4YGUFPDUpedWE3gUJRPsXoBdW6dkwh9h1+oRw1xoS9DVkMznTMUUn
C+Uz5TkF4cHMO610uETby2/jmRRp9hw1WZ1w4GsE7vE=
`protect END_PROTECTED
