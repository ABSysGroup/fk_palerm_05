`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
msTHxm2TnvvUzvwU2GMSj6iDslKp61ABW9bP7/hoBUY5OfISj0xtW21Am8v5cDfY
KKHpaNU1B/r8qCIAqCYiwEpNrabIFFoKor3XdkQO4ZohMwM+xUccjSGHy1y+5YUW
uh3KGRYH2+IznoxlyuJ442YN4Tlq9UguzDrEIZ2evhfFy/lvIKWTLiBSw1nzYXWb
E60fEd7EZSAqvhAZZJGGjankObY0z9SFGWk8GHG+hjhPiX/FfgLWW1O+qS+/BGgh
ZaNn5U6wuQnti4Zf0FF+vC/PkaChxH9jeu20ilIS6AyOO0BqhSVfy3BVwkLEJ2qS
WJYq/Z3dzrtQeShSdEQspCAgeHLsB8y9DJb3m60Zx9/w7XtSDr02C3JGS2jfSAli
l8s4trtACt3IbwcsKbtqLYGyxoKOQyGWkIwVkkTqz0l4PLYm21CSSaswcgMAJUhI
`protect END_PROTECTED
