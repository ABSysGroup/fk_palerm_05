`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xaYFgk0tt+nIQGCcjWqg1EGIDsz4pwRNCQY+8gpe5DGcVBQ9qsTPDNsC3i4UmU8i
J0miA+ET8j2C1p3SbmozW0RC4/JI8gOvHp4Mfias9PqIv1VM5vJBMmqRnG2D0DsX
PwEoazMpntMOg372RUcjhkq+Yidksn29IJTOzJpDuExa0m3M8tGWqO3j7XEwCjek
dq2PsiAmiAWBlTf7p3RuHhlgfmnD2IlMR4fBornhnHQFyzmL0i9LZbp25bG42yd6
LnGwah8nFB1Ri63Ug4zwwtguKmH2oPNC9wXkcvGoiRXm2esr6WDJ9xgHNkON9aEK
9jzKhJpJ8wB6lzz7DXlZMQ==
`protect END_PROTECTED
