`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+4mtO/HDr9Ea5+OjsAPsw4yIKWqFgGp4PJUKNwdvhUkXfhUbnSDzHR7BsIr39zM3
FLgraYbcTPvTGAlKuuoWaZ8hN5z7S6jFaBGx+39/tvuDR9dIXJFygf/YtVX3vS0y
dtlmi7zQpiwSidScx1aOWMh2PfEkdMJLxPVnCwI/tyZjeuHRTeBOowPN/sUmus8n
5dhhFRDbPjfrVjj+ZedA+JGzeko/gJrwjZFYPEABXyLN94FnpJ+0OKe2g0b7ZAvb
/e9OQlers4XmENcZh6XLIBE1GQmY84sq5+l0YEfbYS/R35omrcDYe2HC9YCtjI1e
JzzBF+F7AZEoTWCR3/Gu92VPb546QQa44n5ZPXpdjHU4xNv7WaRn4GeKgEkAL+gb
6JrpfYHKnzJ9SR7xtUbtUiYnFx3SpiqpbN950ooUtVFTF1P02y+oP2WfJav8LO1P
lU6ipmonaPQcS5zHR9M2T8JAERXvB5bU5haF0T+wl+aSfpZM2Ex6FRof2WoibazN
OJE2pCaEO1rk2LKfbn50s+p1Jw/EemJ4q8zRR6+A9cdvrGqgxtBRpFpolim8XdLk
5nBEJBpE4rxFWeNKlalbk5otmUrBSdrGjfgnmc8bQmG6rXa7/Aq0y0/w7EXidH/E
mCm6kkAIrS0mg6CUnRjtKQ==
`protect END_PROTECTED
