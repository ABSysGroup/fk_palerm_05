`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y93iygiXlGJJDgFDwNSdMV0E0F2qfEMayGMxWtJ43jP7Gmimd2JEIc9EN5fZOqeG
87DfQhdZOW4KpDTaaR7SmiS9Je9LabRyvUWa07ZN9aOl2kPYwmmSWejkQXmX/Z1f
1zGEDVFsb8kEKJ/63UY2/L8HsQVa/mWt/+sVVXEBauUzgWgzyCya5kecNwXoVYmb
tl/L9aRqLv/wnjhJORt6wK9q+gCytI5httfDtV0CwTp+XNNLMQPHpoKejY64Ys3K
crxkXWBPvqBVFakhD08cmYUeVIBBEX66ox9M4fnOZkzFqzVk1ekF7ioT6YGwXKa7
KER2JX9q9BkF7n65UkVTHP7ZDqW5tiBfQetlcgyJ3jW3anC642d+FucVXgvsZCe0
xZWjW7ExvxWCnBWUPbgfR51ShKwidxj+UgQh43iUkB3bYZYZybejuboXoLzI+Hio
oV/ckv/PLhf8lWsalLxXuhz0H/K/SBKYE5pb62Bp2deZrAfJ+GnXGs5F6ehRQB/G
cVwauMeQp6Az5xwxnBltauFDOLmtAKJ5T/tTXfuYB/cZW1RxJtYEohb+G+ezlVBP
u0el4mvXD9HD5GoE75Os1l07zTFUk5M6poPBDbNryYWGQBGkuaAqisirL4SucaS7
4CupzkazKyPKwAMF2+xvZqqJyz7zIHybj0QIO2GiW50xY7qLoi8ibSsp2KJ1GYe4
kuFYDdI+2HEkk7zZ25uT5EU1CMcZO5cPDtnpv70QRH64m+Znmuw+8wRBsskf5b8o
og0o8P/MDQYJs3XeJj9atFHYaR2GcLdKuDniXOuaMfA5SqHfOKC3E0W+NoFrvax9
GxiqkrEOlyR7nwKYruFtoNsWWDKSpsohmO1cefQvMq1mxs1mwhuW9NsOCgTrtkCv
6OWXLLd3dYfZ5O2A71gmzrBRovRMu+dg0x8UmRhFcIjl9B6SpT5jV+IOklXiOezZ
`protect END_PROTECTED
