`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2JeX4AxgVaTx60xGNtrBkaBMm+qHpScu1dut7vGpQAKnq7aigR7O6Zahi7LdoCKt
50FnWcR0T10VBVzzOAKxniUfEPtvrPrIUv/RResKNYD+ejwyGZmazAmOah6MDImf
OPhXNiuPCib9RgVN6Kb4tc6YGR3gJBn+SXCN52DyT9LVwWE1WGlkxhVu9svqRjPT
SBvlLDFo5cqg9f3jvWKvVmYFzR0BMbmYMu7stTGu1fW0WCprWj2tFXDUVgHghP5c
93+hP5x1QWDE3xxL/oMrEAAepboCBkbV/p+m1LfcdM442/aWMK22WCf7fXb0N48k
lHflwxmLmA1T4ioZmyGp5g==
`protect END_PROTECTED
