`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fCEaa1uJqfd7QCOdSEUZl81M8tx/icK+CAE6DTHtkcIEn2UCXS/BLFW57VGwoa0+
NJ7qmvgN96LJNk8bMQWlMDE8gaDc3I3vxB+czwj033/o/GFAs9A1mRH9xGvzJ4Ll
WEWqzXGcVvYreEOWV4QiaSXz7iVepePBldeam6TqWn+iKQk/Rtyb+Q+DKieZjnBN
oflCdZzYdWVfB4EVyRzjyUQGpzuTQc0b6bbeYG4l9uYuCxuRpQM0LhXLXJqh2s0M
qRcwaB2J/LGAVjLqv2uy1ltZJlliDRdArtjs87xr1dFOL4uMVfKAg1CGjmfkauTl
k9I1TiEhaFToo7o8ZPhJAzeV8S4ogs1Ot7dIypFmhTsOgKvRvmTupg7J10Cg2dQY
oAmTi9ufcDmakA6LB7XymEvE3uAt7EWhgCKaDxQ4gXxbT3fdkITcElqDTDpMXVag
`protect END_PROTECTED
