`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PyuuQbT6Ugvfj/3t79KhIFjB5AlojS3D2QhA54HUxwGnVutMYBtr2vzMsSQprRCC
XLB0B+xZVtyE/9aq0pbJnP6xt4yuXR9BLAAfWscESJW7AknXe5m7RGtnJyJkYTOd
BibDfvqzKh46pXYpwign0ZDvAS5ioWennW/H2AECDQdtuer0KIs2gWU0vOcLl14M
Q4LCapFv41VRH2SJckVYAA2LiXZjNdfMGJQm6rzAbfhR1BCySWDuSkzQlNQPIuLK
nGiQPmj3gZnYfhu8+z4bvMHa3z6ZzBTpENC5gZQnbRidOGJGtLOV2y6DbGl16Esd
5zFAkaRHEAmgyzdVAeXjQsH3MlaQtTtm7VDLjYfsSjXgMeK14i6A78ygXarcqx5a
puUiPTVtdU4LE9haxOKHG+oQUxqoZfAlKwBmIncoH1Hc7cKSo9R6/2+uf+faDwE9
5+Lzaaq4dVfqrPZLX5sSTVK48zWZ2MBBKPzIUU/wjZ2kFUS6K+xoi+/8bE71xjNQ
oKR0gwIgCzr3W7ze6vhA/FGjVj5AH7iJqwKx8Qi5znrjPNpzUe9SSF3t+zpjLQYW
DfWsJ2o/RjH3mFVY7sNnkyrmawM/k2L+h6lG+63wl7WaAaMO34ggaJkuWv66b7F/
F+bxpwqViEy1XRqZUcfzA1HNicK8e1y5D07YIAUjBxzux+s2WVgoiL8DSaPciPK1
rxpkWYs6YHgthRr1aED0s+x7yKMI2PBEjuWQXXTy9r03zrcNp+zHsfhiUGuxUqQc
8Wnr6LvuBF6dA6iqepl9ZFArhEcgLM6/alsILpt/TiqQkYM3peIHiHfN1q7zsL+B
hZuovnMWGO0QtmbJivBYhThvChiHU5R+jY5d0bAJymEj1lFF+z3gcTsKCnHhL8ZB
4juEq4vZo/PcsHDO/Yo3uCD3a7XxA2GwewQRYeDyPfjyXJc+UrczRBTYiKB8i3Rk
ZWKXTPAd2uF0OTSygyxuaNPDwt2l/F4vwehyXtIg2QCszkY0gTrEH6jMfeBuLhhO
7dWE8YC5xN6vhy4eDB7w50tLl8IfaaBBecZrIa+WnlVc8I8wPJJoGWCCvmBzfqJA
6I01ojuTa435eBYE9Z64BlTbn2bugN8zm+VVDXSQFVZS86ICzGsiTsJP+Bw4oIPV
xnoQcAE+GrsA9nr9id9mgBpb1CbuH2fTZjw47SQZm59Wh5iO3GrZT4Y5xlyfNChU
qgrNz5QBl9xHbT3+jNRTWIOSPWH4yDUgTdU2ky1+E3fYgZBozk0aEmEEKMDO3VAx
uX/3E8ECvWPsCQw0CDD8k/2wT8UlTYe1dXbLLCzfNgGBHcvB/9F+5yjibE1XnXXO
03l/j5LJF2l7gwYwwAzIrHxjseyaPrJHefO+qttsdMsg//vHpAp9i1Ut8q9QPMtU
kjH18TmfHLPrrwUJDFLjxN6K/bsJHe7D/myX7W52I+f4cQ9nPaRFbeKlmOQWNuET
8a0OUOPc/29u3csgZPaFAjbYZB6r31/Lho6yI4K1F5UmVaSpFyiM5gczsPk+Lx5Y
Fdt4o/WSdHXloXZn+A5wIdSbUEf3JvhZix+r+choSQLdXeOaWf2vXap82r/KNY8W
X+vxJaiozwkVgXxtwC4eLeyXO8jOchr2JyV2r9I37aJIjm2adDa2ZrJmC3gk1Gja
Fm+H1h1bmCp7qh9HKEarR0YnGJUaNPEd3FCpFbnWbwhyP/jo9st02bBacyQgNjTo
DFCzsbRCAje8gsNkkHbQJV2oDdTNgBB/FNFb9+R6xhB3F83U/YhN3Mi+ANqm5P5l
waCtTRVWbrp2XvWmY5OGJx4R9KjdxCYEMNb0+vP+sqeaMb5kTSlTGXaaVSzrwpOm
3xZV992plClHlZzFcNNIgd/wg1FrwXCDiwBsR1/ZdwCr861JW34y6poJtrohFVgc
uk2cElEVWIBXBa1EA0PUyxPvLAQo2zxcaIDSTojZELiPomwnLuE+X+0ATRLzibNH
aaChakBKjaYxS6z2roukNgXvsloJNakM2vUHCLthn8m41Y7i1TQkmTjRv/jvRk4e
19BOpSUerirqwE41XKFzC29xcib2gyYRMfRDSjzqSuwh6Gves9dGlNbHkoYDJ8q4
oB+IdallgpxhbuEAlUKJ0KUGNo4lkDEJ6X7/kT2OTfzRM07GmhJ3nzzzgRyAnKJK
8ism4j+c4CftipmyyDVNuADp0WVbpnhEH7oE7OwLB+8yyxpuWSNlePja57l4wCYB
KRnjgUEfJsiCSwb7mohZcDImHPVqQhRq50CkQw82gpFx7ERgV4rOYmP3DC7zQN8T
+mEhgHeoV5QTIrhBDVAy0e7mPVugPkMAVY1GpPkrGnnyPYeZ5ifvcqtZqMlziZAH
wbXnjrRLi67+7lFA1NbAwm0dCTPfLCX9QFU0UKl2Ytyd1RFXHoRgyQaXM7oC5J+A
LB1oduWvWR41SxzgWuQKRlqhtv66Fwjm1kAKFJIdhmVedL/f8Ce8PMJtJXn9WH9p
/gtJ0TRHvOs80X9ttRCt8ehTD0sjlhT9LReaY1PjJh9wLa5u1HsbAVThT9D6ywqT
c6wjlhioAuzadwEZjM3oEuYBZOIt/fwOyQQuwsj1BgAckVTCctkaI93HXVwEjeUM
M6KG1sJecR99rlE33PqPc4wbYUsk2KIasdRNtuSmvjn0NSTuZ5S9b9GDrTVytZkr
9QqPi8gxVEIBp2jYy21gZqQYjqXoKtMiUduTe0Ft3/S2iSEU2f8FaCz3+V7TBWid
l1WsQdnz7suJUBezT53VPkrAwlcAtoyXlXOD5qpQ0apU1eJoFl3H/CB32yFSSh3j
GSAirDIQheBEt3jZ2U1BLA+Foza7BekWeQON2gIqndTVwIzXA9GYWsZKoLHBYR9J
cjMbDlJiopwY4DcYipEIQuGU5cEc2ynnYWIZKkW1AvJSWI1QiveVzZ309/ORluqn
eidmq4tOtcq8U9z1e8IyU6AP/UwCLk0X/b+An/fw0+UnrKxq6dVVQVUqDBEaPnDK
oRZwHhgUYuuNifvhwl4HEy286KpFKio72WiYeZufqOpJShB9k42aDMsBAUX1zK7Z
pSWAYt4p1XAxwIbBDXJByQ==
`protect END_PROTECTED
