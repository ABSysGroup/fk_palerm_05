`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WzTiTd3sdoI3tyyjxhUMr5qREmhnwDmPg7sibhvLuGgoRfos+Q2NLSSrfan1lN6Q
Y2kU/lChPlc78PAslhLjlQSQ9TkttjdPO2qPU0Po4/18bBRwfczqPONGOZAU3sfY
axANQCilkX6pAD8jL8Tq6KgqrFDGgKW3F9v0w8FpTSNqEZFUt5uyuuM1e8IdQMe0
QzdpaRYpvto+zcvfisESAEt9cfVc0rsSvndYuGRdBkk=
`protect END_PROTECTED
