`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V2/xj/bYC62UZ7CKKPxogPZsYP+ArAhfb1apSGNKvQEEZ3VuiIqql6Z0qBlQ3k8A
giAT39BNZ9tRTjcmfSWbkorqbcCwV5ZDBm6H5DucSiORJd3KfVsVfl7dqo5vElC7
3oVILn+wjWkK9HP/6FLOOMw/GTX3DXg8M7coMB1OSVzDLvlIINwXffYm9JiWioEw
SfDrTUX0vkZQTkQw0QVRaHMBE18w55LIEPy8ENzJYevQKdUewEBJ/8AOPTLNdpgV
`protect END_PROTECTED
