`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qLho28fN3I1bH1n696nzR+vYJLQokw6Fo0J0x/GQn1dvnkm5e6+lc9RDind5mGXO
khC2DkWQEKqAx6GjQEyvfCOm+o26t0as2twIW2a59N3pY1UZQmr1rtcJwOha734v
KavkCGG1a6oEirNc1r0FkloDg8kfxjNKULB5zpdQcee9R08Djw251mEfYQH+efqO
IBb/0zgrHApw+7odl8MdHXqZnL+C4LisGAsLjxdVwUQKvVP26eDg2XyJ/ZCYlx2J
cn3CqQBPbbUqikTuzW3skYJ1D4tUuCF+n2TU/lihTywP6zS4R+vXWssiyA8DXaqx
ExiFb0nkBoz3hl5ncbEFQdeNCtYrKsJhkdRy/kSKN855QnNOvwzMi0Tjwp9I9zDv
`protect END_PROTECTED
