`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JbhOn/8nX8T9ujKHDjxbKE2BTqlLT3FxRrm+/g4WQbYb+b0FfAavvpyFyqtY5gZL
WY0bM90mxkwRRUM8sPilc9MBj2yeHTCiqSCSDaLjolepDl4DnJOC07Bt/Yh/ThCA
dKiXMNRgSr5akG5uydG3/Zm0fFIwAvEKZS4O7M1NMZiP6T9+juDzqQJRdKztrnG1
yFS2rX0ErA9GtpnuYrTzp2+1oEf+5SvHRaQpP6eBypAKpgLfZI10SEPqjnObSA2n
/ucAZgVUXokJdfB+dmmvx3FvWUFxYRVjxOWwIm0jrfl6/dB4OEHlXE7SXb3GHJkP
TA6HWvJ7jw20iAGjGz5a4aynfAziqOjDX6Le5azjgQA=
`protect END_PROTECTED
