`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EI0bwzSWEwCQ18rK/kta2hGWA4aKYsE/CbYFYwYzozdNAvuimV/3bwi+6xQulGAZ
K2rxKajbpIhriS7gfqCiGfGPPC2qUHSKdLpeHOWUvwB9zf9mFgT1DYG8FgspVdYI
dU02VFrmYB13PARBd0V7AY8Kpab8zrzIxxVqMwHqVVU59N8ZZNgVPhut2QQPlFi/
K6mSZXdi6DCyXB7NIxNjhX4ovQ/PegPXTWVEA9CUsQIdR4DM8pMaBL8Qpl7SFu1z
Y4410V9tPZ+Mr+vd/jiQzZ6hqf6UTTW76t2uhmKLIFCyETh7Z5yBOGVtExrabaUG
qC7j3RT7vuwl7SwC46OpZMUFDNWw7Zm0GMYNHFWHNXq3nttW4OO8KoOV5EM3E/NG
7UzLaN1p93vF88RddH5aMiH0PCiUkNnEcLygaAcDmFQogupNWKLr0e7aw/WlEaJH
W++uH4khs3E8/TWSh88dLMQdSuD14HAYBQ84iu/eznGTmht48ghzDp64zxgbvA/r
lqw0ILgHzZXyc0hv7lxN/qjBeZbzdlkgErRc01OxAQedpae8mkF9+KFW5XmCJs1O
5Yn8saInfkN47sPWotDj5ra54r9Ojmj02tS8/rMbic5dsKTOWJVum4xyC4Yk63Tz
iNDvc2f1MGgNp5GlGbO8DZE4cxYFHwsZpefHeQXlth/ZXEPixCh3rgoYDeJ9MQeT
5L5p5cYZeE856mOri1IlYjvYI7Q0/LQ1GzRydJ6j1lMrY+Ql/oLpk2/wy+ft45Mr
NT0rAxQvnb9+rwBCzwfG1O3t/0zAKH0r3vAJgdkSOQX23x0Gb0JzQVpPUxNVYKMb
1mzQjKc2DtGSMcSiIHvYeYxvT1WwDQ4mS+v7R8xWn+9JtSoNAJ4YJOu+b4wGgJEY
WDl7LsYzhJyjK8w25u37wUExS3Xdg5qVS+Xq6QHOusn0PvF4tJwUdnVQDYenjq//
FDIL1BFMYicCuXZ6jWKPeZb6dVVFJReJh6cnvpqXCl9bmIZGOfGAryqMJ2q1pNbT
`protect END_PROTECTED
