`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gPeuBdk9+cfEHEUTPTlrm3kJCKUh6KQLM40GwvwVlXIrxQ8bp/jVW4mfiDRWVYZR
fUAWj49rgea2vzDqW3aiwS8k1vxwotngycVwrRU2CiuL2sV5+4/hCgf7X1mbJnWw
30KPaU7vwaaL7EY+3r1mQIJQUayLAFgb1RugPrnr2+Zi33cdyYvYdWmK+YKrxCqF
wOV/MjaVHuaTqaH4WOxMkHxRcRer+7ELfIDiKjOEdG6LxFtx2zMTosd2vUOqK3xH
zNyEHdRbLacGYiT6MmtJy5eesWf5taXyDNLK8S7beiHu+NpAndd+a5eTxhClaRaq
wMnE3TSTOJx+K5PknBqrqz4ngkKy6JwrYkiAm7dwv6gK72DY+XKxfb5EV2zRQ9g6
2U8diYKAsDXuXjS8+UlM3Vlm4VB2WDbOdyFNMtmibwlP5krCWra+zj/oMmY/kHVd
+Z8gmIdHOJPAw4CqV+MFT58jml/2IaOtAIgsjyOZCyBqj5pzslJqBxAHsFGXmTDr
1dG6mueJz0VLtXyqEsOdEE5gxX552Lo83C6f8AMdwARWqb5lwbe96xnMPwMFDJs1
GchmVHFb0DGHhRzYAtHXgz0eYb0XoMCWKWjppzqcwUYVXDBaXH5NSTbXMbuCws1+
EUWc92k6OF6wqfpjtBjurgjAAaA/MXEw1UMlR0e5WfE92L38GSOeGT5t69rTKrnV
/cT25YMMck6bv4Lzi7Unh1bfQaLgpTDpsvhYvfA8MgnzE/Z3j2n97esUs5dd6i+L
6hhMpZExnVRKIhRqaHMtNcQNKUV4+fRKD6mlA/q9ASrTQsXpcZp6svx2S+LP8DzA
et7I/cq8NhZ6ZFDejNLv1lEBBAISmx1RveQwoCCesEIhyNLc3o3usXmZwsOighAW
bdNh80FaYRp71Uyp3yl7siaJ2Axj+Xy7chsiuD3E7jcuA/9TeB3B9GS2vS8nmt2g
AzW1F1wxUi165ZEDlcPCrNBpwBaFNdgj+E86XE+QBbUohHD51Wy5Jyq/w1osQJmW
8vfsgvwW/Htp/3Jvro8CUpRaSHSR4OFyQCsFB9r2vkQPltIXO3XldW51Robr63jR
Pl8qneUBYDVVbl6K74IZDpe8fVxCHEj+0CbVxtXnDFs9QnVZnx+zRktntK8Tk3ZV
SzfgLOZeETPvTWSKIv2/kjqf9IGpQmwTHqVS6JjLHOqXxUCuNwjXwGmtY9/82crK
DLAUUkPWkjT4zL6F6hZDnTsNeRdHTvWgjhMFiU9kJvKBaSPiJhHB6roLFFh8LjEL
q6Bn9/9dzMF711oavZggIcttgMwAfVQo/MdERRQ08T2dBSo5h8InaCR9p6xEMta2
rbwvX7du1Yb4ulH11C2ahAYmh7WcnTRkdqvVvunlfixU5ZJlVOx2K4N+xmhxEfxi
ZjP1grjSpXLLOTfYvyEh4lYQXabHwtdJTGLxNaEN0pc=
`protect END_PROTECTED
