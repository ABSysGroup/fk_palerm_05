`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0W6ZBwrLbboR16m1Ae7arWxSlo0SrWsL8iupAkz22e54XKaqUainB854hE4tZJZs
ddkSeNTgCO1Vd7LQNvEJ0GDIj+Bpk4cYOqm+CogCi6kdDm6w1PqB3UjsNcbQ90jq
35cLWiWlzX6FYCo0dzr3HnR5gaGwPZyxwFoz4Nlt2e6+3QdUqTIrhrnVCsbppT5G
b+82hF/SKqVV/5LUfCPkFsFw0SDeNN7Ku+OPHWeAmk8FcccQ4/oZ0dQrkJWywdhq
GkS0aHAY6G5pClx1a+cZAgvGQvbcOoYFIrykhR76AgHf8ssX/6QvdVQ5ditemVQS
Wou7UqNULn5gzeVVEqJF8eUbbPwiMfaJdneE/7YikTEBwsy5r7OWPGrOwkRu1OiL
wLCQUrJhCy/rpaupqJsKW8ZViCCabXWa5qrRWkxlz+zGt+xXfgy2LqmAMwkkjn5y
PYPxbj67Ovik8lGvuM/O4YqM9Iq6IeysChVkmb9Kb3eepcrkyQTAW/3XUUm/AfP7
RsdTtxiOwe3sUYHA0Durvtv34EbvHi8hMFCZPxw3mrr1JtAnvtYhrlXACA+UsTQy
V1Ch3bYZLGxS9QR0Xi2yn2Vd29s++Gvr7uphNJGXwq0RBXU9uyzlToBoak304Vlq
AbSKZ7nOJMfd6okmQt/WWDkDKkuRDW7kjdTivMyLZeBdrZCN71BNMWBeixYfrGOV
mZf8m39RIY01IOY8g9Nq60mUKPtbz5EtGKroZ19dzbh2+vra0B7TIbJ1cuKVZPza
KJ8G8WUp7I+P0bNSj79McbUX3v1yiJ4hO2rmizKV910WmwuI8KAxwVbxwTN9P0+6
kkvX46SNUEAhdaTUT6Kyegr5JnC3zas1WogNNw9PBf0eBL0GlOFMbStM+tNA93Ba
b/+/7i6u5ILoVdFQu42ixG6HXA0U/cDiNJuklbD3+3MNobocbEeMatJVyJ7/M1Z3
7Lc6W78J8tDmWbm4Tr3V4cGplPSywALdiOQzGusquy+VnoCWTJmsMrTkqfWyAJ2n
gB/sf9TwNu6CS39RvZkfVEU2ecVaZhGITfPJjlve6zhf7J52ZAP2guaSv7xjSOVs
jB+/xo1UI4PdSwHyFQtcwfBDXEzLPYAkiSrXYyJXIfZCZOsMRFMlleAEG9RprxXL
rUGKO5HTJ6+yn5acrDIym4Ky6RDkUbUB2KeBSUeLpOlL7nzg2VWRJGtjfYGTJAf+
zKMGxHZD27yVHndcPx3EsK6cVxjkedI4Qs313M4NWa6hzwO+0lGAqWHlWu/gPRio
uZwNAf6xm+Tu1CQGvTmycRpGtOVc4f5ZTRhRK2t3RHjBIFQ5Sgo8n0xOTJ+XT2Ry
CvEBDJfgrH53Xn90u6r0eon56JYrYRmIYuPnAIfO1E6YIruxf3QD+sTpWkuhluHS
2VwK97MVVPtv37Z5VO3c1WWxIG/gb7HeVm7hUTeYNPXw47KdNesYbaApmTlWd7l1
D2LY2kfpJ6YY1ozMJbeFlYdLQtaxY844YfoiWFpZ6oQyOyjMj9WcC6hrJzEn6ZUX
Tb6bjdbgE0wyPJ+/G95wbxjntPTQN6q4aEZ4WFr9o9btRN6XmANx+Mf4rIKncrGS
WzrNiWDGnlUcBTzXVMe4SMDFxN38DfaUO67feJ5zreVuyw/EBxK+mKrvB8/r8EEE
k2Qezj3Ziu5S6YIqkqd0w0aL9woFHVd5nid8KDxJX4ft1qixh7DExT2MLedBb2sJ
b6Ff+zshmWZkuRXlQOsuMddD+Nu9TEkLfPkiqIJDLnJZILLwoY2QyZ7WmKG0WHaz
Ul4+c/Zllx4AbHr6vzgmHtIxSieA9m++sExVa+p3Q0OjcHdY18W24ID6LaI1EBB5
md8tgiMdrVLJmC+CDUj1XoieQS+7/vriFg2+XiWUn+a2pZGUDKbgz4ezFNDQjiY2
6p39IHzbnRxiHKjvj12ej5qxNH0kglhXHhXv0NVXBu3Uts3Xo60CN6FvDBX0ITVJ
EGkztSS+yh+qFe8oKsnI/46gTFWjeF7rGsv/DbbAeVq5L9qvFVPHyItcWRXQBwbj
8c+is5UMZ5og/qZ0OZqbpchrtZLVgy48ssBOrLpJHo0fnYhRzQ94BQHbjyAebtSD
UHjduzg+Pg7bCLHrYHHedcZG/u8K6rMVCmjZPePeA5GyrRVWPq1eiUXa+kVB7SEH
HW+096g+p1EzrEHgiBnozfGJH69zsLMsHatSZShjcjMzePuVcU1rxJ/tFBzZkToh
nybZbLtocmtEA2Ic0EDVjzn0YjwprYLUfLlN+hgEmgT07mFu6Lu8vrbtrBfuuaEV
E6TEh9b3D/idaE/pDcictBPaY5VmqpfEjwNafnCNGyC/lyM5CNkI6hLnDkbo2DUd
Pd56sVeGF0gWfdnkcgqkHRiOOKytgcIaaBAm81p2hxn9VR0EEvUaOAee5sN+m8N4
FtCV/DazTuwCl15COKb4RDa7DQNDB09FRplKPTYUvSbnB0BY6a4p/Be4HWSm0Sy0
V98B6ftuJRV1OuJq/JGZLAkmnen1WNCOkEm5yYOOpjjRpyIFYMRU8wz7aiGTp5nT
3lA8Md1aBXXox+bEgw+9M33EA2lEF8znOKDeY6rdX891GgTdd89vL5RmZudfFlXa
JKHYB7vu7oeTpvk0mhpUjKKrcUOCYdaCeXKU05Ploexob8owuInTA9dun2tVOQ51
U959xgXSiqnMbsQyHPx9f8nHNjluGOdmKZcQhsihEQY/rAzl4uekMb1RvIeOlieo
YM5NVafq0YDhpUZkX3eEeOhuop5TZap/ca+nzlm12CWRD5vxk9xHYwNHqwC3T5be
wgSSTCrMKPxuMwOuIk3r2K0YGDfhe8W+c2s5UM6CkwNgm0znmSqkwXnpyII4ubBg
lGwdCJK2ck8oKMJbRAHKt0icite9z5K37pfLHgquVhxzerZBaxn4ZGAiYPY/jVaA
f/fl5uOJuNGV0M2SUVpkMof3U5ngsF5o+e10eGBoWSq+1LL6On2DCjKKRMngKM5P
aOpVwm8fO2ykzhtxvGwXLvnSx979RPYAGI4d1Hpl3yX6jIpsaUEjHHaW0V5kFq9z
IOGRZjm1ylBb+CmsRJP6Wpquff3HB9IuOWrvyL/qD9lDJRom+gzOjTnOGmCRgEO/
Gol60kjoeo4PR5gLBxxylfhNkU4nw8Ax/OSOINeJfVWJ7A1nVwqROngLPvk8Gu/C
Fxg/sSYfHs9QvBPEX3X/z8mEA1yyWdpH3t/zUBWOI7Ae+mASQ4fb3rE/9SiKHSNc
Unok5mhVnhxeo139C2z3Dcoj3EFtia6butu5VhR4+2yxJsXkXVjiWL4/pIrJKvX6
oYw3HtZL59YS1dNvuFQsrupsB3S/aGEsHKMX0ryQXwTfH29nHsZaCPhJLebJVK76
7D7pr4Ta3eDZcDhrTTb1C/pxIQWSDdtZZXJQYBfiYr4FLrqacUTp0vN/bjALr/vc
0LBrOjddtPkaSkf5f6H6EX/feZ7hADZ9r3Qv8yMs8x/ILpTIZH7OkqqEbvvWWoIv
2tNDOOpjX9q2SEs46p2CwOBL/MtDXUxljNKBFjG0csIXtOsElwjKCMdBPnuYpLuv
M4AwjP63H/No0YEYnLatFzAnBywLIl/XtV8B4/kXgH6qoIs+2GRY3JINcA71Ru9g
wvwVRFJSLbI/uwo24o/64v4J6zZ5IQXfIjsPhwtjYnXJiPcfJfxAeZjqW7aOruHa
lFzdzGjXOuKGfLGw6KjAxq5TywgiutV4mVUEyPb71K8K592OtRVZJXS/iijz8Icp
f4Vr9e2jzL8ru7hQNarrGxrgJP93DVdnwiwAjYu78DEqZiJn4LD2Gen8trAty6yr
Rg23MEprjaU2onW7/hYfbamDfcs5p90EiyFvyi+csxseVIIXr3erireaZqYXhfbm
hU2TF0zHhoKyDAg6tLWclaqTbX/LuX1/NpdGxCRpI589yCIQlMxR9y5KR+D+LOxe
JbiazfhsR8WtwuJkEaxuSCvDCgkBTCgW96FwcyJL51FQ9WOc5180BGgSiKiwLRlk
IyNQvNw2Njyu97C+2Wq382ny+WTakfszQ8pfwwRS4YkBqSqHbiGQ3wldRQu3WgRG
elpiTsKZhgJEz3GmwiTPZA==
`protect END_PROTECTED
