`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3f04Dg5Kxnr/nDp4GXYuiSUIiUZHvRA+wKzkaKummg9Xxb8tA3zHuxQRzlk2SBFW
M7EyNsZ6uRf6YXIdWhpK9VyFB9liZPaoH6hirUPjysC9C9weaP8cX9jkF1M7L13P
50HohXA2f5/JUrXdkzdwBZAYkay1ks6jCmRNu27QiGTIZZTKJYy5+rCn+ZrTcLb0
nSPqq5w8nAw81pSUA3b+rAAxmPH2F8YmWK3Zsok4k9gQ1+VBU4mdX+TFPJn02ZT9
wrvAqIQFxsTAoWNUiUHjBhDkLBwjtkaAEgxIA+dxJC9rqSjMU43c94zxP5jGsMgM
7zIrlYPvbhG0Lwp2sNzF13xwUbAtJz8NTCpqtLrADd35Gu3tX7AVuFnmfo9KQ0uz
2VNmXeLMt9UWn3YA1zimM17Yd1q0Bj9J57vA4D5qQKpaGO63tz4XbDLUQ6l6ntmw
wgL0jNr2YvkXK/QDq6G0aGOj7stX9oJfWKU0WdhEkH50bpXSCnCiJpm8d/bwWlPk
QbMemqISdXKBLSa/VrjAdv8gzJGxcAujvochjYjrQF2ufXCIgrp0iX8MATOV+qac
F1sbrQuUyriUMNdVavodDgx0+dtL+18jrtCiNXR3AZA=
`protect END_PROTECTED
