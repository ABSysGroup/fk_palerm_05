`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fvsywfI6bnbXFoXm3M61hdRjjV+kVc1M/65rMAWdM1/FscBL5fa/cldcTFIW21RM
56U2OQZZ6HPNwsA+KSFCIagAnZMsGuuv7l5C8ivmGlBjnVwa2SHYcMS1ABDGav6r
D4ObPd9nY7sy6DrYUEO76fEjXLGkC/2tx3jFFLMxLfs0p96HtGwghB09YWcg+V6X
AkrXqFo4zC8k8K1ihAxyKIKc2JAtkRhaunUk7eNxfeUZLqDit4RtqALZpCVctQBv
j4+IzI1/INwmuH0Fmm1eJVIefqu7W4d5ZVNKBvSAic5mlWgHL1aYGIuGvHEhv4vC
NhL58KkiKHmTNgfJWY6STS4+Vkp2CRRo7sXAXxNk5d8GeKlp9GgsxfJDfLGwKV9N
cQL73XZBvWGf7VjP4woLT4DP6sEJza/itk0WwRz3ttGAs8gzB+ChlaOz70lHFHQp
Uc2jlH0QJr9QFtoaLFOEpBZCFRK/cFdNqSRuzTNoZq62WpsfKu1UiYf5w2PemsZS
wr6eEfvIEadHJzs2rGs5Pe4X5mlFiE7a5op7ZgNIHtJmdEXiUYJff2fI8NEOrdzE
s0GHoBhCOTfvc1BvBjSByeRKFUc7zrset8KATihEzFIoFpa00h/YU1UpPYgWWev7
5LPgwIMV9eX+ImPzE+FTHw3JpMY6QhiLN81BQB25BDu0cifAuEkTgN65w3BPTZvb
UzhH1skbjp2Kxdr2qO0axVslEqvMWadJGQB6YSlFnEraj/LivfH5qygIRNf50vEg
UXNxYm3MAEAw6o2lmN/BNh2kkwB4rXVpGw4bNMfTPqAvyBjwLI5R3n5FF3tnujMt
xt8PynJFa04/wDtDKz4ofb7xB68ZTqHjNg8UZ6JegKpZMB/Rfyo9xxyomvsP3PkH
lg2G2fldGPTcDvYdEzsfLIGZXDH9pbtiGdPi+OixcrTMNW/usHf4e46sfRpeMK8O
BB2BMUbu8qon4sYvusFEiXnZA9hbKiKPzesBA1fpM/n1dQNjsNv7D5W5TI/gKCn/
Acum7zFzm3aSGJizmy01EM5z1hAjIsfuP3KFnhOqc8ia3moQXITCf4I7qcJgrUnh
7VbzDdd1B5eB5BY+GjkdIghgFL69W/DtgKxnsI+OJT8hbWwwzl3BVYIdWNhw5vJG
OrpW1FLUwHM5YHiLkpDeoVXN26FZOv4PqMFcO/To7VrX0OxPf3mHLQX1Ly9C23jg
OlW84AVPoKypJV1f7UhkQ14flMTuqDgsi5tlcCQ7kKOabT1jPtLLZBlHDPndyikV
UIOsJQwut6IPvVMI4vEKEDxqmruM4i702Tk6NE53CRhDFPofX5JUTOeNi7X4DsIn
obd7OVKl4mUDomEX/2tRiDbtPsoW40ux3L9X3IeaOLvlH2div+dXrMI4/jKgAViT
QaS58iyNJKfkkfbqEJ+qboZyqj4dzrx4Xs/Mp5GtMGC2Yy3EJCNUXNhcux3yLsx1
GmBlo4I3ImUXLB0eKtij4Q8L1JsRNkWCZA86jqLznfQCTvN3krdbgfq9Idi5kMGQ
rF9pZekKj84JZb5ih1+/UvmJbBn7twYA+5PEx4/OYwbsZkdRMyZoA6Q9uyIYOzAg
G3apbh63bZeqC5UzrZeWAG9hSdSuZjU4m+bGFJZFPD1WVQy4oZitI2znzFwrsNl2
mo+qZX4D70F4n7ry0CrCzcp0nHFU9gK/4MGBZMAjTO3Xp//EdZ6VZaf5SOJDO4NH
d2MeeICUJi/7QlKmEgtnZJy73YeFShUAc2omxHsouUK754aEOt8Rd1t/798MOrwT
DwMCd8t/C1iCWXui17UmdpJ2YbOj5YKHUxqYQu+fT8v7JwwaGfMJ2Utru1hWjE+S
B7nZJryu6L4F4DPIYhrSTj4CHYVDiZusgQuGEFiyyZypzjSh96ZIqUjCx05JEmeY
iZaJ1WvZWOavbQta0BFm8aja52swPQodE/NoNJ6Z9zVd/cer7I6pppboKtScoNyg
pqhP+5Ywedjr/jNhGKEuE57yHdNxwl8v4nmnW2x3BHpIzaHzizQgOzLInoBGma5e
SD1Q20z8Z6O4rRqaOq82ps/xr+YcB9i9q5WVB+PzfNf7AzhHAgnBCeEK1jMkHZq5
WtUEBtGkEl2+30HqmJaxX++g5RSCTKczpjD+bZDw4xaOtdMHuR/4meSnUwdemS6Z
VmH1j3qjlqMEznr+eMSHdpNoeOL901H/8cDgNzORYYNOpO86R82F6MPhpGW8z3TF
JZ2JUxuX8qsbw0I8s3Q5LC27MhjB764FFRMzGgyo6LwmT9P87+izgI5gJvwEuV8v
Yxz2mRjKuzvGHcwxY2wUY7L66gL+ULHnTRJ/f4F6yREnMegx31YJo0aC7HIUo2bE
OvHOZB1d4W/tBeCam9g/ANaJDQRYyCY9D+PhPeWIR+ZeStTfmeyNoITE/Dmg16Lt
l8WwBHehlFAc/86V+tvJy3FUCis3nJk3qnJF/sdqHTo4PvBUmmRj8BKuuWG5YURo
q14YhhZszEagOAhMsMkMVGlM9CZukXXSTOd4b0dj0Vt0TAXKCT8D02YXSUvmpgiw
HZNhq5xZhE/I4jnIDuyVSnBrsvT9V1daKZr8slIKDI08VOvs33T+GWrTrRlpRYM9
tEJncH4huyTMqy4THJ1Bp+YZ13rolfeU74DFEnT42I5MzAEsZkT0GmLl0hlqOT1u
0KfXCEAt0BqdWfbRJvxJBTJGwpGqBJGBreuL/ffZ1PGTQEZC3eyw1zrFUMuAXVJW
roz5x4da+4HjWY61QI82ktXFygShO8wOsjfpWbuKkp0jS7hgjLAVnBDrO6886vtS
NYzIkzKFbQrkBcQNiI1AdNkDL3JMKKu7D+jsTwpKRQfXX7uGKbttEdh6UjsrFy6U
5K0AtwG01cVw2F1eiCdNf+1bhVk055owcO49Z5YpX2d2N/tONsY4el5XFnaPEJcw
BqWGJRsyL9jYnTUaVAIioCmqLCy97HuUMuAdYz1TqzMR8hSSOjsYas04Cl1HXPdI
XuPt+GDYY5mscWSgq3QFo+37FNycb4JQ8DwRJno45hazvgBTwRfEUMSYgJnC5lmJ
I4hccPTQSlXZzScjHQaebZAti3+wHTIgw5EVYmTCEb1u4pLNbsKkHX/d1L8zHvGR
VavE9FL7zsQRTdR7JA2SrhBNnZzl0gPt5qx6u8AHAjoEe+Zy8C7rS/cmjnquO8QE
bo3hmv0McSZjy5QN0jBUp28u6dV2l93pr2dSDwLhdUbIX4nTrGfUXWrdh7+C81Rf
a2eJRmlXvJ2jqX5FNl1J7Qvlcp1Yb/+tqEwzu/fFcqC9o5I4ruQWj9AuKYfcGllM
9nHdRzt7KEwVYMgYSle617E9ZZ9Y9Z7CAIF7AeMlaP0yCYBQIjs3MKWuninmAEiN
mmbQ5iHuthLhi8FPDW/96PIXY+t4ibLh61tsItq0ZlT6hTfsQKjxUSKtYLuXA4rR
uElYT7bLjtsmhepEZjiMLy6Mg+VhUHI/Ba9rppsUnlIzZ+2+kol42Zm1WJ8U63xW
zfFGeufCKtECb7Z90xSkrMvRxJgiykVh4SizhNB8RDiahF+qCDVncFvTH+GRw8DQ
en5pIVA2B0jIOTCSL4FgYcmGzKx0fMNdXfJ6sWS/u9xtwDKZ3pjS3rv3FQmPaXG/
MNX43luSNgEvdw+aztkyLDIzGlll5VqD1D9TRm49JABNwx4XSdsEwb3cQaOW3euZ
MB9E67+j3MBZgWz+yR1po8oOrjy45LLetsOKl+QmVCzcTdeauCn2oXNYtTcfItZY
EXJC8/lddNzNlCszbXjMdIjU4KZMP8/odriUP1UBjh0ihlN+sa/GzYcbbtvzhDO+
0bWoaYa2iaHtCDVN5H1wZ78PIsxDc0oEYRU3KKv93uVZSSlVwiJhjfnKDJFu2ukM
Sdf328vTMPTSd+lgtMJbhEnCzgZmefOz9iO7K9Rg4LeutXe28y3QLNDaXy60MSw7
FH3K3uNA2p3b7DJt9ZtIkhSwdbhANhV5WrPa1y4OraW1q7QdBvmiELxP9EIRLcHV
`protect END_PROTECTED
