`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SOYPrrn1Us8YsWLSyJYyBImMgg5T9ttyKf7skn5jeMN/MMhVIUBkbGUjhzXZIo1Z
NR8+yVZzAF0BeM//H0GLh5dj311aa1J3CjRs0pZ9ySq6gzkDSUBwgl4OmK2LDcH0
M67eyojXAVOGSxjwjHwbdgIqGS7Td7+GmOguxZYCkhFLFK4RZ4E22Z1FbxgtRZC+
/BBF0GgjbHzpmOFTmwulsgq6V2NRG9MkaGhzkgpxlLMmh70SM7rHd93wYMqVdsqc
A7qmAYhUc5nfFc7XV2YmGw==
`protect END_PROTECTED
