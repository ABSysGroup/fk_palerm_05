`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BZ+czgW6tp0aAz3XLV8dLIXQYDoVnWUd+JYGtwmifHguLbc906tITuGwvcWUdDDI
/85NJMmfIHgd1T9YJIP9xz3DEJzR/0fRsT1Scz63GVpaDWzIWUTw8RpHhh8OZWz3
01Xqk9MJVuculgcKJ0HlroDkI6xA0qGSG/nIRKEaSc2Uf6WeLoUVQtU3joA+jgav
QawW/mp1Zzg2n3AxacND+ef5Oyz902YgmWz5bdobs+3PAhSf4urWsAoy3yVMDH9R
ZwzosPymT9dm7SeqmgJV+9UhGIcdYe7HNrAujUbyrA6XECTisri2P3D9f+5tNCYy
a4f4M84Lc/JaL+eiU1W8AcKaD1MdZGDvaNWmgAet+AyV6SuP+t9P5OHKB0ONnGQf
GIpB0dDva4cMoEt8qu1Tmb2qyT21XxwPbl4Elidpa9+yvPRd9sRyckMk7DsdN/dD
m7jbNZyDYEq+xdOixTa13XaaxEcdxLtSrEJBAbow4lvHXke2DKD5zR1fy8qmnUoJ
NeGfUdtugZ9+GAAwc+fvDWqdy0sde2sINv/gTwqfdBlH7Fb/kw17osjEuIyYL2yu
NaTn3P2NlIzVMomLZcBQRJNJcQmBPSEeYDXkeK7e5A9/ADQbJ3FvtitXv+al/+/z
hUsdlAqlxpFYtfIRR16jMkgivpQZA4UdwMvzmhYiRNnPLmNz93NiuYoCepNqaNbr
2iLUIEUHcfRxSnbxLPiQZuwEcHHGAd2hFh+IdhbOXTD5DGD0F5c6a6XCZMHvYwXZ
UnCoo1LAcd8dHUAuq5iPxZ3/QsmlpF3efZ6ao9czLX7jlB6hca3KYTUJ28VmMkZo
E3x+A2cRxXOa/h4niZl29kz1El9WHIKjbaS1w2KfoZnJqbwcUati5M45h13GYGq9
qOkUiFZW7UOY/LiUN7Ek46FjnSesGlMoyy0zbPyngnxbGdKW0syJJMb8kwv/Lngn
/PcUdF497WbRIsuYdmWEiU7N77XkvQ3KEItcWue0f3ZnczGbs/zl8BQVH3CHjc1q
JkQtLg7+VvWT/ly6ohnwuuh5uCyy6mD5vkOIDTvvrkCPSb+SmWKWZqh/xelR+Xxm
BtLFqi83Njz1oBDYrj1hTYf1jse3VjT19wT9c8xZhjNJ3bdOJN59BE2QRQO5YBTS
Jc540hzdNSXzpY+g7xo4r5N4o+hK3B9DddZ2OlyuC8Jfj316BLB1qMIma5WnBhjI
ViSCsuo9DpZQwwLJtBElHorkmMe+NcPaQmJWm8B/VsL3RZGMvvUoKg/k7zEQf9qC
HkJjPpEHLFTDyn3e32kDZhkdV5dL/hdEL5E6oHynWM20KFpaf9yCxoFAGlJDfV/A
mF2PVdBAnao8kgAKvFTs1p7YG1wtQ9Mzz+LEJtSpKVyYuOx2+HqJ2rnr/2nx6zrv
gcinY0HhZ7nEu2LhmbmvaRri6NJ/0aNfcQ8/2XFxSnkx8Kp96Yaozhdo//GFC5a4
QJoSdYZujJQ2Wh8a6HrDiHcY7yFYGFc1XRzRrudwmbaH3pnXEPUYbrYMTtZ/FJCa
6D1A3SARfIqDX6yR3/f0UwBobyMno1RUqr9SDdRozLolf7V1IFjJcPEcAxZPajOm
GovDtX78DOasMemT2s09OPuEMwrTOmt44xYfiFbQ4l8z7MXt0xWB4KvUIkFn8zeI
Dl7zH7zG7XLzU1WDpNAVPlPm4C5d3bavbR9rLzPUmJCrc2/Dnj2RzvRPkFTOlb0V
lYGlNzjdPtMUFbNLSK09L5ZdDe/xsnENoG+xDgCMdIzYbM5/n65N5R+owiXroOma
ldtBPxVuXSj7LZDRwfUtiwROI3P46ElPy1DUD8dN5aFgf9SXVM4yuipX16thg7Jc
ADWR57j9VFbzwSVpFy6gMUthgV+exjZaRQxL15CpIe39drleBvEz0Z+IB758hG3J
GpqzL5V8OneUrS+awEDTVjqUmgXFmemxTEC3caCpgT/A3eUGHI4AOOCrvdexE6oo
SR94oE9jqq8RJiERTJu6yfIhWizGTH+/f7UtCC6PjtNsw9VawY6pqWtx4EdMs2+4
2WaolLdBGaR7V9ygWU8OU4/Gou4a3Ko6IooaZx3bnyNa+uzf5/ZVxqN6zvRJGxPZ
QulRqEpH1mN2PN0JbCpGDmhqi2v5GfOgINNyxrf5YMcx7p/29MY2aoZeiyAIMyFQ
J4LPiR6DT4YVQC/P/VkI6NYEJX6i0wHQiYr7DQZDAVC381Z7GgP44scvUlMYUOo+
N2Q8FKLEku2XpEqT+M3HYGqXubmG9xg0fNF6FEUZ5Xe681FzOrTIRQhlifuc68kH
CIBbFJ00cvvTiriG/Ioxo7Dr+YAlziuckp/Bt0wvXLlcEbltqd5KT/AGUY3RaW/f
P8Uq8d1ask3vBn9ORqzK4al5WosVqL8bxnES26Er459BbUxqnaE8X0vtuzBCPZdE
zUk+8WTMrMuR+sm7/IImehjVGr1sKOytRibFO/VXbJf0Z2bPtTI57Bf+tHzzmyNJ
cnWci/MFGG8/hah+U58vvdAyaPu0SO8QgMbsZxtqYViZOSc0l2iCkP1dhP01s8oA
dieLrEpWUlPqhZ7khG974T1NGm8y31dJrHvfVogvXDnWZqAHi6aW3aVVF8uvtdrP
PTtZ6v8iB/qX6Yh5M/E7jFdo5HMvmzsxUBQlkazWFul42HeknXuZlPJ6vpaiVFJX
LCaNkcGrcc0IZ0ri5EJQBLay9ZuzEEEil80RO1/0ub4kP1V7DbmQgatRKHUgx2eZ
o/ldwAjUYiTvAh2d51vOMpARvtQvaprj7vVCy7xytTghjA1lx1263vE9grfIlPMh
7zJpYpncPHxtan/75mnf3GR/6bSt83kPKPClxIVBafBIFz4clxRd7Sg3tsI7cygs
ZC34PUBJV/zAo1IXBsxPJVl0UT+nKv+QQLp5lWFquS8cOU55F9bFgSrkYbOKPFkb
3PgPZzLZ2d/9bYzDtxT61S55gkc2BktheKKLZ3Dz+dDcS5ublF28GX/QgPxJDM+I
ujtmSH9ykfpcAT9eX3np6oTRdaloRoync8Ok4PMtRL+nDgx9sWbOIwWlcc2GCm/k
FtYCnoh9gs6enF1hYNka7WQkOk5wnAsQSn4UN1uMsmp+iVMRXsr8x8YaQ1bDUs3A
qErveyf+QLmqPCzidIahOOMjRHkuZsdoUTq4rRABcnfhrSNq4Pvaq5qoVfdLOp99
O0Oaak0RcZ1CjkN3X3Af1SDPzhmR6JR/uj520c03dfwf7/GPk/EOKfTfNy3cCVX9
MPIPV4Fb8JXBpqwjeu8pKcqEOFgF1sYSONCMieQ8L3uIsE1Dy1sWrx+f4q9uWXnh
kWLPNqTFaDnP6rMQi5w3ke7Lf25wz2QIivyA2alJnU/hrvq/wq5HtSTyhJ76kV9x
dKT4gOiRjMqfb4ClXyWE6XVaKVJjQhnuoog1CHfCsZDgb1craP8hzliBykyufaSR
O11tlf8HNO7NWipvrCfCbJ8DAxw2JAfiW96fu8q4+pRdKBRi2lDBugv/M07H1x9z
QCfzeXx+vsko53Y7wuQYMNMKAvSVCQ3EHVq9WOkN2/soE6kk7rcwnFvhOiV65HAY
1KJpn0445CUPhkUSoi/iws2c2z9X+DhhnJj2cMUVnrjG0RgUEBvKIi+AdCzTG99Y
VXxKV4P/MVH5tc+PUbx3NZLoxbwV8whcUg9BnTJytC1DBGKt3c8xy1LTYOyizgI3
i3xqYfNbIeEL9CIH6eM/18HdXJ5F7wmpk4aRs5jx7oSVa4bczL6HciLLS43IX27Z
iD1yexEpmuCHdN0VdbUqimiFMhBa9OxqqBOdf9hFHz3Bzudwj04fEP0Gfl+pY2lI
3taEvtYsjfJSXK9bFHwYv4Z4KiNWsVfUNkjmjvaODeTIQA78Q90Y12Y7Db5+9fsl
tZo+5Db9q/STa0Zr4GF7w7shVAywoAHNnBCZTPoFAXW6oNN2KU7V/xCtcgDz8V52
cNxgRovL6xMYzazo1ox/GzEuDTFJPS+MpL/h8CEjoNBJ5Q41tInY3WvgD8VWoYk5
1G1EaeXOjHfjAynu+H+j2yf1/xAaz9s8g4CoUWVCkyIHZq/iSU3cyW8SKPlTydea
cmPdONLucAGjmVAVSzhlFVtbbpCdR82eit/NiN6iAN19B5UjmKpqA8TjAO9Kjdt5
gKurS7RfReGoaXaYHb7XURmVXCdrEjxRanuFp7f40ansXXcpwq8y9qiJOB8o1yF2
H3Jq7U7g6Rd1t4fJqfXGdVfo2iXGRvZ88cKKc5GMPT7ULGrq/uf4AuEdXScRgTab
2SzwF4G3smCwY92TsrimusVviOeCFe7MbM8ssdQuhcaCHHI8f2JYxXDyZCc0MXlQ
KdXe0B+4tLWpnw0lZctpR5oZkHBWhyy5LQLuiwwN5EZfNbjCMKBSEtMuJx6pGJo0
xTysfsWwGZC+1w/mZrV1wcLkVO7XeTxcGYJtK2yH/I5mejjb7lTHe2o5tvq9AMIz
RKKELDzod+lytloqlcbga5aaMUBKJWTTS6LQ8aHerZSZJFxxP++MSgFiBPouLJBa
W4SAhgSisNqc16dB7moFFUxCpFtNLMfRIcm/uaNxklqwkdWBw9SMdW4G0rnIiEXa
BqvCkYe3lYDzv02+emj6qbdMI2CIofFG78qKaGhWSNmEJEmGFwVDrp1I4gA53F4B
Fs8oEjb3+FjTkXx9AcYYpKb9rtN02thVS3vK1DG7O1FtHa+0w721Jktf80M8HVwe
RYaaVbvhBPBEEpeXDGPk19iponZE6Kdhqx4aWaU79PWaBNAyfp6PvvytsM/Y2vOa
XNsILwTc0BCR0vic861S9SZsLAcPq05gLZmcZZ7cvJpsQhi4BJJoy84gbyFnpJah
PXJwRXe04dlLxmxb5gGcEA+ZZtSGLsQVJSd/60vdAiOdk8Lr1SWyclTLQBgO44oO
kwk33VdmnafeyQawCFkqX2zAVPQ2M8V7NlOVTp+JUDS24wK91qtJCr76SqDuACGB
8n9NHT1zrwvSGvEbl7psVpqa84KzL7Da1z6wyJKm1w6PVPqDwDaFli2BqIcl9cO/
v+X8x9hVZTEDe0L1+t7367H3fK2v9kdq59R/Czk7Nxs47UVJl1gYVrPkLcasbVgH
MtWEtFeqccu6W5yaBSk67BiXMZVPvl7E5cbyOhi8USxqinhelTdl+6EI/ZEEZ+qO
OIZ2QKplVcJvu9J0LM54qBXqJItq1pivVi7EBkrPOk/atYIPdH/n2LN92I5SafFH
LYGfyy7AVqaNohyh9JoV0+2CHfHNhPvbteVTmBEcvAzBxGKOBsKtjYC5V3J8oA2f
E/gFiHxYagf11Y7qk3wl6oCvxRZhuIfLkHm7kAxZmDnMiUUDtsLNQL1Kiw4giQJF
n1UNuxAfx50EIcwLHs2vjgiqWk7w8QeTXKSTHOjrZulvskt2sTBrbB/k1TVwZhBN
PJbBDkBGPtHkqMBjeyBwYDjl2Dw+Jy/+vE9APMMk70b9nJF+IuGY7bETslarvxvF
PvnuoMY5NVzzb/k9s18Sr9BhlbVO2WX/BjN+/Sd3I8upfgG3m8unvTj/7jZURqQA
drlmFaJOKRcenBJDXSq02e5IrAJFKyeBhDtBV+uh15KpMssqMrbBCS/mUm/ra4S8
CAfGZHRy/jYk0RclkBI8fw1+o5JHxuOW3JhibjGJpEOIPgPfcMicCsRHmgD+mMh9
oC332NhIAnLIosX7O7Ko0zl49JkRUJY0tMKMyinv2xvVHp1U5IHAPmoh6GymG+eR
aeK4PnA+qWM9SiLBDvRQ4A9dk9GZPH763wZHr+f08cwthiwms9AMAURmTUi1LVYH
vnKquRYgEaKmKc0S4BswZgXzYMuxvklGMiZ1qJWbeERBLJrtVQ0IsXRefBHQzLZC
xtJg9PpUc00HyHULv3Z0xS/1AToW6L1sl2YTHrgb7sB9kV/d5B7Hk32Rv7B/b3RN
5YF24KZlF/em5n7kTYI9hXmoqMl6H1zz87ZcvVjx+8OeJrjClCbaU8JBioXKIsEr
GZdQQrJ6iNl5eSNBaWTYtU2K1MN7wSbd0LKans7vL9/Jzv0J9SUemVNbxgX4V85G
BARh+TZqgdOhW78+wg+WOYJATWWPEyUftrhJLq1+wt0xfe9LaZH8XbeYSZI7VbIR
QhxQTqBVWQSzApBM4JF5geSm0lRsm2QgNI7+5g8AEgSeNcoyaKcQDEOfAS54/8o4
ei4B9GcScqyA3RXNztYaOSO6TsZHnsBwPZJTcx9k53BL3CuX0FLXvlCk4/dG0PbG
b5dkIaVeDYXr4Pwgzl4vKnRAC+71/t3ZkkF94yw1v7URmuRA2zzz+06Eoo04xAdJ
41Vv6s5Nj6FQoXS8/6JaYtQ6aH/hvSZHYgk+zer6QvLNLRlfumhAfyNPuE83mZg9
5tMv57rvfvOEDj2yNUID9A==
`protect END_PROTECTED
