`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fiyiG2uSleRQk5MukfRsqNYanpOgQD2aPrdKY9FVJxt1jISQjbA4rq1cFROimhMl
Uq5gOTskMUm9/sGjQZ0MfiHwzDsKff0K+rL1e9QZyG2XpaAWIJh1cJhWgar8C58E
BtM+im22VXHD/CF34ekP/9Y3xZAhwfwfcfNcrcEHliNf84eNJmDiGujFtGY4SJex
imdbsAmsSxT/+GVOd2n7w1Lp03cpX/R+MGw2swClGpCpK7EajI/VHHo7aac4ezGv
VFvkiOwq210CdkbpKcW53WzsKmcAG17Uu2VF8VKGaRBZau/3ncLULNYAiaH8dqB6
CuhdFwnnuyd5DkEbNYorcQM0aYJ94hn0+gHgDSM25p7Q+rZGq6X8CJuIJnx13Yay
Hg3U9x3b7mmgYcfywAowdCgV8OYshX3oXdupPLD4zPlqvaegoFZywWnukp2TRtCk
M1anJ8e4m6TDo6/T67DebVwqEFinO33SOVYqHpSLITUvAgNKLAkG73b1EgK4xyPl
d4MTJm4K5hFAowNV13vMYuFijeQzkwFBujuvffgvdcP5HFeH5p/OhFTRAalZ8k88
`protect END_PROTECTED
