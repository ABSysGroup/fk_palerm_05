`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VRE7DRyQomQJLuTbVe9A9WU9C7Y62P6OfQLvXxWD2jDUm2Wpw5XOfPEDTvoadPsO
VcfdhmcfE9/QDkxaOhldGS+WBBf2oQIrL3/wjsn7aq8uBLH8rP1CBqnuyqWGe1T7
WntrYBm0wAlMu3vPce5cQ3op45HEwH0uaauLSLuWx4Ztrm0CN4RCubIl5pQbnIkq
eyQ6k0jNYLh9esxJjtK4kIpkwUT47sK3mgSEnF0bjbGmxVtpT8a59cbOO9X9DVIn
wILktK8kKiRdK+8I5uLt5oYdR3NstBzIphXZJfVk9X/D8yKyHKdi0CU45LQcJBvp
O5JZ6eSHFIqe93a/OOSi2ES28t5GeLm/mM28IxGDUUvtWRIn6xKb+lTHu6O/pwt8
tav9yix+I3TVoAZz0y5fpW4eTugKXkibiey/d5jYVQ3ah34BdLa6PQEK74tLM98A
zBJ8K3NVToHgbKyMrY2rA9Ws03X9SIJPwtqcGqqNBI7W9N3k/hlimgB0dF3OKD0j
Ba18xLVjxmWweILjhj0WCfTMNhOGfYEi2LdLVveH9cwQY3msCOIsV64ee56KoPjW
ZGhE1X55IBGCmND19j6hc2nIzA0sWC9uSubgR/FlNcE=
`protect END_PROTECTED
