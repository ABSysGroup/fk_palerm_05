`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lB0kGfbbVZsEPzeyh3PL6VeC44BlRczMxtFxtEU4Nx5tLCuJ3dDndiBWvdgMo0yN
ioqZignxDYG9zByOG6EqiI3+01REaHEAXhkew4txUC7zZ0GVFSA6SOIFk51MIkbB
GNUeQZJsNV2w2/rbYmhODbl6lKD7TOtrMh0V6VR5yUyv1Vzi7MInPveQz7F7iQXf
Gt06TDPmvDCxXhV/SW08awuOdBo+PPuskRqmoq1oNYD1zmLOfJzeqqzux34kmjZH
HlZREddqoA2GYwAWNLObBVkSzfbPD2fpo5oZkuitviXLxD+twruE/gGEGKInLV2d
pDkATyZ40PftodpBQgjyQrvUqiOxcLTVIxTx5oYrnQ8=
`protect END_PROTECTED
