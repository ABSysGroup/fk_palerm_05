`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i3j75ebFbSOilC7F0zWUoO5jnxZaiLzyKiR+w5vlHmYsMw7pw300O7+CVXiSksuv
34Igbk8XjIf45G3qzPkFKYCXv8G8El1/ACwXrTxCDYMqsh2U4crKyH/mrofuMF4I
cdexN5/6dSkpfS/4sN9rtlvm/12MXa7xsE6sMq7FECYVkBzHK+4JTaEGeT3c9EGF
wI8gSUVQD+hbgoVNM9lyswFtz+nEVKk8hlK7De3DkE4+YL/ma8o7OweLlKNZTu7f
BbelzCTZ1z4X0myeBcp3RYJrosbHIhHns8xWf+C2+kFqiBGuq8CEquWk0CDlopQb
u80P4P6DynKkpnfkLIfWD5zTK/mIMmduL+mwlad7QiYrVJflzbpMuOjWWT/EgmqF
1h4MdhdS206m3UV5IAwCxJUwesDDNhx7nCM47n5rByuF59s7q0ut7Efy5Tr9DNiV
rwDOgDuvucRLeQP6/mpyJHsip835mB0xMFWJCW/Dhn/OFEoYvZRC6key26+VDC7P
QR/j2ROBLF/jD0zCWeGuNc0K1pyklJPcElrSOCE4Osznsxao4jixHgR18uwZTnXT
9HAyy2Ebpdgg3RYi6Cf+kzo2YBZCUn/7vb0uI+6Pt2faJTOui0NCszWNlq3OAxPi
wAD1BY3dIYCxdbpAtpreArHAqFrAJAWgHu6O5DbrcacVy2kYCaGAMfgNudnCauz/
sCv4taSiKqnVBORNuyuD7E8oj8+AuKGemd359cN1+aOZPhBOVUQ5EX3C/P0FcUqG
NKfaMv6mR55bCVka+kzejGLm5UJCFiCWhmffkHCpFUs31r7kbYzloOWKjRZ9uaDc
PmD53Rz7uS2LRdK9d4CebZawLJ6mLPtGD4xKIS1qmT9yh91u7WaHc8EWdRVbibVZ
/kVH3YCTo4xNjZWp+relE8lJO9EftGxm6MWt09TXZ2k8SrcHdYvFbjNIzShatz4K
vtDj5vzyRykUUFuzAgvZhmyw2G7x7V3DVMnQYcwsCEObpg3EpMt7AL26IBwg8p1C
wIQ7h+mT+mChIC0NM/N5mCX+nHUlMe6TNBhUKejjXhvPQbQNHYEZG1vDsshObg6N
N1PMFqY42EZCO6F2isTmMMZViLWclErTwANn/W5n+ZtZ4etHlpgo/d/sH/ChujRq
zg+z4WSbUd21Ny+SevxJ6hU3XiXFm6O/GSULqeKvtuSyk5W6kcjlmeIdvbiszFVf
UO+g8hkzChbNWwx5oL7foY5o7PsijpEEV/teO686jqaUO1SOWjn21sUWIEViNXIh
P0qWzVVjU3uZfvjT9CL5jjLSHop/ceX8D4Nx0eCWTYkafeOC3mi+2nAeA6gdoiW3
PIlnhju4kLODzPwCk+kSH3tPleCxcZxs+s6i7EmRYEmZ4WF1JiSB94zsGlg4VQIV
`protect END_PROTECTED
