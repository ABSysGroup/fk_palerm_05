`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mobi7UD7W+iAeu22mFQfZExcngefg7OjA5OsIKU1eALxTcaEgZH6yyKT1ELiE0wQ
5lPVT5UeSEN8MXfahsWVSkQjx1vi1g/ATk6qkCdPFsnsVWBbwUXK8ne0SK7razG3
eUF+eytlcfXdRq75VVLjwp65GJSx8F5DPZinwSz/3ZD151TyJjt37niLZIPWDyXy
nhZCcaesZeSwAnCBkJpf+qyOUF/q12NkPTvn7s8fL/SV5RZw+zZO6cU4bMmLl+is
D3TR95Mwrpmcn8T5MdXq8Q==
`protect END_PROTECTED
