`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qY8gRIAkxdw0v0UanoZimF263EgpdioectiyGCb8VZ+1jfXmprr2kdjIg+h6zH1N
VKVT6UKNfqZNeWNI2dMjvR9r+nP/y1ZkH0unjsNGbYlkWHG7MYDMeq2n4sm/ZpPV
ejCEIDeJkpvu0CVmHOp37oldYsjJ9Jq8xsGKN2LJdPtEw6I8mmOSKH32M1Qf/fby
krFb42cEVklIKhO7OrB/VwKFBDINyO60GPuqk11nEenpoK9fm777hB1cxgEu+47g
HonOA/qAsa2ksyG5b45GpyAggZI2lsv33kTMDKEbt0MJWO8RoC5v5HAnRFg+zt4x
n/bzOyX+BlxUJNsZxvxbz8MVbG1DrvSqK49Gx+JWJjogO0CxDxvzblzwymilcDa/
u2aLN1Kep3Hkwaa10phnfT66ZBhxyePwWQtbGp8m7oyHEE/DQ/PVs18YPl1OEwXv
5mFOBMAYpe7GPpEqOTc+5HBsTVixP3c5wTiSyjGDzEgfW7dcaEPbXxZ2V/S4WTDt
eVeU/gUm9/yfVnF6RQL5HzlffYYh2CA2HszE79G+TLo=
`protect END_PROTECTED
