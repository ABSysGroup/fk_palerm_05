`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7rTJEQCiJG6N4UNrobkxZ9uWKe4M27Z/Q/9BBrepjWcWcWLsXukHuYMGEIjbofSA
fLFdtjPEiYPL0WuoE8L+jIllF/EDx26rdVFrCPR5ht9GeabOfDPE/SRo8PWb1LBT
5PNLXpRbtR+QIJA4XvYoNQ844XXPYFgJZ7ZO4/tv1l6IvIF3sb1KlnNP9HKITUtF
mg8gTs6JoxShquT6bc3A5iBRUtwM7bPCUKd5Z1QuXtBWQpuJpol7Ss71s3O3VuAJ
osHdAAsv9OKxhnHVFMkOBPf0yWysp+9CIbU+HfZDG4uc8jhWrcgl3hents2ThXQb
yTt0GVUZwv7prJKZfHHwbtj1qMmQ2Tc6pIbCb5gmxN8=
`protect END_PROTECTED
