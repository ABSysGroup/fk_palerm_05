`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zYy0BZE7ypy1eqBzpkK/kjlBTmIGVzEkoeKFKdMpWwxs2289Hxyyr2maU3MPFrpr
1CRyKILbmx1tjCdoNWDQfnJ5pac9DoNQglCTG31yc5rtr0Lx9KIX/Xe5C9JJpQmD
AicmL2tfnPGImdjWSpemZqRGVXnvckLKfpSr7ko9xfHufyA9swf/+yo2GGipuDpz
g7vmjBbkrUtI2VjWyCuF7SgAN1MigUr2b/Kumydp2FEybqUZZfIITofGIkn9zFJu
9iMVnkJHb/n5AjVmAAy4ZcP6XuvopwQlF0r8nW7ZAwS1mlJmp46WtJ+vq8t9D439
/I3K7+CGh8PkWvdJxecIaj5nwrsrmEBLh250/AEc6gfJs+LYybpv7EAXL2FV4RbC
fpaKB1ByLxbwQMx/aGFcGybPTUdn+GwClhO5oIcyfemWg893B69dv08Tt3tyJJst
ZIBmNH3DJV/PZ0voTENaV8TzhGWZxDEqvRd7+rizxLaZNAaeaDfW7gh0MNWOeYOp
SFQ0xVY2TEAi5n8l1T1K7sGA4048r88PQ1wusM1B0EbQARdpi0DdVKq4psOFpckI
vnfHoSO2FSLxFEiob9vivtUtiyt6icSs6VPO6RG/0QSsxztsd8n163kXrX4xtLuz
OSmcSRLDF8DNpOa41+qkAA==
`protect END_PROTECTED
