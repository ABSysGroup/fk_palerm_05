`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bcrzhBCKTxeR+6sV89dPE5O4UpvXTBuSOchqAruysO+VmPucZXitMUH9KwxVKyGF
uHRe26VbH/wgY6ZK+buYy1cXLl8CDADC8LUtAmFPKHZWEFyK0eTg+dNpcq+JkfuV
5MwsJkY+X/wn3ojY1s+bY/AqYACdocr/kxCnHfE9pf/hZID4WTDQa/EHHnLChhKe
NgP8r3N3BXggGzmDIzJGmsPea9ypTfwoMNYTNRQoG/s0bYyscQM1CFETf8HfkLKS
nSPtUiorKqUWo4JVzMN5OZOeA2HvBybjy/2cdmi1MmPa0YG2k5ENEOw5GZ1F1g2U
opKeIt4spaq1vuK0+clb12C2cKg0otrG6LMbh5GrXmeutalU63rlqlgVp7kMlhai
h4RNJo99O9OwO4707Jg9ow==
`protect END_PROTECTED
