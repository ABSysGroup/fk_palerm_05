`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KCdbEGk6eI/NVlCpQ7VUKQrXqXCJALNpkHZEaXWAPcb9Y6TgAffZmsubYFrwESuF
nfWASsq/i86yrKwqfa7F1a005fJQB61wwfE48yZSVrRdpErR24fB2jtutBJk3oWz
GN7Z91n0ynH+DnZkOxaMmSEBkTwlPelqMvVaHjyYuseaXmvVH4QEbVv6VMOQHCp2
L3COKtFnyfNy5YW95lM8Plwn8VgiBJzYJGca3a6HjujyUnD7Cv1pfIiiDSjftOhK
TtmAipwGChwj96lvmhovV/fKgMgg+mW42wuxTTnJ7pb4OkM2MXDqRQWOKkGIz1CR
O8BKEoMYWowwSefYlbvt09X+SnOC+Ze8euIDLQomEI18jaY4M6Ff83rKwA97deDf
O5gmgUzXocDikxPh5107/L5E8KKQpV0bxunH4WO4S70e3Ya8kRdS2G+PkcscQT/F
oewhNea5KRMkfAzyLDBE4doRlrxRDPkIK35yK1Zih8qPbNESSz4jTyZPhTVPSbdI
QmidXWpoTkW/7nvG+eeg4YrRv2FiZpQdBGFmEc/L6h28h2NVF/CBn9QhotMFxshN
NtdT0HXDdrMbA1XBflSw227nQWt9TQJhO9qm7RI4OPaPZkO1m1FfHW6M6ffxVxGj
ihZVnwvxwLb7g4r5sZQ+aK2rWUuUocT+xgZJLAiHsezoyc9OzTreA8Ny2V/oPSmm
f5SXGRUyIXWCx/TsoPqwy1IhNN7Adf6M3tgT2gRCapbr0qqN8WNIxHFGRlA+i2E1
NHs6RKgZiXG0muUtHC6xmlhKGcc5GMyVklwcNU1aTT+H3WAUBPCVTTdzEpuxHS4q
JJKyKxB0legL51Bdpt1PrlNYXpFEUdb5pE4X9MfbAQJRruI1DpH77hAqkN9wU8/G
RqexuOxKNHwG97M4EWNgylJy3fehvi2rcANkYqj3bk13HeY76oIRM0ABkUOVBXeo
pp1IJINNneSS1PI1mlXmmN/U2u/ACXNNCwxxsVz58Zx5BJajsb1OtpvOHYpsvytO
pxvhGTHrSVoGsXLU8S+zR6CrKcBaXayokX1/LAv5gVhQsF92sE41S0J7rhtN0BNg
LDO5CUPiOHzCeXeiw5BEfOOOVPn1M8pZMFYgQtCmX/80x0K1fljhhbiASSyjryuF
/CRoPa4j5tXaugB/1FdubQ==
`protect END_PROTECTED
