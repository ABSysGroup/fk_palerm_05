`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
omTHWUK8J3Ub8esAkpHle6oiEv/FJxNFL6xSnnWvtSane22vtxDTwHnDmYFGb6Ii
oqF5zwflqxNVn0TrrNXn50czIwyNRMGAwn7K9b3bWcuzD3izoIZNSD6+n2xCgcf4
hS/ylXkR9FaUkjfnx0YBmVm2Z8QdM0qQLOjB/I/Zbcb/+3K6VVu9O+QduM9G1R0c
KYkfaWQxslAou3mQJ2wDodVOQdrhbhf1yBmMzoNl/b4oyFJbgXNGuA1iFhkK7wV+
h/eSL45u2GPeCU/XVCYV7QxcJTh+Hyqz7QYdCBknGCdvuOO+KCTUMo4a+HkYpD1q
h+0q29wTUyy6rZkbwlFlbKpZ6RXqZxLoK79cku/2h5Ra2/9JmCEL26ArJadRVkHV
InuLRZzFrUkKAr12WnGgz5DX7MTt0H/nKfTY+Y33Ma8xwJclEEv0D5R2IbXRgngf
sn9g1VWNgoVB169UM5R4vLD1PGpq+JsHJs7otiNQJMVIg1j5DQJTqPDXB8PyHb8H
wxBbtUBoPqwysGjudOjeqnQgGMREIwwK4B87MOvyKnhXBe5Pcw7b56bPQbk5EjEu
x+ISYPFTlzgwDsO3tp1MQ8PKzNPiw/4abPwKq1wi5ALnn3Pn4FRGVA0axKfrzlLX
r1P4mgmPVIm/IA4G14ZKT+NxnXWOcCqt9dK8bwL8oS8iKgQOzAaMjx3+iB1UiIHf
V31jyxCCzOz9EZaTLfcjDDYXiuj493mrKuwlCcLrY8GDrZfHAV4juub/qJOvZii/
iVrm/NFeXOW+lj3KO0yixIty8ZDjYAVeEZT7bxXJB6Z1QC+wBlnrpj+U2bEmbgdP
KnOnEXfM6WtwxwZioErn/BFx2JknEIwUBl5uXp9BsH6MdYnAaZSn/vlIci9aCWsg
xNdyIKGrNB08joYzaT/I33FBTJoJfJUmrzQFeEUPOBf10I0Z3nqrftKq2LQ9INzm
5UZHZg2DzEc21jpXbOVlxaQ7IfyyCYdZoShy55yELIO6bZ8H3EvmBV40p+gvZTvF
uTdukb+nMrfa5044QkfowVKMQKtxjqfAtMa9P7aN9rjYxmy+lZ6rw+vkO5Cxw3FM
y94mUCtYaZSYDVAAtQHZWA==
`protect END_PROTECTED
