`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BuB1OH7u32JjtBwkFx31xq7Vrj9eXzxVpjV2lgz0KqwivIHcFSD6h2t8t+mIU2S2
mv3cJnOptUi9XZVqJuGcwgEE0BlyMqPhaX8bh/hLw920OmA0EQOu6lw2+vGkmk4B
eCMYyCpjk6ChN9PMyQWXki2R6D+LAYwt+G0nYytVpdF7T1zQZfUoyMSGWOKADcHh
RWg/g3nvSuvvprudMJ/08hs7cORBVcVI4OEGgsWkRlxPQdgrx/GgOZXbFay4Uvs5
q5wIULRjjn2bEb1IDSFJtmCruzkJeKptIuWOLEBzd3Bqa7GBCdv093/pOyxLi9/z
NkEG4p2OfIhJx5yMOeUDi6rtp0PMY1Vk9CzC/ULpdp1poH7upb3ehASk0vQLbEsU
WVxHYl+HkrWuty+PiUQ1IJuGA2J8qcuKx9TAdl1Pn5S1QOlRnJzkRUBVZmJWxEDB
E2A70xxsU296Q/nzHGg0j54sOsfC1Xhvm/ZasDUmiVVGglhdil7VX85xNeeToJ0N
2rA9eWV5GfabGhvHupFYyI5JxsvoEPSQx8eOnw7UHbTqWUM0pyl8E+wYqGKwy8uc
Xm8wUVC0JSrTi7lrAaww4XjH5kTJq4tFEIBfwVyRNql0V3Kg+s1X5Gl3kU+Jz8hI
/UWMTJ7l0LJVBlnV7C8MKUG4btbTRwYR4XXDBV2ghbyDgrxcNrNrJNdp5ryv7dfg
uVmKuM/y7JJjzQrQ6PxxPKEHOAFIUynncFsLUDBmEPFr5R2dgjk+YJVHLaDhJgBL
5dNzU/dF4DR5ae7BmEveY2CE6dPwo31WklmLDhwrVY3JhgPVHvO0em/XVf6dEcXy
tyJ/uuu36h2kvWbbPA7BBaXu0laYjnhS3/a5k6KVmh5DLMSTA/yXAS0hqCaSgseM
dvoIHQUuKpDmQkhco7gaFrqFtW7WfgwS1at1JU+wOPI2/oMXtBB3rjqW8ZlS4O0t
JVeBNIwocew4BhGNjVhCRZt2Egw5StUnJzT546rbIOeTt8uHKKfgHfoJfyzoPhQM
gB0I6eO0rVeZ7PTsrDgvxu7dhPHSnVVcYmmn+V98QAiqsJkRMVpNpjC5EMS6D4ny
P771N+DjOH7/u3k5qpMgAKTULmadtOI8oTRe0O9RNek=
`protect END_PROTECTED
