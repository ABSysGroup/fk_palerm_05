`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YpRAlfTLTeMWj0JuigQ2Lu1Jud78gVSYKru7A8klGDVTn8o0B6ZtH5k7XVWuy+LH
MLpbPGy/RKcnuBg59+Hz15i1vPnJdzvzlamgsJ6P6eFk7LZsVFypoVNbBeXXIUce
cEOizASDxyirJ/0XIu2M3uAYep99KU0hTRAryipMlBIS2yRx1HbzqTXCU/qv1eBd
+4v8q50GyK1ceFE+M7pzv2yXUwU27SbD3WK8C7dLuvWCnJMw6jK6iHFXpGjTLEjI
4bYJqOx9s3q+awp70DiN/xSSnj7bs8zEU0bI5zVd/f9yUTPgu61DTeh/mFQR/8ke
bto2uX+WHbyO9qdDV4uttz2WzM68TY+aYAsQnd4yrYQ3zECYrawE5ny60YjxRuHN
kBYXVxsp7z0JDd7n6XKB3nf09tFWnZZ7AgvcL3JYL9w0b2kfWUpK1NzMl+X/fgfA
bjIIKboFO/2DabI31YExbZKqSzGLgwOTU26VGxs4BFe1wttILVXanMA0pNYVaG6+
utTtnLADuPb2Ql8BZDt7aWjrjPKjBUPp8OrLckfmv4pgrCYTib3WLHK4W79vRZgg
RPwIHD3vdc3PGGI3qc+Mfe+EDJWYsR8ue0W0vWXjZoY9g7QxZjXfjIak55mMfa+j
yl3iPKFPG0rMz0lhsYllsJSNUcWIBtzf6+QDqk8pBmLsLvIIP2k7WH8xuGgNOG+f
kSiEzjAh6+2voAcqc9MrgmvU1/74n1FiIUc4YRBcDo42VcoAztB2NcTgdyHX0VIr
PWUJNJg0LG7vz2qXXcVcxg==
`protect END_PROTECTED
