`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JvK6ifJOiVwx5Ciy1A4wpqNY2xksEpDCQ+IZWGdxFptsBLEvClw3WHJwloocJeYo
T4BtGUOablDIvk8BSy7s/e6DyWdoX9M+NeQWdQvshV8bHBPExcmZ7bN+MuHmLtUq
3uAg2Tegx9DMFtTF0EvcRVi1iQPLACrGjgRHHGgNyvpti2aQLUIi9V33dZ1UBbcc
w5g+PuNHstNgKT93ZFdysm08Z9atl/DdQh3wG/bTAwq8mtEXc23eVc3u8eVCibco
6Y840qEDPjUfVcGRQLyVZQ==
`protect END_PROTECTED
