`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n93xvGGSDFE/dI3PqvSmRE36HrbQB9A4VmaG9VA4eH5UfXg6CBqXFl/vracqWscS
8Lxkipj+SbHye7/M2MREbiYZyNNLRm0Pndv+5fHbQmYOe4eDUfDmxE7wah38RpxI
WT9P7GMg6QX8w9oq9lr6poioF5hPIkBlom4k2U0iPzzjMwa5S0fkeG9HfN9HGQQ9
yi/DdTat4LGuMShhy6iV1IB4zTVmKOgS3juB2P2YOsT36bgnoqBCJ9gbl7GZMy5F
DI7NPM8WnyRIH5cCbh0qiUNcZuayz1gatBZy0JmDjHWhbpA0TMVeaTkgKijN4t5Q
DMo3rHQi178QTltdg+6R+bq2+Sp567s2Ktn2V+KfONIrAt4lsRnWRUlyes/wsg6h
KQJjGEZ165lsDFvnsXrZPrqPZCbn6Sqffvqxud71/CIs3U1uXNpud4oylxHIXmXR
6LPOiopBYx7k554b7tUQzC3vrOvMO1quDjY+C0eH19l9+d37GJZpDzpBZnuZDmJR
BCLCyvqv4MbDFta/x/elY3CsOI3OvmYQuJ+qUYNYU5qtCgo2F9JFhzqON3PZIkZJ
0sLca99MyWpir61/k9iwsEDQI6TL+ez6Wok1hsSnfIrdRNokN0FoxTREvUKPWMc/
ADJIOLq0KfwwIT253SWXrj82nXu7JN6nKHzIYs1hvbZpj7cQT3EY/nnBBSajFgSp
0B3RB5cyufbXAnD2iAYsvphv59/r/Uc7lSZPkqtBmzomJdB/LqjzUhvO09Hc3QWR
v1dP8t/q2mE2x/uwgZs6IZmAkJB0oMhSegHZ8L8euvibHQrCf5Xb/hdERWgchuKY
BBRvGAtAMWxL1V31hyhpbKRADMmmVy9Cit2AP6DbBo63Jbb7pvDnP4cluMZhM062
eveSwHtdGDrC5viNyN2sAcBccVb60xLYj6PRlU3hoeI+w4Q1T5xnYdkS8lrIIU/f
ukQr8MTa+CSdVYdijU8dgnqaBerF8DSA8MVLmNSjDqVD6f5cgLW2YOcWz5NQgQ8J
qPe6Bc/DKxv5wfSB6WdCo7YO4Rf9/m4/YvId10MDLOvmbjWYaqhZ9qB5zx2YL61H
QHXIoL1kb37ut7xF+7qcs30BKEl8PO+Icmht3lMiTog8yRx5CaDIvCV0Dr8aLDWw
53KeXie+Wuw9yXoXcnm/M/7atebYBp7qNLqwXuUJSgNlRgpqUwa+BCnjKvJdz3JW
MopDgSVeIdeDAqD+i1H48YHAR7imm6kmc6dWz0at8rQT0uDNo86p/RKRrWFebT8C
d1/EqjJCmzubo+HLsIjsNCp6jEuehIAWv2TMy0YhGSwCvCzT6wnqN4gIQglgIQN3
YWHkCzhT7vzZ9cv7Y2eJpUcBhzSe7XSIeVc9as+fS98HnB3KrepRHRUrd7SYjNt9
zBVatFTyxTFoL3gyxnbLqLxWGiJ4hcOp8XPdDUY9lkMPgsrZp5/vUIGJwquM22fX
nO0jc1Q8KNRYMWUv8qdxiw==
`protect END_PROTECTED
