`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0ZhaO1Dt9BrZjCz6csullnLrWxOhMJ9qEgfhyDM5WLL6imwhndciSk/dA8zP1KBF
jZasknWgIylolKom7cQmfpWwGlMuIAooxhQMmJxOvVeWLfVWXSnLuLtaD2HpVbBk
VEaYW/nRtWOVwSm1Gjz3WfSdx2HZMPfpFdrJQ819doCUXxJYjgiNhclRkRvYFc4e
PIvGLYSQXIikQZTQAlR4h3rHXnEMb6nvxHn80YciY0OR5Onosq/8ECecv0xTuKFM
DTdPax+KWTO/e3w4KYPB5cQVXch5liQLs8XaOmxl0JCQX0If/oP8bAKrUGiWjFB6
50XFFIk7ljxFKhLlIixRO1Wa6mL5DoQ1jZdOyBdllnkJSHZEA3jBxGG+4CuKik2e
XVhPaQG9/ZMeem7QmiEdzy6o2vhYZx2cnKQDsooRAvaXHvjlE5RtK7ytbyzIHGjL
TulvoX9Tk3Bj9flxxdlcz59aQSPHRKhKO3owQ7MU4mAZmUzWOEoVTM05AIz7G4Q8
LLAONWAB5rG2XpApRe+dXQschq75TaVJPF8r/uF10kwChc5VhNM59DCJlpGdkKMi
k2sk2wf4ZzqZJUUEzfNoKYve0PHMu06mDvbBZEtHuTPdjBUKmDPgEIixHOGFMXcQ
ijHUpI37N6vUWB90fC8E7k/cpvjnWSBNru29RgncosWQW5BDaSy2G4mL3n5He4xk
TT4UAoiaxs6a6c3MffE1UrLyooRrxcYled+fGNjxmE6WMf3sv/9mh/ERYtp3l6Ok
zBI5K+z6Z+q1AvlUYPd3+Hi1UQl4czi+m4yD027N9eKKeJwt/CYnzQwddxtnFUAK
yxOR6VbXUvHFoj0sf5HkRK6g4+3nIjwHATdrME/X7IEF46hhLiFjWDgWd+259kbJ
UvFlPMRCjmpFC5wJB4p5b0pPYOC/rNxJfklScP6G8N14wkz1S1FDlxzSzVdBCbCJ
mJUBivMOukA7Gz/LkauQzfpwgbMYKblZ4RWH1JACioj/OgpqwsR29DunadmmcNuu
mHweDtgiUM7VdLQF4Pn6XkjFlEjtDBEIhwHjRXtfv9nm8Y1APPWRq2GmlNomMGft
163PySNasvydqv2WLAV0g83ZRW5XdqqunuLQNzA5sEgsGodFmWdk3B6nh8L1yiHk
pAUIkr+6k3b7J0ZagUpsKaQGuEOKvCOp98ntUKLXJIKYEouh5sQLPY74t3W9N48K
UX97gnXz3s6Ig27Uu+Z5FW6FyhRF+3SU3lX7MckOT8SvCQbFNN2pyUMbxfR/7ymD
v6XlqwsvZF5K1MxXcqbFSIfX96cMAdW4GrDmQqciNbofI3v30sRk1bQqrdMwbjwW
Yx1Kb4mA0MnnWJ++yxUoq4kq2StUb4qFqOJ0IxvIvRCLGvOxdpqy8cT1Gzm/zQwK
vxjNNOMD7mPPlPJLVG6QMWN3pw+5Bipz6U27meERS2tmPDh3R/2lX+Nnj6Cf2t3K
D2HyUvYJycvx2g8G6xAvFc1tFGH1Z6cWEdpUgZAH8sNS9N7Jl6mJVSpUfaYm5myR
8KmJlZpyafmsxnnY47JefolDyPbpVM47Jd8MvHgtl2G5qNctGIy4Osr1QK7KUCa9
ufBipGSnRHcgvHgHeWaKLtIi3AqMOa6GTZwcRcH/BAPv++M7JVkj3LyTM6Eqyunv
T8V5ou24TsonhusofHR032rdwTnT25iG80t4usudTq+YEfpawlHoFMY7aSqiKRgM
54oyXAPr70HoMfsPfaUQWjWBRl1isUUWcAt9OBOP4xEjC9vLeG9942GFPHhAFTN9
K994o7NyypZkFUsMBhIGM8pk7j8oGoWmnKH48x//ckm0colpezDgCQZIpK4g7mRa
7xQGAMza6e0MGx9y2iBFwUi8tIQl/ZmOQ0n7sqg93ZjIMSvkGMm2fGnHHs769LXE
4B+vHk5/imN9sz0cU7ijT748Km5qV9eFOzPis8xHlhECeuwIwj6jJrBTAgk6veDR
kZK1s971RQzJiZ//cTdAVIbuCOmuETO1AebMdaz5yVpJoqWJKK1m5J7L4AkANunR
CEI1loKmP7RolapHTyWImc7xsqZ/9G/UgBfB7x+o4xz/nsR8aPjpm2lAKNfjTiPn
9swDr0hW0MA8th2SKdl7QMMh2Y/ak/NoGyVIv2PO9oBJNYEoiV8haiHcgvo6g5Ks
SHhol75RYygbQl3xpnWEP3C8DHVfhSqzM1+E3vGR0FsYPFUfxekiSdQm3AFLOiTg
oPu0EX/cxd9FJmG4cRDr4Zq4Qont6EepSjNN+18SQhbmrEq6wq8+jEa1Y6KlViKA
kJn6VTIVAmV6i1dkYLTGiiy5agRfRKg3+bemiy+dB1F7P0KLULv8WkC1X9bk9ex5
jRWaLqkrstlMlTohmZYJwWjDdidv7dqtXSD1h6Nu8EyXQ+TfI7PihCn4BEsrEoYR
8hAnqJNVnI93gItaIteols5LcDBOWEYbvjNaiZCAi2g05Swcxplvjz3uD4LILlzg
r4gy9d2AR2KOLzmOekAnVW9EQMKzN2dS7ry6UkPeMMq3h8wuk3z86Mxo4lbUPPvx
JrcfmH/1tTg/kQ7+tWtTPeAfc14RzMspzp0JuU50wNoVNy1owxuKelBbr6dT+CLp
XUyEaLkGOoKedjx6iIQ8MlGVFdhTj3me6nNYulkzHJ1ocgQjsVrzodvKYJvFIz8r
y/ooBviuNPCOcr6gAHTHDMIxrkQw/nI4w2u7QbcBd8bKFboBF0XssVT3BlHQCpnG
8skUq6AW3aBb+6EfdFW/i37gVdtGEaWAPE49NtedrUgC0eS5c5929yc8VKdSj3jr
LcGjSj9Ujb/ZYRG0xOK2oBaz6q3VmlaNUATajXJKi50aDcCUfx4/ULc9h59QK0sb
/4v1T4WM1/kbuAZh/QAXt84oMqKi4iHC98Q+NDTkNdwoTko7njCjMZSNgwHo5eIr
ZeRJCJU7wn9eimZ26WesQep5iQInpDG/c62omhjZnuyOsjeXE8aC2qv86FRp1gCW
5mwkGiuzRYZgjJWAjbiTKpC000HYjeXaKDgy2PkfNrbCYfpCK+TPxeGJBsAy5H2Z
qYUL88b/InmN/tCve9lhzWJ1tAZyYZhiG58cAEKUzYuaWq68mh4KL7K8DNhnJ4UZ
U+kZNe3upv80pIaRoXK5OdKB3HBHAm0Z+y+yrNcyY5hIBldOnyRR6lPXEK47jqzk
Qz+BKV6z70nVqhkrEhgpMKx45GWZE3SxgCBgqWc7iJ3FTYpL9bZrM6SluPNAl0F9
ku3iZdWbJTBsJ8nCbJsORipKW8Q9bPvmdNhedfPHfDvCtn1WrhiVvs83lKKRZfo7
L3dJ76BDHs/HPDB5KtTqS7tc/LeAewfwDxG3jCkC8C0Sog5WFFCEOAhPxZgJ/pbV
3z1ekWVLJ9jJKgNZ1DWfFYx+D9xG3usdi3kZ78kQiKKdnobP7nNoFMFCAe30ilm+
7/msIygGWTDS4cSixRBT/xJiClKv86QFnAioXNZuIU/3pGDfGtDref/TYifvvb0z
ZXOORYNkNoKfRZy5hAUDMn11Yk6R4zDajhu/B8c1OInDukzzvoFXRpDLdVA1lXqa
HGQ8Cts+KBG6XIxAxfkGGZEhb3jccmCjj6qEsaWNRoR2oeCmNk224+BK37ONBDSv
Y1O4ZWPMi/kkQGuf6rEQrwqzkxj/Ef0laLi+mkUpjlSFxI612aOX36Up8MNF0Cn8
LE+/Z3XC94HD6f8fvbc4xDpQAw+rnmCUlK6IYmueb4bfHwpjcy0eBenHM4Ao8dHK
LNT0rBdWEYlXkxFWRDJ0VlAO0r6Duv9gZq4uPeqgsDeFKN44rfCb2OreGeGiLI6I
/yVdoEN0tI1Om8fQhe/dG8UVkaiDEqQtIc6O6Ig5iwVXeC0J1ZjAsxtj+3QUXZ5k
IuPSAvfrK9iaW/EKmbhllE1wAd6z5yeGqeKXQnmVNSqOyvJ/0EjzFAW+zWGKB4yu
F+E4tZrJUu3fWT0IZouaFL3nGPJgXamDcNzfLrvBpjdP92pnYu01OXrdg8gYyzY2
BnUbTY/3i19FQkpmpGP1eQcVfi+t/lA0y1ARKJZ34FMJVIL3I13QYIcbgrfIj709
MTMpMH6c6aVsJzDfoufyd1QDcmYVSAqjcU7wLaQ6aIEAYJOgeTdUdKCuWxulrNa5
hBZ9sVRXaL/siScbnpA9sx204ILMOWl5EC34sYjwCBmXwi0X+EAG+K2XUfRb3Xal
zD17RtE8Ki1oTvDB2bXlxsfyy1fCUdLnnr5iOxg9U6F0n3dCUMuS1M9x7A/Vx2t1
Q88P9YHVq+BXbX+ZiCTUAtotxHcdgpcEFXedQ2v2W7eLf7nRWep6MTUBRgAxahPf
rJqxMpyht3CXF+zOucxAclI8AMdfW5dqkDTQjK0+FfKO7iukKC7oGn+wlarN1SHM
u+5Hbxg6qkkEJOZ+Dv+zOA==
`protect END_PROTECTED
