`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l5ZY116u1addaxUK9ZvXRlANbnAqQk7hXB04qncibVGwEeIlJQrOL0TfZSy5Q7WD
hRtAQOOsfKFFUWAJDWkWXOz878lcQkXt5/cqowMm1yfEnm3rIux5dxf/IjV3M30E
WHXRulHPlDHNwIAC2rLqTh+nrNk5ul7gCeD4HhUPyEJ5UzVWEalQijmkRDc5kfk4
i8FJrhdV2T6rauBwSeL9EUEVeVvSd8b4uS+b4m37o9ecnGm0c1s5m/oPGQqhv/I8
MsQ50Qqi9H7WFWj0OvkLj/ipqQZoopiP70HFH2DMEhF941hL1FtMC7P5V7sSzkk+
xBcY9BU0i/Ud4m66GicI0EvaaAT7GAcj6PAAs54zsCvcNaHSaTL2Bt4FpdomSdm+
zuZ0M33bMk+8D8uc+vBOElT+/KHWC8iwPe+kgxi5rNCv4NFPDv59E33vKW4lNeuH
2jdoWI7PqJMJkIftADwxeBAbQWezPwyKzV5pQ2qVb9iGQzBukUAuWG2VEWMevtoU
EQOk5X4K1nLlE3eg1bTQUiCAPFwsuQReFN2t0Gl5g/xWYTzTcr7ZL9M/7yT6en21
ZSe0wNCS/EXdbBPQv81E9NYH12jLRG9Zr+0YQZf/cCuLsssU422f2M6DY7UUH9G4
+andk+8DbTht+jPyC/5RJQfL8X7uEhYqJpQsd7fWUtbB0T/DMi0a+scXhywHD404
T2sc9mdr5c4i9gAChBdWGNOyi/bxq4KtuwqbnMQNHf0=
`protect END_PROTECTED
