`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HyxDCvw/l1UhdMIiws/Db8dyTNWRRdBiSFgwxtybNccYXEeoT9iixkAzACcU/8BU
d0i6eWXVEDeKyACH+vgVUJL5wp8iEH141Lv+h0oOBzGCLJBAGNrTPaD5BTVpNM9C
+m8kY4fNtKmRPcinfDjjKYFFxONFYXl5P3MyiG6tV2Qt+sjcvIMo4HyHdS+p8FEm
GvCxHMX7HM30GSRM5vM6hd21/uiZ6bgeyeh8wTGzfGEYjrm0x5JgRsWZpaZyw6oJ
XLSV71qqTqYvvTb53bmqrTP4SCcLTWazA9FJ0yXVH/u5e5lZ3XZ3J9F8cWwmbpR/
/++acXfzQP8XXkLC+iOpK6N9TIXae0P26IMcRbuk56kuR3eAe4w0uVByQQgIdaTW
TK1RX9/lbNrqFVscC0NG8S9hrcFlQEOBoYKHpafK2IyOxDlI+VWzX5hQBCWP4kCK
c1FuS3VCYthGPXcqMo5hxiEI2eYxSe0/dPkhB+3hHIDdQgp3jyVrpEdwHTenCrlS
uJ9Erce2IY6857ODEk5PGCr/Zfm7TNX7SM/zcZqtEe7bETFnJ53dF4hN7fQ90iTK
aIiYy+qUhyjiKGO5cLcRl4Elv7hqs9vd/wj3AvChq68sTN1P67uO+CtFhVq76Jb1
sYh2FxyyTAUtXkts0cSj3oyBm0LJudWgGJm7YaPx+z1pQE66BReoh4dze/NdaH7E
YZxj7q1LAgwdjL50ZVrRTCknBmo5K6Jm7pzzbOXL7Cvkf7L+lK4Lb7ZkHauMvj0H
w8nOuTZm30dOoOuJwYCNRALBsbWyxOXtPCWTQvq8H09uXnjqmZVKQXnElOG3etWV
RqLXJR6dQlfEeaboZ7clRfzlZ6m471NM4TwZxLpojvq2mGssqo1Xl0qZ9If4DPIa
`protect END_PROTECTED
