`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q0jvlM+XXJwhYvJ3QLUxfDFhQDTVKNbnEZS5ct7swZWeD75f6XvF/DAc+p+tdpUm
4qTf/MSo5efYlM71icJeIuC8aCcAdX7A+CIdvtdrpFKmL+gZydphSJMi8YIsbcIc
tpcWoQ2XfpoSqAGcj4GyEr1E4eUDMUW8IkIgJd/3xjlDqZ9vntDtNaw7lYf4mqtj
bwCLwViP1imh3IOTwQzLJenXxV+UBLLxxY71TY3qtMHEMXMNzp05KIT/woKvqZm/
aoHYGx3z85W3ss9TirKVTSbD1jdras1dI4u8D+ozqt4G4ss0mYNnmI3PzA40hfmq
`protect END_PROTECTED
