`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Da9RwCrY8EEnOYzYi4Gt7Ze6msWpiSpg3VT+UVyYyZzQ89kkKudNsCwosfiCyYcH
SrFBZk/z05WAt4bh2aIU05Mw1kjOL5omeTdqTUcdqZCn/WvyKTBjKtlCNGz8GVkw
v4H3Q3LN9KcqJkRipdqF86kshPHTgQZtoJgterb7Jhat5Htio8FLOckDde+gIZ3x
Y9q8NPmWWj577MTe9EmpeDhY2onIvZjG+fLPHHb2GKZnJ0b9on5XeYKB6FNXdORf
aqdDJTCceq1V/8hGphNgBaPjMlT9huVc6luklskB29hV3EE/UQpfqAHE82BpbYy3
PbIXYTPLhhEi+xSOjK9cEFu/K/RzeK4+1LPi8i8j9GgP0Bf2RWLK5tW5woM6sm+9
mSXz1o3rnhWFkfphhwu1885+M0CO/0VYQiAlwML4SEQAvq+JWILxQPIy0PBcLc2U
YvsSklKHOCqgh9C5i5aHaSiNKe67iiytNLg5J4UhSYU1qLSHrOwYgnmc37dd+O9e
bKiKgK9VP2Lcq0PCwKQdKi4YW8H9BPHleteV5INzlORFcvbU2VcapIpZlxlZih1p
/uwT9eK3ZtcnhxmxTIqjTQ==
`protect END_PROTECTED
