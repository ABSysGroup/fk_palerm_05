`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+PaRwoLF2Rl42XoiwAvfP05MuMoUETp3mgwXwGb35z9DEKQCxstXrGzQm6fPTJ3y
wxLP2itY9KkRSLwpV3qfldhbQbw4QckffJSDPTaP1UjJ5LAlxeKLmhsly9Bm9Ka6
fcpsUlPsnh6ikCrO+KqWzWdlWQ87r3ZowNkM1oji4tY+8pAooK5+nyN0kAnOkjf/
mqGew7c2woBiWTa9/nkm0X2OYEJY8gR/TVNASzNRd+KibFfXIJimMkDqS0sdWI9T
Y2BXeSaDJX9E3HiXToc9hkDkFGOOIGpCZTSUPkiQOZODNUiSlOwb7E1Ai4eEV7GA
uQB9eWNiJW7c/xMwHQF9du/CNwbHWmhl8amM1QJHURtWFmOQX7hFj64/q/inmJix
g2tTs4STlVNu3pF9aipntsNX843OPJ9DhXCWhfe3iT6t4E/HT51U2NLXBiN27ahQ
mVfCMzFytuCDgzTGFd2JXwYQuynEhCspSMTCrUmjq1KhoTvbDR9dwCBP/6Jiql/5
B1AISt+k9k0Ud5YpVObr4wOAjMjysyZJ/5sEugwSK7/L/jpTscVPXh+qUPRBxeGI
kl7fLslvK2QFa/5noYP3/o6wTCTL80HgCqsEi6FY4nO6lzd6sJnhWDdtsMWAX8+g
1hZiq98db5fmTxzOXI6Wjq8MGcmvxqqnafRljnN+pC7mGR/0hRFCqML7PrwZO6c+
Xv/iY1Ft1Ct5yrR8/nMIxJPLnGSb1PG9O+Ifjy5Gm6c8L1TUIQrSwUh7InY6heI+
u7UA9f3Wzmz2GGy9gV3WvGVmABf5eEWIJZzH/I8YpVkZjZvesz8aI0J5bF/duvk4
eC8tPweZp7eogUbKfIU/nz8fDbix3Rzb+J+a0gHpFcRdjKz07UcHS6IuHqrYa//I
QDVulzQdm8AR9TJjIToukD4DSfyLtiegmd8pi7il+pL2QrNoGsn9N/eH7W0YxbT+
`protect END_PROTECTED
