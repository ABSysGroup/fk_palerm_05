`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U9yaynDWoqXrynx5bnevXl9ZtlSJRtWZmgzVko1m+Dp6cMNOvEVlTUKhJBNm0rRA
uh/eCGQHiayyby+jQc5A7T+LzSwIZqi+PikSUFCF+HzqOQx9GTwJZTW8VErt8UXW
8s39nUIWmLNOlSMyReTeDAMYPnOgCqQJ+6dYww1nxlmf9qWCZX3+GxbAGSLJJXkH
mQp5ICh8bD+eNZPEq1tqGzr4pCYU4yBLjfotoDP1xTyY8gBu2tVfPP5QRCcHVGEZ
C/cHGKfcWJ+tfN0W+QVQZF7QI9XaXSveJ6nOnrH2BLRlplznMBDTiMdItHMnPe4b
3T1vjfxLclsn98qehSaq6JSt9d7xINuAObFZyAiGKAuMSBWlKz0hWVoNJGNJO1in
U6q5ila1Fplv/Ar6Ib63WA==
`protect END_PROTECTED
