`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RbTfJ7xpLuf3Qdxf6i/pjroMl5eupoQHP50dzfklK9YWAto8rig3ejxOkS6sVdYx
uA/0mps1Ki3YVM1i+lF3bVHJ1sUQZMmJ6pN6KUyjfdrACYNnr31Tz90n1Cgaatq3
QSofz/9/LVjEKmTaTwBr9vNOkhVheGNjWvJ/+lRid8ArFHMC/9hjv7jOSS1S7MO+
IzBPsLrYFt7+VPog6g+KgHtTG+P94i7ud1PHD9Cidverjln0byCgEWoS2CqA2/5C
lkDA//F8lggR1Q4mYKX7P44XcpQVLpfhxwH9AJ9HW6oKSREXt59wRrg5ILjeEr0S
Lodq3wOLfjOPsTzksfH0nWfmFqZjE6Z9dOzEuUhUysu4dIjGge47ZUgyfqT26oVm
yxlyUZDajON1OW1KcwoIAVNvOTk1tSmKbozNjxIC1UK57Rgn4y42oE2Jn/AlHOum
zHBfSZU1FnAp3tCkUdPPpVpI1A6IaOF2c6BWgmQ1d5NctYfB87xX1jBJhlSD33mF
2lC5Upig8Sh527rTIyMMp/WA6HBX2JKsGlHJQwuih1U6AyS6BMv2X/1GZrmdtWFh
BtYDXfcNL8ONKwclIYycTCd0IEoBvZbyKx9Pdphry6w=
`protect END_PROTECTED
