`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NjvU4q8VYz96YdDkqjwtnderSaqaEfUHgOjF+PlCe1UJcmuUq1qW3eydPgOvue7b
7jneVF8JW22Q9iZJV/HSjTtRE9W1KSckdUBncgghiygqyuFoq7bLnCQ0AMQhDtmN
KQpYZpMuwtvzkxkels+IMGBr2axw8a2eRlyr+tqhY10QtyVT8Z/AIZEDdQCA5LUQ
zhjaUZiKrZGHtF+dWKrTKGsqXuewMp0gCS8oPiThFyL6U0jVwglPDRdxtA54fvgZ
QMbP2ZOQx/O0pp98LQ2d7K615iagLEiq1/ARlTPUDJXayzNNLC9f/uN1cx/7ezSK
NQR9UiE/r6M1TWB+nZh5wrD2reYUOWTTOc1dJZZ+ptk44GhKmoo7eWDsgZPRdaPa
lGeeuIy0ASDpeupxK5GU6sh1jnL9dgEr2FwDZpzxy9tJyJ1OU4JX/euj/5JvGFL0
llwkWgmZev1ZrKM2o86Kz6bhNt3dW8nlb4+t8kWg7nyGguXrUmKQttoZKZ+E7+gD
wMJMowfFnBbVSBerS9WWSjQqGtHn97h+dRCInI/AkS130giijEhA/PashoCK19LZ
n+tjG7DNr8TDyWYnzfeQOVy8ogBPbAct0bf/O1xwLaDBx4svfNsKY416tvZfBd+4
x9VVWNkN568C4QN3m4f/sMKKxuX2w5/nkYXh/w43kRxX+x9tMfzIUm9FKeeKa3jX
r1JnbzQcF3SYi4zvouXlNzXbeXWP9LaN/rZTUhHGSqzBEl7hEqhwyH4Ds+wImXpJ
fsxbNGMATLla5WzVm6KuzAM2X1ekyFKX1nSgJWGdOoxfWft6s4ffg4msCZW+uVzI
lfm+7KW4+jDnWRgJ/XilQ8yTIppW2bWmb1F2ReVtGgCcbnhhH33kqNniwPMVuYKX
l9ICqHlR5ZRVxv3S1Gq5SS/vi/0EON09MQM9b7Arz36Bb/YOlVpOlA3OKgREr2JU
58LIFfmh2YPcdTQRGv5g3qI1g7z10ugjugzQSCdM9o8NkZS4zwaoQmITqm2klD79
BWSBtfyhLNlw74ZMyAmsTen9VMxh5ivwubkfospH2had/SnJbqtgta5pM6OvgCJg
+KCjQyjDbktppeFJazEGgywrEJe3qu4MJh5/cQXkTc3gK98olA2OEdHMk81toLQ3
b33TtMJcn9GDK8OXl/MU+liWUq2Z/DdukU+mFEF1yciqOxVCvQ/eflr8FnSzg38r
XhhwrotkdwVUWzPzKs+qfOjIXqR0VRPbf43t48cPkRGKr445ny+0HOXY4I1N7UTc
HypHqfFBoDrT3YJJY4otLoTqX0KL6f5saQX99HExyVMUr95loiVIRr6AG70WR6uj
OJi4RqqdAm9A7jmusJTOpI4lQLsGMrwvATK5zIUiaBu8uDnYoRKNNzHYLCf338Dj
alVpI6nNNqYRtmdHohOnJ31p/X4ADpJ4QedP/4WF3bk8abzxNLFQqIocwpn3oauE
gaoGlWQcSpssSRty/uwCAYM2cY0d5QHuqF257KW/3aZOMxSagXeolAkF2N3Rw3ke
ss4NMoKa/r0xmSEFtFma/EAWvM5P2iMlLWn3TQ1oex+QJ178IUYsxgzwUFrZVefB
fJJGQGlwOySFeGq/ILUodQl4bXVqH/ocDnr7yBcsqL8wveJ2sKRWnLfwaV6d0oy+
+eFTH1lB2yg0d0dR3b7u4LDDh08QDy+h5a6dqlhnQtlBYxBzla6Jd5WDG9RPw1Bn
OD5pbIHZvbSMrOedXUYURlNksCCwnhXaEXLnWlyWKTPru27ZYpW/BWHyc9E3C+/a
KpjzW7HxVRiyBbJ9ZHwLgGJ2+gu/kxKohVeV7o8r9tS+SQuPLqd5dK7eM4c7Xbzu
B4GLSKlTvFMNOd409hZACQpvSoeir8iHLlT7fce68Jr5tkyQTlMElus17wQT9C4P
obt+0g3ljRJcxugy+0UIbX7DvWs94EJCIX4TtoLoio2H12RqCwaXjvgAD0ZfR7u1
N9oNcJzCK0FqLNH+RFx7RGr/zZe8nUzmPDbyn1qKaNfRW6A2xbTjHQqwkgA4jTPD
FzoaHiDxp3Nkm3kKUC7v6IsTl1rN/3Z+fEFVYOX7eOjaFw63VNxz5qM4iHXvvzaw
Sdv6aPh+BDaAiiPGvjZYKijlOVcAJgJl8R6fwKFWNJkbmdjQhF2kQc05viAPA3ht
UF9IHP9RlmoIbYIIUQXt4WVm9eR2TRJwgQhg1ILNmrsTGQI+v/u5DsiyyNRjMQR/
v3aqeQkJPdzu243LkhcpXIVnO4p1As9TEmq+Xt9DO1domdrIQupLRk293g8Yn9fA
oj6hBZ3UOZu0bTILayKnMI9oBFc+79/5VMyv3Pr+RAurDSwPrAxf/AnhK9tx2cnQ
dKcEOblfm6PSz0rojjCaNcjUjnKBeiEq85k1cilMzvinAZCaZ0Km5XaGgVmIyQUL
sRjvM84AVPPoPO75KT1u3h0zty8zmN4M1PWXtSMqHZVz4b7c576Uc+rjHeA6LSOq
X0T4SCB8zWsCHg7i7rXVrAiczzPZYc0D5Y5BdDQHWhVPc8llI1Z4putDntTTB/St
9KHLpjO4j5E93GP9HUcb4sxey9EL+AksdYjWfGVXtkdFhQDbNrtaNyZb71mCxhkh
TYjT9+FyZVW+6Wlu8c8nAPyfvCxuIRh1FpHuFbOsh5zb7QqRSIUFmyoYTxcy21BQ
Qgp0cbRUpqKO4I+fqhY8tHBmRWczABS/CoOfcFuxWv5MhhwEsOzAP/FqApvjGWPG
2g5RuVolSUlWhnB/EC1lzN0XyNMzpmpDhlBs1tofsdTl6thfJjkpFF9HntcGvgGs
/D9703mZlpEVOghGESmo+8VqoQsp1B7o9XaVx/qRRZjMVmbZX6wPWlVeMVXODg+e
E9/8QplzpK4XqLNw7hMe59HtWArw7JU4zu8+FlLS0Ju6FHldTr3tuRhFofFbEx+7
C5LlxgTIRIUbSPuQBrxAVN0ahIkriFYqQKNAt+DXsUqSs2UyhrxKsXMSADzzY5F9
BU2DFGft9QQKxW7bdYjHF6tBOtLNrAA5GdaJQJFmsHOGjGkChnbNfzk4IntJo5So
JoS/EMwslz0r4Rpr21EyFBWR1QN7CRiVT87eEBTr7LeHQFh0IZCj+BBMYNFXzDbj
8SMnoQCdslKW+shp7SH3zgtaXCguApxe7oYYAKBe7ATe9Na2+uOVWGKS7ceiR04E
dJ4yBvjc3/ozIeIMUxTNwUEeBgKcPOTIbwQsPnF/UyXU47fsQ0OnDSfbTkpS99++
SqxYRV8PuReSL6l37rADUOpoDFoT2fkrCY3u9jrUMDu72S1k0SvN7kjDfa/zN63r
kDzDB5/AbUDKcA1Uhh3OSmdBBZXwNSqr3d+PORNL/2NX8gtdQZ3fbGNJgbVzfkMs
DFtvIDv9LCF+yyn+cOkCXvtZjBq3OV/33z1/ogKbTHTkibJn8v+GCX24IEzq7kVv
9w7dAGV8tzRbv+4cpm5zs0/2ycYsviVz+N/NCc1Y6HCygziF6ObZEbe3TnXoOxmI
9pxns6UlCHS+y47dUZWb/DSWeBQnAovFRFHR42loz3HIF3L4SF65uz0NTzAu6FKk
Aid0zowDRudzXqj+KfMTmGSSNrZ3Yx2CCCv1E/bRyi+D31G2KhR6HDff31FaRf2X
`protect END_PROTECTED
