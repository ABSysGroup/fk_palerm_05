`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gtRX29yGxUok5gMIXFvcf4dt9xLhNksccH5/R1Tb5tqPB/wOR3fV6I337BAQ+/vW
lR/Gd/bAqnj5bp5/AsADsSnfEOf67sN/uND1KOiEOyEkwtOlLG2Hl6MdCOJ/uVal
9NAiSS5oM0I/0VI7i6oyMjHG4Xstk31GrS98aLD6HVqqBA4YMsEPFmcqhV/lkoUy
HlXiwhcn7pG2YnkxC0gcsAjw3prwA+O/9cIXfdd79k+xPO+hmsKLSdsWUeouE+Us
CsDSLqX2IUAcVgIhyuRPanQuqKTbWizRScDH2JoPU/Vo8hq5yi7igtNsStWK2WJO
f2SoUjy1Gkqw2mC+S/zwn4Cvv+Zf+sLlxEEca4Y2Ctn5oHAUQyQ4Wcu+0p4BT61Z
3Qt1qAfisntsaVhHAn+SiW+e4WzzwyVE/j8XegaKDonBYEeIRsxtOmEOxcHKNSDj
6XgYRHk1DTv9KqHZ87/vyA==
`protect END_PROTECTED
