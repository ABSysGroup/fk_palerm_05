`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3T3pgS+uU39U9zwPueUt1E3ZQMhsiewcRtyiaMWIX3+8LnrqFVcs69kwH/tdQiut
89KAacGU3l0xa3zK9JYG+5nd0wEC+LtbpxgPmM4M0CeFVIOitCep8ubApdSRuqb9
p6ptvfSQqREAGRXtUjYCU+rKJ8TsOXnT7RTeFQ4y78lkUpYTP9UsqkCuGabgivLl
DBkKRCTWmQVFypZVfzPhM/j+pRAPUiHEPx498Tco9riGhUbtSLG8CuUb16RtvKCO
lAztPgY09QHoDxQjYgZHyHlCO3NNwzHzawd1nQvs4Rs2zvraPVoRBvE6vHU2S9Pd
2c+Z1e6P8Nnhs4Am9fMit8DgUGPJiEv5iUD2OsRiLGk5t1JT15/+2ms/5OSyDXw2
w7wb5+RIicPoHob/ckV9SIr4GEfuntrL98fUFgoJRt6+G592oUtBmI7JhUBNrBRr
px7zSx1vrDdMB9vLLoI2Hg9YvtO54FhBZW9mKcVRdcracHvqssxxOqWZY/9Vdx6f
RJWPu1yqylVAQPxNsULW1okGhKjdYmGzHHkV1LHXvZq9GSUhjjZuprqZruq4EN4Y
6WltM5sTBcMdf7A8XTzLZMMGoBDdcuRjpWw1Xxhl5TruKAF4XCf/5OeHAH3T53fq
STbsx0g8aQYv/FUlvKEJUJlh5qVnNdWCc0ISV/YNqh//S1qsVcZ2fqHOt1k0HgUx
bUWuDec2RLOprw297sgbYDZHsoOwsaq3RtInmlA/+rVOJsd/O4N+Vq36j9wCcJSR
KjeVJ/xdS32WFkS4NNpyikobrGMw1i0HGq4OUzeW4jIokRYxGUEzeHxZWEw6zWwP
1g9/0r3hk/i7xNMfsmT1TIoeBrokrg1+C4pHw/RSuW1qcbjhVFQeZJCRn7oVva0F
rRU4j+pwq8LrClBr2GJIWDJnxDEIFXlhbxTV2mBpKajvCMIeAWsyqR3TQ3tbjfSC
dem0ZJpabxlc6/PHnqxlwAhkz073Ycoa20XlkZuKfn3dcm05H2fr8rg0UOSVb11E
GHyvo1feNS+JoL6vEJg3wD42uE0Rz9DTkPVvimBKyzFv22LI/Xf4M/8l568okqSC
KchFYlNnOoNUN+vPoH9yjblGL/dZYK8hxmHmAsrsi82zbbz5BssZmYjKjwK4Q6bl
fSoyif6YqqHVtipZlM59eCzQRxv2O3io7CsBqJx5rOGX7bPUZpT7sbLnpj4Fj4Hi
RHuVA7kM3ahvkOSa1S+Iki1IvPzUecoDjKKM+mME9/W216Lf50lRHrOGOxqhyjkw
kLG4Q9dcOaWFprknEkNKfMkZiVV6kgpniQ5KqObL8qXYLwH9ZqyIOgZocschOw45
MeQ7qRzKMdgKFhu7SDoV2qmDAJXB/K7QmcVwi4JD0BbR0Wm67gjSkCQ2eZLs1ZvQ
6PPsOoPg2tLwQ2tHTJumGW38NM5AHy9REOrMkRy2D3j5shZHDWzvVZ/2yP22ArRU
pdgXSXaKNjCTr1KG57UiySSMJygH1imzOgMqGsQFSF//nRNNLWkmajzT8n8MRUa5
dXGm5dCYfHtn1IOQFO652MtiKAn+2+Vub+T7HQioXbQSoyGXCFu0JWw6NKm4wzGw
hi368F/mg+10XqI7wmFCGfR9eYaAXjA4nHHrPi92D7p6lKh+xh743pU3okXVXk5e
vO+L5RAOn2sm2nLH6Uow6UymLpNeyq6BmNuWk3zlHX2sWtMCYvi3eoNYCJXjcUiB
+kOX7RsHjXQEd+CEdz3ChP60Luac+oegcq7lGTjE4VWNd3h2LzAX+n0AmPu8YG0b
Ul/zMnVMyoRu4Q2Wt2IGzudxulLyvb2r8C6hRnQ0kZZmD2tdyUxYVKScfxVePmqT
ZdF0CeBCv5efy6mfwotJgxRq1+I16+qxGuuIm7OwqQSS/OtL5kI7jo0slRAVjTRl
X78htsmrKE+fV3Zv9Xv3xr0CLYAE/3u2ACT2Hiz8ZzAkZQZQXzMFmsgQ3xo0/uz7
dCDoCNyJGBHZHIPBvJX3n0XIikKOHIJeVfYVZcVmAGQ9YEaDSlbW8y/gxbEpBKM0
LaitqzqWhTzHONdHTm+cf6ANZmBHL/YBQAe0YV4MiELCWS31kQq+Ac6YeSTOQX6b
xb0K+N0gLub0TBDidGSRdnn5X6hOsAo83Jbtpd7q8/8WO//5uNeXpaSqEbbPX+Y0
TMYIZyP/TWKIglRUWvDMM24P3NjfUi6UhZyZnhBCfhtU/xqkLYgKYlDmXBexgYB7
bMgGMQ2ug1q1WnFebqlOWco0R4LPhzV3S6Kf86XjCKGgJHdh7k+3EsUgn+szHn0N
ADio/CGKh4S8Oq2Tihy/0scmppUL1MEZCJ2SiGIDLIJISh0ZD1bJ9OY8m2iQlBZc
CUgVK2t2EbfV2QGlfNKU/fnAuNk4+JiPrOoMArhwEuF2qk35vK86xnQ8ZIk8kYx2
cIL/yJtTl198VGHKJhKFQsZzo3BjczY/RmORHi6osM1Lu97yoanzMMVA9TSu/Ovh
9gMZ5gsF/PRW7kTyynbGw7f3zcZPeheyKSbCkCcz9cTq1bU5mpBrC3EHJ+Rzu+4c
kYNeDFcrWZ2lgEyFdFd1NMdZSdV85zZzKykuA/CvnGuEAZbFAE1hApzuPWEmXJ73
LfUR9b7hroX2f3vYBgotiQfFxUh7Lj/H3+IlOhmmr4xY3i+um9glI0GGCdylEaWr
IVgd0b/4N9Yh9U6mAu9LRuxwqat2CPi3pdbl3N87jA0IcczIB+H5z93MNz40dptz
2OrGf+F8KWMWf8qZkYo6Q4Q2IAxvDBRRxvtWNub638JL8aGZSd0M+MY2fa2OklkI
DcNw1ZT2ri0xvr3pwA31p5znOFfTuOcIKjkcR+yEoeRfi/s6qeMarVSiij2nPDGd
7lxUmeU7YAhFm3EZWrKtOV1ajKdYK1gNRfz1OxDFHwucusumw3En3DUT0frq5nNN
wF+gjTmEQFd5wmkcN2ADou9TSgSle209XIOHD/Rweq5jod5OA7UTzP83wupGjFzN
tyhT1cKFKV/CFUSvaHkdi4r7kTLazNrnMyScvvMXFWy5xaOidrSooNCN/7ZFvja3
r2OY9O214DHwR6iEsCHPnZDm56Moe9P+nF5XK6sSaLHHhLG3vUcVDnQw3Q0UsbNW
qd7kTcpAb7GcH8UqF9HP7vxBnrPRTMR/olFh/4i3oGS1emORTA4d6F3+Qh+JDY4r
eHVGDGnMN3n/2hhtDwg/bWEWBzfEfkY3w/MwP3NogfLY7xFPn4NU09aTtosrMV0y
ZyK3GfDjz4nxcUZRMKdOIGMRvtPQul2HuKr9h11wbR7j7JDaqakJ1gJ4/opE3tP2
qqCrnO5LfHgUXxzblaOBH3G/2YkMuls1LLEs0HqMtN1yX0ue6p2TDDyUi6S3OFof
vD5fxPC7LVIaRCSWQ9akSWuVYXwG5F5NKd1fgUEJmz+BSzd/OWjPHNx0Ul4gEs+P
0DKBLddVVQJiEBhnlkea20m6iSRozeeUjADBsCCeUq8mHT66lVA+8zye/YiLshtj
nAamQ6V+9F8M+w8fQeyapW33ASvBcPeYZxkTB22LFsEf1bRnghIqWgtcdI3P79KI
JP7h/vptGILtkquoQ1qXQSwN7Rns+SYtOBFO4xdB6iwIIxPED84BJCIhQE6ndzl1
L7JG8BeAlCRu5I2s4F+qgGnJEVgU112lvs9hEU0w2UtgxJUijBxaRQEfyY8nfdK4
+Q+IG+fRL8dc4G/moJ+aKb8X0g6UjAD0NUFtRVlfLZI09tcTz5UOGCHykPKyXjrZ
ri4hAdz4f4a0grD14X8Pea34cZCISMqNOxstX/1cYFV/wNFxMXZftEMTIN4JMSY4
dJ90t3abnQaIyRN7ovezpVIJM5+gwVOQFx1jc0eC1MX3hVSBU4nyR/L4vxoDZibj
GiNXCnlGbMxWahF6ytFuxg217F1802dRxmkI62JY8wCEE8v7S82yPA8CqYoBFWOz
bqssgCjH4/+RqvtX2CM/DkCE8h0wzvntPHZT+D98vG9kwUolvw56YMzh42spUTmb
ewSmc0LXwKqIFW3BuXYKQLw4NgE2SZRtANGayzXkc6o7fbDVj5W/vwj3Zzb1sfHx
OMQFhU6yTLbqfJsMuUNzafnEgDpXlx96W9oncd0rRddD/LxJWRnsp+BTn7EGc4QZ
/jF66VFT9xOywPnCLn73YOngcMofazbb4kMnguQCeKsMub/YglmesEGm9cvOB9r2
qfPqWFF44bFl8zbU6zJQcaARPla7aX8ipuZC77b7ybuVGu93gMYQBFFO9e38cuOO
H6htD+W4uMzc2HqF/oB72D+AeRu5N61MU6UWsWJTvTseKzRsT/A38jFEpoi0BZJm
8yV7f5x8OAXtrCPUKxzunPr2DPWbYz+TKoa6RuZFSwzJvlz+JKu5tNUREj77VpQk
5vt9kpcIXKHcd8+DWtDdqTOBViHvNvfd0oLr7+3EWc1XBVTSE3q7g1IDvII9kBB1
ZOeCMh8OkSgN0fQyHwzC9MGPveQOg4I8IkcKv2xp3iDD0SRP4u/rUNTgFbVvilD/
P5iJB5wJEXn09FngPQB6dYbd95al6f+YQ2B9V5L3MsrwHGWsa5MDxcaf5hlY50TI
bK1SSSrStGbh0XTcF7cmoTPTr6t2hIHqQqN1q4VolbPZFIUJ5Bo/0XUS13J6KbFO
9e1a+V9nAYJ69R93itjd4Tn842ayATqGLntgiQeYCjvw2gadoPi78GECqjqKiUnQ
u3OMURLcKUO0vrQ6EusBhGR/zfvMbdMPP8wDNXET+SyqVL8++NtjOocRLjW800uZ
jPjCYF325MLRWfNCEHVQzpoU3SOGT5QQqzpwBQOwMKvA6QEyqwQS8aJ25/FBhM92
Qp+twiEQbAFi3brvWYBNz4+4EHjsEwDYNQ+XchH448WbI/icfrHx+q1KLBZUbK/Q
BsrzfxfFr5cj24xDQvpKdf/jETDirPDbyEdwuvUKKK5ILEed/lP/y+1doHIQQM8H
t8WjcOS//5/CsRXJzUls4JAlvAYJyNW3w28gZ3gJ7ukXx7DRG+c9GtDSkbCPTnGo
jkI0iKJm2BRMPHUH1N5A9A==
`protect END_PROTECTED
