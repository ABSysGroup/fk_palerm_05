`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fOd3cHM41u583b+Pyaz5vXsToc8SY5lWz5Hck4VSC2ujuwmRg8c4yZvrRPK7sYkK
vu4hqRN4OkwWdsm7wglZcuR3nrp91v5M2EH6EFAvCJ/xKAp7dhKcsbSKe/WvZrOq
7BljJ1OyaAfwzFt3QF4NCVTJc5lDYjy5kOlFqIpPEZHAcYDpXiDJ+LP8JpTppFo2
CY7Kg5Zi7XHdr9AStcc97YxbVHuQ/nSEa4Ff7udInZ+dpgLJ6NsgQJniKOh6VkCg
TDII+o82q+l4lGC4mhkrbtnFy4WqfJK1pbmMnLrjhxJ6W4JbDcx3iVvyXu7X7auJ
E9b+OqMvAMXPQkXSqVtdblFucrhjiVYQL66kNRN9jAdsl5UjiYsqNeBrhUVn6fI9
wELzgR0VHHL2W2GGjWQofvnWuP5cAPg53wsCjz5eFAKvcqE+69U25ugGuYiBp8Ne
kCoQ21L7JpglG+9BKO9ZI+cON73bJyT+SYosBpIhsUOSUzPCOs6Mz2Pi/aGDWrhw
1mJuZ8cvK8L0/HkTGKV8Dobyt4Dz7slsUlgYHZqUdzlgqE7IruDIpFiig8KJpsle
65tR12CzbqNDpXHYm4iwWTdOpLhUbUh89+gd6silwcFCVCMzR5WkI7Qq5JcJATRT
JBUpU0Q/aNIKrny6vjuYeKQZA16ZEaP769ZeZdbk9NRApDIIGF8mveOh4z20TyIm
AAyb/6SgfVQX8C3NbRzUN1CJOos1FBc7y7JSILj/S7xgzawAbbdfT1sJswFRta8g
DUjKtKzqwGKzdiEokaXCqUxBCosY9tDez9Mw5ugctC+mB/cvsDCxSPfzEyi7s/if
XvQf1XcWrklccYNq+R55c82aK/jX7Y976JhRAjBfUT+WVwQeRyizpIu5Z9qO2H+T
`protect END_PROTECTED
