`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sjypfu4cdgeQb+8O2tlM2evHaxW/jA5m3hlI960md3VWoITWyDA5w4SCE81kYjeR
2EqVzmeylhMZlPD/lEy609cJxc2qDOcKc/okXqqxopHVVm707G/87CiloFNsWPAQ
yIZChZb/lYkIFvIvLRSTPpiXStIifxHNPO3lDs/MmifGxHBMeU8WOeU8UGos+Ek4
4ivUXgmdHEBsN1uelrRc3KBi+kdYkbV9aT+UD+a3ug3rx7HgswCm/yBCi5sMhHS/
uOg2UukzlQdX1Kig/hSpuipUAlVQFG2N+PGzl2Pye3E3oRGkLOLi0bu/AgvYw7SU
NGYPNgHlz9bAE8UjeJqe5U0KbTyzs+pMjlsV6ryumFXmizDiGBGjFlEA0GlbPDFB
Bc6FC9yx/mZkv84qeIqTA5+TBbaYLyq3lEuEXkRC3y/LuPO9EiAkoCf40zMw9A9T
fH9GFaAbEn/pFyrTgB7k8g==
`protect END_PROTECTED
