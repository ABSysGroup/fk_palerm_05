`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o9Od75E2zdgYXb0cOwxMb4prBG+Bh6bzjHaKEHRxtttlCOv1eOJffVZPBHey+NAj
d7PhRgJyoPMmI+kHQtUe9CoXpZqFh9JqEUAJp9/01pgmhV0jz6GeOKuug85fZgiQ
vEGtOvGERj3KsrjFjD7tNKIJ+nUmj5zeJuDVdnLrgWX1tZQ5gvEvdaslKWT15lj9
ApHlMWKFQsbeu0jSA/Sis3J97DRUFxA40a2sYEIb8yx5bdLDoUS0pRCcYss7Ggil
QMvszm41KaaDbKZMP+nE48aJChcF3KCfFp6m44fXYqkF3YISLaX54qfJRHJtQIB7
`protect END_PROTECTED
