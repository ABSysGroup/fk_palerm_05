`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LhCCi7Y+opjnKqJvXHVSNeJu+zOcZHLe7mamPGPR0eC80w5t8bi0j1SHPJDgelDO
qKrPR8vLGEhqA4bOd9HWANPmzYkakmWOHbiDjb4blO0+kaQzZhFh6hkNeG1dPAcG
15TMK13V5m7a85RQzFTkw7AKmcFtBPzAQJRPEFoD9u6Xp4ol3FnBFElxEV38VKg3
+6ySWnTNMYO1dGOqTl1G0jBEl/onUXxE7ttptN4F3S3Gl1y+N2/hT819bm+Eg4ga
j+E7u90IiBRRTG4YmcXhe2k0X/x668t4A8TuN0h9K6+Mebhmb/yFybbEq+XE+We2
6TmaDfPJf5OrozfJkGjX7FRWXO2bpq0SF5u45DmS244La5RSz3grJEUnJ2etLVQ6
xIHho2toDx9XioVj+8U2dcDMM3xMhNr7ZlcAe4xX8D5Q9zNY9S/hvimKLlFbvf0N
ziBzLqAOIdRbIdEdFDQvfjIZfquKNumMpljUMtqKBFAnJ9eOmjaCLgCOIovgROA0
Cgtcoev/o41OChdVmIJFvf64GgIl5SQE7d9TngXZjDkG6PnAI1yHJ+rjrxQzifOi
LgLz/nwNzIZs4fw7+qbUA4y1b3268wxjU7F981eJtY++xRhWAqREvaw8x5A+bWh1
LpFDVa9ooUYeoIZMgDSkZc8h9alAjtpingvRUadGJB8z8FRSHfT+s+2fJPT4bon0
dzMTH5I6aMYE0e32DAcelScgqSzVlY+0A/V9OemcMkROTyaDv/bNaMN0ycgGkzvx
/mls/Defh4Ori5b1lHGmKeGxyCOgPWimANSjWTIMI8XJ+DHrbrTHpVhu07v1NWnj
ndO6VdLgGMbDfPLbdYveLDKxfGxgNAuCC+7Ja91ip1wxFmaIpJJXH/wNPxYp/cw4
p8fX9wY50yxS9uNiQtzJqeiFaJQw4KxpcXmVWnb/XUlkeikgCoL8uZh+0PDLh2ia
iefpL/kEMLhIeisvEGA9ZNNIZ4TT4VrN8y0NnRwvTwYPFQxSfgN4DBGi/v13ZD3s
yRVuj5fiOP5wlcozQtyumcQqCplzerhboeC77EQCrVY2rJQa/hy9Qz8fHfKyX4Os
0+EVL+4Fk2EZtc889CCt8XmbuBu8N8RkmOcvfXYAu+L7cN67eJoqHVCJpFeEPkYG
RFMGhiTnTc/v1fi3KIlHAkjUL0oQqk4hmyzsltZHhilreXyrosUFy6sb7jRgnfyY
5pyPRFY9PhNZdSSYe/c5L8O1A2kbYHmiHdGItzf437uvx6RKsQf8+/qu0YZP6677
k+T5HQv+duG3/nl684sOWfuT1l955fNtN/yUYoyCfC2FiqOMAIiJstZ0vyk0Ob+a
xPUyvB0riQ750NNcnKR4lTT1SA9w06avCV06lYK5yapOCeSZtHSi7cylCrLh0L0G
zCWK6zYHZA3r3HWX7AKW9tMorY00pUAM23lunUBH8r4XXP0jxNSHkIIg6qBcc34V
/LvAR+IpInkiRMJfPwB+YA++Jk57dhxl2Obys7hnrWgAVVRP2kayS3TTKxZFOUki
75gIk9MeLQh2UaTROoHvXTeIE4dMBsk2KbqX/NXpSt+/1oKFuKMSUCl4ESlVNBBZ
2mDICtehZT16PQWaRtC3XZx2Y/Zgizm0EhLhogJNYOJkHaZYay2fg5YZjQ+66bpf
lEOcdhg14srOexTbNKB3ikW6NrMrBGga1g4BkbCjwAABaFw3IFWa2PQTgZAwY3lI
UO4pGrBIrw1HtnGXTs1O2DBf93GSka9AiOj6C2kxXmy07nTg5f7k3UUhV5Z4Trg8
WucqMHGTNx6XVMoit08TiuzJ3ZXerZtFNY6HQ5fvfsjNKsM0hnJiVKCmLtsQiFNc
XrsbnijrEU+7UpPiDiG5DLtsig1kQdpRFXJrcuNuuiMRp051u5E6f/EZQ/HTpFRc
SQU/tgULuleODHXFXA1bKHjVPhtPdsAHMm8iZyt1HBcsKU1oUa0cvxRl6SYlXdxL
TVmxmr9X74QKz5Hi/Hzr1FxPQzHOm66b+wJhSHp78JAVhZHlniUAg2B6jpD/bnGt
KdSqwIn16C6GJMQ9cvSV1CbksiHIKzAHCtVI7gt0BB2aDpMa4vFzV4YU+s5YrWJv
l0beOdqfhQmzNzI3g3gavIQzX6QWQUKmYDkmKmUhlHXQFzxmzGgh2Xcgw1sAPXwB
5G/VtGV6PGP/+kx5MB6nWs3RhVKuoRMaxF1uQjmsWbMG2Y6yJiQ8v5pzddaQwEkx
wKM/i1FBi2ZVotXvZ1WcQTv+lvqT1q5zDgn8gg5/9ml8xfMFJ0L5MNfg9lhNXP+m
d91u/kVnFL5X5dynNg9dWhl/eIouuNZquqpxmNn9yA30tlH8hoyOPNP0/2b1NvSn
kgk90wHWioV7M5xVK1tD4TzD4oivLuGUIxNTg3UoLNxnwFqdqWJYXo2U/zqkhjVK
NEaSPbdJUUB3h/k/z0X6Cg==
`protect END_PROTECTED
