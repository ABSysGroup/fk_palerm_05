`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YHKOLqrbAOZbmgiZd6iuRLPQRiL3887ZlwbEdPBHs9fexO6hJXgVKQSql35mMnkH
2YfROzW23HlGmmpfcWPwrqgq8uGjoXqguBHa4iKqIqmxsjucLwqUqUfhX8KbY9A9
5l1IP3YOHKgK03KcDMRJbMi3m/eaGpPx+LUFvIVRZ5UwDWq0cpOfjbBRrMmwg3S+
gPVeeiNUfBS9sZlNo+9cTUfDKydGDuvSpbN1wiCNBjyMstwInGdhGcfl4NfMJHvT
DUGCyxFV/H59QonNEUT6QilMKzbUFi/Cb/tpczmjF7090TJISlAkcdJd8KpRitWE
7NELIhKISKmNO+qksM+3/bFJPRT/kauxGK8Blb47/3schP7MWW2XTm2JQ+1Au0Gx
2IfqeoQSO6h0cQbzRHL2vdEAOm+SpuggJJA0+KJ0U2wGrAANYd/iLKytI0n9XRRM
evYE18IskpBg7W+PDUDGS7cWlSxeFebUg9I/SSgWSJlevv2Gpvhn6n1NiNuUijIg
XcZ8oSoVsYPMy/0FKZSVgW4eb2xLA3PblMHUNwwLdWGyj7lteM74IXcVDE3wDayd
3NNJgBU1oFzKAQGMJqDAXFBmVcHnGjV0Zq9GOIkO/yL0icCzQH3uTkB+AVMUr+SU
KsqYYMDj3uDe+1AhAp+kIfCdyhMDqlxBdGzg2+HAoQwZCmwn+fwAwKg73kSTEP/e
PebrjlyJv3pfQY1qIdFPm8fmlqakxsx9OGvUhKcZgoxcZjTHSH8NWIQeuKSxBfZR
iLdbFtYL3yeQ/Y0gP2bh44GArZBFvKOXJvwXsq+YL06qlrB1PBlaFF8emR/QoOo3
+jWc3omx8HGjD+QM+nTnCToQC1KhRytVtdUB3niJssE=
`protect END_PROTECTED
