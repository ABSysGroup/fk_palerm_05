`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
43SkQpyvl4/7EuCFGJZhgNnO4exnCBA/9sHI8AZM8SrassGGu1T7Dit2gP0NpipR
gkhIgH9petEJTLBsqjQjfW6zVJsLGsEmNgEr6060p/BacBLOLLnXkaq1MZOLNFuY
hAX/qvTWIe7dIeoIErGbWuIWCxkaaAv/UrywAQy3jsfcaw4ThzuS4qFNHUWX1Q5L
pQLAX3x80LWe/2g8wu2S96maXrWBwuVQIywbbKcZkaoxX/19x+l8aEzNZT78Fv2z
`protect END_PROTECTED
