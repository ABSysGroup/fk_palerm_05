`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yu7qGwXhU/AI0YjbC8a7j197z0GKMuVBsySOzmg6V2VtnAQ6hoP70Jh5wz0F3yaW
Lm/05XKfYgUJRBfIJiaPp4bgGOvUGj2pH2zL9rar1msKaTvcBUtHAGOB4G6S/Jjy
pJ+RYOPcOVH7MISHyVtqMCmxTr0GJ96J1rfguUlCxrt6wdaroTzbt3KaSrIerSpC
T5XCguitRxs+WcC5+4i3e+sgINgzkZiXwWhCBD6kDZ2c6sZB6QhzAk1dHvrWuQJe
XFVH23xVPpwPd7wTOtEw5P+e4hq6eiGbCIBb5qcm8cRYUz3esrdTOTtAHwclkb7X
QabVDiFrsqWhudyuCgkMFJg1nYlB5BefbhXr0SWbuZtscxuPHk/pCA0EkFpKFzEE
usDOUwTJYmFAhvMEkwrJLnFcm0qoc6flgXqHWtjnn+lVsJuWY2ssdFJCrYaZu157
FrZRdY+llg8UR+YhadSqUnbiKMCbXkxRTD5DiMSWv4ZRY3WKYbcBUFwh7ejMsTBe
iG+sxqIp3J2HbC373kuUPcb8cx2Z8DbN517gbqQcqVc1rEbtPj7d4dKAC36v5V4f
5hwXZ2IZsOe8y9G++6/AfDnzu/M63CJ6sbgg/us+VnTynIsMegEgmQFqKHdfs6Ul
2KTW6fvupqv4uCSVp0k2SILroWm4PCwWYm4eRM5SNKvWLSWdPt18hUamjtEWakuz
cTIAmcFPV6u05me13SHL14BxLB+PkzYudvbH3+LayN/C4nfsnShU1X355LeWfHbF
Bp+hhqpYytqnChY4/1xi2oOeOccPhBH1SurtR0WC15n5Cmr59qNuW+YRz9lswJhP
yvRh4b3GhzaN1Cxw57vD3v67QfHNn8SQK7GVH6TUIX1MeeEnHRYgezobEAUGcq0Y
Efbqh3uaJo7HM+kfzQsOY7am2g6fVvYDR8vqCKHWQigd8AmXgLtKhmqKlHTD9KQB
RmuzKT/aRj3nNst//d0Lv06z88/uxTFYQCvWPrqLu+2aM/KPBWUqrzjesOET64+t
kiaMfHrABKr8DuHksaK/+plkP9uQ8wq4YgSfhY9X4XGhVmObAR5zEeDzhbkGutvX
hKDyF4Zzv93EMZVFh95tredCOPV91wrSBZ2UJbcO79NdbpOxDe0LnYlfOoWq6Pxr
hSl7pvrHi0Pg8V6pfr4FXRSJ+lpwIjL70bqdMF2TSinDPh8Ks1j1Pgb69h0K/sCa
G352ktMbbNoqVy5FomiYEZ+3Yp6OMvkoow4ozaS22NKcfkAsC1XjDygcsQfZRPtg
iUeccSjOoFge8EGnV20vY/c+94v8lUsDLc/Or12ExfiLaldALZTnp0tEGtrzG9Yc
ZYLy0dHCjJ1tIF/cNBqTZWcm/QV1uQLnbJqD4iRriKw8YdYLV2NrYL0TtpRhDex4
Ha6GLWLn93O14lMIcvGgZJB13ihGc3gEnL7gwcMiC11vCaw7hJdYfJUlJtDztqx0
ln9LR29aPozS3iDKR8l19sXssQ5g3K7xbad+6irMK1AVAhmmjQg1hXuUndg3OjE2
Vm/5rHqITQInJMsWfqIBcgHG5uI5wIuWf7E0kBerDsmnsk+mZ4vToEoR2KavA5Fm
q9GiZRLCPo//+euM47y915bFtC7DwqGUfNUUXkN5A73XGQj/4TOlh9vuLnjQO9F0
NhjquVAONUhd82IpAvLOvp/dfxyNMAyp2oT8lass2Nn5ASmV7uhuKH1MI/s0cIt2
Y3Mz/IwZWL8N1hqVCRgMCAUrpWILdkoSnFu082qy0pNwH7cejevQM7kd1LgBQgGV
5wA1PcRvpjJOVbaFFQ8K3vLRWlGlhn0Y5VUMIvrWS4kI0zeYKgxdt+RrnnSwwzsI
nwykLzq+9zOg6fhF4bakHa+xBnc4ZlPS4eDzM7eNW620x0sv9tpQJ6/JO9HJdvFQ
0lCOH+CMqgG2+2vMqnfsKDIhf7ESLQUfC2/CNpjY9DKCi7qmumckSNMjSqgBDhrb
yRJHujloc5vEYyUN9GdPoriFTzW2WZztZBRoUpGc5Hq24nw6SIfhO4Rs93ZTaiqZ
bpJzHsOko3YT0dtNYhAJ2/sG15oDFM4lyPcZhdYwJMUCBoIoz5sCqBJKodPIz0Hk
/qXtESsahEY5jVQBmirFM0GG4N/X3eflEi+eF0KlBkash99JZmM79yds4hg7X9yo
y8yylrwn2lHaL9FPEwa+1tHd+Eo1vHrTnLSpRjy+ou+XyNRTPA7wShLZt0USv2PX
mFNUlnhziL5luL5iYU7uzbsz3JVjwLF82bOlVJ5+MLcXc3hgW86xzgrHOyWIG5ng
bAUqri1nxGYEhKwf7zlRq/E+WFkiaRe466QCeZ4p3deC5xkjiVHHIoG6YnieKpK8
9L3V4Y2qB5LT8ZKMM/qUGkRh0I4m2LdNWYT3EUAEDsgs+WhVQ2iQVs7e3A50b13n
uF0irG4fmK2PHMw4CN+nSu/FVsp102wWyINCWeral6dhJmqsoBFTY3zR+PgeRWQj
CWQvASUezzshUBQQsETnDHmncdjKvo1CHu9NXhuMXqEqfxoPF4ismYh5qcZBh3Zm
D50dqNGqc4lynVJCryVgbHo7FFC3hbomfTB+jtT/Gu1a4+6Jpaf4R0dqNwWi2N3p
stXVkuz24vJX0NeOS2nn/qNib8x3bzcho5SVJJA4hpAZjG+4H0WLqueVNT9qxLWi
WdY2S6LbwnWxcjhvgyrTkVCi2MQr7OMX2Qy4prSZoZbxRX/iefph7BdVAzQtLnrq
xMgZpNmMst6K1jzv7TWx7/d1k/5/hNRpFPNuNrlZqczoeauUqtyFrcXdi5KPJ2Hj
Ddy2XTh78SsqbKDyogVJpE2qI4MtJV+ITz6HoxlaZQaz4siM/6YmTaaLXprXnxDP
v9vIY4vKYYXyIRjZj9sQXeC2HDXQmQ/rntWuFcst2F2l4DeRew9VcfuQ5mAQmlDZ
col/cLuMjO9S8TG0avd2ADP+yodnMQ1jw9+JV3pvl5McNaGjyG9UbptP39FCpDpk
37JFsEnPhKixbXeGmRuzzd9ivEFecoIZeLXQkkERbiKbMioGRZoJQH+D0K+TcM31
wtaoFTo9oZGWIOE7l5xVRRdsjH/h4CmKeWnZ3Uf787KX3SFSkYtkl/c1I0TVmG75
mE0sFsSZ09w+rG0nkqHflTzPXRtu0MvE0qOLMDpsxzKmXHYrh5Qe83MdF+fRKQK5
vVeDQGwMxh5j0OsZgPO9JD8cDtnrawL7pplcsOAeS+BfEmhNrkLY0Nn3lJ8fXjLj
lgQ34rWRKfO30h4njHo8s74x6HvpqH2VjvCTzPiRKlqJtlBujnhrekFlqe3+W269
`protect END_PROTECTED
