`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cmh5Sm1qAuUQtS7fzqpJFhwLzHq3GUkoyC3kowgC/bxiW79RwxIiESOyWOyRp9JY
zYgHsHWmsU477e6hHtlutew3rXwTslKqfRMZjvg2dn1S7AcjZPDHbXrczrvj/IyJ
7y2jsXaY1H6XTYRdlmo4l37nNs+MIs50pnhOHO37iZKv8WN4rt1kz1HUCxXTI2Mr
MThru0qyQNrI6Yw0nWdIYokHeAJvOf8Krui5gcUd7IiNj463GlpqONsIBpfku4Im
0FaWEfwQzlxs/9p7csTGIqpKRfG+cZAiKM3/MTbqIU9pFI+O+KqJjq6YZIBydGm1
35i+BfMPTgbsUuP+3jESBB2PJbB/fA623Vaz+f7fZeb23y18SPgG+6bAQ7kkz9Ai
qqLA6OUF2iTMZfffQm5xog+0sVL9NJVKV/jmwokw1bCf+Hz8HPc8SVeYt53bQ8T4
jEVssQd3qdXO+D5S6KCxgq2yMs6eygM8/timUkhYlo1LNq3OTr2GuGwHw3xYVuxQ
7TOgxbpEjQLMUD9T5hvtG0rwQiGvgi8K9VRwRZ1/mDWFBfRaupezmiZbCh15RetV
`protect END_PROTECTED
