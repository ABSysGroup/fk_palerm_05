`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LRm8dfAdH+fFcvjbyAmaupZEymAHXScX0Sf5+v4QGi6Vr9fp2fZ1aRuMKEmXosdU
KC7fBQMVEk7v/p4NzUjJPa7gaLCl4C+CyDZOt7BQGvf8sHAm+cRd+fzpR/kP5bGZ
8nuwczW8OKKXraNZI4L5jDq0FqpEaQ/58qUYFB/FTjWtZnXpOD04A7/TiPpnc9em
d3Y3d/A+bvX6mZVfdx3kGuVbNnu0QX/NJrEyhrHB3lNkO9osGB8pb1GPOjOxN1Gm
2+6tgFf+TjmaDSWCVqgxJUzQ0GWHYL5sOzfWUsHgm/5nhtUwAAIJBPiK6dPWaiDS
WQdrmLpnFLxPwuK/6isQLCKZlNI5jJALzRoJV8E1vMdMx6C9FPcV1PkzYKkPlvwf
W0AWDHFd0PhPVOTeKa3UbY2DLYjwJNs6vu9A27U+8JjfUwYBkAS8x7NC3M5IWO11
uBQk7VGlItSEqSoKuyDk2TDp2Q30Bk5/bPNHp0gHWMc=
`protect END_PROTECTED
