`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LocI0nyJq0rlAPgze9PcQCTJWz8hNr6/yLe9SgJsuBJqsQX5SA7txlvuozCyBcZE
N6GXPPMmUN4Xaejr3zKL+Kgc/BcpSk1sjd5ACdnlan2y5CtZJWGYLb4aUpXiqZFx
MkrTgZlyaJleRVqnX5Ble5+iE99t7LVLTcFmzCVw8ANhSz7wCmBbCm6hkKd50t/5
WGB5JUpAiW6ZoXqmiWUENKlIURHKCccoVfXt4pw5xPjUmb9og/6mnQkfODWfmd+b
QvUZjnOoVgvfpCmZ/Sgc2wWmJpv//Hp97/eDRUiqzVQ+WlD1WuMPgW+4FXyBMIR+
BcNk/IBEDB2r4qdOiuUNHLAtOzhFqOIzz5TUb8SM3DEmgCiI5lSw9UdfnczxpbCL
K5Y45zRlmWY5XGu+opagwHWT4qvHKYKkrTxjf06jTfoekUxAjwoN4GditOrIpCPo
zI1CB4bp76gdFdpInqKuPagd/Q3Y+Wp6H/WerUWMp4LgC6+N61pLLVhTyRVU0QeY
BH5D7mqwB4By1V2jFenG+lsp8WEa7MedSRYvwp8sVksw7Cxh5T/Ob7W7E5I4cwxw
Kcr2vOMVfF6PNE3WfMcpNTBUlcdDy9Qx4s+qfy9KJgnCjlGmVos7OuVEqYax+36N
nTSab6ISgG1HcsruvZWRSXzrVpLuLoaROvw3UuwSaZwOehtsXRrBMZa5ENckomeh
pCXYGRW7V+o6l+DWZBWiCfv7Jzfw8/rKSdt6z0CB2NHawCCH3v3qBS3feuDJrN/m
dyyQhOY98jLsiyrjupuvxtiVRSNXrM82TUzL2seVEZI2GqEbIKCBHwhLc28sRo0q
CYVwIxJ+opsFUuO1xEPwy7E7ssTOdpDsU+2454j59UqIgv16oaD8AOx4YyXnbKGE
NlXzlJGGWEtIZBSmGLVf/4xL4FUC2wcQib+lfw0Y/y2C4cE/r1bc8EycgWIZRAW4
G32UvhdZnIV5XEg0rEURE88T5hgzFfOer+IoQTxfs3P26aQhXU9I5lFf80AcNogV
XjJ+gdbtITv7RS54UzLIWdtGOpeaQtllo6lTX8+OHepCX7aQle8axEkp2PcPJ4oz
yBsV1cUXddx0NLOcpmsACziF1TT5jecL+L0zIHCTo3O5kkxqK500J7ucdnAeoOZ8
ACuZfKvkFXqsQftrKtLMkSN/584V7oblWzXJyBHwURzEaiAvMkKsDe3UgwTyT8Ui
Iy3pyTSlZL93V+ahT4O65I5BkxRTwOYriSTzHMpHE8dNn/YjnHWGoL7VOJ+8YNr9
7IcaJjkGDmKWRpwpQXYLwnaxftKLUUj/c2kwBYXITu3k+MN+yfjnLh6OY8oNZpy/
J691b1kRKNjnAOREs12IDhvt279BTYH77L6mXHk8feCxuQxcJhkTcPo2WTtTGf+g
w/LurYgCJ75CLylY+Rf5ppRW1GTUdSeLMRoxw3Sc0EsWhbK5B4vpErtjC08atou6
uhKHApVB1AwG/i2LQc9CZ0P0CzHu+zbfWOkN2HrMrsqwbkL85VBlAWUTwlG9bFaR
jbXqFVDz3d1aT1xeOQWReWKvhBMD2QPWl+hOejhXX+ctcRSFzMVP5l8YzetpvgHL
NDZ30Kwvv5EvMsScDL53T/MKVUEwuq9oyI3/+uGtWLphqJWmDib8GDljKegDUg29
BLV1g5jk3XeJlAsDxmqQun+qH1wfU0Fa+IX66Gh2eOkLgsIpTLi5H8nSbZEIOmWo
j+tYvj58GFzDdNwrb7n5RpYrGAastbzsLe+bPX+2azZNaAW1aGTqjmaKyz1HpbR6
AfmWWC3KDWrqZYZBNDt2TfjJUqN8khEewD9Dl25EE5QAaFEHnOEJqaYNJ/4smHOZ
FDR/WdrR8Rv4damBnf+uTBFac9B1jH6aH7MQgJ7Gc4RIlWOGpp2wfOZHIvnUTkwM
rITFp7+QMXNQuiuSvZH5/5j2okSJN58vQQ8uhZ1M3s1ZML8bwrz+clUCIsNlU26A
0r+4RxUBPt5O7rv+bsg8c+AzHgFKUZxVnZNaVl7qJgMWGVarFeakvw8M80vY5G+p
VLhxkHGsMetQ4/4heub8+BZEsS0+Sif7FvTesuP48BuyNAohl4HvMPqL+HqyQvJz
edj1nkBWIKBLdIcXIc86xeqcoyi895+fuo0I/TvJRXsiLfEWh+f2b1awT8AbFvd8
TrsAR8s61nU8CUON1OZzLqUJHBcs1JyuwE892qGu/93wcTJe5b2UwZB8Nxk2Xm5T
yqf5U7Tdiy2bT+r19vDrcEGN6mLR2LyUbV1+byaICBUY5/GNZGkenh1w2XkSgl4b
kHeJKyAFq0lFpVh6Qve5l1ATajkCAjclnb7lFdXd7941SlocNi+90kgUWEa3+OJP
3Kgp0gfUxpPkDnqN/AXXdjgSwCO3f8HvbCM0Rz3/KCNGjH82MpSyBnepBNbdIRKP
qBkaqAs0kj92cSEmVw+ivNRMM4jSbAD6+lf3djBwEzC6smMeoH+I7dVAsewn5yzr
vVcXt7j2VSxSKZogYlAVoOnWLMQpDsl2+DonFkl9ti937X+CvVtkTcDV328ZuTuw
+pqUhU9lzZt5ZbXznTZv8PwbNGzyRUlgcR9i4aR3cbo+DWkCzSq5HpDvlNXlsb/4
g/2KYRGvUvrLesPk2TWthG02J9NHaDmz4H90hzcGu6DYuqUMVtItdDJYrw67fBQY
n1ttjQf5kOehAQ4dph2Cnx5AnS2Tw75C5Z1O6LVRwPYBsHPgar8cDOaAnbYySWEr
3T8YDeSfZeKwQ0WY5/jcvoA7QTv/uOtubxvDtaP5+7iQ3qQLQvamJ0fywT3EI8+Y
`protect END_PROTECTED
