`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Ai9sB0FnhuePyYrI6o8FAa42dGqy3pr8Uq6975yIJqKH7xivaa/EAZ25m2Id5B7
WGAC8f8XkRJlueZ2v5htRnWCaeceqXY0nvDbbqOgyVMkiLyC8Pp6XhQnKgazSmVa
KoHRaSe/PA44dpkvqK0gOszQ8ot6l0MlHQUU8CQWqu69eDg4r4AQ0rIRm94d7xKb
SFmaaqd1hMitHzJlPKqYUwTFw106KWZsvijMHCWO8+2B8JYJdabe8j7IFY5qM7Kr
vIMKUIMigNPjWu8q4c3DmeZbDVzJmfI2fY8RDnxqHiY6K+bFSGmgty0K+Ric37RV
VTrATctnmpcRDyVQrAF/v7Klfk9vGX4BYFaim3Hn+k35FBVAieL4hcb+OhizTIpu
Zhgr+BB8iY46+tp6qoq48jxIu/bLlKjox9AA6qei9zw68abDEAEVYUetScZm6Sv3
rypeAx+mg30VskVTDBSaRA==
`protect END_PROTECTED
