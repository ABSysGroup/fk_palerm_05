`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1I1BgkgghNj0PZChHLpj+p6aPc6w+a7+W4JszrJSoaDJjbs7PnWd50B9wCHvSe2d
A+9wmwl7Lb+WVf7uKDYCHoLL24nw9QbUyMO33nJQyj7ug0Ap7PKEJtFTzjd0dnfm
Q+hr3vlgYZW7H5oojADKNuUwyI87Ry7s7vUjGR5Zyri9s1KZ5aILk009hddWjoeF
WlL1JnQGY5KtglRR2YCFtCil+WbSxY4dDQzQnjQVzOAA9XH95koJniKb39U/wfZu
jx+wBIidrffy9GM0RKGb5kAekKduq0q4U/+E6LBoBcZMRY8VRC9ibDK+kwPgogbO
`protect END_PROTECTED
