`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NHhmkfo54pXt9MicQsFTQJ4KTwPMJ6V/Mk2dXQtf2c+JbmubB9JJqU8ThYAmJDm4
Pwr4s+G512wTGy87QGct0np+nz5rpF8yyy/eR7AwlVPLsTsJ8jhC3kcF64CKamdd
oMi7cFeEo+teSOHAr1xCqTr/4PPoRLvwXvwyItwEXXH4iRMrXRXx/f/MP4ci2Uvg
07rLpyeEYadmOp+7oZFeEg0g4UubOR0eR2Z0sXvxEBfZwfwF8HtJ/30w00nCwv15
DG4xj6dwMrlrKIS0WqCCoJMDtPgJC7OznWw1X6qvEoUCFeXfqBuAKFc5yZA0YxuB
tFuX0lTZ90S5y4qHKeV1C2YVbJ6HVlWhffL/RgRDkb5EVK5wuTG4oVi+lZSHvJZu
9AquYN5t7vdiQ003NvPNK4NmqcM09eoMxxJr2k/WX3OY8sPkO78CMk3CV5+RNy0U
F/XEy2gsbIcUD8Od6FHBIsXAGWTqwHUyRNWaXWf3VUM77aceRhbakMp8Lt20q1uu
rIxB2XHAPBB2VhNR8QcIML9HmGt+cYekmrMzlKSLqzz9EFdoAJJRXfAnkBg2hYt3
9wI5iLaqtKqdZ6GU6TzlYg==
`protect END_PROTECTED
