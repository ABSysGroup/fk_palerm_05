`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2bCIGqXVbQ03xP76Rbi1fUwdtd812hu8mrLkLHNHdJYip3L1X64MRL8mywj+z9GC
l9CZ6xyF5mD2s0LR9fQKyWCoMZcMF9HrS0kpuxR+JCMiWZJHpRlpIUl5/Qo5M1fk
g8ZQhZWnuBJN2l0hLtQCmkSJzJMtWArg5xZ8F+6cb+Hd4kslbdOPnESzM5YE7hRQ
eXNh6X6BD4lOBYDGQ5qQTTAkZmXa8rWoMLnvY1QN06wrbHT20FyJwrGtHzre463v
e8qcz6X/uCP3QBqGPPWs9vOhW/+cYLrud0+7ZGYDE4MHLLpJmkdy8KVwERRjnxXH
ZE8DtPgmLPvq7xnl+Pc1zN/ciItTPmxDOdxVW4SWb7voQitpux8tniWPgpivhwTG
lnlgJ3p8w83ewVFGjmoih8zrRe3EyMEzSojK+jCiAkBvmMcxu/uzCqVqLkMBrcAA
L6hjlDf+V7V3MxiD5ya+0OdxX3ZK/2Av1yp7J+J57IqWTJ+dozf2wqsfWxDAqoRC
yB9TPZ3J4YF13K8RO8MokIaO6FMGRmI5UMZSXuGBa2WLA5vVvDfbZmCMpZlYfaw+
/diDniQJPAncr4GbzR5msQof8m3kQxTcJpLvXj2WWrRAURJMdWfz2YacYwJfyiPr
z0U5nLWRopkUxqHmgCPPieUnzuK3uidYRNZUhlU6HiAqSchYRD7u97ZJXCwgBnde
9Za14oF7Z8CUhnyYJ3nVyCbC/769QURalqHHQBgJY8w+UPmhUgH4T3k9/jt7oRNf
D0g9wyZxJxvujco7d22uLDQkQg9Uy5QKvljX2JhWygaQG+VQn5ZyT9T0GMVx3jDU
p/ymP9rFF/Dtk1+XeMGTxdm+pyxYXodPzSxyZJbtHS2UMZ9W3wJhPpA0zTqkgNz9
j2Tchg56YZ0LZzy/cXo+U7Cv2PsrS3jkd3+LO2O9JGmuN7ESKXlbjUfGIvctZbfN
9rX3Btt9sqXcpU7uRwJMn8L9eaghXVjSExovCDQAHJpuWS98AStgSwW1mRzcoVGV
4ptTuwe0YYTDb/ToNeT9lzkdX2oQCZ44wMFg8TxxPeLmhUqWHCaBvaXmPYW9nHYM
3BhkDbrUziSbS7PkIV9qJw==
`protect END_PROTECTED
