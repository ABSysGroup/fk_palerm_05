`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D1cubzVRhvo4vhs8pCPXxzPEykL9j9xKEmeAvRHS/oJIOS823VPeLD5BOG33UNUq
skOyIIV0WwTBBMH1XIthBrUoqXC8YN+GsgihHaceYkGBBpX5Enwse9Rddf8lXEvG
+SUzkDuaqfEXFlZOMcy27lR+jqLShTMIaPGXz2vfWrYCOJCnfrkKM8cjxlGr/S57
LLBoTr+Md5gTMWP54D6RHpQguRY04APjeyvVwvBUDR1xeOJsjHQLnw2DcQmG/bWZ
DGsSBhU5fPa8b6BdCMVEQGnxaNeRG0+5b0k8eT8M52tp/bBqI9E88mJ+OX964bJB
anPRzRhI5DbelJL6JZSS6QPrgitIpI63BzrcCKKb3qxbivMmc1IlQx0GuCf7bLmw
2vvUBzU+uU/8N/wyKrcYMFSJ9k8zOhhkIUVQ1WeELKmTisTvsxgb33cMacmPoExe
53OXyttl3Jeaqj6bp1Dbp+jxi9QieBZ2v65oJkdAuVhx/P2WPv5JoLEhEiontCri
+wmKhvEkjP6rJ3MRn0XdQXOvZ7JvZ1W7cgg35xys6vuWdivQejH55vFReU5Rajqn
lFHHbZpn/XE3GphJFQjFLsCaT6/4fJD/QJaatDP/1RXPneLJlFqG8y6BcYe/tHVj
Sci3wwDqC8BbuHpAXzTZWxZDqTVQaN1ZvSna8tBfuGs=
`protect END_PROTECTED
