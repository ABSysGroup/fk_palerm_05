`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nMFWU4h/z7W+YJTIe6fAiDRY5dDnUEhNBOhVUxf6pa3RmzdUYcIxVMzA1hYlwVy4
KbdGFZV9V2o3uFGGq4abTDRCEafOx4ZFSY3mr2GTHG+NAevoFz6ijq7vK0lT8YMo
DZfHTz/ngsXnNbriJqD5ftjFfhIQglFJiIwhVpsP7uWCViqi/x7L/4VrlgCHQezV
adtC9G51fCCkznjnOORSeksEu63ardx6TLxIBPVhr2tnPMXPqybYOXN3yf7LpT3Y
l39VmKoSiTUyhkxP1vCMfPwX45s4iPcMeP7KZCSQO2gUpGaeawR4991Rv7BAY6oh
hO0K6vHC6Ez35lVSvjzS7A==
`protect END_PROTECTED
