`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UqQTzORV+ad2PdhyGST8H8MHj7yDBnCPsldW+vOT0htM+/hYRxmWnimiLRH1CIBf
DVZ/TiJUrL94gPLAa8iwyqcCgE0P23/8EvVnbGRJBq/+v/vVX8Vs6kEG6ABDOBq5
hMUC4e0CvjYfScJJRPvGceu8yORkjTOgd11b+rcWPd1ggqW1nc0Iq5d13bCBAAWy
podfBjiiRVLcp/4hJhx7idZ0mIt5MU4LlU4vqghB3qfCVAtAN8GHa1KxOO0VIr3P
J4uS8aVVBj/iSUdc4KwIN21FbvP3Z0NtoE5j+AV8Rf7dCuiQYM7SUzrEUNVAF8Cu
H0Fo6Yl3vorjVpOozY5GGQbBvTpCItMCOMe5CigSuWtbks0spTX+ri2xvHCJi4OE
UIaDuJ8dMjxeMjvl/LIjjM9gv4sM+b5Mnb6KbuMLndye1O9tBEv3f4i+yL+EB46c
Q8Bj9kMF7iFMzB4KtmrpfTA84ZLUbM+rwx33lAiB5E7fQ+mvs3omF/lWfn3hvYs+
f4CACyJx7N0VfNwzcZcMVVjToYPV6WAD19Oq+rrXI4pzlUsxlFI6z1d5BZqpPRgh
MTuXDZUGXig+yTVgcf/fHCdlAjGg9Y+U8TnyqxAHKIPSEtFC38oTHbd996iKUCQy
cMhA3nQKWsfkemT5RRGTb/12G+zRU2UuIXzk6g2goK8IxtekHCrYaqZgqQEmFALd
CBWYuqbGVgS+vbF0hN2W4CHIyYBwVSGXFmjmgrt3i8Tm+TNJnlkge2i6UnGM53Sd
zwVDvdDceGD7WA4haHSQb8+WUM8jlfR8dFQZxMlz7LZTc7wSR3yNMwV2oSxpP3yw
RWHnnO+VD3Ck6WGRFq4/qIQfqAxGATJJjpFxWzSztxMeH6PDT9mwSjy3k0qg1l8l
8xhILCtLQFYaT3EptiE3AU3FfNdB9OTZJLZvXc58KeOKA21EZBVvwedU1BiyBIJe
mIREGDlm/KTvaSq7LnCdJYS31xdqtS9/QTDK1l7eOhQWHFoZKe4m17tgOvd5dl1X
XYhXpG9vWV6i8G/3HmWwaMwQyi9qwNLwPQbuP6R1eE2lRVwpQFzyXfUHXYIP1GoL
lADdYJyGOciEm8G+yG2MTLgw+saz4tYOv0TepdlD7wipjz3Y68AbO+frs4mu58u+
un2ON0ZoiAyUqCSfgk9ONFmEhqn+yaQSCG015vBuTn/MtzXs+ijf47pHU171JK13
FdvcZh/eY7EA/onsfcxK6Y8yWEaUFlSmuG4gUKAN/uHgypq3Z6pB6nNLMVRGdwwO
/WD/dJVb4hVN0757/22X8fsJ8pdOESITG85cKKPG7f+iuBdql5a4AGB4dcH4vV9g
KnAgGVLHy4gN6s9rMC7W+Fgs1kq7Mr5lHRggwKIM+Yd7XaocLMACc5A2A04tP+Ee
l90UaWpTGN9w3aVjWIH4WdCSnTRof3vY6kAd0QtdJE+UPJSC4d5P0VgKpRu0eRS/
A5waVw1MivRrN7jic1GVjYOPW2qK9osSL2PUIdQy3LuL+T6ZN/dzGxUz6W3q/brj
1CpzJCQ1QJ6btQ2svxuHJAS0Ceufh+NhvxqX6xmEhd36QpECb13f5FwA9EmVXZJh
HwT6Ax201myP+em2zbsFF5ptfRxiMs1cRGDI0w6Rf15xKUKdygYda7i5KhRqb+Oa
vXcRM26HmwvsRLuev9r0Boc7EhOlpT+0+aoJ4Nw++6PEkFtIdlf/L4nbDkD44C7J
TCMzVLB45nM6gffwPmFTShg3AJXUUqPJvF/zRaqJ6D11uG8NqyY8tSY6sVer4j53
ET1yBv0Vz2Kt1ZonQ13J+8nCIlr05mNNQ3Pf2BICk5MaXwgOg7aLY7KCwfO6TX0b
sIa30zLFnOGFQjX+Rn9kxI9twhUxYTVt14+qmEnueVeIg6RwbIgpWoG9kWG16dBP
tfi83TNgHmfsnV+69JSmYnk9nSpvjCQ5IkllCv5RY6719A0Sl20VY1xo4WyamDuH
pxT/v+MBIRPQopjOlKGCZbcTQ/RsZ9GH9NRMpICLdlJnmhXRl9kzSTZJnaVqNFdY
TOce+AwECs7rWU+hx9KDh/ndk3+FVQY9GqRgVwG/jy/vs81mXcTjmJpHPM35sogs
R8Cnvug8qBkUxcRKwh+wELkmT0NzJa6OmG9qyzyG5ZEeXYMtTeNBnFeEVT7JZgmp
J41v9CQZAwDLrxrSo+SZ3XqngEbtruH9HHulIDf9p0Y/x8+gd9JcTn5GxpZs+BZN
4Bu66B5gwr+DyEtfTaGhob6szkQKmZUmYhylrC6HBjWiS0Q+iRdZG1Ueixyf/Eqc
C+0hYs9bpbonUWpW9iQFg0bv5D6cYo7XVEwVM+YQvoMMC5d1vc5eilyX/Tqf6cwi
2ti2hoFm+dSTspLxk5GAUMlLG0v41UOA0TuGGlxcwNg=
`protect END_PROTECTED
