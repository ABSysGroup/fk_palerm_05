`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/5CiWNUjUesz5ZorG5NWfSLHenr21DO2+QxF5KJQu/Y/ACkoAjzUDW9zl89EBXrd
fs9u8LWa1K4SRPnQuXcfCJQyfdynGW1reXKepSclhHUYqmO/83wTvCiwfMaieUvW
RzELOUTDKyK+KmXc/arRbFNt3l/GeL9vyCgCIppF+gHXyXkXC3OEx0VReTRn5fI8
Ucc8q+thtoKBLm0wR0rUITzbmmn8M2uABMo9DtqQ6onPeUqEubOU4n2j65db6GPr
IVgYavIgTYaMuJe3913OUmitiwBwTDOTnvKI2YYmO9sinX8lGdbFUlwOA7PG79Im
bRhwd0LHrk3+tIHf/4lVtQ==
`protect END_PROTECTED
