`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dShYKXcrNQlHyJTxIwZ5UJidfXRjWCK2khqoHN0FyVPLQAp/wkKJ5YrsWQZTTmMj
QEMBOZDkXTnnrWydU3pxczG3LOgr9mUMgs4LxbhlkYy26j8ln/8/d5XhpCE2GoMP
16+U1AVmmy3ZqIL6qYuwktVdEE/y4yDCHw869Hz/NGjBF3+w9AgIugFIelmn+sXw
sp/Qnggty1+VTxbdvjKkb0B9Wx3XG6VnBOA4uFZiOhXnkhnOPAuNdLPkackN7pcz
BdZgrTigWnFep1SG/IaJGdntuKfWVzTIm3fMVjrBBzs5Zv7NCcVPiLV1+ovAbZ6T
+ybw1stgq/g05tREEG4EypSP0kkdJfrlaYGGrzjNgG6dNYOCu0KIXYhKM9HT/N/v
tLAH0OwapYxbvutdPbSOBffvyw52YeMuZPAKKPz2QtxKSkWy/ma7AfyYxV6hYVDZ
loH44ExPuVZlfUTePi41KRjMyvinjG7pDGEMZps3/SF/lhTiqzeE1ZTx70/xsZhw
G2tX3xFpyaHHte82A1RD+mh1n8gTVP3IvZUr987cDEQ6v+bd4Acd4wN412YoiufS
`protect END_PROTECTED
