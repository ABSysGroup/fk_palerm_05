`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nctNoiECUz3g6nBrjFqXWgy+SdMjuRxdkyNm53Nhqj6sXHSBToRtm8E/vKpkE4bF
ndEdv20gZGztTQwipyRhlkLxE4cmtaXG45xaNGgaG5NWyvI0zr7yip1k2cvMTkS2
IEFxOosprvTFfNMJJgTyK7GdKXLHtNMlnYF3KzgEGT0p0XyYDO6gOZdNLJwxOjbL
7KMcwIBj9KLLKEbZHxiTRBpY3Ttssl+ZLaAFi6u39YT835ccu9S3rG8f7rO6bRef
VZM1XRYxj+xZVuXMkmVWznk6kFVsFKKu5EXurhdOVDUCXMNwF0/Vf71q6JH73YGn
llh3Cz2ibhYozATkMc+ntF4tuoQkUYToQBqumPm70q5qgfXoZBDSzwz7Kb2a1LTg
mR+SueRzv9Y+2nDM1/oyROHsemhqp6WC7iOIOizRHd16VFxztjCdR5H1BmmQyEo7
kFuH0NhP5Fkhng86bVJ9Z+j+93NRUK0FGUgkKCXNAYVq4F8afqBKiRgrdlgAX2T5
hs/P+udZoRdyV4hT8ab4fAcdhnCIekfwvTzesp5g0jyX0nAxAe15eRJFrmSrWvA5
EuwA4tzSKKnrbSj1OYAZBsjy2Xu5osvjEfpF8vtU/cKl6Zik0qiSZ8zIgJ8fIz54
O0pgqFeAnLkdAd4Zzjw4u24f/Fhgy355EMfZyJhppXxBPsBtnxOdJvjvZ1xcwWyL
xwGnPnkPcE8eB2nKjA9yQr1pOp2QA9qEcm3VB6a4bPN+6dIRsGuIwgn9C/hO1xk7
6hBNABmY4p33Nniexn8mIL7cE7HsgpTWBjXNW6SSPoYtXzHOyJYToHzoPK5P2zNd
I9HnjamwPmuflRKAHO+To2jwMVUr704vpvSWS+nZ5/g1WKY76WFsp9p/ztZxgg/I
kuWrRtMF3vDVFVygwTIWnJ/mhoJaOXgJi8ZcDBuQWWoV9mbuyvv9fbY5mR2IHdDz
refwxrxzYSHwK5Hze73JdqPZe2E2LZTmsDb9fGHcFysrOVTMvRIxze5BQJK1NEjX
uv24uAsvBG9lgGbPjojizu4C9z8/HsYAdyXRLmoE2e7FVHwJB0fTfncZqsDFsxA6
HfT0xSQU0VCPo3Xl4eejN/pheUhYB/7u4gHgwCAjlF+Mduq1hvXSgY2aaCqXqiV+
tvAlX6dEvqMiQyAgVZfzSVqO1crIA7WfY9WudjybAISG0rmN+aNB/JJ0T2UGnKJZ
qICK/W70OBgkBqnbp3JIXfIiTdHwVkv68vYTrPC0jC4Di59gDER9YFUxRES1Z9D+
vQXrCW7weK7c7WXB49JQ+zXqLFZO/WqphwVSLDO9ZhGtN11z89Iz9ZWbI8gqlrPO
hpnR2s7XVo5zn+uTSCu+lWdTwhYi72UePozhBxxuiZA21qsAGFxEQnNWfa8QldT4
c8UlQbYFCtSeSInm3FdigINnJLfcR8HO1LdUh0qUeV1IqjW/7LY0JW50kBe1cekd
1w4iPac0yD70v5IzmROtiqfAyPdmDq48ARTe9b8haMLkK9uKFkH0nXyRJXTlIGNB
Pr1os5d2Ji6d/esb7k22FVoCvCBqEohsW6/qwIcqXvRM1erC9ym21yN6bxuNf91s
J4fGc7abX0Yxqmz0ZzOA+sjxPKNoCkDoiv12QD/mlSUdkRLgbYD78IoBC97Zl7Sz
oXDnMF58rs65fk1IDayLu2uP8YrS88usZ1098x0aQlOSOxUJ9sm33S6q3g1O+jhY
GWY0CC7EsWbt3he6PtUFYDKTRUXOKnZ6/YT1poyoeU6ILAOHuCzcvS7uSYHaHtqb
bkKFxU+sejBDk8EYoJSQeZ7/a6pAcM9tBIA/48mYDnhcIDFRl7Wz9Xvuf3bzkvLO
uZoEdkWA0VCmaNQbm4ROtCjDfME4O1HqZaB/ufb+8FVxykmYfFme5nPjstaKb/NB
4SZUHGQBqcZJaOXa0kQoLFtVx5z2itqgONZkXvG2+a9R3boqD235BfSy8z//dnax
vu/OMBBhaga+vnSQx9FTYO8BDYWJnc1oOfhyEn0PNYgP7ubnnFINiWQA/96QBdod
1ODRsFGb0CKERGT/Ml9FMy0q7AQNx4jjdVR+T8fAzmz62leMbc6fop9uQ+uFthba
Z1CaT1REuw6g6SLhJOLgkf/z3IoQ58IQN5+Lk36VPg14iXhU6ZU2tshcn1BFllUf
wlCgBTIFxgzpDjqhRPl7kjSxuIwf1LXtYPjM+mceQpN+1R+P3lHSUcCpVVR1pEeT
TsOa6Pvj1tty4z3zqhejMldg6VDmYONY+MO1VPLTtWWL4NkAzlxIpKV9mCoMOV2M
jQ0xZqpAV4XulSd6BNQi5J/sSaqO6dbS6GWA04VHTVIvM9bGpAd/RzYDIDdfbnT7
NGoq1mlq6SIFQyGITD3QOgbr1kZoIbVqjDRMjZU4j1AFP3pEvyWtcrJOAKkERflW
kgBGhylDOQI1yUlYR7/R5k3DNtRM/NVfiA86QEP2coY=
`protect END_PROTECTED
