`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zfnx02fFoez6S+famHhwKeqahNlMH3sEE9Zx9/4q+m5eVZI5kwZQjy/5IGH5p8C7
jQwORhLetUpRm4PqAWUQVyHwkaK4uAe4Bq0GgG7XStvHLXZUTY9/IdGWyBiDNSNP
f5P3nVwo7zWC5gzLv7eY5SMsQQWgdD6KArUrRNF+HUIOuEkxlae7duNmwyzJmNSM
WA87ji3AiRTaYpIkcsDhayOJzUy8T53L71PX9gjzxdPkPE3UJNsKWjfXvXsii07J
fBtbhruEjv3DeBiF3+EskpFG/4BOSQLwkit60s2e1qbCytNcU2NUeCd3EwiX4Okh
coVdyOsz1UyrWDvUFa+kXl8tugvLrl0kEONkyZXgSJIHYr+bDZcuvzMcVCmC4yv1
pU0XgcwrcIpXa0o2ZimlVGkuMlw4azvOjdFUkW/2hVCgqlUn5CpFaHqNMHVqpBeX
b3ytAVMor4h6/YUmME3PSIjPRC+KvDo450wWZL8mF3bT+cRIhbSV1/TOrv6jGPio
FBgT8XtN7X9Z7E8kwagjXQLp3HrZo4nQ668giHqEVroKheBpJiTY+bnNN3Xpg2aR
zBqAzOVgfDNNx8BBfggF7YxVpmqHGmdhjOQbGGfTjBIdIWeAwYhFF6PO55AnV7d+
kDIAV6GjOKpGmixvG1BICw==
`protect END_PROTECTED
