`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oR3GCD4tNCa3bbNj8EwU9UwER23paF81OCGPhg0vj2YLRmnyA/3HLvWKE+yYul+J
fhYhNyjmizVP0etTH+RgOqFV3Wu2tVYIRE2EtyX/1S+gOn3dH+r5994Ib+TrG6tP
mSNEtcdOCIKc3/0SOwFdN1LEgGxN7bH+01E7CPhhTwKJ4ZDynXRX1Gx7uowrG8U1
F+B+olNN67y0Ha1Vq6cVUj1VZ+e/DbuLtK2ki3UbbjQ6ckxXnXs8yCvdakWh+ojL
83wpheDTjhRH/jHAFXBIN/VZ95HC8sfxnw03VnowlfNVJsSjd9vBuVZiLcHK67LJ
a7d5soBtwoNkrUOxVjomwFWwY7OWzRR+cERkd7Ej2IJnnZMqTJ6P/kqm2nDbO55X
HrFxYoTznj2s/N8iZd+q4ufN94rnvBoSTqpSKDJnlgjKC4uWuRFekMoUOCQnPS5p
XteZ+ugdw1SBDM/Hb81SgdrIjQNkEqz8N2RRwUKKoQg=
`protect END_PROTECTED
