`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O10WGokIoK8MioADQ5FpJ1HFuNNrDeEhX7jdqFomPm6uZ0ckvrBLLMGNsarXLdOm
Zhpb8QezBdoUqOMz40ne5YvSYqXGSssSZOLH3XkgbWDu3QD2m36j2XCbE+zmPmyv
UsrJsBmobyotch7VDxk2uSjkBFRIcTkN1wZcu1J4jz1tG8SYZ/Wx/aVLx7DhK1Lj
49nZFJ8zahXP+llaB1JADRbvrSYggFeI464brADkoxJ9GWmMANyHMGhyWhOXtRoY
aRdoC4JUljy4TJLSKpbDjQ==
`protect END_PROTECTED
