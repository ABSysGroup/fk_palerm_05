`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZcHWGR8NfR5budxfYon/dFTPb7XepJFoF5KtP2aOWaki7f16+ht6bxn/ue8PcdYe
IdeAkppoM8n5jJG46JtGYzqP72XXlGb9cZEeLjUGcl3a/wsXqIujSHHqs6AThhb1
JSFUhZcLJYPW6ktoMY6rw/CcIFXukxPOKzSNudk4DZWvZQkusTBYChhJLObaqwd8
3F8hrhcNSjBy8zm6BNXE2n4IOxQl50h3swPmWQ9QWqBmyRQyqBjIiN+2e43zqJLl
NvD2TfUQvV0Rji7Wfg5sTP0sLGdfLyFNrADhPnTP3Zq3j0egl0JWdokVqDohLVGS
NYGQvTzhlHPWlFd5e3DVsR268JcH6oppLRZgt1eGYLSpaiLmoyueUewm27N0/66i
yMVpxk1WjkoAwBULoIkkp7AEOTlcgUf7NsvM350yl1EXcDY0gL1WAomsQEIcFy0U
3VTVuSq0IfImqA40japL6/zt2iwcfaOjyN5TQbe85UbsbRzUOj7sut2f6QJANrRZ
ptAEXrefsp9KIEeuBR947Vz9gviabuLhTaWrCvDjmIhVhDa4+uf71DbmNeDk6yHo
`protect END_PROTECTED
