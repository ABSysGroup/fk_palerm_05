`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pTMLzFJ4cLbY7dd1XcalAKspehS9buTYbNAR8gwbEdbS1djoKUSKMsSmx9XDEfzz
QaAOAKNc4nOjCsEv4lB7Ug1In8HtCuh26x9UxOlC2uTrnuv0zjUCP/u444jkJ1QK
aePMMz3wO7LA/zParrBukemDg561OFMyPUcHYYLByeA8vdIigl0aM79yT1VE9aoP
SufS1JWnMO3yhUQeW4u/VgHTVIi73QTbSQgWmAEsSkpncSYzFsbK6ahcs9U2hA1K
T8xBNsmekknjJTvnajDNdMH73v8BPUV0iNq30qi4CS5Nct6cyprNfUFtcFNyrBjU
DX+iYr9Kni56QIM3qPMdVp2QbGDXXiNtIDiTC/b5qyHCLF/VC1srBgr1HtnPVDRD
ux6PzjEYSuBqQhRKoI3wdUCzJU1GZonmGe7CDdUR0QG7xGRdAEnL1PqEvmnrqsen
wTMGbSclqRc+YkPPYso1UFThGMuXu5kj8SlRfBkWo8c7B2Uj4Eq6HMDF/qjj7Rxj
YCR5m/yqtDwYOnbL72YQhrNQRqwMIOlRfB25Qf3W8Prk8UJUKr4FlneIcQ1Vfba1
w47CkC6nj0imH6sAKOMoRX8YZ7raPO+OG2VEH1Ze8ASCsKIwdEi473FTKNdu8Rvq
oj7qyXcRHIetZy26XsuNmoCKjNqlXuIxk16/o/X6g2WP9Ioiq3HAf7qUUDOSXwTa
WbLXJcKSrtVyMJ/w5TCLITEt2IRr0yKlcABmg5U823lSJm1KV6JEGKL0dTy5Q6sk
2LkOKTGs/tG54jZx9dY1sYeKaVob67yNQ0uRh4Cu3Eivi+NfBms6RBBnH4RwLAkS
+Vx1hvfOhk6+gt2agkVxrNqLtVFTrwy4IRcUHbCDJlL+czNbFFzGTP4U1n5O7y0e
K9mgnEI2zBXrHPRSPeIEjM8TjF6ShJGModq7kbXZZuJoh+FXLYgWKR4ilZ6+/Ok4
TLplZeUmKjnHw24+ZwCs/89J5ZsPfguTt0lda+ostQLC8NA5+w2Pslq2x6uz+Lm+
3jTEDejJW7zm3KCSAQr60jza9ZwANxFOXC1UFGQ66K4o1tbLq3iMAbNsdxuAoyQP
e+ni8BdkFzjI4OHZgdxsxr32OMQ94KSOxYFfNOQTOpfcnGNdijIPFPzxGH6NKtC2
dsC4TyJaLLvR4HkzFaYJ5wUK87Fx6CJKsItAvSZHgt8yHOBqP+m8P2muUJUrb5Sg
CXFrIXIgWZmHoPFYfjRaRYNZfj6pHl6+iabso/+WJN10lqtqrrUOgfjBjguN3AIk
0vEA0i210kFi28AEeTm7Nq4tU6yIXjugAeCmYJ8PmgQJ4QmVIpo/YpHoOMHMyzrA
6Fiba9GLhx+CKg68aDr19/UUuHCGeoi/Euc1FgByQ3UKlTmaLuAYEWR8iM7c5ldy
RenFCLMIt8sHm+lJ7zU9XDbdNZlELUOVn7nsG9bmiG+LOV6D19lEDdt5UzkIdD5+
nhL4U+zae74tH/7zqEl/fK1mT4DX1/ZARf1a8S4UZGc6CQ9/5kp+sJ8DZTzJIHNB
Xf0AaARqJOzU0VbdK3wMczFliNDw9x82s2YODGixjmn36pajP17MqGBkQrMav9Ye
dpcJw3knBFuxncB6sVVigU6BUCG+EbihzWE/G7CCI64mrJLln5uqD+WwLQw7e4Ib
YgzpN24upe+AVMWl5CZ8kZ8FcIzL0rQG2k/CpmxcZFFZ+Tq0cy5LZ6no+8s8K1RZ
ySXlhNuTq/47j8prWb0JR6haJVtkXEYa8fsvQ/Owg6G1tM9fjXuy07gjFzGj5Ajw
Z4//nKLK+VVCsWpUyUWLyB2+hjjpxPJmMpa5AQfyMo1BcLLFV2iHa2Sn+CrHRPub
7lVm9nUhgGo4cPGkIppwAA5kGoMzoJmKCLmIU2PXAo5E4y5hiw0f+rbeMOPZdqPM
muyfivAyexXF4ddfzfH3ojDGobQukmDysd2qXuwtDrYMOj4/icGOHYY/ZqlnBZ58
6+8H9I22oGOACw0mkvankf7ePEWQs3g76j9qjcmjekq6Pk9+wqu2trOQTTg16ZxN
4nAQ219z6oh2SkPOKaFPNW3t7ziUtIbUU+VWMZ8GC4e/dgKzBvOQZnatelB1I3Qo
DfJnxvNU6wJ2crnG/EwwaAfK/jMXzppUFP797Oidg4VK9JSol+AdpfxYn0rSNotv
TSHHW8RPlJKZ1/Ih06LO9X9SoaPhfYNTY6xmhJ6EWoK3OJBesQ+lp8Q1z0Id0aYq
QPpepLsu6DP8NZmuA7EeKjptzEf1+PQfTlPj0G3v+ifenNyqg2jYXH/smH3A3wyF
aAPbUxTomslB3w1WjZutJxaw6GcduOY7HjUDJKVooOz0SJUxTOefqPPMTPkXXp1E
IfliUyrgF/ojiBk8pigOfBeycBJqCLMSrNsWhL72/oR+wuAaZrqqj6PK0XnVL4HH
Ys8OnUOzqdWXO4INOVMc+je5l6pxkIzPSqOQ4PlnrjhR9WrbPijr2k8/ODeL8hV9
IE4khIyj7UdgPBasqMt5Xbk/fxRHl7h/6JGxWiP9iPxIL4940n61po5fwYceGjzK
uTj4K/15lt2B4csLKAY/Qly5yXcAiNJiAvENU9zEqUEk8Ae5ilHlGye98JINu3tP
kyzkdty2CXcBXX1NptXUwC49vCIxq+k6gFP6/taf7pxobYlhXiogpgSkYaBiDzmD
h43bdzrCHhTB6ecNW0z0q2egOogpbzxQjB2/KEotbTz1fyNXeHscgAwnYCwP31xB
tlQsJhis8/5k+4JWQiVozyh1GmIuG5WKw7FD4Q906JAxU2JkF05Dwrezz8rF1cMx
LW1zEsjewJsJVdU/afO66LW/wEymPPfjbuQU+4B1ie5TYbplLFFkgYdaJuiHyYjZ
Gi4w8sMzkkEmnu9BT2VlBEed1H1U3tBaH1TyMfU+rArdCfz5g2gaN+9qKLbNorKy
515sWCWHnsJUrfR07Z2rdtvcDl6wAEt+LxKEMMDj4pvQ6/hZxEBlpUQeF9Kl8tL8
VrPAtXmPlFqzu7LuzcU++ev9Ctw/SEoJ5hK1wafFSSv4IJLFKfqV3OAbyPNIRypW
RpXczn61NesLKePp6ztfkHCms7LQoSyXh2t1ixTbcm6tXO7lXmDfPb9qfVkikpG1
9kLqYXYdnsnpBu+sKdbGDdhy7XPzepauSJquQFfSxhXLOD7/mQG5zTubRTorS9FH
vGYKuCgu9PQusAMa2KQQR3r/Fq+SrYVi0RgijLqBQIl/sf22U/v0kMwzpPA/gVkR
Eer/Hbkd1ipI8FW/Y26r/KZYVMkHJyxN/JHTuutLuW6rZX+guJuYjDnNsHo6ikXW
lYkRwX37QuHnNPc4iMaMlqbde7FYE2GZTkAPIDYsUN6jtqjhEvYMEik3MsnxACTn
+PV1fRiKkJkz10erAo7+yl6h+iXW/RLB/Ks8yTk1us2kpuYAhGJ4nqcznPQdDC5Y
DwgjLkOykwCaYZ/N0YvaNJjKCGX8Ru/MDfzmihYUe93PEDsfrrsG2siwNSfiyKmd
Wz9+5DJxL5XRpRhxcDEX9Zf94aIm5BgWHzizkLk7ONkYnZFqVa0OQ3EoEFyuCK1h
hghdCwzyL3Qvbrw/yPWBRd+yAIMraS4e5uY6LuHjKed4rlUWvsRO66ZQqa8cqjFf
c4HvhyaYLsbli2Y3N4jsfKew0m5IHqw0/0TrRgJwJ46ulrFlo8Ssba7PgMNOCu95
cBv0MA9lH/iUX9oAZsD5/HKGEtXVVxQM/jtGlAfx0flW709dJXr8UTx+mIWeDiqo
UrziSPzyVpxSsiE+hznKET5TBZkKl6ujgTwc04CG0iP2LUiADS9m6P9flXYybCgC
HuxpTzxRFp9sp3HxgJHx2vqhcR2Ho24xuscVd+iJrEgJrS8WBF4kezQBkRqt+XgQ
YMtd5Eli09o84x5h5JI/X9K0o7HB8wA/oGJ3SLeIMQmLVt9MOrMCEzdj0wPJ99KB
LSywUkyMJQ06yff3J2rFLNN9DCrOW8aBFRRzOLganpgNnxFPe4KCBess0q65Ty+V
AJpR0d1fl4vjQPEh2wG4Z9Q7RxQkwsb7vV7W+PxYJshQDEGb8uj4ziARkRumTe1e
S0V6B+sqzlnxZHLY1hj4RzndR3mB0SCWjlXpeAtq9bmUtMZU+vCxWncZ42YNWaeN
`protect END_PROTECTED
