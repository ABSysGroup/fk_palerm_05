`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rLlrMcYl0mTxSQPv2Ux4QXJy7+epm9EsQf/8+0A8bgx4sYtPfIW38Q76IJ0cHYTv
7WlL1ty2vJbW1g0JP2Ku4Lr4roRno+d1obH/RBjzz5UmP7dwgJZbwJ9huMBIxsNu
Qr66SNYsmxWd7bvfbgOzDbptgptl9dc8A+Dp5hD7W2tk3tl3AUCclQtkmNv17wrD
B/RQqJle0EbPoazjdPYPn37xMz3XJQlo62Nrb1Q3KCCw4r+npgAJwWRhUGE+6g4Z
rTjX5sd9wrsVyVN0PCphohdGZlsp86KO0ZPOxmHCayaQINfwj+vt4WV5X9DUtOl0
TPVDnkzrLayGNQSE9DwqxAkTxCaqzKgCHSXbziZ4f+m9CNXsy6ybdgHILKrhxuGB
+h+dpiEDKNepfO8qJ26tww==
`protect END_PROTECTED
