`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mzfKz/rNTMoVsQqy+WJRpl8l8vbP1vtzUZdJAMSSDDZ2cKKu/ggvQFUzzu815p/E
ez+pYyQdmyPF1yo+fxwSCOBCZZFRwk2KcJbQZ7zfJjgf5Lx1Uuftq9SmhCpKCEon
Tb/BNrDzPGdF2Hv2XdphUDQXkyd5x09MSlY1Eh+BsBZ358Lr7OIkOBv6193TbtNA
rgXlSRS6aaQV5eV8zcG3g88b9oeq4FUlnylXKq6Ibas0QyOE2Nk0m9Sp06MwJmHK
9Gv7b4mQn1no8gNU2KvDQcd76puiFibex7N2jKay6MZmbd7RsZOBvotyeezRzTo+
M/S3lxTrGwe1ZP/8AEgCoq1hEsy33IIjN7Y1cmlfromW960B+emy1illBDiBnDu8
qTQSUG0ZAiNF+BOZ8euYKp9qrIszPtn5QsvL+MZNqHFza0wkglLquNWkCqFTcus4
H73eVGvCuqurlt4I5TTRL6fSahhZ7RY6GOvoNrto6OlnO8188cHiqF3oI8xBHU9e
3KM3setrANFAOUq/orWGT2YG1+41uFlp/FtF2f0rVk5oSYSGS6oTJdBmF41NKh3e
rrWko1sc+MFhocFinDkm0h88o9AuHzp7kfy/GwdHZ7M+jUzgWLrr8vSg99DZwGuJ
E8zuVrNDiQtqfVQqP0LAoji9qcPi8xdKSN615LLP+BzvibRHl2dhts5zcqabmaPT
aQXGZl8oT67+YWDntSIC7kAgZaF2HedGeIotSaVmcl2kl2Th9igIoWsJXBfrGl3h
mjyc1tsCkrfB43JN7AXygIHQQ7mBfWlN2gbFW8kQRE4pYq5EFIA7aaF3g+RX1THq
BVEvkizT5P8dBYW/BonXuRyjttqyXNaf0vEeH1PIi+9o53XqgHPlRx/U5jiSVtqa
5AHK75OBMwRIZdoiX0epxbHZ68sufjW7y/52iSrLylfumrsOU4AR0Q7ISR/1S1Kg
yfl2hL39lhbR2PsDqVbiMAIUBF8M2tBM6W9lSguZmTAPgiqKrYAzfPnP+asymaqn
/MHwQRpmaHxU5+2FVO2C+Jfsp25XiQ0ER4UbOTIPMv37MPPVB3PhjR6h6CYckquw
CdfE+633SfNOLRsyuS1Od9AHjhsz4wThAbDUrOHPYHoprOjjqnjWDsXvlcA0TdNi
0ersSkR2THCj0yy935ivLUNpU5sRAOSyg8oAms3H7aov2RILydHrvh4otyib3rbN
wLuqTUdYfH5pZ7LntDu3TA==
`protect END_PROTECTED
