`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T29223hXdk8blCb468z1j3PsO8/L8FnHDwXxDJtg/qhPO0Pvs51434y5MJxQDbIm
BATwBvwPENmzJL34yO1VoYfBsByh83S1TzbhdKR1cIWcm/1M79t/XIh16yYEj0hg
VqGMu0OAfLdEcg7Vr/xYGPP+bUZTQWI0vtWik6KPZxg8m/a9Y0EG42LOnhrD3guv
On/5NBxZZB32+7cYtlmqKwUC/YUrwSMmYYzdRSjmQWPOx0TEN8Xw4oqvP3KniKqy
9vFMrJsjNLd2KQRcsNI9a3dmjnYxTrMOBY+ZQk2OIRUCu8xegJI8L9/YVxqyCY6G
Jmjyt/LAFshs2CbsT8oTW1J7G7O5JCugYwVVlUeKbsEmivdpIWHIbm05LUyin3Df
/S3gp4Ypg27M1AiN8HnmPiYg6WeRxUl/JpcvIC1eYJSqLtOgTpi/I2rYPON6wT3+
ZRFFQBWYXoINylWTIlzyug==
`protect END_PROTECTED
