`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eqeoU0kAgKPtxpXQNdStHYmrltBWa+TRF/S/SyDZIIBmPXcnFljSpJjI7tK9Q8Aq
r9FCXTHb1gNghchI2Q6ipQ/bTmlzZOq3k6lvNQjTsJQd50SImyjx+0/SDoIIIlV6
bw49f2bmi4LUqxQjGY+GUT0girQx1oTir9rBU1coJk9rcOuq9SIZtPyNi1JHHPBc
lAVoEKU+UDREDv5Q9ggdxyEcfUchoQFFEBYm05hTc2Z+mMkhzeUkL6tL6xfF0BSU
AUOtyWq7IR9Ew+mlYsNe+03QSpptmM7ngSleDFGcxLCysTLMs1JPe8kJoxa5U84w
tJZkK2Ki0qX1Fy5wl+7YwMaDLl/N4wTuPcVc4KG3WxItd5KoXphdOv5W8aT0ZMP+
+DgJuWI1eckbz+zoRITpNDRZnG5R0QmEIRTZw9Wqy9E/FHyH/28dg8H/6pJmXNSO
plN8OutTO8mvR84TGrpdlFJi3/pL+Xwh9EQHgqgB9ivq+d9GSrZZOcQkTWdEMZAF
M+uuChddvyaT8Q/dMUXJlEijVkGpx0QxfbcHvwbT+Mfeq2Z6ptmlv+0khH5clPZi
4SoDBoLDnL+q2q7Cq0tjqREvz5uFjZArbfTK3hXbEHmar9CPdFlqEUqiARqCRNl/
E4EET1WIcroU4oGoAUaJ60zuAlsvsGwv/WbBigiFWzoaM4BAhaq3YhgVLE6Zla3o
GbryuhWCMbHwGRJ++XLfQUM2oDOsxeXFu2qplSnqlV+V8XFTLugl6f0O1I6zpOtG
pvFE4k+kUkvAxtVeWQglRToFK72Xh2RhZ18ZMXGq7GykrjHyVsXQmnOh/7Suwmmw
8J3ukbCHL4s5rweMRstTBirEu1YhGZAu1tB49Ix02vepE0UIPn9CRcCZdb6dPe2x
YG5cdh9rJf2IAcc49YjirQ7Phq6SD2y1tLVf70kB7wrKbU/YDT0uf0xjKHb/OeK0
`protect END_PROTECTED
