`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vR9EK35txUaNkkE1S5Nu8TQ2qFKvGcfchj1C8ntpyiqDNgxa1ze2e+GyW8gxhMoK
vEaoQEeT6TdW4hDSR3TqW1wkqddnhe8qz11qHkJkrl1EjHygs6zp9oRkts0iTmxj
uxE6j/X4NBMJmgT8vu/XqIDIb252dCaVAgZ66Zt4Q1biV77nzFu1kuNam6TUeu04
MBifACSvwKKKEJdPAk+l2eBKTlbAb18NpBlZskvNZod5/Sgr8iPH0p42XHs3sA3k
O5kqWxh6Wf8unhlgzcpftUbXRh/yWcrARfjadjF0UV+V2oBIKNH+wPttgESenPrr
YzNsigBV3IxM8PiiT9OpOYr2j+q+Nawo0d6ZtbDO4UGIJ6z8L9Wl4uDyN+IoAEp1
qDtxjxmeXhTmUwDcPb9DM/10x1AA37qmXz2LnycVPjsuJOYu/ld9jJbcIBM1ESGb
1GAK8ZSoUsOH3hk28h9eXpnfOhdXuIN7IkYppPO1ZT7XLOAODAZfRaiaocBoiwrb
Kc9MDp/CTyK0zKNp3GRisdYkQ6wbQnuiI7+bkBW4QOqS+8hzUITYFFTLpJOVUg1m
gq19udesaIcodUgkC1C8CLQFBLWyldsgovg8QB4eUT9qlVFvLGzuaLXssxuNoK5Q
09gj0xxqBWPMo7YAU+GsNEnLw0061/r78AGYu5WvwfdkuQy5AS6mVz0IRatn+xcS
Bc2nK2Ig0bEEzus0wIf+tYFUVT4hHS0+gj6Am4GewlbofE/+NvRH7eebgJD3VXUn
9ENSeG8tDaJ6b1YgJZMawvylddGXKOcgJjAC2c3ANs55N+FvtAmcSLtGwmX4e6jx
Uu93az7BwFGb4+H4iRWh3L/hs4u7V9tew0tH8TyKVEcFuP8Dp5oxvL+H5dh4PhTR
Aoz+vhfYgy53pn1U1aGAX/lCutS7Uytx3/pjZwnKBQLfH9UK2lMMhYv9zkQel3a5
tclxvHp6y3oVqVpaHyLgiB1esfmf9jdmVws9yKM2gNHIBVkSMVxwE+IaCZzAdDI0
8T2HJkMgCBymjFWMfud5vC+FkFqlc6IaXNQ5HRxPVZpCFWTNcXq8nXmP/GJMPjpR
z10PUP+/NWE6JuN74Bh+pZB06JmtzTgj+1r9racUar+wAIk98p29Nofe3Y7cnOe7
xYW34D7XW9XN20RUf8aO13cSCllL0LAPwO4/UxG7+T/eJgfOJYmR+mcPAeiZrrzY
5MwNyi9GCfxw7fZq9U96Xhc7YHanRl3DR/LoCKz8j3sK22SgHguID0WWFfPd9b0/
1rS1RqhZnDLBCZiqxEJ8INAt2foSi79QByB+rCnAfkGRSRxnXOhMXoMXNMTowa9B
MO8sKI/4VZ8hZ2Rcw98lPTvYf7eJWjSBZB+3rlBJcvcC1niRexh4k9LDgNhU+6+F
6/FDUW2Bp8Q5qUiZCsIhmxTxqN9a/6JeSQ7oBZ8T6sBoFkamPTFg8cTIdbq6PdKA
cGLo6cuBylXxBAzaIVuRus8OnXF3FXuZxSjlZAgmsfeWqREO30HsA/xBYmqynoqs
aFJ4nCZCU6bG8mdgS97MkPhuS2a8m80OwCLOCjaRnzNfj9dKPyh8L+s/JAVvg46x
rPaGKsnjvuQOljFpqTGU8Mg0Mv/FoAeFN7CNjybMrJGMoVM0ATWqe2zi68Qt7CSA
YzCP/aSeGKaGbfhUEtE3FqULuJ8phg92qcv3UlUUpfirzU1JUbh9Bdv0sQd1Tx0k
i1iXLGbNAvXlN1B+4a0WclxVuY4td3pz5QJwec/AEpXq2GsE6PUoqN8/rR+g4x+2
GzpvvprmPG+RMjepElmR3hajMKse7z30z4j9RpscX7Xp3U1xre0pe3Tuz88yLkDV
w+LTbCQxKoCvk7f8TA7zYZ2AhzR8thE68foWMbTIDXCGpoIv60onD+BfW4T76l+y
6BlTboOrzJ6CBXDfprXAXkVIKmJS+a3pW3ZETPEOgDTgWHioLyLGrI6H7GjD1tTY
56Y2ULWHslBucmPlVfL4u1j4bZ7z9SyHxuovfIuuhNNLSG8UV+ruWrObiFmaPAEs
ozrsYSDkxQBxu4W+HhEvdUXSoM1qWTUDkckHdqdZI2TlPF+Jsi9OJQ/w7qn0Q0Xw
l37fZDz/CjbS7kVLJM6+V1eXuIermCV55LlrQhIZOCLQ+kWQK3gNfKp2IKHEjBr2
aofTNSa4EuNwdlEXEBptBDTREVKCqG84p0+WdNXB2aC7znQBzQ7bjN+55HT8a0R/
rcwgUz/6Z1PZA17oRTiWNxEU6J9MArfI9RlPgG2tQ+F9QiRNjvlii8Bm5QOAs8+O
XCW1Uru4yy9VELWls8gLzKnaqxURi/i3+2G6bItBCSwNxRMdMiDnfmaWgHKfZcRk
gMd8rL1ouBXK2xyyp4zbbngY5UotTpRSvjthlXUu99DdjhzWf91Ot+rew8I9coV8
m9QMHBpHfHDETpVkvA1zEDkdhB8xo9I3r09pA0qkFAyA5+o05i/ci8Hul3sCvIRL
Ve2iObOlCm29rbWFN5BN1/ZKM0oKVLPjA26SRAW7ZHXP6PM/jt1Wo9AhEVfTx8D8
inI8XOYm7x1UJv0fm/9rARrtyaiHAuSnJ4ogEZEe1JI447LEQ8KE9SHptzRIO6p+
E3VA5+B9oi2Dz7osZHhdtC+aGhfIIghxYYzShGY/U8PeBbMGJ82iBQOBW55u1NYJ
scjJH8AFP/JHNt2KwQW817GR7m5Zpyo8RBabd54quM0CgI1lh/KD9MOgohDDys2v
nyZ1SqCxdD0HELAUa1+ps/hVgKZXAQ3rQZ/X/vn4/RXmO9k74w+LejQ5AVYcz3z2
ZldtHudq+xYGMcyS+05rPxUEaOJCk81qCj1+WVgby6lyImmTh0hxHSIonMTHoWFO
OmJNgmZBSo2pgWvKk58V6GNuZRoZOjKfS51t/3ihQFIbp2gGiKM6ctBtCHeMq70C
5RRqSytMXSUmS/DbYwHIsZqIBwEyFY4MVqXFaRyxE+/wBqeIuRAmYKvQ5e6hCEyQ
voi/uENsK/WErGfImu/ehAGkbt8wIPnWP8RS2xduXVz6hskAPvuAmcS8fAnncItJ
giU65L/QqpDqiYG2BR08wz467CBcWH1TfkgT5AtdL3LXH4lHLQgO+TUVy+FKvy36
si4X5UgTqLdbgJsI8Lcl7C60Q0E2AVNmCL+2hVPhhT9vl+fdqL/C2DhUrjV6VeNN
z3z6arxmZQT7Ck5rAobfXseTyvXEAZMaxcrGhlt65Bgk+dgJJybTE5sRERpa1quk
k53nsQ2H82eghf+69hjmZrkrM/NZKCPHUXufpOYKJECf3cIgnp/DH/xtkmztp4+W
QNHCLxFiCwittOlbAbmevRqFnB26deT4KQjHGmgDPkz9GDpREaqE+pLSo5l2oKpi
sA/z45vZpUCa7xhtcIpjxQ4a3z7AlcaJqHltrCJnXVWmjGWLAKbqV0pCUGK+DIfo
y9wGn3t9h2QKMaV5B43Ea2QZGP6bpOoDoB5kQTX8ClP7OjokQzgEbu4ehMbclIRW
MhoXaQ0+CjpwEhkIqX0HTx5TNtPHZ50ljjWRf2DBnwUuE0reZs4y5EPyeHXN5pOw
qrcaOp9sdWfsVLUFzNnacPrVn1heXHe8DFSn5Nvi+f5xZhNb4fhVtcBJHsLXDjI7
xAUJOSDjjD/SRSIefLFoGv/SBCI0GMrPeTGfsCNy0BXfrhvcTTMoWVGeLemly9s/
Ly8kcmrriOsJA1GC4NF9pW3yXQqB3XEdjfkiE+34a9yDWMAH0MyYLpeHMYB+yUFJ
4UlRlxH/jIu35/MwQYRWp5fRlCbsPK6axOBDe21BTLudkNtOG9vtGeQFjW6KFwSD
It8+aFPtRPg56l+1iDP1KqW7hjfIDIGJN2VhgJqTTBRWOAdEESXele2iM6Aaxwni
VtsR3LDOM4L/3M8m5VREG5wjhvLTgFb+jkmT4lL2I5pP0mNZnGwXDuHag8zmlz3X
25+ON6wWshdrH26p9sttWq45cIjThbM6ouXqwo/xSfaWgNMXqfJ3fqsjGBnQYoPa
REK+eGc8D567SEDP7NANHEoaDEnFb66OdXcY8z5+LI/kgwh4oZHU9VgCa5W1hOBM
4vPT8YDoqEIYzKqxjxRROWp8/HBs0EHQqxfl/CVytZG6pdGTVvc+EtcD/adB0hZP
5Rd4K8NZ0A9uB/SrztWpNVrBAezsjifnMBu8uNava2yjjVKQQbvaw7Y7TFcJoZAU
M90Gia65Y80JXGneizPtF1ugJzZyCk2qA1L+DgY9zz2dZuR0HY2f2ERFQFOTMkl3
9KoSbTtzwGl9MoAFCTuZnBl+rAYFQE1Lr02ZZYrrS7LahHKQ4AWTFKoKzrjCcRNt
CrYxkpNE68IHT4VTDjhEwpKURF04xwpMGbi8QBwbMZMioDtnTpDDfxRvtsIK7dof
uMaUERR9cqT6aLfCkclmzSuslXt1nVbAIqWC2ep7oWBWueA1g0WBSBXTCKA9Wqv5
TIIDmnG/WDBaWPRL+78o62eXAUcE39sSRdlIz82i2D58rkUKFA3HKj1jssOKQxR4
0hdIDgeYJgvZ1ZUHL3eQqhQcd2wB/jAG0vANYwlp4VZzk/dsm9mXAszfgJ2wJOBh
gU1UddXxiuPo4V/pdiUrULnv+MBFt3l4dNnmTLo/ouE7WGfBmfNnL3htq5s96fF9
QfKr2n8yd68XRbtZD47RbKFITVg5XNtgGr82VmIQXykkNmSlioj+1xKJ9F8Nv9uQ
P8QFDVq2DRzVhX5jY/3WujDdoLpI5HtCxpXPGXRr3V4DLKlH1/rAxH8oLYzNCzip
gfGZTVmmMKFdu7uQ/UWup5LcTt46UhtNs1rNsp63mVq23q8Eqi6fe8T2q6zgFcaK
UOxzFkZr44j05NtpazF9HGqe8Y4YRQ4yFC6AK10ZaaQkSfc7FjyISMaPjT5YqqDi
IvKgowrtDw/2Bin47fzG4IcpfI5BnWhdYR3heH2N47D/GzF822/HN0rmoFmGsI5b
HCUNoV11iOPM1hlDgTVgvvx3cIfD+8aZ6SaCEnl+riXIJUSlq3nzFCb8XNg0cxAc
dEBqXBOu+PyXNxCeTRFxPRHg02azm4l5UiaZwiV4LTY84tz7T0aYqncatrj1YViw
rwtS8CapLgFCbz1uPlUJk+cizudlxc9ohew+1WO2rlv2Zn2cuCgwMSrp/5oxP+Sb
RR9A2AWY9/U0JhH5k0iVk2Pa+ZUBrOf7dQsM3JLfI5h86dJHkXTCiewqWPznrOmm
eMe1scqXgGD4mGS7AWd37DfD7mYpI9Q7MM0bzmUyoQCBeQ/9NnLUHr4dOZTr3Gfq
L78M/vRYjttoLUwBIRHG6ML1o9FAOIKLd6t9lcU0aisRBcHd7vS1C+jfB3p23OOI
Z/Dw1rteyoSX709loqL6D2kRdc+F7gy0s339Q35cabzllrET0eKpn+xtMucI2tNM
hehWARQUgGVX6/95qjvZSn9wddOQw8L0mQ8D2d4xSR6b6y+yQyQyMh0XXMBvpBg1
/8zmRejGDFKxVq7gj86IE1Hr3FuunOuXc2Ter74G0mTFxtfNqXejD5GB1Q7/j+ZJ
BwYL3/7HT22Dcr7XbObQ96u3ReQ4MpfuIrAm0nYuvQ7b0xfH3idmq89Jarlj94Gj
0+OToDA+Sb6/rtZLTm5q1vJJQQ0UzU9ZErRi4DdiM89JZItONwdAU83zo5aBNMOj
JFFp3qR73jQGPSBorlPblC/nkwHaPyjSxZAXPfXcMFbBeHW5dtkHwWtcW7/tdSj4
P1MNKCEYpSFp7NWUA7PUn5EEXFJyHJxhVuG9gRzipJ4jF4+qgn8GNoVoB1h+Fcrr
PnFKHPoelrGi30kphnMB2CAKjb4Y9mlVDUxR6HC7p5YzNMpptKpU5gmUwTa2MVF+
h69wENfRVK8PQzMmTu2LU73/C8KaooQ67Qw+z/zdzIVygJk/Kb1h4DbRqLj28CSz
y4Per/DdGL0bYHnY68SDVToTP4sM7onnAAaQpCqeO5mKmrVukvmnQU2hioK7U4mp
y7amIjTQqAWGq6OBNeThWtnzQFJTAgMWV4iW7FPpPdrJRWUfOJgEKf2+mVJ+pZvC
+/XBqZja8YfUbG+tHg4gwpW3Lwa0RtnSQNa5xNOSI8qx9CJa/m9KZ19hfz9jPZ9h
jQrNyJR4gFcrvr3pw/Dt99xc3ZWJWmcL1KSGII70w1CxXMot1ewXu/+2uy1/Hzr7
dJgE0HUfVuPOztFPsB2OYv4htfrgas1ZvgQIc/cZFaKqTSyyLxQLa9cIUtmCddeH
gqauiALP+ZLjovMmmiEtGpCfw/+DhK0d0lnEdXpx/QsiGMBaE/51wiVHLt56bWI0
H69RZyZ383mZeUMpw027Hmw7AlswdQrdnzqR1CUWvscbjV0l6XqFRxh76lwJbQLp
yONug4MUSQ8t+IzqweHcTFrk0CJSReMIg8k9O3SFgg6i6sho2oLwNxCwAIEDn0Xq
aDfuQCb05z1tiCALIusasaeAXoSHAbn4LyTj2P+A/uDkKUjPQz2OmwV+y6qrFjbY
MW+3Di+8xx7CFHr4PEsu8MuWXxnyHEQz40lxGv+3FBeLEWO21NVBxYr+mfpg5ZcA
eUSwYQOe63i9iYC58UeR2Try3fxpKE2fbgnOMRYBrdyYrcGFGqVJB3tr2fD5Qt0Y
ic//WAV8xO+lRR8EsF/+hfRFawLXv+uHOT7f2Q4UFdy8meuV+YyTqE4G/bG5EHp9
ugulyg4IFcCReBzWmCfWMvFMEQEDqf9Y+Le3w+Yb4pE0MnujRk8+lzHJ1DveX+su
ulk6KT73B+9RwQQ3MnmKvt+1UVEyUFM6VvHv8yy9UTb8GoCgnAgI7FfWLVAvmPZ2
ft+Q0pwvU0HcyZ4ByOganWKpQHD5pmzT/axTqRCzVLdepkYDgZPgYM0pUmqhZKxt
DzM5WXBZpkCnBEN6dr2UqLy90JOUh5yFBNxD+NBpB3hSitE7/6cOSXgmlYZeb6zN
KSnAVMojmuojh3tBw5nQ8eBASVH7X1quLFw+JCAGx86zZXNjYYAaBMbYO0OckEVD
nhWm4CtIZ4rCgq22XYk0jxbrkXz5nW91yU9KJ0DIbbiKNmQCRsLm6D1mG2yMfrgV
1HaU/X3O159CCFzuF9rVi3J64LcHUWKrvEtJODflkT5l1eTaGZlc5mA1uVgUtrz/
RsuOpmrR2UBOo1b0LtEckPvua6s01SN8cWcq5XygjjGLrWU1BOv0aX5eDkCylVL4
AabP4Jq4ivbuOAqs34BLfzSBiAgxldBN6utsWlLqVH9kbBwLoqWtSLm/82Epdgb8
Fq+/7qZ3qOBd6+sSfenGI3ch3NV33eLQdYyomlGFnYw+f46n4K1Qm4GqOEo8WP1R
Abo7U9KO0wWy3w+2kwoRPc6XE3BcacyLFCAcOp5A6uALXW6EpgR+rqNGNfZ1mw7i
78UH6C2a0hrYRbRWV1ddVDT/cvCFS1DYYlHVKlhhV2s5Lp36l1YMjj+yHVtw+tgr
aSvE8mKQ1wrRqlTVTm8ryGf9qDsmUJ/iRadK7oyuV0xj3Sox1hGeIrJ9rb7G7blE
fcR6y1Du4wq0zYcFT2Dn9D3VyOCkW96J8miVZDT92z1gnpAZpNbD7fqSEeX35F6y
Z6sm1BVMeI8ydiXt2XiSf5/uQDJ2FMF9o39Ipk7NELopfHvfiTV4QTZW2z+kIagp
iZjmOIrLa2p8nmQubA8iCKK8fSLsIzSv1qmHLBalCL5JUQYNDbUxc/uqcnr0vm4Z
cPw64CbIBgOeaqj5jq/PHt3VZiL+aNMa4jIy1O9r84PxnOJP+0lfYxSxVQbJlJz0
98l+6jxNsyXBij1Ef/DW7FH4CKW2cMBAW5h7RvTsyX4wUxCkgd3oz1HlmiakWdW9
IPht10t4V2LNsv+2dQtxrLfwXLaU8AaOrz28ffElNl7d/0Isc3YjrQ6NN9ji6wtA
UDyTaUAC7Zn8fHthLRzj1CIx2bEuwcQUh1+6frFDOhnVzl9kC/erXVYgBeCUJi40
vK/hETYJjAIQyBq8IhMuAAapuTdfjho8biAoiO4Q4JYhWIaMJ7cAGsMkydca1u3L
Em9L7ogM8/wT697Y29bJN8MnrtJ9UGONT+lcyKpwTtr4XuSeg5znXQBV9raAJkGA
VoLUX8waqNbA4PjmiqB6n4QnwMDQtYmgcFGnAm4Cx0HwgkygtFaJix8tjUJcjIsl
XuFaaqef3pZndMM2337klje7kykTlWnxZAJPaskrFBSn3TtxReQb3i5jEODTT74+
fRMLM1g9PcXUKDgU8lrlYJuG/VDYaEpOOUdW1W0YbMdtiIFbPrfOTCEVOyP2/Gky
mI1T/fHBhlpYQi4mYN3xJcbx7xUm0pmXstkcwGRIEXtnttSl6KziRVaxR30DMZTl
lzGRZpUsGb/DRzAwIMGS5omkuF99nGKdq4ThJvHGdK6JuXgzTWk9pNgffGmS4Q7Z
3JVErV/ePZrb5cV+ED0fvbGkTT824z/r0mZFRhpJwqzJ0O6SRLoAgdfTi83kYlxF
q3p5hmDQhZhecITMH01b+iMhoqZT1D3Ba0cwuxdNcsb5VilvXQykdZHSuFhdEqck
iPCfjx7XGfwyXQT6w/mnApZn8cfWoIiISkTCPKa3Il9ZSm7oPgkgVMehE2wWoO1s
YAMQxj5WnRBfxYZrYA3A5eOmWvMpa0v4Rvmtq+kGRvCbZNol7jtvlucJ9hDF9qgF
WRvY4TU95n5zcovUGk88LTtdN3XM0oTO0OlE1lNxL0ByxPFhUbFTcNT59VgM6yOX
Qmg+wVQrH9X+gIBRjwo61LXlWSHOytFsNKdPBwIwzudPVWOx9I+Lvj8Io3V/Z97M
jy92AZWwSOa1qYsHAuttGaGUPkAc6/xPWiYmIImrSVey2aBj7I7+FuWSWkP4o1Nn
VFoG+tLIb4BhZpn6+99lp/yOrStMgoyVqPq70mJq9RT7+w9hdg+0iZeqngkKY6cR
y1yqQlsXM66xKEUxv75r+HS7K+73EGOSanMLJh/6uQMkemTHk3pBhHso9UzRNK5M
8KouNzziaM1SgArofgg5Gv2voi+KzVacbXyeysDWswZPKI7K5zEPWliJMrruOLaZ
JWuy383i+ik4cTn9Vj7n18VS2gsqfc8qvVZYFusaTUIcyoHh0jN8YbL/h+sVSnwT
C+jbDsXOAf4YF+/yyLG1JKNFOjMRF73tqeFYriUyc64dSk34gGnmmQPH+aXp19Kv
XordsAVu5qdXO+yhyKaZ5jfvMAsCBzLTfB6Rl6+DkJ7qQvN9Mzd8dN6PKk/jVADU
GT+Y+49xgfDn5dSqFyJHZ6nnhfeoYuqyTYP+TQZE7/JkQWcbt8r/cbzbzl9B4cCg
m1VvzClAexDwyPs6kDK+fzvQfpTyvi87ubVYo+0Q8XUwVWQdm4WUm9wzKM0kqceO
6rm9tJkLyrbbetRe7t67tAvOkwXm3L1gbMM+UEZr3QrGf7vB7spyPAa9SWacP3VK
vGy4WK0XPo/iSqLIM8HjuyuQiUs+GL1Q8NjKdcv+tiMPUOBBT28QHE8Yii7nxIyH
Z4zyUuoNMXj5Z1x86fMzZ/p5TQo88/LNpH848mceSSCePk1wQzN4kIioZi7qwU0E
ysieVK9sibXHqusoAX5glT70D6F2ep4dQly2/8Eh/HlB/RTCOHejdNs9EWW0ow5e
zkQjg3Bd0hhaYh3lSgtC4KECzgTo9EJDQDfSqkMTRtHeBhXxXBrdgnyxD65160pC
qD+5m7J//3QXqXZ7eNpPdxwjFAKY00xsCFQjDT+VFR/WVyi5k9NQ+6X8Em5o1Rko
hxeZpVc3CsPeHaYay8kWvKbGy/smbvBm0Qi++pwIsqg5K/PcQd9lChwn0hwoBKkz
fkrSahE40D6pb3GRH02jDK86GD9wpKyRTUg0ZRZEOwIIXUbZwDGCLVaai9fra39p
yGaHMKyvEPaNnWRtxTCCK5FPNB5sdiaMeUx7UR96F8ao42t7G4kUOVL4qRhSoVGw
s76/fIz8MySQ8BvV5G3t5Tv+8MIjvZ8MxVCBxFUygWTLF69JQw2CrnDXxXeuCNLO
vJTUYHsYSglZl1eN9Svv1CP+ZYG0kQ6CIJXs17MlU+qo8lxRd5/BI2xcE1IX0Vsi
oCcu/7CQ9qAUK5Qfy0wYvPvXMeOBBEQdxMsea4JpxU2Lu0e3gArJDbf2DqdoqEJ8
Xw46TrSHS4UO3rfYIyeL9YQRP19PMtMuEv0foYZkZR2m+hne6t5SWxuKlRVJqYhM
NGZWl7ijYJp4ju+U4ABCvBJ9H2vm2JuSlPnS2x+qx6VCxUrlMsGA+sCs82eBM3Wn
tijhaFm1a0CSdy7HZcx17cdwDV9zbZdcYHIxVlNbockD0biUlxM0lAROT3vAltDf
pQDVpP0Y9oWCmV9fuQiV6G3bzi9xu20JFOh1AGU6zCJhwXHTnNlr9zQKac/6vo8U
+fY3aXF2m5L/Le+2qXDO/c3ZdccwUz1xlNb6KaNhhIlz4grCJIe3Y22LTC4tkTHP
CG85CgocSJoKXH6n9S24l6tWmsWhrf8tSkNwEea7Bl8RCnmfFLRmG7rb7B4Qxa6L
0AAByW1JNJi6MWNEmmId8fR5oL6HlGL3unoUbxOnH6BvL+FUkZEU4ZByVD3aX6yJ
UKh8bPBcfhb4UgPp0PhEVoYPmKjiCwSIK7BQM/OG2AxraIbP27/GpzyThTO/JPWC
oEDo6VYeZkcKaPgL6sZwKiX5z06wGY0IdbrAxDL98fNszFhIWN8qMKszHsOBTt6J
nVvj+eG8Had+y8Iw4DLB82DgOBs3jaVlZTw8rZlbso3ruqF5YvAw6+gbPHpGWWZi
wxbVsqjK2Rv445w2wJ0OGuAUQEO2vPFLLzdnGlR/RjIF0LQA+u5cp/GobItwhC5w
nvV4xAAEREZ7IsUHJ24R4Imlsg8vdyKYaBKS4JXHDk+ZigceSM1wYzjPxZHma4CC
GZVIgM8utB9zXmD2xMB/MqfiqauMVg+B5V9cq61Z8R1o41yj+HV0ykDMkvJWaTbZ
x7y0pkgRMmeeQDFk00egiXiGif87yalKFVjRGOiaW1VhTfFOB7mpmSOR0FAImUx7
oESPg4W8QlG1WcEzfAIALtu7MgdxNHDCxSo89kStudwK8hD/ng3ROXrHaRVe7mMB
3ln0X/NE3l2FJNL/Pqtn47xbsZuiSAKxThU+84uKJkJg2GJjtnW4BJyuM6Kw425g
jU9ypqlUZm4YsEL0JTRxpALXrVlie1KAuHDMUeYHCbPsX0+nADimnINigLqwv4YP
y7W2Y2uqJHc0i9g9fqsOINj67E6itCX4/3Qp4ka7UbVQwYrRh0AK/lJilai0NjGf
IKqxsb6hnHaTt/TNJ+YowzHCBrP8uZx08eU0vnxg7VcelUeNYJMVDinNzbKUtcZE
SFPnQaGoW2LkAo6zTheXwCMP3SQbd53zefY6snEAaC8cJEUjr7cW6IQDTLLokyLZ
DUBijTOg0aw3O58iUczXMj/uVeyRtvFDA1/kCd/k/f+ujNV9eerZ91Ulk3A8he5I
/ytpuJyO67OI48r1jbE6VY+e4YixuCJPKxq5aD3E+P1jrU++DLo/RXSv4g4KEwdW
dM0otSiBCZoz0KkeFfp6gJ86IY7Y5gUlln1/5EWEy7/Mi+lEc9uolkpoC9sETrdM
lAeLEnoLNXX+vb7We/T7qC4hzDb9r/3MtbhGUx5lT9CScrFS3x7t1kC1J7XPZKl4
VtiM5VtCkwUPY5mYqseM37ZSVqfyAUdfaikvn79Qx6L0cSBKq+uysk043HQNKy5a
yg2ePvagARY5AWGtuRBdTu772WmVpjtxyoaU5SHbFkazB/G+pW45ROZzejo1Iqip
qn+2AVBHBQAovPeSM4mKEfuymeqBEWQ4v1PMfNjPDdbeohEVh+0jWbGi6ECWJc97
LOH6Pq0vHXWgL4dyq8viHFr4GQNrUqhiAQulBYh6kPkiYM72slpJrpneIFDx9VSc
xkNZNfh4fC4dyzMCQ7D4WpfCFFvbnXbR+NlzeBIrsEcqdoT5nf1XF9cRlSdLm7bL
b//LadAbsZ6uCVxIPv4c2DEuluVdKLuZqLoFhSiRwGqMC5KNvcY9IfxiubruNZMk
8j0lgTEba2tBoQpHzsZLuvyD2rUQb2kIwYBE8K2iBfkYi5Qp/Mgpk82m3xifQAm0
hsRCxwKoOPKeDg+nUG9RiW2Um+68sMmaHCCIfXCHPcObOmWQkV2zeoJPP6PRUEbe
VG6OrudjN7+uSMJ+KE2olPEVNVpnINZqHU7g/xuUerCgEIBePu6OKPDJlI1b8OPT
Y6PmRkKnSHE9dXc29KjlfT8NuvucZJpuE/L2oVrA5L81cakKBbkLlJE+PFTN1EmT
E5LAtniV84m+7SJJNiHOwCUE/h2xZw5D+w/AyGT/Pw3GTmU0ZC3Ic5FpR5QE3q12
fogUnjWBF0WcfsOT3YBXpdjpCXQLDNzaPGC58KK8OuRfj7nzpZi7sjEk+xQyfJPF
uFKvrYNFfAjneJJCQ/V4Gg1S4bOdMXKDoRdQMah51g+0koqJwnZRfBZvLHACKlS2
N1gbttIJ0qrbvuodmX1R7rzgE8bkG/vb6UBzNZEYD8k6b3hsEH8q2zZXY1DEHME/
LlWrBlOTvVpHnF8+Hyjeq5G3z4bodqP46Xvbvqufe6FeM//G2b1X7eFdUpOCoweG
hNSv3tjCIEx952OOwFyNEI3YZ+WTVHj9NdYZ1nCX9SbbCfVWbedOAeOYeQ7+nxgx
WIpOJGNq4iT7SDUT+ryqp/5o05KFamumLN4PhVPiuQYa0y9w60gek9pZP6D6hQee
W8+EGteA5zY9Ty62fWIJn+qARmIvSH6EXRyDgl2FSYR2UXW/WMaWi1aL3r8RV4Yl
7H+v21zAe2cd7tSybQeTs6gYM1WLbeKUX0LVX6qU2Va5WA1Dq9eWliXu6y1ttL0+
MxySMnUzx02ECkGts0ST0y5NOGI7JUqWXo53wZLWTg1luvgkFHZNWPk8FBUY7E4j
6wnuGjumvEBwWji4c0Cy1tIcKRNcBAx+qUvNbQbAVAlUyukLT/Ff7xbukVfvShOr
fxfBqtZrb4a/Rcg9XSbfEaPNr8aJ86jox+rYf9SxgCOrJIV1olQCBnZ7/bqcSafg
vC7baB8BzzvhC3IBCr2Tys8qpxhg6Qzw+VwRSTWrJxNHb4P3sGVEXpgJUoODqydE
N/xZmsyL/V+70ZGaKWUdjd1l9kOhM+E/thG/Xy1S5mNvk1qAqJMkZGTtWGnlSEXg
GFx2TZszvifzz2sTMQmXwZLA62VJJ97nUxmM5hLGVYSc7GPrnekxSNK1UinJSdSE
GMdkMNr+/0/LM97JYOzj9qxp4fRaEExnfqYrnOEsDahXEGh+7W3wmhfMWQQHAjMH
NZY5t0v+l1kg0FaZat9KiwlQuiXf/50a70s5FapIODHt0OrxUQ5dxZRHPEBgtCnX
ap/qO77tWlrm2HcRM0fodl/WZBei0TiPoLqXBvNvEI/fHM8SDF2YkcvQiPPM6pUw
WPqHrj1JPiAWST/z081IGYu6dFEknzRX1Ey17eDHquNwTbGiG5Z/QJpQFK5B0zHJ
RTwEK1YlwP+KQvY8wCU5I133uWMDPUqwe/oks+VlZhr3+15zRuWFziMhgvtnQx45
rms+mPgWU0NkzH6sODMGlGxmpkx45CIO9GrhbQJad2XqqrxC4+71e8Nanc6NvnAG
JjLXoh9F4z19nQgixcdToS2PgZQc+Zpi8Egw7eipXDHy0hukt+6kiUOxjqDD5RdS
/wR9px6KisIVX9T6685x2G8pUsXp6B13M7K4CRiIZ5J31ZsC8BN+NCb54BCmpthZ
dmsRUabMhu2jmXc66dbi53BpDcDt6txEbUHTv7yyzHXUNIlkVkFmv+OH0Z5fSFQd
y+ib2KJUVjeki83EWik7ctxe0SzCanWks1tbbNqxEivhxznm4bvcgZUr3lTQBYIe
Dcc9rbDh9E0nh14cQI2rhbfAF4fPFqyzO29SvB9uA0Ppk4bIM3gdnKLIH+s+/Jz+
Es5O4whSy5mvKyf0NpK5SzA1SZRPxgjF7qXXs/TtzBvNejUXLZtlqbRihlz/fcuA
8uKD0+sL6vmjOT9UwlvQzGFlfkpeBqsK6H9lNFBH3HtzuRbCSND+AShhb12sBwtA
rWtys/Eu0CmP9xV2KELOjZiIqSjCL2AOnjTnt4EjHIl5GUMm82cCWmyplLj3KlCu
gpTOmwYqL3i1iiL1CTVRM7x8irX5OyCZSFTFq/6+rD7i6kAVA4PPJgxwu2RBzt9w
dUxTWeA70dDNXggw0qM5/0B1sYaphdFOkKgcLFRPzMh0kVtW8ihknwu/w0RBZHrT
qoNudtDxCk8Az5pjjzzSHgZvQ8LfXgYJxkfE7et1vSOIXLk8HgkZaMf8nbQTv+CH
oM5GTTf8TnWEhj8ms5JJfxqPXAW8dGtbOk6DZD/aBkpzYSbyicrCkfUTbdWXMr+a
VE7OTQ5llRhGe55xNAkHMUQguzxh68IH3kR77y+MTGA812dW2VOP9XJvdtp1x9O6
oygdJubSCJviH8+9nEP5xl96WM6QM5CMnUsD6h19ILOFWhB9be2l8nHxKv891yBA
k3VH7HxyOpnP0d0o1AJ6HYqJTW9dJhDtAEG/A7KDDvS7JT4HXqY8G5fnkT2sjNw6
1o0VyXLGYcVjIDz0iL9bkO1YSiKDIYlG/7UFeWi9wSbBJf7HGTZS2Qb5SUdSyKAQ
5nGWrpAk84/MuN1Lc+VDDis+/NbAuFylpwx+GL/T0veI9d8qccHfz3L7GcjYj30W
PlgAykGzozaExbZ7w3yIHclMIQ+mrwLfGa70iV8MC/IvFhEWPZscql0FPN5efs5R
kRhWS3V7baO+ySWKcQc9KK98zNyVYWF9TTr9cZ9lYDBpdsTRah4jfKzF/cXeybwV
ddB/TMz/JgNDC9UE8BZVNImQp6pRxjhJqFbm3fX4Ev7kF+GatItylQJbzC8ar26U
LvbLVbrbUSxmrB/rQ4GzWGwqi4Qbq8F7fRfKLwAHVUF+2Y6kiDWTBehHcLxGVcfy
HnaIYy5lvagHnnFfbjY8uVjdabcTnbZWJooIg7hCGKfLg9eRb7ehkQrqpdyrand0
zgUL9cbKRde7NHEW7sAIetux40Irjamxogo7KJXti8NKK6rdBs7eNEbPqW02QzkH
6QVfN0r6sSpy0Xc2pK5bN0I02PD6nrGSqF16nlTVOJBmMAy5fXKBtCjeN2XA1JXV
O5lCBwdarS1HUOqHHnkpZNFT40719ndjbO1cQ9ulqOlH+3P0tXpYCr8zgnwFvpf/
vfpK5H6CWATRhAGGCxf6NaJvvLBZjddyOtEU3OVfJSSqLmX3SrQpizL+mvTnof3j
Wi/AbnD47KkZP0qfxQD1OY5l7INrZAVUCrv7tO4XybM6i6pbn7YPBKIF4Uq6jSAV
ij8hOjOUgPAIyvKJcr7gSFg/TFN/5yYXQaw/Ex/VmcuCtIjF+AsnEnvvS5JEEC0N
PE2vE1tcNY5UO75v3yOazQnvRr467swqkW1P9I/qPubTt9FZLT6/JqdigCu6d9LT
IR9RPMcLE0W69E8/RumbRpA8LgfhCoiV/1yL2u0k/ALD17ZdUk+8B/1qLAsWg6v8
bVNo8WZO4p7ORjEqr+MIIdmSl6fXblPF2jDm2ddud4S9k/o1t/WR4bTsV4e71BfN
tfIoJoJ3adXskZS9h7lIshnAK4/9lOWbGmSBUKAN0xrYPseQzByfPqxpHyBkznmL
7BPlqzQNkL/nR+MzzjTwDVtjjKdwhqQcRlxyp99m9VH6OFX1YuK39HXi+Bn1dVF0
BOm5f9VEHrj1Azp+ZwU80L2j0/lXAfAZPVxKMPbq0JSxc6THv0SgZprKICUSGwdL
nijaH1gZe1JSuXCb8DXM3nL94guK5Lb1zpOv2tLkrnotlBeXvLfzaY5Un8YkNP2e
v07Wu+C7Vz5RqXuIU0meI3dwcjC2YjSjLWzcPlsLUyy9xJYG86OYO8kN5tegt8S7
x4vLpJLBl9LX2u1UZuOOpBbJzqb6//OI/UmLu87M8cNGZS5jgmIE4nEpWMjJ9OH2
8XRqv34NCHtFOihI+1RYaBX3KrWzx6I722+hgkfwfs0pZptKodEhPUt5528HdiPz
ogilqNkLdNSYMzwVXHbOtPdiGl3aC8MxofWIewf0a9KAfe1RORS5vehLPoRZDWQi
Ts0RggwUMHS3kJj2yz9aa5AfbGqfktNYuKK2s1Id77s0go4bg49tAVws+4xaOdMl
EmTYxewOLkbmwE4g10hVvIZbeWejWZNJFnyS8TYliSobAgMZQ7Z9lvblYnKGR8IF
dK06CL8lEsx8PlnpkJIUFgYWV7accJnNLyE2eSbpKYGvTWGbvhZZV1eb45nWup/0
iDzLwmQAk59yWw6b4iQPv0pJejD8J1OlYFi5HWKrhi/eDDJbzbGCwDXOdh/3ft+5
f/ntiAP6+Q2DDwxnK6QM02Kfh9KHqEcsS+8UXoW02+dOk1siTvih7xsIf1jv+sJY
5SykhuxhfndfGBSMQpfIwCSe3GERV+Dy1xVrl7de/cq0lRR4zan+oAT3f4rt4Mf3
uGhGSKEguZEpHtyR6H5ITQ6ujpIKGvG3nqFYf6Ofuhr2ytg4MPGHbxJBpKXaFRmg
4oqQPIEbPPnXIGUXu/xeLKZeV/QZ4seMFyCSkiI+pKjr5eXco0/iiEEiVE9HQTAv
NPcpLCirhdA66u+27YZnn5F1E+oIdW42HWZLDltdeGe1rbYItru984ppm8ErTrUo
sF5sSvn9wWow64yFAWIFA62bt3TxKbNIxlGMJj7F8FbNtyuoHvwh5xP1oP0M3gEP
lWxcIVDB9JdxrdXOEwwBn2YCZAEfoBUZoN7vu0wsO0iXeClsB/EhGw8SvmskDeYv
UW+pTzn2rxv3B0JQUZEv1j0MQavlogXbya/lH5GkDYjgkQPThYO+TGNzela2Y9Zk
03XIbSaYejwuvTDtP9X5sA6w18W4szgHY6xc0C+SQ4ewXsEBp+trW7wm3pqBI31P
gUfGJswyaIfoYoQAf2cJ7UjIO9z6xkHlZP2cwJk0jh+8UyOR4hSHnyExtQQznluT
FsFiuerl853p6qCNeOO3surHRpk6AF2le9aOvvBCwN4fjKeOXqheRGEAiDP63wM/
XOK/Kd2ZU9BZXe9Ih7Nz2AwXssM4MqSrOiQYCMNZjmT0cOpRhdsmMfIToXwsVDOW
xwCpvIfI6afg6b/pQdVGmDP1rNPxR+KpUpWmpJh796vqazFEQW3NuKjrGPELJene
1QuT0SxDCIX59Wg5mEWlMkHox0gMUB1kUrHhmY3xZPIswNLgET1eLljq7UTThzz9
DsgCAjvCDOSp9IG6216QHC86QCWnG+P/BCKoqqj3W+fwgUxkzG4oYF8Z6FkeoJJ3
QKJQGsY6dmQAcNoe+eKMjJ+y3+XbYXS8LGhjgYk3vFcUWcInjXeffTkCc4c33Jgm
2UcHPlYZAFsmomkW7q91r2wj3yBB9Yl4CL106J5Jw+K2qX0+7bAJkuaq9/iutdUa
9N/SJaHrvYlfH/NigAFxgna3c+iD4tv7vmbcuZI7W+lQxE36HxPhvcsrZ7sSAxki
k+qajkIyJ/y8gmP9x841Dl/CaQK0GOe96/EyDkqWEzDgIcgs+TjvlpNeVrxnKzn3
1D3zEjxP0ePU4FDADZNufa7WmE+pcOqsVx0iJugzle5+Cxq3t2GQQMq+61zmD73g
e4MSFowFMJZpjOT/J4gQ40Z/lSt05FrRu598DGK/O8coE7W4eyxrtZMnY48fvvWT
tZVZI1Lkn06DrFZ30V7GsFg591VtmxWD4p4W+gPdKZ7wofzO9vVxWWCcuZYJTp5C
ESB0ZhjZ5guLFwxcJSdPAOHCz2ZiKxCyPg2WTwR+mtWuBMmx1NMsdQujdgTgj9mY
Gzg5AKBbK4oBueGyz07/Io64+Hn2dN7Tbr41ThZbi1QumNr0R74y7d+i3qZC3Qoh
/dn/9kxvW8hmYKmyew3A0qQ/UYSRwQ4N7/ahFaKETVdMHQL9ozIG27Lbbmgx1SIN
8mzHOWpxQzQ8L8sWcRrEa8hMpHUk+E8G+red4RU1kmWMqu/f49QpWuCVRhahnqFY
VWKuWu53MrnrqmpWGCMHCTlc/cOH7s6uz8ORkP1U2brgiwFbw61ZDxAsAuXVwhqj
OPfIfZAb82EaZWKeXccSPUCZbDykf/JjrdVeuX5oitm8h1M0aV4pEOIURhiio/na
Yp3mZLF8XFQCYcOy01Wxo/jA45lur+EdtNcD2MadS9WYpCCwI7BEOuudg6FQ0J6a
INvO5WvzinqCciw83ltiFFNJKj92FPR4ROSHnGtr0mvSWFScuHLBz67oaxyQKCXM
/ZpUFJHOjvltL8IjU66smjys/uIUSv8w7ZZXWv0BaYBjCQ38C97lh+11jo6RSTMU
o60InyferHi84IUhadxNQF5p8BeJPjHS9sluTyEFHjlNalXj/oF6V3GPlMT4zg3q
cVv8PoDwCM3YsiP7br3FwePj+g4AFVAYb9reaijZ7tu4yY0DhE1pgm3V3T+ZnOwd
m+Pd4VrhM0d7RJZKnst8nwn7A1APjqa2m4MbRTpSV643vVYvrC7ImhLSMNAOC9Wr
O+MFVLC0K1/svVx1Q2ieMBoTQjPOf4mgJ/O/XVhxsGjbqxdpMyrF5TaIO5a7KrzM
wDv48QkvlwRGemG10ZOsf23TPpbXIBE5odjv/y5RSKC5/dIaIq5ypl2DVZuIbNYz
6h7ndXEmZmsMUI5vUJPigzRBwWRTLYZA7POG0j+6Rn5t69+fPF4NfS+JW3Thfoo1
W53BbeYIfJ6pI2T3WEWqthddBujB2Ltin/W8Ca67l4UaJzF4ke1FzmbVkAMVq12S
hi5evThReXNGHZxUYH9o8rFb7e/5qxGl/x5zznPJF33DYbjrOVEItSG9GHsU3Zq9
fnAtO5mlKfzyn9+Zejo3DzHPrwiVjv683YUgfqEb5GBWOhvop7PfGWtSWxISw0Jt
`protect END_PROTECTED
