`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AdzHKu3DnsI6f24vd4jxCc+jCxLuikMwVXi9UhP34kx2DPwd20CSD3E2Ft0nPbVf
k5NP8eY+QWis3gtQIWfHZC/yt3EaHisFBu7KyzCbbrcF1N6JkagY80GwvvwE+ixU
Y1ges717MAqxc+gLlY7bMc4KQom33QcKMJ9qwqZ/F61vqlFGPdBJxn1mQiEaRsBv
wQX437oIjeuguXT6rvw+v4O5IVLGFknOGMOziyKayO/byNasZjYfOoLMQWg0MbwX
fwrmpH8Sma5NmJycxVq3/A==
`protect END_PROTECTED
