`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WCPKIhA4292avlceALXVqZqhJW2B+avrGRtrxl/DrMNSFu+DsrQvx51CXfehG3n8
dxX+qjQv6EYbp9VXsGVlOdBDFNTENN5oKYUHQ/HkERs0zG3njMyUVhQMY0ZuWQNH
lCKN6JffXfDIHbCgLd2migH5xOespBlyt74xe7JkIxV8M9BLWYz9W1bEHyyQ++l8
85qMP82h2IT0duAY//TgZg0klu19BttEvlNtYrA3TUwR+NDVfVM036MshI44Lb+M
+LUgP12tvPfGFcdJK0b4XsK+0FNx98CoB74mJeZT0XjxncjiRvOYSzFhN8eXfy1g
G4zIUd+YBtrYvIS/QrADTTU1uI92DX9EBrOJsqwwFzN5+bdpAwD22V/87JsPgyko
hG0tRDlXoRrHcRUukMwGHIgBRRmp8FpZadqECy5pIbTVC50CvHFEmo+aATStkzZC
gIxAcxEZtcLsLpYv6pZaJQAl9h8yrY4rwZN1I27emGb2TLVSJzJqYifKgUN6qzK8
Hf47OaqUB2Ng6UuMHCDw43kkrGgiI7V7H++AJApn1wgHb+h2oFSQwKZ/z5wKitIm
Q+qcluboeUtcw4M+VdjwCnIYff80/Q+9jYOcDoBHx+T8UCn71uchIWXiBY+4z7j0
LQCT6Ow827zvmI2VsaW9RiXNfGlOzXHwy2ObH5cJoQTxRTUooTlvDKTLMu6d6VBJ
UTSNlL3pjF1VSiiorMBt87XJKCsF6jJ8ItuwnqF2tdjctTSVCQJWy6zTtdULdJi5
5r+pGSBrCAeMnuyIYFD6lnwoCCsK55/e/JYaC+M48YT0N2dF8iDmym+Ti8h+JWKA
8nArweP/aorgYOUqwEiEyBJ7eNqzQyPva4k2b0q8i2stbkksEOF4gfpgDXtw67CS
mCS7cfopH+V9zxb9snO8h8enygxCeUaQ+/wb23AFcKFRo0B8Yev6NHhoakVliC0s
AVk4NhcyoZMEhbhPferBnB/2/saeOFGgk2rc6Q0rav8=
`protect END_PROTECTED
