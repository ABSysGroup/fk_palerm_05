`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xPsaxR6GEY6147/Cez3D9Z+ojWXvnAmT2mmg8GPiGK/YudLa59VuGkZaf1j0HrlW
mwyO+nNYIm8+zJaXpEi8hhMoeiuG7UUtNMjkVJIRShCM9M8efsv6WCs+eRtKiClL
wOKnfcskNpYW/lFRgpBQb2rGDRl2oRsrm795dSR944Cr5RIiZNOYan8gZCX0pyjA
6C6XX5/jmFN2TqYQUEml6skBlkuWWMvPqxIFVW4HYYFClACEWoZe04k60Yzs8eje
e7Te/VPoVIqaPvxTl1R8TUtlis5EuP6rEOkUKPfdUKAFluEKXjNc+YiSdD4YvYLs
0w267964lE3CDhIdQYm7sYqQ4WbsHiAJW3FswuAHsWCMWIh6p4B+m3nf23CoiHvN
LkXhTZgr+aut6+t7Yr+v5O3i2AQA+E3WfU1Fpddm2a0=
`protect END_PROTECTED
