`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AJUKGIYqlEF/7NqGVsqOhfma5xpYor0Lu2C4mY6xGl//D7P4j8SiAH5HGFCm9GYW
tX5+oq0QMAuCKpsINmvip9gqrjBZAk7t3ExhUWOWxCRll2CullP2zCL4YAX/9vNZ
Fhygbk7LTn5C9Xom6EaGkPosEZiSXvOMQMZzhi3pzcLMRAjaTKcxyqWOUIAK32U3
kGO/1hPx0xmES5ZR+gYtDhT9vtBnBCa+4MpTBreYPaLIjr1pTeES9SuN4oHJazBm
8VBCXPH4TFodD5JFs8VSYFg+ASJZu8bbC1Ur5gT98th/GepevPfaDJ2OgSO1nqg3
Go5nIAaBIg3wDSvcSYfJDN60JRV5Xg7yWS8I3kJXKe4/VlkkiIPj/ZRnyLprmLsU
sUcCmvGNUyf37Hpz4C8cN8qlPK3H7AGKhFtuPjEmR2gkBcMCLWXmZkCFAcpgeIhS
e9gCIhBqHJTm1iILNUnRPstfx1zLR4sz/yE2sOApDzuJUWMqjOjkoIOO3CrpxZfa
6FNJQ1RcSRb371r5h4YzinzK3FPFsf1PolQ3yWnDQMpZB+CADIvLK1iapLO3waM1
AkyhPNIyPKbLS35f5LCtrX9+X9CiFG2WlMnyf1/yHtlAZYKnoNnyo3vdFqH0rDJN
lV0v3+V9rv03te5AiqfzDEzAZxO6ba3W5K7Ry6z8TQZf4KRtoR8xBwVEre2Gzgn6
NiXlwukHBesp+epbqGWen4PKshHNrLNyr7dUvHLQs0HzDUIpq8YFvtqWM4ORZZ5G
ddnDmtDIzbSSR/cPaWEhFwFTr6HYjm8vp5HsutmvHO9TVI7i3CFeOV+gXCXz/5Ay
bTEjLThaLlWiXkeykfXJkG4tmk1rdyjOCJum9O9InYnIvM5CPv/obOd3Drprf3jv
P+h+8zg5cI+IIzzZUDMd9IyoE6x/5cirFmZNKq/d2YpRXhrcQB+KnemiLh2i2FE+
c5r7iHkn6BrtgrbGLFPglEeZb6lSVNbdoVRHDOVrg8g7R8573aS4P7XKJF24xgi6
vraWfraLdJiM2TUr0K3PIGjjY5fgBra37oChMvf9Z0QvWU0JtIFQUg97YiNfqsdc
3XCd9HVprLoSFOUzp2aSeQuFHOejMyP7sTySTFgebpF+QmRtK4B6CpP7x7WUwX67
laSj4iCcgVAO7P75Wad/5sQ4gTeyNIUZlezDeZEEfsRysjfh+IX5T0qXBCHIn5fh
a4TQogLHdUbhcvV20NHT0fKn6GYJQ335/eOZ3dPKcTtcemOgJd9B+NcQWJNvTHC5
`protect END_PROTECTED
