`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
30C9gu146BqdjtgAQKvngTqRAg6HRm0l7f8o+Mk+Nm7e5o6SmvUbG0Btv+Ubl2hs
fVf9Gd8/KBP+N+tsde1tAYH+svM8Ln5NY+CQFdHxDs8cfDd7HUP/YKI6N/uQp/iH
6e4dJFvn2KMTjHniTsrAwzJPUFDKn7z+V/f/mVb2a6ZWcbCqnIO+zePXgSbOWrdF
NAMEfiknVi/O0FG460uLygLCm7zGj962L2tn2HExdmBwjRY0jWDjou84SYkc4yag
5bjpKEGZXyUo3EQ6u/c8UdKp8bP1J+lCJnuWDn8cmFflRGglGCXd7LbDdrLVHzSR
fZZAbjHL+wsA/uDh8W9xlA==
`protect END_PROTECTED
