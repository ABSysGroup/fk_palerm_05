`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zepEgDAhRLSkwlbS6AUufRZcLuTIWRTi1wJvK0E5LuvV6A9h7Agv9c89IBPAGk5D
JoaGsDFbunEwk97BkB+1Nhw3arRsI+iv59hk/qlGSS5TRRXrreMFVdkEZBV45XCi
jL36ecSloURJvLyFvp0bRVMGxSkKPoP2uBQbzR8FcNS6uop8VKKvNIAoSxG73NJn
4cXu2N+V1QKL9yqHarS8UCEyBxceZVHo6pikJHgl4T+YwtyJnCk0CTxHhB1eJfPl
WdYgD+F/osMMd0h9kTRHT8/oHGm0OxIBeHyEvlluOxezRsK3p+n9U7xWvjBDfk2n
sHj7BRh3qUCgMkM0aAtg2AxTTUMhLp4ld40i5JmwF+rtOcwcMq7w9M/C1DauJAN2
+ugxOh3J4pNHJiz6jiR9eWzQIUa37w2pUj/eYObXzVVWn3qVDeWdBkt3NamdkkrW
BM8gB7DLjuv2pLlFPJ71/UCe25DHJXov5IdhyOFm+ZhTeAHPAm35a5J9FvBIA2li
NgoKsq98p0Nr/oHVuOKg0NgTc1wWY/AODYXFNWCr4bxejLC/mkDtqAK7qV25wqUQ
TMdRTx4e5TCoMpmNPwwNqAt34/6C0FfJcoARo+Js9SSbNfiD6SRDcrsUEeJiEF8P
b/XZrrdJMXxsyWXwKzqzcr7gSnU8Kp3ApxnFkloXV6FLY1IyJ5R6KFDt2seCeLkM
fJz1ygSNUH6btkGP1FC+oNvSomiw9jl25NOXUehM778bkn4h5cGtCizDQB4MDo1Z
VC79RLLK0CI8PcmiHVWD8jOKfCET5Our6ojDDxXrV4modE6FzwQtaPJmq0BZtEn6
PY46KxSwrXvuBk//jfb8EXTCaOTCDYEECzRrl1LNmH+LGFvSDx5zwa8oU3LgdHC6
z68BysGGkG/kIRO5km3ElK+APMZt5lmcsXkCyJCn4l+TvVa6iF7bbLOnoL5hYz7Z
sv87P3Lo53DXFn59m16RP9eGPpoOBX+TVIS2cWeEqVyI7Oz0YUrb25EEyZUQe2s8
6QRyilumXWg+OmQgNzSWovw/RDipolZmNZQXHu8i9d8pc/btZCjLGTQ9BTt1bVdY
g9TdQqxkq7FP83Pvf/EJNdLiKiDi30ZACJBGJGIG2PKXknh0q2Da1X8J3WF/3O9t
jfy0p81/KWNZuWMt5TchbZCibRfAjgHCH7m/FTF2NyRlDBRPs9TBbo+lqctfoq+M
fyFGVSGYQ0A/ul1kZ5ova7Oqbh65pxoyYywcW+pC7d5HoqYLG4EndqlXRgFDBTu0
t0tPxqpg4sQftQHsh6D3rNxFC44ofZVSZAKa3dujKBdS6Z10qG3HDCQV+ENLP5Un
HcnbDGFQ+KyWYHNQcbm+Ttt5+vsGMDm/nVo/oG59HxiS4lt2rxPD2jsq+lOO6adF
c3pcO7VZGpNWTktqTDbrKw6j1gdkUii94eiX//WofIKEG7LXxLhShPZuW18L/m28
ME9J2WM6Mhd5IqP2sCKW70P+z94kLCyvbT9pb4fMtZNvWkwoWoPTXV9yFnuvkUeh
hXRmZjOzYOMCbIiOIPm10qM6P7AiXn/Fe4E/U2WxkbupO2hCW9CLhVBnw+9FnkKR
hVPd8a2btE2WceVd9wz//VT6dWz5ML2DAM5go7OWkO2SvrTyaFfU32Abk8DGE6Es
Bw2hD3kwQDTliIxb1Nc20GWRSg55Rj/fsw1ZQ7yICDGw/QjFMaiflCayXC2UVA9k
GAD/++s9WEwbGe0MYkX73Ks0n0SvS2gtKrV7wTkbrBpwU98Oh75Ymc2PET4i/Pcx
Osb967CcfzfRzISpVRtiXWVX+V4KAu8OlaEiWYLmrZkRpjD8Fo9Uc1IJxuovCyw6
iO1Kxb3GjwwlAwJnDzWiYpKBIRt5oaQpcnSPP9eWldLOYPaQmHQcDulG+jPA2Vno
xGooKRUJayGRq4aF6EKBmxQiubZ9Y7cPxg9idtApqiSTBIRUhWqU8I1gQzTv3gCj
Hu9yJ+nwUhxVaUmKlA0g0nZ8f2Bi/gLIHkUG3gyL+vkvMhJ4MGNzU5/mFQPKLEz7
vh7VqivB41J8Mk7lngsNlUlILX8+u+DUbEQIVzcIM+y6cWb9hFPQV+FWSvWQIaaF
kdgQH3Sz6BvPpCs+Aaapf1lSiz5/WQbX9s5WdZoEYos7zYLtPanNHeXOkrHQs4dy
Y8H9EIRu3aWSloTkB9ERVL/3IVEbLQlHcKXxWBRLy1OAsFZ2Q9E3FCe1+Y7xjc+S
w+HqLcvE93kNivt2lGr+5zXw/qStZuA6Kya44klmAWERimB44vJs0MmUKSDlD+XF
UE66VmNVDJzrWeyU1UcSF+hCP9Az7SwEBZxcKjF92EG/wTzbZcnsjETI5bnPAR9b
w1z+8iJhmNr5+JwGONGZmYNPg/2Bne3Og/RVFayUp4eJAc32iIvSaBOhdRL9EUwV
jHr5IDFVfCRHE9CwIUmzNbibNtLJc32ERoBj2Fc+lWOLF8PClP/I4r/sV6oDANF6
PXgkJ0Ri9JBb6C6cFYnCv4mjH5dTwM7UsMpqCI8G1i5YFeXLRffslNT7Xt1wMPMp
jVtuCrs3PaeDHpr4vbGsXoQoSIoQAePSq5DqvBM0A8uFpYtmWL1lLPsj0Tfli7/H
85UjqAxXvftQCshQvJpkRBhBvlRZSNZ+KMkbJBggbvr23AagwnT2itY+GdUzbnuE
uLBBGyTOQDO4e3URP3xNwkH1trHHj/B+UlrrAbq6roY9Gu4uWKyYQtLg/Z96fR4k
RdkclJOsF12jhw8gTYyDz1XeEt5/U1zwDZ4KeilioVYdiBHo9hoHEzvNvy3MkVHy
/tA/1w79svwNn9l4y3cq5KMWKJ7zhKc5lYmg7vq2hafK4pWpRHSKgbMNlDSVL6LF
PC+0gwF5hmbsh0jcLQ5Sc0FGncHMghCtjjwGgNZCPefG2FlVLTygYXkYKfzW7Pb7
4zDoZ6srvfbGWX3FQqvtEeZXNrnc/SG9YKPtK78mohqLeqY0QTJhKxmB13TxOsn2
l7VzEsZTc9OBFZr06CvYCUhzbFcQSTM+cUL4IWAyGKl7PmQg+v3GgrKKQpAub+Kl
yVjGzNA/ZXqMp++gAFzZ3/61BEKP+mqt/2GEk3YgHhx4+Ga2x+vHW6ORKmO4LkIt
4SXo35RDFSkexA6jI7Umrif4TGcbo35u4QUdfVPRXvtgMkNZtEMkqJU9/IAfRN41
TpUycKng2Px9pKl+GsTQTyKLfbKJo8RNDST98CDM0oqlcnxEWJ173aZoX0JzfnoV
XkkPXkjxqSzHwdpkis9YJZaHSIZ4dGpiot9J91YwMofCx1FDYsK517Md7HmHnhaT
Brf9nReHvp0HmJ940q6Yk/q07be9SXNmBhpiLlzBx/h+b1I3UdvLNp1DrQow+CKM
T2S4MfGS78PLkVCfbkXm4CYIhY1hiyJr3huHTPL9DkCY4NXakvGxNF+F+sCASTUc
qlQ+J2zloi3H8Z0p4NitSKOPyXM1zL9QzxG4WRrgrGdWGFYUtRXV7htGi5oa4CmR
A3AdPfDX5sEJG2M6R/paroiYo15n/y061jWsD2+tPnwVk9uQAcOjV9eBjlWaCf5g
8UR58nJ+7PCIEGU/X6uqAEy0zCoflldQzZ6dOpyLu8Z2iGQHbkmLv4EAZfINE7Pe
6ZJ+m0ZOdSA691iUBW7HIkhPtt4Jzm8DP3sXnI3UCEGT3m5j2hylwFjO6RSIRCya
qfCMSsGI7xem3FZRa6ETYrMUnAegAPXr1Xbtg0CEtkqmYo3EfKew+RTdAIdNEyrQ
Q7KRax2wAXpVGYlWaeMXbWWWrgqYVCKRhxzUkgKmRe/T/k4iHmoIwijGVXBkizOn
170IZe6+6nKKt5KpJuvsFnrHPfbZsxMYowL5TAHarYUsm+iG7Nx2RuNG++ok+MQq
NeUXluxsWHbB5E3JUMS43zi1tQmTK4wvviKOWZVDQ/IQXOJVNbvmq12A5DzB0ElW
U+oz/CRlCteqEowZH2TxhTTcQ4xYdO2gFe/3EhW+Cid7rs7LVSLuvexpQJnzh03K
Oa7gjtJGN/YEJnlU0ydAFBtom48RpaT0DPfqGoWEWIylexr+khUuu+ks3fcbS94Q
/MkT25qGyrJX7O7PhVj8mE9gyaFfxdCrTYPT2lmf1E2VtitizBe8DD55IBLxh9Sr
2dCEXoWbOSJB4/MYXvTLIbebK5tTjzNqcBX9sWQeoboGGpx9p/PAanZRVhYaC/aA
AvtYG4Sms83wknWBL+0MObYlzG78cAT0Ro0uB5yb0nAYtwkehGQrmGyc5GRf2bph
DFInzRVdAdQvd5LmpwwOl2LOcRdhOL8yF89McEaS/GEf5jUsZS2kcGP47ow4/Hq5
BI8bLE/7BbtvOCEif3C5FnjOtOuM0uAWtTHnkSXkzykwP6KsKpdQGxR+kpMBALzZ
9d8LlgKLLmA/8esdvvAWz3OneGmJJ5Fv45HmK9pVwJdChFyJO59dGquvK+6yqw8S
MzeZ+nOMiyghph+U1M2i3pKkwpe6UG9VTIu8jkem2PMw1oH2PombYw38dTPOk6gG
+3P2tWtvc5avS8cBV5yTpdpf7VjBIzv6ZhBQ8ETmx8yqYjLP5OG7vNV7NQx9CNrO
rYx4UInicjjwRZkxO0UyFTty2/YwJxil6r4YJNtanqnZooUUIBXzX2yIfsyyK8f5
sMynfhYCdh8/fvCz2hGYKQ==
`protect END_PROTECTED
