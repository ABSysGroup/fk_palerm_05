`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+c1SyfkzYs5rCSWtk+FRUrnKtzMzjNrH9f7j3hgoQmrumxTtCyU/pE1kkoPMZlv0
MwoZXJIc3xnxsBguvFE7QuxqSfmYO+HLGetifrufSduZ+gbXEHU6mxXIG8YGbFh4
tg7OojHsXrgnecXMmWYv+np6zkkzLAbR5xjOAdE5aKI5VNixm27d59Px1ZkID6/G
ZHenXnDIFVO4uYs3tn1eynvJkD2nJN4aeAmDozWqaERErks9NVvqGp2IKRaFFaz2
b1kYrS9PC5DRtmhiqRFReUrLwGbpkfNedj2sWxuGFl3hwi/SAh6UijjF/gS8FR+r
d7rY62vQe5cjvMpUPkSuIkGdBu3M6B/cDpuHLDWv0LZ1qPkV+Sd4VfGdNmLsRdCe
`protect END_PROTECTED
