`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bVu/piQGb6YkjliBZ2qsWBO28EWZGoU3UNV0pZCsmsXeMoWoR2rv2iUJyh4+dymd
Xz+4bGzC9/ZmgdGyaxNSRKwemqqjmgAdE+X/I7Ux1t9pX8/a7Zc6Yrv6IspSRrVH
M4OhY6QR04MQELU3NmP6K9A21nTEZtxP0XSnFeS2P63e2zf/cf4L6XzJ1e5T1W66
ne+N+L9JkJ4WSOQg8ruAMNd9UVfaQYpc+FC3pO43dj/E+q9Yf1Vhf+oMdOrNpb90
aJixf4oMUWzJJuXkcEY7A/K1JwzE9x+C+bovNWo4H2Nf7imgElVewA6QdX8KMaQB
OeAAk0hfQdyXMlYUMungqw==
`protect END_PROTECTED
