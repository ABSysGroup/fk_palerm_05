`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+2unpmFYfN8lUI4gNHJ07tgCUCZWSAlabENRqt+o6jYn3RWaWbYG2Qoj6wVVvmn7
YaFfzwHpbfO3zopKM7N8F1gz+WYY8/jrwH75oHF/uMQoUgXYc+xVQ/YO/Af0E6tJ
Q4fhaAzmree5xD6HBCXEpTesWe0td6FtpaZLszMfXwFvtoTF0cI25Qt8CfUin9CS
faIr8CeeJUq5WnCrEWp8UWBWBH099Me41se9xqBenvGjGuDv8b/sOaFFeCdLe/JS
v1z42WRo1a1uhW2YeH6yBy01BY3r7APs1ibrakSghU+LhaGJ6NIYp73nEaOzGjen
ppldKaJ2f2IiJVEor17qMMosOUzYMrgg/f3dTBEqp3Quqs20ersYJB9Oo4vWolLP
B5BvN/DZubBk/vLhiudTN8Fnc13WqHiUvHBoa2y1TRiNNQFRl01Pp0Kwqhp+eQld
eDwXpWvBCHL6AzOXA6OkbElpfFLGLnjwmMJC9X4eXG73AD0BrXCtj9sx7QF0gQu7
rSuwros4YBZJFagp36kvpDZq8Pk4SHx86r3sV2aL+N46G0/DntEwKxyBzrjs0XhV
UzF5jirrqjWpJGZwdRneMnrE9HrVQvHg+6bi+2gSTQmNqq6TGUsY2on6PApxqDJT
AlaG///KEkBMxdQyvy12gOLaKhfmupn8qou+mBKEJD1Qxcfbg/XPOwQEQ0E51AEz
aInWh+jgYvlNpPkLaevjPDG2Pzrsjr/hGMU3uixvAE1pwgz7x9eaTg8VgBwPgVNT
yI6oOCSmxbct5+ILDHlMQA==
`protect END_PROTECTED
