`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E2U7riagk0Y+nTSY4Kh0ZFE6rlWEGBwgWUJomMmMRQi3DmDIfboxoCMCLsuYw8jC
c77IYUlMIMcS90JyRwHIrfldMR6lE8ylwDaedBSHwciya3h4ctMGyi0fgmVohkJr
rwvRt714owUoGuvhaa1oCPJkIBljUeiDkCiZozoHPwaO/WMZYjMvEgyX1SH/cQil
4PWF7YEqjPg2tBynkhTClJ0rESFwyRfKOU8TmGCV4wIYaoldJiGs1bgvn33wngKi
w8yhbxgZdafpBqssExlQBZxuFoOhpoaR8UTdkO+y/i/OYjMwxDt9MhLiMEVPSaSP
g0/axucSQRCYmEIRLjQBMk074swd+BqGOQSK2CigOfJHXp0LLcLXGIsj4KuFwUSq
d2nW+GOY01QHYANNPs8Yv/l9Cg4UFXpuoQc3sFjuqRyjzXhVBfIKqOBI4YjPvzTD
pt8vH9sit5YIsWIGf05qDYjLpBslSCWkqZ9L3cAT6WZVLn/vddVRSxadM0CtINFD
3QKbmUToHpP4qmYJLLJjhsLkXOoqycMVBHPwgUel3fMKYyAKpo1ad8HbZl5oOD1C
bwXjfweSWyIrjVllx2mamVkGG3+aX4Rb8LMtz71kIHUBVN8YlGPTBaBkZ/EwA8s4
SfKWNf05uUmv42/lwq2/1OtvfyGZ1/U7tfeFiU30D+i430jSnsfAvNlP8GM+WSQj
EEkhpNMgVd4S9qpnbVs55tq5dvFTEfywbzKLAhwRffOUbtnBbQ5jo/dp9NckKc1h
zIONMWj1Tn+UftfBB0DfLxXAUehxnBEnW6xkwhuKZWZJAAnzPmFJHUX+x++IG+1c
xzn+YQYJBhDftk7LvzibWx+sqgE+iZtJtQLkAXfa9XyQKeof58IFWQcDM8C3TVi7
cOuxHe5+lxOMBryMZnDrPlVULvkiZwOS1zbOtCU5vJU1HCtBGGQh10GJa0UrQvez
ucgRpILFVE/nCsaC5mfx/1PcYdKETIk3mXseHWP481fB0dm65lCARzpp8Q0AIRg4
J3ot0bsz/ekHRe0btKtLlTR6ckSroSVqSQMfZcL2jeHdo6BVw1xbFiM6xWxrEmq0
k5mayKTNSl9kpdiAJMlm5Qr8YJk86HIeJJoJHJoIG0kiGyLF+WbuuP2ICRZfmZ+E
q3W+isp7mDgSUXC7WTR35tV2JFocJZ+5P7219Rdq/JqTp1x93+hTi7+9kO9pB74q
OV1SyQ/BZPVWDtn0CxUixm1n28U0+4uCB6UAKFmr/KXE0ATYIQXyS7VyrFFeeSa7
MVR0HTRoKOHNCkA7toEbtWNwg7MkvtEWV0e9ixy71EzhuFz5ICD6mCL+b5ojxdTD
EC3X/PNYCH2AkyaorO6onCs8pb38H+BhOBV8h9MU16iHZO0YZsm8A0Yzg/m4PcWr
eQVmShjp+iwQhQyETgUlGuaI0bBKJb4IfgN3dseGIw+URoKFuPIEm51VujO+kO43
iC5riSQrqUDFfLRXMrfTG/qrL/VFhevZazPFvKH0lmqkneOiE0K+IbCTB46/ubqe
rbl83Ij0NyyiuGqP532rXcOwVM6jvK34ufxxvnVWACG9il53raMSsWZW//arfusN
eVJiiif55iHu9DK/ddRt9z9nW2J/eef+oaA2KUdhmtqi4JO6SvLOyQ7X+C1YipHl
oce67DkkAGtyjEl2NZVqFREPvPZLL+Oir4Uigq3iAPKGPmu17A5pgFUnSflml0I/
i26Rz7bB6LFR6QPfSxeES1YCUE0jzApqUU6aQAns3/fw6zP3/V7zHIHdFG+4Tf7c
q2Cvv60e0Pw1MHBGzKCH8ry0rTFVJCSAf4YtPu5w5JqVLfn91FAU3fF3AAq535Ux
ggTlszyd/JLSAYzib4LMRqn3M3xhVuqvDXOU4dsrTEDLMAA31DuXIA5XUmoBP/Gg
gn+O0+v7QE7vJcfcyLtRfCGr+iDKP3joGCC//GbVc4s80K8eGji7a4o0dUzeW258
FD9nvgUnGCHI6AH0EOT0et/c2Mev7HCIPyJPt76zPLMaoubm7B6lJ9C7xNhARzlD
ZGB7dcChwehhHEw/22+b8qxC9gINRH0gFiqoLO8szGn6u4ICQ7c34pmz7vLmqiST
9U7ilrcWNojjqUHZS5dOPLl4HmQt5nsPFNczAO3zXd+bbRLDdjuj5RRwL2GVRtbZ
mbs+ITT8mSjHhGzT5Dw739vnSkKoUVoHi0Y6hQh6ehGdA6udvGFZY5ae4M90MaTM
7s3RdiokvZf84IZyLDpt4KmI7V0zQNxUCxqnMonApMtTAiKw8rG0q3UizXbb7jt3
wQaUWTIOpRObLwc8e7+6DZ12jwkNkfM40gbK/nGHzXH8evyfsovl1T4ERleuLL9v
EaQjOf6pCeJ23YSaHzSlutBWViNubcE+wGijtIq2v+qhMRdF36zRiCP5i7YjeKvf
XWTqziQiP5yi5GHyTlKAMX8amwTEHEtiqa5CZQv5KSJdEJ6wEZ0nqW7/ETwkE0YR
FXA+65G/pfmT/WT8ic71o+NW7VxwPZTQSzGHM/YGDEccs/mnRbn4BuJ1Fh+WQ9x4
YCt6a6CizmlrYuQv8NAFgMBxaAgZv/UUo4EUS0welmrAi/rQ5erAHl8oezRSXs07
F65pioUbjmK4iIDHlZepa0hBtjJUpk3Xo/D1MX9noSoMsQa6OfvhAsCsxYBAf7La
2Tpp11uKf1XmmnEBcMoyzjvz8tP2QMU4ASpCb7E+iADDPLk8RjReAhLTh3q3JjWh
+7YnH0S/nQYAJktx2Gj05mws3lm3q/dxdrBu8de7lU0vjBY3Ab1DyN0z6n02Swup
TSgPVCfSgLvzv3zSdIUFv8fVa18OSBLWydHhFVnlL94+3ft1L833opn85XeSxgG+
3gMAcySoq7IXZrXtQiyMWD7X7v9y2lDINlQr5f2uIcn7YfKmoiNXrjyyjsKMt7sV
MwSvw8I+xktZZJLV4oB8X5wR6BBNLMYyMzkhkBzwRocSjD2o1KNQjlQgKaRh8V9K
nInIJi9Y02oINDA1DZLcgMdKTViaK2OeHDuQE19kEQDYP1VstDL5PKRcVcpR4LnD
AdVf6VLC1WtuaVGpx9rzQfyYGnmAq0XoaogJez+QZR8kBdvnSo2s0jHW1++3AXfO
WC3SJIPD4GVTWrrPx/2I1uZBmotyYD5s4dccuIuKyNxB8wwVFtqe1RieQC6pA9NP
BbquvNsK2lsrEwkOB39r2MEEhuD5G083MEyh+xq87Dm1l7Sq7gGqEKK/Rs/aqgut
5scnmCNUDd45emtjUzjNGQ==
`protect END_PROTECTED
