`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oNu7oZn0SYT8pAVP2hyVfz+6dHK5kMSVryownPDCLhXjBG4DIkNvWG7wTfwk8End
+KiCOpiP44gFZvIt98m6JrWqmDoOVk1tx/AXEso1e0kT35WVnm+J3ipCtBhicfDT
TTUxGLWSKcHmkaHi5GWKV4YSwrYosTYVrOMkvS7HduGaa6gcx0Ena4T+GAvrra4u
PK3WZXM1CiN7sy/Cu/UJbpSmbAQsgCaIgoUAAAIvHv1VT+yKCZL6Ia6zZzCm8700
tTxdWFycmBOwNYL9imvcTFWCUSLx/RiyKvxBnHwWS8CJeCp5lwHBBJ3gp+eWIZCm
S/SD9O7OxwJCDXdoa1MQobwrC4i+iDydUINEEn0ffR9BZyCdrvZtbmmWW5CmLmaQ
aw7mILBMf1DWbA6cyqC+8GobBaCnJRU5QPLm52JWdpBKL2mVNWiUTtLh/XE01AtH
opkYaeTz6UVSwx/ajvwCo4UcmuConDQLceNB5xw3EcfHhBMGGj27Rb+Ukez52WhQ
zREskWOg6wxSUaM0wdAaL1hmp2Ljegqrre/M0YV0sB7tKDBLip3rtTihCJpI1zZ5
IljN0s7jbpNq7UVs79G7kpakBSVNh7h2dVRO4PToD7g8JLijSDybJFOzGTsIWGaS
8vmFUf53x+4+TIrtzsrs/OuBkZCl/pK2+Gc0lEXGAXMRCpkvIjshUdpvbIEWvcrF
3+VeIFuxxEqnQLzpUOUCSwHby8ASEEZ2zSnR8cKFk2U2fagfUpufoQxDUVhK1oeu
ZChKucq/AS+KKQlK7mRMeaTCy3O8G5XyelJ3UjMPIN7d4NiE8UkAaAdEmCjhu4DR
`protect END_PROTECTED
