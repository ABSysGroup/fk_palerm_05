`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
teok5ve2sRsvs7aBOj7yCeBU9mXRUicUAVcHAgHk6iSBnnd0wNXu+/i9bt0rrBSt
J1WT3ZbigNp/SO2btH9nqINiNKgCc7gmcoxDhL4o9+EmlUMa/T0V0aIs0J2vRKhQ
utMl/qMF3Ew0Hbm+Grm8bZh9XT5FJvD4Ly4mgrr5n2MEGigs9lN35gt8dq1jpFoL
ECnwkG7aU8PPNkdwP5jo3fqMU+zXb6OT/wcvs42aB0Z2RbFYc8wjS703VfS4adtn
THVt77nbdmTE2lShnRvBe/mlzUcLaCuskHl1nhweeSGpUDYAfra4CNXATECOCCqm
fukCzqK8nX5bD98Z1jzv7qcvDNLYS1QXYk2c4QqasUr+hf1T/g+MyYEEgAox/a3q
F2z3LBptGCbuKG6na6U5vQxsR0xSFia5e+WMNpZhuSE39BePvDJkxajOX9hvAJpz
xzJJZy8mD30eQod+pjdFrbOLBotFXW3MBJU+cRu9W6F0S0mvafmr2+MmO0O/2Vey
uF9/5hSPtyPkGI5+rDEsH3RmxeK10fNhWa+cNCbxN+/TKbEZhqFKeioGK70Es42D
i4al2+E9oCKQ0h06IymtYZM0islCgRDOgXkhaqRfqgDK1kml8ik3FE4hXzT9sx1S
HvvBStBByKGsd8+AGHPdDuXlqgxoIkALKCo20DUFd9cOehi4p7qulwBv2uU0ft+k
9tSJfDtJ0NE4flSOVlBIAu+6I8EGZ60Npu6F6fC38WCZRzkzK5lunNiw/ozbfNDN
8ntJ1ag0AyUsXX/ACd+XbsOD558JKqJWGfyzxrzj7BI+6SAHMyIicb3Gub4Gp86z
DXh0qraRwdnemB/shSWVTk7ti/zsVep9XOun1RE9OiI=
`protect END_PROTECTED
