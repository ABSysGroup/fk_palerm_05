`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oowEjxy25Wr46ETwnI1gmByvWP/AV7+BiLQFX/JVPwe6AgOSJKHYokAAN/PhvdIP
PJMhptkiozVcqIHiw5ujkZ4A+lhbGu2ymzCvR0EDODlPAlkOs9diuyToBDZ4zBlw
X7Pvi5IqSfEB9vlASoW7u8XPTHBGUvrgKinG2iMbtYzFQbsq02hvvl9vUpMTsiQb
/WlkSYTRUMC52zY4X36bJkJChKoeghasUJm1A9sc5x0XLdm7WvAslbw1LpVLieYb
ugLI+PTdL7jGuhizTt65e4E2ngbmaV15cW3Iic4rvvEoWQx3pehhsFOfz+mVLycg
gD/Xn4cWEKV59N2i8QxNGLdAraOS7jr+ySwOTgn6AMAMviQN+YjRSsIexvAOEQKn
HS2voQinB7/Sj1zNYi2Kl7ZA1sPlmO7iS2SQAon57ik6ADYVTeluDgt6PuwrofP7
fPwjPn9ekygIEWIXe6mYy41b+VXvfCaNTh0If6EIrwkw2Hj/feLpc6g3QQK7/vKf
3ql56sorykw3KAP4fveij0+ln0p/vdtOU7wPpxGx6hcMqJ8Om0w7QxWebm44VZ/W
oNlR1N8kBDwhdaxH1ea07cCQnPgPikMdfBMib49rNefKlFb40anYfoTmobXvb4Ou
MU77w9/7me+YgsaPi9uNryLlTWQUdoT9tvFEq0c1kjvkEukC2rcsJ+4TYpeyNj9H
yltNXXMdPyUMu7MaaZFqf8RqseEIPo8kNZNN+W/7fYr3VSXquh5niN9sCbH28wh2
`protect END_PROTECTED
