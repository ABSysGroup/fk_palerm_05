`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bkiw8ocgSl/l79V9h+wtS9JgJMKJ52s6MnRa+dmdZM4CqAuNu2l75rfRryshALkB
u2W1JAWGlskkAd94R8TCy7eHlnKcQI/xKoTzG2KMnmDpnX6t2SrJYM+vHdGgPshJ
gcHPHIzWyMGuZcyZdVgy87EXwM9ofkA6eh2vokJYJu1DRGRhSZINt3SvDG2KeEHm
Y8kgazkXS6A0jEPmE057xvM1x8Sbm74CiB1b62o47R+gF/8y9X59hWyhjDeZzAQ2
a90hMxhj9aYMd6hE9zGMnK/nTLlEGVyIglivizjrx3dV5c4GRXLjorv4dAZ98gKH
`protect END_PROTECTED
