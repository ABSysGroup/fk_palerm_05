`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LhFwCBd9DFWgEGsHUQhOieMi3h62TNE5M59ibPaPYmAk5APCPtsq0Ky9gbb5Ayud
K8cnVMJHPqeLRhxjJl0VlWJtxdUJ7lrLqj0JLBazAXUlUt6TR04VmDywcOuIRdoL
EkmZANKPfF41w+yc/UMf402HKrwGWerxghsBBFEOXOpJuWm+IlsrOlc9XN6Vhtvo
ezPbviY2WHXIJTY+FOKAO9b4yrAiNiiCoD/1CSyxBabV/ghy65zHkSPyJe02lfMf
TpDEBXKsE4XLyBmIS/0J2RURR4jHsAVdCycIT+exR7+NO3gEj2edVZ+7BTYGMPE9
lXHPehfZ/XQ7r5SMNmaObaHAzXfqltXUyM0eSlCswLRDm2hsgc/71rTM3a0EP5mL
5BmHXOf1dWj6XjAnTOq9S06CeJU9xzUZcZzcvMwHXMq5OIBUkElciWZ+AA4i5n2l
7L2FT37wMuOmo7l2ySxuunmrb4sm1rhizelWFaRXVJfSdacGwlXzc1gyz1aDSvif
DNrtVfbBl8fGqZ5VEqBS/0tkRyNtOw2Z6ljQFo6SrsbeUtLVeLEIGqg7X7aTQPwb
yl1JG1d9ZQDXqUn9VbMcIufs8eO7VHwx7j9oRf7BXKVoGR+YOsqPGizxP5my35jp
FYEb6E+4BW3SO5dHZhrCNA==
`protect END_PROTECTED
