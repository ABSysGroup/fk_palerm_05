`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sWazIa8sVpkofcPSJKK9tghHtveYSX1umXqnB8b803PCmJFYiI6v1WJf7Ps7Beie
uwwSjf5gcBG6UVnZKbsNYMlR8SYaMd+Bw8wG9TMqIWGq6jsJ9ghZHwHarAbzpGVC
C/9iwseyb7BbGrApBQtaGc0NLdKmMhDPrMf8qWSHOA0rlFRCWtWTThN2tGBb49zX
bzdtzFhqsBTCuQCHtOQxtOMLuLW3kjdqIuqmv3e6Vpq22fmycXYeOLHJv/aDe7aN
B+xolGur/3xdW/CkgmAVNlhU1ClNR6UX+WAkeutUkUFlK6af2ecfhvVTuo/10HzB
h6Uen2FGMU8NLs/JqvsLIfc6A/N72WtJivLquKvKTLDC6WVw3TxX3QpIzzGBNe3O
iuIHGh2JpDk/iZ/hgm5+fW6DJtdJf5Ag0xFfsygHKhX++9B/QVMkuYcKapGzY+nD
6nA53/LAw9Srp20U1hP4wC7XpXLEU/HgnR+nlqo8HCiynAkWzXfCFyoGvjd+QPgO
FYLRTJfFq2q5amc/uXLBeEnlAGmvE0gownWeHt7l21/8c1fGWqZjy89+CN7uK+3d
mSaKGQEJgKsuyP8z8z8NoeVjtITkX7JSXQievaV3xjG8qmh4JdWmX8orRQOfakG4
PDVsC1l0i3APY6KD/2QNKNj7zkisfDrW+L/hspH1aQ2/OogNkflNVEYh+XewA1G9
CVxO9IBwenAhFPSrN8a+QfojB/PKMOSngXGO5gInUR9Dhl7FW72nmM+i9NE/5X5M
J3lDubiC2PCqOsXHM3U0ufSl9ZhCo6mj2ZmCkEaJSsoydnSsWDkDo1NkOeMMqG7O
xPgir9qZKommgZnV0YhKg6EMTY0s3j9+1s51njvFDOS1+F853q2jPc3GbEdUapah
r3s37/RGZAtRr45s2VeumHsibnOlX1rv8GQ+82DLH749G9ypuUfHBl9/Sr7tjNbk
Ar8V8Sa8ZwG0YtFWtjrv/qgqv35AP9AmU5fOfAgENP2hI4LMr1x7+wdxFhlus7Te
9Je2eHKj6/ilxnjdkXIYHrA/2BzwUkkz8UJYx2+kx3URz+A0XXNJqPpkX7AhEvzV
M5A0ebzplV3mQ3zv7YGjyMejDnTP7dG78KABUCdreTWrN0tc10++RarQECD6uyan
qNUFIPc69G5I0U0muTL3sFhxyGVITGscpHX8LwLP1foTEmapmf22qilf48fr0w/c
7uWjqaCL43G3hCoehR+YnNyGDgZw3zsQuhrolaA2A89saITIL1eyYpADIk0tJxLU
/70TDX0w7xaicRWKucQqBLIf7kytRqsi1A1sjmsFGxaymTeCqwjmtHiIUwck+s8X
2bwlslOfSxBkf95Rcf+oxyhwZ9V2yW15dRTOiYYEfGfY/yFEX2LaB8Sce9ntZuTK
dFUq+ni9fnmqouojSqsN+QM9IoF+MHcTY/+NXLaAQfaXyaWsj8ChhxCB01M58kGY
hO8KOu/QOAbxSe6MuyE+p5co9uUfszJ7C2giyhvFSl5tcUeA1FPfksvWIOjncHfj
L6/kYhDAj0qnHokwuCkaPGJJntumsLYlyzOrtN8L7ikqeMOiwfK9H2OAcEiF9fC+
OpmdcNhx4RexiTcwguDb2OiDsGj59ddt+dZ+db1FF7Z0IZry5V0Lv/SNqT9SPYb2
9frrhdbTB6HPF38xiH/1r8AK22yjcu8IULjGiKgIPKkw/A5zea68c2DWv3leL6en
wFmvJNMj10iEj3KdTlI7UTnDnEZGzWRsuOvBKs44/LOwQR84JwDyNiPyQNlzuoMC
JqSUBP1yv9RRTEz7gyI6yHWhkMObilz0+tJK+zmX89z3WyAvDMGgaPMubIzoTlML
uCYSE6/RcfXpUS/+Nz7qbKT2l2myAb546+oWB0SETCm7J7mKgbpcF1NyUTXpN6QA
PvjIP425WgcdZ6F9Qn0qHvRkuc/9IUw0NQraxKp50Ws09u0qFAIZKLOSldzrLKP0
ge/CiN0MsBCa2WQvIDKhush+SthiTLs48jlRjOLD52nntE0k4x1A7vl6AHtn6wdb
G+G+dOkLiYigSIb7vDirWzEFX1l96d7aF6mIBXvQr6ixBEfv7rMj9nM9UUqClew9
YfP+6gojJM6WjM2E0LgaPDxdO509SUqT6+RMdhakt659hJEZWQRFq/VT+oJgHabD
OnopgK1f9o3AKL8P3dfiweRD9ywVd73yfmcWL+i0dO3ElACqGeZfTbYGc0Y1foBK
Hxp2JG0cN3nP+KyvH09FK2YaIUEwJRcAXibA5LtQkTor6qXlUWTlT05sxyxR0+/A
/dEnQM98PfVNz8jztt1qPhk51m+xErvJ0RQ/uuuFT1e9kO+8YBFJPJqU8fcc9XUF
oxOy1d/H+0slWY1yCEwM+nsFjFGpU8E1ID3bPdLJFB+BY02i3MSVhMXxqxLB7IHO
VZ1o5NUFgwuCKr7zMUKjUMwmxJkGOd98zYnaD0DCC4VB+oSlQnL1h+anwNB/P+Zk
QqSVC1bbZcTx2tweQMhqceiyxVQ8kSA6eWuPSkgyL/HFICdxd/3V5VqFbEtzqu4y
LuUeNc5rjpHU51SD1L/yi83ih+4QrrLDfKTOUmeZJkWDkaj7t4WsMrvij7BtZj0Z
MtvvbY4fc2xa5LLvMjY18jYjCrS0X1BxOUwoVKzUQvZE/NUep/6fmlaJK7CrxeJw
gXTHAwzm6HO8Dh9bLVknNHczXtDVCcwQcpdePd999I/x75/10rf1i7Wv0VRGZMbg
v5XAffLoz+Zy/OnUW7LD/QI+Xxgo4/h1WzBWe5cmkGtI1a7pzkE5XNR/WjpLgGhd
cJBOPZ+OnXpUwZLI3iPWnfhT1QgglA0OduPaNvtFarEnkLsw3wDLa+++lBcdrptn
Mv26mH532lheZhbxYDBhFUYrOZg2ivlPYsLl4WwVHNwnUTLB1h+aVop+tNbZLDmr
iUp6CGwTJdqyB+IOaDi9y+Ni4zO8o+ovANtlzlLiJt0Gsu4l9KkJ1pmHgn/r1JBM
nnk8IHlfv9XzWIuAhrVp4BqT1h/CCQ+xAurfn6BU5REPJ2Ds1E3zdTOM/foyBrMD
yt3xIO+QdMOBvxMT0/G9xB15wQMVNyqqImr1TItPgLORAme1e68o0gEGKNDwh/Tu
RLUiitxm5RDpEkYYNsLKRWyaV1mkqL4Lkz+oteqzL/XzChJboxz3zexDfJCtBqzA
2ZotegQlw5zTB9fdDK7KLLB6gmb58y/eJ6D567I13uOKlJNdcJtfMc0Ty0eO3TsE
PaMbigeC4mKEZE0aNeLo+Mk/TTCpuaxQQ0TLA3pAStqE328PQdW1N7wmyeg+JC3N
h5m11Li/Pz5Mk8PS0acJjM+JI6mSMJhN6iJitDX1BA6MdDn3qWotXQldvAldt1dn
7oEw2jeIVz7/shi+Uwtv+erKj+i1YOjMTiGUo6eTiwPx0cSq5JvQkuG39rmFDvjm
u1iPv2zRgXHw3SBJCbr4Bgk4Liv2HeOZOn+Qjy5cY0voYqaVKV41+HLiNkr6MXk1
qE2NQbwJ3lDx1+bAj23AK7qrXhNuvNAYybaMxKyZI+9CTXgAju097r5DjkZoTYiY
D6jnKElDzdU0OLsLtaFhbzpBEy5jvAIM+qGOccI0WvqD3MR9OGWiiamthZLdl5zG
JuVjp7CoxZ4MXBJLNIRP72T9xavAW5rD9XC8Hy/1G0UAydQyA5KQavIClNaxd9Ft
z2ruKTclGrAQMFCDDRU7eBpbxEN4ToK2bpSg2XEfnRZa5BdlxBc8oBL4xWZ4xYwt
a3vaV+/gA8tPGXEhplCGE6G5KGVscem50vQdLlY5eI6YteAJF6CsECVzKXo8HXhk
/0nDHjBY6levSu5qi89gviym/47fYGvBGzZbeeIa08IT2xrPbw+bNB+CsewisAJi
xfgHN4a/Ws7dmhjT+LyNzxmXAcLLEGxaFFHaWCrtgk0Rhs2tnwAFEeKyoqdgSzaq
IBTLqqsfpFIHJXPFiRQW68uNtdLBO7SHJlzjkmXWc7+ormBN+BqUz1QDXd58PXMu
vumILt9UmXGiLT0UQVNTDQucwcaZIky/KCipacfigS9HAaP/9TvKcUWyTsMnx/bC
6U0R56/+VnfXQuN89B5L2gAQXHADNOzguEavZwhwby+lmKhASE7SAF/KaVNmJRtS
8B0o6SuZO0JhJfzz74DCU+D/73hBUIH5TjezIFn9CRH6LpUgWc5XvB2eExrrthas
gv3HzZ9gE/ug5sEPOUmEUaQ/Wa0BP8hNEJlP642FLmVf+dUtIdQZetz/el4ywxJl
jUhEXiW+2HUr6KKPNN0Kie3Qt7ABe1SB4DFjShle6+ILt3aNUn/JVB4n4xwmj9he
D/0Vzyepd1wQylN2YoiDG9gJgvJAQMiBymu6f/ZrF7W5l1fGp3yzitJa3Lq284eU
/rurl+YdMnQPcg+8m53Scq1T0Jx4u7vchldSEeVOd0njxYIO+0yqg9Ncj2okUQnD
p1zNUMLWuLJ3fhpQbq4xJkxnfvpMNKxuSRsiKKRqbDV250lxW99/E5gkTutgwBtY
Clg7AnUGjxM5+Ht4rWeqBSq/rnGT8aSs44QqD60tR5wOz0FnpWohxdL/5lcPGY+k
/zM1qtE0Bi62akeZ2jylqZtPkdEhDf0B388SUGWIl1m2iuMAjexDaNNBZuRDdKu0
eD1I65ZaCfHvAHjkOO5AK9MiRsDSW0cTStXVJShTtsHVrqZZ02m3YmGEgK00upsS
QeB07De45hAMgRbPJFGRIpCrvUMjLEQKNyKb0zg5yq8/nA3Yskgg/yYIlmPB3LBp
cTG72ghQesGQ9ILi4jtApDoBzEAqF3oxUjOHy+Ai/Pz0cxMOer6v39x09du0djc3
mzZTHwi3k1CAnK3/sY/EJkxJjBrIBeQKo4s39h6WxLeHQ5pZ+0Lj2yOOxRjEqGuQ
4+NffJPso5sglc74oAEPiU2x9pTKv7JVLBFI1jw9qaUnZ24v9OnZKRJsVQ4uFRpu
5I1Nkp/Wo5tSqWHpRXXnnXKDcEUBtnhE5LUk0I8V5NUrm4CG9zHY3fZnsY95/1M0
xGHRns8Wp+rkefSZ/ttxFNU6kYt9ZrKI4CT2C8RrP1AqCGt7Iin62ikcIkK3wHCl
Yk4Vwjobp9SpQDe6C4kPJczQKQG6PpPDN8/eE9/uBU3C6kzl3mOHqnwFVwKZmXZE
1lSId1VwrRA2slpObQFsS9Kzm+FuduBKLp9GlDGqgTgKfQ/skcsBEwNRRdHqp5FU
1HhcI9ntA9gy5MSOlHzIyMmDFR/BAPQdnRA+CdsYmAJF3Kgdrcc0ExPP1PgyjyMb
8Q+U25NjbG4olwMOxYlSckxWjxa22MBc2qbHkcbaiFtNRjXriBDqF43WTklNFdu/
0b7dV7Lp3VZi3cjaJq22MzThgpmptekfE7ZZ5CUXIluO632BYOu5QbTO97sxm1gc
6vWYFXIPXyq3baUM86mog6my4TifcBDxFuOnCFAW0Yy8bVG9Nz0sgbLvqnvnkhuB
yxsEouIxjNoJdofixWCrMNBldoiwN72wHHC8Bw/G+LYCBrhBnN9KwipohGPIbcbO
1uoH7Rw07+1Mv1QTsPHojJ3mLJvWdHz3zs/4PEMQqyaPGUFq6fQOAFpB4JVXNi8s
fPEJZbdFLLZZmZjWGO60Lr3sR2XhVLaXldzk4QTo5FokRRN9D2gQN6gBHyYfwwg3
8IYNyX25xMXo6UR0P+56H19EDQDxJtXXfvJPqMRRONbQmcRU0wIzwKOIhIA0z77s
nh0Poq1TiK8qZxdqPyE6G9ljWqRtcS76sZVxKDWJ/RYLyberPaMCaDK1P76aCeRe
AJhwURsMxsHag/5lOsVdNv39GS5QPUUl1G5plzoOCYJFQC+X4w15pTUR6CeEU7dN
Pi8DMp9ng/wPskigRKp1HCVL5LxtDlI1h1NMMz5iBpAP0uqJ/8UmMxBVFD4czLOb
StlaZYavODoPgOIRlWUCCf4e91iEAAT+YKM2/VYJPQxx+8YDj3Zza0vh8SwMn6CK
9sVZRzlVLk15P/KLGDmUrRUinjF6rjurbbcNOu8yesopdeg+3OPRYPvrQHGFA4t6
/3XnDgk0iJAlUQjAhvKOF2pbAvis8GgRHVz9pjvwU4Zvg1bhpX4aBTwdRbxUC7Ld
0Lg2thondBR56Frc/j52UHc7z45MgCp4P0l6FxwdZWrhtlvIdk6Pv5n1Gy3iRLjc
KiXgYkP0HcJsAmzYEPMkiBBfQkCGR01d+umwVztDVT140cqQ+bauAceEssLDLfvd
sdnXvHC9ZWiE0t6ZEF3+EWiSABiAjSL+FYY2XPhpMIKIp186+8VAAgUoUuqvo/tW
HKwNPvEWs+d0BqZvmAAvjEbdwcdSvB9NFKSRT9dMyEIj3jzkbJgwCAXX4MiHjxv8
H8xR1ucp4lyXNQedCR1vPUuYWbYrnmTt2cfPoTqnIkWU6MJqSCsRFLIgHWN+3cF2
xcBrGjnSWbyKU+cry5FOkVvCAfTfDFa868GpkWNbnaAaTEvSgg+5zPrJcv1Fu/A8
qYm47dpApg3xRDFO2ys05uROuHayX5XUjJr9Y22NJS0QutITpAzLlsaVx7Mwapc5
uOmPf1Ay24NCe90ZE22YOJpA6njyw4JTUDCZtverE/FZwTV2VmfeLwW6DlEAW5UU
OXTijR+acAM24PG404u7jM5WoQOe5q5qNmbzbX7T2SuexRSLALmO46qWB+4dao2x
SneE8Vi1eljq6W9ZeH4WGPkNeu3Uj0WrLAmluJK8SRO6LmIafWq+AU1hN5f7hRFp
dX3bHBQzwGMMRenGwU7mAZybxCS1MfJYp4ocYICCEPGgfO29rlJa2Gqx0lTJMlaQ
dXzb3VC6CDGWnj+B728pBoRY2yq0Q/7P2meERQBSOjeH3z5ILPI4dutiVzAI6B4U
LlEDzcZfZD5yAkE2+XcUYRa/zc4cSZp9dV7TTp2JowIPLZo/Y3NVogo1KYuJdVCu
06aA+rAPW+VLQajjx9NJWH+Tr6MHHRlKp8v/sLvxNqE3TYiRykixXjPch5ApE5QQ
oXZv+xonE0X/8Et6mIXbr9s3xHeMcpTeH+NsAb1wwHKH/h/1ooTfcYi985teRJ58
ICPyDIPBcmetpalyCDRHSZoVAXXzBLeu3VhJgz7JOKnd89wFThb8LM0AfKuo+qv/
MNbz6KXD11yQL3cLR8HdfXk3y/Njjua/Yy3vPj6ZXXvqUEK8X6dWPDh5ar0atjA1
A0CIePG+DBhXCPajCAm2FoK7XccaGNhKJ4G6gSAh0Ghhy279gis4PEzRb0vQdGws
h+eelzUTBcU7ngfdryR7niDUozLYoiKDACg0iQ34099DQUMtZzk4Q1anTma3lm0m
yLJTE2TQG+TdnCgVVNl2ZoXe+DarXAtVUvC129F/YiDpC06sbaCfDDORvIHtda4+
7lUGPxSpypNM4wwqVdXBI68YA+tASlBl+rrUDKq9A65ZCgPch+OJrap5p2keVN8I
4f2YRVM3eVU1pGQdt2ficmuUYPcFcNdLSOUifS4j2xnoHSjI+0b1q6rHr2ktfJD4
yew2ry9VlNxLon9mip3NXeJid2+TES018Qjcj9458+hY4y3v7kEI6iElAbmkY+qq
PS2hzG2/Z9KumoPAzkflA+tFw6Kjx4jqqf8wVuShEXvkYYTw0I1Pz4j5VDON7khq
ytedlKeCCooOktqi1WpHwsvsPe1nA2AqBxddWwdMQ41aQfQCpoBTuomndWSMS7R9
Xpw2PjmXr0ImbYO30bj0tOTIH/uWJr7TDsWJyvyc5T7BtqtTLC/Vx163oHD4TtxO
DMcBwmSGS6PIkIyM35ETEbR5ZBShKjrKuku3bRJqp1iTSAlT/I67t09QyaFA7Syn
Ulug8JVEeg9K05kVeHaD0ucGYAbVjFJgyB3I+HexB0hRl9LEmIVvcVpxNwxMt4OX
uXITILJ+AG9ocZCE/Wc3Eucf20qJVpAh541tmVoGDA6J3Pzz3s6h1CTf573eiLxj
yR/32VVaWayq8qhU4AsBRUKj2AB3c3WluNj1SN1giTzoPLM6OJCasYnu1AoVXx9W
ApczYO9/e6957Q2lCc1JCSgLre0JbL0Sc7qu4Oa0Kf55/tDUeDGuTyf80oMM6219
WbRkqawOSBMA81NyvOfir7MPFz84VitdWaGf8zJfxUjf+r5XLXe8zjvXaoqSteuO
DKE2RNzm2D8EaCXmsiz5b4pYauAYFBjpOtUrklyIlBJwA4wfFhzSRxt9lw40GhY0
A1DIna+337BLXfrufj/EraEKFrZR+D1el03n7FD2trFLPC3OuWDEhO45kFYkoeyN
B+vLiummCHgefFHxuHeTs+XcOVs1hwiHjlTvlT298OzAVLgLJp2Y/i64DCqgwik6
s3WpCYQpnZWJVxaMmnUYCszYDqqBpx533mwTdefMT/BIBdPJCFlVK9PcAjuWwz/n
NboRWMRi6zmSsdh6EcZaEnDGEOzuaH0Sw6s0T4t4XprhdXl+B7NVn6XXaYaesWm7
rTHtY+w+AHsgBANvVBetX3iX1GglMksayjc8oPDGf0swOeWfpifvbAO9tf3yqzE/
/tPN8Er7sMS5XYZnE7olDDZKxN0DnogRJfMmud8wGOuAKqUMEwvfIrEub/10+ExZ
9Uk+bmvs1MCPq9VVOUxgm6ONqudQXVHi95EbDQqZLAWHj3cGJfxSdrDxFZNQdO9g
tkq2+5vZ5Zq8jZcGfv5TXXfzagvDyPxw2GYa4EyOz+I0apXZOkvG3Bqa+Mw0yCXx
z1LLACrRQI8/equuM5jRU2JXsVeaEJmsmgQNe1AD5wCHq1h9GrPQ/A89q7Z5lf1a
BPNmuvk8DscoNCuqkGMO2L4DmBGJCegmRiB86KG64XmIhlW54vPUiR7Y9jk7IRXv
2/yDYh5qRF0mhUY0/LAexBP2s5gPBKNSNruOxhhw3IDIs2nBJ9a0Y5rZMMjBK6Ht
5VnwN1VCFqcqk0QqKiTntfTHASNwORCt1SwkLJPi36MAKTeAZNqGSMqrL3UaNRRT
hNlxFL2oMOBzeVCtNiyuGFmHGdyN84TXPzpbfEiMoQzwFDnpvJJfIPiJLJuga/qy
z9fQDqOd2SzPehoRwPCHAivEMgQyPjUVpKUGhLXbwKz65M32AP6goYDyIT7RCk5r
I3SRjkR+cpJjaE7Lms3QTG28a+y6Y0uckvCGYgEBWKBWtwdAe+d+2+m1UxpM8YFq
gWQtIOP7M+KczUT9xstezUfv+ljI3ExtZE0NZ7IuptGLuELOwbgqsnkEqIPtQKuG
QMZR64tRFacDbvLeNrD25s2b2Phqj+85R72olCPpW6Je5E82wocwfrvfFUsHeDFy
R/vgZUWMp5p95tMnaLbssdPN6DGp4Y0Cp2jZTi67oe6WZKVhOm+YeF395CruGp7u
3HY+L02pdIIE4L4s6fasItCxve/cOnh2Bp5acKfRztRdPhg5Ef4G0kxohYyApJtx
aXpeXGRZN793YdG2ifLYUDPbTWwXqGEhdGvETR2diPJqM0DRRXFa+CjZTWJkoMDY
FsCU3198FegnBuvlMLAo/xhqI8aPbm5TbgmcETIx1QCfQW75/Pt26vXRLw2Rto5y
O62PbKGYmO+qpEsxinxc0tuA3epk6C+NjS2g+U3kItzca62vTb5MIUYVgPN56xfB
1YbsDkZTeVqGJ6NOYJzYCt0khI3TTgMU0wyW+P/H9blO52njOb+8Qybk/WtOmPbs
SXmM2NUOLb119eUkFv3+XvR8ib8EXngwwLWJqIB008Qjc1XOqY3wbSNAivmsoIdy
cnRB0fsNTlk+LZg6Bywuyl2lszoGD1sOoOLFPmrhmUI8HHv1Iq6ndBv8VyvqAolQ
KzwuqcmVwKv9NP6tTve+U2VMYUCM13p/Na7s/rVH2JccQWx6pUGK4k9rKcWiivAL
R/bmJ16zjJbgUjnlvGbicp+uzf5EhjZqbQTleBVq49o2SQruR2yy/Kz7ON1d8Jx9
3A1eSXzLb/tZVZ2KvxImLq2up8Eem9z57/D/WPIN8aGeRhPcvQyOq+c9tHgARetP
KCBknb3or5Mq4Z8mrDe9bEQdYCKOxTPfVhPsabG+MvAXPsCfQFN7NjBGbEkjQFzq
L9lUA6MlhgY4XHfrDM8KgwYkuw7UeaL+5YAOQbINbwi3som8PQ4721zoo03V9ztn
Q3JYnMzRL5bSk/cYpqMbj1rD5ttJCZMIE8WwopEkutWJEHkihQBcw4IqT5WDpsjn
mcZsBwxbDuqtnZmp7d56gEihiYbCYIfG9LrUS8JU6sTMdgXUoxOwFHKA/dsjKN+P
m1TVzmdp0rJ3Axqv8WOs9wsyUKmoErCRA4SWrBqV3H14/p0H9vDVmz50uYfO/nGi
/ZkDdSJyM3o0sgxR2Df2n7EqO+5+IXCeHg3hEmcoP6tD2gEqzboAbWMh0blThEEs
35e5rBXZdrf0inYNy2z+/Vai0+4I1dzLAWFPwPO25tMqiHFArdcEr8HWZgIrHh0g
6jhagEu6M00zxHiHgCxHKvEA+nPRM/HVXB5S56B/fm2cObWnJJpQvM7cGtI/1DW+
lw8iqQcL/5c2bVyeN3GWd3J+u8QFjX/9Jwtbk8fJOhwZrbeAUx+uF5n1+7+kmYJS
u2Gcj2c7f5QXhCaizUMbpWiytt9C2RdKSgRxRntCEz9zixpMA1L8XABhJfQGNin/
PXeXJwJbj4NwErUyFkMYKQSOWX/8j0YhfMs1e40QyUYVDN9ugIid4AE2zLi+on2q
6S8dNOlBbboD19udMjWwg6S8sOgQ7UkTky4xRx3+mz1CkVvFLdQOHN9Cpbp+aD5R
+KKZnLBaQL9IhBb7p+asD2skG4iB3NdzAP57AE/HRv3Wp+MAOiMrWUk2t0EtkxQz
WPPSl1hlc6oj7JwYxRtwnTEHoFNxvoGJV3bl6TQ7mj9C/US7BF0lYUsSPMoVwwYO
3zgVP4J5nr5OC8HJYWexKe83R92BE16mF6bda9wu7YkuPIDfJ4z5CjSdPTwNFUQO
r6xwrykFr7KNS3iJVDJGKsWAsquGwChHLqlWjMYDmDYzNjC/vJ8ZJUfVvC5JRrnZ
ej0CQpCLbOEBO0rrLj8+iyclKRp3Jme6Y2NeXwCTEx0JCnUO9dChplST251+eM49
mD1IbtFrCOmmucsIuFjhLYQ5XMBoZAXXA4wQlMKHARWKqKgulLeAS8aKz+jsWOCz
hae1MNh0Q08kLgBhCtpJvCuMHwypkCuiyM+kmdFOyEzX3T9afNNCjtd62SWskpFD
N0DG5GXdodyUMd4dbxJVh9vQN13N1TVfaQdH4OAEDDWHEnmzC/eO0pw5N6YY5FNr
FY/jIzT3wdwrq8b3idn3fjF3snKTi14o5Velwho0qgil+ZanWrM7FoXqQaIzDnhY
M4ofFH7XaLlv17odTarABm9X2cgjbzkRso+FcCK9ep2jjMrFMFc/Ks9bvNDEPH3q
p3E8UPuALZGbdKPNdfy6IKVIFrH0T96LIGBA/UT0NLwIaR17MjXK1bQQ8wKLRKma
BmGNGcMYuH1wZTgDT8kZ5dKfkfypwtL6MCN/UyhxBBAli+5Kcp5fnvqrt0Un4JG3
uNRHvJ74PBtvrVnlKqZTUvpsU/J+MOgS0E2EMeiLiMg2TfKXJnQP65EH/BwK68qx
m+sdaQ2/BROIrBoMiPQDO9M8VM53oDOogr+wdA6Ux9Gz/TAElI/y3N7wbL6kViQc
4nNn8Gct3ohp9KU5WTuHySY1xqKXT5STvSKcEcN8t2madldZcep6Ewvn7KBSVBnv
udG3KZbR4btcyC8XZwrmGl4vhcOCHj8Rg9NsusRF+Zr5znF2AgNzD/yzOg3MzOlW
rfgp/YY5jaxIRSDwdwc3EZD3DjSFSbSWFN9SGVaoRNgO0TTIzes78NoILj4q5+Z8
IANKMqHNdzYs8c65uuaVPcxgWj45RkYDv6fIDcwVYg4SIek9nZZ0pK4uH6cYrSVu
58jgcL7NKK2H7DW680qB0TRMkuVq3iJvaNQp4nrDQXFn2irBLXDkpRbiNqXEoX9x
WTMlENeT3X2U0JF2MGo/B1TahQq7TFp+5n62D5uVuLb7uCvmdIdBW9q13vfD3rBQ
iDqKksyp0/XmFi4Vh4G2DU+yWdD9kILJ3c8gyauCHFM=
`protect END_PROTECTED
