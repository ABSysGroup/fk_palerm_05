`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jMxPrimBklu1om8qTnQufb+CDZkM21c7xob7vk3/P9fw67L5eoBqiulDKmvSBbB7
r9B5H2YXw0l1r5iHZ5OHOEE9H/jWYh/Y83TtUVQr7HXpq0hY5BL2tOj1Vu9oRzMQ
dpHJo/ZvEq9laxOE0kgrvdoDCovo0A0OtGJIgbd2aEYkwvpd1a4Vntnl70NUZd/0
G6XR2AmxtLKPwSrca9l1aF8N9JOYvzyXQvHDXpoNec/nnEwbp1VL7CPRMuS0em71
83cOzsoX0h/JdHmkNwl036eVpOdHc8zlKhv2h3iKI9/qT8qnJ7HBZ8f6zPqgiNyW
ZtxJKdn70RlY+WdhLsQiFJx05teyeWpzTfyXhWexVJyLTxq8AGnJzKoPsQmhFDuv
/zHxWiIZngaGvj6vr7bEM2U1KKkyHTDsg8SGszMxaDksbIzTvwyefuoNyEhTQVZw
Is+qLQyH9macfre6FvlnexHxPPL5/0JJYbQ2uhUEqco3Flgpf22YiezPS2nOSwXc
Km7N2u0ZRCPanG2WZuhclgV2p8NhuSc/yVWHrQrpk2qP2Xej98oZ3G6O0Rdq7pDo
Ek0PO2s7Y+w7rKN6LRlu1zfnkuCX1DDfE04IxyabcRkhCn6/HnJGCEJGNqDnEIxt
MGLebwJ4oAV8v4ioEaEAUwoyPvazuIgt5CAnpNf8rURcWv7/AVEDK439G3cJD2/T
g8LyAEnVFbYJIcPzE14d+kqgrJD/1V67kabj0eprrav+hMnopDhSYjYxeTHibo1G
KTDCHnhknXOiXUZGFRTD1/244xDXB8+nKS6e9rlEUsvSENWH+9d0LBZB/i2Ei9OQ
Aj4sJ7v+6+4UrlCX1+jPFkz8Woxq0KnNmjbufBNcxXEZjd+lUTttwOEWYxpGSc1D
EaHaQZYfBHgGi1HQVSXmbg==
`protect END_PROTECTED
