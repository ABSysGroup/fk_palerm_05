`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wm1xBfRVeiQUPgqKAFKOfK5SFBo0rtb5S4XRWtX+7fqIJxW0M3P6GqHMePjZuvfQ
CR1x96ryq+stD7uhzJ2+S9sPgx9TGNlOLNc3fc30PTLoMwHDqMG2DanBi9OBwVOE
X+p5h050uMMya99CmfDk0Blbp6EIpaS87vaiDt3XpFxvzfi2xRxc6RJzez4eMTC/
GMcW2NvApu+1hDEhLJnU6aUbOYdUlZYxYyEwm2l6XrdszC9FAONVAtT8snuCDTMq
zSpqQQzg0RxluBslOWJBH9ioP3WhZ9LNiRou3FnO4lIPM3xvA4aVG2jdZeqy1GHC
nLMJdEp39RgYZnnuVSd6fenlrGHTzC4NV0yXX9hNr4xpn++dwfP7lQpKYt4eespM
+p1vC0IFS0+tW2HjpzJ4/LpMEadDl4yQxXtPIXpbTNDYyLI8flYJAG3ASLhQ7BlT
ZwZY9zHpHWnjvB8J4PXFFvwX9lD8P9JFWq8aI7htL7YMMM0mHdCsD0J9eD/SrYt6
WmANXHcxd89x6CPf/tIOBxv7/xLYCsZRclpMrzcSn6IhHthhgaopCTfpSTyQGYSo
0zL4jnF9R5fR+tByddqhk7nOvMQk57/BUtkj5Tgmwsr/bQK5GkXcscB+xVxhEQXD
b/uNbJLpgxiqZ0bjFjgR3weM2BJXgUNm0mW9rBGYRe1CN2+2hzaXdHa4gffJsMYk
cuisWGb2oeONkmuGpocInfOkM+596SS549yjcVC8lfbJNTib0Gw8ZNqP/Qx5vPo6
ll0Z99vdg8VIEjeJccEUAEwOd0fGvOjnK2wf9ikzq7kNtv8TOhWW6rpNYDHtfKxV
Yrsdx+us4Z6zrU3s7R99qzdYCh/RFlfYduNHDVZAfmYRnAlqZOaEd4OciT4Vq57v
iWbM9yi5/myPohNg0sqW2KSbtCgfwo/NebLtEhJfMdTbN+wao/puevI/GUe1RRxG
a5pC5LxUX6z029DsKN/LNuVtRrZjCEAitJAuxWfwO0t5C/1sU6Imbobl+bbCttTA
U3Qi8TXAirjuo0ej4mPjo622hJZw9vc3hQ0RGc7xmenDvRzb8C1c74od1bomgLzb
Kw6uCKrECSRTYIXEjvFoh6RHdW+wRansTlxu88Pv2sNDmvSwIr+fUhtWV4XP0tSQ
lR6hOQ0IDgEh6i5L8wXjgynVk/TzZt5snNcxLrG6p6NM2AIOs1PjsUAXOX313eJp
atz/Ob+vo4tDzcZYcb/5NkVLIjvefEiDx3+VIqwBURUMmnoZKr1/VlQmB7WJMwfg
ywQ4i6xMaaIHACqBukFMM3paSCgtBY9JDWhZWlmLgHNF0mog61IWATzmJmar7Xpe
Ei7cz9VPWenB551KdoS2wx9/wjXz3s04uH3nI2OCxiOOw3X01JA9Y5CTfhWq1dcl
GtqFpkC88/c6vxBkvkFfb+7V5EXMCP5CkrW8fKe06bbhdQ4QnvAPwrSjVgDxyVmU
CJfQIuSq8G0FinVvjD+ZqK0XKF6qT7rPgXpn+WTR3xq9ojj8P+uGcKXJMT3LAfj+
1k5gL5g7vAHd+YMUqPMb6+5psWT5YMKwIq6WE0kGQjhQcVzHmuIsDYu4bkRHQQ6Z
VKvGWQXf9VmOPxwsasOE1HOQVBTm5d4Ypb4lY8FwZHw/yBjNI6TVN6AjtmNQlkI7
c+0o/hKQsmkX/Naxxk0HHGJVV1Ijh6YEYCEvojMtFEKa7q7ObznzUNXoJuekjkGM
u9KQuCzVsERgcqvketgbE5w20CyTBHXjQEve+knFLcH/KLev5FTySLoU2OS4VACY
EJYW60sgmz/KZUSvBPDFVdXzXMhngt+RmVT1YLBXHNtlhfrYJwiIcobllhTgIEsm
ZJiOzPPfDex1gHKGa4cuN4fsjY3bi+04LMQW7WIMhP5dvlQBmp9PnLsEkqjKLPYP
Q+Y8C5855voQbQEDi00anMl92lokSXVwEubCyDf5zjSoccbBdoJW8JeE23nwBfSU
xCHmPoNJnfN4DdOtPEGOb+vxhuRzIwLdqvpBmmY8C2bzXt4xVrK8MsaBEypx8pIP
pI7ayMlXu9XauSN0kQpZLYYqdluWuGCnvKgfElEJa9CBL+Dz5Dhbk2pMOX34G12a
VCsDnHZ9rQMLqfrgdbhqEpNc9rc68idMdUhaf1v7fRvk1eTxir3MkonkRhWrlo4m
sCIFHuYpBHrENFE0P48r5Y/SqfQuWwFw9KotHezoZjX2RPo+LHiAMc/aVVQuMw4i
7VRA7jghRyifRV8fYRPi9KVlgSa5Sm2AOD+CDjfesDXFyeEdNJgUXdVlcEQfWvVb
Kl8y6yhxXjzPs3kUt1skhox7EL5wlj0I3Me4NxT+MQA=
`protect END_PROTECTED
