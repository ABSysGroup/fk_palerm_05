`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eW0a9EQJnDDlCTBVFbxRQGJXvWA273HgGxyzJ42I1uYmvz1Pv8ZZJ8AbNiEGIkN/
mQVELw3C+nLSkAdtkyqnLMy/mhXgPjFr20t3QmorVqFaqQbXAB3ZX4ZFvhQVFo3S
GidgIJDjMY4BLiqiH7rLREUnYYPX8ApZh22V5Jtryhfh9iNXK2c/AX4vJ6JAj3Jb
DK3U1RaXoj7W4pUcphcrdU5Sy/QJCwCJPTdHw9pOFUBPIHRMfaXUgttXn+wYH2ZA
`protect END_PROTECTED
