`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Og0vAZz+DXSqEPxHFHWGPzn+bC1OXQjwIxbf0w6DQUT8xJVRTQ8iMAvm+rBY0ppo
top7psxENj253vniudW3lAVwGv9hZSJceTlnHq+qsG/ATDvfu3EiyWxpHPaRkBcy
dDKqML2X7xvNDSo4HitKpMMuLWEBGoIuNo5wFd/eSBovzpwLJOpY4QyKsHB293hD
uRWM6pB8AM6Os5R/SHGB7Ohsr/PiQk+evtAEr6PnNVgVqiLPQCxJNmSWD3a1wP/u
X4L2oRxB/vTSWnCI90XWYx8T4gK0WZN8EdgIt2W/m/NRfh/sN3B/6awkYkFPpchb
RnVDjdVKBT1KM5EWwo/iXLPlh+R6tlSZG2Wq+xmHPO61LDP2gQtLtid+oyl6y2nN
OsJX6PjYkaR0iGg9o6seT3b/sE5OwTm0O5cEcn+xGAuPoxh7vad6YVz69L31Jl9H
ebDdrqkNQyaVbXG/9PmNXNQ7n+8HVFhsPMYOrlhhFlM=
`protect END_PROTECTED
