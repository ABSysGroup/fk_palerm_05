`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EisL94ExCCwaRpE9Y1xVz6N+1wjrgVWMyowDdrnBgnJhQHjVaG52FeAL0meR8Fw+
lr3OKzoAwUoTI/cLVwEUoZWcLT4J9uChnoz1E0GS2c5BgwHyqqGaN6IxtHaPhN3S
zvtOA0CNt+C1agLRvvT2rsYOhEdQb7TfCSgKxsO2jM6CX+TsDKc5VEnGRfvW3P+7
0pfLm1kRw26erNJT0oYjIzq2xPexTv1K3BWioi3LM6t8XC/GFTdBLMeEAxEVgS/H
FF97CvZFxayKHtAykjSQeVN353ssoROj4MQ7e4otLn831qziNfovGHd8g0pVYhfv
PLbbEA2SIg0EPx9n+Ekp5w==
`protect END_PROTECTED
