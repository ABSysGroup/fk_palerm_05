`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hRyqZfFusw60vz5BTjLBoNv4bmpGbwrzlFX+HrpCINsWRgVWil6fT1IZSnQ++JMB
Mbpw86Aq+/+VUeiq7ImBGz9a3mKJao7In/zf+OjW+ESVORZC4ijBdeEaj6l8j8/n
qIk9/xa1HZH/+XgdDaaAUakiwjmUNcYNZ9oyPlMHZ3djZZ/nUMqLe777p7jnRf7w
hhb0D0Ac6MrWRSHEc/O9DfPOXHxh7hb+hO7kphI6PvdKdQV4Y3+8sbQ3tTWa8VUy
6E72JObduBrfon4r8pnLNRqAHcA1HAoz6Cz8Ecuj/LWzNAosPgO0S1Rcf34xB8P+
uU80nzZ+ZOT2UfjWIB2mXli1Bnc6TlgBaW2nRTFfgVCFJDQf2dsNWu4ikYp/cqu5
2KSNHeuXBZ+4WAAv/2pegKmOozV79b7MMy0eWfmmOe6VrStER8V3QONCC12tXoof
`protect END_PROTECTED
