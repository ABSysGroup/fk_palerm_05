`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3toSbzNk0pyS03G+g5RDqpZTs0Z4j9WZtFzKNLAb+zsWqJ2RmZq+qdH6KOE08TNI
XTKFC17w5swY3X9duOqgRHp1WHpa9WMUEOYeSNPuTUsFKSiker4XRuey0YUQPwcq
gPz4T89KyK72vlhiGELjNlCz22WlAoJLmMGLW3rliFZ30iHwZFTrUcVr5TLQR3Cr
Y6OJewiC1BwZUW3o/cl7lqXM+QCF/+kp5vsxb0L0RORnnw+S7rh0xE8OUY5Y+Xyt
TuqvFj/7PS75ulu0PEgPk7dGHfCq9/X+UGvzFoGI72pAX4pYjSVo6ii0z44QE1n/
AxJX5fDXdpLX7W18LHuGcMKfZIEH/Si+TmFYhflqwPqX/3kT9uNVSqCuIkvaiGXh
`protect END_PROTECTED
