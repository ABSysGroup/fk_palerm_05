`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
20dtM9n2rjBJy4rEd+lydP0B9ay1U68De7HosA7+Ks4kvQFWHAOQ5geDHadIC/9l
fg8u53FtENuE2S4eRi82l24T0qLqgnImGunxAuYcxzVwxVYYGqHALCT7kT7FIPQn
UUeFstLIiKiuuRFWl2wNvk5ZcHmtONQ1ajVQMW9K8zwwFlo16T5K8U6FDU7Hwa8N
w8f1HRpHZYHWonNotRFTTOnEPNiZYXiSB22hgmTSlE2GtMOU9TwsKqpxYdKNFyvA
6zlMRyp2QB6A8bal/su2ERa9KrdADbpalT4wlAuR5s6FUDKcnVaphTUFr5vxJWu6
tJ3fEgIgmUlUbV4lRf/rSPDOTHG92C2tXWwmXS3M5CcnlSdEsrDuZJgTdDjVXdF1
p92QPhG9Wag28U6Xfd0oboMGpRjJBkYgfXJJftKLQoNJ9hzpUyjxlMA6OwwmMdFT
9w/gKC11l9//Kp/qbUUaw8GuhSWG/S92nc3bxgpTZS3hG/Sak8Mce/wdZFp+M5hx
RdLSnDQLrVSVXXtEWlVaZL9wpe/KpOVTL3D0xu6dIId2pVJsqokawyuSDEJ0iE7O
5HMW6jGtE9EutjALWs43MKKxJFUE+6TtsuABDnowxu9HSOailb9J1SbNWqAljXrm
rveNxkRx92tG/lVVWeoOdT+9bpLXp7WtCO3XGMtjvqeqGWJfKy5VWk/0CzKDRnHf
aWPFtGJyEVzoL4Ta1+XilxrVyylatspPPIHmmrPxAjtS7y/DYODNVZxDhtg46RPT
5K/ovdsAQAmiHhjsRGrpzChIUbW2mJMneTDYDosLTilyrGXc+gn2u+cxR7CCv2U5
ZHaiSczXs39YjTu1ZKAKR5car6DVVGxYndXyRM4F0wVsb+KDuth6b8Wp/S0BAT+3
KsaxLfY3BR7cUbXCksaO8yZI8SnpdtdLOvcxMXIAYQc4KymTVSAmiMnpf9/9cFAH
plrWzd/XnVY+fD7IqOpixpitP3ZBucEQ8ehoGhGkp57V7liO4QKOsAD8375pIqNo
Wm3B70m4nlx334TZwQXA74G1sNqs+YuLd4yiyOaNAskH5rjSdod0wcyx/CApJixg
xlYTovfx/DkocnEXMqrWEiO9iwL5B6d76sLWSRZXVZGuF7mZB3gptqcYJT6mOZ/V
0Uwjf0kkTu9n7+KuNiaf+JJQnbO9cTxWgiIelpMr7WNwfvwjF0vfuRf9QsiKgkYr
b9HF6YU23OangghWnlu50+K1PHd/MpL5493KlWD4zxgKQ8JrjtZdr8HX0IAc9wRI
KqZcKyR5aYcqyWoAJutDX9z3PywR9cJEDzOd04NxlZ6U5kK8VduHIba3JSCPwjSX
pOyoOTMm7IxtnqowYgvRtOm0i3raePxs7hHdYLUhGpQ2OiK7Cz8BgguoeN+Sw+9f
8Q/6OsgRByvwuZ4Z8Zkvh6AB9iCEUzxXsuvBO3QAofpOf5taHfYOiLYy3UGaAnur
P8yA6ZUOa2NUfYGChHKdhLaxoaiAS5J0xA+5in3RolzhsJRQwy/BXX+Du4jvnmWM
4jU3dCY+soLwKEcXeRk8clb3hcF7pnfApFhqHlh0iaJQ0h9UNwVkvOWQSSgZ0F+u
BWDZxLzZ9PT91O12lYM5lISJbOhgFpHXbydHaXfWhVIlWobmrjw9UzAq5xBqldYT
GIdSHKyyPL45qkaMwsIWWEF+XQaXDaaqw0P11SJqKo260zxKSgLl9iRr3i+7Ezh9
nI9YKuHDrExnYpXCcFfjsj2q2w79FZUxjwb/4Ik9FfZOXfPe8E0WX86NfaUn3BpL
+35AYBSGIatNwG4r/aB4tZ9WtcNYPVnZ6NWihyuhj+o/E+dGLVkk0y8QhSWtyp94
jsvuyGmQYuasKV/x0/iB/wHBSn6KTSUSfCllLrdM91QTkfiQCTjb5zuh4M5BFAZR
WlFUaB1j5DdoPVnpetB93x2Tkibu98zF9/HG8HO0OPJqYGk4WPzHEaQ8q9WRZYa5
zp/erCS+oeON/h1PhpuW8DIVcPwkDvt+5klcccZ+obsRCBdCIOvfZpPXzNTg1CFU
1+OxvehgXWueSspSdeLLP3euTKZxm0Xo12Jh36mVqS79sfxZOwgo/jSYL6Rgb84U
PeeqVA/Z1L+q3wiQiu+HcxSopB7oPFsWL4Pu/d1EFZmELN5Q6mxwLP+0d/p30Xx6
Dn7KhZjQzjPHnWPtjBfYDdyDGZABIvSBLQVmwbxjSTGiGPD7xaX7rsuB7YJujXWf
4XwmqHYu6rROaFMJNvV41Fcg9KyJG0A3oxnGm/mjeir7ye5sAOK3j3R12LLd0CC5
SBFyiMlQcHyNFhqq50gNBeqmP6aU75k1iWwunk7HmyfOpH+e6O4BZPvghTImpTJX
OhVL9IkanNEH1osHCSVgE8kDHTTRlRoYGJLqVwmmKTRNyKTy+9UV+Rs1L+Tl4aRF
lGHGdHsw3bS3WnBGQrgh6v+vqihhdeABE41pe57yNzyknd4Iu+FMd67hB/X94q7C
AoWSXh+QMyMnj3wOr3vw0/VydqDT3cBbryRKJ9TcQnSyLap7P3ppZDIcMWoHpNra
e/Xm1j58p6YIlXsx8xzNXGDEKqB7hvheu+xDHRjG7rV1aGsQNXf0I/OHKNmNJcAn
MgETv67Eh3woJ+tRuQBjga54XW90vYVeKHbdJ9IoNnuDCjPs1HMYKjyvuEDZc8F0
0aoFhhzV+Q5oU2JFsBqawE3mbVxYLPqU9iPyOy5uc15KwodYySqukfe4PKLZb8Dl
tn2aGOcCjVs18DgCHJXS2y5ygCAEWlZLQ00foHcqs3ORcI3CQXAAPPHQycWn2CSv
UEuEdLC9+aOmQajl8KfX05RifLtWNtp/sYcEcgFG1AyaGABUPch8UlggHXUJqSEm
0hLFL6Wyidti/kwgYmNbTmZyOJ7jBQ9pccUiuIvjiM67oOiTJyX/g1pZM5pjwQUl
aeKEzmbrIk6EIsooRcppB+mXP7on8zAKR6xHFMgJeQ2FmLWWabh4mNRZePIZRfCf
sheCdI7HOh6mZ5Hpvmf6KCGh08N4gAxPQEhiicz9b/moqRjvyOtDzFvMThln1zHp
xZ/XiRtsq/TbN6gC9rgjmo9mLeJpgIOPBbqa1EUbSP9z/N/2RBDaZyQy3oRCWQPm
O5CpMI/2mM8S9FhLdeKRBoEql077FHBFDa+JujB5AnwH9pjM1r6zKdWqnlvjSC/F
tCbcRjh+waLRGRLLBwIGpqiNpmKhDiFozoEG6hQr2iWYNDtZSwtnt9f/LhDZ03aD
a6W8YGK5XEfY67RMCtT7aCVKta+kRIHXYRTkgwA/NBVZZDEK84Hyxw0lZiQpQz5l
2Reox0Icsw6AlyHMu0BAk8HRJHAZsNwDkl+0CQNOADjHRqifZ+6ry7yuADg6Mf9X
HHofco3TMrG+jIJVuZbQ+Hxe3xEBW9+s3DqpUhUtaJVZgJnCeifUd9WGVCX4vvYp
OUiwrkAnsUob1cXR31KG/mnrpM+nCyIPKqjYCtSL8uesOmJcv42b9cuZ5o5+vKIL
XlvTGsjEOQL1ws0FaT2tXub1y/lcf6Aqrpw6NhoMqWUpYYgo/iFUL9JebO7KyGmu
S6rD3OEK0xfeKzCiiPZhNoAIE4lvgRZGrQdvoQxYk3tglntlZE6qmJYJHhbaXCmG
pINepeOnL8HncCCGybaMCUtSEToYGk6iDwjDFXqgTqNBR71VqWNYgZMnQqoYC5HP
IlHyxgOGqxT3ZfWcUySIXA7mvA0gci2ZHELGIvaMtdRAWi2EhnJNgEl9pNaV77HM
3ZlPh4DsLSB7Hf0mnRr6RCssgjpR/HQvyp778FhPtMqjRx1Rn+I8HvwIWjFYgfBb
28dkEw5ypR/uohiKCR/FNE+BDPU6aX91OWuttZ1TMDgF24DuHEqSgz9l4r0XN1hG
uM04oms6pihbKssl8m4wuTrvW9QzqezqN9aR9zQuTZk6QM3sOXSMBKhmD8at2m3p
fPA4460Uh35OOqBBu7oGgSRGutabadOnaFJH5COmhEn6XlobSxr9HnrbXKd+jAvx
RBV0X2at285e/tL2f3qY5IOVEWjvINw5lw8qVMy18/hkvEqDYBNLb3mQl+vjM5Ws
`protect END_PROTECTED
