`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hh0Hj82AkVj7Yf6pTaYT8Pey5AhJZbuebYNIcuq7aeqwXzn+voC+cdoUFwcRV/Tr
ogPkC1oWFNxoBTpy8em91H7Ho3P2WCFnilalfaZNgNVQat8n+Rwz+b1AzesQHyI7
SysQDfqMZwQIUcRRcA3ejV7F5VicLz/OGV45q/Fp6Y9Hno7wIpBPUbiMJxC11GVI
2KUuTGVzAhDeqDuh+/K6PTP6IvkN46G+hbIhEsTsSbyusuHO0PWI7TcqjJXmAqAt
3vsaIhAoYeFCt4QpTp2UsqnTb77LPvWllxjs3RtZbWdpQLlCP0b86m49TdFaFAsl
zxt8qzco71ejfEOr2ZNuYh+13LfXxrMDsAtFb986MnRqLHW6LNkDtY6DAfo1SH5d
zOPJHSPag7+ob2R3iPQQ30QljpmbcbE420UDbnarIgLY/DBL9Td2JgfMS5UjT6Pn
1178SGnRGr2IX9tIP42kBjwR8xgMLuEgOS93Dg57/n9s4GgR5VQ5ZQgmD9hwzv8q
vCve44GjoLE+pvhq/ev8C1+MApp3RMUw7IiU1DLigRzbPSY2JBma5cdiEA7xuSRa
MVuWUPMxpEYyn+i3RLR7jbx3guTgPmcxi6vXv6rjDxHEvULS+Tw1WdpsVLSeTO6b
Ioiyjw+Y/dvqM+yFGbuh1pTltTf4f5EDShxIrZ/c7Tov92sAQiPmw3X+3pMyADvV
cEQ5wwgrYgnd3j0cR8b23xZvnt8NBcmlWW/XBglQ89B7XmfRewJhObafKyR7gHUU
yAX0u8p1K49AnhmymH1HICuAHmRThDAMaxKUcdPa7xXCxCz3N9zxsuEyp1b0xA9k
pblBrGTj7fo7d5OFWFETG8H8b8hbJODtmGq5w7q2DQdk4u0QgxViitj2BdUWEr7A
BRrBKA+8dYslkk3KuYCPdHsmocW9p9RQjIVVoRrz5ZXcds7ua2xaL5Qtiayk5luq
4MGsTg0m4alu3CNI2ygqDpIh1vleYGoIIW5hnCPJSFasHkkVfMn+vOJ0YglclfGc
RVSY5K1gj/tCV5VEj3GWUOkwNKncEPrDeiFGPhuKDjBgkfSZlws0l+NLtB9wwJ/H
0ZWiqy6zPKZAbPjj1dvx7vD/dSgvW+crpdueYC/E8S6Q4k8Ph6ddvMKHsoRMSFQI
aLQNfin4UWCz1uVcNgxcjN6yV8r/+kOEo/kQsu415BLpjQdI7O3dhkOvVbZ1ASBf
Vcc7RHouqau5pWoKURuIqTAdxYbPxAGUAcOCXV0FhcJExsw6su7zzWq3/tvmK3ZQ
fKrlQpB1hCiWNdrbaZ+XB/CFrASwFeG9d3ba1pCwiE+EnhjlnbVtlgoppwMYNufN
0ymWGb2KWGhz268U89BR8e7hd1RHdYM4w8GlrEEzmc/yjJ3zvZYP+N/Qg/UQNWdw
UwWFd+Owyjfx8FEEoPr73mwi2CLmGf9wnBh0EuDaV8cEvw9WOhQNifyMOufmzgGX
6M13Trc2xZ5JF5t4VtMuUBMHdcJ+LOVMbUKXWUeWaZJicQMevjKslkMUAMP8ImGD
XGYLFTIiuiIZHrB82reFFguuHPGy2gNZLnAq1JURnW5oabZq1wZjf/K8Ju1JsaCK
fx0YQSctZ4a6FW3k/dulhnkZzmCqoMKGEDoGvuEetWg6IPJ/y5ZGkNXtS2H7Wqa4
CkVUsQaNOXwtsi3lVyvlXGwhwDX3T58msfn6jVng3bK8naO0UsoclPoIAikKgYLj
I5lB5v5FHzyd+ZFfz0tDQkkJwyX86Cv3DzaL+beLy2MSJLMYahDiIv3U6+7rx3gZ
8w0KVZqKcedtOQlcYSRdBEtiZ21nGK0XC5Dzfh2ZiJpGlHNecnyXuPd3q1jr6t5H
DyLb792WDOjF5YFTl+KizK/jJMoSbIibzHYIjCXN371mMb+7BZVSgwWYeuShaWCk
zUfmhMrDTM2ELRguXuJeQXGkJFXaAycHoFfpWCJ8N1dZQdm/OfS7b+LA6cZ5QNiK
57/uYtZX+ujv1PtqkBHU1innkWcXokQQh7iKULqMbNAGMceyudHkObsTfQDdKp+z
Iu8enPXxbWxaEbm+tisj4dOO6CKspqc56PGS05tip4roRCeuaxruauBwchAZxSZb
DFwI/BFQ34NeVg4QidSxqN76iQD6kxBJTead3zcJqiMeZyI3/LGo1KQ9Oikxku+R
suRlKHFYJdwRnGDWxp733gh3qQDXlHY/lo+xPQc8iQSP+GfhR9zW62domHNsoyho
D7/ZjmWvrwRPJoZhUjQh3/6tHPHpGoUqHfz7v6AkukuihyOhpNlZOsx6iLyt03J9
IWVpPGkfOf5cemSgNMU0wWzzSgS34xeiQuFFLY/9sHrRUc7lSEa+d6m8SOVeP3CH
A4Rormf+/UogpUKbELEHXtxB5qtfGL+QIla2Fgg5yQti0IsLmo4JOU+TnPy8vidH
LX9+WkefN8ON4TOFmOWmge8S4lhBc7aGCebLeAi4jP5YXoXDBKCnkmMVMqh9AlWj
T0KfAR0rNQ8UYILpoChWVHXjAN4f8YRhu3ci0lsuBM06ro20uX19J2VgTvHWUKSW
dYN16IE/LeuDeYzjG7e1dV4NXCuPzEfQyDLFCwtclgKJN0eIUTJIhtALmjNrFRBm
v2xp+uuHMWdfWO1yPg2jq+yeOLCNQ8V/7hToXAwQVUf3+BLkqrum2RGGx5r5Rbq0
Q9450vyvEnVXh3RWgUjDMsKMjcBtg18STwXQKgRGdGlqjv+zE3uEIu/j7pu7pnZB
Sip1XW5ls1Zxtl46P28/YsytAi/YHU3Av9Amw7tqg097YS1TVfCp6s/OcOCsPC0P
tuM7iN9iE47YvQvcHuQsrTXV3h5fEmZHAfE0YpJ4BTvP1S22RLFRkzwsDtAp71Gd
87w7Gkc5QBnk0iUY96xeujA7ZhVEWKy+YgJ9i3/akLMU99KoeMWNCKFpj6J5OLsC
WS/cFygK20VjzAfyZ5ehNRFc+AovFV4tks+wke5lmDAU9N/sclIGEmXaMDYfEC4C
lGZWwkZc76AVSRWsidiNR6bJBBvSBq7yDiQ8D1T89/O39cTFTWu6PIjtKc1iM1PQ
2JWg71cjW0ewgkk0o7ymeSkCT//9t7ApzuwfMHOtf211Bc1dU03mMHVOnI5GXfdN
KRRPU2CMfg1O8o+Vsqy1WDxP1wDoKV05E/K/yt3/MIsnxgVVp2wITzT1kPJ9zmfP
NJcFQEVlRClX8SWh13NKPk6jbfTerhA7VLu2m0K+YnYDdR3tKuNLBctdXxfjRUzZ
tV7+KA/kgkBHccyZUMCuHg==
`protect END_PROTECTED
