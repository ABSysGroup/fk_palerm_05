`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YjFp7jkDAEvjcJU99Ex47V0ACqFfBwreUQ/mCy3mXLhBN6ppIpT+LhD/RYPiLnw1
0/BN4RfM7DcDu71SC1iNosmlPNMcXZ4rgTWUn31a9KP3EW1CBxp8nnmQ3pJjkrOH
WoyLJtQgnjbfu7pknZoB2gMUa7pzkXg/2snupcfnA1eCGcvZIy6TD4Y5DAqf3NXk
3zXIs0GqAkF5U4psAOkP/IApq48Z3Zv9FSruSyGr0iev+L9LDgqoUGJpMk+HKWyV
UpHnUqCb60uMLMjUDj7LJM+fRbypcXBgUYVH9X/mvAsJbSjpwwO+VykWLWwHfj10
+2+s7/40P03Jt7HI159A/A==
`protect END_PROTECTED
