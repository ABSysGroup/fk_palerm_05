`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dGo9528t07T2dsEuu410Qlz+ruV2wWps2xFaIreD9Q0ISs1c4AKehL6+sscNwE0J
awWbBWxqaFpo/WgA8Ngfq46xRRXaA8MfeQXfTWpKVlaWX83ZbFF6t245Dr0SKBT2
9PmZl7YEUc0TmRPMNp9bjoNuuN7iKeGFaBP6PYOjy0NIp8Co6xm6IkRnEvfb3tpx
wHaVZc8320s8jYiafqyj8lPIeEcXgaGpJjqXNl9cqKb9D6LIuBh6tCrC8OofogTX
3GgcDjjlXZ1xTHOLE1fWEgZDs8QhZHrzs3zHBowMystowk8bSzYFZWn6IbVdrwjg
7RxrlR14xa8Wk8KW33Jny4PBkKE0/Y46qgGB1P90Pj0N7IhyiULknSy2mnOjNTh+
KEuE9jQ63SLun0UULDpCr/2gq0oShD3KZzbULkVl5K0IJm5Aha2Mk+nPw8W+01qX
pRA2feCUvvNdzrs++Dm8MAV1/K00V1ArGuEc4zrgRgoj3W2OWDkuD5rrtH4Qqwga
Ibu8MWcHdb+BQO3g6etrIokl2eEzPvyl+u1Fv/zAdNc1f3eVU3cfEyMveUq9IE6/
VjUWsansiNANjThyXh4YfSDDINKbA632whgYMnXUChdaiRm/XuM20rGP/TJ9usHy
ScZXdiY7tcikNndbwHqMfOZ+El9ln/d/XJiuiyXnWxNdHIyYP866+2MaBzUEXzD2
+nkklDU6KDQWCISIf0TGPLdZYlWPbXZL/N+/eCoxfiLBHBjxj/eoOzOJh9agepB0
m66bJJu50+FGZ1hFd03IFgMujJhYrXnAdM1Kut76S4cUV85SkPwcLf77XZyeg37/
7yeLvTWZFtyWlUpNFxpjokI8Cg/lViv9bKjfaxeaRUrtSr4et83PStYR5bAf34J7
b+gzMLUzxmVNkJe+nIR/lnvLUp9vJyDLhSFu6pzE02PZI7/mJio774/jcNQnyQAh
ickHfxCMNSyK68OFdeY9dtxd9U6+a7WAl2horXOzWdXg6LPplr+i5wEbyKhgwJA5
Z99ilnLjQCAY+8UMWGejgTrq7OpYn/w2UaBFQgSie/CaDwsXumiLsbltg7J/kHtt
/PzyrZesiZFxq5QYqWJK9qq9zZ+6TNUGgGgoeutUbyVI9i/Q9EG0xZM+4UQ3HU9a
n41xbfHJaidBpYVWRfwbc35NvLLTL3zGeMni0hmS4pVTULGJ419cCdRZ5hmkO3+V
EDpsHGZ7g+O/Uvgnot4830wfgTVzQRLQhw87qSZOqs6nMusKa/Da8G1i0AMBCF+t
NExtLLk8O2gQckzjXkbeWf93gCPA4Xj1vhWzoKvZUref+QCBBwMnMYVIkbqLZW80
zko2gEf8rqxWH/WMl2pYUbX5l8Fc8BRuDhjV+7GXgUmmZtVd8GtETp3s6uUlzM1D
K80Yh33ujeDdKiEmj07c5r41fZJNiXKghaxzjAs8ykKRORBPUeLvUWk6xEc4mRSC
DuiyWDbEzDrbkx5JneCL+zOVByZh3Yo2GXNBZO+dFi7Gdx4M8Nzk0u8ooHxuXL6Q
0kT5NF/z36mUmUpUbioKGo9Ezcp710StquxI1hp7FGv/yQl0gV/7HR4/LX9JE1KN
Id5QzwskvYOCwsQPVSF+P/K/dbTHYstPavbOdB/TS0BOQq0+63St934XCKsYB3lf
t+CmiHrabWoMJCNaHqQjNg==
`protect END_PROTECTED
