`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
25Jkndd3yRPFfDr01c1Hd0i9DnRVXm4VdpXiCug4qsFrxJ78tlJycBO0OUH69eA5
rzR1IE5KatDXzw3U0zv5KdPBXsX3DbuP+AJbWoVeMY+wus34I01DOdMhKQ5W82tO
GFeKlWqXz6hMj0DTqKwh+UHncctvdXG0ET1AsWkSsMRS3p/3glfsU0RpKFbCaxkq
u1jpLOdiAXSkXGkC7Biuh7L4KkXFlJSg5YxRS4nUnBIjM8TpUrvQshwgr5v4iSor
`protect END_PROTECTED
