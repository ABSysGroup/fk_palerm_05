`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MRXxfSKK/KIcPMIo7lFMvXok2dpBER57daacTNbu+qaKD7C+JZl3iGFYAJHPV75q
rRRHlqBlGG6qetu89ZjC4GhzVTExEKZ3Fum9AxSBvHmN4NMbAn+vLfMQ4jO+VZNr
99am5TewiNsvY5ifalYeKvjPE9idD9cwY0huqIQH9jKS0szGxLlXbkksn36nIbMO
VWoWRX0XBOGdF2+ouekHMX6CsCn2obtM9Euvgk2iMEJuohREAb4VXXKi9uUrk6CQ
yT8NuEYQAeRLGzPsh2uGXihaie26bl7rFP4lfavFoeMqezfFoprI9axkrIBqQJso
QFKLWRw/Yape0yJVPZq8tOvUFUPJJ8qA8q1uwx7HSZsG0JTtgkfI3xmbbrr0whCp
fpWD9uTuSdmMLW3Ar+yAUAac/mnOEctn2/0ANumeVQtPZdlxxt0SlAkImItXJRzy
lkT4pN2KDpRhaTF7yvdHe9df9TknphCUzE8WSUZ4FpGySOQ9jOodvjGn1NYRgwZH
lZnTjsWEyYDVP9hsKMsY77KveHkcIu9w0gCcKFEhvwpv0rrnoMqucyvGC8RWxDdZ
Ymc6CXjvmbGoOcpvToUEKEu06nSDHTYnPNh5tNduNua24ZW0W5gpbopU+gVHN9uw
khwA4TIPy2A2re2R30azBUybswvM783AJSinRyku6ja4WpzC/SCN+9vK0e9Hdk2L
OiecKvxjRKjAHVaYLk+s61AR4qKgKRpOm+FU0G9ry9LCob3d3uk/IbA1aj3UVDM1
8W9GXmRop7tno2t2kHtlkLuF+5lrzJCJ6UIfMG6q2GMi/akGEFm6ZDiqDy+0HP/n
YwMT2LE7k7LmNubFTnYx9n9OgL7HisNKI4HK5n02NVSsc+bOoEDIfFE7+Wlmo60y
mBQc9WHmVzapGeJlWJ2B4UXrVDNhKPs9y2Z3V2KTTj7qlSq8ca0RR9t3gsiQAQMs
mch8huQ3KXUomAfsFE+iP3boZJhdAWs7HDKwAs9DFGarAQVaKsu2C/J5M3tZ/E2Q
mZblf9EuKwgXKmGzXZSlylOJfO5mfKmnP0L4oTGzc05ZWM3hSo4YDs0hJOYBgAdO
pBsAllucQ0oH7melA8dPIEPtdfvYxpRm2s2vABFhJut9pF9Nk5eq2S12v3TPZrQF
vaKQk3govUIWot5njMbwauuSXb4Teyjfl+r5Pv/1FzjZ6p73vLCm3JPQ5HpqE/jU
77WSgRj5MbgMzEK5YAclwGc4CKBRzKrmqW2c8rUdSCokSLoSx/Ltc7PlLbOXViIx
saiP6Xighb4gIGHvRH3i+53LWNUsN6DMAdepDjKh600zLt2bsyNoI6yzFwN9I4Pi
Rp+QlBAIpJwLjiSD5mIlCfj8SDnMkBPqriYrz44iTKBupgYRD2P9RsxyEiw3nFdu
MJcr6M7QPVI7JSP9cAWETzN+XEeOE5ynfwvIGaPWBP9wUMjvXn58yGtZK/LB6Wi0
HW4kZ+HhfvTGtkFw8levMmrAQJQTZXwodjZHIDTvd1Qd77qGP8OJlj/SeqQ5y4/K
nD7CBPw7aUlVfmCHnFZDKtC6YMOKp2cACQZ0DiJSCRxOEL7dVbXdVQADWlfMhH8g
TxTSUuZImKEk2eY3CBXYRghlMiW/NjqNYqjxFEnTSZ9U1igphqAeJZg174+8qrxM
smVYbO5es8b5RO+NKFClV4ccxnGjkPLxBEmy7ddq0Vn06RLIidaDTOl1NIYkXQ3m
CwUppyHaSaCqsX5rIg71cuo7p8znvXS1Yc2CZkjn2Jv/iov4tRPY/LOSjaiaPqJu
uyR76TxygXIZvS+HhNNWbJsPv4M1/porpnrFeDYNDlSeRF+UnCo1Kt6HmV9h+oyZ
yA7rsHXN1PWbdYLZi2Vh3PzpPkCHYSwuBUqQnbzdg/WcRg7ObkyJX+mIalso2wVc
ObYZjM6lSu4y+j2wjZb9onujy6RJMZjixsSPW8f4gWeechagaR8073XavjybYlff
NLqrKTIyjmPHKIiou3k9UVl9RMUdeURs5eAAwkCeWn3Y4Z9KmDvWqDYm5d9BRCn3
2OX7XqRTLdHIjQoDxl5SaAsjeNkA8axWG2H7jAT3CoQaeROv8/OBCM4qNBs7RDZV
vNmbSF4PXHTh6nN2ZJHks7qxDVMoL2LhtD3lVACi0Qjr3lPbHlH53Y54KDNEgpWj
SwVj0qmGxS9f4rjnoBwrm35SBwNPjec/SrAjBNDAKLAbBcrOr0FcijHa1cNjd+b1
KgE6fjwerAE8KTC3gTLbvQYZ1SSaTi2EjLSRYytiNPtnqd3cr5EsRNfuwQp/7gpq
RBMfaK57aMjh3goL3FHXGPTV+GOqgFb1viKkW22VBabSDgpUuEMrKDWwy2EiJwts
QqDrtsgMCvtbv65AL7f6swOH9nxSBR3hcuNirNJYBKp283bDqYw/djy9xluPtb6s
V/YsQ34Mq/8rBH9YvtX1ASCIUCxGQDiKnfzOVS0/U+jGMUuZq9DrPcXW+uPN4+uN
KqD9yb1C+h1j1GKhx4QS2dCxqHG/kZe014e0fDE0ER59LMstxTeWuRAkpc6gM4uc
b5Cg4TCmwIO/yGOgewr+ykl+Ue0UJL3+zsRC5E0+k6c2wiuEv+uYj5uUuJx0DN1H
HNIMp8+PNBDFnZ5p8R2rq9OkezzD7D+FeMNC8eRpbgyzVnBTzdYoXDpjx8k8/Mw3
TssNA12vcOCgInDm30IE9fVSLDHFdhlXe1rfnY8+aPi4T9JY/Ff52IRnLnvjS2WT
aAgKcyNns+FJg8m5QmzcLTtzB7f9x6kjUDAUiD9jCCgJCH0lbGjaPoNFPSnbPHNP
jnxw5fiy8dKL++zzKYf6SSNj0/o3Q9B8lKbHAmG4GyD5VgcnX13RYk3Se95jIdE+
85oMK1O6W68HbY6PqZU1vv0QE92O7Kacq/LmHzycRONVaoaj3QlzBJopDiir8jGP
ZmEgvyml5m1O9U8518Ye5Hnw5ApePcmS8r13qZh2yFFbLew93//WiSdVtC36iwr/
xWsQjxgG2pn+RHKIOhitzvuCrPMIW3UQ8//06BrG94lM16sWURF0pSCLLxvFf0Ac
Fmc1hVZ9eKYPvQO7st96C9+U5rFsnw8B2oiYsYP0c7vsDCsdQRZVkvHzrypZPuu/
hEhqyxahzNOkOovT20JiLGzrb5E0/lCh+x4HRL4qA9dA6IGdIN2cdF7rXUFPfaaA
bTqF1/QuEX3EXNx2rO+kzpUw5kJZwbpeYc9qpWvTCQmbpWwMwelL8eMNXe6fzKVN
kCXEnKoj78XDMNJOfLEFPFTlZhS3gmAmEaHBoHysodw0j8nDkW30l/tw2x7+xtT1
zoOoH3XOtW8saoewVd4LTQpHmuQsUJs1D4ERrnRjEETd5UtHSo2FlZ25/vPCQbzO
pxC7esRgFO6RuXVY+Oa8Q8tQy2yotaI8FRV6sOE8kybtMdW49jePXJipaxtndzJh
dCv7C+je4jpB33jgL5ZXL0OyFdbKGUBIgg7vYs/6vb6q+AYvIVB5CauZbk6e4Zlc
SfW5WYddLTRmd2kiPiy8A0SuHgs1OYhiVXVb9K2qu0JRBrrkYVf5EupAzNtsY0bQ
6G6+Z1Msq8S15CgW6W+9FlHkHkmlRp4pcm4iN8g1hYHEMM9IZII0FJZXLyuaywjc
4M2M99AJH1+i3alPZq5MrEUmaJqHtuOgxHUQrIK7yZxG4keD0X+E4oBw9Nbi7jKL
9D/9wyPBNloLfyWp749vnzwEo30uBo+Qa6lNa/JgpC0LBbaQS+GgvLf/d9cHBUej
Ygs0tX+qJ7tVn7hChpu7YV/pcWGsd4MZ7ZT0XGO8j4J4Zco5VIMyAhVLTlwZ75yL
RaiV1fxA0CmAXjrXJB7viaePx2eLCmqelytj6dLbc/76K5f/piRR+bkPb5VBALR6
g7JfLwrWR047Mi4NzUuE8wPGx4Uu9CoKxWcjogFctmzbDNOdhxSLX9w1R05LKqhr
prLfL9wAlNrN/bW5yNqRRu/W7Mog1ufpbcjPNFO7NgAZoUL2fnrp/oHGiRPYY3gk
DWlHNJBMynWmteP8bAim7FHyxoR4Hj7g1dfFvZrFSsobSMxZtBCuow7LNI+1Hiv6
HJSSVaBMqAZ/ZSAp7jDhyOq3xWP+MBAKMCaXO4Xoi/h12uAkBgRbgOLYEaq2Snnm
OVzp1r5ISHvBO7DwNgpKRhPuiRFTKe0aAuBHEeGT4cIFneHtS0rPuLx6/iNWdwzN
pwTwE4pCTHs8TTYmxOswHuP639o7QBZ+NlpDXZeaWJ7cgPZjgk5ao7iynvzxYbZZ
xZJQ8MH551hV5bmLoHUs4INLtlfHYx9pH55s7UOzDwh8WRBan1j2hwMO0c+Si89+
8rkIRZYtsQXE7IXBr1090Gf1oaCCquDKfxLd7seBHK5KGRlhmniylJfupap0/t3J
93wKSmN74DDkoz+tZwAD1FP7v7Nt9lf0xKQeW2u51BAu/bnVZusvUyx29Kc31qWS
sxNQiUWA9xXrVFxw77QR6c6BJFAqrsotp+qd3UJJEEFGpD74LD5HdTjR5c0LnWDJ
+UwIXPOHn6n73AaEud9UPsTxjdvewbN0DdjOYd/tJDBnArcWxixWVNSlvw2cREYB
r+yOvEVBMeY0RioMo1LYPYHkxo8jh7swXlzxom9Yu9BB0NATyRclAxWrCQJTM9Qt
8xaPhlfJspZs7cLlf8H+To4IOMti2Vp0HC+3+q5+WHcI71or0R6wtXTIayXgs8O4
4TbwK/vUBnodIcYhNAAP0VTC4+alz/iUsB104gr8xocInvti1GmP1MF7A6zLyCQ+
O9Qsf/9nY5zLYe9DJPZr1QpHHKzOyzExvIZg+ekAHPHYo/eK8GS2T8TZ9ebiHdl5
qJ37mOjQzh3R67cLyusDx3t9p39bGbnuEEhMb2V61j57Nip6Aaa+yhpkRAdAP/Et
k6+gOsFv18orNtrCNI64hoscigc31FXuQ9OUM69fU1WB0kaedJto2XmwdMJiBfUT
oc+jVfNZWgmSzJFsvzUyqkg1UanGkFjfPq4JhkfdOUVHhS31S58xT7hhcnME3NtG
xdepL6/IrTB/MUBaYC7/XY+vur5ZGYliOPOYxsRF1jFYSd93gMcUGEoUGjvgefCB
D0FZS8ifoTzybH1XGfamDHTguRm/qDr8SS4EcaBcGKh4cjNsuHsoU6nxzM5+cH1/
rZ8z0dLMzNm6joQVnwWv0Lz5UTqMzutRa8Wi6q6RORlbvjwjYGyw51QuTc6BZFsB
5OzcMTCZIXgZLRQOi4GdV+LrpGVc4YiIkr6rCLfkucPVW+Zlmw4QIceDxodBh4KH
7rx1EGt5ZcCQ4puqf+u6f/Y5YHXbVjObD309DH1FI0nJWGh1Vr14gZlHYNQ0g4MZ
bGD+tNiaa55Rwybx5HdU15Ia7dPhKlb9PcWjKx3ufm+BhZt6veTHcFeDfqxlozVv
i4NLiOpT07N8Iq8VCCiKsLTkVYbFayPTx+IfJxTcNZzFi8w5URa5ymCBadaBmcxX
uNPv3ghSLQOVBXM5onBAAP4FG/licUTgevciQgfQOz2zKN5GKFJe8OxWmZBHoRvA
fWjIoOna/H4++UN+2dd+0K4DvQoZHTiTZtdCqcZmtJ1+vIlBoLcCBOL5ziWLaTtu
H+V5qBvk2IGqQ3gJSwV3tOukm5+4WtCX9OasEaV0Cke5coFpgPdcQqPuTY+WLPjF
qELMtU3Qtp0T0BqGq5N9X6INsZ0j/Nn/IcKTQorjc4XqV5N3xhabYC/34ipySMkB
/wIRVxEvQPt9VFVJx4LvA2gXWMbJFFlmt4aj6+CZak25BO/fdu+7dRgOTQIWMggY
IFRzYciqnQAgdfEmU6rsdpz7j+OPVuRGtpVMw14Z0zvOjrBDttLh4WACvRtf9MPm
+/7AX2XKphmryqNRJXYHFOXdd2dRyTahr1L372xX6htu2vGpBFMBIk6sfoyAwn94
5pjn2jAYHv40jSr62H2GiQfJyAq4o0V38lgupeSDO3O9ox/CE79am+91nxjaUa6e
5/vMXBX5X4kM0yTw44zZdviJhyP7PObHSstvUn0Tt7YsLg6YRQaB8kk6WFvOhlPv
Uj9P3m9ztw4ROo+qSLeVsrf946vU52YK1W/coP/QMSWA41Rap/69BLl8xLSpzXCA
umbrHUaclGU+XxUsgm5aGsH78KokQVCCczpOfq27LcGC7+usYG1Rg4Fm01oi+dS2
8Iir9nZZ2rO8zTCahJsJgT2OE/FmPBW7xmjyhUFZdy3XuP4UIbE/4VYlRdCj8Wzq
+qWUo/oYLZSxns5yL1gOmlV+ub5y0jBpVnYACLzyKn8+Cr0Kbl+1WzQf9k9c6nr4
s3VwCGrqE2CBnaDr1rwhcPHtJjRBxOk95yJQRGr/KRzwETEsjzeABSQV0Eod81TB
7HGrUr8KJsZy19H6lJdKIuva6Q8SbfBWuLnh3/Bvs/HYyPAkkyTDrJ/QRQrOnODn
HEcofdPSbIRpgU2SW03D8Y0WlXyi7efaHuwy9yYGHD7qSjLM6DYnv8A8QfmHaw1I
xWQ47KcuqQvogXMW7wyQi8fPm4CPaMEYluk6AgehD2xzqAo/FnODUlJURM25D2o+
aUd/M7OQYmglzUuTrmsXzVXxtAt2sH/B07jFeSgPmunZq7RgIaGJIEpjvFK5UcBo
m/rCngJWoYGrv99I0UsW6o1WT+Tfp9tNXQRh+Qy5VuS00q0GctTBhnt18/0FrtEG
cKbBHZqf+aGPgiGRvodoI6TFfL1MYPgfjNJRzAzp2NkKut4KFJjAFw7oWyFgnx2P
GGjbtY2A2BZQw0wYXiWcNKqvfeGKu74EfMM9pMFD2H58G3Wp6lVRXAkYdty/WytD
QjYLiXejptDdaKslYvNP15m72t+dbOEBdAZsiZZO2L4t8vEkb6DsRE50/xIwX6Y/
syN/t9MA8e9LgoidiCyKARZjiwtLt6js7v+R/vMk5Hj7TA8vi7RxJ3cUzVjMMLCN
DdOJmCm5OukGm/sM+B1wlIsX/sMjkO3oqd+zmb9q+MIRBFcHftBoA4F4CTcsUG75
iwr/cq2jeR0eB+vPisiM3+Mdc2AxwwLvJxmjFty32BDCI8Cj5WX+Y/rP+egoEChx
kwPw/nOsiJpsHiY8YTseTGd2u7eB3h1ztM28tnUTS9YJuxtV7ciI8nxUvQojYXRo
NGpi2yzuWdDtjMYTglkpaeG+Z55tP9jGnTmVSxBrUJPfPfbSK2v4kCLhIJ6cIoa6
99yDv7m5zRGqOUeAvJZnaCRr+4aRHL2v0BTviGnOnCRAgfdAHJQO0RWsP8oTaruw
UhRfLykn8ZGshLM7Q64p3tpgtagRwD4PlttbOZGs8RjHbD8dmrxP8VN5yXgtDDP3
tqP3o9S9bnzFILrUgI4OjfTPlHhH90e/nAhazuwsmxqFqlwuQo4Prz0omHszJ82Y
T2UAEP63ob6BAKpMRBnpBDILKdSiLFPpRkkUXJcQNexGyqQXcG11hYsmS7P4S9gh
cq3FhJMP+o029C7iSSCJZyp/x4ueczwnUJwJXHVRsowBDfpEXTaYBSsSg/A/rAjt
70zBJ7u+P0lTL/+V/pQxG9uwr3qALzHfNsyFMRcmgo0iISb/cXYKn1xDcoOv1ee8
T1wRsQK//WcjdMFo3KurLIDWTI9l94RqM/+KirYiZAfPZ3x8pzMRxUwnsOrlHImi
5ZwjOxpwY8SqbHcfwcSOFhtVquDXQmIJ8Gj2uExgSRcSRo4PVftVOh/7Y2Wpm53u
3Aul49u+fX36uba0vygpHd0UzCAK8IuAc3GP7EuwxoWuWlWQtgv3hNIAOi7q8hBk
cgWMgld1c/RJMqklZRGRW3uxEvbpJgu5b5XUklUzfO7iWEwc1/AaLBWBjEaz7i5p
vAFU0Gg2sGqmx69uL3wu2cziLjy05DhDyWQqC9TORmz/L90Yx6/EAUczo/SUN7PZ
nNl4FRF0rsX019WqVUw42Wv91qKw1EssAE82R2fKU1E11VhVv921vr+LR8zgfAfz
TTq14mIcr6oOkqQiCVbscRxDObngVMvWGliucKJNc/TizdIh9EpWyGK2vaERdOW3
SfSrOx2KSLUPHRU1bI8G5TGTiSoGPQn/lETh2hEg3RImlwkhnBc+yuj2o2NfNd5V
o1SZS9carR7OSdcARpXCxne/cOlvV7Hvp1PqGgiDUTAAZ6zoZhHq+tMnrewIorLP
sb/YMRo4eCcAfV0zCrhc5E2AKfzY2RxmhIk0NU2XLnBpeUYdfuZKhffRgVL+1SO/
9ua7mVzPXezWyRic1tpePoIVAdlg9B9ASTf69BIWJHpIkgKGW0kjUVOy7S+JPTEf
nzOf5SuSaWxxPeGdIxe9CnPF6VU0Kr9yiNHtvABmbpcpNCEDt+uJAX+f/MbMbzZ2
9cgtW4i23+l2EtIoOPSsHWyGE8WyDcwYSoXxXVn+d5/jUoLR1cx+nQMcuTxvoCEM
MY0NlGzAwXyvM7/ZqTWNJLnw06uSJGUK5OYk5j9TQdG2I8Efzo4E8yu50zPyc6vH
rnHy7pNqFBbrQgKAsnNDLjlAMtfVLsmGu+P/2L8jzCg3pUZzDgzBKYcqm6qMl61f
/7NFWZGAqhDVyfHNqBLZDOAFYWr67G1qdHIm3UVkcxUqiprzzLoy+3aX71psTbt7
4De7cePTLX0ZOAln9ar1cKnjM3PNQI0ydbFogV7HXD76SCPk1awOE968QGippHbK
fAT8PsiurDt6dsPv9NdI+6EM1ai8y+Cxpuf6WPp7R20JNq0if87/2pTvT3/fLq59
M7W24PGmyn+Ok7bifdhgoxR+339rN4iCgcGAgJgr+O18HnR7/5DTatfVDcH40V24
LmvdqCqKjOKye9gUDpt+MILsWUxbQsvIyhJPkaQn/s8Tjc+/lcCQBCfEn9EmzkmW
7wHId2BWut9uWjD10oY6NVyCx/IEHADtSBtxx4+wS/CqiGwsUA2fYIFt0EhCJ2+P
55mLrPVM+XLhUHl1zZwbjheM+JTiYHkz/yNivX3KuZUNNQAWjoF/id69x7mW/W3G
LK3Ev6ITH4o6mOJannNLos5jDEKH8hPDzj/HHBtlGmQzKm+Zgp+tmpXr+5ZMJfgj
yDelB3TtlepgDAqs+MF5g/CnapO6mo4DLJ5RlrdRaY96E5SFr4NdLnJ1qbXk+54B
1BkmN6AaXY8UqbcTlqyQkCEmNJ1l/Cp3SQbSS2m4D5Icf4mbVQPrnsJw+VKqAD2h
wiagSfR1pdDoRC49hbBfZdSkdi6+vPG0mgafdEB/rBUY3h5UyXzLMOFCurYWW1LN
pKSo0jQ2MtycuJwWNs/4Ft6VRihjI9rAVZ6ezOkxU4sbzXqD9dJIv4hMx+PKHKPY
pFGPa/ujZEOHw8PKX0XmHsOgw2/8m26C3lw5PV0jQGgxGjgIuBl4gq2+i45b3UdA
HcEnAnJqGkTN3WJ2ySd/EONS5VR7S0zn/pEGEWSiWdvILKKa9+KtVi/lJR9Rr3Qx
Hv18+q/4oVAUbgG9i1xImiSC3rXXY2K7b8lnSDdgAW1LYahpCI6tJrh+hXcu9sy7
/xB4bRSFpVFl3PGWIukBYwpzYUrFqNY/ic8Gx6DBgu6vEbifd/9apndapDc6DJ8p
pE9gYsYOcOhpXSuzwa6Ky4H9Mo5hQ51vXsrMhRtNjrm8jPyluGBAQlSTLOV8m/xS
CT1N2mZ2hfnaIzDgzf3laTj1fYPOIyNJMFZxkCedljtt9KnZpFecS1VlWzF8yCPr
/vwjafOZUkaiPXN9K1jC+QmVVB1HPhzFHUT2MoaMvJ7yFQJ/Fm9k3YU7UiaGyZiA
BcNVy2B74Mw2hLO5utlYY0KmU8rWkAtrICw0z5a9ofO/pjzBkHQrBdHlwe3Qt81e
YnUcdbJRZr+iZUPi5QukVE9JQzvuLktyJ6zi9HbN/hIK+ePQves2i5mAaxNuj4nj
SCDM8oVzdQ9Fu5vFXH15tJsueg2SUz8BeQDnfv6iizr1lwePjtLWY1rNGmVmrWyH
2HohE4QdV2g2+DvGyX2WO6yN7DWC5f+gzSNhAWEePdPA/P2GyS0UqLIdibsSP7ok
kFjfuzmEuLeER4mAjSaIKwcm45hYwcfWnB5CcH6rj7lMitrrcAmvoDP6xge4tVUq
EjeDCexzuXnrqVjbjMyo6cwB4E1nh+ACoH5UlJ+UwqPpFVyeZBhoj27X+uqUKmbJ
z6h11ish5KfliEBMGHjcBlKVEaHrMOkP+X2YhTh1vn4NtkjwcuA+6BnhSIqyZImx
SRUuZ5MQHMXyVMAcLSz+hF3ptjwhNnl5tQAiToF8gUR+IlLkMUVP4Xn6TW4C52nM
i/A9XOKLyGepsnLhylUzxBNpX9on4PXoi3SqW0kdaJ/oIQhLG0Cw3GWshbQkOc+N
tt5YJmyG5zXnVlL+o6B9lc0c5wa1YPGyPnBgua8xR3jx+yFkPaIt26Hu/g8EaPnz
bA3P5syTYO2fYMUWPYQjoh9DP1xMHEkIhixErs1LdW06RIIorgyt1c490ytuU+Gb
NlitFFgesMxqsvnO5h91syYRt2eT4ys2JBi5UJlqeWUQr0zMnuyIlQs6EcyGQKUM
nikZqPrLD4HUn6E9pOmbJksVH44+srMPMxA6e6NWVZ8zQPhjYJ3NgKNxcCAFqUA+
GyCDm4EXedJic0OlsfXGDpjRUjyK3A0cak/0ABG8+U49rZbwWLQXnV9va3guRVSs
8VwUgp9uK2hJYgBpvcPPTcWRZOJJiqGWvtcP7PocGUDLkO6jFYOUPbFaZMHh0xMy
RJ2BxnJxpIJ85IKZTqluox5a4r0AUzBLJ9hSGUWs5mFngqhN+bnBS6+HtyksrmrJ
PP9qacgeagekXekpvmgV0XzHcC0LtM3Deup2IbFc5RH7Ht5OcxAleQ+A8KXXerHZ
C13d2wozaTu3Ngy34HZHmZ84D1LHs4GklODjQRTKc96fSbdvkOun5G35gNiqqy4F
fxJQQOza9tVWYJvN2a2Ucr6M+QCGpSQt1OctbYWj7PKJOCh/jHRjfTKfYvIYcz49
mXcTrdR1r/lBPtUFMqAYZaPLwk39/ihxVe2FfnS781WaE+bX8cyi2B+LLbO8WRGZ
So4ZN9r/0hKHv4XDQ2rXlTmBlwItnzJgbjr7Xqwp7W4rj1VGdgL/6DdeB382ETLZ
D4Fae7TLVdLYKrJaIH1owaU++zC5JH8Esa+qU7If+yCJTgjsy3HJF8h5lsw+y596
bN2g1abKHo8YEFC9yKUW4NPUUYdsKmrwtsEXLFA1d+d8kHgM+WAJnoBBC8mr+HCB
Jq7YXqjs9zjy7M9vN/LRNGfJySgogBItoyR9N1RGKLdfX+r/9Bov9ttiyWhPqDCe
fyiKms74tvc9axV7H+ZqT7BABbu0T0DClHZWu60C4wrRY9KG9bXTj1An93nCVcEL
8LPFKvedwjWoBHsyIlJcyfcc4XGbDWp0L/UUV/DeDdPRH2SFSGWZU5WfFvODrDS/
C1rbyhxZekV9UFH8uIhV+maqW6xjItcxyeKe9hutR+Tnji4axSIFhARWyy+L08Ui
SCi65+lQ0fPKVA0QXQtw0uarhwExeWD82LPxa0VT7BG/ziQAsKCCLyNNZM2hYiro
A7do9orJxPTGrefJB9e+/7ojkPPihFd6Ofu+NVJUpmxIiiLJRElO5kV38ReDzaSN
NLoCNJV0+RB5lVtSu2jEo16ld9wxpobw/ux3EmNGH9+4/0EbzcJUhijyHHWFFjmn
kMJBJL15ZRqK5pzKZp0bUbYCy+OJsQCipIPBPN3DstAi8gpKuhG2MNrXwQ+X21Za
ZlcRIKXjMaTpRX+BdRLxkeFhUq6RtCl5iq9tmfLPytDn5ZL+XLp+sfLitqfRkxs4
PbdsUQFxlU0jU8sL+4+ALScrw/E/pflNxTx4UO8Uhs+WP/HiSCkNWUYTluDwn+LW
txoWyEv99qqRTRVWVMbyzl9dxzDYlQ0dhDg1z7of7beb/AtknB7L/acbT1jI0b5v
8QEJVsHmbTC1jRj8hqbEjWGdVBI68rG1kfjCt75G5l7VTkUGfmzhU9ojh5WQT+ci
RUaIato3JInkfqBwVduVTpNMEl6Erg1XPv+7LcuXA5noNPEN7vQXufdNYGANU/vD
tzj1Hx9DOFc/xssvKBwQCTfQP/pkJkcdIVUqnriME6hEsv1GY4CaftLMAyGiXu4g
IA/mF0wV6hwmz/3AkVYnf/KHb4LRatEAgayJCMmb9TtywXEfqTYP97lyesMzD4TP
HWS6o8VDiBC56J7KQLupYj0W4VyYqT7zCQzOhpDI/w8FqtpmJhnd73sA2DO13XNT
dU4v9m0ZWhId7k78T2BVsmidHJPLszyxH0KYBguJhVEagL0dj4lGN9ZEoOZsqtAN
g36oLiGK98nltyEhefFIKve6FEeoYk+vrDCXdVaFp/ycNtRhsRxTQaGGhCYrxGNI
dSMNg1WD8nSt5OiNXhnzGmw317bWEwi5BVMkCYXb3t03NiIMIw0lhkh+4D31z0MJ
KVVWexbgZB36ScD/p42cWdTwrhuPn1zOcgu4YF0J6SPgt5eZHfkatiow8/FKarWH
7LwPMr9yvK50sgK2RNOkYrLdR+RygcLAlqo3Ay0cQTbM1/yg2FcNAydcZ146Kd2b
OeUX7J6rW3ez+Ts3a1fhzyFyqDqD9ZIPs4jn9jmMXLAyphUUf8AyXqqB1jSoNH1b
szLVTVPeJUXCeZyw2fFBqWMwXuL/9F1kQ9U4met+ESOFautUtbVM97z5Gk6xKo41
vvL6AcgmGkZmjrIB8pBKglkDu8AO13IOx2vuS+PsgIlsMpVyK6O4ATv9z1cJcQLT
6z985ppjvakSYDqQetLI3rEHv/xPbb2F4DSjjIfceNfpaAkad/B9aGgQ2lyDclMU
fAukxF97No5A0P6cOzOk/kl25/8fU7M21sYjinO2stFI6KVEUc1jzUqtEjyJrNdz
Z5EXrChbInTc4jkkssxH13Ia5rSHuRSeqXu25WC8pSM2gRS44yWi7IwNpXa8eqPs
d37Jg3Lk/luNwRtxcUCRyaWSi4SkNDJZm9Ro14GvIOgiWSwDyp0YMufqTvXPAgjv
dVw7+/S7U0k3o8teKc1ft/yzMOP1nMgrTwHY2DLK/o+8rk25YUFrsnDhWLMgL9uK
dM5rFOliX+yOnPHWqih4xvSEy3pd3KrBnMIqkEz4opQ/MovcXSRKva91FbYuOr+i
cbUBNJEWkKPXpqSztN7FqXP51jOb6db3bVfGJyWoBl15RaxVxL27+XRG4ox9C96T
izGO/XiT4tvgam0ab+DaPdfxpqxT3QfK/50T98Fw0l9qMtv7boms97Fq4kJcJLL9
ru5fUr1rUEFn2y21YDOEayiHGYlRGbz6DM8bEBUG5J3WQ+6JIdl+CQjDqOdS2yQ0
x9t7EvvKw9mv9sPA3kqPtXKgCSXyXhWyqsk994RLqHBslvhGQJ0TdFMztPIp1yqx
BJRlPF7mW8oyIWiXhA3mxarphLk9TSOFutqhPCTGa0oh1wLcYJYghjV+jkFjbiQ2
vIUUyiM6jLBbuIEzEEwfCHXDCDh9jLUnU5m5hbmp+vT4yqSkBdRhMpHyzXJ12yNK
PLLixLPkZK59Rq/MrhGAJIOmIVWsYlIPrB1ep+kQiUlr78GwvPOcZE4oUKTFCvM0
ieS7eY2XkRU2+fErMeCJsEcdHrG3Pypfji2yzPmc/wyCnXn/3tQIJ7o1Bqs4XZyq
4R0ErKHNqKVJxPuY5oAiEPGuyURS4FW2La/JVPToHk6Okc2IamZzt0cCQpvAKwyn
d/uEyjjESwdOidYFWvs4T0uuvUO/MMJoWjU2VejDcm/8BN3M64/IheZ1+xYqaFyX
hyQrf/FvDHxOYIZqqwdlhEnEz2V8wUSSKoGpPaTh/BGlBfoMyieUQ4Qi9RivhRA1
dIu48cTWQdh1v7FTEajV2Pk0cxgFKvranyrsh/6Ir/euDh23QefWqMFWef8jhDkS
AYJ6RGSxwjt1osvKD4Be30V3sxNI/cetvEFXgjJ9JQpc2fqiLSf7TYODgqSDlwhA
Ek/DmSzEHTD43ZV5Ou0hoqCcP5GxgfMFwDJXK8OLk2SS2JLBXN9ntKLtxSCp0Xt0
8yaI1O9o48/rn9KCGoVy5ZO9u0mTtVTe769zJYTOvVrpbqOKdeNQ5x8U9JIgDFhx
/IcbpKiMULrTeU/GcQanU60Exh0THBcV6sQtDaq2RRzGC5cZZya7gmEXQNbtXZ0p
nEuMLFIuaq8kE7XxpYs9VuJx2CG+k3YLM2aJ0iRM0ENgXzwE94Nap3cB/ENhGW1S
RdUuoTFNMeufIk070W2ioYVNH81syyQf+bp2GX4KSUOzM1QFm+Jdjtsqxu+2cRXS
ey+87c4sTFIeGcohZ0dtK91Ov5cXJtYIS467HgFrGyikvGPVyHDiU8MaycYdhMze
FlgpoJswBRJai0JShY8o9FLk9l/BSSoBJrkbKZ49Dtb+wSqC9nd+n+C2060JWMfR
yDrUyFUQRrDmq4OJDbf0GqV++cf9QRWEt4pbzzvFhjwRCBwWjMLswA4UgUhlpEva
o1lIcuneuQWjVcZqlF28XPKKPt56G7qJHQjRrRI+0FGFyTGCTbg9IpVlX6t/46OO
+R7M/kCFip6ldGjI/tAghk871V5tPd/9deazunOqe291VvNmBvqj/FrjcXOtpP6+
t7f3UD5xwBjDCnD0dZDpnfoqOYK6pyWJP8mnxBe7QakQcx/KCqEGEgi3Wn2XbUN7
9G2n3FGm0gmvTElWVuzO85rwl+Im4SYmcJ5LAPrb/1R93P9wFARZV44gqvCqPNdL
z4GLg4Q0RAXIf/ygNxAXHe9P/D7kd68AZVTdZbOmIVUHOaH0eWdL1MPR/frYjhbJ
QW4aWA/NHL7PpXT7VDDLQKgQ7vFE8+1ijn2P4YG1OzkEPZFqT5RzfZAb5o+1C2EG
jzC2vgJh4OzAwblivWYC6oiNIOuE7iN1lbv9gVUMJNL4N4BD/Vw3OaNi2nZjcOpf
9PPWiZ7PEJsCwvyRFEVtiLYF5IMaXibUVFyOT0/woyH3SM8OqVE+l04Plh3ow+iq
dR48TKJsGByIDEUopajtPwpyMT+AdkYpjaxVyufxRDmIp6hdtNtJ70t310LU1Nkt
qFV14rtTd6nw030eJfSInARV4sR0qlMmK9eV4Pk8II7nHO21Y4bd8jgUgGBqYmT6
LQAVu3GIVUlLvpyKec+ykhC6AK7xQI0FBGjuogsyRUN75QjaAlklHUv/MzBwpO9U
rHQyexFDM6ig6WeLJikB8/ffhqK3c2CSozl0fSAD9WUBYIAZF0F5D56VjYe8eSg2
NlXLu8+LCYn+o9hOBXqP/9siWYtgNNdIX1pD9/SdQSDx4Y+3PQlqMZfvGKXB8g9F
lQggNcCQWC5++nS7NxnGRia0aR4b7dtLve9aA1JrZ0+6DMJZPTlceaFJfmTdg6ZZ
InzTL4jY/I+6J0qsIjdz6bivOrsMfi34Bd9cMOp4APmU0bKtn046tNQ20mlnc/VV
BRotJikTVYOoFaCtibsezne6nmQdR8IXe+dMemlQT093zMhARRPC80ATJTV6mP5w
17EYHiQl5bX6pvZItnh39fo/eqr7buD61c8W9zOnj3Dp8esbBY0lJJNLDOWfGBQM
mIRj6USqZ1HJ4p8tZILaqNJba/K9y6HLRQRd5XpVgws1rhpZSPoN+5xYXshqETQu
u1H4POr5d+yJIVjqHIy4qJa5WFcwv1+GQxzMgx0WObULBJNtAV91XMmmSLlFTisa
GT0YOuisIb6Rw9tFXPRY/465yQoAu74zvpnHaj12ILhQ376qFWKk5uuCIZ0NjUjR
b1qajaffHMwKeZG6qSzW4f+4pJMKtImVSe0CwTFtfcPOY8VixKtpze2qfCmwqQRD
MWAr2t9GrPnsh2E9IUcZCOtdgf5IdNTMFwL3APLItRymXRCETzoST0D8QAPGVREI
sm8DeB83nkCa+074uc2NwSYZ3rh4xwO6hwzZGRXgt+AgtdJamYGaICEZR6KZq1+P
q/uA3gkQN0D8XdsVVYwIaPhy1ldSIK2WG3VJ0yFdiN6oR4mwSKNMi67hwnF3Wtoh
sQOYl9TKhXgmK6RJ1c7VvjlkOvtxb9Cybah+TWZalRItSLNYMV2Vns/jNhv2tLt7
Rr1yUbnh+9i2Slu8JPfuVsBERaJlf+XJPE4heHA7c05vp4MQA42j+zMpHWNLqeIy
YJc1DUL85w97LWXFmBeIuMekgBvX0bwNVBSCxN0bUwz2+HZMjAa344R17KOwLL6O
e3pa1JRYK44d2sY3ajyVhnkXPpyPg0UR8al2MK5nmFctwaNBal+7ehhm4fZN5kMb
CHXEcD0ibXoZzNw15lFYpNHqU4lAoU8k/IENs5Mx+bF5mz568CcnhITc/CkRMpaw
UXTyzPbFleNXjYB7ZG8n4614B3IZtex/GMRcj3fuU2tCEZnIOm3yBEn8DYVqrZLL
h4bxeGad7j+vD36kApBjELqBt7yCk/93X25fYWcU9wI64/+1b5LRqnmGF1Jxq4Wp
vGJI6DQNVvHDgD30F5BdzzIQbQqodUTSFCP2WIPa3nTaQJE1I2jZZGF2ijZBjJl7
LX+/XKkPdQe9kGWxJ2cEH2q9bAL4603OuxahBPcglbP8eSln/Mt+seUj+PnhMp7F
iyKQ99sn/Q4ZS8eGEMeu4bmuDJ/Yo30kLwh9qvb7MBD2OGmIi1ShVb39NxhL/6uV
Tr9KHi9O8qgCpgdvUJvnlpFu070UQ1UjONDsJlUlk+HKoAj+5flvZt/qmp0mKzhV
FvxpM1fdd6AyNeM81csi98SLO0m5s+m/NwOyzFbyTJJjXbKbi/SP0RDWPFzIkX86
+b1Ui/d1lrdCMTkoAoh5rhpgu4tMXJ0lakMUHBEkZTGdeaNZwnJ+sbzvp9YGnvto
uqzqa43WfvLEEz7Idgpq//XJRxWlBYeK/ShJ/+n1/vMvgnzoiL6ef9romQCFCet0
E5i5IsrR9390c3VZWKACp4Ros2jRzh1A/AXUC5nsvQWSYB69p9GGguazb+HU8MF5
UiMnh6c2HAJdTTudUjMtjDbppLQoVfukv1NeLdfhTCsks/bCxH3PuVCh/VDc7wRu
kRG9+D8hqIt9scYYiCh1ylACkECkGQktCwG2Z1E8tZ5FdLcFuUfytK3KYIrA6bRl
TBvqYjra9/6n4aVbZGMgRWF5TQ2ELcnfGC8fsupjVOVAWkQi5OBlxfZ/2EDC7lx/
Kz5V8BZiTH6NKg2Dv8B15ZpFha5fQOgMeCCcKnVRUscgANipeD9BcLIjtMhvmBem
6NcuPIjF73WkjB7nsHDCCfGheCxvC9r8EFK6/6cnvzyxhSgWKVp4WLLXzxv2WFzf
BUdmXXackhIw9lq6Rb5uMgwaMzulUcHinBGIRkgJ6hD4anKO5El+6MCCizWKtoSV
w6gRHw55bLPI1+OVRJBQFV1mIQWmP2kqttaAT+/Hdpstbaw5YBG13BrGh5/kpAcg
rmTJqntomrTB+7bHviIDNfi231MIngR0ipW4rOFy7iqcXgzyUZO7kWxtJRab6wy+
3eAuURN4vcLFfHEOScmq5h7BH8jBRjpU2v3KuHPgh7ZpmDqL1KmoCB1gprlag2VQ
fArtDndFbmIYeRyIK0xwZ6FVRJSrL/sWBsVZJuDIzjFbtvT6tUx3dZTAYWcRYouC
dyc9xNwk2ff4BeY9sp73Nvr0ngsobID9LejKF2BkGc8Y4ZKIqpoliYuF1jXRAHao
RgbVGEqn2ZbMi4PVIGzrT8e2ICDk24XQDAfP/PvPEVSMqdYJ+OR3Nh4mj0EOA8/f
+qGFLonrORpo9aByBfcp0Ne2i2KJquNymvIObosZmGNsdpNp/V0liz0M4ygWkZ5B
EGyiEzeP7MPjjOt6cxmuUKBwiMLSAalL3m0wsdw8wCsMyqsHrM18YK6NWThhakX9
rmz0fTQs21G76axcvxq6oXPYFQpFatDlTmYWxUJedVxFEvfYt9xLszdXuw/lK3R4
7FEIOFWP/YkOYyUuuxrp8uMn+lIMaarbdnGA/r87UYGtevjTr3xK9N2F3S+i0n7z
mJmfH6c43W/a9X22afOFxvHkI6Eik6Xz8ETpr0Na8OC7ijwUgEfcm5tytva2B1xZ
XM32aRVASl+fARwxjSZ1/zIauT3k2qv3D/voID25uSkhnz4pGFb7ClE1NO87mjqC
bYTqfcDttJXbP9JQ4Rl50ou+zdk41Iu19JuVuF/JpoW/e+f3HMMwkMon4IzMi0cq
40e3G7o7JZDqckXIvUjeqKBLNIe+PfcXUnb1WcKlOlK0BNT83SeKmURHjitZPaQE
rb55C/5aiJ6afV+i13BIqkXZQWH23pWKCmRR8m0SKTe39r6bB5MEhPvx8YqAbbc0
zcznQ7u0jSzav5ArmN2CUIPQS1YwXzaJCzdt/rur3bnFmObznEGYovNnDr535e+d
dbHOVyiXIdGLZMW7ZOrkxY/RZZCRHD3nm7gPshjNpAkjfN6w7ubxFDjxv7S2QGqy
OUHNGfFLkY38Q0Hr0qIJQWexvFYwbHZo5JN4exHie93xfwtYm4gyBX3BbpfhtQ3N
Qg3wlBCdnKqtWpqBCFQ7RGNtEthgP6wpKFrOXzsuabUyh/KE7oJAZQPHh9T7SMCS
BZeo40pQjsVGI8Vn62tNbTFMW3Ez5sjN7HTWKoF91bXa9M1miSCl5keZSj8uAizc
hC/uNjF0g6YtKzuEkXRpXQWDYBBnSbIQ87Dsqp6PLjvdVHJRX3z/OyELd5FMxJqI
Z3g2jvenqH4TxdBi7uZPFLC5ua0jTX/jD4JPzdiXlv9ps0OnMNcEAG/USN/dnMVp
WbgblBCyAXAIFdQTPmkrX6A3WYeE850BITLV3/e5CiKMgnvHrTlPNzMPmythZK6j
GSy5XMFrW+JengP4uBSJ2e9WzEIyGn5IiuFL2CVflpndy6ySBDFfyg7NF/JIBu8t
WO3Vcf++LvekoprzcyLTwrZzhmNLXlsS6TTP5wpVcIzfvbbvUMLwTaCQ94Mki8NQ
kpQ17pBn47bqbZLZChaOCSl9U7A15rz8v/JAMLMBQoN3b4Kl/B+o+SJbIC8XSa/P
CSvJteScbFqfGSUU7hWFqPgzdLVW24CKZX3p25+/fTxOw6UA5SXTBvzERj6pBdJ5
nJnBrK7IOTY1UsddLoX9nZWqGOo8N5LhItZY/zgzGUNg/uU9Mqh4z5ZTjgGMlmBt
p3ueGrxi5mgdW/IV23fYopPDfDDqgjySZjLqPCTSz6Dm5bssF7hK93SR2ylTuzoM
sucEEWI5ZW7vMYexnonTpJHSh4+4MUjo4ZPAn8jbwy0NrAnhg/F6wRLOruVNPAA3
b5TKvceGPJBIJndukq+rTfX4fqhr2u54IfWkmrrjPOd+E/kWHcYYnGkaCZYJIlLG
bZ/AsxVwtiv7f+o8bj2cixWlKzVbo5jCn1iTRn83e1nfDuupV6/x9i1JfCw7VLXK
5DqmPVO0P/WMloRCmn9wjnVpp7z6zQ7kX/I9h4UQE9mocIZa2K4I3t1jXAcKg+3n
+avGf0y8rVogreA0fYN0j6hEMeNRwVdgRqbrr1DsnSvIxzijmLCuAnrLcLX8P8Z+
UQWPX3n+tYiFDbCbX8LZqwcyW6AY1FdAKbZ6yDtMI4Gp+amRYR7TAJGp+Lzrztxw
2WTd+AXt/aFRT4PMvBJRrLXYGBLn8AwkYZGjX1eHq0na1nQco1M1H4Y/lZN3wtL6
G0f8HkpLNwXx3k7AKFuluvblLbwG2RMQLTddjcdCodmBsqPXqGy8TusmpACIj915
isvOpH+rZ5PmrQPJIqLLC29PL0xusih4lj3q0P7EzFZJi4i2O1EBCFC+SGystEek
6y5Uw0Fn9FLiyNwzhmoFHcU1NcxYl7AbhU+/xMJc1LQgemyDVlqUvIxRbnr6dNYk
IjEXTw7iPn1vIhpFUjJucz86e28tB3HoDKIxekboGRYoiZvhJ9w2QTBl8o5raZPO
B6tDZygW93Wlw1HMoqEvmPv45Pk5/S6gdZ1n/N7I2Qn+9kqQti24vp1EkTQBaHIv
mvW1RHptbpo5TIMdod20263cleivnaUIF6mCiHjlmVt5It/nuWjbNDXJiTGHcReH
iNrDsUxKFviPWYo4i100Dm618gwC0yOkUUu4D7oXxfnqRiogIiz7E3lIq8pfwhZ/
Leny0elTmyzaxq7h1HnOTlPLCT9fFMAvDDSnRoL44aOKu1DR9J6gK6fDJwiRPn1w
avRZpivmH2pCBv7p2xwg760Vk/klQlsBJJOAu3anM6D4ed7rnIqPhuvqzKpNxjUH
fwcbVjDR8E1vgI6LBsvHK8QIFqmIcOQiB1+gpood+GbkYbnWIii6LOabsVN/j9De
XoOQczf7MlVI2b4F9sT3hdOCeMGqeRstdjrEh53pfwQxjJMYEsKqEe/a7Znn+1FL
kXLw5QbSqD2GU+R1WFPBI3vyn6+OvPxZvAAXdi7vJWjEOG4QfwzS+2l6WSzrQDbg
54jUZiDxBWPTOkPgfZK9fTPzP2cPbvNsO6Vf/cHV6mK5b14mbB5V8wzxuh6dDzqP
S5NYLQ/6R0/PLndjsQmci7i++mnlO/WJLIWBAL6sw1Tajz5O2cz4N/tshNJ84RA3
B8+1eOAKHgMOj/2gpZMKGW90pk9zH6j+KqJM16xhNu2fqFjfBdCdPTyozdHMtyxl
4QjHlAD7nEQK/psFsn1Z1IjVhUTR+g4WwwCZyyLD6J1iW4jqWw8ZURrtwkoJXLc3
ob1KVKGrh/MpTSxtEiI16ayhAN43CjeUBfW9v2P4gjOhJOIxkIhbCApNvgNg8NFh
xTSa7uP/YfiBqQSIodldw+E7Lnyv1raODKFMyfP2bdYq2HzWLi465pmSWcGWYCq1
CT4og/RgzC2I97E1+ti6tXLAq80S+oLmAcoW8GX/aZp7Ep6wnH2sFcmLknsW4vyE
ewyAeTkbK2x5VoJBfKuTbaCmOcFYE1GXhhTl1q9LBvf9HthYUltn4CsIqKKevRqi
6XoCs+/gJ+5IyS0EN6lSfczzG+Y43N+ssoKDEYYWLzzV+C7Yr4GMtJuvBhvDKH8M
5dGYBVIxUiTqDOcnYT0kFRNkpMuFGTnTXmRV7O4bLrhfqNfT4TRcnarE1ourbU9w
W/EdRMmfHlGMO7GNv8b+x98ZWPM0ROA2EIEJwZ19sUICUEJXPU/PK73Nk4K/jXgr
YZhTSpIVeLvHRB3e+6CwtrsniInISPdWw3IDEnpRR/A8heaUPApAMLPL0QZ+0dR7
qHHsuSFvN8PkZGM08MuiW28mOUZ67izAtRh+1RaMl1zhSonTnEf2ziDjks9CHcDx
aIx4kIc+F4B4KzG4hR1GjR0eV85JxSw89pFDe7bPq08Mp9e7KhmMzoHOwt1htYqK
v1vn7bCs+wtfI3HSO5jJFzeM9fbebbKkAQMHcY1aPMKdr7z5XxBvWZTXn617nUZ3
G6DognN9HxV6O5jBZP5jU4qRReJ9u1HwTyRDGhsua2NaJkd3iu8eb9c2dWi9VGiP
hxbTo9iTHBew4/qWKA9e1M7L1bJqEHfoZxSOpRy02IsG11Gyiddjrjymo9PaLFFf
mK7Pz2FE6eJQGdmo+8RsjKILN6ecnYF4xU8FsY5gQ4/7TmaZ3T45zj3BDIkedacG
yDrz86BcR9XkWlLborYW5BVTG6kOyradIOVWERFLWc5XBRH7cE7MX0eL8t+HacmL
/GYgBbsJ7/BRJhYGBPp+Op5F7tlM3twjSHnCkYPoiXtN4/3LDqmTi8b2JN98wPz3
Snjn8GF6D5sbvvuCXMri3y5F5WXGX3Z1hS88u0QQ/J/0gIRzzdHcBTayPU05iFS6
t9NHHnGXqS14VzTW3sdIbci+7cUAtYS5Ccz44abj+3b6yW0mb98KRloLL2yWAFPg
wefUJssA9PSzh1ZM7M2dAPCWR2UsomhKzjMRGOWk0dWrZDIFVbGaf3m9kWFD/M28
Z20Qg3VdFOBkgbmJgls6Q5vzwFw4iAmrsWNiPT3j/uHustkcyhsGc9M90AAjHy5o
gFihdGy7Ym05yAAkDH2hR0Zu1rn7h3XYxSLKhwWAdPINyKz9/icgA5D+njJulEme
4ncDFvR74zxNDQk+5y184moFZAfqsdJtqKlzET+zHvSdLZQk6tQzwlW49sM/dTUo
knEX+n6jiM6Czuvms0JZqc2yZ4cFKko54drv1iIvhQSRRw4Ty0UtubIMJNu9J6/V
jIiiuSubbj6PG4G2+Thz1wMwGTYm7z0HUYsW7TSAXwNWbllJi+6F8YXrg++tuhE5
/x2rw0S2tfKui9MMq6w2gZPeQoUz1KsZwx03CYgpP5lIQYCh652PZNzEH1GyB+jd
0iZI28rPF+atL1ZDR3sgu4BXFz5G/CGvpIKxwq9AThWb1Qh85Gl11hO4sXQQcUMG
VLpZgI23HS4+q1TGDwpEVABLesEo7ckH3D0bteFuecXJLjLEh3PGhWwXR5fIMek1
SGpM0tGPl7lOOIjV8ItbYQxShoUACcBaaboZALBKIxHIUZeUGyk+Hm/tTH1kos+5
AKP9e5Aj7kQo/yZ8d0dE6mUEqSWThrFnxpd6J3ZYCgRdJ3M6Mq5moGo1+RIziJOF
TSKAmXbyNaAC3kPSRET0+6EXVYDiZq/Nxy1jo9d3cUlMIDYQ/hRsyLXi+Pr4S6uh
3dWCyYs71qjGuZ4nIsiPdWGq51b2vjvEF95lYZaHoPg9ujInqLNj60VVNyzdnWkD
KxSv3EHghv2HLve+A/ilrAbMFwK2S6Iyfkzw9M8IRIElQObZjYGct4HIunj37ezm
vYfCvR0AxXVfVTul9EZubu44mOXZIasHI9nAiCJ4/pHilBCMcXv/JctRnpGnhwf/
AfkLub0ukygyf1Al3NVzoKwgsec2Y5IFyhrmaA3f0RSuJXSbPUl0vvlS73eK1RNd
e3Td3SNxQ82qHHRgjOum/VDJeqND4RWZ6Y6CqFeqZeyKV0EZQWhrIBT//b1y7hsy
dQOpLXlTpBes99GOLs6CaJzofU736Wfap7IPl/mq0I/j9x68/CtuV6e7VxlfvJqV
2VnMkfV4FY1khNwhiPrF8kEghh1ELs8gZ2uVSFelfpoKI4qLAYCVEoG4LQq5rx6G
efvqqe1NmYHAb8lGAjP4ayXum68CH2+MJLP1JIIyfQ8C0+HI6dbxX3sQeiWmNDj4
34FopC6RMcqQKpD70ZsC3S/Yl6/TM8ZNfXItRjWoQHrukoMQWl4a4Ukf5ZE6AVRl
T3ARBfhXkWYi9B+tt2elz9b3ekoZfr8r8KH8NHYLJw6N93G6LilwZOFvFsPiv8VK
D0w/QNTd4LnCH5qKRwjOi6hGLchD0tfURj+RfL+iS6xnOhka+H0cHwswz3hdSlf3
Srr+dkIh2rtANM4ltXYm1/Ka0HrUHoNjOgIvRwSxnax+cBBn5F/zj7a/3sUeJowp
iwoFQcbJ+h3tDAplGkFrRtPJkecXyvwt5TyzFGlXFqYDDBAkCveU8RzLDbfFOSCW
Gvlw7RGnouQuoPROvds4UmNi8xVCzBhYyIr0AVOfLAfxRZpj7aMC7wDPKVPRNqU+
zOjsPK5V1N6HOjwfJuesfarPaqNAsY1rtgOcZ0BFiuoYjytLSn3UgP26kFycBVIp
kv3vtY44ykhO5yszKl/o2wGZutXikuZM6DtKaalTIXSnUZ9QgjMNi6rHEFtQ9mJ8
twPLxg2huqfdOL5TB1MddipF0F63K+WJacwzjnyNbcHToGfIm9bbNgg4s9+qVrkr
+6kTfV7h7Lp/IX6+GWofPNbi8bppmaIyB+1yw8VHB7JmQJqjdT/TlRAyzkdFWVr6
XEZIkuPwz9WrfLEndc54iBEZ8G4etSFbTqGHhPH9urblO+M37QtCzZGHvco0PL4f
iRrBHFP1mGQIH6Hk8i2fip5rYdRanWhq6h/yl9s9YKQbiGPglrmtM9QXrVoHWZzH
GArsxlHHucUunQ7qkeRVcRxcK1qOr3Ps1ddeLyyBw71CPCOxxuigVgiZl8J/35BW
gP9KSjowQwbmjzTxjy47A0XWIYdJjeWzXzwtQANwlhYRFqPKwJDAz4xUi8eBB6d+
UfEg+llmjAxtWmbex+PcFM+2jh+v8/34pL7jgrotRAuxyv5Q5X97SaF03xc1avsT
3C5DyynOskGk7sM0sxijXr0ANFUMugagjZ6ldHGI0JRK/63gh0Zq8ic7PMXq6MAp
jfDiTNThNV/Da1qWXbILEvNrxJu5SbAVjTEFiuBfitaBblt3ufdJSw1If3HOyFlW
AdKmAizWUgboKr9957Xe38S4IDYkgJFUgCjPGAgzaUSHYe2rTvqGX4KGLXEDsoyW
qu1I5qqQC07Cb4oV5Q08imCelDp5Nob+B5kRkSGs35S9JjnVkRUwWG62CfDOo8qc
jAtFk0kcSHxqIuH6L09B368GrKK0IXuBQ/sm31a99fTWSOTroaA3BGHvkLTeH3ip
fpAyIWwf+BbY+Lh1dq/MEuENs0wxdDBKqH9UJlx4yF0bu6tbEikOaG6fIFgx9lex
ZSEaxEolutJ0te9PwBFiVVypnAGQ5vSebheUzWtm2xTrM/kxUHymxeI9XGDA30z6
THuI1EqG+S28wNvKkY1qSOsICaMCNDhmn048datjkrdPybepG7I1SAcVo1Vt39sT
Ca7IyQqZH9yALE8EvLScf6X1oltQ29WK7F5OiZUzOPA1DxzeVkdCpR+daigXXYnn
K1MYiNu319Q7KIt6v4e1fbw/3CtJZmrIacQueAKMGrIHdPNjQ1khmrDam64Djvus
AjP0gRStHv+FGXzOF1o++RB+sMzczFo6fO1F/WFSMRv9iFmbTAzxkwSdwTNpfZDI
jVtEXYQyDx69NItY0NNNEnHfRnKK5PDhWVfUXjMYFOBFmhzTFUB5d53m5X9x72yA
EkX3LEMrtKZ12VJ1AAcntdmH6YK/nLbDv4wR3CaAWIdSOgp64LltQmCweujJ/u7J
7EszZPhnbeYHF78Uwrk5eHjWRh5FYvpwlqvW2WJs+ut34+zqzjOLUQFFXoDXhVt9
kr/FuV9KS+Iugx4KHXfzccxaOY7MDX6w/b4yuIkMGgjG3oT/Sbqpqo1ypGs5DbTi
/E17WwthjKN3TkPWBnqw/IR/kKaxtF7FuPr9K4HZAhdXrSHTcJoXWGbD7fZXemVw
FVrMySJJpDz4+W0JCmFOOcvUy4+rdsFASkDmyWUUk5YvPpCw5aJqKqaP5/PBIdUy
gxxvzmQ6UO2dHIL003XC6HsbX5TaS9bURaNdfDVYfOT22II98yChKF/Cl4xHStiM
Y0lWBxK682peFKg+tWcAhfaXqHlk3d4bvs/JkPhf2r5nbTOmOkLh8QAvXfQu0d38
ZJqL09fbsbhdAJUe3SMhXBRClaJzP1d30BTyeSg4CLaZiQ5jTyE1rLo7Pd+XCf1y
+XmCLyr7TvyFcMMtPD6jBC3SPL7gQLQH7+alKz1vsPKUVj1pN97Kn0jGQJ0h9Nvu
wLU8nYYfxl5MmQUpJh8Ouy8kT8mbRN2ChzwpZRWkiifIf9Bv9CjrzsAY6MjghEug
gOr66tJ0WSO12EdmSuv53A2wQF9S1eELajSAyKWqfio5zFgtGECnWohc1madeQBv
A3Lg9zdt65FnrIJYWxCPT4SbJds0pk7/OEXdiihqWlfe/I2BsecnckAk0u+2y8Fv
DjWql49pq2tK2DuQNcLdsZxiZoi4CrP6W43YmZY8Ita0HohYd4rMnIVE5GznL+cw
Ttm9AM/xAh0k0wrW7qEoTNZc1pug4/XSIJIGmbsmWAVrZKJWkQ03nNmls2AiE3+K
+exX1k2a3Pde0R2NQG3LHWoIyHDpJeOBJfSkj88agDNq2Htfsv4g++vw8C56yi29
iLGWLE3BvsNIh0mkydEEtOqZqrO1scDT58Hkt5IYHTgRR2q/djcN8i5l+bJriCBC
XA9itbn+VLuuLOpl/5lCGUXWA6BwnPFdTttPC7uNgNonIPT04afa7RRiLsBSXF4g
Vag4SygoB/hfjfHBlyFHHxXZjHYNyVgSTtAmfYUkjeDGMVzj07L1vCaveIEqZqVi
zkkc1I6vFKubBQ3eXfR3JU8d6xHNmbecDex9vDTRRvPF5z60Cnxc/7marUSQ9uVn
sDPywLRLFabYmYJKceJ6GtQAUoJuQi4wxp5Gp3gwEXqg2q5unP3oWtfiM6bvSTPu
sm3z0/DydWk+1VrnsWXj+Rb+FsvCfzVHQEdNvt1lRmunKY7RGJtVeCCcAyAgX0rn
7pEG9u+hKiAXjIgL+rMfG3N/BM/qrEgyWPew6WhzjpbT5PEPwAE9pmYDFWrsUKUu
RJn+PYzXGGiZz9PJ9TmODy2Rxq7w3NRyTChFL0aZ58VtW7k67VYR6msxtmjOJmLU
8YAbIIS61GqwR+A7K7Aa/sKGMMo6yWESqQ11TZ/HQc37faEtGL0S9xHevVsPln9R
tAKzFd/S8Y68KGrTeA0RtQbdzzz7rmDUHBQRy23rC11HQwXggu267rlQVmw+6bG6
yNvV0lmgSDsjyHa7SymtZYs7277kTIuGSuo4PJ4/EJCy5hjmStdf7nC8Kie58Wrb
eyzpB+CbqyH3kivsb5wGCBSn7MeuG4jlIVBOKfZVzQ9+oN770WAlNMrO02Y+xIlR
mnrFlTnAAkIB30Y5pnfP1DT4miJpacmbybOvcnGplfIBgPh1iWEfM6y7xo9z78dB
ehqm1Yxbg/nRJ21hWOOrpUdAlz/it9blK267aCVEbx5tIckS6QHE98tjWSVmnLS0
1Eh8tFkis3dGQn3yZZpB+XJnDZsYt2rhQJAk/Aaxb/zlKxHcUJxQ+kFXbzrXVQI0
T0y+oJlHZROE+NVYKERxjdtElUB2zVwV9petO6USEDiooEpslLnPhkjV52HZjI3H
jmEsz3MLSu+mQ0hfLUP3U1LItPbWUw1pc58JC9irbk1x6RcjqFBBWdiMEx1kpplh
cdWBLFR6Eh3EAjpELb8OH8Kfp4jwQqsOioGkuyZGJwe9IQW4wddKWR7WzJjyfnTo
OWPPutw8xnoYK59v1msBlUM5AUpgzVqqsWb9aHjiQKxY6scUI9kJPyxoDtx/9ApJ
UmuXTy9sVOr7kUf/UxHdUlBCjC0z6w1SJDGvIl+ni/kwqME8augABs3Sct3rBFyc
KqaAs85ls8cIliWcr4Ll/UbiP2PBWuqqj10OpLGfcGwkhUq9parJyFPxALh9TM5d
C9Q2O8RtKE/9lZASTg6ZtStEoavL1FkkuCwlzCQcp+urCEKQCABFfRdJSb2DE/ax
i6Yb8bUIO4NaPlL2l4UONBWDwlEPBEP08WD/RUWEG+NMdcCM0SvO2AiKiPejFrqf
sf2mOjXqZFi/CGDAWuvTXO2qiXF0P6323ZlPafDa/w7oMmTzBkfhTWjmKuvCeg2c
5BJbhPID6tD8nFGntkl6J5t0BT/H7SMKJiDAbE8iBapFNaqtH00CVQEO5qqic9YE
9khr7d3LDAR+jGyliW2bSdQJwjIGgnsLpexA7jKa9UabzpVdroQtD+6aWGZoN79s
Z3E5+WmwH64CMKz7NrY0tFCZpY1CLkydLw8SoFMDvMAG3A/Dl5ahmI5u//OXvQur
Na/y3NaFTOSB3hFfmJdZL59M+ME+k0osHbeLsq42dB3WVRZ6Hg0xtT3LZaUx7aLk
B0k98C3huMqiknAWm1Urqa3hjTzRRWOJ/ux6CgSP1E5yKfBf3RqCRnzuwCZqCdrQ
0XVI3bnapCJaYeRe/bN5+3y2DfyrFtc35D+/GCR4+eHPgJ2guVpOcxojDAfWc9U2
tCMU56SGGVEjgUs4cQpB6b6CBzgB8EUCC3CvEyP2VjLTe/dhtB9WZRvzDklBj5J+
lkwu84z5vpH/eNFMLxgyEzPxTtMZj5ymMGJNziSfGFnMp8Sfcy3s+pTSerODciyx
+19LVPfW2n1pYlNr0hoVDtpQU5M+3TzipOlZ2iIKUVwRw0BQYtUztBsEJJ2n1raZ
XWOKtAQHYBWM+4z6M1mrU0Y+TIC+/inZzSG7LMMFv+B9rqWGNu7Tdl3B9jW3EzYF
9PwJwy8h3VPpebwHeS6XsNoyoddboKBaCwBZBaIf8mHSOzEuV/QGyZ21Oy72GXMI
/054PeOAiswCwVMAbfBOt8cZNU7fMfdAz9BkDh8ZDVUhOeGYleasjSzVL0KHVmfN
LXBHX8XoIbIR4zHYO9Ln75chJmOqeWNdq4j9z+K81EN5pm3pM5VETiuYrtTf6U4S
oLBa3a70pTxhEd8Jb4Zv5Bb9HnLnMMN30+rzUQdI+8XN+Y2Nfbl2jTz2mIAtzIPG
hRqUanLeR2sN8PTNiuGI2gbOXCikWR+MSvdjWn9O67uO2oo9St0wetUB/mHwtWt4
UWyFd+AbEtq9+UHZ8Nh8kgGYyNckxBVp1CPj4dcTuZEXjR2QoUymIHD/EcXq1OZM
IbEwyxUB3duxGpVypOHd83HIm9iSsgpFOpom3FZ+8ND+oxjwhlGxP2/EGFkVD0fO
gNqfGRktBJ+sdCdgWgrMxoLz7i6B7HBi9sL+MJ/IUXoslj4aHoH7XNzVHOYhcre7
LZ/jEpKsocgzEpWcnKEdpfGU3+UcJJm1sQsvK6pC0M3O5SwOJ8G6jjMHK8wRYBYR
tGDm+BHa6w2eVk7skgsotoxqZy9246DvGN39iodUL4cO5phcgc7AeiRsIs5zuTYL
EPdHfT1cLy/hTmWWVeDbP9t7OJij7C+kSbQUfBHXubSXFsZ1GeiyDz8xkykO3MaN
DWhw+vNx+fCu5YyHOuVVZ5emd8nJf/KLPeyh0UZT+YmfAvpQInc1/6VYtW1xiooh
FXgFl3H/6dv0CBCmM/UnXr/jZmnjsreiBFB7X5P5DICnuGMgCZL7jphoWFdrmyu0
Diab/dJR5CKXMrLbdz1zEek9loUO+3h01xBJRCCZKO46onH2Qz8CHVIcx8rR1KJH
ZjNJFColqvZbMggs5lnNBsk5TstnY1RgItD+7idOrta5ggzs4dOAw+WzjdtkfMKR
xzI2dj73uCRybnInBC+kwKFTzOEPOFr8l89rKMOseBI6Gel0Uztv9hsnzsLZu4tV
uuj8g+3XiRzzw43gxaYen0rGkFv5b+AdbRT/KPoVtwVcbWEBtutN1jp17oGv1mT5
iBMBAvkGxoQ1mPEueiqiMLEwoLIhKOgaPvj6HorpN8NpfhZb9eco4ZjD08yFigK7
1UH/1HRFrIXc5njZyvCzhwV7SNbrDDBUz4VGbqwCXepFeJmsfIspujFrcC+DjrJf
XPwEoHqD8lCw2IlZSxrOncfvJ+LQ4K5lnziYhGmXLzHrVgDN5vcQdO/yyH/yHSCx
Ag7pUtOO6iPAjKoVL1PH4YJgfSITBifAXLCUI4WK+mkgTmlek+kxKTQGndoVVilt
aFqns2CjQFR/dpZRnuM5H6HoAx3dRwK6WaGB6DziOvRBkBiYZhTP+Yrgg31wOE2K
7Ejk58OpQqftAiySIpNiTSUx7LKTrV5ngCINtoKXsBYT+vhi5xRLRezYrZDgWQjj
Hvu1NSRUHYtoqsAYMwRNXHFV8t7iok+o4PrSw2FjbWzDH2JFkJIymH1ZxEk2T6R1
WgLQAvVAwMWly5UPg6oqmdXQpS+wX2AtvZVrlxFHewyHlIHHTa9u1l+LkTyAao7X
TLmM/+cIovxHDKYQ/SxZZaWwI4SbKjaKA392TFEWpMJzBOVmkqxSvtvjami7Iclo
vj6u4xAOt72lMEPz2b+2nvsXuXTNbYxtluYsLpTD90x2BN2KMNmtYyhZaz0+7O1c
nH2aky3q0ImP3Jwax1MmLvwIIL6lXwv5ZrWNnmtRPQXALb3Lb+W/7JdOzHXs8LO/
k4IUwJxnAcxDGaA2scGtXQGA99HQuxwClc4CBJiYzMo1N6NPfY7nK8DCX6DYDmOS
MorvSxGqpCzz672aHbbqFXyBGLSVVisqIpjThh03PvmwFBMiV1gj/F1Z+pXSCSEF
DM9gGCXj5kb/oWvRecCWS8BDJo++67xWer8ds6Y3H5+H1OA+PvcsHulCKn1oHc+j
VieDvZzeiIbhBa3j8LXa15hcQnlmNDhikWU7BzJpjVjMaSG9n2qtcwAMVdaRvpo5
ivd8KgWNkYgnesV2qre2I6BI+gJZrhnNhsEo7X8oU4cIiJlGhhZ4yYvEVaaHXxkO
I7+5LHS4OUjY9xIZvx3bnm7zIMAf6e6XALupzplSmwFSEPAEymSdEF75mf0LR8IB
9V7q+Zm+w6/yFMPg6AHdztoMH57Okc/CMYUJC4Wk0tBH6LjwfNWse4WLTIfuoLGv
urZh7nzJzwqa1P+cKXIRibzjEHF4jsofOvUSRU1KcmRNcgKRvczvtFvkBJ/h68tZ
I4S7xPvxG+N7HQkC6K+Gy3h1EbijcIH7C2UjSD+8iW9ZTVHgo7Vc6OzDrUTc+ySG
OKaFTRBqja6rQEEhZrvcuEMdZ1Ru026t1Vwss/j4HtZRdgrRk6zglU+RsGxXr9JS
CtN0o/7k4ZKHVJRn3kw6FzRavJrOYZGHZZPKWcQ0ZT5Vl2wwP6YxqB+C2fjLn7Ri
LcT1MvPD3Ri1AHpCvxO/v12MrxwZn3gAIXOAm3JN7ES8B4+Qe6VcZkOLiXpF8JuT
84OCKy2u4qrFHxxTOqOUv4HGsd7sWDVxxVT2z0Wo5VhP4EeYcD7JgAGAl3OF5u4g
PpadsvcPaptbyau3s/3mNrHqu9DCdxFhajafMteOmP4NoHLUgXN+AW6LVUs4gN5W
enI8VNboPiwouc3PTzUR3vP2hKYD+tw7NSOFDu/8y4Ryn3VwihLSSwRBWOwpKjat
1/0BRgaku/v1pH5gAUjhh1ozVO9gNjOlpODwcVMkkHY/j6A5apuFvt2ryWX2nwzg
MH0UypF7q97sU4XKxRnhCKGRO+dN7rpGcfmZf0MGfMYhztJBt2gVinsxHdrlxwIy
tQd/DdsUMyISs0CKNQYXkd+BpnnWGeN3+kJ8iQ615oyA6aatdcQuepIreZj0MRKb
MBS0GrnwnWdIfcjpyGxWi3H4nWyqDBbn+jsXE9vBFJfzEUVplzWFPhYlFZK1Qlhy
0s4ztPIC1fua9lSdq4HXOskew52qPl0IzDQ7/jwaEEyT08xvCmjKR7Z/q88KaXsi
1WXFxZbENqDV9xPWzhN6Xn+v2chcWngsDxApaU9PQc43t5l2j01p5S20qPKH1idx
7Zi4jXb9eAhy8e0Ww3pAGSxBVDIPbcs0eLfZQOcijvQbqkxk0GTsZgvFDD40uatp
avsLfhx9xGRIvMY6y/Qc1zqc7sfbqS8CbDMzK6GlgL3Q/RvbUikD0w3533fbNqd5
kaSoWKtsaKsRBvIld5XHLtEH7XbNJfZSdyz0SMlqYkc9BrK9pfZOPwWxdei64Vcb
QJiI2gWsH/sB/P9Rm9ZCz3LLdLdwnJ7YBtFkOeIF0u+pqOVfCcsdPn2ipUdzBClo
yJs6/Q5EcwzQYfC57gWPvrnC2R83K4n9b8i61ZXeZiqpkdomg/+6evuBQ6GcMb3F
V9G2NEzuG5acPKF4GwXoZhCLdT0+ISH/iKJGNavDLdq3iTfrnFZU5r9N+Ab8GbwL
STO5vfH0G1/vaGRKhna2uerukk31MEzX7p3MBaeZP1JVHlGMzO9Xcc/4HNmeA8Q3
rj4WEr6dJ2y40jQ80kIcXb/Mrv1hVGUZez/fFgSPfLE4kGpsTpRCxfMAChulBkl3
OU5k2io4oFObA0Y4QZplPXIomdsxEprcYpnaRY2WhhU3O1uDHcAR2kI+YpJAb/Mf
3oolrQnnq5MXsgmvTSpxd9ZmmogWiMJaFjyYSdb7RAUADL0R/l3eXtWWgGutQHnV
3GOreNsssuHxsQ7enYvk7apIGqa/79RGqDYMbgDSdaSVcDbWnJNcbEIkz+/L8BXt
DkHPmTdJkQkWsq4Q9Q3tfi5S/Togty7a/y0EuykJu48u+xtW4Be5y4fNqLr9f92g
XcdtBwwUePppAI/L1FwRWwqPZl5C2dKzqQTnRg3+u6mrCUpKhd4U0t4ZIqYTR4OM
7c75V0hWNvKxSy+5rtuuZcm2hfVx6KLkmKtKWW20gQRryBIaJpvRsaHKTl3DxyRd
gro87wUYRcNU4qff7vOxF+jbyrQfa7XKXeO65H+26EQGZygfLoNrV0aFyJSMKYcJ
QhBX7ZY+db5RCFYQv5NW8fWEbWe0wJkK5ARWNxKtpDvbwztgaJ3ETMCz2zI0ox3X
9N7l/vY1TrMbOcIgzlrRjQMqH2gnX053xlorzHDJ7Hd7K91ENIGpTJSQkLL2KRWJ
CktDsLmA2hcK3h4I9N0H8JuRXP2CLWBbAoCRvcP5A5pht8eyUvS61BTRxBge3Yr+
aB7IN/ZRZvWU0UN4lTOj3DQp5AWGIEIcA3cShYtGCS/eDnlT12mWZGJQJcEf6Nnh
O2/IbsYAq1aP7hMhFDDvBm2lVhDKStDqvFNa3/T3uCfP8FTvPKpPDnUnfkiQyTGj
q/eR0ZekwI3aJ/1BBFYkRPmhuOmhfFPmK5cz2Gvm7nn5HgpJ2HSx/3TIT5XjV3g+
o3lcXihzdVj67LqynBxpecZmGFscrTVnvoswJgqzonL8R5xKYPny96NlP9L/DuMa
/dT5w27kRonsF/l41YdmH1rhDl4eDDmpCugh2DtobvqBH9UD5driKEeqKrCC6rwp
41TGhV9iENNL79og4RK7K8PV0z1reCEAht2zsm8o5w027ahFz5Rcg8ST8YZCNqjH
gKcpmbxo2QyS9y2qFt5QuNKYbf9em/qybCJwTVzzlXYSPAnOP0ib0Eb6Zlfd7D6s
NMGqMFryOx0BJMSL5iYu13Kqw5Pr20pMzDKBN0GdtprF7CLOU5hLA6jeT/7SAjho
PSg6b6K0gzYL8UBFf5y+4WFsHUYLQY/iZWPtzXsTev34p2fFSBGNOpE/If/wDoMF
W93RuMvTrtNxGx9cUhC1xlWoqHU9tJ8ikDjDTihgN3/Eg4C09ePKTWBvHnQRprnf
yYWTPHgAkfNUamzNsnl6z+H0vYk+8UCfRyPtMNK+gz/qM6VAwmuAuyyuUrFB19nG
dgdQxppmiI+6D+5pH1MsFV8J4tKkMQZFoOBhnAJUp8QvK+ugfGkeG0W4Wkl2Wz6w
7aVyz238QqWn+NXtprL5WyvsKlToV6mnyGOCgQZ0Z8plYGckOFbi1XwbwbS/+pYA
2X4beMIgPoPSSLE9e2ZGNQowQgX/fq7+HJQqpoufycj0bHSU2ocfaTDTNQdh2nC1
M8v8uYhGmlLKPVtW9J0Rc7Ubqm6LoqJ/foIxxo+W4R5/CQxsZMC+QKkXCBRPlD81
tR4FgM7pR3Uf88aDV9+GGDqjbnBVA+Z+Jg6c702pRTFun1dpYcLkYpvbY5F1AR/5
tSh6ULaXUweYlxVXzhS3JtvNbfSwG/4r3ZyfGBTzn1T0ghXRbzqdkrQZoSS53MZg
gYV7Wq0Nhd3cqsz25YNy6snbxprQbRb2qkKuZGz0nVMX0V5AHGtKFlk9xFfiIoO8
0ZaVfnHpbrhtjk4tLR/HJPxAd+g5BGNb06sEbCL+grlPJH6XQUeUrYSIrXYJk3FE
Y06F9P9c1EWKZzffPUEvKGVftPMHtAPyaU0EV6Op4RY83TcCons00beByY65b7kp
HHgetHh03GKxhw10aENxxeGCSQjfViOH4xq3joyDjW+aQI7JQ1/jEHWdDwB8QNQS
4v34blod20TLEEM8DzJQRhGJXUfUun6+4WmEl7kRFn+XN6r0aPooE8fRVDS8cJ/D
YrNolCKm2ZMiGriMGq/fcFkwpSj7kiYGSJrZvnDWKMkn+pplCAPlDHPAoxTZxXBI
5j9FXdykg7Iw9ToR5QMofIUZ42rP2gjSf/6mw8B3BBQ9Wj5fGxYrBnTDQyb1qe2e
LIsNMrndZVKdPskRP1JJWVryzzFN0UlMLXushiveNBCZNfDtQhnZtrzI6WSkPpSJ
LqXnlzbm9VC8LkLH8FbL2Pd7UscTdoLH4Bro9MnSEtaFEGsNbuHo3qcgEAZTdGjS
0OIaieOa2KBapfQX9KsnXWLO65HLRWk4JPeQjUQ9FEvuFyWcEUu3ncx/EcM7Di5T
Qu5a1M2/1U58R6vR1WG5gBSHsV8SmAFS9qxZ4D+8ZdrX2ApuvAZp6kLbs1ynxEf0
bzfqNccHsVa+RdpUznOGxwwdPw85sV9iuj8hrc4YcdQchGJxe9KSuJOqJ0sM7Ui4
zpOcfk414kpyUrOR47K5gqoYtKqTaNGiau8hc7KE25QVSIVXPaFUQBjYkf8KotPv
4iHCya8S0ACr30ZgXqyulXR8x7Am1vn8aqiPpKFm9XYqQg/Q3/oQUZl6ms/PW42+
+iGHcHsVSd6JFC0/Ga/T1B4BZkO+HtUMm3LG/X5d00uT1dL1+YC6cjCYKCm3pfqI
syqfuajo+VjPgSHs0y6THeY1rfDoAsonEXRNZZ7hR3c9OAdkbVKEMUe9FTJVqyfs
a7Ucphw5LHr/zr5uVLtZME+ZO3QIcfjql/4a6znqG3LioxSxlHwIeOX1pUVIGdyZ
3OUvpBo7ERuQ3mZLWiRd7bo4DJPELsqwdjqvPRcf1h+8UhfzGsQ/PzrSLaG2vYMu
kpZmiJ3HVko1BMFiy4F/oVGQTaoOBKGKp6a+oDAAzBQ6V8EiU7f5TFt1/vGfNeBP
UDJoK19Immt6ncEY2UbFx7sFxlQKa6BmwAnHIUB9/ZXy1xz2e+Mis65PFTMeDPBA
ur+5NaHggjg2/ZgRvOK3XgFQc7vYChtzVXZTvAC8c3xa5F/THnNDZXt/rVTUlSeS
LmaPplxhkxfVltuWt07f9KTxyTMSEHo3XaT17uYC0QsQSuLjaw2E1hmotSPte9vE
D1a4xj+RUZgOsOVsz7UjgmpBUids4NTthyn061ODgMCOgM8pfN5iJ3Ik+/rhGAvu
TBexLAFIrXCRVLJ0ClQfnphLdIqUgU3mylKesGI5+6O7dsis05AdJz8lFARweQaB
DLCikoeCItBz8SoK/k5aCHM33Hu7gJoddx2k00aDBW5e2+Iqpnq6ATzJ7+2/6IQt
JHx15b/1pCQ9/lGvYVma4rEyYhIs19huygb5z6t7AEVGn2ahSASSobG7H8UbZebN
cTs3PTxlsOKshPb+a4kts1FCKmewK03iApljqwkidGuqgPCf7gsVjrOWa90kWo0u
8EuQd6Gh2aeCwxy+QM/jGwRxHqdBolZ4woDSxZ/f2irkvBpGdRDm1vViln9+GfAG
8Bm+PXdI7J6HDJKGBQz6E1yPh+9x6T9nVQiF6kIbIRQeVFg/dDOajXLWEtfozNyw
AeYv+ehU7dGX/3E+MHu0P9yfIK8q9bHHzFQ2E0UHTvqxkGOs0aDi4NVNiJcDABou
zXdPx1YWggSE5NWiVbJL2Wp2rJxEJPYl0dAb5bUaSg4JC8eOweKd0RLyQzanHdkK
yG+koyZSY4NAuFjMwE9W5+TRueEnyX+UPLG/28a7S6qbNn2PxppUgjMB424nbax3
to2s00vD0ClAh3dbdtmJDNc1kK3fzTco8FY5I5bC/4FjFados39NPCM6QzBYTCCo
5xl5dOPIMccAsvFSNX5hFMH+icW0d7IFZ3G2252rKwO6JtHdwIubduuUH0+Ye9L1
1/ZkyrUcI/WWigelzXl4uNbRMRbiuX0V/4ngAtNHCnxtrzdXO8cXUmZaLNbnYRHm
b7Chg7EJe0VAfKOyBrQeGWMJ7fnEOk4s0laM615X6n4fem/FR4qdaoNh4q7r036n
IDdpqZ7JD0zl5xh60A10cH5HDZSDlls4bK8AN05RQMUWfT9FDmOTADNyBXiRY2nj
rqiB3rNuJUr35W610m4XvevSyxtdZca6tu3cm24lK2lPSluiVlcl70hz6rFFQT2X
0ZsyabMlxlqooX/Q0Zh7vX00HKDUaXFrOaLWWPALV+Nmk4g/McHzjmIsLk5RRvRW
bBv3sF0bdj8sXJKYtmzNmanSKRdhYtlEQWtxUkPVyqc7madQENho2krtR8jPpUk9
NEB3somg5gNP+LQf+ZOyoguqvZt0AZyRe2d19J+jtvf/qSRiSkynqalwZQarnSj9
wi5edMFtSYfAmeYi+cgp0N/LSxSPv6CoJcDs+ttnVWLNB7Vth5oYELApxY1/XQSB
eAy0Pm7IMPJ/I9MQnz6szR3xZUQxA8ORTVtDx/DsiMPlDhB3dBLOXKYm3MO4CFyB
nOt9dfYD6WndqJtMCrgd/2b8GLAhv5Au1yDqy5LAEp3q1mMSodFLMxY8SqAA2AWG
gtNp0iaLMSM98gw4hUpttOC7V4F6+tz1R+pn9DzsabR9sNB5xIflkycMtfbZJQY9
467ji4rJyrcUUl8ZUysCTVM5VgEC17x+QPZUfm2/nzH5QQD41J5pjMEPZVGrRMHu
jakMfMeKLxhYymeKmvXpRsgjUFgEiNNhihwklqP8f0YbmNkBRXFgWP+xe1m4i8qz
nlMjhRYqS2QCx2lcY8lYwUn6LKXOd49WH+7YCm0/si6D3PNDK5VWqHFdokTCgyeD
BlIWl5GtJtkvYXjk2RkfAFbTssGW33pO9WfrN4KOGDn7icVJQTeDA81ja9eU1y/7
NUz5YRg/sFMP3FW1y1ye0TZsc7k84pzRPcwq8bslMxLDO8HEHIdebAS47DE4YHB4
xEjEva0BHWi7bjvxV9PJqU45IyKGfT72dnuHe1XzC0w8NZf3RAMbPkQa0hQofO/q
jyfLJSRiK3uj6FxHEoPmv6Gt3BTNOgGCVuQDcNlu7OTeS85qwGlVxD5R2xRtRs0q
/Sfu5UCD63ukYjhhoGa+EKqYycEI15zsTB43txnEa06sV/NR38HF21sI1Bh7h3od
UMMH+TcXGbSicsYnM4Gl9FqMV9QJkOr5A0tV7Us0lgR5cd3I1Lfaw5iDGij7uO28
dXQ0u1c+s2AAEQhhSxqNm/V8s95oTQc5ba+nsUpG9NLrW80aQhRSkZTVGolOk8xb
nzFERyKiDBTlCjmSluCJBr3c15m7zIdHh/hFUSAb13zRufNCsvtUyOx5ZYUKbk7B
Ei4KTWSep/gYRglWf0E5WLf9eR5a9mZKIHgmsJBV/hwKf0HtXfR5oClLkN/Ttcc3
gNJN3YgqXhE9g91+Q3tSMLQMcv5DQnIM6HJRKd2Gpn/+f7lDAVutFwosMdW3Q9Ll
JW89kqoXGofgiWnvRWa0JARLa0x8K8n45cbjgMCytMKlqbHXuYIumKpqpZB1LOkF
nMUZqPzcBj3HSOLNAoFicaPAFqhs45sZ8lcNv0B+x6jdhJPK7zybZibSFrEbiy2G
qUFajkLLAQPXwnFAG4lJTvx8AJfjq+2NQ/UElBL0Igbe6d+f4zk8ronG5kC9Y3JL
jvAewu2SGCuuuWCoZ+6ZCCmDWsFllhRZP8kmKwNTMn1XPBiO/7PnQDEw8J5z0Ytk
Bqfk7btD8rfTSKsCbIZc55xVB59Sj1XKobGcUJn4y9jTUKicEMwSfzkGRXzB90kp
SrKlXT3dzj0p7xMfoDe6RgUHeavFoMi3plVj9ad2Ucx80Ll+fhqwYdqxjWWg9hz/
Qd4j8Hj+V8qmsIx8qNZQZ1L/1zqC68n3dyJzn243CR8ztYBYvYt1oeKC2+Yp54JW
gqlK8QILC8vGd8oVywToHFUcazmbRFKv4fnrS7xs8cJWV/y/IN/hGT1N3jti3MQN
hXipwuQpZwJywoDwl0k7jAXYZa44TeyR5TaJDcpNe1gamDltkPephYmds7il8ieq
McEURRQIFGO0//jtCybWInuLqWPrnQ2vUgwn3Jn94SyxUNGnxoBtHu4e08loMHR1
8Defi/y0cgawQa/ubYaaTueYtnBuMcR47cRg3iVJ01wDcoJ+2Ynq9KILwVA7y/zc
YZ5JJWUB1TUNLE9n5nmIQC9GTtOR0xDPF98hktE0hXUG5RTO0L9tVHaVxIWBKD60
ZfrnsxAJFln00C6HAOKbM6xR6h2u0ZFv8BDSmvKVn6M/HDOmStM6f+ykQXR/VFVP
FNx+m/XvF1VUQ5LfmG3Au/9PxLONLeKCUMi7XMOnnEMx7o+r/Z7VNMNWn4dxl5Ah
pcmCREOaNO62SkblK6SRqTLTJFiTzGlO4PLEl6kNLjOMsUJeS8HZJbLjXV6rCU3g
Y2QsuIHha3IvwLzFYJjfOg/7ImtzNJAzkSEm9sT9xGKr8U09cd2mgB0lGflzVrVc
FXypgA8TJjk7E+t+AAtSIdwJ+JFNo9g9nJspuVO3JSeSRmsNnvqtHoQj3uZb1y0J
HMYl+Euw2mwRjwbWuHHX3HTmWlgOhdHODJiH1vQ3FPngM905IhJhZuP/qwLpIOlg
AVcuIKQuRXlU1YWAZCrLYBwhxsqgoZJc/l3TtYUCizQski6W1mrwQPSPyJ9cfdhs
ozZV2BflRlyUfE6sXJZv2Oo8bGRhVZXVcpAnF7JK3dtpPnyDxgZApcKcPEFl3xc8
hJRkmvSpbm31xewP08VxjzjddGWP5nXoacDWe3fV45hSxT31dCEfQ5G2zawaQGRM
ja9EN3wh52FpqIML2WLLU8eeiE/ZcMOoQJtymCYk9QRNpHRuMqpvgXW6waZGE2cF
HzYz1sJ1S0lmfLKNkf+osfuEXI60AvOHGMbkmkQZ6778ZtnPAFHzMuax56mZRJ5f
SDyN64/VXP6AF3jOTVF4tBE2ViU+O8XUu29nQM88ItK0CZanr3tGLy2Wm2CGAKY2
TKsIT23NY4DUH2XqsugVxRGSjyEc8jpxvAwuK/y4V1m8yKTUfji7jfhTn002Tc8u
4qeRr5WxAikMO0nxy8bqsXGLlyqmngzVatBnHlnJ9kpcdbZhJeJXsO0eI12FLD4F
mb3z6HpDNp4WsVPpjNuFbRc3BO5LLFVgYS/4mAIbcuYladhc8VEWBNiUzK7J56Yn
tDdAMNwE7x7wEnX3bFrBoK4NLD0VeBtSY9LXpW9KBOuPDUcI3ZbE5nz8QklFFnyL
+EL2DmrUNRyMevH/SnzFXBDpD1bkGNnruHmbZRSXJ+s/ouHkvCCbiENho3xDENOm
EM6bELW7pdYAQiuJuYhYlMs335yQwxD3tS1jEpReHqHxieffrjo+BAS5APvE2UtS
OM4ZCD/55bZF5QCuPQY/FrI0zo3YK7byjPOGMJEgFFvGdDLLEPTupZTvC/SE6OiV
fTGjo/NvmOhthLbNXyvWe726PUfXNeqUTfZv1c9eAAdWuTlHk/pecxkCX7QICBbi
iRHJU8Ezohg6xrKaMvhsQ+iEiCwCFOQ3tVYa7PcHDR87UbzGd3QaJ9UcdyrKY6+g
rhalibmCaMlyIeIvMgwtZlAC9Zn8zJP5y6nWjIADVXAlim/g2etMyv9SPRcojEI5
bZJbbUjYM/667RtViVqSndgHnIlujcP0F8L3WMV9GIwEglaieyW7+unWORincv3L
4JxCXVmtQ+TYfyJJKJAo2TNPi26zGNoJwd92cH2WcyxXRa5PVFhC9i4NIKfXKIpf
PGBFh8tb3JlGPQJLf1fLzRdkrarTjCnWc1k00qjseKYAiUFzXMmhpm9ACiAlXaIj
i9EkjpBgrDzYo6jLMRsAudDiSwg5VYLkX3kGs5KC6BQHHmCdQ7bYcvEjR1C8qxeW
S9nZeBdh5e9vvUm47X+/rfu8KHudSGG2ZsPwMCsoeXX0d1pzowiFFxV6aYxBIzi4
o7wXjdquGOhNePKS02Ko/ySikdg7ll8jMNHmpDCEOEkg1sPvUBET4tA/MZinV0i9
dkV72aHRKXCun1Cmq28+En9X4T5uMGjzhT2o9YS8ZKX5INy27TGUj4sTdELmcFyz
FB5FIxRGmWp71W5qKlZqim+YDInW+QgtZw4zm81ypW291BoGxbRNpa8deMU+EzwW
lN6+CfWZEi9OVyJYZHfdQ1oZRIXGnp2fqkk0n2k6mSipoqSjHADK93xMWIAhy2DP
Zhv63jUufilI82HyJtkXyCu5P8+aDFzpHahaHC+EiiG8W90bVkcDm4h184b23E2r
aCCUDs0xcPsjQnQY3PX3a25c7MaMhNIRFc/po/bPEoN5oxBUD/MidX6CldllAYZ3
VAZ78jjDUG3VSOP3qr8E3EK+kMnfbe4azl7uoWxMrw7JoDapGY4sz4VDfruEErHV
OEvi7oCxJzdMNbeA+mChOcz8GbhcTqJ94L4iYQumUE6HXlqXmPgiqQ5YOomxQ1R6
+ZSYxbsTBrjXFZJoxvJKjun/eQrbTb2Yr/l5ADbkyp6RFoMJvwCkZESCrlzX38tR
FAcVEN539YwUw6dFyPbsMFpVAB/uuQxC5OZJBy0AxhF5cFOdOpK9WJU0LP2FFeNT
/LzChhmOx2uGE743evuf80eIQa+PA7ckHH945FHThrwu0l2KmhpYQu0b4vw/tflX
k+dPF5+J4oofdApfXHmoeFXGqinmUC+zl2G4YJE3TCRBCXA8Uc6A0jmWX3YR4QcH
dySN4NSoB14QCkMLresaBZUhBi8x3hOdudcZWb7yW17XhqC2mIcjLx/OnL1qxy9e
HUELE3/Yp+k5HtbJ1UHe9iluLhnFbsq4kqD+YkkJbpMPT0g0puT3QVh73J6oDZkk
U9cmsZF+uwgjc3w8kf7QtXys37baf3gBsbGVl0qyP6mox1w8hRKhMGYCopOgeXZ4
A1b5rmZh6FBg+a9e824c8eV4LAL7FCKxleQheaBjJYqjp+EQj4H8eIqqPDcT/uop
2XkpdQyO8QLmiq6hpbGVp46WiEUvK4IQbhLv2EnFZwOG2Qq0PJytmjkvvHCYr1IG
KpvML6en9D6PsvIDlYvmhKyHLGyqS5qghOheD0lLN00anrCAVT9Lc6W46jZlY/+z
Ii6vvc2e1wmp60XsXGdjTb8bGPTUyOfMS6GCY7TJ8LREz4zjJBjauqGpX2lJXMPz
sUoMlzRgK5kSjtydWJu+Y0Qo3RCoj+2PxgmoDkhcFW/VJjh/peZQR4++LTMxz2E/
/XJrtFz9KvGx/zoyugQUfdbVlbRSsBRH2vDwoQ6UsGWhNSLYTwyvqiRttu6kL87p
bzKCbM9woeBtwJDPuXwLuqXelVk8NBfw3VUvjDxKboQ3HV6RgxpbtsM2JC+LO+Wb
qv8NhNYwofjg1peGgpqS3maVSApLmsRbVOt6ypfTVrs1T8AA/B4LzNNdeT/3abkg
ZPmr4FVJdo4I97WjQ2FdX3NPcpvmDRpHPYB50X8D+Lv/HGXFkwXZSvPy/sn4xIEv
z0sab1/2Qydj9kbQAC8h5pXPkMGZ4yg+jJG44vpjKuswtihckZThJ1h7oW8k7Q99
1Jv6xrRCqGuAnXFHx4VWwVS57TZB7WuqUpFjicZLNiDylkV4V5AherViBy5wZj7R
qOr3lRESDjvsYdrumd0sWJYEtvbtwWVnWVfDsqSKN+Y8mQiWsABhD7DgS5JNDZ1R
uZkDaJzFn7hOnBAc5hBP6aoLaFIvdCfBbvbeEq1XVARE9+phIfG1+fiw+gSzsF08
5JjyfQElTOQjfsnCiQ9KR5KNviwlr52yDlz5W8A5sbWv5Y1Y7RdIVqiITRBFBrrl
tE8GkOSz9jAZTyGYEu5EYmfbd+nQSoTz00ks1pHG/bN8dDmd5iRZtYt/zAidmWPX
aW9GxZZ9OigLHdXNtinRtJmAd+gYyhwckxC1MwiwiO3az8vj8hL63ndrTR4DlzSM
ILbRO4yxT54y2GUCWnYWdmroeZOV3fOxopZww+dFfU3ZnJPTWhu7zzSW9inMlO5l
jO759zAY4ioWFN/BRyiyB47socris5rrkm9x7Uq5nv4O9UCuifRAWmu/jfr8pERP
TdbaoQwnStsM6rdlUzdFZssJ73qi3aD9Te3aaDQR2SWA5OgKj4r+MlTcMpOFAs+C
yVQVj2a4Fc33hUru12wD6PIPXIqfZ4/BOq5Vc75QJw6feLSY0qGxneEFYcVYO/z+
NJd5amaM5a37zVo93+GwkcUAz8RcyS1Gv0Cvbze+M8uP+r6+FIpsV1q2eSs1j7YN
nYYIiigtSO46NQ0msFRXi5A3zI46xxCV/cXulUCBqDbvVjFa6YTxfP0tLOeNPlfo
akBRDT/EzfZ+o71LVFT/dFe+cvVybTY64uNT82O+eJrBklMi7RyK0eLjsIvmsC4K
ki8xJxEL+wtzOgtJahyms+BMrMp3rQ+aQfjV9QDaM0H0sx/1KnqejNLCQd8cuTBJ
z1HvG9tqVsf6X0GQS4ORiA2bLsYwqJDqDYBh1O59SXY+aqqPqv2UFdi4mYhEseij
ZoTS5Hpvp7rjEnGfwov2h1U7Ne5FOggf3p9tF/36HMTkW4cxTug/zw9xb51cnT02
149xnsgxOqtRhRQcjZ4NpyCeaVuL/bEZS6GiWlDLzAJ8bjavcZvNwXWxHFEamcrJ
dnT5xpXWrVLEgEEu5deSZgqy0UF9KG5KH3+coqvuaNxonzH+7MdUc48qOwn8KKyG
Ai84b/7EOQjpKoSR/6hcRPO2QqiQos2tMVhRXop8c9lzOiIi+6ktzrN3W3OIZbF5
PyF1PczbRKz9nMW6wFNPgNaJjOjTJO/G/u+FseQ3sqZUWsb/cu9EnG7bXR8iINMt
+PAldfySHSza3TFYV8PpnbvFNMlvXV+y68Uzy4DntXnUw1rHXpn8yfmPzOWnHuXJ
Yu0NburQaY01eSmVvVJcplsNAgs0EfQtcrX1jbZnkqy3PcAPXK73gSOt/eY6WDA/
ZiP0WwD3XcrMns6E5Vknkhf0UvvGvCCiW1uEU1eSKKv4Tf4htrKbjmfbRk8obr0c
HkvpKcq7GjoSWL4r1f6qVFjKld75fjiX+XvicyXIXfnYeq5BI89PHocuMDXIdYAo
oJnqRvWB7UoZTfGiUfbHbHBe2s4ITaTR0dUSGCwnf5sUS0rgQvVF8Hs5G4RNB/Yo
gYYoA31OqqzV//bO/12D0s/xS84L7rewvGomztgKP2rfRHekxmm4A/SrM8/a39lB
LjAppvmkYlfFtVP4NNlZizypYr/wzAjf0FPnitiPTy+9zqGzgMHrLu/kn/Zr+a2r
vlL50Waj0tBgXlMjNiP5tHbmRdoHuioK/IOFkwh0fKh+UToF3vZf7Ca7o2T9XWra
LSH2dmWo0YiKn1hpdrYB9zBbPpW1jfW6vP38nVtpjWy4tQjSqOtgaeVGi0mlf/Ha
dRiXO5bO703XfoDj/u8yKAXZxt7UFq2cwps4JQUDFgG1+1gumq/u/AAPg9bCeHuu
Nx79tzBhFjQC2pr1pTiHBWfIRMDgVrPwUFbtzD9KRDdMZlq9RUTjrQKupfi0CfXw
eli1AdY31LJA7YIchcPubJHFvvy0C9ebd7azznkOTdYzQE7KxTofDHuzZ8mGJIx/
pC+ecWtjktUqKADRYtAEn067pHwufc2shIsOVwZJErl9BW2EZYb1y6xr7snHlddT
Md3MLkZYm9Iwa8GG2nzdlTZUUY1RqDmlThQ7O/sGJkP1qlEAQcKywOZ/3x7KOJ3D
FYqWSH6AmiZGg13PI6cZDMQ6KYnFjRzIRlzfkxy4qeMCrm5M/TTYJv4ZhLzxlrGn
Q5W3lwCfIIp2rXvemrOwZHZzHb4dJGo1QOCGir8qpOIlcDNMBRdpXiEhKvdMTko2
1gaxe7Pe+LbQy+2GcLA6ISDJLCTEf9trJM/vXdxVoFlZ4YsuGFXbTuhEuBiGACH5
67Q/HqmFwZ1WaFu3NTcNn9BHrlx4aBSd3e1SmXcBo7mcOg3CUKPNZXaMmRT2A8Yi
t8UE6ap6pnUh4AAmf7YKbGLvXcbzWyLR6v5EzRV/Cacec0aAxGaOAkz8eVRW5lyK
LRAb7CbE5Qx0WDpq5wyCtQ4aj2GjY4s8YWxmD0mKjq5EDWZCptVuJZXurVH8dJbM
L0evKhcXdZ7rDurPNwZULs9pqk8kDGOZ+lYEqaHXu/oH1E4BB3b2GwLPhnEOdPdo
NDqHfztjAyR6YgcSmh1kXhnAYRg9KqyB30XJ6TNyICtpIPliJYy5AwJCrykm4a0b
ohQ/xTMJVUl6n8OTSDwG3MIsjUvXd5z7MWJfQDPgVPF/nioFE0QZ2sLRfeyjLkq8
7D0YCanUqlHPhJ6IrHK1wURrQDV/L325DKDaTgobd/xgCIJ2AwyrNBhNEs+P7vNW
PzvldaZYTg98R1nFfVHiqgvR109NxJriuqZQ80cz0yG0O9DtSYTg5PmQe29947zU
md9bRbmLjWAnUCWXHFzksH+ZHbi4HdnOlnMqZjyJNtGorYyJpie8t3nIn9xmeF/v
F8F2yCfec/6kTedC2za+m2iv6PtyuFA/57gbXnHf0IlX6KeizWY8OhjWGLdT4Yuh
Gw26SmW+BjW+GLdYKQRQVvqAp02WeebKxItI+PeRNOSR1Wd4DscBKHoodIV6i1LC
62arEvqrHIwmmsYEEgnTJyoxltpcinQNgbLs6DPFqp+61GxO1+kN9nHapDbqIj22
niQMENr0oK+9n4SM54QY6ignjGpRuQGd2cUYvkY5aQr8GI/39uCrVfAqo5nu9d1R
p5h+3TQUVo1qSszAQ62I+vROf1zBzYPrpnC0OJ/2LlS2PwwzAsXy1eCjyJl9hGRF
nFnFGFBrJXAmsflbVy8zn/K4X9ab3yyYgyJVa/y2DiZEAJkkgYDtKo+PSnnPc1wI
JmW/W6IW7xQhPr6CGdloI2xgfFE4MmpmEn99qQfES7e8jE5Bosmj5o8g9I1N2rGN
23IqVKFtB8P0WYVzZ1dAiLtKb68MG20BphPbVXKgwL9TmngVscJWvwRdpPuWW9n7
xYrTFXb3LcboZOJLdPFQ+ssy3ogoeFMMoqPJzI8ImW4/JdNgeqA5RYPpI7FphFKM
3r2jpvSBuzB/z0EtW61/w/bL1BbvvdInpn1xuWDFRCyac9NfVsH6JhzEJSY6e8MV
mcbSuLYHSwpNc4LR7GMuCz9YvuyqNnEodVUbes2OQnaSHm87SfHMxgxe8AiTq28X
TmNRmo1z1mJIW1i+EmR2cp6PR+kURYw0Bf7xVYlgMguwsee2UniLKdmpMuaoUAgn
zB/MuHuCrNtchOf11omR6HBWO4OfzegnHLSTkGRLVEih2WvvhJjOwSNtzynuB653
LNuDlwTNlfRqB/2971o45UkEkf8LUm9wpPrLD4l+pO/77PRBd1LWupvSiHMtt9vL
Nq4z+aH+P7eIqdlruxi+lJCO+LjJIdYnWCpWOvKK67dalBdeKp/MOTjJBY8f+vON
YS2nSm950w42FT/iYKuoM8kBYyv2dfYJKuPjnZCsQAZoo9Lh3vo1Q7yj5vxh++ty
HJcOgu9bUTTOEsQNlL7eMH58yJdkL58oPK9Rvlk6VOARX7qS7pO1Eb4DlbnfN0sV
2sMy/0x7jclBjKMLkBdv2qh9fVFVnWhDmp+Tr4PDvquIuDxagTeSSmkQyBgBepSX
60MaR1l6uLAlyT1nDwWLz8znJXVyR3u3H/+pD2jBoD9oF5I/cvVsHglvg+iWKpJH
Zu6r+1e+1vPlQfchIFxyexdUy1HoRYvrkIPHPvGpfC5rhXaJiFV5cgcrOlH4Ky8L
+gZfFPXbc0PWWrDJu4c2qBlWQQQha8PLFUV8VIF+WOJ2dImc1oJrB9jJQTpdsBTQ
hVGoSVgf3X4bdBLZ4nGfOQ4UUFI9Et0sobSTbhztQE6Km0v+O9k7bOBeH+GbW1Q2
0VQd6E55C8VLdFIu/U23+WZunrb9f8c/qKox7hhFwGdut0iD02sKRRfneaQwVN5j
HWc21HnzQ4MGBApSv3CRiKHBjG6Enh/jJxR39s4bNWDgMJhlSiS9oqLeV54sT/v0
UCyuHSx7gZUhyPrTzHnY4nJ/dhDXR9DnCpL2GEnT4P1mYM4K3ThpEZV4U7BCa4YQ
778pGdN0oRRdyYRhlqCRNjQqhoNHZwXAvg1P/p+RCFJGNqAhch+7BVy+/5MPIJue
Ir0dkCLTt77+lVpHfOa4DN6tAypEOLDJ+VDH2I+suV3azdKAVIh61VNhMiqwbGxp
TnCe9zIJWd49MX24zvQq7uoV3HUBnXE87Er/nhIf0J2WOS6bjJf63ZOHZf+3PAzP
4rKSA1VT12AsPQbXnY/o8Hwh3emQPTcTOhBD5VcJ+SRLpwJCYb7Pn059CYB8eDm3
hpgx5IKeFXb2y2w2sqJihrz/0se5Jd60Ca9dtdQbF9HFgEHUUkLScRKQu/iCSJ6v
AKwBEpaFDiA7M7YWTedNRvCPf60YS5pNzIv2ROLVSLNlFmkV58qDX6zHDqYFf1dR
I6JxMmzg4Cr9l7MMH5Qywy332YqKWN6sgb/wdxfh4ZYVssNIeuaSw/oKKqQDLtwE
qYj0VmhKt0wxz+BSHvrgPONrRZSeanQd2VuxDy5g2bUUXaS0Qt2NTX2IM9srg5L4
XsqO5o7zZIp/VPHBT4ENF8OaQOnKomYxadDEtRsIPUYuafK4EImTcqj1Gti55C2j
3tRLIv9bFpwcn0NKuIOr7GKzHKRgv0D5GwM4k8peAjM7HzxKwwI11DvNd4lvqSwo
rZm0s3LxoiaCOhNHTjujmz3KbqibjYNtRnDWnYa0w2y37SA1wH7pFUB6B5ENU+uJ
WnJVLcCKdCSPoXlM/C4fgYQ+IbIv9M0pbXbFmhkgG3eve+Vcs9I+3WAgh7t6joa8
Y6a6UETX/XFpjH1wF8RlmlTJ0APQVH081dTNXQahW0NbTrQ40SlscoLrGxGxqhk/
P23pC/kk2OWAjEVzjnth/yoT2TPqq/iPoAJhz+kLbpxIl699SRFhVdYbbMKY/Ilo
emHBdvZG+feRhVWMwpSqCoKfMSN3UE/OAY7MT4l0ngQEJIpiPiFhqe2igi/ZxE2F
PcDLNBda2k5WGjIzcSB1g81iNVA800eaJdfE831NXQcswI5/vSxYiff0v5bYcfHG
0agQqDCqh8NzgTn7ru09wSVmQMW6c39/TG6H5SVkk76H42W9t88GQf4ItoT23PTm
g5VY4WTg7B5P2XLpQ/G4BVGeub6wP+eUPVIfV5LUmJGQZgDgUWuvNRIvE6MbOsMR
Rf1xpHHNF5gzW20h7NRmSvh6NndAgJCL4ADy7F3ihwQrLXI6dEgH24DkEwNwvbtn
2vLmBTb4C5fmGji6U9l+3rtxiI0WJU0xMzC3W9qSWsdlIcb+RuA2P+vEbn878FAr
bDmLYeA2FjF17dIVqMlekTPUIPcsBHPk7qnCViKH9+VSqg1IFq+lL6m8vHLlTMHz
ia7j12VLnPyjcJ/hLH4cVxp3ThmltEu5D+jYorJiIFk3xxg7KEO0a8VONYqqP7DN
ywlN8biDWRXBfImr9ArAohlQmGUTk3QdP+Qa13F+l4lK+VEMzmHO/HuR+p71lhnE
O/9tSy7BXo2axhtRHsE6diJ41BgvXTjbzMOkofRp94khd1PtI1Mxtt/DGy3MHVSb
rEBoVHzJFW0q1k/3WWSnZuL3kVTZEVF4dwtMjn4fQP6IiwQcimRKX3UzgWjdB9ZK
7o5d/8JG6TkmYfvdJ03NbPrDvKxSSBUu3JZ127HXd95Cpv/W1kg3R+vioTgMPXKB
baYtqq4ctkM2/jKxQrv66MXN3j/QJ+0jr5nAB0kbpqbrsMusR+ZmgU3b068vx0Qj
SsKz/nCvrkHGjZR8oBvviiB0nIxpQ4RfdBpISy8IXICmcbXfQjg7iSxSwNeJcUcc
JE+Ok0xR+TijE8BoHlaeu7tJSe1kb/gtVYc+l1XsTNML+NSsYUQxG6+qB0u8qhIA
EXLXNYR/hk9Aa/ksHlcJ1eQh9cmAfyC6yAPJdWf+TjWjIzfqJBsPsfHALkecSRaI
wLE7q0GVjTrslQVKos7FvGw62L/N7dcNCAHoTfnjb7l1lZgw0z5/8LY/2DH18496
EwPKrzW3aDWjY6jjd1X/CK5H+OEu0ED8OpV/YKOjxNxc7WIzX6YLeIgFQpGP+Msf
eTxUtQA5idtYHSZPxySDV14TMmaJ9VslOEWX8IN/EAC9Tio6MBhdfNg5/gbgQrFV
4AXW/N8vJHrN+xSWgP8QdxF3HL2Vjgg/CyQ75wQXgeq7WUwRQlRP1M5Ii2Xnh6/G
LNCsPmfB66zd5xXDNZk3/sRpt8lF3Yucy2Rsy8cO/U7vd7M4BVP+hy/RYzwEjh3g
gD9m7hDEOJGMAcNp6myaxZspFIgB/tGgl8ZzCHwFUOnrJrZaPovcOV+NHnCDRWaC
vTBa3qOgE39chVpw+xsL9oI1CZ4QWmwwst5ykZJiTVabGxTVNI5ff23HP7PWZmR8
wwAkObMg5EedyQKJLNHztNnpeM5OoWRazSJ0ey2f6VxqcLsnsc5TSSf+rMLSGfVr
MK7g/HiHPz2XrAoiLttmZGqGpTHUYMfL2ukm73tdeR6BZP0lzY0hyPAH9vD4/dK0
qJG6eFe9rbzSsGaYVR4xln+sw2hSzPKC2NW4PFzO6RnPhZvXiVDdln0TvcTmIy5e
jjbIlywD5ZSk/bGFS6EuFNI/HYF/s9CkbQ9OCudsF8POAzkVI1AUZxtXadhRnxWy
Xwu4UuKQ2z3g6rPBpNugfOIRvVXFKXrbBOhw+ymSwOMxaj7PuM+7kt2ZsGJwI4Zr
kxY3Qc4TwkUumKih8tWD6g5kucati3BAFjxwS/NdLWectGFjXFbKuWIVIJsePOh1
TMrAEJ2d3ASa2VlpI1LfZRcRR9lge+elm5d1hZkjdw7ySM8YNjBq3Aoms/Ar0rrB
OG/EAWtT5meidAzluCzDv811hBdM6cYUFI3lg3eYUY1KwfzOzeJyE9La090EJ6s0
Jm6fiYk/0Pja3vwCRnUks7jt670U3HuqAXZwU+7T8Takk3d/sw2RDzbpXYhUx6q5
hZJsC4O9xJCPljULql3PLZZQxplHklvp16N7/s4plIw0cVq4jNNHTHnzhsA9d7Em
C469UBoLprYwbXGXmgLA1+AvkrpZYNj4MCdyo+uUatD8Nkbd4/6W62FBlq4cZwK8
x3zkdVC2JskglqN35iwe3jsPYJLSrt5c5AtThhGLs2jHzbDGaz5O8YIh7o3Lp/lb
ZgoZDBb/B+Q8FDNj7Y81fV/jOw9eMdvAdT91fn/lZba1dmv5I4qKb7yNPFajeqfa
XvB5SjNabbVaMzxQfoEwJbuBQl4Po/VT6MljDjMpXDqbRE/J3D05qNulDv1ug/pk
+84MkCFXemph5TIboIy/JWsz7ivigxpIKuz3YRcsVeKvJMqfzQsb73hGR5svwm0C
OJszXNssiWkj1gIcSxjUjzGQotKn480w4dY27yh/hoki0e8Tm2Vh5oGWuy11dKvw
6vzDf4M/4+98xRsuJHR8PwIxLA6hkyJJy5xZ0tCS7ssUH/SidihGC7UswiVhhgzi
tkaSFoEj788nHS+muzyK3qMlq2KMFQVmWvu7XxvKPXS+vOsfVzQR0MveC/q83T3d
HVo7ZgFjV1vKdsiz+qvFsvyKPSs9m8C5EiOoIcJltMHacUgBJbnuyTxrx0Sc7JED
QnRp7CNk+HIhV+3i0XVdMBL7mduKSj/GRIUaEH41gASnr3Xya5Yz7KgIrhu+vP1v
f55aRU5sTyGFH43gWT8QnbCWmtIhEaOkyE5+f49gTdWPnxn8vFRMSY9eJ+yMvmmF
dQDotLyG6hJRdV8J6K7wZrTGagfbn4j/Aud/OsK/FFUmpPJ4ks+R08KLE+Rqf2FR
+ahW60w450gUFCkuhLTvQ2IkauNv7ZZxtF34JMMeLi+jGNWZZjmVML6V++kfnEPx
iAoO6Db+RGPN03dO8ljobnID5VlvwqAmuiosLXi8ShBe1XJRgI+Hby9C9UBwIvp0
ZEKTGv1mMhXGMLBFP5plPOsywS8TaZkiT67BHwnliOUjZOX6C6bXlXAEVU/d/Bta
xJ9291sAbQyyCHJCyCUkvz7Bp654Bj42Mxz8ju4POS0nRzouzTaHgz52kWolzV20
/sqQ4zMq/NwP31dZshOkPlIhszEcLXuxlir3a4J9nMPKhvriNKTlFiqOcD7XwXRB
HtdAAHo2mFrPelgIit/wxPyNM7B8rqjvLzoHOA2aq6VFtyvsqWmXVNldHcZme9Dl
NAIfHWhKB5/VFf5jsQR/eYhfSq05HeIIv3CcNNesqZ+QUYcSsptP2eEQjuVwx5SU
8HriPweOwQ+i8SSw1QYaAlRGlvI94Q4E0sJR0sKEA9Ijh4UJrvtIK4DE57uJIIVt
JJb7ydXjIsyG9o3jo11DhRmci8in1/fm29/o7CqibyB/WwyRgfGCtAup2O0Wm8rs
S485I1JIK9dAUedp5S2DdolMzcNyyzbkaEehaqFzPTlR1W8KzS4s306nDV5cvzrN
nxbxX6OrwLqinAFQ4ck+uAVHzyN10zeBB3E7x7AgFl1vl7IGhy+Z7U0OT5AnrixQ
5+Yw1l4/jstUkBquzlOxg5dYmzaH7ZUPz3PAXbhcFnAzX1L5itUPaJd4ykSA4q5R
wGS9ZXBcSNWwh17YVpNp++fmO4KxM5lmwegkpv1jqSk8nXs/gv+ryA6lZ17FY1gO
cgsJ9d7YpPbBYirrBR/ksh6voUKq+yl5xhyTsvUA/QjKXSCdWUkZRxPDH/zuA/WP
R7Colpzw3KiE76qq68T5vleq15pWBP3l6FxQ+VePSRv4GZ7qI8Wyl+QdFJMGZ+Lb
kqPgFLUUmPfEQgkSkMCeLfndX5SvtZMD5h0K/PI9V1wtC5DelMrhJCCZGEtrFTWE
bvR1+idT+tCNxF1uOy1AD8HvMgPCnNQbGhjIy8bWtTa+5lqfRfde9mGWKXPl2HGS
XthGWKPnpgyVmuEgS8G6HQGHV3cxtEdqsCbbaxjsxpBxlgMrD+EeoMEymZkDhwOK
40AQQ/AVnX3lcdRlT+WTutyykE2Z9nuDqNbSNKZ9JwvaQm51V6+50ys3ynjJ7Uu0
RXwSM8nxjdBq7daz2d0o1GKYcvw5vJGP8QVOzNHj/BCLAYb/b7Xr0fmwW0LCPr5B
Rmq4OW70zS1s0dYYHn3LVPVEMeccWpRvFBRo5K81MpeWed7dUi2AdXby2cX038QF
gJkjPIqZGdmnU+q5zgIY1FI4zLicSb92I6u6RQnJr0JyQ4Uep6TZ60HNgCFUdlCx
rsN0WptKKkLtgxcL4ioI60L7KbmT7I2i5DHWASrE/imYS0p6zaNHnckMHOHOm/2S
H8g9cOYxpOvF6AeB811eZRDikLN+aNpgsBk8aLotcAowM+GkFRpZbB5mSRyynghC
xpNqaalC15xXESFCsuuVw4CxfLzF0MIElyBhuBMMx6BzZdGq9o+b71iWU3EdoNCy
q9Tq+L0lO3BW0xglnDZIhnclNCMP2M3UJOAOdqb4+kYhksS3NHEPyFIGUP80iKLt
uz2a6gglMmVwwTjUPsDMH1LTZ+kod6/NQ/iaxba8NeDplwmYw6z0EtKl70K8jd5G
ixuuU+wK+eO3Wq1VS9latAtLYs8RRq2pqMgwC86NnQuFpUuP2EzI4YYXMAlzWajN
GALhTbPGTTZ5r1gw99tLhqoEll95BcYEZhyXAT7U0ECOlioeUlHm4PNVpUqZXPyr
aKfwJQ0ZEaEDGAVXJZl0LJf3aZ+pFdgapdmRlVop1PXSWT7pHSapc015yY0boWIt
xc0MI3p89isSKAYQMBr8/lWv0//oyaqCrDOyMtEirwCjIqm4KWedjjTLVdSkvDGn
T1ee+T3eR14uXII5kdBQGAhtM0qqiulQyipXooT0U2bxSe7BxkrcSrvuZnuMm4Lv
pcgtn6Yx8h/PBnBMbCJHEIxzLhRjvc/qMZd+L5O7gBOAIUwX2TKpcn9gcPQ6b4Ce
KD+qE4uZ8viopMLlEvTw+8vy4vBZC00AYNFRi5O/JNVjxjt0jq87q1NGeRKA/SBU
XHpkJWg34qA5r5MVlhkIir91elo6CXwkQKlH9AWZPVODfWko0GzKCwFQMaPrJZZF
MlGZvI4SwzHBSbGosEW3ei/vBlBJncyx6gQRkV7LRM6VZ9i0J4E5AwMpRHoOX8ZI
bSRJyXEYRWkySoY8zaGWxKaEXHkDWh67Xrb1yKmbF4mtGXgYJM82ufH4EkE5c+RQ
YpjKDU6t2h6Lx3YH1eqE+hHo+kmO0bFoUF3/VE5/ZXRh7xh+KrdzfhNh3wO2ACzy
qDO+k3He+4/7LgjfgGZPY50HbsSfZSlKmB9pwUewlxtfiGhHIQUUNTnLcOTDPyf8
mwFI9pPEsOU+s2CRhnYJODf+XU9pSjTlvMNw7WbhrUjE7eSP8P31ORcyg9Aez0N0
LfejoXI45NJLmYBBRYTbHMWK5jSotWGgLFRcKednSENvdsgsopef2lAPurdxYn4l
J39MNjxxerSsh4LEtlRO1+e5MsKXj8bifd0AOf6arFk8wgJAyFXw7eTEYRydxcuk
soSQkez3nMHeyO3Dsee66Dxa8A07Ns8j+OJQETeCxDMdfu9iW7auGVETsOhaSyyx
zsUjZ/KzEjT1qvynajxNQbbiKufno7G+vmVCsWavCRYgnenX9DYXp9w4Xeucx7Gh
7Cd7hB8oDigZWH7fQAQUKopjGo1uKMTkDdpnp36N9O4mAh+11HxaHG6spx8ao4v4
rr+6KlK8an1pVfcQhGy2t5I0ESfRfMJHjha4Sd9vI9/tnQvkdXPE6ERPv+5Qnooq
4tcbC2/JhxfVCsu1Njc8g6ghR0CnkNdDlNuPrQuG/2sE+XWCxwpoKg2L87LWqFo8
978UtUQldyxef5ULTc2jJkYQ9NCqZ2OCLes6K0mWcaRzcM3ofVdxvjEiiQVhX+/D
ZSmTz++32zJADqXNwXAP76XHnVwZj90Uyvzq/iddDap7kWynqlRttVI25aTUEk+V
6o7/Dn+tiz0hW/YfOmyVXIF9IXlpexthMnNJRa8ef1/Pj7m7onMOniaAdxX3tTMG
XwHpJCvXa4bmGm0xnweKSkvkJ3BH1iLm4MQ9oo/Fmt5xmzXaYL9tLtDR/PuvGf+Z
dXCW/iFDvc964k1Mbqe42YS7c9sfpYZJ9YfjIk0IloSetJCQ73355saJUa9Qn1Vn
OB8t+i7+ckOSSawL0mLbLmEux31evP+kzcS/eO1OvP6dlXtMwuOSlY/QSyYCig5b
zXlhmRh2hf9mRoL3CWmPcdLDE8yp2WT0w/MQZS0+PZrhjFTY/rlzcG7Q9XBmzzMR
cIL5nY9joYomejvwQYeiyi/bniCrchWQr58Ozzt2UgkE51AHpKAS7EFUTyvNtpSC
ExOS1RLf3Nmntue15je8D/VQtd4lVyiweFBUsdwN1LDewtgKYjkQTNXq5WnW1ZtO
Jn240RAeRoFhtjtubccaXCdlvuofBFjtF+wxGygyslimuJTb1tODuecptBhHraCO
rulsH8MJLGAOGsQOm/Nwoj/2VC02An5MwhgqIzPpTPDdJPe38pCG5I5wYoxcMcxA
fyyNzJeK4ET24mT5T8wsXfU5rv5y0lTFvyiC4NZQxv+vD+YIcmfpKkmQ7s4p0jZJ
S32S0JMqrNHtmY7zexe7xNiyqvx7XfzMYMORwA8Q+zi33OZJHz66QtrC8D0R65K4
XcFAhJ7FFzUd73k74BLwNm1slY5gWWYQk/ot6wIaK0rzg6iHhbrcJL7pv0MZm9zz
Io6fUm2SOx7xn1PCjyHcqN65FXMInZdeE6+VsQ3Yj9tUkhO0I+OizyN/kt8cueQH
mlV8JVYlWTH4YFkYiGEjSxaoaSGC78P/hnpMSv+qBOz2DrlVpsCKaXrt0sIGZkvh
MrY5LzOmSr/qx2GCua38i1YiTKX0r7C0rhdj9vf+q6wfnOQOSa6RvR+PgjlU+RhN
/zis9266qnyOUQ9RqQNu9KRYC+7Vz/xXAQB1FDjZ+l7rpy70UQIqeFqgolWpW2vS
GzccgTPxVspzG5+UJl5vRdXjNFErTci+yeOs4X8wEY4IhipEmryqkZAAkNP9VUpS
t9Cmw/lE/Cw+fC/7/Gzl2AHBzcO/Xkme6k2w+JbWqYlSNnK4fvrc+CZz9NTfvH6D
1dESik9zGq9/7MShks4EIDudUQudcsvilEQuweKblKnf9OR+NjVU696yHqG0b2pl
JRb51KSgjvi6ETN6/r8wyY1iMv4ds7I2Rco+2Gb1h4wSnAHSTCApFgA4qGlFogjs
gechUh+8tuU5QFIMGlYBBr7M/VVNb9gYElx0RYwVDwcJEgHs9eZH3DenJANnY84A
SgGY/P/llMmXTx7fQjZevjCFB+BCuP1vIlzj3u4HE1eJ0QC2f0OnVxjZFDA+FDuN
kSAUP1UHLS15vi4WO1e18R64i3nNZkJw6GgScFsBR1pzbwnCCEtEsBmi41Mmh1yi
vN5XNh0n3Nndygtg/5QG7zou7e+fiFBWwsi6gF+3eZKcOHHg+Ig4Z0+CIgoDh0ZN
ErYdQM+S/3Iesd1XJYckWR+v36CwSqe7F07yGTHp6Z9NpaX4TASuEdMvepeB89vP
49yd7vW+QM4/AcaW5edHcO3eECKO2WZPxuDjB8tEDm+Sv6k+VY4ipoQ7ztXCKsH2
h71QsLlVeEPdBQQ6VuSkw31M4InSjFUfhED8H3C7KYcE3YLgREaDg6axCwKqbR/l
04RAdjVtsogZiJrIwjuNzNICyuqWNg07sckFiDzc911azc7rNmnEX0iEFVWoMD9H
uNS7RrY4vfXB98En5603yXAnCh268lBkpYCnpHDXXdhYKkTH8evk1MGq7xklXsIx
pTCe9UMHVA5Q6apQxVFkivlCaO5d1CjOlC4LukRGaAWldNbli6p6vpMxQbzOCMZj
I9KsvxdT7NDPDo+oZMpYGSh5uCz+516lkrHy1mlq/sEZu7M2XpsMqXSYGE3Ax3Nb
h+TG1mfSlPB9E1tsUBNodFlcK5ZT+7I145SuTNtKRtAzzuSy5mfiIygJxvOaxqcr
R6sNyOSrjktD6BwYmyAzf28Tf+BUgoJG0ELB9mX9vmoafEQSu5zqEo1s84E9sRQ4
A74pNBIVn+Z2kZ2Sei3j52ImocKnsyRvDtXh7xXaprSgFEGtAOq+/8dsAhbQ7ljn
8wh//2MARU+4GEQLmbSAHb8oAn41XfSfw6R/cHFWXg7TV7xjFA9mZ69pneb1llHN
hlUw8Wgo5YyxFDuCux8mcqjX9MAGqgrI0gpW17dV0NDggfk6jaQjboOoWqigQxcB
2qdSxluQ92JNqQUBJuBkN/iYP3AYQN3h9FbiPvNkAzKVu3iyElQE5wd/dGoSiq6X
GHi5QO/BXiMxabGKcov3K3KLzmKbqYKXi51Vbu5FFGEZ6FmgGGUEafLThKLiky4J
yC9yaaM2Iyo2hKQ5SUYWU0n3r+rWIDpiagdoUISPSvvgDRiOgLn26ECTFZAqziT+
IaB8ipKCkpr2KvLAEK/SXD/zP0Bg3veAKlk5DZvklvCBANFWxOdpRLVdXxfMelRY
6d7mrQpFGU7MhU7GWUpfqYQefuXEotF8BhFnI+gbT3UuZ8kKEbxRtoWxdPpid+NR
JtxHuev38EgqZvHXbS5Ux+O+N7fIYnU5mb7F4XNjk/FOqFLet6Yn8G7qzZjs6SPR
UMfUOF/ndyNMLWhaC0g4Ko0c+hNav8ZpkVbjt9xoWF4GM6MtBgpuxmMfA2i2tHMW
dRaZgSK5E3zYOIHSUsMPosULykaySKM8KABE+2+U2oztcR5/K8QmbbxhTZb8akkJ
c3DFt4bOX+eLbuS6/ivxxOAn3C1CrTkcMGuH6yenjlg6BoXXyDtPSQi2JOzm9haN
GKbgOFw7Jdut9ma9LakAuZ2+7phKJa6QQS85AXrjMhPkCyDREZaf0AVMn8Xd5VqE
Jj6m3xuM6xjpUa1Vd26BPsbnQFyne+KIa24HKS0kx2mZ7//Yd+j/ErY0gfAj2s4G
crbU+Y/Hl2C+2DAV32beKN+a7sfZZdFvKdq2812LE9DDDhdIhg28KMPaoCM21ExY
h8uVBxFuAkdg7UP/GqWnoYOJV2YdX2qpGud6KBDPIxingQit8SR2U/aVZMPN5HRF
PRvQf0xDz0gGYAKA+/swDfiMU+tvK77pNla7ByQfj1MNmXzSmtXmXQAKGPGJ7m3Q
m4eJk7vLkyurY9NtK7lMtXPvZSreDcfvUaP/zzemGSxaFdE8ShVpyOh6RGuKgVLj
+4bRE28BkYTg9Nw4BKYNoR3aFIdMbj6Z/ThyqkdnZoj7kp8Ig9cm8zUF4T8iVPll
zS1BW3z3mOPE+Kk4K0zmFm92wFidZiTfkmKkXFx2TbljsHBu3YyYIW3DU4FPa0Pn
kj2B+sHmYwdxCD5IDo5YOpmbG3edzw0HbTYdF+DVybDspjLZEAZLs68+n1cxqg4F
WtZK75EnUf+7O7BaRJH4g1gOeWlN8BXue/gGgFn+5sqnFKajjkWH/aZ/smPPgj5g
Q93cY9Iy/YQ93TTrqT8Q4UStNsHtCpsOkrrLNFbIWybTlYTSJR9HdIadW+T8mp+i
1K83xZDyi2+g7qn8T3TRJ41HSq6+FIfarm6v3bFiDHChZOmcBUD8G5D2qxkq1uJg
VT98NO1FTCoEQaytB3gWRUIKWBXezuuev7xI8xylGugW8x4jF4pJWoyil1yXNRT9
GBQFIjG4fRoWmUYpcTedadEVkwSPqlnbY8raPcHBLEPETHrTiEGEQUvk64cW4oVc
9ziniyfVOdFmvXaxTAZ01jbmlDAe/e4n7wUkkplb4XKIr9IDYaxjAeA+V21WedXu
on2XrXcVIF4sXh6auans1Fj3UbLiyrdnuI4BY1q2JtOQgoSy9YfnbyukgNiy+gZB
Nqjjg0XPTybsvGS9+8dzMMKHePUHSSK0Nex6K4rcovThljChJ0U9SINP/HFYcns6
Qab57QgxltbZavfP7gyHuVt67QjOjd2rDLAx9+bI2b37jDN2ZOEcYOve61z43+fL
jf58c+3JQQX5TpQmLq0cVlTHP7YSMy1REoyEwJ7nSWp87mqAifQP0Ttxmnwuax8O
A92ShKuWJH+LxSRt/0FERkuaZHV5biEQ+iWG8rgWW6T3lQzEoGRbGObCsql6/OtF
gv9ek3yQC+vic7HuSiFTWLXWuHYLoiNV8KUROJpLNpiPp3SrQt09peqMuBONEN6h
eVfw03GTKUUwkmpa8CKKm3XnPluwIOzqW02Ox91EuaPzwcUy+a7j5kFSqasxdlD9
wsxdzKnvo4T9tQaqB0U0SPmcUv3Pp4KgHkn3/K2wVPaHDmgreyay3xkZe9GE6TTL
61j1JGYjtEqtCSrTRy9p5s7N8xQPlHBIsUmxy+l//ciIZlWFwnlPrBh82wZfi2nl
17A7UlpHadMhIJd4p4mO0DrpVXtcR8kyE5MGcnvQLoxbrNEWL6+Y9W305uIeaSDS
6lnBzOnuzuWoDA+eMJc/mqSzn6OGheM4PISiwOGG+7CsFyxazwPV5cRq0BSXKlPI
nURJVgRqc3X1Edv+4FtYsHuQIT88IU9ncqfoq5C9IAdv3Gj/Fz+bFS8emJp6riq+
PG/NIIzhq8wUFJ/NBpVF0lFd55IsQbcU5DwLPAN3DqRFx63XeCHruAJl3cbMm4Rn
Rp+SRkRUQdoOUuTaWFxutwf1IT9+PvIjugZntd+YCYMD9zRwqbfl6ezMwF8K1M+z
m91GwH9TQYiVCUGT2kSzBgSGn1uNAcaZY2qGH9mB3/pC4uvbOKe68Dq1b/I89vjI
Qfunb/vbI/eBIGr0mFbuVaLQ7x5OOmolqK3Y1PcpCelWqgUiZOD3KbfMipguu8hA
x3vrE6QklhkbXlpcRF7e0G6uqDhoEM4vfq/BKgKsThZih+RFunXoWteidhdIDJar
cb75BBUkuEdiCCDEhaeNo7o9KylNIHVu16dwU+bpg9jb7pDwdVH3dRAvu6dVBRnQ
G2ETIlxznK/h+hhFUP8gvYK1N9k6d7ptouFk34Oq1LH9Wrk5GefzKCWq47hG5VZi
XYmizaYPtXd4cJdQXOWTcUBFuEiAX/JriEHg6GwXa/RFtBx58cLTk52NgVxnF366
bieBMQ2rWpjfgrYcMQ/9lhkD90rLfoYLkp0BftKTLi4V6SD1FM4q1utAytbGFeU7
ywVvBNpquAxW124Y43Sg7EQPt7EunEFcLnwvzswst5NeE0phCVAw7krpssWnuEUr
ZU/FRL7BGqMi2DH0OICl04YZ9QYh3jwUhNy1II3ViyVUgOontQYwXscxGqDU3Zz9
ueh5TFBrRDm126/8xew8xtGokzciIXaTJ/b00iW9kgh2DoNOyxHYUJaY6RBYVccy
LpUoFClzYpFMGerd8OChKQ7xNdGyqn2+HeEMLPTP3T8hW/rhIryZmlr2c2GTgjlr
Y8+OGOf9Vw1oWqLF3BF+/x3vDilXigdN4bIGgSIoCTzBVQgG8iX7fFyAb+KzV3yb
vvKWSz+jlQQi3N9IWZfcuBXmyNubNusdHCVAMM4adGg33ErcSFL0+hdpo+OTPwmW
KPiUf4wvBgHFzH5u+kVxIvLgVsYZiJ2R0pCQIOy8AzXb2YD8wED5MtM6zkgTqpXY
YuSjwI+8PzggUGPM/u3s9ZU+KGa09EFSLKzIzf0YksTyvzaD4emj8tLWqsz7AJ5A
d2pNKRSf56MJiHLidtM51bEdngHDeFPtXd45XlzAiyvrc1VAc1FGHBxJniTF6ne5
+3ejqLtg3AZ0mWQiB8Z6ykW9dZ0wVZ1dIYusRmvml0VhDCMgX+nUHAlee+2c1eiL
wzQo//6XBHDPvDXLuvZUe2ATDHwFcbUo5PCwlUlmfqwau7RoSFjTnN+bm45/5IZF
eElzZ2RGEb1mK51MXxvElqwFDvE2kKfCfC+wX7nHqeaByKsencM6cqbax4xTLpBN
32bf62I79bmCtdjJE8qh7uFOUYB5do5RTzVNGpirXYBrIlQ7d9mqMXRL0bNApzcO
ZFgxw0DoHPPCi6xY9RAdpAkdYe4q96o+l5mrx3fdBkd3tNyqHXpjXw+zkozg+VM6
tILfaSriNlKC0HYJsf+efiQWzhA9AJ+aYLInh5jIaVf8ZdRdgWPaIBdYffM5zif4
G5iaJdMmxA9jLDPG0OdzU0Jo9d/DKOGcuFrr3vdahKov+Dzs1sohlA2PeO0WquoN
4PdWkv7iLNZzW+8IbZ/K0IC9BZtwbXpyjYGa345Khom8jbTlKvZlGMJ9Ud5aHWnE
UsaGJjZJ5rItbPZnb1veQeqCBhzTXJxm2GoWDgvCqtFXkh4LD2WW6EYkCKMzdCtn
9lw+Tk1gpBryV0V8ONSDybh05egl4Ws0hqob/KB17uAIUqo3/qUQveGf72uUnptG
GD/w1vm2nOu0ABt+DHC/P1kIBZRv8wU9aUSmaj3gEDBR2P0roF6xrBFu0Y4URngP
yILRyGZiTFZrAy6sjlOgLQ6azG4qrhte22ICm9DVpnYP877HONNARxdDQG698KIk
0AgdL6PhUewYZ7JNGy0cqbvklNRWKpGz7wogS/37a/g+A2sVwAcfuNTF0NBPi7rT
IOcjUtmbQo0A9U3Kh79HEd0LPQ2XN9mIvguPPFefMR19ih4f1LrbKSsSt6cAFHzM
nn2WgiEEu2uMtwD25LEgJy3SZO398NmcS0aiXQGCBVmUJ01KDOwMCh4xNpBn39bx
TqPYULbg96hcB+nhNjXPhw02lWFU9nS1Slpla2dQfzQ+Y0zDfOHSfjz0DfuU4qYg
GqzRLB8Sf53B0GOMokSWrV2b/7N1vn2YED6lNeP016IhZCjvs7esFN3m5tr1HB6I
WfIuNRqp1jLNT6QBAvpFwTkDEqOZ7eIeD8ugbvhzSt/hw9NoC5/tfEqcTHz6pmyL
xCV0AbTkdfDqjAR5FwDW0zUCSd4F0goeOcmcjuiGgU1iDhlmS2TSuAUntmKBlM20
HrDdfvOjCzSKoVkIBPW4QCc/PL+B6lMbut5SXl8gQ3aDQOe/yNpbb6Vdp4S9cwPe
hQIe1z/Ra0/0v8JgWA/JbA/yaVMH/+VgKZ49Q+zHqqIg/keNnl31b4vB9wPB4ZGs
RDg2RDbW1PDEdFF2NlxYOkKSWyjFM3cw5St0vNitUogfXHNcblijkjIy4S20Bcns
Ge2SW0ZVr5mHlk0Cnvi2gqPkVN1W0WRA07tnyFBatKpwCs9W67yGTJIUqHdpBwFq
PpsEDvFG/Qg++v9v9/nwYTge+HTLDhuchd5e08QCW1BEvtplFj4GQ8KxS1G1xEGr
F/sjz7d+YJaN4zSxwh5yUz4GT5ZO4HsNNLBV8oPYmcTGJcw06tH+fJ5tbRKOY4Wk
lQ4APz6reIQjHKMOYffiEEdrkRU+RUILfK1HMGM/A2NSPv0gd9coZXh0Dz5QocOV
PHWziwfGWEwECEcwfggSfo7PfcU/lAItWnp0dcsLNlodN81xNSPgen6XV1dt4YwF
zMfsg2KH5SPzTgjOmj8xZ6tQAL0x2oPbFNH3MRs6l8gEzdQT8vkFVwfS4EokN3nk
hMmgT0g7CYSVAuYHCyj52WOM+OjonuGu3vabRSr/HaSHVRiKeISZR1SZwYv3UTK6
2kzBtDz7HsIgNk2vFYB6c95GlBtZ10yT6pHJ4RqdzOLc02044GQ1edUn6a5/jdmt
92P1SdFCkMYa1zJr7ES06NML1zArYOuCamN+7uTT2247uwtDW6b0AdDRONbOYxtm
kDvGAhFn84l8/BkKuvxrjrH4t9zxBYLtsUk7xaXQv7zrL1n3xBcg/LVZ1t1ORV/W
sj43gK9vELv/PdSLV2S5n0FomlR9F9/JoJtqffAmOF6vQ4JNUX0fzrp9TsaoftvU
ZXO0nNqm+S9XiL5F6xX2nR/ixhzC4oxTDD1BMfdJmu6IpjWf3zutCKiZUXs5tgj1
F/0AlFuUDeDGsKRML3JgtEG9w0UQnL65xvptRMBuX8jUXHcu55htHhJEqo9UO9r5
Yb7bSbfCK7v3jWOKN+W+g4F0uc821WJsC6ngPdB5rHxA0/s5UPA7xhh4Q+w5g/Hi
0UMJw+Ws+fWvPJ3cC8KiRerMTsaGsosMyED09n0wb/Ar3yOUa7FwkBrJfixWqjP6
hhyV+xbGrcCxP5IPoPZGtyN72uoVHJ8iakAmAdVK/3n82x5BnwF0bXE95CYjlG4E
x2reWnxWQueMunCauofqfWsQG072Hv0Nke935TgijvFFMgsSeS57I/4UMcBqePhB
lS5Bi6JRGK8B6/mej1b2t5l5oBRYtSfl76a57LnKtar8zCh8mhtBcQ+QPEA9HjcV
ygg2vRZ38lPOAdZSQQ2ZTbHeKsuwQfBWWhx0DRETDJqLPTuwegmUmhgE8/eskw2a
Y1vRBbZgCFmrLh+DW8GwRUWpNmMqEFn4BCFvR526/RiX7XnwwubpflQQWDXES+rw
ggTdvm8k3c6H2URQ3h8hpiNlPxNWWNYVsXAmL9VlVtBAkyKPn7ZLK4/lnr0YkxjX
YDmpXMQ184vJh2PMDVy3y7yL1gs2Z4oorlyAVvghN3rC0N7AL81qt7UbOzROBxET
E7KXkSIkPZyA12mBIkCmec8ba9bY5zTY9wPndm4ajP1fnE8xLzAj+U0q+DhjmHNH
pdGVvBADPMuLYzrK9O+PhE0R29gJM2S0KL8+DclyWG586mNifi22qGM5AA4IlvHb
pBmS0sR6ZLAvyHTX6LKz8tFX77LCkba3+vTwFEmP9BqbqcMxnY6d3wwWh14HrIE6
L/Xde6J+0Sbfh7w+4VxTCdywKRlNiN3UMXQPKr5OFcWzwtgvRiFpyBlkmTlpSJpm
1Z/wQ6P8l2c4+FnfDmdtSu7zp78bm1DABf+KcZsw+xh2197DSV+E4xYnWZoreo5P
3jB8mJyTLQx0WBFmKQA4E+GSpdxYZqyB73hnz83qG7YkhRvEu6F2ulEyV1WTM+7o
Z21e8Fua67C7/kGBx6MCCMAVLXg1BCqdcacgWKUwedHfGCFHZX5phAUP6yQAoqCI
/3iZDkHnN6uNLIgN4zsPG/lry5SNAmSv6P2KUbJgGSPmOcK36Ij8MS6cuCVwG0AV
v4f6I+v29AE4dWp3IwTtIcLsVQGZCM0Gr/28mF9LooegTxKIWTd9IP1H3p/L0knP
JQyPz0syvkkFL2CfH4qZlnF3n+pZvZam9vcVtCMJLrSVjR8agsIT1OLj55iq00xi
85B0oBcKvJ/0pTQcxBMLW8DF63c56Kt9P+K+HcZpTHtN3oZyEek3/uSYTKqyG5uT
wC6KHPEXPpXCwhtRkIcOJWjBJOHcM2CLHk+VEmxmYcap2oCEqUC4lI+q5XMzm+P7
RC1mXFYdkRDCG90MYNPVIiEhMU8upL5T2LnfcHrbKqOvLTMxTpTj3TKp6xkbJQ9K
aNX0VwvUIwmukUPcadlC6UUtMwxOnuC3BAM8PpimzZziqaRNWwZ9MbQiAG/1n5/3
dWv4is17+N8jm7KLHQQXJXlNG0+RgXAqSCrJTkgySQyv+5z3ZNNovsK0sS52Ufv5
6vvBOeW3gSFbHYEWPEAV0ruTciIbvRa8jiA+KrfjxLmxmFHLH12BkIs4+ckRPcB0
505ulswPr6L3EXHhbIsJmsPYTEflTdn5hNCWiA7oLBz4ZsB2UT2nIcSeIMppHYzt
t0nKamAegrNxJsScZKbo9wfcUoDh0DY8e2V4uxU0Ol4ygTGQ3or7jt6lWOMi+q08
VwV7XQDz2210FVPWjf5jktPILhI3n3sGmLKhxT0Kd9UotHpGIw1gWzeoPgGa6UZX
5bCJDtuC9ZRq58XdduRVRq70ow13ufwGTuv4Woll8oDWDvXw/4/Oko6KU0x7d9pd
0GTbpTS8s5dGNV072oIEZxiuZgzrhxo26hSGoRf4Ot5NFacbr3UkWIEu2fE37738
qUBG40jvPkdMLOZ1riwURPXSh82RUoWwDbxToofsuO+S20JhkT3JjdSt+E5bEhUf
mzxyhtOH41tVXeUAn/AU8B4qFT59BRhNYIIqRhZ5syagIYX4ceZB7wcIsYg4KkZ9
2rabfxJzjUvpO0mvjtPKRk32rdYNBJTHYOhMzhSr+d7phIB00TgOt7ROgzdlFt68
odz797pRqnDSWY37mCQgt9hN6IRwXDzONoonJtuD9ZW/DnmHkiUCj+L0viqngZhR
moPEGI7EcMZF5CUOuYCyNt8JPKwbOU9dqF79CmABmGLZdTuzli5C3yTv/+BCNam1
NIoWZE9s6MokY9o0kzyNDXmkx1OOeXJdoyX/rf+jLU3je6eS4tP3E8joriJmCcla
eEh0zkJRUypwilFAgOYSwZIdwg4+XrcBQ/mJDu9g7Ksh5A2VWgBxLUMkkDzuJQ7e
ybmGFDp6bINMt0pOeHt9zp+b8WRoaTYGlYyPBceAIPXLP3JtVImjTzZQ8Snempix
6vyxPGw+WrkPMJ69A4QEdwPZxpHxHChPRd/B6ygX3pAyfgAAHcaEDJefcO6MBTVQ
vXoQ1DtvIVYZ+ub15DLsPaFCaC03KUYgtoDV6qmZZRnARVOP213yJ5hcxXzgYGnk
r4GY7OagIOlky1pT1nOVrMN4jqZ7/N67TLqf7cYoVw3fzGBPmZVtsegLJh7ZKYr2
qnM8jidgTzsmF5qAm/JTIQN+YiTNYaPrt3kzHdkWU6+cBgKHJc+7ZQ3oRG6w09R0
THgJu/OBFAtc7iOnb7Z0tjRCo+M81K56l8OjplS0B50erMepv86gKpPBJz50t8vp
TF3B3JhdN97F+w6Czk/3IRJiVMOiFUEZxvIcpLvpZ0nvgIo1IGPIflhPb+p+9sdP
Hf23mmNyORe/WPWwYyrLUc4NnUxzXBoFzCd6U8avW+JSmZWQ6pgPBzIWimuKgqKE
l+f9b+QbVHA6dpM5k//eTzumEOiBaDdCJyVaX4MTwvD/m47Rp6USSbWcjizgLNXP
8SkmS8OTi+IAhf+xwmYSIIK36zQI/KUEoa92oAUsqzMxPKM4VA0vSaluFroVonc9
mvxK4XCsPNdtHe9RI/tHWLbQlCgZGzL1d2w+j7y9PY2mvNe9+cA4xa6PJO6U8G5R
giNJmmkqsgfpB/gylWF4pIPKzTOcc6/lEJ8scYrzz02P6PbAdrN7ntkffHFIhTCg
nsXbcVTXJaxL9CpmaBzqX12NffRTSHswLFFQH0SO6kYdDccJ4wSApYGKMcu72eTv
oYcJElMFrECl55K9qSXMfmFMvmqPxU3c8a8K2+2m02SB/eqGsE9VhLXhNOJCVdXu
AF4Ie9HP2KBWD6e4Z7MnGiFzwbCvFQBWhJOHfBpzklGG3BlDDnPAY5dpB8bvWPcp
CL5EcvIjQ7Omo7e5UXCtV89JdoCRYwf1lnYJ2ruc2h60P6c9R8ZlHrronBjCIyWD
Prvo+OWdVtDJ6Xhhnu26cI7iRfcAc0+issTWRhZCHPzZGckqpX1THFm0iIgff0P1
eEJyGMC47WB9IQzGIjFJC/vwOuDO6BDP5xoRISm7N2flk/spJOgmKET5DUkgcIda
ZCQJkXKLcJU50dBzsCAEAqcqA6/H4pvdJ6yT65wqT7FaGW9cIDhU2Ws2yZx/ZO5h
1oDqp4QYH02jl62Cb3iooecPE4Upy4RJ9Y65wQhrZ9Kj83IzZh9ZI8PKSG0NNFLq
jWykTRiuD7CN4l0109D9vj2SwUfaQhfa1RDpwfRozynsZDHti+ehA/4oxuNv4JYs
LkmClonhr6PW4GenMhd61kRsAKMTcB/qzGb74PF/ZCYt7C5dgpaevFIh9KV3CvGq
/x/2uNqJJANTA792zzxKO+27vnWqUBkIwXhk4O04SZJE2HcAL0AsVZs3oLH/JBuc
D7hG4/+hPY0BipKlyVApkXzhgk4Q2D5qYnN6b2/110RgBQnVuAgEExI/J18NyWJi
0ET/abfac6KJiNwRpETsD3ZCDITphP7i864t5QztMkI4G948vezcKOByuP8jMjDQ
OPuuLrK2cnMTgpX/4nAwj8XehtjYKyHH+E7HpyqNBvDPAz6/6FsUG9yEnjaOwaJX
P/pDAXp0/gzYzC53A2lcuTus4E/TUwv8Y5pMl7Dg28U3DCrnFrGkXMq7C9Jz93F8
L5Jm1uNEqkxi+AMguJsHL7WFlbrBRhtbImYOMdMI2yS7turbMuEoqgc7FN7WxmvF
nl4y/xll+9w28TI4Y6OJVf/J0/ueqAo5h8NjI6l/S6ASGvWm/Az54cAQ296uXTx5
KZHvElum3MXLOHmPXrll+zhcD3Ysj9p6+IZrIfG8oB5EeDInCkWnqsiewyXWQrL/
Zcw0wmz5U/e7z4E5ByL9ukrz01P/ncoDMUPioDAvD64Bn+ZVI5p0eLPUAcxQLUOH
3SfaDZ8eWyUbF76kce9FnoLD+byzvv1i7UrvqfNTz3Nc405T/e7uQClPesHIluIn
sFuL7ZmWz9ABj7lMWeHSG1djo+Frmr75Uhyhg1GkUT+uUnbFbn9/Fk/AA07vzCmc
OngThER0G/8IQg3RKaQAdhETuu/BqCMynpfI/sjj5prCoxCAhMFkDeAps02gBp+5
uJjBvxk5CpR1L7tp2FP+XHpk+PRWr8rn8V73VM+MJ9807tT8J3J5K4X+ln1UcGoL
yN1fb/+WAMgVKzOK5HvPQrczfr8n1iRm3hwSyOpwPSRQ8Xgwrbi4BbO9/sAeIbFq
kVHE8Vt084ZDSb5IkMHMVQo9y652XhRaNFcUpwqJw4jSP2c4glJKyagSOF55P/sA
ObbuzDR0AXtvC84uJSeoSSNY35BlY1qT3m5YpZdf8AGel7oYHIpTaEhj5zdhUzf+
b0kTwUOGxLSdehc37DuqA7w8D0631RYy/mYpdjr25ds//0Bg+xrqhY/6Is2uS5kw
du5VY9P4lW3ElX6S41F1tnVMUINFHKbJNukayJuqu7JicQXWJ03rDCMXHdNweYq3
LSnLJZLE7qnVrVtUB+cRPs2skirQqH8+wv20vuqAhBympVb9E3HEfOZgzaodTL9z
pBCa/HGrjFovcfbENg6jSKyiviGGwzJzPzEXeBIAHbl7ZJZEioH1pI3KoDPRVuYu
JOs9ZnQ/GCBlReeRUgp50Ao5MW+241HPREONgM3L03fKhS2t9BpmVqocN0SMUNjp
hM3ukFHcCUn6sWQO26gYv0PVq0w++es5FO3sCCsSSmpVrN6KTWToHoc2GimfoMh8
f55rkhbUGAsqt941UykQXM+XV8xdngp9cY703V+/HxD+QmDGV25cuvUi50flQP21
4qRX+JCFPufpNlcY3FD89sWiOeu6D6ESENeXdW+jnqhjkVrTVjSv60VTBdccyZsu
8/MX/nrc70GE6PEfwo5QwLBBPcU1DEVBhiImb0eVA8R8Qc75r/T3itZLH73pEvRn
PsfdY8HPaQHGm/IRHAaKET9UcsMqntnRzA8jYfNJzLYqwna1OrdPc8PCUkWaJReJ
0kC9RELSEx3ZtwJGb0d4CvAwzuBExYzZW2vWkgEQ4GuXJXiAVYnAD83NyxYHYJ1r
ltRSomCg8vZRvN3iHT9NAtXvHm5lL/pUFcHukscKierwCWHT87vCM7sV9Cl1smXH
0FNGKjigQs1/w0nHB2Kh2Ly138jeC+QHypM7SgoeXv+T8JDjI8/P0PFjgo4b8j6e
JYJch9VJ/jKciYph5FR+ma5zJ/INqVj5tCTZ33mQ7q3eLurKG6yB0/U/aUyb+XSE
dw9g9L1OP/9EDBO6HSgaxNamA+aRmXBXhlVVxCzCWrmTSy2/5Mfwqzuuhz2xs9x2
tnhsPTpHbPtm2EP50Y84G/w/21E4kZvKf6/TAlGaf3DXP7MsN1bI/UiwjaHzxrQZ
FR6UzgJO5H3BFE1BAMyvDEji+FPFXdNqbB0E1WBC/2jhTg2BhnWEzvv1JrDPjowe
5jfYfD510ndOV1gBBVyFCciLGvryLLo1eSTKh8sctxyA3fm8HgitxwIDGJ50oZhY
hYTTSendNAKbnh9jy2dgOmNgbSIeNuK9dDG27B4ovP0e9J19ZkCKiNWaM6Fdiw9f
OZb1xnJf80JPaLu8UnCAXONh0IHaEG9tWhDrPY3hODUVtB5PmMvH4hyjT6zh1fxB
FdfDXnLnIF/My6qfPhXzvmZ6BZ/MF2UXZ2q98rH8mdqCMrqYzBPgLqv5Yl1VF3Ob
HyhiCFf/+37HMb4t9FpVQXS54Vs3TGgPP9AmVCHxypXhxQfzgCrqmaGcLx2rpzrd
vQwvzHZgRkOcwiQq19brBPwtutizOqDFoMUdJy/jXxflHrATuznyi7nv0h4kjJg+
YhBui0+sIKC+0fLdDJCEFvT6zHAQdaE9bTslJG/9Rtfzw+xYZNcWEKkVDHTxOYnq
jLiPKrtpuPtrv5Agg30ki9PsVTx3QeW6sgC2mc2qlWbhzSXbUIM/aVnA9fkF83fB
CkwLubgPVTaH4qGA0xv5gUYByFCOXjD+rjYf5fttu3/o/3jkYzLDg+t7gY6rtbXi
MpcbfNTeClbckqQCJOeXupQ/7yW0/3v4uGD92gz/dH0RqcHVNmcaf3MOBtVcf+Lx
K7AMVsVqjzNRq80PF0i2A9948xj+ZOGonc/IAe2wGMllJ2/NeUaHuUgHPpfrnfwD
ApgGZdzYiW0AnO4/nCruNXLLqZZtD4qr4ZWWqFIIVuWTOgDyXvGqeuDaGu98y8+p
Nzcw0I5zK9ZKI+OmI+06j4lO9ZcIkXtTew5gAHHCuPT1wI5l9UOpv1wU3K/bwKgs
ONFEZnkW5UbsDjjsCqHDnEsMsUOqHm8HZpQlyKWNRIQT7OjWodPbmJbrJNIvGcCd
wgIIuXHzodbL42HaGnilr7qFFNb94tZ19eRPVCgYPcfAV43Q1WUNiqmRGzPWihN4
jP3mrPjmZZ/sqv3zcwtwr5JO7r7m9BS91iuws4MPhimTXpjocGGeO4kQrlSiHvgo
hOHxkURDK1EPHTlvC+LjevNzME19/+4osFrWW7UKstL+rfKL0Osfr9Mmn1lHXXUu
+lryi1bDhML1GzKwV6ElSAMz5kmrpM2puT7P+BVQJaGkbquW+iUvmJT3O5IaMcDs
9DFaxIzVaEc6eZhvNodl3xscTlQY7N0inO1pYrDMOHQNqRVB51Ww+o7ETCMAJaLc
BkwrRZibCNwv5+YT325o55NLEkCnAvVCmKhxjEcfuus1fEXLSiwKl22bYTDIHSz6
56Olnpms+11GQAsKlHjMpqztQUCr5R6upiLEJe94eRfKCYBCoxgptlX0UofhOp+J
WFWhxnBDDu6JHo20sEw6hfaAwradkA2wUSeHYe/s1rCDR6/7HrhRhqqQTjBLOWZh
0q4c+S2l7GO+B8lk9WhpUlboacng6yfw1M/obcOAeqh+C5YawfI50RJEHPJ6z7q2
ifav+WFH1JFjJnVgtPS2x+nsTdR1A6n3MJPAjjXpw6cd6dx6cKjncbA+/JpP+3zg
QnRYb/L+zxhFQAg6009L65LPZGKy06/3Pfh+vG0/pN9vJgWZpKMwDatel3TkQF+5
tMFQFgN5/m+oz3atrDAGFUjgAzi6Z2fLakVVfBBAikZOX1Vwudnh+cjcPQMIA5h3
/xMn1jnElJ1Tix/rfrSotki7/nvsp9O89/PsijThExC+lkXEMxe/DLo6N+921hyR
m6HLHCvvmaN0oTBgM6D4WWIAqLMI7kqVafHwY3W0a167OStgchyRQdETRdm3YeQ/
3xboGGqRmIiybpH60q9r0X9hG1is7tL3ldqgZBeo49OFi8NYErua5cVKjYwIudss
ljlIuIetDOuePUUitJR97X/0yzaYfALrzR+X+rcGNMY3F+B17nYtFwT3T5XhHoUz
a3NGBbKy5Y3vzFHad7Z/mkuLAxYD3WRXABkdMpmmy40lZs2RaVXyivJxEmS5+LMD
Pkk0VUMcLo8/cr7Eho6a8zTvldG8qFbEou8Koz22/+Qtk9ZZLb2Dg4XPLZIizNi/
t0CnHwXUhO1igZ0qahZ4QiQ0yxnTTdVuOoWVVCmHHI6po4T7jilHZCqBBUZ0+3pj
elISy6pmhlRPPcNAWt7J4urwgIh/eqr5AkYzO5qVemeCS0Ap1JHQVKt7O+uKGpmw
uKMgmBPUpdRPLqT0SLChfNXePgpqonaaAsPiwsqygfhQpjggmxX6meoFfAZbvxvf
hCgxgifRo6EsDs2CzX+fz1fEp5UX40qYOpN9EBtXZj6P4d9Fv+UVE5CyMhUNnV7j
mSWgTZURkIFLG/ih8Hkyqm4kN/hBbdIXH8zAIDEtcyfngzvW3HplJrsi2A3LcrG2
tfbBp9zqkkP0//dxnc0nlwvlGDNmbT4G+dmlhBHkHxtB+AO51S6VzCjyiWDMCBwQ
rNXmbGfGC8otOlc+VNSUXc1R+bcO3JRq8/RMI4xQ6n1GyMLN/bZVlcjE7iK0lWSO
g199eiadI1ryruVQ2FSQ6mCGQtdmQ7sJdiMz7qCL8FzHQB7dDAwWRN+MMuZigv2e
Or7+BxtJseSQPI/8Tq8oeAxrCu087zT8/OX6pnOnKqDRRb6pE4cyi2yCTrq6urYp
ZBu8KzHvAQpfD0WehDX4MeM4lbj6bRqBKVyUsXquHTNpGHngJifDEW/D9Cx060U4
aU8sg54/izcTnAWKl1ExGvnhsI8GsUkjAQjSMQVBcWoy6Go8/xVnDSSgEweBri/E
OXPqXJ84RtqOCwb7BASZ1uuDKrPa8hJ6Qegc1LMnTvJaKkFlOJSVnLSZKIS9d5TD
9NtxvN+jjSg0MHPA6AzZJ4KeM4l+FSNNmA46gxjWZL4XjW7d2bwKzRR9NQCSopkt
UNZBCgTU8MgO8boEwCwOoIvIVY6hBp5GPm1qCX8WDQ6oQUAJV5HKQoiW6dHT/pdg
IreIT+VAE2aeBaveQAP1SAjYCKnYRi1Y7Wx0QNtMXICr9WkBqqt2cJDuuBC5WN66
dq042gyhNvEJbtTKP1nhXcq4UKbP81KOeXqxj4JyuPZ67PmljfPErxOJahttg6//
/001ABSMT0atL0HCrHRn3P88yUCX95Ymo760lN0NxY1+9rGusXyPZHFxAz/mamXK
a4URSmlUojuhUAaoQWnA7k34SZ/cTQ8QbVVSkqJLyoAMGc/E9839iRMh5sBCHNfi
ySddQYXCoXxbV2G0i99RNzPm9khJ4hf++YWyDNXk1TRxTVdfLbnxQJryEgLz/cff
hqbsm+D+Is55pCY4eU2ljhA/dVDRkF8Eid3srLfr+Jqq+z4Ct0HDMSYEdnmlF++A
fNDZvMc0dhNb5bYNldnWF/OBEyhDA8I86gl0QQ4lzflepL7286oXHWZUsp8C4cf+
bqedLuCv2Zpv6qbKIjACk1STDfvr1E+sMEMVXuRughwKWtn6JbN5TV4rWOw9OIgI
kHeC0q9yNnm7uHOivaQKsTbHnLhThdRe889wL1F434eMRory2/Vk/vw3ga3BV2YU
EO6sIob3+kNfKl+atpXpeZbD+bra5xzoBoAyYLBuSKFbfYbqOsFML2tmZXRu0i2w
iwjg276px7ubf8U9jOkbI/m1RV6znhuQDv7XchgVMrf7YsUgYjfmd3mNTWsoT4Ib
QzQXudhJbcQtK2LIjJUEx7Pt5jmqL6Ak2bboSYTu1FPDTLmKd8J3eJ0jOQ14AbfS
Y90p8g/Dyd9EfD0lqVrj3x9WWMI9a+zCDArVoj9+2Up1MVZWGi4hgiMwFplSntHB
j6viXBpmtEWrPgoJ81MFukmGyVXdY+CO2EAZGGkazRk4vtNLzkcwf4yB1nKhPI78
xRLdfVFdYq2AVfI/A/Gdi4tKJjblqFFc4FDerm2Mg8Pzmi9RRishmGRA5tvkR3Uy
+pvl3jVbGjOpVmaFs/6XA1AkpF9dWQjzZe1g7KxUj/gVGDvOZqgCsb/iQljR3qvr
X2BWJy4NkHQm9K0Ep8GlI2RUL2cs3amXWfR9eR+CdOGj+a0NyWxjbpS/SidifcyH
ZAawqY+gq17EzY4KWuVYZ+ul6B1suFC9mAp2aXa8OalltxoV0ij0aU5UUKOvD1az
HqID4PZthCfe07UPCUZTlHJShHmcLFBOLBAN/oVtvxSeW4KVh2npuxiop5i5ruxE
HmgxPQlcqxwdj7wwcauEDODobGLBJ9HcinZW50m72f8d5b1t62VXkoTZAw7wKD1Y
v5mh6/TDjdnIUjBLjGdV5VJWiQ89d3KD9sHUBnNHvsFA/NLKfyJ/+aDbOs3Q9jDV
lm2QkaQQU9feleRaB7yQAd/N2CVrHuFGpdmJUIPClThssDC8mtWMFK67gjYOyiMs
cNdzs0KkBRfcfgQbIQOKiwmeYl71HR/bpFroZF4bQ6Q1ix6BlCXZtWfqX/MITV9q
+nC2ZWMPo9VKUgqUuuEyqC/rmep+wC5ZVq8X0cHIGrBZqUUpch2T88jAunsDDoMC
04F4S8gUDLC5P0q70udDd9Fl1fM4HuhfpHGjr5ALS3aqsJQjDxLtFfFSNYf5mZ9y
b3/aMtG/QBM2TmdjocoFPlNkATywDVnQnMC30d8UOtVb4ED43aA75757Td/z41Ev
0BU0E7tgFIM9L+5v8xXeScDGSNFaHu0hI3EyBpuvseoK4X102parRiKlxkW44Tzx
4sQnQ3VW9SpCY3ridKrU6BtFBgUDn5s2F5omEdAMDq+99p2iea6FVwLzr2k4cqCr
g3QEVAlUCpMCLhoRWwHlbqgojMZEBCks32RM0yxnkZFeC0inwfZdm+FBm8Ya3Zuu
1gLpb871ppehJ8ueUgAINW9GvNRGs3kW41C4MkiJsn8VNm1aVff8F76KtCJTVA2q
vsvhHgUhIE6w53MHq7SM1euhTNxZ+wMQNeNPOxq2WuAn1MHWPqTjKrXC9NSiV2it
EDTKIqoNbsFZVgTYkl+N3YgwvQ7leGNFkS9HtS1C4b8jZe/DMSgG03r9E327ndq5
K8RBgVBfCows9kdAN8L1Y80jJRLUxyR4AgBy1ovmEaVYdfqB4WYJ/nvJDfOvIkGZ
EjX4GPLs4P4R5cZPe19Z56rGP+JVTAFckqlBHAx8fJR/ipxyLRRb8hrSGhxi1TXX
nwyO5LzrpZAb0loVhqtdXYmDsMBXyEfLUlVqRoCPta12ubW7TLwQvmWm5Rbh7Jb0
6r73UQpodMQ+uuBmNGU7NDuZzv5vWdIdbwRutwl3FoapeQlsqDmjUbkAKLxn517b
0PigMfsSTIbpV3OiX1CAf6FRdsOA2LsZbbqr3hq0rR/6yp6fYaDzTqtOr+6uLLsa
NTkK7e5lLgxRN/TqVlYbB4M3MS9nTJTViGC+lzEzm1rJ/fbEVuXdtxuVF7huon5B
XwBEr0OP/NbhsBR6InIw5ej0RSksbk+Ap/yAEVLOHh5IC0uSBTjEmdC7h+nDBQ31
2LNKmdMgFbAVgRIvH3ueja3LhB8rJstpcNAfM3I04wvvLGalK3Y3ymTuot4OMxbf
bnSSs7p2I+TwMufIw7xzkCuPo94GwNNHrmefvJnpAf9B02ctLK1bGpmbCWMEPZZi
yE+vE3ZmrYzdc/AqW3yo/oijQbnzquTXFxnvjz2iE811SbhRGE0Rlp3TONt3jGnd
yQRTjBwD/An6QzvuKn6oDQCcZMqh8dcLBHL27VOyqLRwE2Qa8iVEWtdptFVhAhnP
d2fPqBiMvZGzSKOrvtjG2wHfQk/vzT067y4ezR/cjwA73g+tgVxzKo63rKaDT2H6
4UeqoDQcblBjafulWglkg99flgPuiMmlDgOWd1CZFoNOfChjgza6ShqE2EO+lg/E
waxKWGZL6LG6rwIaWJOZO8W5Isv0rYcXMbK+CjyBzjAhBDJrH7M8Q6RwcTio8BaR
xfcpWu1fgEzQVJBXDO3oK1Hec19ZkWy9NIfZTr9HFguOWGDvenUUpXU+Cx1FyRKS
xwNQLRALOwqmpIed/wgxs+cItt1udzkxL/pqHlZtrQgAmzBo/78auyfFyZOfApKS
fq+7M+OjIBqQYD9Od2u0cmVHQ0kTg6/duYpU7shwoJwKnbvLya9waFo8MgZlJPMh
fWqWpJ4AKPd1EvrDDux8bjuSqUvkW5SXAiC1vFCKzL/cZtbaZiwGryosUCh+G+82
bH2tDzvfKkLFwhxMtdNzAwd17Yidzxc55kkFZsOfrYFhYGZXWRGzWDX+wK8P6vPO
PueehBjMSRdpTcPr242MIGgiQ8RBkvCB09Ea/Ek6I7JCWWr/xc72RdjA+G5Uc1sy
XZ1yvVNEx9GxHR+WTVyTT3YrF0ssadLPLOmKGJKLOsKXpII95Ndh4z6V2Eqms3zb
Itsc9rLEH6iC9wGgyh3QwMClTjoMzyZ+nXvYsqoij6SaItLiBe5RxYVv7CJFkNNq
XtBVfRBnYylEusYNllL+SAPJloecZqctYQuIAVsL7peExUIsMohjFKBjdU68BOy+
of6R1yiF9Bg3UjHTwVsSrrsLlIgXNu968X8yWT+Bz4WrKUNawN9ROI5h0zATXR0u
BsRR4CEQmQdqXk6oyCW13gz5h1f01otAGAbRSG94Xw9JkKtfdKCUFfApuACs2y1f
+3Q2Jakk1URA+y0wJI09hcJhmdhJi7hjO4MzCQX4LuEVBWtt0vSRWy7KgqXlmPY1
WVaxc5WXDF8mmjaG+C8rhnGvWpw0VOHr1b0eXYGcuKmBhlD48vzNp2WwfS0yM8oc
lM4E1tqdOVA6di25vRm0AVpHGV9cKj2+GvCXy9AYyZhV5tu+w5a+c8Sj7BJGRetV
zS7CQasQzAju1HqzCTQL1CGx/7hBzzrz7x/QgMV2MiYLNNjRMv/J3YlobRt0Sys9
03NU0Ok1VS7wZaeT0eciuZBz3ZJC9mjEKGy7Em1Slo+PQ/3sL3PCUZmftOggFFv0
FS4eD65Nq7CefPbOwyE9f1azgyhNF+/cMf+89/Zmrs0cMFqHRG+w26nTkhWND2uE
UgZiiyRSwTLZTDUUx6t6kWR1eRdgKspJsaZB/ZHEhyAeWwoL9HlLNubwVtI0LKqE
KdEWyDhPqcBd7cC2dpWIB8JCyb1TJa/SZW7c/MhTIAZKTCO0a6VvRyzxdM+tydFB
2HCZKbHZbrOSdxASIN4Zrey5kTvsU/g7wwOZ22AqyMxqQVNaQWmrt3C7xRmBa9/e
jLhA2t0CBBkKAizpRa2bFxuwGjBs/TsQ8YzCjz6c2fexlFDfGynDhPymf/eR8OUY
uCZjOB2KoTndTZsye24Oah8B7HhvQ0kBFQNb6UnDyJMGYaG6+SxO/3PxyrBJZpM7
CkHCNbjY+iayXSe+xZ18JGdJGseMdE1SE0qQ9alNm4zS4jdao9lr3Q9mmuZxN5VH
8MGokQ0nFGN87cq1hRt7/GI/DaxA/eZy1LCcg7fqa9mwUwXp8I4aI0UhNxueBdxE
U/r4aJ8etEBT0KPtvrSiqYXky+46Yb2TFNZV0SQvZy2p9wEg3VNdo4J5p6L6OQx5
Lvw5Y7S7xzeutZIeJYh1w9yD7yV6iT7Z8kyNS1+BkJUvoEgw7UZFoUbk6hLTEQUe
9Y+fKUwF+5Wcom4dDKSlQQxzZBGl4r/yeiUPsnlGXw3gPVZEhzGhcGLKf5tSNQcS
s3zh7LOqz6wUU0334Hvd2cgg0x2/mmo2GKP6ECPDv5/v3oDs9mPXXlgqwMf8Or5R
Gz1+RrjfPMRTL5icC1LEblEiqt1zHc88Misso8DV0LdamxjifNubWpNXnUivQ6lu
AYIEOhrBCksxyB2otSvyr5qep8//OFpa5/SZJq4jDv0y4NatYd+NYQLWMbqaKbNs
g4fOOSrFB8naU5hDiX/uBg/rwrk5WaC19PsW/QV1XR6xaca4Krr+ckzBCQvIQcPf
04enNflB+midsA3u7aK/AJXfkZHDR03bFM0RLiAdHrsu5QPq/LEMn6gwzp89X31e
6fDhUBhhLEGxXqXuvRV0qgUMoP0OqwuPcqFv19vvw4Lp6B1ttOPhjGO5t+WDmpxQ
r9f85TBO9EA7GQgqBAjpYepdbvnAKPc+U2tsP08BHUs5TkBu8cK3cXomaYHk6/+5
SqRm3QWnZoSVhK0yDjYSiHXPVhbHI4YxxzcN29BcUufDxADcgfIDhOlwX2tbuAGo
OWEhJdOJGR9LZ32k1NcRYydN6z0Q9Urp7VrB8hG1mrXn6i0X+QSS1KWE4r6jmESa
6Gz2etE+HgNzYde3xPss4jjO6O+UBeQK86kbJB6hh2Tx3tYXwqrpN9x2OvN7tfqx
ePqfxy9YRFEBpZ3JNgTUM+abgXB9XMLjeg1BLKI4bnRBt3HgBukHg02/IaKV1QCZ
khtb1XgLKicF4Qlb8ch80x4Hwv2TpMNEDdyjQBADCbHzTTw3wyLr1zS/+0Qw35MC
UeqOSAvFn4SIBUb1GZPNbOXv6KP0ym0gNp9t6kX2eKHrARPHKQ5A+BNzyvLvHeBA
qZb11ZGqAf3uHVAtwJYEeglNCBoY2vn9woIWtFX4+GB5I9WP1/wlPwpJpUegLxuj
XVSGh6lfoIFByoIJxLFl0AHkYwmab4+PIZIexQdWQ3BtHGzdPwB/yTiGnqWgvOQP
BIz+qw/vzxXQhJIhyIUsK7AsbkjXuwzSVmcry6codQvZqCAoZ6lbzvlstEUvk4By
SSxWtzPSUND9/Mr3bkxWLEOydGm90IW1v/e2sWp8mp8TRhDwuv3vA53BpnSB+96p
XKQediCq0g9eiLgsnG9jb/bTZuSETwRiDBPtDxDjPyHi1wH8fKSXLAlFbYzhQlC0
82h5l/jpEJjc3bzIiqWl9V7tt+iAMFPCtKrc/gyM8ZE9J6C0Sm74UpJ6XXvzyO+7
3YePApzUD/IC1/WAzPAscRiybY4RXORKOQ+nZAkwU25Iq6oAhM5bPOZySH1DEgY6
nSx2hvB3T2YFztnbENlc165QBy3+E6wK87Gi4wMX+zWKJjCvcHZv1Eu+DprgKb7h
OdRR/NMzjD0PEclkdTyl1xTY8McXqlPZO9DCAd08eC7MAhMZ2+OFt6KJjsZPb65p
TNJV/1G9gZ4TeZi5lA9MNrBYXp4GZ0eiByB/oViKmS3ZltOd3GgfjsRPA4fiMDbS
L4LJiTgi40ehap+q9rNzuEb0pObCIN+U8A5DUQyRUzeY0ZyhZhpKLGLCkTHkUzB3
bX19DZL/t3Nn428xDO25M2e1sTJRmYsQznVY24oOVLd53ycuUKv/AHS8rW7rH6cn
OmnYtDQ9IKQWU259YlOtnkmexmPEDt5fTEIIIPbkeDSfo/PMXrqGhgYpcemc1wnh
AFGg/Ck1VioJB50MHXyV9XSg5U39v/MOHkS/10Tc7GeGps817fjSf+QoGrRM/EEH
QYBiXhksYUeuAzxb++q/iJi04ofDq9Rb6BfOUu0ps60NN6Vpd45XN78igpXODfjO
`protect END_PROTECTED
