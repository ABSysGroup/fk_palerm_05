`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xDm/jwToZ8bobqqwfq22BDrtpxEFL0ZjCrXFQU7aHi2PEkyTRQxKm1obI0hDQlCX
HkjfnSLWZf+BFGLfEjJ4pm9f5nnBFgugmoos16jaH7AlO22j2QDNDxF98z5z1sAK
IdzMykTY+QVVdOsXn9fzlMmGU/VThiBzCvjz0UQZDBraFr1jkvSev79T8SEjSEWO
BMNL1tc+QHwVkqpP0QmtMcqapjVzTOnuZyiZiF9GlloHlFZFAPPagMGhU8SAIf4W
220g+TCC3baBNvtbyLc4zv09oYVQQkblye3AG650lunjve2u5aXQlry1Ey6dqpJV
0zhVEsn5lI6P8he6vUTOa3yutw3P6UMN0rFGFP4ryMqRj16Uwui1eyD9tmHVRRI3
WI6jQEksVqUv/VrX2Wwod4gyKg/DjCG8T8pQ8e0lID362Hs/Fj+kiqsvzqkK+JVe
P/4zsF8zIDFPQdTW4901gvL+ypwfw8suTHwC7MrSe8us0M1n+6zt4T1229cpB63v
1DI3w7WMrEM0O8qUTR0jnUVejvKUyot3zy/sPSVm5l/d7voeYzDZTTGKiwDzoT1p
ArxBqC5TvfuCueHvkK6WTqWAntrDDFzP3Y40LsOaYyXKgDVPJei00Lc3cj71ZRZR
jAN1xSa/k6Mv1+egN1CpCN+xwEbjx6WqrJsSzrq/aqGd4ShRyQMFkon7rYIHcELD
7z/LT3xJ5jIQUMhu4NTdZi49aHCVe4PGuNv5w7fZQhYzOhw5jMRVWe8GS6hshgWr
WFhNi+/XAcixU1+TDwupfg==
`protect END_PROTECTED
