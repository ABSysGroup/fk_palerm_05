`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wNQ7IWG0kQ/i1PRewPCJuq8RC7Dhlpato7aznFOxZSDHDu5qcz+uHyQWjib2qcNl
S91MnbvU0uOvh3w3RDH8nRWuNXVJXvp+P95WR9SsrfQDei3PMmqYwTerqcFqaX2O
xxcG3lO+KNWfVOjV1rKG1C4mQr/F4ya5CM4TAtI6OyCj42SvQr/45okrRgPkTJKI
+bCiesUZRJED0S8g8fCd01Bf1RUR5MzXIfA8LK4sOlb38N5FCIdpb4X3ZMFwx72P
MnLTHKIANguzEEIT+1vguyD/fQr+SrxY801ATk1KeSQmbIwCCakmo//l4cH4y/ww
Q9EC8Ggj3pFPZC7XWhdnQ+Bugb4gRijfKLrbAvUQ7gnigXYSTsyBx0/sp9uFMKlh
QWOxM4spmWeHiHEW2iK6IHudSBt5kWo7gWKwmURAjOvv3yUTtXcy5cGVwP16zKBk
/8Zymf8eJX7+HZPBtyJzbE4x0jYDxowXRGJ83/oXsCLZJKGDx4eAA+Nb70/RqXQA
TMQJ69CQD2Uk8RL3PAekL0Xo2xnPZ4bynRGvZRCkofBbNH9Hxo6DR2h0W4lB5NV6
SxMI57hHD46Vypxsc/vtL5VHpUnoaIBOi6eeXcZOh5pUGRU3pBJepFCPMS35g9Le
fCmNcX2cxSSIO1OuVET1JWnj9cuhECzTbk378yFoBBs3GND/UakrH/Q0647RuIYG
0mVpIAdvcPNnzxTYSS42LI7qa/bvpC7NdW99GAo6JDrSnYKbEwLjuZ7b/f8fvnOl
CVLUfLhnDcAwR0yKfPos/Q==
`protect END_PROTECTED
