`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IHTVftaFgNNDkhHUHe8dZZ7tjtFYpgCm4natRvNtHCqY3QKuuYa/SNVbPWFTpV0p
B8HQy/cwuGYsLOfCh4zDaQnF7gZ6y4XYT6AFm94qCspus6gBvUOoLK8/KFlK6jBM
CtYdF85kdz08GILoVqyxfg9HTPhAXIecdkGKClRJKyWKEadgsgD8E6y06u5zWQxE
R/cbrAIdBneMZShQRLtNZpaHH2+CzTg41pN83twsevQsIDVu7QWQI5B1q5enDsS9
WpQS56qXO+Pya41YPtDVa1JeYXOxmnmPpbgf6rCxNIJaVJVPa9Sa1QIb6AKTqDTC
XOsXxucw9sCE1XrYAIv+wWhNmeCmumrZ70u6qw1Oh2qhBKYTfoKmdytQVIkFPusv
0Nk0OBaaVHpb++aKXTg2WPTrahppylGK+bbB95gdZpbAqqi5z4sPNJgBLZzcr5UB
qBAhgnEeG688hBZAkFZ1lWAr2zSyX3RmZRjwxF3d1dHQZ5xyOuy5YY4CIpYcjfGq
ISNgJPf7kz0bRIXpIJHNCCGQrIr4E9X/C/rXKqQw3NC4Xs2nF3hKHmaZspF+F08F
nZOYFwjaGbAl9dp4F/dLsY1kix7lXt3FZPyn5CRUWJH+UGmDRzPTK7lssv8LFga0
UoCsetdvF+S1xykExi1+I5xlDcVUiPB1EofaSYe9IRI=
`protect END_PROTECTED
