`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SnrOsNW8mq1iRG3wUWjrzj5h7RIhm6vous2ZpJLCUZrbDgIB7y2N8aX51tjHqWal
e9GPE9qGWReqDTU5ejBX/9ukWzzbveKArYPw6P5NolrHnyqhouqxvjybCDAIM3iv
6SVuxaNOiKnGB8Qn1ROtoOQJhmPLXyZnoeaPJXTeME9aI+Cnu+Rk1oBfTavfFc9T
/lDxmCCDVcwi7oFK1sMS0A+9Wq0/BYSeNNRoXLq2artd08HmCVCHw2xp/9TmcadW
vn9eFxE0RoGyrTng30nMHQ==
`protect END_PROTECTED
