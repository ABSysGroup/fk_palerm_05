`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yPwtdGDbwhBkkvSfbfzFOilll1DhtMs/CpPwf5urR68lWECGq0xtFIppe42kjg2F
cCJyOtV7wdj0i1H34dq93lGGTa9o6vjJwcXw4t4SaCxwpMum2IfHzzjitQyUub8g
KeRw9z0VS3viqiMXK/IJA6ih2pzosqCUpjTxTf46YklZOPvd9g6hrdqs0iG9UIbs
QXRfZhZTQ37XKjclBIVsDTV0+bk/8oSeUYJWV17c8AXStZ6YALXWFXrMfCcQD3Gz
jZMNRoEiE71PvxpcNJVlHcx+LzScSA8U42ix9Fhw5d9D9yFar6yVwBNljwuJs7oj
KnWBPg+ch29j9zu9rlSYbEw6X8rbTfmRjLtaItCEspw7ewM73dTW0u15Gz20B+j/
JqIrk/oAxK4cJ137dugi7lXbMQGXsDEqVMjrSBwaC9eFv8aCIX5dSuRBc2ThTqhM
JEN3PvWWex/E8pjRGeR+qCDDXxjqJdjjAcVpH1nHIP4DXg2SnJZoAM2/OCTFvtcs
m8swhjNzvueJBfCSj1TnwFQ1gAtzDfF1T9tA+Jk7CuMHBoyzryAIIosVosDPw7Cw
w5DM5T10GuxkqY7XzC7vG5L2IXhHtAWztNzW9a3GmHqOJZ9gWRPwfN8XLEDTyWuu
BdHWBP5MtYcfPoR7QkaiQJGtHJyyYo2JCmGidoXGaeCByf8Xoex0bq1HD8JOZ/I9
Pglry+DUGvmwc26HRV7YFqQq3pIkqaN9tp4Ly4TcXRcZeF2rA+k7lsENerdOfBm+
O3b2zSlI7nXEkExUgL1fvCR0ssnDmqy36oWVQ6w3LgIXJv6YJLXQbTYwM1oyJHOF
pO/G8oGVXQdSQ8HTfzj5IuuYOQQL7dnv4saHOLWDgymJahmgZFs3F9fwleab4xUo
s7wKS+lUQqpWWnZD8RT2tey9PO51fvBkIXYZFYN3iKUGDGA5gPvbR/Z+y+MNQGL3
4BLTjNpVdZiOiDOedPztFi8ZAFw4eNldE3c3xlS6ia3RJWHkqst8lAXb0PMt4u/I
y9v+ev+j/Tbtv77PRypj1afPTPkLq+syQsVJW1WmUH0t0GHbft20ZhTIVlRk2U5m
W1whkLWJkhnEJbTC4w90zD+eF4NHrB0etDPMdOI5uDn5Jax4bqkhyKu28y42Admb
zEitQEBj4Knc04+me7N0tqaKhQYvmchvyCamfSy6b4ORHQW+16wuJTaOktGqZf9k
VYlkH6RR5i45FQDRaNWaM6nrJUjbBKjHaoxznia4Cpf9uF08JsdiPb6JBOx78Xsa
O5IJfHzAQFQDvpXQm1Cw253oV/Yj/ZYzM0On9pneT6xwYR9KdUWVORadCwD0B2ul
zLzF5t6A+h4wbOhePYmY5dlXjEqz9/SLa0aKq79/h8J0eS1MxesTd3XH1q9/T5o1
`protect END_PROTECTED
