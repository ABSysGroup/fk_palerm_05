`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fz0gLPz95ur5tVgYuiKzbTkF1q+zyc2AQwAFpmscAK6OLLigkddgpKkx8g75S3+d
UTfaA0Dd8v/PXrSB+WOeuDFLCmagYhV75S+qMskvgwBil4VX6DgmwTJ6CvvcQy3j
3KVp+gJ6b9vNpex1eX/fs2n2oB51sCvaxDgCj2dl4zkTCae6Tzyhm283cJG2PnYF
CkEMIuV2bXljjvAaDafdXDEqwVgJVgCpUCijGovzvx2SdAe8k0qN3TEkxmiMsDp8
L14Ah5c+poOh67PvOuuo8toLQSTi+/Wz6nn7+Ytn88LlP67NEC4vDJ4hXdTSRMLL
I2NdiVUnEUnZ3T8SnuEFx5yuPWIQn+FXx0jP9vD5Q72t4m74UYje0evTrR/WdVdc
2E5BEJNLvAFqh3esJ/crSTbMB7SxQ8GvFK1ukNyR5BMw9696UXWIr2OWPf8XeNFN
jjDfF3hx9vhqMwc14C/vevcQC0N2a7lY/ysSMMIsx1roE7fw1Wps3J+kwxgeYpwH
5JTsZ9DAI4vBxe01CXW2zz3XigTGZ5VI2vn5MpLlUhr+MhrdEkeXto64GVhrl75n
ES7x+cy1TpETGfyj396+UBifIjkL8Wz5HCqsvXKdbYeianpJK5B0DhW9PIwhgk6W
qePrFWAcTfgRz8zDNNJ8WMcTeIYgBf7GV3EL08qIj4A=
`protect END_PROTECTED
