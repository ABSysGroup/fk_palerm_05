`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qepw2eYwUCGXCQtBOCDfUMCTVZ6Ci35SnFjtFbasoy1xZelihc/HkZJb2ZzgbKce
7X6aafYpLEXfCKtoxx1XP8BbnrLg7tHHy/mwfmWUQ/544X63f0wUrKtmDcQTXWjs
hz63/L84VlDD1nzKqhSQnTU/qMpUeuU3sHWMr1x9XbTUZgqksixEnPsHd0TodX4y
5I2xx6H+6fqrkriPj3tiuEQ9CvPs7++OFoO2mk4ARZdBvavYu/gee/mvPMCpLV2I
`protect END_PROTECTED
