`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d9DGNQAn7obyS+rf64US+aMLMAO413cjJpsgw5HC+gJN9SXpicEuLmm6+sdzEW/z
BvZCdTFY2R5uVrxrW5/J93vtHIuUmE5ZaECstcIBTRifV5aQyaEEnOEGhoMfOQYD
8/6HZwDmYuNkus2JsGD43qWDCkVaQ3gjPKvOwZAC0YKScm0LW96FC2Yyc3fUl7Qn
9/uTeNxVmPAe6XPRQLvCxZBQuQWTBBIHnLi9xXXU6w4WtE7vqe2TmG8BCH2LBNWu
AhgE6ft33eWXrebzFNSsRg==
`protect END_PROTECTED
