`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3ivoPD0zy3bG2RrRwlOooJs7HtH+Zn5HprNybTR3Xv6folUoFsEX5RX5/iiwVjka
NMLu4jlPDFYR/LLuuCkCScsu2wVuZ3qomwSTczp/dNM/NyzI5GOwCMLsbyEdTnTe
MbaWW16mhWDMYADUgAcshNZahQXm857+LldmyhN4ZYycimaifzSMcl/VjlXHBIr+
t6CbiZNFeFvif1yrbVRmqLaeZ09LArqll1Fah8X80OlKIZlLcOBIixGFV7dpMZKz
SO9Ysm7dC4Ul3zZskw8lcUxQcEmGXaK3lVh7BkGv638jTiF1TebU/zPAVLQsX++p
MTUngNgS0bKtOxV4SUJ3Og+d8/K6wCWFyUhgrA3+qqp8lc9ffvmhpJe8htow+pdU
bsnyhcrrbX6/LmV6lVy23C0/Pw8JM6fCPme27cy/5SNqy1GUnF0+G6KMLQjUW/Td
jaEnCORO/Ypmomj1vnxTsOHqGcYQqzzWBN8IkoE/uVDbY5LvQdQ2ovPha+q3h8Va
pK7AahYLXORi+vPgsOVDJ2nAc6N+Jj2Oo4A4GULXIRpFhh9CVAOtZpT7PpXTyEP3
BWajFH3A2Y1qlBr/zqR/4Sanw2yGJGa72mHvpLgDXHgPu2azB7jIQQLCEFx96e1k
VthgIVYJm5fEDQAKoqCfq9HBefZQFaRu1tBbCF6QEHTTXyn3y1JMe7oU8YG+RUcm
QweIr6tkNUoNF+EDY8XiWCRO+o6kn34yiIXi8VG5Ez+PSBf4O+DRrfuLh85YyX1d
em4dzBOSqWOeeea5SUoTT9lwsdDQIrzrCUTOI843D2NjUUPfW4aGQxa9k+NjT5g1
LzZjnoPwEZE90bYM0ys2MJuXXqiaXi5rAFVirSWUhJ90QQ5wM49NJtiI8nzfDKrq
K9e3H6htHMYBy6NUiM8kax+Uq+S9dh37lq+yZga3RUc=
`protect END_PROTECTED
