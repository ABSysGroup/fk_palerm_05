`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vS5X7iqUEJ2XJoLb5Z9RYRiwGK3zqp6xvYVLcw17MyRZzA1TqvFG4BSszGA/+/mI
LaSsncwZ9n9Ml5Gdy86IzKHX8qBeD+W5qJSOxQPb7o6qlcNsyRGmFI7hv/Gfx351
uFj5pDulwCdnY3o8Bwb/OCgpOsFGxMRJfh1IFQuSm05q1l3x4SJ+yrI3KA/oVVD0
uTzH4wQoFJV0Jv7+hAPPguf1b00/2olJZNlZraasACXjMlxT1DaePMwD3+/cJGNG
dEctUIg8eil4vSs83Pj+gLpTZBnCbmaE8GxBDWHusH7vO+ZuxB1xdoVbC3qq3Uwd
aYvj315Hj7KSOjp4LAFnTwPoOoDEMbKK3eokQFH/stYLM1M843J8xWbDKzf51anM
HZJz46J9sRow1dR/GPbfzbn8XaRZsMrbcgPi+ij0iW1BBl0U8oSaDrGzQnON9KSC
tTXN8lBB7ldmEbakreyVkY83dVfmMkONfx+Y8Zb6crzIBaKuuUtxAD16vmi2L91d
ektMlRno5vzvj9PIGTiV60NTxYKMBrd8DWUIIVjau66qQywc+sKdbHPwR1MKsI5O
ZfrkZAiWdDlQ7JSUlqyOmt9DGxIOYFJoOg1Dex1f07vSKjYF5ijsNeMHkgD0YMPO
lHZ99bNEEjHGu+iu66Rb/g==
`protect END_PROTECTED
