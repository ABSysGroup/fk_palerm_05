`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8eLrn6JeqT8lKizrTe2NtqhWXC0T54dBupQo8PZ7HKU6gsxb/QyfachvrMP17yD0
pBzURk5NPQVd8KSK0ZuCe8ChO1Y5fhyz/OBaEQk5zFXzjYGBDU12S6HJlVW+ljvx
D3j/TxWkuomhKyh3q52DGhkla9j0fDEfHVonvU5NBbCgiS8ixzqueDKRtnYam/Jq
8BGzdYbeibxtENVdFlErrMRENNFi5Qz9k88yEMIeIKm0dw8+40I8NgEVfdUKuD7Q
2aJncHUmewFeoMFoVfSV0EYXVHD5LhGeCpIXVTpdDJuWxzPEIsySuDE6JpqNBlO1
PYTZGFteNhhLwrv6vMDF79H1D7n3JM2aT8oVVKMZKy6vA4zXFAIXhmGzzpVcwuea
OFYvKonyyUuM9f5X+kukevxWO6m18wrCs+85DLkaNQ1hPSr5woZcbb93IhYTFK50
IniP9/5ScblztLZsME1gXdGJaiyNnSD5nAdV3M7jaQx/v/e+hIkk7EF/sBSnxlmf
Cw3KUDjpVpZ66cE20lvSUI1NkHHBGYzP+/8CaZj01NakM6WmGImAiUBL0K2Di8lf
NdopCYT/GbatoLHbkYcKqYdl7zhjASJ/ae+aPf4WUX9TPfKVMj5NUlyv6K4L6o+s
rC3Ba/MLCtRsFJnjJgCdp3xO/hfxKTJyCqDaMgK/HqFNZH5boTHVm4b7IeqhXzhd
fXixyAYwtExTbzJBU6NTrvsQtDp8e7QFdfIt93skGPGMArGFcdg7o5wv2Fg38ec/
IV4wJBsAT1YZp6HMtK26UFbX/bcmx2utk5grMitJA+/gS+cs43C6lDvTer2Xn2U9
THXu9Iae1VQuKXPsnZhoy6W5bYyDec6MIYWUx9fTVL84tJYV6dKq6mdLD0dDpoos
xgmtqP+A3Oo/F6/IjR/ehy2lDp0YrjAfJdud0MbUS/n2platEQwsBVSH+vKb247c
8lA9P49VDfGCNG4xe6AxC43UHo7DDeYk1/m83QVdbJxMwx0SfmRZyUFpU4bU4hox
8KQMJcqrZteVbtfWomfMuazbYpzNe6HG5u1beoyl3iPPA0LkkA42NtJNFU40iJOS
nIo7J/uwyqmvXy6rqSfEJwvRU+t3op5IA3RgzEMR4ymxSQ+jVuKVZz2WiL80HjF6
bMxg43sF6YPmXrZPm7cfSllGQhoCE7pFHAy+cmt2wwg/MGTJxj8Ryj9jzYs1UENY
+yxPnBVzLruh4gW6wPbyVSE+9Ulghn3m/XFZwSzn2V86BbV6wDyVElBRVnxNhhfR
re3R+LWpKURUBBKLh43P2ui/cqxiv6L41aZKF7MJdCYB16vFN5QEczmCasFjDMQ1
GnY8UlaSyLGZJD2lwRUjkP3fF9Sb8Z1bkOZXTWAxP6AaqSfIK59tnvnEY+Hab0bf
QGcbVKZvMYi40fqWOr5wBM9kfMGC1S/4XuJv4B2pJZN7NIv7TmBIeG+E/G7iG15s
aP1wOuWKeSWaIioVdGbFkpk78TzCmFhkMupX01QO870BIPmHEyk8JQbNJRxMZSEM
oS199XX/kEt6p8ddvirQaRQc7CxapAUfujNiYxtCCcfgKamrw6pHAIQ7aFy8dnJB
+rsoVsJTjMiQR8twEUGsPwrukYbKO/yZdi8LIEHOG6c2jY0/mXYOejhQNr/8RdTS
vXFmN0/dcCSs8+9V27A0RmVN2sR6ii93DlDZBSXkJ/rDbqGM353AcdF07r+mu9/B
+yk3wYTg/Eqf4p02Pq7zjnGYtadUwCMyrafkZ4hAtqu0gCfHFt7TXT7sSdFwOMUI
/PT4e4+y7+5ss05CNEG++jjjTq1B0rOStu0WKL//L0xXWvqv5EyxhxTV7AX5OtWb
LFMzNLb2HZWMArSNFPsLf9T5IUmTkQHbOoSEkwsSDtfjQwEXDmVTIuq7h0Vy/Rqg
PM2F37lG7ri7++wnr4AVrbqH4gbw5oGKKRK2vhRIfy6pHUH/oUTtAazpJPUkt8Tq
QTJxr5MjkODVK2SzaUugDuEoGST5P36FJNl/OORfM/EJIaGBkWZQpuO90gvhp5rF
/rVw8jjxz4PqYFNO9hKwZM2LTJOLCA/S1da4PdphgFXhy1amEd+mwnQ80VcTl7rg
`protect END_PROTECTED
