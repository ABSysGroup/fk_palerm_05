`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nGRYS3X5t0TW2cUtR/dSkLoBxiJB99o0tAD5x1HFIlK1WsTvKKg4UU81SzpkWWOh
/iLVeHDskv2Q6tk+rO/r1K01kxWbbFkXp7P9klvqzGJYnJNYnMwnVKjYC521h/s4
ORxd7javyfFPt8lPka4vpLfafD51c/4tG3yBPyqWaKrrm1svavWR6DOXoYobgMfc
BHALW/wrTbORv2rUDzR7+o5PKQ0gE1VImLM1DIKVjJ3p1ZUEZivg55bb5DSb2fHV
oGpJLbflToCpKD9I+BgpHepcs4LcPh5S0E7EVBsCpE+cifdDXbaEXuZPr8gMG7hl
d0cNQJIrUu+eLG80T1P+bQzX4aQK6yUwMkmMS8USwjsu1ZeZtKYv1mvdFpVMmVg8
MxEUWiOYOQtlqTPPzJ4OrVRi24xwensOAls2y70WbLFccFDzEnpHPJiDQp9q/exw
RaMzcu2zP5CKOMAu1J3qGiVx0+eqVgwKVPVaPOuTCMpG64FuUMx3XwgV7kVl7Fcq
xjjhbfXD0vsVzYThUGley8T4U9+Pl1JMeaqRDdrNsGGxv3e5+1Md8XEwnqAwVUHA
YGBRtQXe6lTceRhWFfexGpJJgD6wgROdLfwLQrsKPj+2vcVbUKD/Sa7R9BSYgJ9A
FM1+r6jJMo0mrVyiUVYfO8RTTNqr0z++/Q7EjiZnHAlMEOPGG3D+HWmIVm2sQbWf
zSx8dPoGKtpGf4KfNSWCHldiBNDkKsld9yqDAYIZHbmWiMFXts+PyM1cn4yKidEl
EheULchddYI6A2QEeSDrQhko640oxb41EfLR+j5OEmdPgVW0QzAR00upqTjMTMJ0
zbQfCFAby6EAp6+zisoX9S0tPknENn82otL+bxIylM8KJiBEg5zXoSTXDU3OITi3
hBuMRQLuzvCsoQH9bPjNM/59OwNUjVumuyXQHZGK/xKmcF8nAxub86w8L6DZru9l
1EpEw1eRan3iVoLNKAi+AOsMLJLa5Ou0ta8lIgZZuAjE2E01Zr8CpWuvicXcYXMu
+denRuNdvAMjxjg5fsa3YjmQiw42CUTLJmz+LEWSOB3W68kLNwSJPo2kc2sa7+e+
oR9ABFtV7lHV5rzKvABEfeqPPZICt4dtGPOEgjKuh/UaAanTompbTmad4X/ntUyj
fbbp5+U4yHrvZ/fQOzldxJZbOgQS808kGPG04TgXgvRwCd8DDXXqIpZdze24AhjU
UhHQDKHWUB/5EETeYIGbWHhOs51TDJ5JLsi9FmQ8A/cHEM/kW9nQ+3p1zUFmgy4v
QK2XDbBv4nrX8vTTotwuaMOH/iwlW/od88mtzIjkdRPotu/jMbmSbPsH/kyb36/F
4lqxIAz8DNPGIwepuUj4K4bdOWsRNeXPiTIbOGgs5B1QJqRQMTZ/qXElia3sFvVl
Jd7zDBKtIV3I61jkLYF9LNxzpyaakVOgLRACvkNGWzM04LLcIRZrrpcsgGQ5ZIyi
8NWJhr4gSZNXd4p9YTvQgC0tv0GPpCEuq9Fj6XZ/pKiwWjePessFJVZNFbM0XkCE
dEWWt/0+bccO+0p7T1tO14YH2BQS24L9lIuNQ3/bfcYHIdwkTEUMqSqMCMEcn+fm
SwCoBkl2CQQjYgOn3ChBim7x5QlvdNYaqsXOxBsQwKAAk1WjcF4RABeylJ6DdHge
uK5xKk9wvFh8KkpsilckoxhhHzcMg0P2xwWSutNw+QKHu85WIMkmVq3FbDY92Vpi
`protect END_PROTECTED
