`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xDLYbcyfa09FzPQMy0eF2qtLNT5/rOWSw4Xq+tsBrI4c5OdgvcJLMSAp6lCb/cKd
p9gI4fh94C+S09eoCGVQ59Ibk7rIoo/hQphqxowwnTvnMST0y3XcocZDqlei3s7Z
Xs1mBc8H91tCkNNgRz96m4AQcnv6apVqjxeTeW3njvaqy/yBMpaqoOZs5CaB9Ge1
E7xhpAd/Rsb8GaLKaDA79u70zvv5Owovtl5kpcAeZyZe4OtjNO9Spxf4ArU4S/3i
CNq8FI5NU7kVG6G16GUiu6kCb92p6+u0WcG5ZHhokTwRAwhXvVFYzF7rRhEt65s3
X56it1dbca0rf60zLgS/ysYmHfJJbsba+lAeO+yQQ5msQgWjN6YPOrL58WDM6vgN
uAmwldXzRRyUXYoUineqr6usvX9EdBP6Q5Li1hWHwLaeDsbpSDd+f0DoEJ5Ldsmq
f55KRH0oQwSKnH6nUnba5IMD0hzzVJCIKTPerFiwZINNeIj3HUj6pAv1Lng46XYb
VpX2XGynXnqGsIJwhI0Ko6gfltkD1h//qsBeTSSjQ2oHHPWrCyfMTso4elYfNKst
n8Z5Ud9sp7jGELrvf23sES9ap6RgplL1NtDQf1IbaNIzvOFA2mCb2pggTq0AKgxF
JzAlVxqxwgPvsn4MtXXrtiRa5vElGZfwc20LmW2olcyMbG4ZvUWcfpmr3DD7VeLb
keIeMZbWSPYfHZhXouI7wXXrebDXjbp4wMo1shc4hpkXQu70LWEzZIxmSIcpecc6
0r2Riwv8JsDTcAr/eLq519zYgHAgmTK4KO6/lwxOOhF3jVeeFzT5PbpEqWayiB9D
kXjUy7HiJIw9cmHYK+iJsGQlCcx5DP5U0fQw2HaU2fQLZSiJ7f4dwqWOTeZIOahK
R0Y8W95RrSI97/lqyM/MMCRhoTr70CzNexadPveOmcCmeSZLUK0oKmdUWFCE7z8D
IO3XVxRmW7dG28er04HPlMz6v6jVvqqsrD9TjafAdj3uceKl2dolFyikn52PxKyh
7TzQJ8aFA2/rN7lcSXK33UaGVh5U31J7sBcjkwwq2DRvgNB5+BjPr1SjPYga1IqO
e18xJqc7kweSe8a7z0IqiWNj7oQQOnL5iYB/K8h/qawk2GuZCB7oCg3otUuLDN71
QnGsGsE5QqNkW2BGa6bnOigZQswbr/3zaTdgF3Ec8tDI1WyytBrQ3BaeuiwNvhey
HZI0u7vo0E+64o6gM/FIWg==
`protect END_PROTECTED
