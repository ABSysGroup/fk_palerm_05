`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BpWTDisFH7A9jSZY95LsfawK1RNbny4TqTX1S7qNSih3UFoQG5OgIf0LXY9hCCeE
e89KQ2GPwNWHYZ8QbTzuqGobJoJKJomPfiT4x5JV3Rpo7/J7qmHwRDKJ67Eq3i1w
tdZMOZMnxe2SBghNWM0Ift9oA4noetIn1FudO8eSOM+kPqJ8a7AM6g+BePDEa/2Q
rgpMRw0Ck/gGdrgTcABRRtOypdxet2k95O6C7NN0VtUQAr+yZIIjmVko6NhsYS4l
K0LDQo60WwMk0t5I/Hb3RlZEaX/S1ho7YgcU61DGq2lioUNIo8tgnUHRiFtnhmhP
ktBi6cJigA+AQD2e1gb9QrUuzyZaqqcZ5XQfcaG8dHQu3IBRxY7ddqYpDvBIIuCr
l4uzkka9FegHa5MWoy4ZtQ2heO8TSWazVM/iF39OsT8vvZtbdpI+uxeiRv6RZJFc
cyui7z61AdT7TAsH0MBNzJ3oEu95naOB9NidLca9+tdxpsxcBKFkt9ly9MBVqYBy
`protect END_PROTECTED
