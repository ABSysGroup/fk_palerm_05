`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3pngYSHjbWj+iAM5xlJcRFagraiG3eZ8argup9+B+nHjLvL+gm/GeRVvdzYI2h8d
aaCKtKVZxfha0QZRlR9xWZmtLtIgl8VPnhTZ1SGTWZf2y+H7uLbUDs3Qd+AmvOH/
/DKHdRmbYFeYTho2znH03hJnTjwKiknUDpt15huSKqwu2zjA0e+ldkutzE5AjIuL
GbiH2WQ4mBUYA7Ghw8b5uIqEFTGoh6iKYqwMpWFhHIFivChsLGHqS5G2Ocf+0xdG
25TQKx4foitlRlkoMlhhr6JEl70kTV0IKl/SBBod2zqzWVr2AVSfcxF5CjQ/7q5Y
315WC5DVtvDgZO7DoRQXG+hhmQLfiUypJplPTXPGZRWCUbfx1oItKjYPrEXz3Dl+
RvnmOffzlLx4DeKa7LdBbsmV64ZMHbXLGETXAsHFVXIxmFFMLx18wpewyT7AIG+2
0pVpfydBiRbuDv8dQfgt49W+t+0YDPSBsomgrAEwgPKyywehCvEc1eDxbmcZhucF
cCpeqczPK3fi8C8RGyZdLyp/yQjEbRxUe3mXickBJxmcoFmBppsTi3CiIMyyboew
lVWbfZyISUGFwd+6CQXKSC+0mVW1Ry1+g0OXAATuIq2LGyRye3WKxJ11dID/hwGW
783fU9+56wKZ8Hnuk1uASfWd1uB392YNHg2vgPcDvU8it/0HFlMoCJl8j8h2y8YN
HOrAsa1i5AwIGhCkiMAxkIQv/UguIUMetFIQhf+TtRA9YF1/6abAsdkqGkFhpGCO
/ljRwM4MlvYFIps2PBIiCvPVYbkYRVp51bai8cY/FR5xA+douqfCCMlWxDlAUNK/
AqaV2O1IQXHovEvPHsof7u9FBE9Y11NrRamF+gMpDbJD6qOkC4Ek1KiJ1aiu19f9
EKiZCPPR90cRdN0bJH9SFClw1dr4JqueLvfyudIfxDTuNjpKE+NsTcHiU1UuBiPA
Wr2QbFVW/kHWCwPKS0NDsV9xx4xg+LD20Pu+fi0y/hSJQHWw3BpQDDmmguc/4jPx
egzoPQdNU7gs05PYsnL6XfZjEa5Am480vxHYORbt6OBueWVy8H/HTJVRc0WDhU8j
o+NxQ3FnFTixW/iNhNZucXLmKQlDSy2TDKPdOydBmvlvfuglvdRiEh+rYKHYvFam
fXK5rVCr6QbFvoBHNUPOO8AczNxzBBDQHDAuBG/2RzfwKS7QWpV/Ys38SyG8cN6L
8ioxQW+bkvUwZ22Ty8ZVe2GLkp+zt6ZUZuSbYYVmcmnRKLr/NfW1lHZouBxvOULl
mcdpnfemn8KJ8v18fDWSmfISC9I5IX8VJW5ExGqTVmMKuAMXKog/k9/5k3jcQkne
Y329vJq3bUemM4c/Bu4T8ENpPvTI7pEKI9m1nPy96Fv2JY4JhGJUaMeaMA8Y05Ts
wwfRN7X+Wyj+maY6OCqpEo4gibEXtlVmQoz0GdSjGKPhoz/lMdwameDe1U/AcYjs
sa0Gs8iXZto/meg+JuftbbIfFv0dI2Hpn//dheVYUFIXaf8MD3vXC/J7oVE0HGt7
QbZQsJY4I4QblpJI72oxz69Cl5gfewgKaIifctEN5srDMmOlYI7xYy5eAwPOz3i6
IKb6qV8OQJWIMLs+tEqZE2VoCaS8k/yu6L/XWQQFfXs443niL3uLjUL7AsCiXhmA
IiKhybHFU3k0sZyb/nHtoeN4s4e9AMgkiGNxltoRAcTBeFROH3zJiuscYbUX0Ajc
eEKJM49hmyuYbhNohGeSS3CeJD0CcljU6FVY8DuWc2q6mrcUcfJBTiKvO/G+yoel
c7MDzPUC9OIWP2Qb5F6DNrBvVKdtQl64uHi2Hlqb4Q3vIpoCGjfH0z/b6lMxnVeZ
WWY7Z9Chtiyjds0ONhG7prDf/fU53FQxF70gCJro+5LejWvyIv0E0GwPyhDIZfKr
5IlrK0VEH1nI6eeYy2SIWarehWjn9qhHsD44kMio2LrQAcEfrUDbYU6DKUJJtZ/F
bDQmG8nQWKms9DkzPEK10mXSiZR3oPSuw4imJcbZHwUm175BrsfFBviSPcCJbS5S
2cBz8m0WaJ//bbTlCtz7pgHSnxxIqm/+Mqa7A6DrKDvRW+ZecAa5+pHH5BnriF2I
JB/r0P77Lnqem1CRSuZKaQRY0TVeZrlNVnNM8qYcw7EPE1aDDxcopuG75dJeaa0+
4+NPwsbvo57t8CG6KHYykHIzhEukf6m9zQgxa7cH6/EdGY5U3YGlRpeNvN8lgcLr
waBrSHUTFsnecuo5Pa23gmF5Iuhfl9BafD3pFs5KT87g8LZubngjG6k3a/3Avv/+
pi8lJRlMRP8pwc9P6SXRzW3iEHjxssnLCI5VWIo5o/07znMkNkv3s5CkhPtaFb3b
GbuGgb2UKGOAIiy3KvBV8GOwIgMo8tvd2r8/MCcK9JvACf8jL5JmPUA9TXnPf368
o3qeVqlxUgwX6CiBY0r7Dngq7czgio2aBXaWxT1LdZdZ768D3/cC/1VznEIN5Hpa
5o60vPdUGYw3jtr7MvySF8bC6fugAYg15h517ssBDJfWBfwbzNJLY74eNzh79fZn
7nGEZmnewT5cOsMF9X6niUk4VqTpheruQDJ8ARB4iJ6X7SVUpA3PFBU0X7/OzkZS
ARHjIF1E5c8F+rJ3bqPK+T0QLZh78WOFYEClnFaFgcAAb+V6VenNW1sJFjp4AsA2
InBMRKbaj9eaV0TAIOkAMHbD5FG8rVR0+LLwrrb6N2BRehFqT3b559Y4mjjvoiFI
tqh1dz/wrJHZlOGocSyoExDwTy70FOa9irSbehD11hxeHFMzk2hspD4dtipI5R66
8D1oK+acOFePH+OIiIsTc7gzNKrhSNmVBSrUMFViDCDG6tfs1+6PsMXSdq773Af+
edH3EpSYvZ3LwSU0UEGgsXMaXcKNCCId+hxt360x45URkBW1pevo0dMRPGoiv4Og
+ZetYotdPAD+NxxQN8Z3fUe80iRbg4yeE9JZ9Ba2AJRvUwqR2dc95rga8YU0uE/s
ehf5AhNjj64thXkKrupUEP2bBMLXb3f4oaBcxMQ45+eW7J9vO8PdBdgULi7GiZJd
2rdciiywRvRE81EUCf2+Ve7y0foTVmsen8m6mCIt23UBxdczNa2vHxgWG2Jlz9vo
Bg298FtuzEbSAcZoPZexiJzD3KdUTuD/PBwqkWjoxMXMmPWMTuWRgTjTeebCS7fB
TjRtztPkh1K/xk8w9WEfWNLgqSf0URzMhA/MBW9u9HngqRu1lyLswxDZuAuhPUPc
j9xovTF9TWPxe96yYtQ8XLa3RZWoG5g1D1R+nh3mFsMfAz93wWMa2+TincYFdqot
9+NKGRNLW9WoGGQvMuBlPPB36SFVIoNShPcxUeWytwEzTWN5Wee14dEbefDukgMI
4zIfs4NxiZjN5+CMiz4Sxu6scB7FAP3xxIHspN+51TgBxRSyQTbBLWxxAi8DPRqU
v6tP4LnM+h/I2Itn/BXW+8qg/rEyOTO5Y3oCC55tQ+xrfcpTAMn8hoCyZcgAmt+9
QiXGFEixD1tJtaM+/Inam5c8jtmmloUqF5Du2vEQJ+uZ/mEJ9v3QnugsBv58JPOF
DCjnkR9ZPHVTW1MAuoIuqth9FCr1uQU+3ciWyLYgI8Fe0o2umGuzG/nnsNoHDsMj
d/yQd/xAj0BQ8OyKHUankM3o6OzbJ1yG5X0j6P0y0W63EqF24xqc5utD34Z6mnaZ
scTsHqjblV0QvlztGsPHDE0YKkC3KHxCiGgPKmUtkab5QLIzYC6unr1LoXrpxfet
4wTqUI583SXh+SqnDrRs70P1W2ibXn+li0m5N7F/51A1a7UHafYe7jVTCFSz19p3
2d6LvxOaa4aiJjS3H+mUErlO07WSpehfweRDQu4msSMNBQd1+KbQYm5SZjsbJsGn
X2jRnas/VswYi+ybHWd7rpyqY9utJkubMHor7VSnK/Io94hEPsZ+lszzkfH0Ey4o
kLondPGoy0wimGLjfr+F10+fcDf2kGNdm5kSE/Ov5YkL4+4z9yByEB5mcmzRkbv2
T5tUOo93AJvTZwt84em47e4lpxU4aP7IlTuoaS2EYn4ojzwq/2V8ALFH8DBu826t
LTgMj22ZUW8QU0VCXLpikqrpzsXHlVhLCcglryNGz34Lhhzu8dGyRdVsS5ZRlPcY
kY6tcfTNMA+TPz6g+Gu2Cb8n/MOXdAL5AOF5C7q+3mUvFPsPLk+4tdStCKp9dnv+
fUpt2eGbqQDY/LVYnvCKsGRXZybt0zLwEnPyEko5qXA3HTYSRp9aoGfpVGV147xw
2B8x685cOHItQclZOzqCZA33DgzrinApi6QmCw1aGQx1f8Xf1mEeDid+HEYe/GC/
jPg2XSxIJBRjfq/nmUOeUPlvvKLAL7x7J8Z2OhLyUrBUPa3EaEDr9H0HP2CYD5Dr
h4P8Xub9n8lP4hAk0Rv1afVD/6po35lpxHIDG69GofODPPTsOq2/jcnEYdHu/D+B
1F7ZSQpxkLiKjwxlKUmfyqnlwsgHIMTFuuW7k+8hDfYXcixNhQo3WQ/M3Qp38FFK
Fvk76Q5bPxe+R9Tj852tYMf4Mq9DByUR8fHEDEgZIPH9ilmWR/OCuY+/3N/elHMf
1rrVEjTUEjZsMbqvP3rRbuNM5zEF/1cgzp3+dN14RJ0QjVSfC0UKkPnR5Tf7CFPe
dwyxd7lSdHeMVXES5nj31e0zur+hLXYZZjeBWgakRbaq728ShmnXAi6iYoIc+/6E
ikUjzrxXbfTuzNS76/rMBy4ToG3Z6oUhcMQRmEVOgpNs3iMJtIlh4EiG/DDicZOd
p6MMuw+MDLAM4wRswAaKYK5nzAlpYjwUf4NMO6RG7IboBX+76GCG+7/fcx78e/RP
uNa4Ma/daqRr1dey2CwblnCUPytAAchxeXnCx/JHJlGqS2fohpFRz5xwjRubOUue
eH3RZdak6T7Hk4orbwMwaXRI86kwbnQWdzCiO2LqP+MAaAehvhzLege6fPnsdCVS
KVktS2QJUVLuMT+viWsUQaxGdO6duUIf9kpNqiuIWapvqlJAz5F5hgnjDxdQ5EFG
4qFtnnw3KDwwFR1kA79PuS9m3fGBZ+Sgv67SB+XnCN8fKq5OzO1CoqoEgWtnD0jc
9LIAtjs6vKR9kEJilgQDCo+Y77PL0r6tuFDDEctTORPTFxuqJouqnA0XN7YG7Q3S
x9ueoV7hdifZb5hVxlbxAUdna9B2SgPKRrChbYMAoOAahHqdylZOLcC3NXDqdw5w
Ek+8jzzdHQJJ4k/gwPXB6sJEvxpMXz7LlN259HtUpcH/MqNbuHA8TCpGIAIw2xf7
JW17eg/zg4f/VVzoPLe+3eqVLMElDeySPKDzbXIaagtWkRC4+y/NEoAXiv6GHT0y
I55AssGXD/Wdr4K8F41GEEY8w43a3JUay946CLQVP9QEnwE6AGmdtTkdANmV+3+Z
iWIY1fNlH3FsTPyOg/47DPnLxEt01lKZ3d/ccAI27urt3R2getfYupmxidFVmLYt
Bm3EcWiMDrC7ZwQ1IiryVElSVcl9USXudKgWYQcZ5KOobJaIPTDFBuAZAvvceQ/y
Y1AL19bNbvBq1Op34yOTl0H3koCuRebm1nxR6nvql73NE/0z+n84Uf7jNMojHYNM
ZIUcybyrr7BNEgLyKyh8kX03zD36Gxz6XAjnFKVJ0jhw2V8Nx1KXXWs25Ec/q1fR
lK9UQCowCB/9tnWSQFyHYfyIxA5Uwa/3gt6HawdErOZnstdITcBpJcJnCfOFkGCg
Hn+BRoYqcTbTrbNWu2iX7h8ODc0eV+NsvUSL+NDDM1mvwBj3Uf4ZJ1/JxxUBpjwf
DDXEfwVXz47v/sIc248dvgV26ahwjq2R9evDsY+sZMUg8ympTWF/sd54fI1qgEnn
skjCN6+lRtqu91KrykMlAn0Ms5NzaY702xHYc3CVDO4B0ko+WMEAFLOLg4TYu5nR
8RviwknrKcRVIQBS4FQyxcXGX4LHjr1oxhoVMXlbOq4E+1aJXhLtfVWVEcVPm+9O
kw8d+oBU55asg/C8cSNUu8o97eJjImacZ7bwUEKReGrQ8lx8fXkhHmh5BB4qeTFw
1qz1lE/1tFo6JU+kI6OLV1fLLMPgdFo+c34xBHxDC1xn26BSRqCxIalSS+e4v15Y
TZIDMTaP9CO3W5/ky2gJwm6zZ1r3QyeZ7Mkl9/MSYgWhdq3e1Rh+CdZPOi9D+Rx0
Z73V/xma0j9Oej6wKsmJWhVQFWgwCp0LrN6HKuvsonAEjhHWZjxnvtL3UOmk/m6Q
7YdqE1FOnP99p1RT98BW3gXhPfnhUzxs34u8GuZupTB0XPFgSMwbDLlc1cvL5Eav
6hs5NADWPWARW0IwGVYpxkpl29zhRHmmQlZZNjz0EuE81EmqD2qi1in0wPM6gGbv
QPBVuz0/lnCdxFC5uaQLiKe63SHETekU+0eX8yPyeQUn639jkyUA8oAudcIZZYtC
XBHiGu75A4V+EEIzCw2HEo9F2dNKY8Dz+PbvLSxZO8dt1bxKjzAqOXM9+nI9K/Gf
psHBNnEl+Q/NZ85+W8HaOn5HeQxcBxYYAQxqMwa9EeW3CS99AQ59ZXtUMezku3PM
AnVJyB7Km+DL9P+J8cDMltFvssJG2PncROi66PBR4OEVIfVxc49gSUUaAZ3Daxpi
zP8QQ6Xm59+rDrk06E8a8ETsrxGUa5YrMwY91Wznr54qf+d0feGyVjLKV32Bgb82
xQVX/VZapQ76aes00IfzTfjUyBK/6fNM90DaVN2Uat0qxJnoN6LSzR5/bkaTHMjz
zFJ6gJ5U55U/4adjIbUBDDUriu/QsneO221462ErCZqCZSJVCzwMLjnkfL/HV73a
/tn/2tZ+9U6J8AxiNyaMa8jugnDEEB3AHIHU+Opn4SIXV24KmYkeJ+UeucA8M+eN
MCz7hR2/+jjkHIzFiCRj92K4I/rSYRyYi1OWDuR+EG4S54aqFwdAnO35jMEaSrTd
sndJD1220QljLfdAq4zAGiqbNqjs72G1gR8z07DD42jw0PiaOUFgQkQvTagyw5fU
TSf21Af7RMTOV395t4nVxG9lornndQMP8xvmp5Cbq2HynYw91hkM6QiJPuCVWA0X
C3q8jiXBcEgzycDeqRslQdoqOD8P2Q3i8t2ropFHBJDUmRFozvaxbn4RGhnAjsu8
FH4UacQmjlRAjJuVfg7KYk/AZxNDx5abkEtf6fUF3xuPv1h3RI74CNV7Yrxqq/nc
emC+PRn7d7I5x01e+2KOUkSJ3Fkbz3qGT10kJjmcXTXER/TRG02FsRCD+TBCJfIQ
ExMeS5syie4c7F53exCf2v71ffqyMCoXHTwI8f0XWBI/ZU4FSiJsTpg8tfkLB1gF
2CZ8p9jScFMuDmHI3ZGOOEJAooumhX41jCDNoF7HPN5RXo2imQXQUKEyQMxLaZhP
baHyqerdLBd2W++DFeVliDgLMCaXH33z9T+ZrhoMtISM84rOxiuICzhiKl4J6iw/
d+fto6QjVrbwhmtPdfFeI2pz3tXDgcRbnrK+/Pi/+ZAvrWuMcAfJYqHEMZ2gv2B2
YpZRwgc6tIFqDwRvmrjilEPiSX1hRXUYGe8IWNxsM5xmPd5hi+MNPmMkGunQU4xt
kHBZ6ux8uHp8TqlzGOvndC0XP7Dw6cADZGbz52nFFaEe0vJBkTcUjfZNeUmlWQLF
Tw3M3/JeKzFDwJObUmyJ0pPM4GNdUg6ifMKFlYCCD67XRkqs2wzGqgdaf9MMS6cH
8HXh5gxhyYYPu1UBQXeFrjLFknw+1Akn7fngtFEHnqJq7TErwHLpvH/MNEmYqNDS
t8jX+CMGHhKh9VWDYFIeUlbyx+g1eIbqlKGzngxAIcQKtSyMclDpn8DjYB6nuHAu
NK8mLppJB3QpLiGkmXzQewO451le1Y/z7W1xLrER5Nu88tbK5YlQULqN+sgZNK5/
/O9qYjL+dQVolEoBGd4SwgllmRWp/sU/rKWOYiDz1NWxM3en8JLJ3ttFOEhYMGR+
MqFQT72/SToiyqOigOeZwwDwmwUufk5wQBm6r+9Qz/S6t3wGPMV9t2AOYNzFTXcI
xHeq5qddznavNhtrdg/iUZKr/N3wn3+k1GWW0BDWKbBOacvWJJ14XzqkE16BdpQV
SFML299gboKpD4gZu/O98Eowuhz5AGNnmLUcd0LYUsCuzof6htsvHGH3mKVQg4D2
+YwGjjtWZxAqI8J1jvzBsHLC8brNk+GmKw+vbceFHmAroMVrZjBocpsSZ2XXPwES
oSU2ulJM0xJ4k+67MhY3rTEPseREsH+Fn5QdfH98dCpK74dcI2PsfL1afdpSRrF9
k9Ca32HG3YbRQ1pc1eGav/TR884bMrwWuKv87WPgwwYLoTdaKYKdfA01n6aGRaYy
CwLKrckUCVNkHPTXAAVgP63JC++yz+15ZEpqahvHEAFk126SbnIWXyK3gQd33UkT
nsnore/bWoYsGVn2wHUuGHfI5MTrghoaP1v8ULKA3yYI8Z+oizzoa6MbrwgfnD4S
AsVC9IurgUDkh7KgQdSb8qXNczAYiblEfOux6HInqbdvrMlePfEyVERnYQ0D1OB/
nEM4GH5/03QaO8GxjcNFw9pnS15NQZnNQmaNhOAAqGChnPN5APH7lSZ09A7UdsDM
uQHbnpS2M8Iw8IofYsOHPa5MRYutjfCTiVq2AaXwZ3RMDu38EcCBCvAuGvLdzt8e
rQYKvCvuE5ouiWT+k+216Vc1VGy9Lwcko4HD2Ii8swTd+1Runn9bfxJ4EUsaBen9
qcZWxQCT9TyYlNnrJQ8KuQrp2oSCMUHf/5gNyxvXw7+NZtGXdXfOI+GFVlqP+dry
HicwUdWtJsUAzjHVnFSTYcv678F9hZpfCTc2nhE+j1WQ9Aoe57JR51GmFSN6H34k
8a9dsYkCWo/Y69DSUancRh8+TrInMVmXQrSIT2Qm7LBUqqKbPxLwDtN+lAQIfBpZ
/n/45fr3Au0G8dcKcXUawGswSnWjWV9E1vEPEC9gJ+TLQbzXfe0bTg+iKibSw203
A6fRO5ID5wo18dxhgWq5ji94oY0nJgIIX7XyVaMxBE47avHktxaStXO1NW+G1OGG
OVBz9P6itaS61iFhE2GTbiwxrLHmhFDhSOJ84Gcc1DiRN0GktQzFCiFH4slgyZlE
x+8Fa/c9QaMEL28/bvrR9a8Qu1cCONjr3gpogNhPxGxobB270w68TIXKMwbwSM8o
GnfBz/2iZrKAb7CS6pWI270m+2kwfY+YU8G+kbV5/IQ31T4Rh73NopM8riW0UwjB
2xOCXxuNG+b6fvfq6G/30girIOrlxhA4o6JgWtJtg3QgxYNAVPmNe1toAsHoHGIl
4FXgXfO70Vc+Lgkhh3YZsDsnN/7BCX0Nv8E2mosmOekki/fhgiHLCm0QGEmISX22
9ivVtPZDT90Qqzj0Z27TB2hufaeOdQN2yI84neNnTlT8q2WqerBRhy0LkImg+mXJ
079g6NQQv1IRNTE4ps3nWlVkj22ubOWNVR7IqpCvSuUgH7pBBGkT5h0gmPQrlL1t
qS711BPd5LDRe/Qp0LiK6ymI/IlZmKXQp/zvmHHnLx0pMNcg6MMTRUVDYrZV7WrK
yNgnIYOHJAHTLfptn4v+/YvuCZmz6xRUco8iWJdLyPcF7s9aPvAlcsQewAJoKYsu
d0WPAe51qRcJapJdRUAg/yNsyD3ngVw0SbCuwrnMae/Rg7zjibgIx/8L5xzaEdDJ
XZWODMGYzinTQTMFNUStn6XGBWp9pK5o3VjtZOIzQ1uO4UlXzUtmTVEPFBp2kgxW
YJ6tDI9pvn/ul9ERYIA3+NcyWGk418teI3qAwvH8Le/BZJf1FjbeuiCWSDA0/GGI
WJmMNrLe75A8Ji5Jh0Dlrpuy9oOEH/H//Sf1XYGw0g3+s4Zs4yL8Ec2ezm/js+Xt
ZfTmUiqqJb1YJwuSrakP+nfYi9a1Zi+BXEZYnpTssjkIHJdUe84z3uJJOGFEU5Cj
WZ1Q6+Cuf7D5aH6r5XzOzrVfswFrYnfDiBf+MzwyhHc4KV398kyATVtCOK5kzg2F
rfPZcEZvhce1X7IubJ0fASYw1fIBj0JKKKce7h1ej6pVn+y2maSWW8j+XwhEwk1L
CEDXeeEN/CEs7n5ZRqyq4YmX3liwu9mdGgp140HbQ9PRDLp3+r8ahEUx2ZYsexIS
Y1ACu9+HeYgZg7MjTONwRYXkb1mVmZwUOIUdpRcFJpL3EWEI2mNDjbahORA6WWf2
6tvAaXCsBfboR4PYM1xav4NEHsK+0XSvVj18f265tlcp6g7TtS1ZsV/jblJThUkZ
jvDxIqtdQCzstlqzDZizZS7h2m84zNbaHERbo9r1cWiLyPe0NA7pvPTFiUacT3y1
z/ro7dQJZMRIPhozSM7I8v7ZX7Rykpn8XDvNPaJKAJffe22zl+ZUg1Jrda2URIRV
bJZIP8pRrGVHHlZR9AsFySquFt10SVwHAuLOjmFuC8wmbiZgUlMJDaLoDl0Pox3S
TTe//GjYmdHy0uWOW04oY0+N/0mkLSjEI/Q5dm2BzwA7wxSkjjIVkL2Pw8yKSWtm
i9nzLzmz7u2HqMORZh81e/uS62RouVOVRiU8qRcqvjas2Gix9kxSVTgCmolgyM29
PBHDEZPa82IWPLoOfdNqVSrsT84TbTjygx1oz5ka5EgXkvhuAXlQLQ9K1FcqsYlr
WLEFJIKT51/D+0oNImFtdrZ15AD35kgmkBFSdFiFQhpkV02Yb3yzD0cnZBeY43FY
6tuA1J+Gf14Yn15NMPLMUsALiGldpTTO8D6cmS7FNE6eYCNQsqLiPSJYTXGFH+Fp
ScPK6Ug1pv9WW1W7eiceT6pPAYx3ThsteF5uJs1wuZBZL6vxdyIUVn70C+9bLrvP
PfICfRxA4kO6BDmICzovcoo36bgPR+IBeTOU6BnRwkJ/yaQUaITDJrYc62Jtv3Q4
wfgK9B6Mi7tKBbJ3GL4k0g/DL+jsJnLl1570+Mx867eXA1YP+WXcs8mseZN1r3an
bPVCiTuGtTp8o+/g1AncoQ362uKSdLHc+BxPCEAHrqI7dCbBpePWDoRLQMR/7K9A
zHDAt+DBh5cNgI7HdhZAR8ne9ctnYJLYkXwnfXkSFMhKGJoP8H9m5L3CvUXvx+Q8
iGUsW7GQgryezUwkYRZSe5xM0nKaHwn3/7jzCMApjpDCNC2Ty6cIlEvllpDJ0mW2
tbTfuXD7xCAwWotXjp7ZmRQGGoh7MDOkbG4w/MD+MYElLU5Tx5+0K7dX+HZDx1Ls
OX2k+AfNibrRjiJ+nGJhlzT75ubgkp5TXA7fOUu7137IxrWT4nYHlN+tDamKQPyY
u2+DhUWAmHGJGLCQej8DvDTfXvBzrewEx1H7W9dFDiYuoRa8jFLR1/AJHAbojgox
eI6e5phzjSQr+p6P22qPTYOYae05v0FiPmK9uNraHRwBHVm0UIjkfBqI8oL6uXhF
cRkJkCfToDA2Eig6eI70bbvJvh8NGeSMI3Bzmy3lsZ2d2P5QAY23D8j7m+w8Teot
a6ugwJ70Re8FLaAShBwv3ri0Gg3U4r/gpM6ukfi0/+jnui1LjyMIIRGsvHFWufQd
WfnnPiPDMAumG0n7PqLMCpk7gssKdo3k0nSYsz16PVyf0T6V4k6q/Za4iO6y57pH
2NVFCNazsBQu7XEpVyUVXCOPj/W221TMGTzHTBUmVs/QEwXLCG6e3ZPFu87kmYxM
y8vZkuGR0SpvhHZj/W41kWWrzmuOH3JzkX/XMc00sKZ8qk5i5TrAtaSVQWwx1z2n
YG2ZiYKLw8vi0Gnzq165x5x1qOoFfkMfxGw/A05SzyUNEbTkIB7Hafz3ompFy3Fm
3xs4ff9636BvW/TFqxSkICl7aByoVE35+afIoKsZHUV6+MgAgqzMZt8VpfzMkenz
w3z688Qv0/xBa7N8MmXsP8dQGT2k24t6ysLa0UnnnDlLcnO5bjWf8x0SsElXObVk
R5dtpd2M29PQZhznCI5xLuTYx8udWlLGuDmFpuVsFd8om+m+3pNzqOm7jhN4Hyfv
Sm2Xl3DhdHS1XPEdEEo9Juw9zBs/4VkA3RKggMikjs3yu4gNChQ13WFtcKGFJmCv
Mp2mmE6W2NMZzmVU/USxLAo02msnBeaaSDVAc4xKuF0Z8k3Ph+BC/whf2qHxl5RK
o6/xYm3UcfbEDvZxmVQwHTtESaFznaPJ77wP19o9ByE9CGJ/lIH8lcM1J7iJ2e1b
C/cPW7GNqBQDQht3usNPaBf7b6AQSMe6vqlYbv4+1MEeXYaQCJBM5pMFFaeQAAm6
19OTQU29mj8dmWtjsWuxK3aF6hQZ28J1507BoC/vsblY6mbv0F9LDXIv58m7+aam
gefsOVs6fzSGrAyiA+NP97wyasS8kec7RBuH4/0lbb4/CFETkD2lQNDB9fmsDJUO
4H9nRj+taTFHpqlQz7x+HPFLkFstfnOfOy9lvXabb10WMe9i5fMRRMNtI9HM2Iqd
ynMF9l7lxTmM/aObzEA+y2wRQ8Hs58EovZZKGweN6alkw50I8WPBZlBZxSWZNqyO
GELczPM6vx1TzhIUEkJ6jldK8cO4hJ10MVEr6R2IQZdHKPU2F3/yGjj3sKUQzVr4
prPhNO8CRvotk5JUVAAnrfolElofTskuHy3hnaOFv4qm17z6eyMR9KgcRWDzmhvW
lqOuisxrRc1Acyqcd1o+eZOs6AEyZIIzlWKVVhvVjtGQ3hnQOE07lhcsg0Qu8Q9k
s7Zbw4I4gXhYI+N9gOrIXKzitWw0rtSwnxqoYghKAIg4NkNfVw1k3V3G2VjEj5up
fpT0cZpp7ybku5xSOPcWP9dO7AUqNOWZzYUlR+N8xYVxeCUr9uaz7dCZlmTbbFfR
JJSu+G8+WSmcUMs3PT7vR46zeWMMXTeejCMvOi6TKHPmuQ9ac2+KLLwyg88AEx1N
5XywQTQEoK2wTOPY/zQBTo+LiniQeWBjlQc1zX/E6nCwC1yplD1mLhNWrBjHGvGN
Tn7PlshosKAhR5i5tjFYbM84zdIhwZUM4DEWY9PgXHtFSDv1mr3IqACTVE26Szdd
6KwNXU0VM/vhTRzFD3lRKQS2ZlO5o2zim3K4O+lm6+Zfn933mZ0MAZrQr+Ch2PMt
82Zztnrro1g6iaRPwrnTKSPT/nOUcoSq4PGbHvngu1nG8FRGrJD2NJoHIayiaxvy
M61rvThPCZEZJxLzYixqcT77OqpnsoHO62+yabGWNfgXT1qpqNbIXdGJItq5ROaZ
+Yltdmq0zHaC0dhWLKbVorUgx3eVgSbuUZyFL9gLCCuGx/HwEIiF7QQrzSJYN/kX
QsF352WQNFr0HIrOpPPNW+ovZDJRjWgTPCLk9Jct7gppl/3xIPEXA14+CEtTfj69
X2id5m2Fqq2UxjNuqssLeTVEBHTrEo8o7kwxILcyNYlpKJu4Dda7wx3iBMjcscgf
6BpBeh8cUC6VAiztkcm1d1e4HYfw4U58ZZJvkFBewaxBPQvf+FmXW4MhYW4AIGud
/+RbaNThN4mMn5yD62oGDHfCq8YfpvBPpqZrPV7ErajIT/P3/DehJOKlpi2P+Gaf
1YVLnKtkz9EceSpPq37lXNe8jJ4khvrg8TZKTuAxtEUDjHvw983cuDGj4bswYFYj
1IM3jp9/4LYUFKALNkm0S5anlHfcKR5YIfbKKy7gXcxqwut3pqvm8l0K31wiQom6
qWYkdJFmPevF/4ZeLBhh02XE3CYV2rT9cngWSklMbIa0T1quLm1GBLC/FHFW3OIl
ng33crw43wCcNqgAXcImvOHXEPZxwk0W9x0yQZD9BV7Z4apoHw4Zp60VFrgJ6N0P
RV2NYv8c/K/7UnxNGZ1ApR0Lckmgl5UT1mDXT5qRlQN1R6zfxSGB2cD2iCrd+Fbp
chcjYIi7LfjHysYvPtv4bsvLSgFOJQRZ47peKmr08IerL2wITo+qtJU7iEegsc3Y
cwqG/9Y/0BXuyPb1v3WqGezas+NFX1hLkBLzD0JZ/+5Wh/yk9cJHbzP5dsANrYWJ
pr0r2v4TqpVi/6t/yhwO4jMZ0pAzP9bGczuPrvCgs41c+/wIEUADniwT57KcilcE
iOzEaeWSQo24CyDvQF7fIYlykh5LAnXLbcUqC51+VmwmRCpQ/EY6XL2PLnz7qZxk
aD8gCqOC4qHo742C5vqFO/O1ByTeyxrGnbf5B+IVjMzitgyGZeZY3fEQY2G/Ry0h
IP4ZFtqM5DReoVviiAu0rNu7R/IIqM7hwZMC7yh5Ycxb8R8E7ITL9KBjJkurbW5f
z7PBBu3mjz8f1a102rN3Dys8QcOfNWleJj9s/piPPTBXg2i5ZfxOplUKk8Q2HsUQ
X0W6mikQCBveZPcPsFGiSDlbUKGU/BKIVH0rqGHym3xnsH1cZ8oeY5j2NvG62+My
bDf28fFQwExNS2X3iBp0ogksiWMyIfj6eGJiM4stP01orsh+Z5ZSQn/YOzkq0mxj
qyl8tFiLMUGvlZpjbHOyfUmEwm8+fW4U29KOF/CWbWRrMU1j6DGsAxdWKpQbXq76
e7U8r6hxej7jDqI1u6YIVOQi6cPQQH2rj7k2tYtnAeKro/vLb2pDak606LeS2tUO
2xHHhsiuG36Yduqk1nvqq9Qxjm/n1SLf7d3s38xGJY9KNNcm1wPj5wEKXMn4VfJC
dn74wYj/xEcit1TxyXDRGjGSsac0n9dxISmSruzJBluBMhWsScrW54t/i82x8Op3
EEQPh8UPIFU6o6/iUaYcywY4W/NkfjcqiHmdksv9iNtQZp26oublO0LuIdDI5MPF
idnsGyZFvyHQzNvnzVCC7S0CBHhgDh9W5LHYaIB2i8FDLTPtT+oFMzj+WO6d32Rx
RCU2R3UQrgq+vBZ1GUW5CnBAXL3B8yd+/p4C0U9Pqdmhf32HKw9nAPkEN/2sUGXL
aX3zCa+CZrUIKRvvxE7hCed/TVGAonaHEawPTQ/94neoyAKfa3Y9Hf/R8xJ7Awd2
WPYqPmDzVMTE12w5lNRBm4u8RcfX/RRV6UfPWh65QlkURYwWpZXZ7I9rgoR+IXtp
IgWuW4bl20PO2FxR0reWVKAaJ+uITNAgg2/4BFa4TggP1PvwfffKC9ID4gVgpgQu
v4eeb15ZiFRWBuUTEfMB6yRmx7tqVTBt3yvlmAO0q76BVv4/h8dtU5b4X6GF1VTG
TEIUgnNl54L6oSHMyyyIMb5SwpB/lqxeKF8O6g5DFlVjKHes5rKIDUQCuvqora6l
pTeEX1ts+fWArHrGovPn6ZT4VgZtSZJn0ufH2Zd3WplSR4eu2cIOwr3xeRuyoB/x
/4r7DKttPdFkVYjyjLByMeqZuKAi9jf0C4pQug7lT015twj49dxZ1AjAZv6i2Me/
78kwXSYamGY9iFZKTiRvDO3UaVr+pKwEx9avZz7P30lKfx3dvp4ETj6k0HeEWmgq
n5SRSA2CevWjUh/fuoZ5O2sOzyc4ngvXFaS0XjCsT6JQ1w+muH81RaVDNXwqL9u7
nLfci3m/W9/s4m4AuQcplQTjklam+6by+d+vYnu07Q0sI9p06Q6A8xURlm7c1ryy
Z8/EPtjJhkSqvTpyOg2uTI3GwsX1EJEpTwQgFoM6aqmyR6cTKqZ9vc7WCaqX7JSc
r97VlMZK4GrT0aT9QhhIxP+EYnjGhMOf/R+pSFVjpzr00Rmqc/6rJoOUp6RAcDul
HL5Hqya5enjYSoWURXFImMeNWwZ+9yUztiouA0C+r9jsAiLFJeY1zD2rxTi8UBVE
kIXQ3fXAYu8KUBzrrSQNVJVNosIxg8edjAArE1DEINt1JODLvvTXfpKAEJRgsW6i
dgBvOEQ798dgS1p1K5qaCjgjKCpxEtTWU6U+v5C75XcUd2v2b4shMkBnK9nUDZ6R
80LaG1pWJ6NrhNpsCCv+ZlOmg4/0HLNnQJeWU5Ag8vXx5D+AmrgQff8d5YmnfFwX
sIhAi3by0+N9YNjnKOTbYk1s76OhSdpVsaj4HcSUCrQGROtqt09Njjy83HO9faVg
N/g9U1iiNMkjt2umPAAuCzY0htvQIpnX/D1XCCttgj1rOnHIcxcayBkQsa5uC1w/
XWrLnXjwRiIGzDcMyAiXwkPa0ddTstfUYfgLTMgeTADczyBAEQOmJXq3Alap24Ax
PhjeXXrxi8igM2j7KLrUvmMC7RVB31H5MJlbDlRqevybJFva09idqUs3jvECk4Li
cZxyQTjd5DU5VlZ96LLbNe0ac0abGKJXyszWfGWQoPKAiccduZp428EwL6v2vZ22
bnDqcYlgVCFDyYtRTrib46EE38/se05FmpMbi1K+rgrupsGZZZRs+ecemfcJbLpZ
XanT3mwIOiYR173RBSNHTAzGal4xWWc1ZK5CGhSVxVHPy1ADBNr9zaiaOwf1A5q7
Yx9qyzrfeLv9tsY5uSypM4LEipdKXix9V8SjY6QbCJmeAemHnZn35gNpmFbZwQaP
4N0rYoFwelqwOV+jlM6W/Cjc2FoS2zN9f6CwOKgCh5liy/XO7qyhF/vRerpeA0qr
W/BTmNja3xkadp37yxSSYjpV3gOTJOY7vv34yvRE32bhAs3oSASBnRBdl6FqGQLo
F6RktphJf6OkAAfWiTvB1+DJImQLPyb7QTb8FUiFLPtjXOSD1hRloNGEkcThinHL
ERRtNvpp6bMMnlltcokvcedvqis9hvmr+XPP8Dh9WfwiCk4nAOOcev5WLX7FkSwR
msJBG10E+UTWUPdII8MWgCWc3vHgS8XpgCqT4bVsEGci/VD1y8U9KHgktH4uj41V
qorLRUq+g5DiUBTvPBZEmVypTjtItTvRmMZWRBTc13oHlE7Q5/JzRZaU6YMnNHUl
Ix/KvGEzLmTW1NHtepACZi5HKB7hO3JlfmoqfGhPfiaqL/CDZsfOSC9uji8Ebob9
LMRnu4Fdum6y8NGSgpYnwSKOZ+MB9M1Yu0z8uGPbb6DxJgFM44Pfw0U2U6p8MJS2
NS0xH51vImFl9m5eMoR6pix9vQD7lksOAsAQHUTAV9kb7csFw1fyazKhhHoZ+ZeG
7jf0rUpIS1ohsH65PgkEU/7E7vhru3v4KFCJhbIrIPdTYrn5WMXnAhRIQc/5rLDz
GQPyDxCjfaFZ60+y8+0uyyUnFVQ2CMd9GvJHuEmCXCyjXqietw/rvuGcQ58NUfUu
2ot9wiweKJfL1ikspz8Fu/6VAynw65WUzXQC9FURBqQCMArwAn8bLQgm10Qz7Bu9
LJPn1/1iE0bEJrhjjOIeTAqiijF6PmkOYwFJIek+3+cg3yyDGHoDhD/WICKUtz3v
5V+c/PuNBJHZshU6aDienlCBlq3KETlGJ4XTTkXwC3JmtbD0PFmbv8tTczpIIyp2
y/ra36WHQfssyCiHegrvkRvJhkpqGHd+bzNme3tVZej6bl2Z5QdDKU8I2KrEpE7F
v2t1EzVWyTw4UN+w2vnmz1fPGIwtQqnsrhargMhbtRIGIvSGbS1uLaD6F3QzU6N1
9WJs3CJeizXODtzf72IbK87e9Nx/uf77c5E1nqgj3WsT2fbeJHY7swdCwSu12750
JQ4AjC89ILLMnl0h8CDBlLqVKbSOvmoFjtY/S53jdoqK/yXol7pGs4dukEwcILPv
kiWG2I9Y/4WVYYrint+fl6V5Uh8Ga6N3vhm3qk8FNVdtvxwWmd0iIXspR98fMqkn
nsMTA0zXMF/DofaNn+hxQYXIv0E3i/6YXGkr/0WfZYDjdN6Jo2DVvfTTQGySsEoI
FkRh3kyF9r/MtGse7wLUirPRrlN6mRxfr7P4INsN10kr1zdvUCDEYnfIhiVEgrKn
jcl3L4P5qpzrKPRvyXD7D76YTehdmYBUIxz0ok9VJZ7n2rhlc0afvTMuj8kEkYYR
zBbbLNPVGuaqpEnyYDxtBWIUt3Lia3qVVf2ca9aTlOO38zMa9RnOax2eNX6P8jK4
vsFq9gHbx8bO5QAoj74kBe1j/mWNcxPmTx+33hUSlY7ADA77b90TLXIS+3HJXUNg
zBFeeZOij5Nnhw1NEIRUjvnUWuTWvfKUs2EQy8Q3iS/rEdrykVWQ3CFZRMB/k2qW
eAoFwnzriKjpwDCVX/ajfhehisnkBmshB3z2+dMMnD1fgBycCgCvQOkkSim9/cgI
GNWz8CQnT52yhsNDnAj0qn2mKBsFhZT0DsyFR5qJZChgSNyOCFC7dWsT/wOqgXyE
koPae9nK0Gp6q5o2ij1bsUsgiJezzOoOtkTpzcEIyIqKcuOf5EruMueIlMkYWjzh
UUwqhUXTD7VTbV1rOaH/9B1uB801r53tqTCHk/9hcrucYASYjYsNuXWaVywHIqKU
hoZQXqNd5IooVwOLGTvJxBB1fr440PNQxQdXRXr/0LCQkPNPISSHoyQdzuSu0vJd
hjYBKKfUoTCdyjc2kFIAdb6PMrEU57kYf21IRzP3S+fhloVB9hisvJEc2nXb/SGZ
Visl47/qiPZNzXFlGl/SvqcS2+qZH7pKBf8EU7kX7n+IlSZWibWelH0E5CbopGMu
vGY4bc78gkwRX75HEDB4Bu2kmecoTy6b/UipdiF1HBPELvjtjtLkigmlUj+Y4LlT
F3M4BsXuNnsWmtEojbKGTl5thbxkUNLc2xG6j0ssDsbO8ZDhf3px33UuRm6j+eVD
kroTBBy7UeFkst9bWDeLY/CZsITYY2MVRQv2zLcuUhnkxV3E2fBGvWo6LFt02Utc
XUX8JgxKhmRTdxu4nnSRSIZegDYTHRfFS4B8QHSYmTHOb0VWYtpAR5wXZuDyiBiU
qB7DRzdI6ThCrO4hU4nIpdGcSCHfvCYcNup5PyfpnNgixYh5d4WXIo24gVRo3zVl
//f6NfkSPsYEDqwDN6vLw1Zal5OI4lNVGMCKBlfMMCEgdBt+osRSUOdGt4hYKFkL
XHpVeN8ACnVLeXuoc+PPsv8GzNrUnc3YoOG4XYAAq1bo9G5YTDcX/gTFeW1g08ZC
4fXrONfne1IidQuaGcHm8OXqtyOkYmyh31bhaofhA0UgiRyrVOJA9k6XKRHrfQue
RDQZEXe+5z4lsSN8mfoT7Jld/gC4IZhuDCgFHPGy/FCkOL+PnQ9Jk2V6cdMkxbG9
mWMY3VHf5M2hTEgAbh1ayuOQ3kAZsMeqQjUHm/JjjuWF4keP0rLJ2Wcg9S8YKQ9P
q52aurXhRZqrR0KTiWT4+GLirRiJdZ3D0/kkwofeK/H1EdSD45PEvLubNBWI7Jmz
DLj/mIo/Q84M8UfZXt32+PEwknJgwCVE+j3y8F1QBygEiLfDzhfx3Dd6l4xWEcWN
rCQ7GHkvs402aGFKBcRJej/Qtie16bK0krcwBtzUAHyP8HGlg6Lv8ErPUt0iV/6R
z8qm13m/0nzhh/iVawZ3tYTW/XO9laiSJldjUVv4wEwS1YDiGZftvbvGG4xf+OxH
HzRw6rTUlkwL3iyJjH1svEpUBEYgkxGRn/3BtTO10EEsXMn8db6rVT2ZUvkRP6Wc
VNthts/56ZQi4AxPScsXanA5UEONdlX1CyeTyJfMbf2mnVd6zZyhOZqFHBSp33Fp
R48H8SGa2SyCw0TOrLZzGfoBFYEBapahPb74anPuUKHp90wdFmq9fJGGVQPsAF7n
5MVfGcnaqK7zPEgfXc2X5MsdDS1wGVY/nH6xyc553Hy4GEDzQK29MpF6QF+qg0Mg
XgCCEOfYtE75d2NWOJ8xYIisXY0TNZIUiIxUmL75OUQWnMBWghO80prlM+k4hRPp
EOzta9lF8rl+c+zJ4827VfB4KpVz4/NfhqIV2LMAuVI6ZkSzprIZOCmszseUDaHY
qzqfUIhjUJ6WGxzVAE6YsG7513AWAr6TEeq5Q4Rq3oWKK0SXvgo/AGt5bRBvFEJs
oc0X3b/4PPZ6tSA0GituRp8OP62lP9O3p2vKNfI7Y4Hg4V5jD4Jp78ELBZbHHSNv
6Uzmwt+VSptQv057tm5m9+93oV8qZ/HaKwRsdM3Ocjh48AtKMWR5LmaXrxthDASO
4VHCQy8Ss5k+d13lVo0RLf2S50V0AOOOLj7Q5/aao+39WhcBzGqYc6Wr4CTNt3F/
nPCcB0D8OlMtbqctJgDnlSzKOP0BNVcJ3IKDpamZ8bLZY4eQ9X3bVVyybwNKNbIT
WGcmQvy8a1YrU824omu+sVgVd+VScg3GRQVDTTMfIerowwcKddTJuQiWZEFi3bqM
yuDTxVeqD0XyP2c3bX9uJPFc6Wq06dMGefkdd4083HQwwqBczOQQLFmoDJl1Fpep
YUfbN+ISDYfzrHE7+jyEd/aWAL/6FdjSDcqlgp8glrpa13DSYROfUNpJUUT/suSh
TbpBJv3b88dVoqywxCfQksa1LrLjJGXnJooTqCJfuCLEZsKjru1yAXrMtsyYKy1t
cBURQPfg+unE6pMsyXJKYjIk39K0Q3fLKLkRkoyqjVYLGzB7GH1WvoaphAN1gJVf
QW8kjH3VxBW/5vbnyYaweJnafOVOK/V+YxPv2LmmGd2iIo+qyu1SSXxLaRjZHzlH
KOMdgM5HjyKXCF7b/OhsBOQrG4HVHVTow03KNDGdhEbJ3NWW7oEYv0OV0uJHTIUr
yBBo7SmhTu4v8pTbW+40rJsyC3SvfsMPFIuO13TJwF8q+NPYR1cbpn8gA7DV7alB
If2i5MoEuYr7Cm9+RHDpYKo0yxghxqMe7MNUld6h4xNr6kwINxHY+iO33/ImbKqE
TOopCGfTY1IflPWREX33pxwBo49oVz2tLZG3k05cnsG/RavXFoKotUBw2R8bsOmV
LxmGALuNfUH+r/lnOLeg7AwzVyOuHtOczk1Nyywa3ozmE3wlXmA8MAJdK3BbQozT
pyOdG8VlhHVRjt+y1gPQEZvJglJwlM7G5Doindr0NT6P3+QVIdHIdHXEA5Rkpva0
zc92DmQ7Vn+EWaab2CGR/ezqCXGDZDmYw99Tj+dCmL8A+dnKj9CGT9UVurclOkgS
YhgpDKQXQcyTITBqgj+FCTHw/Fvw/KMnGxng1Kun1/NxHmtSV9CwScSl6vskLEKV
91tKNZ7RogG+C7WLjZgqeFECM39wnszJqQTHhK3Ppq/sk45AgAsqqhIYmdhNisej
dHvAJ2yrdzosWjfYbg7asXfnSpnchRrBjaM4ruokqxT4Yks8XhWL7Y70l9Ic+GdN
+IKiK+am/SUdKSL1creOHiZE7xblodYS1XwyHZxfqitgCdoTua9DBSLLQrZAVDOg
QkAz0FTnQnv18Uto42GDDO5WnJ4B1G7cDS5ztSMcjmtz0Mv4cYQUidsQK6oqVp6s
yqGWHNZzG3AtZUoFoYSl89bZgdWPTQdhpbX24OzZTXEthh9pO+Dba4zBmiote2ot
Rn7WLSiLPwYKvki2ZZAgV+XwfdUb0t2EY4bGguJi4IraQahi9z9tQu20qhATfmSF
kvRPcDY4cGj/R9LgglNzQOuIWf6f9zMI0NA8aNmya9ZqmCaopSPg47FJ8mfBWfqX
zdd6y4ppp3qso2KR1gftPR3F+c6AqTomSR4tfD5vvS30qA1ORp1Fhr6S1bXsM91w
MB24zXlh+Gu4tQoLdw7gds8jo1pljvB7hflUeR/GqYPYcTLqrC7RIW8YErX8kmVU
ZQs1+P3/lKuxvUynLkmHn9YwHpYK+kBBac73seSNzriixXsDxuLyXPdEvmdUhVuO
tARZYNHA4yBDEZ82zZSBrsFWBu4wz+VWoM7qoMPcI2mE4A93ZJ4FjTrH+oIRUVqN
QPy9VBU7C2npsO9j2NZEz6Pq8cIyEdKwGBSVcTMC9PKoG8g2ClTWQ0MTlXyIpcDx
x2mtf/d/URKXUm1UQ0DSLyIxHWIk/1ZKxCMrYLv3E1+wxpeVy1CFWoNsJDJ4IeDc
F7j1Y36Lv6cqMaPIj5IhIYwbNXW42ZhaJSqNgSd2dnYFOvAIBU5AtgzNHtcuqyUg
N8LNPoxwkhm+B9E2FEo0Eq+6EkN+QORUsZPnqoeU6Pnu4coYmary/3jmALOzmi1S
X3+nTbZwOn6diOLFcKzSZbAyB46YXpip1rMCcXzZ6DInnNTGsYR58Hz0Syyhurcq
6yfsK/PXP8aRbMIIfvbftlFlIgclxGpc33g+ROxQiwghcXePBEW1VNUeYg6uarkr
V/3QFJhjv+GGlTw0kIexURbI1VnIo1/tmwyJRON6+hnXfy3PqV+slffA7Dlf6jl2
vjG87Nvf+lmeMOYsi1vPUh2ptUD1OrHIoW/TX1n5LrvKm+HyeOXTjfQPpCcvooBL
BfaMkKHGyB8+vq/NtXHiqQ8xd251F7Ymc8OfZ+WGb5zuD+Anv8tibWE8KUuQLWj6
aRLzqpfBeo53MI6pZeelsTSr0TEnoxDoGxZRnXVcJw8UVROYXjUvodRsVzJ/v/YA
geY3JkihJ+abSNxsXzMF04Fm5jE1N1kXf4nSc42uEkiFcVekiskEqxs485XUXWjt
JarRzJ/VvUj3tea6kax9OrzsuLqwgxIAWcQIC66XXrrPQ4QSWUKgFofxeKW112It
wVnrsTY02FUqD/tzclXTButbSUWbldB/KXn/BlD2kvCNQYUw1jXuQ9hTl2mkk7iM
T4yRtgdMqE/+1yDyBmMHSMG58GrbTVisP4kM71u2ALGAzjFY80C6X1Q6jY7s1hbj
q8nxykKIE2BKY8rMvka9w/T1vFytArqMvkwIaeRUYyTcvcI7Hj7p20zIZLyBOkH4
gNq3M3vJ7KGAnCIlsN7nf0A/5f+e5Q8Bd+XbKeuMmntmet9kOkXqN2435JLkLM5t
u7hNyuXN+MYy8trHUE7y/Co2qhqq5qd9FahEiDfeEs+VD5memWjBVg7liOxdFHWH
CqI07R20At1hy64kHCT53XXRWzG2oNiNiKVQrFw1X5a/wrw6gGlwPYlAcMqeibJW
OEza50l4D0Xve9aYuolZIrHWFkATvZiOEEPLVvu1KLW5b9S+uPh6CwVWdZZ5shjf
Odw8e8on73jNgbnDFUPeuVydROtf272VXN0fLs3B0cgUKEtSpv9CWJmvTNGWWLQm
pbZkKIdADIoJKKvq+/rw1E0rjm4jC+8payfCvgr8nh/gZtQOhgNrY+qKXAC6FdeS
AbTqGS966d2+SMAqdAey1LsP1WyrM0gGZgQixtml88ld2iXm8ZNiASflqSVTNMp7
+yL6hhNYfgbyQcY+OcLR+0skAbjULnikBEVYvpkxW5vrYs6z1PMH0LKSBpQWgCt5
5e3G/rw+0aR76W0gVTGmaCC1k25iXgKGdGkhPf/qVdY7+dNhDa1YlZ2bcYaOQYhm
QVQUryE7//Ja4hxFRg8cZMmSvTB8Xq7ZUaf/h2yNHau5oRvTrUccGoM9r96rSzns
0wBkChMDfWKDL+337e+98wO0AuzQE3JTYT7xuCLUKhCp7Sx5feC9PyLimLudFmsz
6x2XhQ7doHqskr1Wh0U8hPd1EKxns/EeSbFbOPlZD6a5NuHt5OEqDT+HLDvA/y+d
xfd153A3sRtlv6/+VHqxdZThWI0dZ8Zcr9cefx7VoY7hMwnhh/gEUmRV9rm8mVlq
TF3UQ3C44knENqiuTKcEOM+EAZpQxuI+AHZijfc3CqF8dQss5RbyzHdZWz+Sj6tK
hxHlx2omajdIG+M3H6z5W5m4SoriiFWa/akxwyrL10XVfPPOgXuOeij9eE3W+xuZ
uvCZZOyW8JZPyUJk08xdPvpuT1HXopq/edECiywKFlvZ7banEUqcYvH7qUQM/NpG
SOchdRcDqfILq3pC2sWqe82/YcHMAlQncvs6TcsY/3V1IQ4waMZwmhe1XIQJMtae
003Pv2+rJu9VVzO7EZys3P36CXJagGqAxNjbUy8iXATc9el9ppwJmhgdBc2bqLgN
zyw4mWpzKMAP0RSWBcfTHhVg28hMo3QF5pDHt0JJnM0Qrz8oK2y9xhNky9LX0F3D
+dmfbjMeAUgQiRGi18EThHTJpjyAU/fp4LiNJSX+UIO1eHcQv1u6ibvBn5xbD1Ob
cwXYBoigzVpSWyQ+GXAslhbxbYurEGpu8EZkWOF1ETgkhnNlTox3awmwFiXksOQp
mCUoMj2cn4kciCjnz1MUSEOjej5PZ/vPmYh0CJ5AA0xuOeQ8+uFiV1UoeEPWf3qB
r+fPowmYijoA0ZTFp+4XofSfLL6TRbk/bZNoD3L2j1FEZyRJiIFhX4NZUZpAhFVG
Ea+cOAv5s7fzFnFge371TodytKvzWKkRePb2+pjSRpL7gsoL2xe14j+hFoy0D6Lg
fRSHvmaiuF9HShwjBdhu4BPvLREUvt1RW+5bE//bJpxcWPeUMyiFRd3EKi8+Pzo/
Q4A87Dria9kTI/KyY4IYYhkMnhVBt+KzcjR/yWEMXOUDRkNoZLYuQj2rpcQqEdTn
FKd3RghjOe0kjzTOEtpjgEoTDX/uMuSlGi3SmbktvgdcznOU8oAVkqn5fI94yTh/
t7KMXR+2vJbineFwLTfrWBkZIe5Bczr2Md8F9qs5aoWwUD6o5WeLDC/DArh4OA9z
GoZAyCW1oeUt6Ket77hUSstSKtUhQLG/LdEfkZXL28BjhXpnqGtBfRPJ7HhHO7Zq
TS0I2phT02TL5kUp4b+mlfoYDU1XIabbFJYvhbUQZX647Wx4sKxIwbq0d3DYkAX3
Sgiq5Ypvkc2zYK/wKyulRblvISXvIzYFiSH/PR8fXtojGjBGJkwPM0u54vWc2FK8
t7SfexPaFxLv2d2W2wJQhrrgDRC6hP5ZbAd0f/5P6nmtmrx4Rau3TWx934/ETuHX
rXVPb9OI4cz8x3tZ+fq5oMYfPkggzHSmd949DwMPtQIrFPRFcOEaJkVxdyg6VKZE
Bc2PDBAGJNlBIHs6h/LUt82WeTuFO/idwaPb7CPFVt4FexAWldcyuO8wJwptcqK+
gS+4+eTmxb7szx8HZdApuL8I+nDnesDccfUDB8wLNcBPtIktQG2XsjoLD8zL7iOM
NRrozxIKTmKUYMWwo9GpZ3xlNxQdogy+r0XyOMLuuPWTaXoKrrwLVnEdm57iyuhm
9/TExuWYISLzJ9h1h5R7stO05uwB3SQJca5IHyT6OfuTVujxwSm4LELgNHr1DGr1
1ljZ4W/agfv9nzDUOZV4Gy1WxWkoKmpMvw5NBlQGvizfbOqMPVS6OTmepJdrrGIF
lRFB/NAQ60Xss5XekrYG/xz0odTrR+/0/6LfAPbiWJ9BtGwDr/e26fjZN4l6vife
bhpZf0gi9ztPeNpUNQs7OSevQCfiPiB8iTg6z0eJNM3yudiaKvEct0eXkPHi6OdW
Kty3qIAu138ViYSyjQ2CODEhmSmVU1JtGkSeMKqfD1meTfX63Gad0rCeynsMbIUb
B2af5e1jd9RfMf3dJh0HzbVD8Hzbnr6CkeVXFHIH1FYz6rVCYU2qoqnB4xWWELfv
JQuWIVU1EBUv+dQJxe+u0imeI5ovEb5vE1YvD6QGjRF//QNRMnRgOWWHeL9bYYBj
xee1FFR2twWmDz6Nrv8ULdM+DW6kILcm3G1WRDyrECl9ykmmEkRj1E7VUEGcyYzf
q4zWcO3Hkca/0/gWlNlzwMfDFp6Dq+S34wQl/GbqllkLhhCINhMfZzYzdrkzi6Xc
IwFpgbWcx8xPiISR4oadXCke1tNmNMl+5jDYd5ytlTGpOGgS/l1uadRTMY0mBAFS
VpUs02Ur+N3IrXHZOQsissk6skBt9Z7OSXdy1UZgDO3WXj4fwqLV2d29TcLxeulF
ILwnY2eZgeIMS7OziGobGrOXWKqEz60LKQr1lTb/ZWYmaqTnKum37jycNImkTuSE
onioPYn3syWGSBCTtOoZgR0oDOUlm6P3fsNZMHG/M9c3U3jg/TjYlVVMqbpO/eW+
64/ZuCg1x9BlIPfL5pU+/btT9ruDsm1Lw9N0L1Jr2MEkmqb84WsZyxOyu32dLzjX
p/S00dlwupuIG7myX4fkLISvAEo5kgwAgk4Du0M81wM0DdFnW6zVZNyF1aRwz3Ro
h76ceEkFHLgthmnn0DKDPV28cTAlFunNG7EkSSnzzM1CUrxLx1cXH+09bVQTcv+v
BfX4mFG8M5thMT/bPUXgzBADF/SNwXDcpwhLbs5rmkwuviGkxGIFdapNEVL6aZtw
nXTLISw0Zmnu/U8RhR9nLBUhfUvE74QYZMgrDFoGGdPMlYpBFHPB9IPs+jWBBb5o
zErpNAr5uKd7wIEXiaeluZI2J3IYXwXFNysPpzucQUo5lZtEycLSt1RrD//kjzY9
Vw3K4b0807jp9mnHhXezqlNxHH9TqaBMFfI2vLdgLoj5BlQjE2Ky8Dzzj3GCdrb1
aeheYuQUBhvZRYCgXwj+3StkvJT7HJr7W4JvEGA+hy15kcoMTDH3uN4MKJdeUR7F
4GE6Hh3ppLJkbcrWD9NsZsulKLtENXhecjvwg+GL4ZMU5QD1ZRjv8ftps4Ta8CsM
iCBmxG4DgCilZtIVGc07lC8Qf4PJTQXjJ16+FmJIBaIX/LXsfNtvE5JlH8r0GEW1
lbfd3Gcaw75JiRxSUOX/vmhg3dmjcSeeuyg5eyoqDcTAQmUnmj5z5PH2DWMUBtiq
r4os2GaLnFcUvTteZGVn0pHR+Dane1u/SdAw/qCeXrlt4fva7L2z7mhlS/JUfuoY
EOksHA/3M2jEk9sob+/gqtTliPiE8HSQI5KOK3b8pMmRtLAGAfBM4SHuBOBQlJAk
C2BXHpxnZKudm3z7XeRsaFZaQ1dtHuLVxRgmU8OSAIjkebuDb0Ek+dr/X8cjT10Z
iZ7O2i7XKEDwSav3fbmHWgYzugbEvl4dom4M0APp71oIpgsjGj9RkgkGRrw8wJNx
EQYnhjh8njD5mIU1Mry0oi5+EmTRYkb22miUFPAbx/YyLgcrqaE8kY1J+w8NSzzV
kvPQw/4OJDwsNBvKcBKPtFRL1QO05/jRfYcDHr52i/Uk14fXKdDLjg9YwaOgWaNT
xmhICdYSx7mdUjHdwMlFkMGLGqOzTrypjori+CUz/Trsw7cEZ8ooL/JYKqsAtER2
D8xwUJp0XonjjDCpEblLKXcmDV0zRwrOBUHkopWZgPhGfwJts2qgnfNGUkfofYXD
pMZ0ySUTFyT9OGb/w9nPGmA6l3hrKw2C+XsZF3JFvgCuRLaOV3K+Ydm4JI2SDDRV
lUVQE2gSN/o/QfAbHo18ysLy75S+eDVB2btU0dqxuQaKJ2LQ6kdmoRbeU6MlQc4y
2FZUUogWDHHJiVYeLYQrnIijlR3KGdWIjfiH4KuPQjU6YFdhfbLWE2+WUhU7JQ5I
SM44tu7Q8zBMG6CS6Umt2+yPUgkD5y9AEuqfMV00bWPI7Nl9PxL5PZF374BTGT2T
l4FLIVaLpHg3W6DtB/1w7eIR1JZ1WEBCzmdLYYJqs85+e2uaEsAWlPhpfvUXJPsf
dMJkNPA81G1MHrCoXdE90Th5glorfT2rarOJAnhQDaFHnV0NbUNpEecsQLpxYHmm
GP1yCzj0nSFcNgViF+h5QsfnJJBY2yS1EPnQI1gI8HGmIeBJHlMp/ewigYXWvJXb
XILg+f32A032LZVuY+L8MXM0MWp/mnSTLX0fVvHeUPvYtNmFMIQXpLj1ZEOX95vn
nCoWKEKwwBky76Flbm1HLMKI7Hp294/tNlo6Z6IGNvWWY9DMBa7LTWWhJvWh37KI
F1l1YcDaOHcvEOKGiNqN08S7vsDoWWgjAXRw8P8WE3r+7J/kixby4WPexevYNyll
LdkrS4MHCHedvOe6UrgydxAqWBaPZffPrAsRAOb2v/NIk5PLXp7OnBRcJ/q8J8MP
ARP9jGFYkDrUVuY/ylm+VirPkB0wNpe9WjYrMV/gw/UVxzEkENGTuASFkfOJ23Xc
5z7Qjuu/jg1q5qx8P/uIfXuAqWdLgSnOCFZ7Ee396rgnNub8Cea9xGBtUzj/aEO0
kGnYjyO6p2ncXnkZ55MRGv/O4bdfRibM5h3p+it8uS9/ui9gTKagoPGkTgIiqQ4M
AMqEoHBxf2EROwdKw9AWlnRJT2sUntp6tzR16w5fUBf6VCpA8rPB/SL2mtXN4umC
rGjtvcLazr+Th2KrVDSGi4m+oz/+0PfSeDqsgS4jfG5GToY8VWwXLcjf2c7ElIBc
26D08+Nc9H6JvTPtzFB+KGqb7EkXML4TaR8ERBsKv/xP5WYq+JWHFQ8w0O8gvkRM
TOfAChLNlc58YxYofepxzernjb2GQWaNdNV9qvXzLbbuti7jeBedu5TNGiYked+4
V3sAQVbJIlpz/poYMQ5FWC1X+i4MIMZ3OKNyjVGdoG0mYfFX5gw6DdTc7Cg/Xv5N
J8wa+h/gUXnKKLX1rEtv65X3GQGcuIQh5Al9EploCHA5gkb4PLPJzAgW09XNz6NS
AjowXuqCSC5LX0ZQB0p2rYuaT1lQgJpDe0ivHbhN7l54KKK2zPsWhEnBhJjtPpmJ
hj/xRJR3XvLSZEDvBLLd71PIrdUfhdV9xdxC+Fp2xPnKOqptmRNOmZ9YLWdO2bcN
SV/sRDNBmYUFV6ymfjQ2CnZ1KZMsap+5Smy1J2ockrfob+itt9quqgwsMBALymPp
Zt02/WZhy9SmEx0PD9ggfCAIUR7uSiBzeO1IfD4k9q89D1BsyTOvAfQNENOHhT1j
vvjf4h6QT4A01iH0XSgpFCW8m3FroBflqr2XDljMniTcHRapq+XPLZnfUXgkKoUo
NWzOxMRp1ZZC9ivuCOJggCSS2TvMp3aY/V4UdFMT3Lw+XI8RtjfpPh+WTxRD0c6E
qvyRAQEHMUnqNB2A+HnPNpnhh7uWHI3jcwR8S1gEqihLTm97vbU/mChBC7to2O7K
uUN3cmpJLHQ9E9RY/xdH7B66We1rohYRq8W63HVAjhi/bYhrxPkJGnXwDNTDhlFZ
VEDoHu9LleUI8W6NBUIUCwypk5Lv+FjI9yhyYZ/EbZXj7HmPxlbQ3ssldkFmxLhm
YMa54kAoTw/aKjE+XXcVuiHUzVqaRCCacM7MSCtErWWrN2B1EENsPHCztC81rbzM
lEBC6JODyLBMf0HkNFKbFgskwm1rveqzDiIw3VilYDgj+mku8YxeAaBKTWFfx12u
THdraecyv9VspcjKA0comKm3vWI8aFhf3ekomGbX824ha5MCcYp2aIIet19LPI3H
Z+YkigAubqAwhCAMIxy3WCUbj2fvhMRYEMzKajHXeOx/veMlGCRbmYE9+lw7l5lm
bA03nvnTUTce9RBYw9Kc9feDu3wQuNSPP6vtM/3a5MnW9TQmw5EYdRDIg1Nf9rec
IcJTjVgY+ao47NiNf7LJjp0Ua18qEB3WEpaUFE6jM8U1X87ATXP1NRxRhNJW7yyc
k9sI83Hk36BNFg9kJbsKeWjcdP/3igM/I8XetEXSHzb2blYuTu1S/uYiH4vMMH7R
3iMHboVMGr78DF2oLwlTiA5oB5hITlQN2iZkSGEpUDKP87r8kdlx4DEtMVmw1Rlr
ZKlbL8HGpS9+Evm7Cj0p7Wp6NocWfCnnpBxlzRl8d9GVzOR/DmVPy9Muodk38rV0
cjUBqDyjswZJLMbAciSLqY25T4CwZJlZjM9qMRy7pgGVGfvTVURnA7dVEKINJf6e
J7IWpog1aJ+5FGTtc0CZedkEBxtYpa5rityaRWl/OeIg47qDHSD3PnmrGHouqlXL
MzWEKxO5nncrAg6ncMOHVsGIA6pakatSpFTopieoPu1SOa4x/SI95GBacDx5fU/z
H0h6vFAx35wigQ+HF9nWUzboGrWYGSOv6Unk4nOgXaCFNB1ypbGy2QQFC6PwrMEf
5vPcyAmOW40eks5AAquwbMV5e+0iHcm92Iv826LjrMf7z2i3KNPfCdtI6BOeV7uz
sa/r2zUrdcA0N19o3FndhNwrogPtQIl9EsFS3bdqwftK1YObAFsw1rFt1FiUsoL9
o6OiR1oVLMQgCL9VuE3flf9pgT/02SQnmgaUEfyj1eZvP14nw4RfETHsPNznq/zj
DzDLp5oUKjGRJU7/ncAbE1/EcwrFQClc+gTANONy9UzUq7VI0u5M/ASv/96KzKok
WJc7fAxxE94X02LkS9PpxI0kxNx3XS+no5MkJZZu6XY4N/ly51bPTx5yCv8Q0cD1
NKkkKFYRKvfFrfkTkSnulC9VB2uZfo+DThuHHC7ZEOnda4x6nO3xmwXA/1hFwt4P
qx8k8z/7Qq9yTTHn5aSxmOTEk0MzuyUJAfANCdg5y+BLFJ/O+dOXF2jEWOKiv1pc
fGH6zn/JVQyveoGwX6CvCSzYq1Epjk9XWUwEWG2ChV0p4bpmyk+2qNpCJfZFK3cf
hXtb1Nxr5J0zomfAhQGkJpT3u0hbt/7BX+rw1ou1S60+UIYsaj4t2/RN9M/Dz4zK
qBOFVGjdFwmh0AbfYfBdUwGF6A3nbBiSeXeJloaEDIX/yPcKyFWQNo2h8zvwFdTx
kScXR9S7897K2Va1WT+tVPluGUpbbAVnb8p/c2TxZp2Kv9yuqq0wQp8XbvoXioi4
idGwNyi5SFu/aOmtkgcPlBXyXgyXK18M7X1UKCZY0XZSUh12PWw1+G8GxFqsp9ER
SoLDWUEGVU9CG4DlP0P6r9pzw49EUmnsXEyPGpKPgoPS3g2OzTyWMWgBUkOUmSOb
80akLR0B0yuCagI8i+3facUSE/KnZkejgmQZZmU/kLiRcCndyZoZnPhZ6jfSDxtb
iPuK7MocV83yylct4sAyh1+cjcQO2nEZt5XsmJTjO9E2TmodMiaErXZf2pEkSi0I
B+0fR6eqj5uvmNl0Drn3P9kftcATAMSx+tQ06NHD8Yk3c7h7CD34sGppnaCh7qt8
CjNmwwZyq38Xbh33YlaVyQOUOvd3AriiIqo/w3vxDforUU50PkhyWcbawumJXajX
d3VNCHyKGArsbebZrlaTMWeI3Z+5V9Q0EndQ7Id+oNY6VUeuH+r2ctD13Lg7DKrG
2HcRfNBlkAUYgtyw8U82InaPB2ZYU4/41P4YG2/OLUGpT7/0vg/eSjDaH3W2+Mzi
N+pHXOsGED6vMuvNgKIwahJQF/CLTGDPq18e7iivyvtl/cGj6Uk4hbhbi5JO4V/W
CojDshtoz1MHM76ZQkXfl6kvbSF7GC97cyDcoHuiTPfnEfkycXQFFf2uRwoJdWTT
wDLm+sW0yqZVRbUnJSb/QgNrMrnaMu7HnV65NZua/SDnK3mxExuoXgjgCxMt+Ns0
FJcDEomawp7wIU8NVLFkp4XHoKom/DyvD23QT9+2iTx/Re1s6Y3l2i/itssIBxgp
YGygpMwlE8PwWnqIZdheetdPZyRkl2tGJSkNfGtO7AFZCh1XGchGiGuG66uIIBhK
RcMwyQsDjP/Hd2dcSxDjKtVHLPUfABNg2CGNabqk+deHDKv5JY/8BxiFuTz1MgkQ
h7urlBrD04feK2jrC0/IOfX7zbWYGLcdHSS4brKpIiAVtCXJeQ8PC+0kdprHbyuY
1CLhaHNabVcorlNHz/AT5WDhuntKDQh0cDlQw9oq4+e/BHfYu141dcL7CPXMP8jO
uzlsaW7jXlmiwIksPvSOHsfTcg0vC/R+NqHyyeetWgek1sZcAcRlThG3QDkdR1M9
BRFBa3Zt5iaHSsZlYV3Me8L1VMdWNbIdyQeCg6iZyg0UEsFdTWjQ8VU7ByR0GO8Z
0eTUJx5C0ycumq9ATJyxbkxaNl55zo2e5ucyWYWyWI05FqcM5hwqqyPzvMK8Pw+Z
+rqx7XrPxKENDrEh6qbc0t0kIu6xCAnW8RZH0/42NFB8jIxQGLMCCYIM1pVrqQCp
yuuJfKR1gqxX1lPS87TKS+TKHL/GBz4E1TLoz/i5lVpwh0ng7IxTSkRBX/HYLn1h
+i8FzWa+TXhsYZ6RTzhwkfplyeU8Vr0mp12xhm7sfO48ZqSRQYeR8+2C+irBieHr
Mg8qE/RihBidnylHQ0Uxqn0pSoafEIfVwLkVFLXAYtrHniHp40+90Xt6cxIjXKK4
Negr23B7bKMx96jRimPfNZoApbGI1dVqE3d9VIg1/xp9krpgPUogFC+vRJws9RdP
PETF/mk6S+eREuoDMnahT18wCZ+jxDF/6usJfK5zO2AmOsAeMehmjay95R7lieDw
kjXKBg16XrreXRs2RCXklE8EiwkyaAHrZzaxfTtx9MFOc/zajdBRSNuWEi8HX9tS
xKrIer0V2QT/iV11Z+zpK8ooGpSlmg+H4E/nne/olRyoHtbM5NqYEC3+ayIVRtJe
bZ/7DEN7G62jbkXc4R9R08cOMoGBrNqAdvva6qcZowTe2A75CuFOQAxc+C4eagWN
LcKCuU6QNSrJJxTXbft8xfYH1HCwsR0Ot+FthycWlfOCrswgDOTTR/REOQRskRpq
gMHuJHzrjKw1gyAYpVLaRJWWu5vgzGJlXNp5BIwRMDpxfT8zOakuMxfNYsmSdpKR
TUeezBK/zXoK0qlY17qoXPG5R8Ii4DwzV0BN0SIowIBX7autXPp91jB8wk0U0Ugy
quK3K3AgvlDekoCwa7Zqxk/opqMoW/TfTgoKsBd2eg7XLx6sXECHzbZhBxjCuK/b
rlx/8z9z+WmjKKsJPcFy7cHOSE7CARwx+kpZXDWRgWMti1NdR8M3PP39beh4cz26
7A/ppMJuCbUQYJROdngeEMEL5LlfAyNlGEbWE3xLc9kVWVM110A1I7nT7rdGNRRR
x1iV+yiGDZEbnSbonuvCOExTqNGHmGZRi94KL7oiohbWURiGYE7Ag/d0QUo85K/g
w+mXHD6cTsZr7gRhU1cfuqHBono64qMN+BGRYpAcnJbOccUEbIQiPsohbFkd03AC
YOx/d9zQaO+4638khz6Qbm3Mka3dUxTHuR5KbcaKynRiVZBRZ3dAyVgZP8lMLA5b
eUCa10mSHC7uBlkaSScMTBk9aTlqKpEy35gq1PPft0eoLxfU7HjflSzo4mEAgvGc
ljK3u3oWnkhkl6tEDO2M9oIC0b/YekdzLWVfPuclsReoVM2SRDbaKfvNuEeL4gKg
vnYRlnrCWm7uQEKsIU30KZTlK9xn1FP7djVFD7cc5c23SaelWVt2KMZy6BxjymGZ
zRafJ0EEN/3uRzDW10rF69oWi0kndFC8vuSAAXVMM4tCV1spfpjkCUDRAcsVXOJL
yUIUJ7C4xwfan4SvUqY/mAgpjjBGP1kzbBxKebEfy/54zND88MKhGQWFMLiFDQ5z
2x9zg/LLmEpz3nnHQm8E/1slSXLSNNCR/pZ45R92ZUDJ8y1m8lYg12BItqlH9Zq5
1XescrJUM5vWzcw/OuCCYAB/35i8Bjh+7ggaMUBK+KnHXuA2R/NISrA7gLZ0/zlU
x/A/PE8O3Kuv5QSDiR0/lWkVjFBnjJpmdHbmImriqP6EdTgENXpIWofftyY/hpye
ZSA7BQkaSxw3FMeLD8Pzxz/H6DSZgIaNy/AFYxHIo2kvyGMCH4acKVAzipekWIiW
tqV9LI/wy7QzrYowuhXKtS8SDnHS3D1pBrMfJwzXSXtUuvv08xqydjzdwdmd2b0f
RR6Niv2aejLG5iErQwgsp3/kc4soFlWAb0mjqi7Xt72i4Alicj/MlTPVdH0mcvBO
gThE9y3seYqSpgCb70qWAozyyJoPgF/BtHsJXnRWak/vZBaHO3TaQGQxvR5LK4c6
btZ0xIkHyHAqo0PTWRN8CtwHg51qrTjAuACiYiLEHD6+WHHOzXQc44rraAtEXbXM
LIbSNQdMbdUHZNzKBEmOP/SWfnbhtZq7xQnOB33/qEfQ577qd5o8Z8/b7smBO0Rd
BCR3Qk1vmFRnen4iX4JT7nvYwFPLK2kl9j96iyfICfwbaLJPR2cKZnen/3WKMr6g
LUIm+hZtYEdAuydBrgr+jX/e77OoVdDqE8UuTrTDZyc0kx8iqUgXvEYloQM511B3
f+TrjlIiwgsEMeRvwypVcGeSqaePNnXnUnfobL87Q7d8dL7Qk8h8KzXcXpyIKVAU
qcq1wEnf4tUJlvDtnNJMjrHmcIHvC/MasnXX4Bi7I6r0hvaRyIprudUHRwNpXUoL
Uv6928cQaWC/TqosQFihSYzuRECR9qILExk8uKpCRqjNCQfkY4xCYffPN/oOwVUG
aLIa6p20P0Hu3GXpF6ApDicFzpWbpduYhwBKd61GKrPbMYlEgjkumbG2JbyEMyxN
VJ8tFUszdj1AesYVAD87aZoDP8xWH1P+v2wLi5Y09nUSd3MCV9h4aTE7rsmdBeQZ
cVHOY6L4Ht9NpHMy01MaLH2nX5rPJH4GOvmv4R6OXHbSljEReDMYNRcrDGXhgifo
WQasFRAFkiNJJ0+kywTeNkrolunULDhQ73BISECmP0nSQwl5MUcDy+5a05kFovCk
mann87HebTvD+fbAh3b7tQaou1WKxgQWv2rRQAL9Esb+qvjbNTSOSVqaHW91drSs
uz9lol5iIajXCRydlfRI6tDXoci5HjkGpEDM+NBNgrQjd0fMo/IFMwGTMjzJxnWU
pfOVSxRHuFyJvVbt83756KBm0zBFYrF2hpJ8D3J+mnwK/alPOedQ4GeN9zZpE4DI
MbeSH7Zcy0KTiqOybJAA34exrqhp7sZ31VpyIq2plrkgrl6FQTQPvTHKP6GzrGcx
YU5xuSVjZjmd+IOBXE82kBrGGIacYmNIEidNtjV1T1HvZZ/8aqBDK3SnBrcf8fX6
aLCFkoHiUGrdKqAwAf51e4td1PDZUZF77PS7U0Uxygom9zA4B71WQ3baMkb/XpMr
0g22pwPFQ1e2f6jt9OLZgI3VVWSKgkZ1Rh60toomb7qVK4cLqzCD0IBkOKi81Hvt
lKY+OlI1TDPuzMEB/kDNAg4PLWrorTS1jk4O7ddY5uYSkUeflQnezqSXty/xIG+a
KOSW7Uf7Yyt7K/DG3n/Ddb5V1ouIGF1QQcKEMkseXhBkH0f4XFP1N0hOj9akAqCx
3OI+fJ1GfdajslVmYupOTcMShvD0DiccYxqQ58NkyIWaKhrlHUKl83ua697TNAvX
Uh5h04eofojCzBBKby6fYGrHScgVRCU3uU06sDn+CChlFyG7N8BDVVD1p69f0EtW
xcgFmrvwQ71ThOYphraKUoNK+75aQWLIDRhW0dGhd2NYTtUlpKKed3EjHlIEZfr4
wDmRJsBsSKdr1/PwSJJaPRM+wC+eGWPBl6ldv7FVgjQGUJy5E2xHWOYGPSWtwo84
D0o36BtOVJGlr3MOIcI854PYwurV9rtbxOEGR+z5qfuk2pulQmlpPoZZiS6fU+qN
8srJ8R8PB4C0RhdCKJMytvu/XriibT6+wrXMkN+m9s1G4Van5w96KA36708eshCP
sMlVIlZkoggpIYboPHNHqp6ARZvEwGMfHT5gMrbTenLQ/Lbg32z/onkf5QIAQsvE
bomA60+1t7j/twxiOz1QGrgNkgujHlj9SpomdcnDxLWuZkv4zKqFJhqiacWuCwLD
tzlhj6/CWketL/X1y93PFuqiPta5hLrShscss7qpb4s9oCVuWwZZKgbY55RITw9z
khnH1LlZN08mOq73EWgcmLT9s3ZRHs+tVz8AnRZCX6Cm1Qo5yQBNxl4nH1y91Vz6
j6Qu2fpyF3LRBQxOuescGSGdwQSKyDBxAKtvKfEXioX4agJKNlBHgBTlkrrCickB
eFfMo3i8bF3c+dVAi/l/xCY5AbnN9mTbGkWjFvrCkxOVlfH+rMK+oPWkZm/cWNzs
kSWucBEPcYPx342p1HCUaASjFWnJsrzUhGheeXZ3RNR0Aq9znBejWQf01Ye0BO6l
y1WPyVgk2OHzJVwp3shMMkRJDwP/uqQHaB2iz4oBtEBElAUQy8SSuO8LlvipxNJ3
sM3bEoPYSdLnTdmHNiq/O+Wyh56XEFtxtSk7Nd/TaGJpeg3ooonswNZf9peq5clT
WuLMaAEBXmmFHCxJbR70rQsWQNZPg+Oafqz1PL92o0uq2O9caxRXamzm2BgDxgKE
BBeT7qNJ7w08zBc9qVSjmBg7g2gBNniDjm50jXISCApMU1PxFt7i44M4zdjI3VUR
JI4i3/3zL8gqqIKzOLCPw1ON/Hhg+kk+2VJWkWJO96vemHstiSiaLbY5k70C4u62
F5pnm//FtsctGcf/PxfDqQu2Tn12IpvM+ke8WMu/aAoEHtdOgyJHdoail2KDYU6a
NWVmkkEJMlZlZ683l/dLqLs+0mf0Lo9sv16lxXJJCu2CGOTnae+Q7c02ErwhtXis
/jYTEMrYgPBauXMNwMffRwClScWRjG8/ep7slHIStwgGCuFR1rp7wDc7yUhTGx7H
EGwLFIXjw79ok+HZgE2MndnvA3DGfjrdBG80snKByGPMXEoce3gToVjAJa9YKJ4p
PaB9cdAkjCg+zpwE3UF4/GrajmBe6el6bAS6+b7XoqegCkHIUbJ+y9Z7rMBtRrhn
gDE2Bh1QZQEsdQn+0JPgHXU/vF8sE8XP9drO59pfxNshikv34WaxG5pvUnt9sCCa
jUYcb1ZXyGuNR2xE4FLlPWoc2BaEzRw00G8CkdHD1EsS4RiSrH2dStrcP2gTep7B
qa6aKe9LVbbmILJ9Ne1yhKzXPcWZmf0A9iWG8RamrnVs2/1bjPs8OD1Tmim3D7UT
lEXmhl5XOZnmfTma9xKeS/l39yXVyChvjbJWLaAfCGKyXB719SF+cn/FN4wKPqGr
6BYO9f/CBB03xDHNY0HEj5E/y/3HWHDFe45ttVxUxc00fLr9MrKk17MWJ28i+TfU
gv6dbvs37rdHXatw6K67QJ0pWc8likq08A5Pqkoie2tqyu4RbZ9kZDBFIK9zajvP
z5Y7zC/cxrwJ367jxvdoraSAgUNOZazx371DKpYXt2MjrEY7PUtA98xA935teggg
yEW7kZlb9SZ7gdU3+PppQj1fK9FNucOn0wMdGZsDjCgqwN5Yq4FHzKHboiI59L51
gloG4A1WvxST+G+XwD1qlJ/zwJD/czcx2kjhAUNIw8oHvZDgpBcFKb0mQiKioUMZ
dCMbYOr4MrdNKMu/Dn9AQhoIxwHu0sbtgIlEuWUMKYZ/fdNh277GlNVDOc//wl6g
qvQbvPItALb/rR7ZcH45s+2USKLl19gTMo5sG0Ix28IwvyTCYGSQdCNHPFKZoRXd
Yx2U2m2pDDB8sIB0Ae9NFgFQq6KOBLzme5LKXfyBcQHV5DIotkyUK+/7GvsKYaDU
wbKjZ3jcYaTZePQIMEvqOWxGH1ZKjFVkp1LOx6zVeBrmCGLtcYTaKmlet4aEMARR
WhsYm2liS26pgOEfVpG8ZW/nK9Q08kQWAFsrueWmNg/DAmBi4mVSuh6yv9KSGlpA
bfVfh82EKDAV0ZnnwpCKVnen4GWa++tclwe+J/qzryuxPQ6RdRwphKow36WuuqHP
8vwXbUi48Tyw/qpW6TdC4ydnYG0AyfdcfAqHzyasEHayk52Q/IdJxasjAt3jtsKz
GPoExUgyItcHkWdSodTbMdHa1U0wZzhPn9dtLz1XOFdcVU4x9+KkJ9lIQly3Ttvg
+2QDxCqKPa2R4REDZBVqEenDiAKiuhShUtvzIkOBJ7PIDoUuJR5kE7AiqLiLv2xh
iysLS2ArAodSIe+ESi7Oz3ujHFbUENHsobNa9mcSSqNzhBkHjMJYKem8QQkAQPji
nsX5KP1JATN0EkQRHOVssod6kUOgVS0c/Icosh2Iwta2QXuGrsKPgrGJM8jaU8ar
ktxDy+hqd2KmaheO2NBZPfZm4uXgbI7g4mHxxciS95/8vzanH6n9l887XBEZ45TE
PTzD0Am0smmIK6QtSwP2kzDKl5bHeLj3GVXZAYDsvnfr8Ww/ODZgYTjBmgmrqNxV
/7tMfmdOfLfHIHOUpnzHe8o2iJ1NiBGRGdqo+moS+DylfrjAkpFkUir8VAy+gxjN
57U5cEV8k96fFAwrxM/Pq9m+gRvdx/lEnzf7kkvfc1Tb1HZbDEhsixX2uTZYorQx
MNIrR8bbq7y/9G7jg60wdlT6NtHWRXPoKp+/Qw3JdINEF157M+CqWPh/bvYDDvyu
Nl4vKoYQlUPlX+2U2NGvAIWUJFCuGjmATaQzZZc3sOGIckvmIztdqzE2cWhssheX
wwyUdRyuMJf18x8PtwHW/goFqhIWToN0gqwe03p7I/F7lTVvQDEFKUi52NfGfTGU
u5+RmRDF5wRJ9i4qyQxTAamyN+zyiw2B1odSBLZ+Gf0V9OdAGQpdx4LXe4BAz0ol
jUc6hyujv+q+6Rdkv1mVkQsiMighu5pZCqT3Y+vVTnfwc3Mrk/WElg6zDXKvz1uU
o/3oqlTnTa2QpZ2Nv0odi6AExnkos+pb7ZwaXLuM9obnAA7jFXBAK1vsL9nqRLAU
QkL485ync0BOibizvD8WVM2TwA/VRzST69WCK08Mps6IsojbJ1yWQV7oVi+OHPbL
/mqWfKP9sm1ZTLD+Mvlg9xxi46AXorpcGeG5VlUOEmBy/t6NXbv3RMQrYePJs4cO
MycdvtJod9qRE8a5V0gYEPUuAd/NNxsWGJDIU6zjL3vhA1nBkgduH/H8QFYcebT9
g+2NOhmmb4cEcT4sut82sp9tKdPuG3f0VVPagSWlsyfKq7jhJFCUWw3cAo+0qgRY
hkKH0YhvJEjEPRDX1dK8ndoQo1aO3CGRE0JAJGscKAa6aY0pRHQ8hvoweP6GdBHO
0UHXnZ7E1wNKcacMRJvB3/YSCF2T4sQekkEeWhKqevRivZnY057Ho72zPW11+oUj
CZ/dyZOcv+6B9b6bJEhntP+LB6Lobo+zU0xfS/mMysHce+VDw99hf+9W5EKJ5Ha3
gw1RpZjdp3mQ4IqmnRVD6U5uD+wOXxmndoKGnnPrnl8LIRiT05bEaQxLbyGjZwiB
co+MGAEjnrv9ZyiENFW8sAaU77g3mCBG9WgVrEfyY7LqZzE8m5NxOH1gEANqBMve
LrMM2HKNhG6GCdQu26j8jR06p58Qu/qW90Isi4is2QHxOSTJb6xEIdchz4UB4gMg
SNjBoJIswfEhPdGv5IwHna1F8LUJaCDLnpwZ8IYS7cErRJ91S1enNXu7pPptaasM
rg2pp4J7UxnI43o2UFdcx6sbowPX1WVH9L+3SHXmtO+kILyBn1OWdFN/ac471EjF
X/pbsUjj61XwATHSFhCktZYR8TiOR3FLKwlR+noEa88ksqUDnUnBzDgIMIVm+dbA
bXIO12ufO8YX9eq0XyIbj5rZ57tjl+pzFlPyPUKst7ogAngtfqvQHwtAniPV2vWa
b43FRtWzmVqawvvigeQ1OdjK3/OLEEvXUmkuxGCvUjR3McXxHfN+mEjLZlGKJR7l
I8W5XmQ7WYuYtg6rBgpLQRLKx9HNFkce6iECvXN1ue6MaB3AQ1XmiDqQvKMyUd2a
F9h5JAJmO3iOUhCdtLu6WxgXxhyl86o8qpZ6nmNiBJP6MB9C6MDv+755YCEDaHs8
CHTl83q/4LCT0hJt6Tt9R7l+nR5VxbY8xsXfNG/G6NTMBauHtIfZhNk5e6D8vIp0
Aa3KwJKuAkGXZUbYWk7hS/HYohBdmQztztYsSsvGfpAh/IfDTC4hCh005S+k2D+0
5R/RgzIHv/voF3QznuVw8YF5VpjSijwy0NBtCT2flXBTqUwKfXqdzdymyOLwqs+p
NFLY+8RDtzIox0H5FvpnLlRYr6r728YtNnGLj5yTQtCd/HFLkP9rOt/lt79i3xK/
2eD/sgdWLz//LuGZ5qwaAZK6ITowq2+Zjfy9IxXxTl9mzta7vA4nWzW/yhb6RvBM
3wuyxFEAhnThVzZbJqSA5xb/c3RTGd7crMs7XK/1a8N7dRXbolv882q3whZzfQRG
8r/KixRXqPXmByrsWx596aFBtyRG82gGnQ7LrDScYv5yaPxZCDW5Yd36gFNEjrqk
lqUaRe3HzNxnip5m4TNN8kAxNfLTjd4Y09Xz7/4dTqzlfVf0+3H2tiZfsVlcV+m6
Q4XUku5Y4RvVjdNZru54A2TCzLsQqPUbT7R8EWCcVcvcuRfapLGJ1d3VKEdVMn1n
+r7r57tZmnFiSr4ce/cfO8W8pdGzr/W3qw/ytSWscUzMNM4JI2TIxudtYI3+rI0M
uxkJYl54FY+GCtUDG5yczhKH4u0yT6l3C89FU9GDm30YYrqSNK8tVnSveiOu92Nc
MMwMBVoXeVuLyMB1IaVn457bAKM8nm+4KAPGs3FWl1eiNjGyBVwBjghFXSkT+gC8
+DYpEgxvAOudRaLDgrtrfIGqPSkAt0XRPKLVo52AehBQc5gH08TAA4x5lL6WaM3B
M7Fnngh5qYWxyyOaIbOjJHE6Lf0lBEeiWfE8lt38D2UlKAFuDoHbsV18af2UQtaO
1sABn6o7QtcsZQFOp0AZGQ8tn3SSIZRYPQAfDRm69uMt3w4gPCupbLKVltLckvXx
3X/zVkpneYPGrdhrUaW4ozI800g69UMGVl+SO4+s+ELvFgs99jmccEl7ETXYq/dy
JOnPr4MKdvz8y5cBiSgBMqGAbt2c/DcYggmLMjS/FewSpvfJ7WpnXETo1Zg0xLUQ
5nsLxHhvTGsmVRjrRBIQA49C7p09KnF7kGEj4RYHLIjmRlxU7CgxQC5dijDHndOJ
/R2Cr6ajEvfYqTgKPoSZaECqX62mwC4KwfN3l9zojk118uPgCDh/l39zjnnVz+cs
bMFj3i+FxSrzzlQhscV95dpflYuOKIxUAYlOdRqlJi30dhhdJoQctjE5ggy3coVZ
moOz4PgrnGMuksq/I55BTpJZP8Wj1+GQ4+Us8Hf+JxAdStUi8kD9CVp+1SyPpjqX
NF3Hkgj3diPTNxfJhjRenjuzUIi0GB2Tu2c6iAyoxLmo9T2eAGLOvbc5CKUpyMar
71v2UimCnAmedojTN6Ee3XGAaOcCd01ooPjcjJcpgh+SeXFOZy+45kBcXT/2weDj
+tAkFsxOnpE4DpIJdnsoOXJOGnEfpQdNE6TtAxHFpZW6XFHoJnw5lCs7sKbIgt9b
G1Rl51taeGWAyl9TluyEqb1/HQjT75aKUjGI5qcZXVGGv3qLH1Mqsob0+nSDOzFQ
/FAr1L/DFmWVOdT5uLXGEMArQ09LxO2Ek0Psu8NsM1jXb+vzaOkU5DRSVlhf7BcQ
AUmB0m6Sbswzhu91sV1U5iD/PdMt4KfI3r7y15RoVo2q552YjxKmMZ9Q2bq37PlR
H40fsylRq9iQAt2vryMAKbV+QNig2m0XYn4esGHJV7m0euzazTlWOql0A1Lzr+al
VHqSEIVhkPVioZF0549xYK5ioGNgzFUs6ba4PYQe3sGMfpNsul2d3ULU7/Drp2ix
2J1Hsi9G2rpPQf6T5NrV+RkGZKgHUjIdf8Y9SSH+r0B6WMVigucAHsd6eWYQQx2b
oGE/B1c90chZ8H+FVAywcEiQDDqE7ORCFtF96uJTc3MXbwVfBxHEu07Fw3iy5xhk
xS72suqcVyBVQMd08bBuD55FghLAF5c6noR4qXGjVIuEY+UIwX5NEVl9FFgFg+Lw
QuDn88WgXvC0dXR6nGgmPcnRbb4vWbJE2LwmpL2kJWlDAr22Q+yIlr9SRO3YjvFQ
gmn0wm0TKTuvoJHH5AgeLJ5mux3aDml6JTWEm9OzY1YmeP2rcxlEJrLidrmdp3BM
pgT3TtBP4wTNIWH68uflkKbsltUwjGwnBb5XnvPDPDgOug7DSarfmKNJgOPp4cWX
6op6ke78JE19MW37D7KHJ455b/qxMTQFfT2kg9GF9qIwTLr7BU1WD2LEYT2pqhf+
SNuAhzj1gqbdt0MZhO6mZj8vIkUzRUMU77BSYUVV3Xd1ph6qW1ZQgfFqkkuLvj7c
qgPm1gZGHkziSnvxd+MzdSf5VL2f9KzkXOlXOHd/W3ANle2U1o1AD5/q7g206RU5
LJ/SPUwR4/DjuTh+I4wH4j6qIvQBxBP2qV+S7OioyBdEr+fDCPIXgpjnSD73aPgI
umhGsi1KT7BAvQCgDpA60asfmRdrS+7rIKXI8aOOIRFwA/4OvWuVCa/VNH/iC+C4
721gOSJt8QQgnTPO2KZFJVtHJ+ITVQDo3Klz8zxzU35iAiCkzrLZUNDWnrcVWsP1
63/uAz3/xG5Eiec7Mfku69GrsmWTi+5rer1QH9jgx2nP9LBB4VHe64QKO08QuQzg
QrmUO8uD8AmzwFYkC2cKx/dpT9N3DxyRY+oGsNS9YG3d0hzyKpBay8GIVB+wPrdZ
bQJlwIZ6fbS8aSNWHpLZ1wx9hxB9eSJIZniJyIKmNCBl5qvy/fcs0fzDtCjpC0fv
wAlsCLLXKroHrIPwPrPzGjcBIbgybt+6EiK2ZfjhLxqNC0cIiwGjWtF4PSTxhy1M
Ca+GzZjhzsRmlAuFscSKCkuvsFez776HceeVFbxCoe0vcvQp48G9kNxrqF5obcgF
t0SYtvIN2kuIsMXU42Mft9dNH/syAnoYDIKsYA22wGEoVuierPa7UPYqdGbd2LeZ
3qFVkpHAYXbfMLz9o5OqZo2cizbyu1hQn7+uZom7s0zZ2EBkbqaaVAjvhtTAgdXs
DPdxBbPO+dO9GBRuRDU0sKTnW2/dMHiSn5jOKd38TuHBtSUhiyZW+ziggxRsKthO
EzvfwQY9zzaFka25qjLfZPoUn+cEBQ2GIt42S8LHB3BIwtCovfGrRcnaw/0nhSbR
uQ+FLdy5EuY3DYNFJJExnCJaap4CDgPa5JwscRyQ/e8nBGppHuLHZq/JGEMge9HZ
FxN0Bwkw1xL9bka0iCsRCWxtPF6uphj6uZg3uk+REr/uguH5Tcc5ZGipzUqDyvwN
auz/soVOZNOdeXq1cyN9fW6VJ31eeCOffvE3zPdwz0fJlSZ4A1ywi4ZOoTYfkcKT
VltCXuFhVp/pQe3LKs+cFZ9Wvhn+Jpk0VAjVziUXR5CRwtjhVNw7xVa2Kaf+oqJT
cKxFdH/HWUZ7uacd/q1BOBWWAxKHP1/J8llM1n6cjL3VSSSXn8NdjTdJuVg5gchl
KKzaRl4yagUROipgF2tNenMCAKGN3izvsor0ko3hTZRg3pFX/0zPm8zu8VO39gHa
th5Y+Jrz0Y8uwjpZimITLQ==
`protect END_PROTECTED
