`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cperjrEspLs9mngFqhgMj4jXwC7SsC1B//k6JHneYJODbfpnDaWCj2GYepLiUAx7
yLYYU0MQB5YBkO5KrQq64MyX6keniyiK5P9Y0rBIHWERdfeJfI18pl18ZAUjXBqg
hiXA4O+OyqEkDY+j3UOtenoUH6VnTPiVPFb232o59IE0hBKPteqti9oCawq9S9IX
76lBDj3ztootab0gxECXNiki39PcP+F530d0FCMQwmc2sZvJUOZfG+MIaLAVQITW
DHVc2AFyncEut3hVBTnRJbg1HBvzjy7QS8MyCUgJH3Vyr9xFu3Im7KbdoJzWU3SZ
UuQr5dE06pZjSX06nh3Zul6NLD92q5ZnsuYZ2Vho/8A=
`protect END_PROTECTED
