`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z2fJQjBXYig79EC01v/9D3ijiKR9hfbA+hsP/HhY8nC5+bu8dIU0izdFaA2CX30B
lalkZ9q7e/nVj3mBDvmJCcYtOnFxw4QQc87khi153BqIfshxIvnWamcguTqjR+A2
EZZqLFRGEQpWqHuKa82xPPmMXLY3vZxLPfgdsMniO/xYRSuzlapoR73KUICJivzC
8BtolNQZ0ofNOobbzKjlEAV72ya7gNGr9RjOXTNwpC4FhYT97VcQ2OKtO8VCczIb
R4uwRhUFoHLTajwVd4dOx6FdLUJInndU7SGc4qztR3saaxi8SA6JWJS2DV2dwwhe
2eyztctiikq8Dva7xegHb8w+vgEGBRwGVC5VLMatGmFS8mNXVF5uXnAPSfkEu7S4
SCv0dThxKeTl+FtdKMtBk5X+nGODH/NG/9Ad6LQw1YQab4M218gMjqx2vpoInOte
9x2eK16XBg2UW0tJwUp6w7AlI750papoLrdNNjoMFez2DZyWHc8AQsVo7pU/OemJ
5kR7BEqDO46oEdVOjS5Z8k7FLDILswtGrCXsL+YNDul0axbkbmyc/RHZLbxiayl8
Y/voMg9eG2lZdEH1MWShHPygO6go69kUzFwwUISQx7hrIYncmneDhikKpWV9fpVc
Gz27j697knuPCSfudF0QjBwkQJJdzRskX/Ac5r+eT3ZMoJqm6Lg6M8WGxmAgSlcV
dYvQ4flsnIp/mfFnto6DZC9bB6fvexsYwjTSHEvNHy61qIetm2mq7dYgy5gs1n6x
kX3HmbrS9pO7x7Tf5/t4vzcQjHt/sQhhQRQHPEKvKKx8JFNy6FfyVMxDkBwI+sqk
hMI3ReaoFSnTi02V9ysOOSUjvlhaWN+sViUnAoOmja2Gwytsc61/rQ5c5g1I3A8J
hzmuAfBNvXC8mf5gnA+3MSsLStFEe/JjiE1JgA2bMVG/Ap7cnBsL7G+qCh9tM0Vh
NwQoT7Ck/YqSQWePSitXRy06U4r/OQYhKrBUqlnEvaZ6iFbWaZU1ob3FhxHQteUE
E2//rJc0BdsJ5DNi8G8yGYIoE1jlBB4/EuQb98mzFUkiYgkPlciGqCixtL1ppUmX
OwiEg2eJnQ5wef/XCuWBAx4HAI+pJewlzUd+UVrxfMNsoQRVbDgZNHBmYeGrB+Bp
Q5o1wNlmUSvj+x6UnOLjKF0lyjj02Tco/dej3iBSuMADYo+9X9TTrdUdQztDMvpp
7DVcVVXH7gqvL7cT/o9vUL4wnkzOMCXzxWv/So2ZLI09JVSDRThjg9MRIK02650d
ajOhRT7bX+9951INA4IuslwFBEaBUKwOfjRTQxSIrvhPAAfqLZ7GBqm3YtYUpCov
F4xqzOt+PNah2mKjqAE5pgRHrFc+iBFvt5QFUbhH0B8+Nua8/SrA1jjARMdySyld
Ay/OwogLPGfC14pyQAoKkjEoTc5D6n1q+5OdizIPbxDuWAetQ5onJAoOFnH9GwIK
oj26F7S1zYYxSUcjzs45ZXbvM0PMmjDa3L/GkIQGj2nFFh7md3nu/P8NKezk6+El
xQzKnjj4W/ZdJLTbG4KV9LxIm3fFXqzcMl9TV9w+yXmAd6YBOoBPvNGC6+les3qO
ohrFizRN0qGUasFp/6j7B+wS+wWMd/VJxSDvc7tB3QZYC3bs6cvjBu0Z/vvlf/Cl
xgQxojr08Hi8essJFEmEQg6/vpVxVdeUaIAAVkuFtwvTaLpwNg0BO1qc2nrhZJMN
GVUEexTPKgtt91rbOahFTjdwCy03spzbl4vIpBi61kdaNQjvHi6r57uzgkQJyBKG
xdH9C4qyY6NqNubZGoxf1EQmNopHgOVu948ZK9hei8yq3EYv5TKSIP4QV3mYXaHy
m86dse+fpaDwuLQgr7D9ggo0nfrV6vfxrqBwjcrXElyKUQhCjNmfirCDqW/iaHg5
YOiJOOy5U4UFbLo5zLnOKgrzLFAGCr4yfoLGxskbpjE9jkBRKLTFzy8gwmXGqwUY
ODJlazc/bsgIqx9LN3Qr5Aw6bC91XziX3/QfI7Sx2pSfMHE5PKe+7Wk9aWhfRr1W
h/+fVwa7tVEMz2oboSw+EkvuWLDH/clRdouzJEbQfIcCtpHDbAjb1VyctFHXiEDj
Ti+IMatcqwBSFtWlmWRaKq9r+DQNePDviVG2pQ8kZM6C5utY9yabFd8rKgtIoK+G
uhXnZrQjVn0QdtuMtr0MRNGgPM3hHxunWA5Gs7xAozV+64ghS5eezXFepnwWehhO
Wi4JMkls9+/tx7XHFsCmxpVwIS8IVbAMfAFzp5UZlNH9K2i3R6STw9ZH5P/uUZSO
HYw3x5/hhqlMG51zBJPt/6IK2GHN87u9XtEhfpjllUdHOrbyD3+iczHKZ2f+DwML
XCGTFBU5I2DR0vg1bEcTncXsokIRnxkCb9Kr6KWyrBBsknc3brQV7jGBoCZbKtio
Ittxgn7CAS6OvvINl7AmfF+nyVgxc5IvkiHylUeHqIEV6CCfSAZaYB42cyRpsLVC
plExx+aUkFDxahlQOzuLyCUKzmtZbxVDZlSfKCjRKdk1Q2gi9e79TnyFdITS38u5
b4RjbsBuDYfmZKtbUCyCzkgBeOQ9JiZFE+lGhza+mAaVZzTWVFZynFlwPkhByzTF
s1efUuo/DLsXZj6Ar0Eiv09W6YmvzWQfNIbKbFLkdXzB3BQWd4oQvaZU27OR1Lji
a9jigqFeNplADk7ZuZIB5A==
`protect END_PROTECTED
