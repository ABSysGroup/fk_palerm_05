`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TYFq03RzyoP9SuxngG5N8eDSLralnOOpkGcX1vuA7Q2LIvFiPcs4G1ENAVcdskqK
1dxdGkfMBck5+SJmVOYmNmg0IGOK0Swe7yMd/FHTVkxNqn5Kp/Q6ed+gnbGlmm8f
X/y2X2snzEqPJcdeYMbFHTT3fE4F6D1O9GnEC5LnkMOayULRYAa4IigcH4VsfniB
jAN/fhETBftMMaRJuqjlLISs8UE6tEvZTCgn0PTcPRH0pZmLr7E8s6AX0YVc2P+J
+Ob9UbKEiSJTxaOrNy1DUJwkRxprbJ6bUSvum77gmVdsUMM0I4hmztv5PNB0QRVB
VPq7QWuSp9JxEVslNvRBGxkGV90l/JTVxEy+EuwlYLkAg/5U+1ZFuyQIRDBlF9h1
B2y1H7DG2AHQLnEAdNmdR0csBbujoNhb4e5Sa2+QrHM1/ja/ttPZMdX0+TOMURC2
7NvAgsIarGgXtFmUHBMBpn1euJnLUGCKyNSj+5LdMcg97STrIMg48OGg+9bp9zDz
I4KXwyYYx5wniJ643wnrbiUHCZPUPMZXFqCI18fuWEacJRw+1RzXEJPScyNvbm7W
5lK2lxNurzpZRU/GkOolH42xkJo+A6RmTpv6keGKuI7TTVkyJOXDowMMHGyvzyBo
5XZr0KqUxmWrZZxgNlb8IaglNmtjBEa27AmecfgBRMdGyUDBTnX/tJKD6xgtfrwf
mnWsRCedafV6mlXBZ5JwrA0bSImfHIS/ZYRuH8406qQClDx6pM7Btl/JlFNygh3a
44cCem5JmgdRtATuqpCjSk44f0klTtnhEhMKp9qS+T/9jBVcWT/37YfW5iQeserW
I5oW7NSBdVGRvm6omPRGKF7lSX1isXlQHDyyS+ktvPbYU6ey9h2wUgQBXtnSfq4h
XRuxQe8z3kTTWKkjdjC/XMIvDy/9zjrURpwXp32jbn7VisqZRDtQb4+LrOnJBqeV
JOB19gmDj9NL3BFxUOAMZ1vANicHjPZeeBwd2U8umxU73FntpcjxXmy2+IzMtzsa
YQgZiksMNHZ5DV54Ccn0IBWAC8viby0xg54ogxJ9ZQlGIxTKfQdI2LUNTn8Sxx+T
VOYQ2psgIfxDulB1sojxt9oRqYETNcbbPnoPy0EXM1HuiQOQue+1Lh8xz81HXTpX
WS6ToXMNlbhwGvJwP1OX8IxB9tKPX74Q+uU50PinbNn+3LleoPTAQ/RgI/o6bzVP
v3b+Mcvv7/GyEPcZ9IcdBFEQI5cS+VNNKQMtwQeEgqOoF1TBWnE9MBCEuEsgEnNH
fry2gdvAjx5xSWH4UkXFZl2mXU/QxI65G32oJaWMXQ//8awbvY8CF0guPlv33PDQ
VZzZAly/zDFcratixqYPFUNpyyY121Z5lzHlcJ0vmaxLiNRluAd7tVWD4Igl9PA/
a1RMuEzM6a+FNW/zVBLGoNQnAnYfdOuw10FEIXvQvzVMLTSv3WD8kZPSh47FCkJM
KnOcjbRDXgSeArt31C7pPm6ZxO6TX2VExVBVRt0hCV9rxWoX9dE0CpXjKDlYqGpI
SD0OfMDihZtBoE6NqY/gMHlsLN8Vh25TH5zbOT4b9N23IBYEdPZM0unyq3tFlasv
mfN2h0uMZULPPRlwd4hUxNfdzYKrnT4xkgK9re1MYVPODUoSc5tzT88YQc0eP/f4
u2p7/MEH/zz2d90fqBaHoyGq9urEKy52bO28bzaRl87arZT+jMuoYxrmqxcofHyS
1yTc9XY3YiN8+LGpdV2kUDar5Gkd0XyQGnYFlzdD2mcwUMFRVZ1hDcuD/PR1EM6R
VYnGW/Tix9myqlPxQX7+iHKcbMIMPSygBp41vL5cVe8gSlI2QowNX+1YsuXh9VA8
EhGSkhnM8TbiJVuzgu+uq3G0rd4hDRMN3G7LsBvzKXfpbwlH1063hQlPGzMeOpVb
Wpt7I6nNSAo0Rr78LE3+6BQmSqM4Gqn3qL+sApef9fhvxkhxFZY6AfeC20vbVJkF
j5HwUTznY4sLRVgZueES+topsTNO/3vrkK+l1Keai/rzNsDsgDt0Mnk2MzP1mIAC
Su514vw/L7mC09KQJ2vQ6X9qGX+ePyfJ1G7JUJ1VdZlHL0jg0SKDrzCxEko1CDyT
LmyDafBxd5BPDF/aLYLT2cNbnf9DpWnYdz+IYjUTgIJBAWJrLyiVkA2ioCsSzU6U
bQIK1Y0kBrDd4oJKc0fYHPsihDJ1lmFT/cnfR6xiOwNeawJMW5gZdoL6NKKVwB1W
yZytGDKH6LRCZKirRHWjFj4iOO/AzHeH/+Pa2dDNiN7qwsSNL1yL59ns47BpT0L3
7Ypa4wHWeaRDFe6Yi2wfuNwwqIugA6vfWLFbWufjR0kZV/IyyrPX7j+TKjEXOyee
e2ytvtX/TCY+CXg66MCLxIb3w/5ZLjlSSykgARNzFSecE3vmjQKkuyKgJ7QG4MJt
AF2NPSDwuFY5Ax0rI1Fqi5BInxVpoLcf514oQvWv1Uy+Wo25vR3oroKAAdSiUc7m
GQ6S9dajD9lLg8vhAmvjsMdLY7WHorT6Hm2d+XYtJA8n/w4pKq8g/YV6ZRMFSn2Q
aWzDmi1m4JFPTOS8elZuC7p3TO4Oug9OQaPOk6jzUFU9Jp5ue0AeTOWpsj/OO0GN
`protect END_PROTECTED
