`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hbMuu3UU9Tt8YuemcxBD4j924czEznAJ/EENqzkAx5zz+m7upLhr1K5rYfqSDhZh
x3GeiR5K2TQWLJ9BgWhqhiiSr3w2mQeaax9V9gSq59wUroO41jo+X7DbmbA/SYT1
TlbWUKG+Up1fy95gHIX/lFtkW0si6lvQL4bqvq78bvjrao5soEWM2ncsheJjmwNq
+N3jLQwXYoM3cM3Ut9oEqCPZJ3thCDCRP3rpR5qpeWsjoeMNC3AwyCzmptEEp66J
k14iJYwFEw0Rfc+EN8hItmL+ZOAeIkro9s2nw+pihnjbdjm5/GNNe2GjCPtNDC9l
ZFdZN0AX1vDZONv0D+xHo76eJCrLMFzw52TSpnroFNtMD7GeVsnTcDXWF1KWoBzr
x7k/Yjhq1kRKa8TjnZxE+5+9d7ASstp9rpUA25d9fqXjJ4E9UTQYIbUUE4xym52r
4DyNNSKA/xBoA+zgqAiAkw==
`protect END_PROTECTED
