`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aLjGuoyTjt7CdAMJda0tvtshbrmYCqNQuUNPJeKgQQESvmxXS9EcOY/8srfs8lgf
kreZrIryfh1nUk2JttMTEY/8ICfPM2/uqLGiPiOKPS2OpxtKQ/HbeH26FGHvxUge
QpRm7Pl/xwkaI1LNOUQNy80WUuFjQP8H7krxp0fVTVpxxZaus3xPa7gGSjYE4jw4
xGAQTXK/8y2Soo7HysvboOcRbeAvBc+oRSGHDmLLEYKYTHdnseq4fcDZlHTmaUIZ
HwbtdSfctME7X0ozevdIFA==
`protect END_PROTECTED
