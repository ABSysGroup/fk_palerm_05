`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o7y8Ll/W95WZTM+2EVLg7Xin32Lc97+zEGmXQHliVsrcLG8QRBrlp0fd01qFb3Bc
pRTXTY2QGZc3jNe4kQKhQPmEqQSt74RBv+stxAzqVxmjEdTQUSAFCnxA7v67Pnc+
MNtBY7jEZuaIugDeVmAtfIa86kZA3FlHhmWlI8SxdGtEMKRPbtXgL/0jqZh9Q2Yc
C1feMXr7tJjjWQYJdz7pHQM6PzTot10nNgjWlnlCfGEy9nC9ppqjaHWAhK9QV+Li
2CYdumT1wFldxevD8q3lg5bTP3F/i0grCE1rW4DuIxQZIyPwbBUsCreJbLYgGMem
rfEFBPuFnDfqKOZDelllvZd1MEM0hAOiubJOWGqGEq9VwDGIi3xjPPEPWsAMWCOp
GPV+gyGYBzfB4GRfj7H45ugNL2QHIMOJlc2l6j3dCTeYFkGIpnzou6r24gzi0cM4
nwAUsHXIQnyBu1GUBFEuxOHFM84nguW7Q+pb0uiy45HLytkfLzpJmJ/67rd6RtFY
fyLkOfj5pbQ8dgdPHwW4sjfDFSYYou3dxqpYUEt/9Ks=
`protect END_PROTECTED
