`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MEiBziwYb3nnkBCNWPtb8GDB+ClnpvkGzRqZxe1fetfF6zmGG8f21Ii1e3sHHvGb
ZOQSJV2M+cItLxWtTHEwhNHIgSV5+oJcP/qIjEfqa7UM8tcZziBiq0z7b4e3u+UR
S2Xi009Ze7KeurtFz1kDvMcuusQF8IYkTk6r+sEjns7DIOUYFSmcwItm7DoJ2Q7q
K1nmSvXHeep1QJ7aIMPr+c4k1AHnnxCMSnygFHo/3PoznI1JQ2jBzjLj6t2B2O/4
UQeJ6xLJQlGNhgNgD/dXb52b7DZIPQkfdSn8fzjV+g2fbljaDaKCS5OBpBLdwCgn
rEh6Kt7NF+4Fda7fyk51wdqPYKBa3jcbW6FOr5XkZqeoXAgr0ptgY31RGSwo5gcY
+JBU7Px6IG7aXR0ESgEYpSqscM1i9dZvg0tJPZvzrmi16tmJLyGZxbjyBGb/io3q
a2z4qoUR2x4rDN8oE7OUua3SW5xnH7jEc1tdfqvQi8YODjJOW4LGr96K0lgTI2Ki
fnpfQI9Pr+/CkNp2Zzc6ot+Z3hKJcZyjzuRQtedw9oJoV9DEWTbRFVZFHy2Ub1W6
V1FyFc1Wo6E1EIfPzXBgYs0pwo2xI+HD2MHEydWWC1oUej8F6H3BT3j49UdrtIH/
QWhXyN8XH7L6yeLUUxxfZ06mjhLd6V/ZInBdlK2KXcI4SN13t6rhJTiXETfaBDPy
TMj31edK23PwrWQ4ZZdf0eGdmgikxcvj0GQydapJU1m+PvMCsxgUxmEqwBPm1Q+k
cmYExphPE6d2fG8M71vD9W/p1yULGZ+v61RbjCWqa9s=
`protect END_PROTECTED
