`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C0w9QmxI+zw7WkplnvFZqaNLE0Jt0Ly7GAYNvQ9AIz830uK1CeFYe2ow6BrpzyjV
6bNj3zjW3GZugizSQt1tjFtiS6V//Fuz+BYcg4O/qPJ33gvopslPugxzcsQzcVEF
bh8jBAP/pinukQpAK0JwmYA4Nl+jS8o8ag5gt8ccNRyJSMdgTgMNJvuIuDtCDlMM
ozHCLQNlbpg0FgyGmD5GCepgInJVJMn8YQpvr9PpHsU2osyKVc8nX74gt1RqcLmf
ingIwNUW3/l9IesOBZ1brbH1ApNo0UxtigZfqQSVleII42ds+77zN5VZt1VGJled
/hxh0NfqL5DPlccT87GZtTB2UF8axU3ochJa+VegElhkMO5JKGG4XGbUZtLOg0wS
JIv1gDF/YtZK0ZRPwD4AZ+i66BN42IaxlECxbnEcrrnDu0R+6CZG5GqLYj0pimeU
vLNcLXcvuEbkZtph72yoqQ==
`protect END_PROTECTED
