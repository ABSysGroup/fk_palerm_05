`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZTbkl2m9JPm6xDcMHy1h7+yMaDEduF3vL6Onh2qz41Dp6sGf+s3H3uusH2LsHONB
aF+Gl44P7VMXbe+THWL+aApy7TrJCiRrzrflVLOLWRg0rctTLb6v7hnQ4RaUKFn3
Gs4bTA9fuXEeDDOMqXma61loVKXcFuRO4YM+E3+qlk0mHdF0YQN8mxIVcSbb/4ps
JR2wYP6cKAa+n2Xsv2VTdYtsW8Nik4HIDOqI/IvZmv1uUuNOkb+SecIu9JoYDNhI
45hhgNqyaQmGHpnSvjkbm27M7VnH+KQ3kmOE7tWP/faYevgggNc6pJ0nhN4HjxvM
Z5W35D5OrwBS7OuZGlf6CENHcSVGLr20TbdScbe7Q8SOS89o3dNPoMiJUkw12fgp
Wx3zG2g0QY7IzFydOfN1rf6acqNELZ4cPOexJBOHpvd1N3NwOlRsVO7hnLlk1PhI
CN5zc4v63/Ag2E+wCvcGkfmhV9VrbVHWhC3qCPITW0E=
`protect END_PROTECTED
