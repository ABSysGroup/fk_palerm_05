`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MYZws+LuyQActhTkLDYoH+CWL1D4qwNflVFh5pDRp0uiYisg3jc5/mWm4gr0flfw
3BlkiYh8GARYpK0eWUpJ0M8qtA6324IA1kpELu7VqpZBHthzui6l/hcHWGzZsy1O
kRsRO/wPHtZYUeHsVRwqd+VNfq0bbn5SmJc8zX0QX+obC65m1zgQeEECS8ylRfLJ
chST/hDR5mrFTIzHt2PkL3yDr1BhDVf5xAfDPCb8s7XgHfTXmk/pqFyIDnRzhEKm
Lq4YzCI2KVkFd5OOkGB0tnzaEQb81tk452EJ5kn6GGsYQtCUNw8Gs5hln1WJ7tle
oH/9sN8s8TrhG2MvwxmaOD86KXt1atQmppY7hBcmuXOSlIlbYDnebwhUwNiTtjpT
LlHem/d6GMixhLhmFKhrMpGMqbfUTshiw6OcBm74oEGgyDbQhJcWJP0EM22r8Ifi
zSK91+XLagc5cstFsDuIEKERg+F7lJNAlBnT+8sqLSu/Ryx1qRmToySJT7kheBzU
k6YivSo3rbmekaSV/WjElkPzSrPDGONFbjr6MevDNSzQMGV+ESQHKR0UUU8DLIHy
PIO7RlIhPRjdvtaNms5Gvy1ukIuHhAAYne7oKRRd6E1de1jo5wTAX9xJZEmtBBKj
imy9d5GPPEn06hpmFpjZpcozgWBB1L+YBA7KsjVr6xcDiBywQNozOEO0+1ER7Hv8
NhLmasSSYaAApVr7bfRKPsttsLoTc7cJwNpVwDNBXwkXQ4FjGn+cSONbUbPOv4rG
rBO9UY22He2sTYpKBcZU6Q==
`protect END_PROTECTED
