`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jy4XTQTiU2is6qokD8lsf6I+A4xOFXA5XRCMA8ubDpJBMEhDSYfc+NsxuKmhFleR
Ij42+cR3CgDR+W34HPvsC2v/EmimaivgHloVAaZCTmYeuYcmHsLZS1meGfIqvDGR
xPXJWi1hDzo9qjcjpFVWfgqym5U0N8mCwB4T0mOk38HpD5ragoi5ENkXtI7PR2E3
QdR3RjZH3NpJKkGEreSd9lsgK92r/AH2stqGiF+YdPHv/3XVV+z6Mecuw5RdkL5x
UWFS/8Fgq9YQxAq5ELsn4ChdfCfV9cscT1d/YWL4/5NGRU9T4FRRyxyfWnLelU6C
ZAfa0BU4bwOdkmxQTw6aYNofYMY93dvaQArTBN9STwlXLuZiZSuPh30mT8alEuxd
48M4A1PAprljn+tJ3Zo1jOpnnApL929gIj+tFnzDziqWlConNGqrOleH+aUZq026
4U9rdYscNWCdykfB69b12v+zlriWeysXU7Wg+MTqGn0FrOhPb5keaKCnCHLpIltw
oDUzOWq2zj8X2NAN+uPr+oXpFA7E9U8cj68v0gKojI/3fDYN+BLKiN0PCXloWEKI
lA3m6zVIE1bpACVxfjl5daxwyqacS2Itb0qYdgKSGGlHU+tDEYRfzCbO8Om9XITY
nHeuBlUnYOy0Ynxb9Wl0J1/ShfevXrBcXvcSI+oVfKWl9ZKZxjzH4QFec3eLRJNs
r51Dy6z40yvn2FCnsA+FvLXWj4yfGPPU/BHdparubde2NoAAb9WlcCffL6HsqUZK
IRZIRK6vGNRwhHRdMET7xAX7ogNX5blSFCh53rBEi+OMPREZAz3znHM9QFSG487N
9urgpAXnmLYRlIY2S9jruZ7v/8Soord/BTw5GNYOQmc8AisTgOdpo2NBW0K/mTck
G4hrAoKAV1PwnnDrENsPQsYldqdW5VAVD8GoWIPL8qM=
`protect END_PROTECTED
