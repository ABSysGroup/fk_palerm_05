`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3U+BT9YXmRtb7wM9P2+7r1IOvc94S4SBE57/JJt0tMJiMKkSZoWnqRd+fVOQwpGc
6fZixhlpaTk5mWUWuUJyQb0ybE7OEa9sgA91gBIOYfAN7dpFy1HBENlDPgP0za9a
0N/ikGuQqTwaZu6broOT6qRYeR54YNMLLRfq2Rwq6wCVQwi/pPpviTmgzyOihizT
/Ye1EaOJx5/cFJXbU/cN8DXExYrUd0/i91WerzsedcW8GoErrueiMq8HmgKZeFAJ
IgOUOE2bHjwCtWRlfwuGqMhZVaIjzxiZDNEON4wqH8FE0GnXH0BykCk6gB6cPa8R
`protect END_PROTECTED
