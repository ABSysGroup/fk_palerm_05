`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q00tPhBlzrhcKX8GxaWXKN1XiQEaDM51pPYxJJ7TRz4XT/3lc1doADAUG6UFhll1
lnspywFj+yO+ZgQ86ZydH1jIpf2G/BVDxLxp5H/ZuStzfVwIsgUfJmOGjqGZnhNY
Wt7e66bYi7vPlCzEukwWMLSaa9Zymp/KjepsBlCjs6NUtVIjdd4Up3aX+Vu+3ZyQ
gMZNAiZKzC3P0HaL6SUDweioxzOfHRVxE+Pn6SHMmWoBt8cac9JaAjtyP2eNkZd+
gEYRlKwNe5MlcdDWHt9xqOxojEk1lFO9iH7s1eddAz2XjoSsIoZ1XdTJGK8jgQhH
oJNN1LkN3r5QqkJ8J85BwvmXTbFuF2q3T9mmeBLhZVrGyYaec5MxoJxwkt2RiO+q
5IUaS1TM1ck5AZntfH06sYH/dL2KkRpBfEeMZnLsG2SJ1U8SunrzaDANDuIzee1q
edjEUc7iDPpEM3FK4JnXidoAppqypCCHcVkx2cCaPqQ=
`protect END_PROTECTED
