`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tsKqRD+l453XsKExXghCz1pIKrcV+qsbv3Z9Ik3OrWBupR+qxVnLap1hGCUkxgoU
fwVxlbxG/+0uXE4LrJthQx8dlBTxvECjWhjeOoWbcsm9xuAE85TWY6Gn+4VraKa4
chyyEtCj4sihoCxoqLVj1RXDrhQyz9qCpyZDk4OZKYD8oAcUZbpoNa+SiojR+x2+
n9d+66zHknqcJYEWd4uJVRyImTA1jvI71na7LUTlQO67A2xXlyN4l/eqJiYLF/MF
sXDRTd5dIf3X/Jax0EEG68Kfc7rYY+PnbGxlBnj/S0g=
`protect END_PROTECTED
