`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RCHY+rDyJhFZI1dCV9xtvdtSBcqO+U6AnyUpRVoyCtuk1wQd5oMBE42FSynKsNbr
oQTE3LTtetyMUG4k3TL44J49pmQ48msUQKvVfwi3n50ilcUFAdkDZaGKvGYmIWdl
cDP6rCVDlz27Ud+ljuYMyGpfJ+nXjBqZ7w1Bnes8q1KGdKqkcHMsY/eVXlW2Tke8
vFvN2VvaHYAvKtMX7FRYDCQU4zm0RCbU1abzS3P9QRLWExAPVBE7iPI1xhHwNKCc
8YANVLzK93douAJ95VrMnPEx0OITDOwMUUzrL1twn9un2myKvYbwNw+XGimAyruE
wsm7MkF48gRe6F0QLjgZLP6crS9iPAxfEXghELbeRVNiQD+QtqJIfrtEdK69U81R
56YbAR/OWJkWsIM3lg1gF017lT5eOm/TYPudEaN6VA5G1gMCbjOyLTsmMpl29qzw
kIs6Od4RoVfNBjSK46HQdbdAygRLUlYmgT7ZYBEUa0HpsUBYCpBzXdTh1u8mdjK6
WsG+tmzq4XkOn0b3yOWnkzmN8RQ9CFugJUeFhqPMF8Mz9gZNbompqVmVC5qp53qv
91Disv/AWD/bJkhXMWvKA/4BwTe8RbPHGFnxGHTjAyRFYQLt+08RkjohxJD2t4gs
bj12lbTGIVEmn1aidq/9e+XJ4Wt0KA1sJfZ+QjaDZxu5yWzLfQa76NVFsUJkwMtV
VkQh/yrDpjGj0osjRwFHZoiygvlbFhouYhpd8et1pjDpIW9X7MJ8E2JshrmN8itU
WVhL4UJ7XZfxv13UpRSI2w==
`protect END_PROTECTED
