`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2oolXry+MDOYdDgql/CBMSEHgLxYIoUC4ngOp7CuAPjE57pqdoFBofY8P8U/Wj+0
oModfLTQSvMAZj0qZ4RTqkOy7utu/K5yzGiB9f7nkSacdG/tfSC3GwATvsGsrhmW
ipaBVczSBFY7ZW+c4XSSdIE13LB5HIUVRczAUnGDeUGTLaCZj/91sgAGzASuoRu6
U4IFjM9tJavKckg1AfISGTbN43OkbrFhcaGoxTOfAJ8IFi3VaPk5I/058oLZ+/WW
kH9ZOahd706O5Bd2vaLe79DJA3TQkjqKfJkr105YZPQt7ntfHTcSMndJwUdafg9s
NF0ztZPUpofemYYmz7DJkyOJMk2TaI/fnprZJMo97QIYjMmlXuFD3Yl2yXzKoM/e
d1jKNHUCWN+poRkRVRWPL9rzEzFAwLc/hk117KcjggEiAThCahXHwap1LIzcZCes
CuOxI7ySNm0J26QPYlAUXlBFyFXbcrNTcbsny3N3wn33ccsCRl0WzOikug6q2YG4
twF465ARpDg7Y11YlgBOhSkIJvW9eg7SKW7uFh+0/sbKITqrdOmWCqPQUi0KFYD4
//dJn5DVgMxGVgOWVbyav6/zsCOTKhzHkZ+r+cxOjFW0BNR3PqNSzIPQEs9wHE6z
R6upVKcahs03F1YASpDGGs7AAMdsARVEuvX33Vz1/Tj19qCeadOGBqjaYANL+eh1
3Aq0q1VtQiHp2y7X66WMCfrbsrfxA8qXYdaBzBnXQ7ZeWUycRPU1Bj6Cww7/yqIk
4mKjFotCqvFzm7MNQlhGqaeCZQya/WyvJykDTyqSFYCWJZ6fOQrZglbEH3AnDrTB
iB1Hb+8VwatoWWyVYddIZvFWjZYwWVF74dks0dKjXsIrVsH4Va3Sj5W96K2vcDTT
NNHjFjzyISaK3B/wqaPh85Mv0lmyqxdXDqnqE/q7zWpGkdovlW5ud9AZoyowWPYG
`protect END_PROTECTED
