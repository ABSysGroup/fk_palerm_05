`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pSHlK/nZrMG9aq+O39MOWofph1qsNZUjHRxSVoWnIivUEAV39VhtkCUjnLgSgOBv
aZQZsPbr20nqrd+o+O/4qoHMDZRPUjUcSE8XgoOAGZNWxv629rwOwvsi5+DrzrTb
tfUOmD36VOdcrcVsXgoCAXLmvAPZTk2HWNi8hWfdQFqOGsr3H7l8sVDKxVfIyLDI
5zy0fvvY0+fIjGMYidqs8BK9A9kZf5nnBTHF8sBIYswZwOpHYJn5DBCC2aHEJcjB
IcvswMBGZBWwYi3SktAbKc9ouAKI6fM5+Idqammbqs+In3lRDcJ8C+BL//+9r0OY
+B3llp8u7EBDS0VjYdwTfjZ9MOGSjQCVZf/p/2egxy3pCJJExfbZZxdB2aeHDnx8
tN43HICmsr10JHvHgktv9vzPFJQipVigC6aIn2aU8rzKxBYpPo33a67H9+YlyyNA
AoQzbtmTxI7rADkjFSe4+MbZKz4k/dKIM4yGmXMQW9hD59ROUJwb60eUJAa9ng5Z
Z/vzKuvcO8TeL1g5Gp9CPFrU6sH1+ch3VttnPQ2NkxR2OqnuW0KvC92dHaBe5ced
9vvpc3Cq8+mzwlhGJ9QNGArwfD1OXKOR39Em4gXXtDRlLqIdYnqH/wrO3SZGRIxL
3JYGdIYaxnkbedqMMwcg0Qh1W1rF/vz9kBIaUE1BLcBrnrI1f/h5vZP2O0rdKI+e
+fdrjmtWE0d+R9FwTpxKP+rVIgbveH9f2eijnPYGcDz7i1C7RgOY+uTrB+29I1S2
pPOy4Jc3BOqe3YxqGpSyZzIFGATY6UZlU3cbwbnzo6WMdcp0V7HYJFQkH7+qp+LQ
Axz45z24aKFoCDO757663iUDKRSebcKJDrpoF2yv4EltFHuKKa54y5fQJCqPwR80
2z5pUGsMzpntX99hgXI1eyMGu5RUFCfJ9W5+49uvTVK49XVYJRFKNltwY1jKiQkP
pqNHXXxmmqWVZ6eT8osxQ56rWE/FopY7XOVroHXgNuyG0u6dWMt4tMR/rMQWh2iy
91FrJiHEWiK8Xn25MBVzOw==
`protect END_PROTECTED
