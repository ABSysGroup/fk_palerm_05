`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wK++zE2B0RT9fQf4gqUjUwUD5VUZNbrqibDU8eqgFyeBVJa5mwXS8elIILTTtL8Y
a0+7eG6IH5fiSVGxtX9HAdpzqgr7YaDbEBtKbpSKcpFNioIkNQCMgwA94PcKNK7T
h8OcHWgFbOI0JMjKH7eEcrxjOWXJxsAVbw5Mr6iqS+8PfqeKSSBvwoLPu+NoRljA
D3nfQ/4fcuCuvZabuydYkJs4rF2bUahqurBf5ksmyzPNJvKlOXLpFPSahsxSK0aD
CGTdzS37e3AnCx94XfQiQs/dOBj/VsvMFi/2ZPwYJCP6iknDgH/UkQ8LcBik7ULO
/lRNu4L9yB0jTX3V51hxPA==
`protect END_PROTECTED
