`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HIuzOWU9LqZ/QXDw3iJu/Vg3IrVV/XRcDZJwZjeIKhBz7wS3dx+IDy+iDCI3zIvy
sMz0IqzdSTPtuXqnLHr7j8zy4LKoCYmxOaevRIeBYtMjoN4aAbljaEMqgiyxSiMb
CPSX1LuYjxNLO1yIH0gQwhhummos43QAZP+VyJz/IHWD4Zyg4VbbtuKZxgWQpXku
u4Xrz95iBlm9BQfoxHPqJJE74wqO+tpRjOgSIjpEKndkelvnH9BttAtv++2iRWb2
x5NxwMBpdVITlu0k4waKBohEMSZPs1VKEOBksk6st15igiiFGL7Magu3NnT7kZHR
2jfQA+T8mCOL5fl24UIBZiIiEEJ70Uccj6Boul0lnaZfbOSEx8tO9embLe5nrLT1
1wCgEGUNf/NtMxXmDMYVzN2FZRkEkiaEnJhjsA1cMHrsUiQXotMSVtDe2X1mNUOP
pPGXDvFLAWFO8fWEQtDocZ1m6DBsKe5oS3QPcSKUXZphiv4xfmpV4k4zf0pTl/dX
bddDkCU4KVe0rfeTSAlVf2L8GH4YeDNog+bCeD19WvM=
`protect END_PROTECTED
