`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Who+zxf/aOx6vpsqH/pGG4y2cvLwAVYun4BXmqcjk2SkRKJqx0vgmiIJsXdKJiIi
gE7h9pwf0WkK9JM3RxTp+y8jpdW1k54rwQ4rkPwqthUYRayzHeXjGXMkpT4xfgAJ
5izR0fTFcq2YUvJ87QehwUcHuwKWu1EBcv3q12s/sVNvBIZZavpJJWedNoAs6h6Q
pW65euj4C3aWxX5ms83e+aWovgkFhHIyIALylum9rH7aY67IMzFrbj50MXhY1li3
N06pTqbEWvgMuITb6UdLj1t9lpv0WIcXdiHL0OG7mm3NMLP9SA6r8+otRGybQ+di
esNevG1INJnNosnx/zrcrg==
`protect END_PROTECTED
