`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EkYTpXComRvfp0bpZhfagBIIR9Lw4VLDu7sqOzdByq4y4BhwB5hzNyLTPAKqYiTl
lQXLQ5mKjSSi6uv7BJ7yZkqI4f0LuvcAVJyd44F7gONakJoajI0iy+Wsdk6CKEY/
R8ogN6dpCth91YVwZZzEyXnTXYnE50cAcYMqmoaNa1F/LzVqOy5ZZljHbcVmpFN/
uX8r9fpn2iKQjvEDSSsI4ktfR/lKyZZ/LWWPHYPwgRjhq6q/8qNBGwT1xubxo1Li
DKF5zZt/yeiPLAaZYFlSyhORjsThZGpGaADMQtVUlamd1eVlwpFBaJC9VbsdcXyp
`protect END_PROTECTED
