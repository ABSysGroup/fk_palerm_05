`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oSD6noIcNmAkz9cDTCDH4XU0Bf4vrx9uQi6NCw5lD0Jg7DgLKYm5x04JpmDcPLfp
52sJ7Yjl9DnL9VeeMvqkNzCI8jzP2OCfi0eqSIlLN2L/YhQt16WLqLUwbsOulRTo
l5fuqtSKCjW5pD5XCmOwf+o0rRW7tn0unkvPT+QSzJskNc9ACCT9s27WcYYFGM0+
NZloWghFa8Jo20czA91xR4PgNyV/wYbRV4iwYI+2C5ayluNeiuCUoUd6Ktyaaa2t
oR3viluuG2EfXQEZZGSD00hiL9vgMxg7O9TKqbeDoIdZZ8gW2VcvrgBFfM+o5r0q
VNtd0h1C/su9Prt9N97uz9SchsrVXR4U3UoZcVSQalU4gEdFy0YE+GAvta8MlAit
ONru3uLlgn9hvqEBhqy5GBAzVO2GUe/8puLRuFHDbdX0A3iM7zJlBjitWhwQxWob
0aVYaX9uAKJu4cy+wJqWhIDSyu5BWQnX3tnlQodvHxU0013PjuMiiHhjahUrvLlO
XI5aSRy2vJo8ggBQOm0muqBbcB6P6HTPhRb/lFQ4IpHsPunEYKjat/kYRvRjdFQE
EbEQtpsauymcHDuoiq4Xci62MSr5zBXYoLp+DvkYuYbs2+MjLyZhZb789fV15fNT
zQDM9sVD7CoNqCQto+rtktH4XeLkQy+DdGZiE56C7RiYLCET4k0hpEq6Vt6KS/FX
kRJ/B+3+CDZSoK75nLHz/P085EW6Hyctm2AxzSMMXvkU5f/bY3svBGCCWIw2JVMz
4BkV1S61bWmPiqdUSdztExNzIf5mVyGKVoxPN+D/xE7jMnb9eSWm820PKuxwLlEu
IDUC6/wqCyTo1F/mvDBvGzD0XCP4+98QnQYkW/2NqNYgxzZWfGVGVrOP9oxa1IeQ
isI/57muMKPO9HpBy9W6D9T/LyjDolxrlWNco8NtgTHNl61SoaVV8QonSVQsZKqr
ctQBj9v5ZpSTJg6dsaB7halryHWSjDlYsP3OEMqWJNXYeWB5pjNOIOCaLtzAwyQN
gPgjW+lX7goTSv8ZUl5/FrC8aTKdrFHcgcdv1+b98kwyU+VBcDMvHuk8nEpBmNgl
v/jcXfVz/zfkATLnn6mp1SthgKbV8KYUH2zqGGiytpNa8A2lIveRf7UXDPMfE5JV
YJ2zV37Rh3OcjLFkI7JoLUXIn+bPcBmcTj0S/XHAPVizzdZXCSRESk79fpPavwP7
+K1B6+vxnua6kTNzIgj/uImCttY2WQ3/yU0I4ghTR206LOvoAF7jxQ/YosQCcO+i
mib5o2ydPmkdmgFqgO5VJ8I3IFG6SbDnfN2ztgMOags86CKK58WanmOYGhJXKjRd
6THSTQd67YGlTv4NEShk/gKHKvy1w+7JNxD9YDbk4BqmB4FQhiMqPgesPouQZzV0
snXLILFRXJGIpsjeTq0Sxet/6Jb0b6SscLl8YxYgsEt+cBxsXayQpV3agDBzGNzU
fE+VvpUmHRXnzYyWpP62TkaqTQydIOQx8wpSmvLO5XQBa2avjIQ0UEIkmnzuXlWp
lBnijheYp/vyX7KvqG36AJjvZvMxq7h4FZmL+PorOx+CFpYty+WUQMvwD1lq6esO
ulNtcV+ZHIvyxkiZvI92ubIpndtCW0Uf7HCaGQGJEiP03x48zBwiKkLGReqLJ7qD
jIoFnqrpHqUEfdu3mZ0uFFQWDLe6Apd7J5NL+bfO7t3r9Cl7VYp5g3TFAdXwi8K4
JpC34GJrLVI6IVPb4eSmOlwuwHh0xeWlrwI65TK/0eoybMssFyxMF9hqVp3ktYX7
V4FsPZ21pAWBcAe9VBoyxmabWsqt/zJhLPRbnIYbLvvrBEvtuLzAF+UlXsv+tqOQ
qyA5QS9hAaoQ9X5Q9SU+Y+P0E5mPJCjpvNKKqg8kMucSRxPKID7tE8H3vwEuyVpP
okcCzhlnNS9nS7aKkYtRl9XznW8vGW9upz99iAgZd729O0qNxRlJE/pW4rDCGCg7
frI8i5UPbWklbOZwQcy9TuX2HwVLtdVdhao6XW6SYXpjtOCkkDD6G/ij+JQOCSTN
H9UFBZnymN4PR1Lgb01LzoLwz545bk+ao6WHTpzhd4qvQH0jzl8kmF/x1/TGJ50G
qPTqWYOH9HxaX0qRSzyCQsE/bwoDnpQjy1TwUq8/ZDkDNU52CQhu8yz3s/u3DkS8
8ZlAi/EFbb/CFaAq2AVHXe4Q61TJq3x71LDQNMpVqsmAE+rlCfA9chxV7FtBTsyB
BIe3dt/XNs1xbXfxU0MXssQYoAyQ6gD1e+ga8IL1AWUqdHbxNHJcbaIYbzhaQZTa
0nteGHLQcZAJYmoDKLk99TuGG1nW5qJ2dRZq3nfATbvP9BDmoKlTKfK9CkUoRcD6
Jo1ZxLwotigvjRfJr66epV5DSzjVPGp1xE2BipaLVlVpuLLOTQ+ADCkO5AcS6FWB
jCT6O8DPWlNWLGrCV3GQa656C1zIxOzCa34zDaklEvJGSehkDEpbKoXXwXPnD3DP
kmJzWjZYo1rT7KcXRR7mpu7+v52PHyEG6waU0aYJcpnaSoeT/CSvNFLFjPD7BTtM
Q7aHYYzaq34AfloKLlf0701zI1N7MNGzNrs9OMHlErpp7u98Z0fSRam9zGZ4Skd4
vE5sIHUibXm2HFtfaK4Xvcp/1B/VmOKTVFKt329o3AlN5K+TbbAoCyfj7+3oQl+m
K5gB1B/0xrBw/7o6iccEqTEZPXnc0o4qAKQiJ5JjiFtdWs3i4w8ldoqeomW5/BJi
fhR8jadoN8YlBxbu8BL9aLgzhAAP4sI8zkb+TXMoTPrv6pEnrgNPcaPFOjRcn0lJ
8Vrinltg2YsaSD93uNgpIECGmf9qGrd0l144a9dwWWHUAshSU5sYm7nzzThKMjhQ
SzBKcHmL0IlWGZZaLw3fh0sVwv0Rs+EKoeE2IxebDcmINKqYNLuGk44OUsVmvFGs
eQlHWEQj00ZUqVA/8yrZm85klyLX3HGaybcAF1dp5X5/QEanhYDzGh6JVZoRLe4a
VvGViKmgW7FThdkqmuZNi88cxD9ghb/vbGrqYIZF2yxdNfhu/xTdk8SVMhJzipxi
yPQIJbXnaLsiWS5Vav3jqMwt7k28RU2zip/Vih63rvfuU0EJLB+mH1FiYhg4gOsE
XnHjkKOWc3c9zzLwmSzUJCPJxjW+Mep73+XuJFthu6u+0Qmti5mwKx218tSpAzw5
pjHhbyU0HHdqsvV2z5r/wcOc2xZ/O+8sGYOA3QWmtzeoqmR4CZLG/A511W5dBtS7
9E8vbib0hMX2G/cRbd0mfT5j1QO6C3l/mgkPGGHgYzsLbrRSVD1clL/koVZkaLOW
yIwxIwoR4ek/Gglk/gsCwzBCseSpWg5d9JSugWKZsWp2cDVZos+XBZPRwm7sMvq9
bRa7JYkfI//WtD6QTpj0RFhSMrvezJWFzSp3SI07YL//u9ldgd2x5pr7sJqhgF+a
ObVzC36jRD40WfccNRTJYpva8FiG2By7NJYHk9ZZTKWzDuWXhvIftT6YtU1XEETI
b1oUdL3une7cURuhENjBYsBYDfhDvwMapFvr4HfSU63pztPvtzOZMl5SmLrWv8lY
z3iDEvtWFSDPDqjqflG7jD/GNR1xjno6bxbis25QAyZ+3wvUOfJ4T6Iqo7bCFkk8
Ddk7SkQX2uE6TLQEvQ/DJVTMW1MqU/LgODVfaqZ2OhpyOz75yOo7eDcDk3Roduxw
s/2dw6EBMjDLrsRzhRNmp74Oplfbe02wWSYwjzg8mWl3J2i45TpRQSS1o+KldK7r
HJw4lTkqjCKHXwxfo9od6ePzFCLuMPp8Ta9EPY5LZBDJR+hMVAfOLrs8CeBZ3eOY
9lb3PwQtlSjA0V9q3RWaj91xaaignIIAgy7LSkj3Mg0fNkXoDEPkc2b9b95Ie4W4
cxdg3+bvhnSYgiMhn/Zk+y+nmqpvcUMXsWHx6Uc9WavR8jZet2B4jp0xAxOsUQRm
VIGafLJrYssiTDrD/0Yycg9nFzTz4fTQt5X6DSQGuB+wWOHQhxBVB61o+V9cRLap
MlTVnC2y7ua8+9iHtBZI3q8+UvpgloJyrOgprQEO64lKcvm6ZtYJuGOgtupRqkFG
dS9cMgI1xowobKp8SNNkQ2uRBgp6c14+zMQ6PDhSeE+BEaFcG7L7k63/VXguKExH
fQAgJm4iTjOG7RHKVCqjg0faF3EsJuCNqqh+HnLkh4atIRe9ExrGW1nVpOoRMv8V
fyPswvSg/4b3U561o74dfhOywVD5ZJKQgjOXlJ9LwU1AqDLxuXgQz/yFVFgHslXx
OkRyPjqsMEb8zRb/bbKveU+cXH8yRIxdrtDjpqb92Lkc4+iE7LLscPpRa0XGbbbM
+VdQnhm7PFfb0ALzULt61ML07HsbnJLOPux+xcJsTCAqqr5LmAzyALIlJPK5K0Mt
0GdzVKwGHXHqilqqGWDSjzorvreujT58QXW2v4P1CqGG1+J12LVW/pubXAsoHD6Z
BMMjRPeVTD4pfC9PxBR3XI9ujTWJVl70SI+7ifEvApbnoWWzSPDLqPOFkOSUISgc
N/t9VxiRwVbdpeHK4ikxfpZwTeo9NkA9xMRuuZLXpaNsokLX+bDjqUCFQ5pqjrQ7
AMQpMy6wCL25cNyscigI3j+F7T4cjiBTjB8LKRkStVXXaABMobw/MfivKRXQz2x4
UiFOkvGjK6m2a4tGXX2oiMb7m0pbU1XzBlHLCpnSARlL3cKPxitZeo67ynVApXAM
zvAeQldf/Mu/G/4AZukwH4Knwln+mvhODfLO2UCady/rhqTpK0m5KamQmg+n5RMD
hXl6ir0FdIxwnHjZ0aYBVCjUswSggowXj1VEoPLkD1QGetj3qO1+g2JX8sHXzR6P
lU8dySQz8LB+ep+thyxptZGitm3V/7dGu60iFjUNvW2Ngpv2fIKZLG0wM8FjT+W4
YF6o7aKNqGfdHx1iNRvKmeNHmkF0V9tEuUq3yHaYtaVARxAePFcPeldxmMYxsDQv
7oOL5XHsNBRz8T9fb6Z1ErFY4LnTgqP4rM51u0Lx3SiHCq5dJJRMvWkI2kM3aR+G
UjLcDbIfwXHLXHeWsub+1DLVLPsxreYdMdzqzyyKVLkJmcKEQGdDqgAZ9/evUaYo
IcVufKa+pLjVhDQDN8v/oAjmeojeuHb84jm3gUhLs2YA+Tx3J3mfCsREFDLWH4l0
p42bWy81R3QsRcHTH4UDbhmuwzWQB+WY0PMAN+8biepAMozM/paayvuZfshaMV4Q
Xo0xTqHepnO3AyMRgEDZEq3JIElRXb7EPhrXTGCcgLP4xmEGtA92+aKEs6xWBIu5
aw1t9KeNf4sVa30s6nuigmwIxaIHJRE29RfNh1lCo9Op3rydHhkTlVAVM8oUTSFk
4Y1tnykCnXXkNrLi5/9FWrmgKqY1YeH1GZkT2feWOguGKHkgpQFUJur/KdSecHJi
xFPNAKkaopFyUP8KVxUilcIWGRU6qF21FvfPWAm+/+yD8MFm/jv5Fu9Q+DMhmGnk
U233EFdWX7tRX99BJbNkZM196aoKkv6e79sEFLVfd/K6Q9pIo/fySOL48ZbeIzDq
wRx8xT+NcTlBKrgoI3HruOd3UtuqJghxLh6/+kDi1IXjeFUM8mlLJdMNP6Bm3OeE
YVCkgYMUdORJHXuo+ilzJnco/qFI4PEko/8BwdxxFOV6XE7c/nSXREJSHVTudaTz
pNpkUICFAOB2YZhfOnpXVv3QB20Zrp+CYxCs510dMp2SB62ibUqiGBofCA7JTHFS
IPgRegniq4wOpLX4Y6s5z3OTXeGrfvCHoBaGkcjo/yXmSlNKeGI6nY/Sr6IT7ynk
cpvtaGIN8aYuFHQgsCQdMBDXPpRciHnlJtC2sE7dem0Xie2R0QltbXCghUVJfObM
wsaIpryweM05C7qhIG3b0PJhT8LlZupCzQ93GvO7VOSZ4ZZyxT6toRrycAhuzZqi
FvTRDPZQpwW+5UygdAfPOgl673kFWe+Uv5D1EF6QwSw7IlIW6G2wQ3a+1dsuegYy
Qc9nny6pz56aJFSFU0m5OPaHMHtLAsFpI4gdUrQ3OA2uOdqSd5PxAymCTqgiAGfB
V2i3kCCjWD1ObldmJpgu0GOiVIGztA459NZrq5wWDESzXwmUewktql9sMWOQsazy
bFILjXkYP8BuPST7l7hR8Xk7bgM36iJKlnuv3ZrQqfDxYTDY3dGG1LkLQqw/6krS
1vhE6nwtovPn5mN4LiP2yzCTfR0Gv0+FBIik9r5nH3A2qhGPdfC7LTm4Kr1NS+JX
G3aZmX4pP6SwWYK0exZuG+1IdYZzBk3i7QLDJ6SIegXAqMZzj1gEXHb3lUGxttJn
JSPL6z1iUDYjWPtj2TMBU8Ak9i8+ToZ9vSwvxJjMs4P9Io5Xng/wrQmjqvxD4ylQ
JGVDeB9Mq1Xzq+n8D069UjHdCSWiBVWcuqrhdSU5KTjUxShTYVFtipiwDb7D/yqR
HNLl/1L8pTKFAXA9zU+N4wts9gtYqamSEOsYCceiTJ2xbLjKawGNSy5hMcLOrnfx
pA9fudYMkCdwBfMpaEDQUJ67jpj1pmkBc/YLA8JgJO68CrfWLj3KH6+Ay3iNyUWS
mt2DzKOWFpO3Z85y5GNEIQfFbt1pr83T0TYviR9cb4Weh4KYdkEgcl/rd25Gya+U
qXc+dZcdI+rG8y8ttj/m+wmAdRbJOdnwhSGC6UCopJvUiZClSNKp7NdnNcWH7rXb
iV6jpjtCN0dPIzhl6q3ddax5+cbCw3YdHsFApQdk2jYoJ/BGUtRfnM3MXX9z5+u/
tVuJCfdCruDl1XnoEZ1MXdOzjDHLgx2lCBuaAGyAr58hQrovpAzlbhiPwzCrADYf
m8gv2w2XpHuhFPSu0A9FEkvlzLt9iPfPHfyRFTrP+274P47bXdwI/2NNINFIaWeE
7TxfseTc3GDairGudY7Tpx9HRHFrHEXtDh7xV3szq/5vLHQw7qgaeNGa70rtIBtL
lK31u83aSLsczBc3Huaj7e7Ojhl1dBk9RMx5H2GmNGtJEi+luMMUE7cxN3B5GYXF
3je4zE3GBhH2Q414ZxwfhAVX9r50oj7PpiLc/h/9qfYYcJV6fgd8WInirZPvltNW
o+CIsI7cmjcR5YdKV8s6i7QhbIZRV8pYtOMkK/CvpEFnC8mzdMSLfy3QqR0iL2gP
38/z4c5AaFC1KWxvlhc6k8HSGc14K52i0KSNJRyuq0uX0vGtrR8LCcMZxld8w8m9
pHkC22/kNCp5kuXwzcF+mjwR1fDk6/pYHOn1zdh/GxBQikvBUkZuzRdnbM2JuHDP
jNoNj9ldYOx7XBxr1+8MfBw5bWe2Qvgk1vXFYNSbOe0iZc5sbcBF/3mgO3hV1pjM
h3HJaT9FOiiN3F5NHLtlY43MSaXDyj66kVOPc9O8lmTZYM8dAEwtLZR3f0hTwjni
fGLAdc9fnP2FCO/mxzLG0SIpqpeaaGmEyHEgjHgeAi7osKh9gn65YED8PO2AFLnz
4aYOqhA/QyRODSItAHAuDscAKQ4x3qSdcBS+57pboSSReH5z1743LveVuppoLCWY
j94XU/YK/MmdWgkbVa85OnAU5m/Bu+PTIstDz3fO3HUrxCAX301Cqx+BN44scfl/
tzopS5MMG6STJSE1vCIMLSf8S8FcgZ8z/wAMi3+mrkQz94WkO3q9ERiPZ59uCJSd
B4dRtGI8dXE+i0te8YzBa6Skd5fVAhzRQk7iH+mria9g9tQNs1KyJewFUuPZJVfW
u+j6wYqpljAJVqInuhfDoa8y1L/mlMZWy9e39o8p/3HbPuJ81hSXeWZNxPWAl/v1
AKqKzLSvRwj5IDV2Vod+X2/8N3beSL1b62kpVk7wRW6U4t6Lc3FvfiEHXB9R73kQ
VrSxPAGgoxicGwqDYdjiFz6mqAR5qqs+46kdcnXLzyQHQ5IBKv9DR/3tp/TXY5ir
Glk8Ku0mlw19iqdFmfh5uDXh3dMBmsL/rgzOilX22MLm2V+9aw41Z8nLqgjTUGyd
dD+M9JbfRRCpT2FygLl2k9A5uErB5pTGz3bI9mdwzby3wlobc+BOp+FHsCGzs2CY
cwbCH2+o/p6mlfN/thg6WH8UvNkhrhBTPDsxlYuM6F6WRTheWYqCnDOmRPlBT1uW
D6aMpBG/Qwc4EvyKcXTOUDK9a453GP7TdPcHekRehgda76mXt8yCrBpjDJ399rgK
M+1CXsNTSLLYJ4TrfGhQrHr3iETvnO+pVjP9dUTnxQm6tT89KcQncMRS/PPE8ZLq
YFeoTmZ7DwhiqmB/W+okThUA3R5IgcmvFVJ0YnqUJNxWxfZVSaxfivM4i+Xhn8uR
MniZs/l8/d5TU/wDOaAU/rNTaTU9MsrbFvMjbXc+q20u9uF7+C8QMoR3KR66Y4Zu
HHGhpIWdLQ6wVAQ8z3hh6woxqJwd00iWB8uatTbhC7R4eiUocQ/3B9MdDMzMDSgv
/yo8HtIg5q8ii4bJcvjBNzgn0A/qtSng68c7QX3ksY2LnDOl0wJ//jvG+9sIS3qs
Xzea7QH3iUkzkr2LqkBxCe4TxPCm6Gqh2Q/Y4W81hL3/qa/9P0a9x5el873vBQk+
Mdsb5GalxoZbSrhY8dTcS01Bf84YW9x/sBxUWZaox0XRGIdmKeb9gbh3GULHrDkD
vohZ9ZJPPhDh+wdR7UGDHrTfiyMRJoeAaRp1ZsZG+CqkCjkEPO6K0JK43HdjXUg7
18y0JXwLxKAAk2swiEkMjqOkS4cZsLD6ZyiiQ51SLRrpWAWCqS+NxEFaNLNBBUcz
n7Ra/vSHoV7XzQLy2p23Lx0+qfgNysi6u026uahdmXYB+EyuOrlwUQfcRAok1+QV
ZUCZHD7Fb0j4gZd9/m9MruKLvcbxNmx1UgYphrgr7qjQIlVZHQyCXe4g0sIS7iwu
ykK/S+Tmx1uFfveTBVAOLdHQRUHrUNKjuObgApfjARD0coAhDV1AGol0eMoMcL9S
5s13+11yO+N5jq2bfm3DzqeTtmULPJw3IvRw0yR9fFYQYt/ItmkBaKFAna/rYkLB
a5GLolmOGAMfrQdzCs9AIT0qAVr/aX+WBhdgT1NvmH8IsTYvitBxkqSvjmE+4ehu
90955laGNLJl++4jBLAGY0j08WJOj1x60nOtw2Qq2Gu7+XddJ9QKaGCBVJ+ZselY
Rsm8Y+vbyt4ePidLbflyw7CEr1GHUgbnHy7qOX5TqY8Hz0k8mlR/HcRbHeg5+ZRe
MkJ00AjeDLe4ug3PA4vVA1yQTCG2dFv0hYA34qhebfKl5cr1bKH+axq7UenGNkfu
6J4gkSOR75myfS8qFuvn3p3zWebBRlD+1pDWHQT6V8iuklBGYKWloAKsB2xEaeEW
TumM6vY2b42MdG1sGe0Xa+NEv2laZiakS1ArAvOYGmqC62XXblhzzVE5IWGHjfNG
IzrBxp4oxvB77JknlxjWlyorqld7W3RCRJgrdYJywivC34Vg27zd81CJhuh27uA7
okUgEAZHNPp7LbcBzLMeknHNmGQV4z3jUufHdRyrDszxvEJapvihah0bT+zkEcw7
JKsVl7Xp4A5batzL1ci+wNd29npH6ZypSOdE4BCielScVu1/W8/qCQKYU7maRkFu
UplAAVymaHXI6YqwqvBe26nuEGMtKTgL/IFqHfCjggeGX58ZUi2q3Y4UxtxLse/Z
aklijucoZ63xWCdRv8a9JEwWnJIaxnxnAK8Nhh3HEBpuz+KgTku4alCcjMhkvZ4o
dPIO17RjVhHfRLM0dOQrdzRFjgQ0SY7KLbdfLpFaGTYiCRGKq6HWcAaZBqj5MghZ
jWNkzU5/A2f/CIkRzzk7RHL16IGWy2KzLrvB48xYpkxSVGp4VWy60kaIHekH9u+O
xZ0pJb6cC56ApM77uU2IYUJleS08n6WRrf5yjuQeV2bfriWwUYJjL5aKZcMevGka
1fT1zrr79KtZJJ2hgAvFkbW17kw6hvllsH8GWHPE6QHBAdQ74Hw87D0XdrOlGeQR
OG51bWyu177wMlH4d4yahV7hQ43aVYhyCaamVxu1YMuscZM8CDkmi26Ux2mgn02P
Jsn3JBmzBnZ+2ZEGHtlI02CvLjJXeD0gO0QDR9zdYB+cQlNk2JlarBkEdCiSmZDO
P9H0RxVTLeVkoUnpMBjy7nZ0MTrUM1auvETG+RPN88z5VZAI3X2MX2/PYWKktSyz
YtAmBcQuhQPiFhrsUzMNisf6I9fleH1L/0q9SpC7nMjUURHn3KdSC8xnyB4KjByV
WP7H8jMNQMp+Kl+0IVLJHwtjA9+YHp3GHrGoeeidyPk+eXwpkGbQWKD/4xJX9Dva
i0YNxbIUX2xbapPUMpd04MGpe7Z8F6WmXjjiTzaEkqVEAGStNSaEXh4ipS+CqXtE
jhFaqoy6tNbNzYuzZ9R0/nlha8NYsIQo7HHbOk5n1arGBs3A6mxniZLtMvzh2Da3
U900T/tUCobijf9R0SUS2bxM6vCzTHkDsZQre5Wx413cjNDHjuhdZs482FjPZ5XN
lB1fm7KVhF6GyI8w3FgI2XsOiU4lZWCwuXQ6h2o/N0zglCVe4v33mo8DAyulmto3
vGNlifcZ6LS2erhRJOPa/vzS4lQqX/XD3Ms+HY7uvV8NWcIkbPmhFLvg49FIgDV6
4dr9xVTjzbyjzERDwjCYzce+VmxQkiNF1n+Z59hnqHEGTjD1sM6At6btCUEDnMAN
oyhUngSUxqRHD63LnrjbTd9zgi3DUHC3WKb8UT1hnXz+5Wjq8FjX1CmaiyIwxxQc
DdbfYWamaPyMDyyrm2u6GGjf6de0MbXzuhVsnatcWeQ0F6MST7T1yaCxTaVLgVb6
gonL2Zd00QdOLWYNb0aZWLDIpfgO+e5N0mf+oB6BuOfk+Aez2n3i+Pi4cZOuW5Ld
0UX2soRRoXk5U2guS9SBx9pDyts+8Lc3OaTpiN1JvvEWRosJ0w6GkqoY3JNJzwBG
X4Ds/DtxyGZUa/PAoGkK9dt1HYVnzrJRAnIKwPJSn316AKFJ3pH3NrJXzjY+Ornf
g8R+7Aj0rCBg7mzsTmF7c3oqnv1r/CNIH9gEEcKg0m5fWYs4jQRM0G7cj2ks2N/Z
xXBCfTmbZ2/QDsKWyGvAjVQxzvwZ2IOi5EfNW2Sm9T39d6Bz83DBPKO2USj4VsLt
IcYNNtqT1DXsca2Rsg5okhNkD1dCLGkugWCFBjf86nio3EkRimRMWvWrGVNoU/hw
E0SD/fO/3oq+wLYK0w4d5FuodSmdnd6gSUiH40OvOQJU+yA2M8/be/8JPCYCSvgl
OogYPUMRgRDO6L3sfZTYeoohqzeZSqDgLUNlyiLDu/h1iL/n9nlGXvTFUjB4cNC+
Z7tzIFMVY7TLLmzbvz2jZM7JbQdA8M/wudNk5rRytXvWw4eR4CMW0WH7ZRkMMoqX
47yHO1QVuHWt5Ej7Hsj7IHxQDogMCwRW/RioZTB9Ncx/E5CY3lkt6phsRzQe7a8a
trzC5kDYNxYQBHYCpsUXWxtSwi5qYOiI5rRuPSqDdf8nfXgCHwCT+YJuu+EUbQe5
9BNjkcNiq33HMF/QzO4h+llzGyeS+Tbta7uxHd/XpsTQFfooGN1EJdjamJPg5BYo
S2nnFUnXxFHPOnhVshA9V+ToVaqfzVdeuHn7ZKtYHxBCtGJ4S8UgOiUg9jbjaavQ
uB/5efO7u6g599arnLJSx8JunvSjBA0w21dkkkO3dn+yP25AG9GNT8ehMa+NDyYk
iDokpOloxnBtl6DFK6TWpARpwPeGy1HDlQQy6ftfKDPHUIGwH2ZWINqk6KYRBZSQ
4vilUkld8boFkw1eKbSdI/5Z0m94w/ScH+ZUMWRlbFONPkgzA8ovrl0AFW8bqs9C
qzSdnZz6W+y1ifSmh2AOD0blHbv8TtNeQxxF1fRrCtHfxxW5xlmjMqOWbK+Q5ERU
JEBpluHrNeaTFdIP5ZipGpDg2iOJdM7wsoXC+OjBsayov5wumI1uCu2YATMFGMuu
i7PqgHf8f/aBvmsLTMn2PEZSO4Su6TtI+gx/pmFDdT8owiCEIoLDw4F8rvuRvIRt
oF81ejwHJvth5VWZOOb7XYA9jAWsVs4KK6n487LVs9Q1RzN8k5IyFgMEjbJ+CRcE
FrbBJypTRIj57wenIceWfe0RxzfgZI1fvWypIeVlyVLg68cK+7eiS+YVC0Njl3La
80xzcsVky8siTXGigQ/7q5CB+BoZT6u99QJ8seZHg95EF2+VIVDimsdvfz88LWoE
KOgp+OsGVbmIwbj5HH2K+1hdiJG25dHno8OF3OcgnaLFcXImh9vCfLUDF3nP8SEo
DlIjgLz3BHfloeiJ91Tpv2O35wBXTRpdFM9XuZtvnEKgExPN4qjVMzixlp6HRQk/
q4zZJtFoyqhL/cfSio16iI6jX7CzJZ16gpYvnA2jQILPhzs2tjeaS+9dvQbVlAdx
GsJsskviPeZz3tB+75SRipz9LQ/fGVE7MQb3Vp973JqPRsCAHEQhEyuUFjh3J8E2
QoTjz8II4PYa2hX5CDB+KjPoa7crhrytN9XIcFXf4V892ZO9AUTb4muyd3yjA2GM
Jw0KHNDBiSNu5xyV5tJoH+VnJNyWvQKEDrzrBy8VV9N5SX42vKnslsErBGRvPvYA
U2qVcnONXHFAqGv3mp6FZwcK96/9XtuX/7t64f2Oi8B0E0c+mlzpt7UoEGEunvem
UJF3lFWUgKyM4runBqp/r3a4ayUoZqa9JEf0KjmaXs2rbLyZ617zSK8l/aJtzBYD
TadfdJL/TlBRcTARqW3IoLF98gxFSA5eZbjdCLp99EoKY+TTfLdqtGOOTEnAaZiT
kqAcJVOd104hTU8Ebht/EBv9aTKt7ypfCnfbReo5e9z2MLVV2i/P+TeoDyshMWa+
kdw2SxCUK3dKAxbzhFW4z1hEjnk8j/1zu+8H+dGOdgYhAlrRTl2QadC05I85x10n
pPed0QQpO+VOiCYcpATRcS0oBbRXT+dryR3vhWG16gV6AcCiHi7r0U7X8nocTd+f
UD0ccGLbtVLoYXZ7fY2D0ZEHrsWi7SnoPE1wJ53CIhwW1KjcRkxOUevCYr0vrZsf
+vIdynHyjF26bhRUjVktNXX8M/4G9Qj3nzQxTSRbuPligUsiuF7uBxJauuqNaAO+
Thx25AUgphnAuBm+P0qqeoHZ9BXAI3ibZ/mFu9gmR0k85nEV+doLyhl8dLL5GXKF
qDdRjPDD8N7GgR+vSBYphqWZc7qQMhP8kizJ2hkRV2eXgCj2WZQPy3z3iAPnqkrI
UWZg+BQM36VlLmOgS0M7fr+trcGK3T126Q9z5tg3gfN741g2sLe4if8K0xYdcWE+
+4wgizAzMjivRiCNhknZR9TcYiwMUmxmJtlpfWwXLco8ndpE+Oq+kLX9wGq9H9HE
XBn+XRonimyF0EDQJkGKETe/sAFDCEOb/pTQLrduOyovvy/mu4Qz4oCp4UDZkIBA
tsDUBQodGgypbutmAcIK6hvYbp6MFpValNwgQRWVlul3dBmuDjSnWFEmyMyIV7hi
QF5L4h+PmUkQhvEQMVaUXKXgoahKta4dOkuA4/v2QBg9hTrMRecoyx4ChLY7bGqz
MrPSoohQCtrzagonWrNmnylDfHmvPABJJO9758Wu73xUu9FQ8q8V2vk1GrUdpW5K
Gh76l0/J5TjR2aPMVBmc+/+LNvdswAcJaMGMCIriOcP3D4suwseNIzUDyOT4PWe8
jzfjJF2i98NI3nU5HGsQXhjnBswIwASlZ0cYgB6s5hniNYoWBnr0186K/qzIKRRl
jO4519icMkipXSpatYVeWYD9uaRllb1FrpZajyTq84xmPPKuZjZYTMHvG0ZiTkk/
gLoHdWUuu8w7lgqKgjdCnzJEPESsAcpEV6iDc9jEZItyyk4AmnFuDCjwBVPu/mSR
ydeEewvwsmZ++Nhdz6M8+jKXF7KxySJ+kpRUJ2/GuWL6IV5Baee3xg5/X1fiaUCO
QQXEoa80ufp+1tRlK/A9K+HlmIEOrdnm9O7IA5ijyj/j1Z1R1poxqgWEmXg5jQeg
eRT/KjnV7ynUt51Ekac2ci5V6z5vRXoShCPX2nJ6n+0ZhKVVKpxFM/T6hZNg9fvp
hPaI2lLWcPiIPhmnvUwz0K1SbnsO1t6rPBZePdHqzuxe8xpUcxyX7LdKDhYXFEbo
zJFKEHd6KgmSW1Z9V6gOeEPSXwGbKi3p/brp4TTqbNSEQKQRWTPGDxEaQg18Odu7
ZsT9z7wD+I5zOXhppsiXiHPleXBzOcmKyCNX1L+e5LQjXl3CIlOdKs0r88K570Cu
THvVWZzf9zHiVFrCUs1MO2KRX5TxnW7tbnpebwnSDfx2+MrX0jbViuia8nOH4T0i
c5hBZRwfDrn2uZnuTe7g2uRkDMlUVTMs+iVMFTSAqq0=
`protect END_PROTECTED
