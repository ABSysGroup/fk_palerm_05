`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F6T793cQmVuF1I/xl/19S5k2qmYQ96m5dYQoVmmSU2jWLsO0I/p9tZnL7LxZcNyz
yjONOyGHGlUci6E+ryrK13gkQxvBQMZx1keXL+x1fmRLbqLsvVtgg7x9HE15iwSv
nDtmvIBf1Co9Hjf0qy9FOLj1Oe8lsSao8WkB7fK93JsprlAT7eKWtGYepAMkDMoh
cUKUVI4WofAuxs/BGYPzX/X7ENLCVaswPwHUFjJd9qj/ZhASBNmS3UYAWc0tJo4p
y4o7VnieIWgeU+QKxSAYMvl22yzQrxqvshbgT5AR6DJFpx67jPUZfKWDS7u89r59
cexnZsALGBmnKVVBDfkqAJxA/xxXAc618l0MuiMyy5WZsMsizNU1tB8J31A5X/5a
syfKJO6aUv97m+wAeP+yVSKptNL3JRjKW+aN1IPOmSC7lh/Da1ZHNblJNddXlGc4
w36l5vPF9xlln5I6kElykQ==
`protect END_PROTECTED
