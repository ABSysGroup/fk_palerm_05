`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c2glwd30zh4yzdEshi71J66tLPvs5f22KW6FxIKX1aWXQj2kqCEic/QjsUbkCcXf
VZrNvZgu6Pfo4MhtEhk1uFptTyhA7O3tBq3gcfUgRC4LnsiT+U41EUstvauJQGOa
VnUGBUMIBjbm/A3nwRlpK/RJgv9vloHzLyDDugW0XoCi8VO7P2ThtvDqR6+VhDoX
ZuJed9LVgiHbfSKLYR9m3JWuPRdh1tAjdwb5zq02cz+ihWfrJBigxNnmh3Fu8aeU
wQBiwrF/34BmX4/oPKS1iKRPTdY7yQzpFnmkm6q2FN2sp3fOmrAvhP9nYFpCOjME
zD4aBLIBHqueVMRKuo6vAJkCHzHEqwt5K9H0XWmcIXTe/q15d2WM/JYp2GCEuNRf
9InjZhJB4/uQ6PViv8BaHz5AJAwil4tH9i/0dGaQJj+icvFQxZ2GRvuoZ4DU1uem
`protect END_PROTECTED
