`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uixdE1cun0ccM5X/LZkfRhZm9ZzRpIAM2gRi9Dvff1HdNqypCfb90hVLb0cn+JCW
liSAtDMOhYr0mEtm/UeZuaj8MCx/KrFTQWSpyglBzWxJJpXer+JRWXgdo33m7HpC
ntRn4tB58xn8BRTYF1+XENeIQJiOnapgLI+DsGtmBGjOSUt/pSOUNvifgN3YVzLK
Wp2zOenGK246cEYGJv0IqRIB2OaeX7fjJ9cgwcA5pZPL5gV8YvlK1iWkqitl6NtS
MND4TA2Hi+jsa0N94l415wym0geO1wzHiDmwPUvXxobudjRkEJ4T+6bAOBmDsXcp
8si0zisOJHYx65ATwzaCgDNGLFrtO2VFsKmT/B8ECPpgtWC2CCOH5ds3VjxO/orx
MjyOuMFTc7LFR+XJdHcq25L9dvV7a/nl/Q9SW/Fzxa9XNkiCrlii2WaoAOpeyjQg
6UgFEJKdX4hAwbtINILuAV0WewLqExwooh5U0ph3qlymsogZ8E4N9r9vbcbQmkLp
IyWGCKPYp/SA3iXZXlb/FCESzsjhyJ+g8vEEtjfddGc3Zz/LzDZGKoLkQ5VPSl1i
lExc6LdTiGIVTGt/AYdzLaM/B97F9BsADyqYA/P8VwQAxidlx/tAD9l/Gt+E/kRP
PtZB38bSgWd0JpuWhzCmyq9SRzZHNV1iM31SHiBsuSJ5lthOpQ/VQAidZaeXkUWF
EVb6zlHj3/YfeHIVVzBt6MhLrTLvUEHxT4+6/1TsbdZyvEo2olEUsHMu/8ppVC12
m7act16nToZkDThaEMdGpJxcsCTJsn7Xh2ZVoIcjub+RMnTXDVnXoOAPUncLiujx
GJyRvnIEl+KYnn3IvCC13qo7biKolyi8vGMErYfad9Pn9XoZbi4B9iqqC2KM9mky
fjru5ErYpweNdcov5aa5xnHL2Bxi7pPnoGqMhzlxWsbqbDTuwE6BMa7ZeK6HNlsH
neI24H4olPXYHaKPgTOmXw3N8qXzNxQuS+Da/E5VrqboelMKRNTaEJp4E+nWDZDt
yhKxacoPGTXI7G8tt5ATA7VOTpz6j0ztr4LZdf4tDB/Zv25XzLn0zNSFaYcPj8MP
yd6vp7qT7eX2gU6+BUMcR8Ik2KwdTr3EXqZYFQumLTmTHWdrSJVnOa06OA3tI1NL
FBaDgDKxhCyu23OhKTt8vpgnp7fE3ANYho3FkheChxPDfn2pDqRt5APG3bDG9enh
0ovl9I7vJk8sKqQCx9FDAdG3ZHDCMzQbMVPnAXTKDWfJW7IU2Q9rdqlAN4SmkvVi
vK4aq7dSrp91xCbW4pTQ7hSgFswy8tpAAAN0OscyI0yJwuLSBkMoWVQVIoM3Ko09
Ps/Mfxoj9z+AShHZ7m2ngYgCKyZUjGAOu/qPGVyTn5zD4tikcSwsm4K9mSqRRgAn
Yg1YOes2rJU4IChGhOcvDBZQCyxTmZs+9wdXKnMGAEfNFD2FOcD+LgD7mUpDv0oO
R+z6T/2zVhrC2scGn3caNrDLiOlNg/x8NHM1OevIcQSY/C4iXdkCqklvaDwkkFut
qnIF4k7HyJjMQnF9jiNv8jibIbrlisjr1kGB3i0w0eNpcj8mqQxayEDeV6MBh1he
LkvaKsPVw69qWGtt5ofG8ocP5kT35v6ty2+FH+vgkSGcSwPSMQvQFpkXIkB+AVYU
3V27xT3g1JfKDLsQ00Rg/mc4GCg2KZC5mu7tjxs9tSuNs6VYj2U3EDTXlkCMgf9m
er6AGaf1lsLiVbinBeZRrUap7Ccen+JGZxqfleBtQ6F60wkgDIEOACnDoPwDUkpO
VJvXmzEH/NT1rT3XDN3A2Xx6xRJPpFprIKAVxGloISXup4Sdl/dn7CgOmignVF8y
pFaO8DMFBqGAwW1k4CGxZf/vvESrgeldgvXF365rCYsYbjm5UeG6D/uQ/ih//DF6
pUE0SFfrDtzUjDuhAa7oxqv3UoPnGcR8E5gnNZmc/8kNNhv+8Zrm2a99YSiLsw2c
Y67DWqvSIpM7tbxH/oqLIusM2qCu7jCJQXH2VYp+JlMvXk2Dwpmg7c6CBE6qscmV
GY8hePNtyigssCEKKViKCw==
`protect END_PROTECTED
