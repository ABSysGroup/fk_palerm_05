`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JEMCWZsPuijLBhZNntcz4WrJ6m/YDdJXGlOyFECoxflfZtvcdeAP55HK9NEVVQm1
yzlcgM/IHttvdaC0BMJCKedO1p+smf6lj19kD/OdRF5caQKSDkzq0SJKvbn0SFz0
m1uYgROJQIhvdZ/rDL1VykyIaZPzm6wbUP0Gp3+2NFxL8/nDsq1ANoXZRi+C8sWj
B4psDtPgbVvDGAw3stOOqquK4iVhb680bvAOVlbmOQMuGkKAjCwZ15GqW79aV13Q
d44Kpa8bmi5JAJgyfUOYgjvt/dtB8PYF+NUCP5VdVutvaw/mRq76uhYRqnRica+Z
KBs7OSWnF4vcX95SBiKvqN6diIQR+wzMWmva3zTznmankcaeWgrfR+79PmPLvH4C
hU0O9KncV6E++iu2u+VPOxCCJbJYmvECv0MEqVP81xUJrnBOK/Ldnftn9kDrWNaI
d5ReC+Bi26NxhV8z9wnAsCgBNyNCWkfCACnk4IjE5Pv5UI1q3d4r1xo6cNvC/clI
vkzfTm08XBAhNi/KRbi5GskRRURenAVE+vsluDiGh9LG9KLQmdfZdq4YnwVVdz2e
3IhMeqq99KNtZ60GYROKbQHK77htMZISgtnUXI30pfuM2Y1fMA4NI214XxYpiqfv
59qv6Ps5GQ86Lxvj4DkBMOa0byC0/kTIC5l65kJ2rWfCCDDrtwjBfuMbbZNTQrLa
JcmszBBK9U7JIIUaYM9oG0ia943thiwOsH9QMNgCfPNIHpy6rzIoopFfLkix3e/a
X0+qMMo/SO6Jlgj3vcitSU/P/zqwMhsfl49cwou2IuDH00s2/NqeTxGmJAtRKLyC
NpTu7SGKFk7pWYmCn0PQPlTcJ1DhKvBlGcC220b2DXl5PEVfa8+wGtvgmgbuABhZ
CSg//5FagaM2+mNGasCAjlYXy9dUi/T3OAFJqv2s21ngAfKXyH73fc7wDHfgtd8V
zPhA9c//ZqGN4PntvBPtFDBF4YRkqWnFoLWNoniN0TSN9h0oY/vr6uu1h/HceelM
PxJ9Q6xley8zRFPTQuWBAj49RhXxHbA4AHO2zhl7Ewf1fbE6niIrK7Wdyy5uB0pE
QV0MF6jFYgG8AutavsNQw2ktdkxcp7ObSm8qNf1tvK8=
`protect END_PROTECTED
