`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fssHIiv7ASuDGzgAekUeZtYF+87jIKUhIe7ZWKfnicQmANsxZsh1wOfvvCye9izW
YnGdakSh7o4nI0G1y/+W7rxUvX2kg0R1NRxe3sQrbNqzAZSh4aX3aYvlXWjDCnLy
6IONiV04MnatbjqAgiwmSK7J52DPHWMy5XReGOLYkNjDy8/UGF4CJyqOq84zmGHl
vC7joOZ6lT2OZMm2VWKxd1f6/C4E94kroeslyoHMQybYmMpCzbUteYT8EY2pdBvw
7wzoMxeX4a6b2oQn4QT+wMThbhNUhI2OEMeCtREGtOjKGxlNBWpXZYd9g4bjNHa4
JpQdSbh3kjiHDfsINRiS9vzWnqK7vhbxCuKsxHmRWGm5Zw5JNnLPlBnHJ9zHvtFD
3DM+w7pQMOYhtre26znB9xOz9PE1PdRfd/us60ZHOallcq95IqD3AHMaNdBxfMJL
d3nVT14A2kEGG7b1laLq8odC5zSfrMXdvgzhJemlsRifjByBG/Kg/Px81j1IPYXG
S05+9SdkQOrW4VuZ9DVupHbvIipIa2HBM2d2x0p98fZgXX8g9AcqzM2QsLfsXJ8u
wjvLUC5yNCT901AzMBOcc/2AdYznKQLIJprUybg9ohH+RNLB1h+1AhPAqge0xkNJ
5wKtwBFh0aqV2fnS40xI2QQ2CtnelF2AsABgMCZN2oeBJbU/aj+FkIZS3Njoxwl6
UhKugLcFv8U1o40AD/D6nEQxrLHTAm7dRnxgjZOx4CRVzeDG1VxZJw3XSqjLBkSx
JMa61xIrVLXZwoRQr9ovbYRJqLRi6e4NOpQuWqZaML7UCsrfV0CMX6plSjONvs4Q
x0KJC7T2CvFO0vkEodZpeKBkAeqsF7IYJCqqV8+Xsu/LF2rJUnMrarWg+L6kvXbA
vNt0NNhvj4/KXUHT7Pc6oHExKR5Z3VGgg8L6ym9qBfwsTzUlftBnmQJZexY1UZFy
X6k0AX025zlwnJx0rCq0+jyYvgMXcwhyqwPJdV2FuPMZCIkGDfULoqn55s0su3lk
jtzrY3sf56L+FzE8hFbC4HHactO26eYbSxhzppNepYw2m7Jl4EfRXwutRxfPwSdd
d2HyV2kKRYJ+NhN9cJ44vQ==
`protect END_PROTECTED
