`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FTHW1hGKx76Zx7aSMf1TvPWpcm18B5GAHri73keMgNzdJIaXLFibNdlutkvItxsq
igRRN22FcOoxo+I3KtN7uSdlZOlh17nvWwQH4sOvFxciBN8bZuht8ZRvFhsvioFx
32+qfNrHfzTvGTd8PqCxzpZzr9V7ZEjanm4zAp/hQVZos2YA9YapMcJ3th1CRYuR
QwmzUrAKSM23vh1Don8wQS0OTt2HG2oXgGPf586ANbj9h6ebYBPSCsneE92t/CRn
YC742+OHQUpU7050GtT/tAsD77QNCIBGPXsN68TO0HTMlwyBf4ks+KyJBOx0MrAV
YYfohErmjphlXZ1JhkSzf15uHjMXc34u92QudSpfQbgFPJtP5i41tj8sa+88RyTi
/3Pzqw0M30Y4mnjowKihuMlZp/VPg3dZ93O0jbxyvn5R1ofU06Ery44XbtHU247m
NtGCBqPHSFbTFDewvZTZASQigjmUSI4xm7D4X2B67d3FFLHjQtALMBWkN9u3KH+L
4E+HgiADNxaKIr58zJDWUrhyDgyPKCO+98QO1bq/lo709+PlXJdDckzT68IYB/E0
5LLnqH0wU83hg8Z7nT/F0CIfIqbKAsor2XsmzjnRwaMWi6qydT+3hC9LWuBxSAqk
BoSL59Aiqx5sPiz5AV/Al8RmoENIlqmTvxLQHe0/9/jtpk6G/wIcoWEcGP4npQ/e
OvxLEG6olvCA6UsFeA9YF71n05Xf5TXZzflyK20UqUA+bXLtoDtVjSmj/I5/icDu
ktIW4T+Zd0ZBl0fvTL3ApZ2HEGVsO61IGS26hNkkSOpPhrVFbQHU9SdZCTuog6pU
4DW2VXcLjZQmwme7gYVYnUjmIK6iwEPZl4FL2ZD2JwL0fARSeGUI4aAfdeAWCgHI
EjG15O14/F7m+cw4RzZ1P/Mr9ZpxFgn38g33F2rwTjA=
`protect END_PROTECTED
