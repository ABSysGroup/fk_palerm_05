`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rxQQcC3eXWrbBCmzFe4l1gXODA37RCSd5AYy6gQpJrAx/EXsC64e4rF+nHJ89Qxq
nIiSRrPt9JsF4itg4uFdGrtIAG3Kwp5FQXZIlLu7KMRJ4gRNzePeSv0CRDBPohOw
uXxo23yWtxqhsuyJGU8l3wS5pxnc+NOzmt+n2tIf/N8YkCdJxsL0m0lRicMlGpoG
KmAO0GD7JYB9bP5eh/eS1gbcQEhcD83WsaO+SjImSxKDovDkgCIWRVJ9BbMoZp3l
p2iGl1lIkw+Q/auq+FrsEYR+ZzjtQPw5rURYSJWBa9i1iSEhFJ4vMakgY6q0QlJz
lU1pFJQiMIGGsbMcyPSVzy5Xm+sICzkJ5dnZdP+sphTojp5bHE7v9MpDXXpU35dU
Pda3SQixR8OLhF/9Fq2K0aOb3dEhM6RCGAoj2p9MyK0DRn7UfKnBYDYRlKDIiK3Q
`protect END_PROTECTED
