`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sXGWIa68hqqzr9Hm3eLZGAY85+Fh7QSXoV4GP/cAdCxBr/ZEp3EoYtmErlacZcHI
RzQZaffRQhepbFFd3HUyM/zx5MxhYKNVOjzqMj9ASEADq0FCrt41yzz/vFJzIzAQ
h2EY2t7cQQ6Qr9XmGJO1hbAxNmtKZbjlChc4oYPUQ1uI8bGm3NqoqBPRRhsUVFKx
CkZkvN0P0GJdXBPgQtOUUvjOaU76HNs3f26w4oKDCo/bK0Wq7E/iVyd1R2wMUHad
VpK8zQlF9G34jZTKWVxSIRI2PtNa7GwBQx7oFfL91sRAbT1AdyoVPgyxKE8EfAlt
lj38c8LQE7BMMTUJoyHc57gVwAVnToVMURGLxlyAV50lbA7jinbnH3STACn35ju/
8Wv40bfA4VX7ObL8hPPROrc+fS0vsODV6lpByc1yuZBUR0XSazap4CYsh0Jpt+Yj
J2snACa1JC+YL4TN6e86iobr66zk/oD+lWQG2UO1xqa7bioR5TbEePZIx/zCkPft
72/Bd4WQPQho1LO46u3cGdKRk9sbB/91G2jUCIgEkrclVUaPz1mg/8J99zDVNllg
kSWrc7rPlPShkqTLl74jAqYARDNChuVfhGQVjscUEb+LwnZRKwi4MZgF6DNcJAKe
Is0Z3tanwcjg2FwSPO6ixG1gdWX8vnlE8SGt6VJiR/KAU78gv7uWRgM2GML4A02g
EKYZ2VhUxpEgSsVm2QxF5VHYuQPS8OgzvQPncyNBMemSxDICHJ9JkHzRSlP+t25b
Bgqnngqwuj4RdMXwVIleKbEr7bexksOy+0p2sHPFrRz+EmCVX4y9Z60a1J7ZZjlz
rJ511AGwXSjsROh268oI2hax7Y0uaxV9bNdqcv/mj250ahXkuQ/Hag50/ENTopG1
mivuTOhc3XTmGQbQzo51OUV/oLuL8oQS1RWPyFqEuV/cYzHa4KWe7SraltRD/O7o
oNrxEC9AD99cmpAMEMzhD999XuPDCicXVc1cUBRTC0FKdWiey3r3Jo5nC71czg8M
kqqqzqXLrgxuWI6i2TH1IvfMRHXtldvGAsqcVN5ETiDdolGDK0phd+H+DyKg9wK9
9M366D1P7rr30/v3lZg9KCL3S0VQryQtaa1ciinxqdx32ZC9zUvNp6dguTIin2X4
bEn5+pTg/nLhmhyKyCLp1OYxp22vg6lS/eYCK1zLEIFUw7zscJ7ad8/MEp1EiKGV
fYWX/rcKTYyg7Ht0d9kgl0yliu2fL0zFinVdd+HMYGUkCiF87O+BFDQTRrc2iH0Q
7PQjxUBxQbBf++smI2AUvfOWEYAOKdfMkuy+RKDfdSa0//UCX7ZGaCeH1N4P4Opw
Dje4Ox2AKUJ5wI9FXSXGxZU/6NveYZjvLKxbCbh0w5hNCbGZc4ob/gzo+NLo8ppb
HE0+Tnh3jXt2D29MG28pyK3sAZ401FnRWtir6p4XO3KLOLM7Nxn24wxjgTdTZw1/
gwPpXfGPAcQF7Stka4Q2OaRvC10kgPPXJEsrHB+khjRTVjYr8EJuaLx5s3SN+Nq4
E0kXHClzqGtUCvotRoTKmVHUAQfyGc5CIkATCYGaE7EbOFl6a5/4lpiw6fp8+PQp
wvCNzsXPdLC7yRA69DId5OUgxN59+3Z10UfiHIHrt4bm3v2gP2luH8sI/KbT1w2S
TVpFTG2NqgnbH1McF7qH811UJ3lBmm4N+aBAcvyC05F5LMix05t1sKNTmHeXMxvx
cp+nle/8xh7SqkMyRYTY01V06Kn9jcVZLFRPFkeeQbsZ71KLTRX2TK7yoTtLBvhQ
k4BSLra++sGblBF+6P4BCR6Nx2qvhlosHXCU9VAKXeY=
`protect END_PROTECTED
