`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v2C0j2knbbsQkXX8fyzpMJc3D3je+7jcVF6UhnMZDyPHdlM7VwqOPhr4A0xvMx/v
cF7QJp4T+MIjphdMX9bUC/y96wH1I/BQP6vzC8vZK86bI9+qLMWC1babuqyOl2h7
LlE1d8HcXUclMLrK2EooAt06sHLll54rv/t9jHf8LsXvApfX97xH7dja57KTCl3s
q/ZHdsFBmPErzalulbsGkpCf+Cs90+EjVKvokvMOs+FkFG52Ejsn3lG2Dfd1NuHw
9dXxWtuep5gs6Ng/l9V8PCL4kgetfLyO/L9tVw5yif597/PVPUZ+JYuW+ij+l8fT
p4Ak1BAjQ6MjTIX5sdEMyCXRSzaaZfiYYcL4LC7gzzThfdOtpb3LGVmWvKSNiAEg
xKIPYQEjZrcwjKXGRfm/0KrnaKUri9lcnBnp1Ss1tMjvpvZqCowHX8gnjUdulrd3
R4hoZyz4gXT3+md0s8ru8tDeej5fWsqUlzO8HqxQrRorEf8cokOd4NcF/QWHgCag
`protect END_PROTECTED
