`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4T5BKXpO5WXmAKFw0SYHW3vQxHq3/BA++WhOciMhYwf3+9rDLMxuRbdIs2BkCXDB
+vZZ88QAik+aVDQpXJTWAFu6sqtfB5nr1PClDtlfl8DErBGDkumdGpe19uiR0iwr
0aW8ck/nAZV0wf2IKuW5VrufHOO9W8BoheL4pV4zoAA5JcxyMxiSLkyniIXBRQdM
vFDQ82DlQmiugpRMVOb/HlQ88TD0jd83u8Qj0dxRLP0DS8kPtU1hidf0aJHSTbWb
Bqpn9dWcT/wMdDEHNvHDhWWU1Ijd2PHBTYGFKyBszMSFYaE9AuP+n6xtRoLctB5y
2v+W49zPJ5g/CcQLa1tp/yjatctuFa2hoDJ9mbevMu8s5CHeEHbZBnU0lt9YkyXH
K2sLOh/DyKZSGViisgT1VpNMf/mpHgauECrmDTxQXuPcy20Y+ey68VV3d+lbB4pQ
Gx1etBVoeFeIZVcwCL8xpBOZRvFf908jafpGHvQ1TsRQ74YbuM1yJLuQsJsyE2U7
T7EzQ4CCdsrfepPrNaJq2z/wimms+s/xfVyg3tR84G5UEUTYw5jZKgDq/vIQ9q8O
MY4y2vFKdehfEa69bADwKBRGEyjBKSFlTW96Los/ExuFYjJ5s32CrW7h2rcMD3yN
LFXGkrTgwT3klGOabUKXFKSZVVjR7CTxVyAwkTg/9IfOXOttpr/W25R2q2v/CgOW
6qipjMu9ImwtHjw6klO90UZI2oZO0hUvYcLVUknEaoNkM87DgzoiY6wuB3G2Sfy6
MKduB1N6iFI6w/BN9wnDhXQv01sWqTWMJ5dpzdN9xKy6Jp5Z3gydk0TRxRyBcOSd
fHE3dPW79tooV4PJRsPSO6Zf8hTDR7EQKVbpHt6dQmYBxGj1EL+reNsgqfPalSXt
mDQO350LcGTrfQ06TxU/M6SKeb/j8IfsqtE18jzH7x95V2IC84ffbOOj9lokT+zY
Te7VoOQBqdaO1Nnyb8otexUvwfNJEDFi73Q6XPD3tLzIzh1x6jZhWhP+ZEh4Ih87
r8WVvfnpznRC5AdPkUDmvWQL+Bq8JTs1A6nfTjVJBCqIKbBTeceikcDxzGvKVRdw
Af+pPhrmeLDGq6I+uVnghNhaqmOU0cYVHoYzIlN8uh8nRm1gAgLdMMlKRd6vulvF
6BIQ4LDHwuSLZjtPLc8qijQLoVYolD8NGPP1dxc8aCxAqh0tXi9hFR/lRB6N4rsT
zdpLKr8SM1/oBqflIeIrT9G8SFMINGpIL1yG/CHJ0xvdjvY4rI49pXzEVN1QLSTm
J/azkHT6DFwbd/+7HrNoMBStEti4lK64WeH+8xNe+UyOHZYiG+YE2oHhGKpQ+ZjM
ir3GOGBa5MInWhZDMcSLbosGQtXsuZ1+3g0x8ScnG2jd6B5KFr7PxvwKQrYd8CXC
XSxwylZZKB2FlcqViNrPTIiP+4h7zW6YqyKtIdptF2e2vnBcr5xMEpthVoUOW+2C
jXEhPkhWy8tCzMWgPExWaSZWRjunm9Re0p60Fmb9bkdzZMprf2G7uhZQhW9XynNA
Z9gUFUzajv5MFuS6vcM6EQdGE/diuAbJqAQH8UnBYioN8+knBvI5o3dgwzSDfuJN
eH3t47yoT60Fv6LiOUjYSJxGbWIPozarT4kvL5O4CheMsY4FtCqIpVP9ONnPwyt1
Tr6+9zHZm25iH3gXGhTfwq8o76tzVyOoQ4bGI+yz6YipWY8eP7jr2D5w/EoBqoZA
z9VnYghq7WXRaWmHlbY8umHQQDW29oaXS+32FI88qvLyBj5piNsbfsgRw1SIG/cn
2D1rAF83Ju+eEYAF+CHvF4LA/ovjxQHHgCwO1DGJsE1Xb3rip8b2+k5Pi7bc4DDf
4889HNc7ibyeWAIqlUd/hYZjEK/dwZ4YKmxLm2411QIl/yYkfhXEkhNpsjNe6VpD
+O3puTRpX3lcASduiQ4Ag7JCkuttZR/u/Z1mkIeRnomKxJ4AZ9GLu+KOYNpUP6TG
z/1kqb1FnsAWZHzJ3BPPXDGL5GbY48bC+i8uXEo4zKmBJC2ZFdvw58ymeyZgEIE8
/yYLKDjVAtHgtVPf1bD0Xuz0vrp7x7aUYLPMt8Q7apTKaB/gSAhcoZxAWRVeYnum
+XDQB184emvcd44Pw5fVkfVKoroQlGsloiFdrbJWegub7wTxAAV1TWpJ1ipOew2N
2h68OpOtvxNvdMCeP5WW7BdBS5ldidicTfZbdzf4DPErj5hKZDrLb8wQio3Fj4oP
0sbd0P8pR5ohT93QER1PlpyUpRRzjafUHzFzfJsvcojxdyZwaLtyROGBag/OIjOm
UhwbTPTN+oes30fwyaohYEqvNu1WQvMElRUSvbzeF/jeSI6UCHMbnyuCyuhZPyui
0YO85R50OKumFflvC1KmbCfR0TynU4JTvhXofzUMtm5akZ3UiQGFOw7aqFCtqGjM
3RhL3ApNH4p4j8UDTC2OOV3WpVR5Y+HCBDSbelo77gj1oMwwRR4ZoAHO0V4MMVub
TSQlZJmuYTCzrujsPkxXBGMrRwTKV7jJLsT1Y/zyTh+xyFRSnzTZsDnuhJLRE5mq
qFF7JKVnTcXtBS72DwRh62b9CeObPh5VnPEEiZcRpBZwKQPo/OeQpfC0BDrWuuyq
Ut2NgLfSiDSLHxouk7pdEw0WZx7U1icN4jSyVU7e3GYFfOnjKKpB7yvbnzmvR9QM
wyUrsa7DJbPqZSbqBDe/ubGMAimZEpkcrAJb+fm4Aq/dCPFtMXhoIPXz5l0Y74ZJ
ZLShHoACqDXpvtf0LkYIwPWnuP8rV9Gh75aZon/KClbwlVsZygwo0P8s0R4WBmR8
iPFfNEYaMwd2jcEgvjjhbpl7XF8HepFrz7NpDiBVHtsr79CH2MJQ0LoB/z2VcfbE
FcYMRt9PxAcW8WtyannZ7JlDbyv611i7rrzrdUAvoDsyvBtRseTLZ2+2fOvyepfl
Q7NkuysoMtOLJPxVmyVfHdAEu2dpnawW4SVcdkp+XOS/hQyuq1VpoR4b8t+Rinij
FR8l3sIYef45Ut558KIDYxyUw1+LSvVc/QO6CDmrvkKnvvYs5qC78QqgEvdT8/X7
hCibjnLLaqFfVpbG0l+H5vhrLbTZBYwWKh1PdZK/DiCk/eg08EVYGdfrdhGi5Sas
61IDV3wS1/7sPhLkeu2v8xzyh+Z8fL7tVi867Uj/+PQz2coodkzgR76wxzruGb7P
a/Wm8xdr3aQ0i2i6HXlHeKZOi0eLudF92YqYekqgVj9VFkgbSiv/tir6wG3qANEZ
7L0fKwT0OnIalyUKcbUdDTpT0u1AfOcWCf9147W1v9OZdAtCbdrm2V9kva8/fboN
yKTv/VkZQ49CwRPIxJPxgCSPR1pIR/n6Q5c0aqyk8NDzgZP4FBQDqA5VmNu2Xx/9
1LsE2sk85ajWAa76i6gVtm4jXIo5r+MKB15E+hFi8/rfh9uYamVCa0rlXgrRfvC/
A+8oNXfJA7dfWysAoG1LxcZMBN5XKEfw/u0/rJCOW/5fbtmM7TrCbN6PgycTBXlA
H6yLPkifJhhQ34n1UDNRC4/osm2GSGL9EYd1kHopJxt6akEvgdCGwhn4E3XzJjBi
vj83p6IVVbLOz1vFbmby9JpNrjpHsdnoi2rWicGMk605GP/oiz1z+KrwkaKhgfBU
uSMta+v6jGoXwC7MzntP1wENohfMaZuQYExYatz/R3lmQhl1+3HX2fj/zyHHg9w0
9n3Z0EzD2eOIZZiFYT6xUYu3g5ArqkUchUiHI8qtdq+rCKAsgpaStiVjvQfwv1ts
Cg9ty9nD3H0LV8FL6Mcs74OY/rPxAUD5Jm5Jisxr7CeGwB3X3KvGehDomIO+YuOI
qQMamhdAEPvJ4+0aLyijZ0d5JlLO3YRRTeuFNk82beUmVj6tY68h1KeRPamSeQEx
XL9soEGem+ym6XWA+Vf8LWjvPR3EvDHqjrm7IHvROIYOV1RBN+GW4pP2EZ9as8GE
udLL/7KoD+etNeIqUlX0ULwKF+DXSitKIcviZ7SMr8UdAaHtMs64NK03HilWtyRl
`protect END_PROTECTED
