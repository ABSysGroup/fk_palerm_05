`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0KRRJZphwjujh6vdnuqV6l2/pnLO364lJ8yH8FM1XdIMd8h73u673Oe7EwHkxfgy
mu0N8X/S1ZQ99Ly/ntOSumiz4sQe/55lYNjt6hJL/jpxqdajMGwAAVsFgaaXo1YR
jK1ym6ALL5HYdz8psh03HrA7ESXECwE/V/kQydTA4yyIo/NF7gZv+/UoFqTsO88f
F9UG2hliiyqprpO0uXYnVFGBpkjDACT2wr9wEnGhrMQ+S9qNrNMO3iDCGVoYYLr3
Qn1VySz4iAh7i3SgFMzZzRX/c1xYRVqWQ0p1Nzxid9/14v/QrdbHqnjrHMPPbHFv
YDSE5Z5CQGvBuppwRSIu5Q==
`protect END_PROTECTED
