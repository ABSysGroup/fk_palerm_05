`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1kt0bNUlWRrs8Kn3NbTzsow4gJNsr0EAAOLeNoCFqwTShjyus3bri2Jjao6KQFbI
EoFeiS3DG39wv4kO0D4oz8WOckFtcJgTbYASvP/HbZUDXsLEvEWyR/Ay3gsS7ZI/
93OIz2YjckRcAfhlw+dFn35o9DkRvRKAgAuZbIm0fTZIJkvVmEgmsbWvT7vIKDUQ
waEWuWhyQZCABWKzbKkvOVaIW7wJsyo9YghTekkgNshS4WYSRk69DSHstANw+Jlf
6qjBObJjFnBW1l6CyZTwqmRdmYX5yTt7sEbuYuwvntaz+Bcj/LzQHTgHaEvN1w31
F7oIy6QkIejrkMAQI1kWx1A8lP/Xzy/lR4ZOB32MA84RmTxo30nICjIAsABJ0f8i
`protect END_PROTECTED
