`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NojJMWe+vLXVtZoMx8gEMOCZ/ymbOwnxUdKWPpKJ2t2v4TgN0gklaxpO+w1QNYqh
lwY9IH7Mx7j+bW9YoZ1YqfuopdXUNehOS4eeu27QpgSJ8Aa8F7CBm74gN+GG1AwM
+DBR75JKntcZCarfpi0UVVfaxqBkgMjtkZi++eJzHd3hk7ceMlFdVY9UKs+XdsU9
SEa8eOHFlI50ujnr84F2vjHSkY0JwonuE3nxms5CmaOsRqtJ4TnIX07I6kKsUaPx
mA7mqW8bhf91XTQW0YnGlOEjOR141nm5ovKeb+AzdWtTpl4J1KbXAJ+6myXa/GLG
LZKi79UaFrF07PzuLx8hG9+JG4EympyvCGkLQWm75HfyTg/G/P/0SO8vFjtxtZBu
pt2EeBq6G2Dr0v5Ki5XV8udAhGNm+w9Y34X6lzG6lgdNFwUGMdKr6N2Jb5beeJZq
taC7wGsxr+8I3jHQNIBRVgPGMWYN6Q0m4Hmi5zPnfB3YbtewqgtxO9577q/MIoo6
pNXNTYIvy8KNnY7sddocL54kIxMinR9DBa04Deb/X6C3mLtE2AbFX6+s9+3SjBnT
fQqG/Q9JN62ZxaT77ot7LClO5BT682nCUgb1bpuTP2mzdbczrIcRnXijBAQATaXG
JzrgbGjmBNrbI4beWWibbBgAkHc9VyLVNQeEN+BReu+C5eVFHMhnM7I8n2/Euqei
G3qq7SR4BkmiA2pCwFP4qNuw99WrfAo/0ENN79A7l95SLvfTwNrWAkealJk9wt+M
0JoI1uzU28WU+MZDRkW3BQdmWkNBxot4q0Wj81W7FcEQssRUypI4pusCd1hoYo26
Ikrr9JtAzJC9QziWBjQpltztbWZmRv6oxBfqodIgGvhnsaHylRzxxLaRuoVt9k0X
uYsG6degI0ua/XA3DoqWcg==
`protect END_PROTECTED
