`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d4AODZcrxX8JKNU47T/Z/x0w7GIKyyBmzE/XmDqlVhrOgJbid8T4n18m1RgzEYVI
swlYgbVRFfZn9wBbRM1ez+6QkHZLXz79aKFpwj7hZiBKpPt1kN3eBrA5u5Gxb1Q5
FuQoAi8JkITD5PtWmr/TTbdvko71z4a8hC815umBc5ojMJJQen+1SzgdYJl/g3RJ
i7PO8vR4iP3Fm0pOB1+LiBdmggRAABsbR+6O/2FpP+ZkBLH8yerC8j3Q2bMa1b3J
Wuie6WEUoOucdYkvCOaK1bPNSfE+O1BjLRXC/2OaqyGdIuPJ9QSiRC6b1L8ZhvuW
evJ18/tISw46r1MAAWUQ3648CNPNupK05FZbXT+wX5o7K5wLSk4rdmJIBzv8PfGE
Yw/f2fek01bnjfGCmaMQSmLXDvueuQiVhujUb8SQSyBpVTZrI+zxgBRIbENEd5gY
Jx34IBL6bs2BYXPkf4nII9N8tnm+smDMpuhvuWYSr500XvTJMgPlo/ELjvuRmtTv
w/0odDf1ipfSGZoOHqfKRvazHVZgqcp7KnlEL6MEVeRI8C2ZDUT1lRtaw9+z0xfy
jX/wfUxBFYYQobMUU+hc2lVo9zmuvcHFRYxuv6JdNPA=
`protect END_PROTECTED
