`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0hPW5KFLEqxrvICSKvIvmMKSmhTNyl4drF7ZKV0hNDQnBIbpEXcNeuMw17igoey/
acdRVApFBxcW83lRWewWnIlg91yxCwC86NzU6nf8BgiIV8VcNmhiGbvqnJ462zAo
dGJSS4yvTQtYgec0xDT61nFw9JqTY5wtlqndA2JXTfeCPBNJ8JPex/m/ljGu98x5
eRZZhuNvZxkduYuYuDXWrwLWGu97D2i3V8D6/BlXYqBe58oZnoixu56/2FaYty5U
`protect END_PROTECTED
