`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OkN4fKDJi1M8Rz8dBN6ykuHhpw5QGNKStD9fEfk1JBAzbIUwRhkX23F419Qb0Tum
ekfDs6i/yazpTzkSv3SH1bSydVRHlTl4S2iVfuG9Trc/NemP95W0xrTCf+ym7TDE
DWWtai3AlDiTfe1w1FX9xWTOM7t16RSXZIZS5Xf9GRUv2mQQv6rceqepJeoPFBjs
sF1diMGIL9qiSmJF+/70eVsPMCI/1RT4Yfp0LlMxaiKjMCAIKoyFDahsmmjafF5H
iogUM4L0EQLX4/URjDdIoPsZZiMg2nmVWQ/4O22DHVUZjd1Du7EUqu0d0OxTUP3N
0PLyeI7ZHJa4eE9fiuVZIZJoZoEA9Le4oLKt1gxhYKS16wjY/oRkQdtyyKX7Mk/Z
E9r89y2SfUWLaRR3ZVTLhg667qtCWAaWnOIVe1eRpa1EeNmP+j8zdfHKH6LorRc8
QA3saxdlv82Uq9Rjqh3II8weRevjbMFY2Q1eduje5ebqjexY1UqmnQy1hTDnBRRs
hZVyzH7G/gJvJ0zvnjccrh8WUJf7bKWAbFEraVHUzRz4FzKajy8cIjfDc1HcBqUk
`protect END_PROTECTED
