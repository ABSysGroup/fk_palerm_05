`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8oli8q5RI7BCQUaEZPKJ6wOeJhU1Hyplmn4PdtooE8wSw7qJaCw5717sxerRO9om
Z2UPHliJ29FmLHMpo655xyzb0IOyZ/DMpKJcUWXwyQXwFk4ntqnYyD/icGqmqMvT
+a7AOgChdRrqb1R7vCZEyCqMYgeKekmm3ukZ9mCe8CzDZ+YYlgg3/9iBVAFWD1B8
j30QBWIHNtthfyKzMu27KseSslS8V5JUBFhIQa466q+5AYe1ZlE4U36TX1YTNicX
Tu9q9qtVdAUBDcTx05uS6l2ukRAAbmFmaVE8AcdVEqyxNhCU/PqoC7I9WwaixTXz
AfnxThU5ibwAL2k8HPK+cTQRPQU4wTcdWpQ/8kthGyrxV7SLBhCFI9wt/hFWCk9A
sBC+WuYkV4ThpASre2sxJEkRdJzJkvOHi/tEuQRyF36uci/KB3bRb2DmJ7ZW8imW
MqARcQ5qRiu9NcWRyK9GrT+fnd9ZckE0f4emYcaHLlwDjl5Knizeu8nFUKN2mCmn
OiHYaj0VHwVfHu/6TOhkuMa7zGvjfWRVdkfHDoi/G3fEKymMAlbsJBfHP2N5YyBw
ph+V19KKvlf4NGKNHReJ/Gqmk9XvfPgpsxMIhv01zkgF7ZJOC/K+bGsEu1BmILZy
fUj08JfPYMvahpNLeFH6QA==
`protect END_PROTECTED
