`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zrrfsgoRglj0C9TjcBbv0YnWD2s6xf0cIG/b4gAnctL75ieZJXF7ouWqh6G2y7Fa
KVwLTAY8J0dEU4qjzKscSHgvK/6PEvqknbAZ1JabvquPzPF/TW2ZPqPvTnhhoLQ5
uY3AahfIXFv/eM1+NBSrEAgSRe/3dYpOmAVnEQFcQOrQw74zeY+krZHS0MIuX+WE
YEaFc+kMXNbwVIe0N0YIdyNeo9jTUdq+kU5rat8aQUzm4WOyOcBpfhv1fX5NA+XI
93BMp/qvVL3njmU2QV7EXt95K3P9fRmg4lyA/zGKB4eNeXMJ4i/88gQvzz9tFfqv
azN7izLpO49a77MUnQVvNQNyf9nxj2c3+KyCwoURg5PaMNUa3BasvLqpYr9/N2Ss
b+rkkihKledoc+l4DXL+Y/PXeTeq8guiuYayOZoF8N4mQlV+gflHSV+ZTgj97/1s
/bB0u/lU1IHTswykrAAFnFqFCb9SbtmvqjyKjvMxa3/EZT//MtyjVRyzZmZTG/nR
J7VlGxvHJ81SnqDyRm0Gx4yHIdO8vJ3eH0jUvwyfswmWudYVknvTscMA4fzw7uf9
T1+DUip6T9v1k/7iXw9B29lI6vSYQ5oI2OtdZZaojMECLp8k3sicZJDITWJxPRzV
RYmVnmwwQj/qopgkrOyqYVGe3m7S79UB1dqwUrjEIflPQEJImADj1Xx1fs9pLkL3
JRiQE8K0O+QqAuCPR9UXADMZXNIBB0nCXgd6Q5JS2GxC0tLRJ+1zdp6JgG3luB75
zpGBrPb1DXazNn4B3VPSeR+v0en1dvfQqDORIBtVQ5GTLu/jyQkBjIDocsRxinb/
ek8SPXzXRrktif5F7yh7cg==
`protect END_PROTECTED
