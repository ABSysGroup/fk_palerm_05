`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ehsbHdzH7LuLYmYBAjULmG1sEMIs/g5QAJ3UZLo7Pl5AidEB5gExLymmUjdd8lgb
Ydum73vC6JAykTsP7Wjr71S27+QEqEZRPaPx+hZnCB5URiwbqvMztINpCe28ZARu
G6Qi06+97yfyXzKeWqPm7Wusw1H/cQbdflOKxcPA4eF5jEdvyOJynJFijjvHQ1ku
eb7M7n5bTjg/wmGbddl58Vs8grdAqwFqBaQngQrlVonBQNxuI09xcRIZdlxW9lVS
7QPJ/qRl1wsrQb0+3jTgWxU+VTR7O7dClKVev4BoAWBqPvh0juSCF5gKVYlcvmJC
RjPTqZ5i2ta2tt+ds7TVZWIbMR5ORf3H7NHl8IARqYbrQPUNaTGvahq1I/iGH8SA
a/iIhjT2raDGakXwjUHq3GakS/LxarU8GP2XuSoBUhZ5iQPquYjCgLEQDNjqb5U5
NjH+Zkw6h4C2Bm1x6k0rDqWiConEpcVZNPeJo3CB5ZSNYg1bf9a4ZW0L0JUiq9my
PpGzw/yihoqizVHTav9kMiybsvW6i7zTg/8Xq4EKum/t4cWA7ZcRy0UZOBUzTcfg
mQsXqPlJSgLGdWtOKMYC0RUwMKghzvMHgIvLcKg9vM9vwjl6qe8GNOjvNlyfF1SA
iczEw+q0vIPGgGhfnIFy89tTX+Ly8ilmvxnXuPj8hbzJulWpJptv4xb2ogpsZtr9
kF89jNuuQc/vK4TRlvMrL31yK+JPhuPDgMOw8ayJrqb779hqMtx8olY4p0kk2nar
N8OYP5KbTscD/J7tnobUBrEjeOLxosGD4nFOKyGMiC7mrHYBYC3jrHRykrtNR6zq
nYyKqsvL8sZZgc9PSFtn99XPD6fe/2gIsg34fe+WBRh2hvjoAuMdS16kdjN/m0gu
flAwlY6sVD4h/sebxYG3e9OF4MR5DeAFWj4nJxmLRvh6msoCcuIsL4/8Hm3cS7F7
JPK8QSRVK3tiPMcixd8qmt5JCmfGNt4IYpYi3WKah0cLLIr0p6CqmS0MfrliWd72
jvwgMGmv+o4/VNdH4zv7jw==
`protect END_PROTECTED
