`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Ra1Yuk3aqfcxjXee+nsNP2D6YEpiT3z9THuVd+WVswxtwtGOC+3PFi20/fZuttt
CrP1WZC22ZYWE+lCJuvqxMhdPWWfxb3AL8O9j4uE8gf7CozfPuI2dRTPhZtlFlgK
zBGAi1ksIkrhVGVn+6m8rivMKta3W/nsBLa7Msrr4iIILrRgVUABmhN+Gn2K5NT7
V2bdyJXKcBW8Za+kLc33gvcH0lBZfChIfk8i4EhwH09ej07EFR+vJO4PlZGm0duS
Er2sk89/ZEBKl5Vnd+sUFs8LYHRQGm7MttQlYKsC3LZA2EkmfT+k9qWFWUUhmQWB
2tN8Ie69SQa/Aw5sJ6NGJ+LfqsHQYaUmQj6UPkfbrGyqqgk7uIuNTRUGeLq6+888
BsltgyxsML1I5PNbQnAZzfjSgTmb3SzxrhEOKjHEve9sJhpKIK/leQHZDL0idlYA
Rm/A74PTZs51vRfFFUVd2PdgwuP1HrQ1Qwcwir3O19qVY0gc4EPQ6or1p3Td1JYM
Tc4s0n9sxlDtzaKWMAdoiiDdhNkAHySwpQuNPE5g+wKkjxFc8TIz1i1seJstaj5y
qMHwSdw4IeteRoZfMaEjNo/B4mPXVuDfjbyDP24iEsX92o/+CDMXCPIG1GyEFI0w
KGuYqMKctvlWUYYIOKWb5Y36WkKq0KFdKTiiRaoca92PoFx/dREBP17oAfHuBu/X
H7mHpDW2KqXZlpUfvY5hY+PJcKZTgcPOWUyItj6pWshLS2VA998hapvP4JTFbBVa
jGGyZQXgFUHSqdCefEsSACuVjPHsfkfd7UxoVcM4UfI1iYkNXjhgFhiJhruR3HNV
c1xp48ZB+4KtuXjRgISr4pWM1QsU7CiK8+iZo0YXATKQlF49EsWoQC9hRveGm7Tt
/Qk4tEGSeiItBnaVjjaJ6ptx1TSt+7kb/ihXN5GEJ0pGqPu3P1yVm0xDsU2vRMnF
rYAt/rU1XHRwB1LyyFJTcAGbZNRhdcbCsJop/eDpSZGw+ftJUc6sb9qa7tEGKM3I
QGz/x2Q3eQCFZnSldKC/NDzKQ3AuHhmlfDcx4J15+YkFsgPIqbX33sq8FXVIDk4z
IW+YFtyTnisxL0d7JkbOuV7zBfIYRV0pWZuzaXrubnVtRLsme0him4MZ81ie02OT
LCu3/Qy+JBsod+184bv3lynEm6RBA/syjw8jHPDvp0VwbKC7hYxK2DbluryBk8A9
0Ih5rTBfKq1oH2Rc5R/9576GEC0QSLC8WGXS1eGOb7fzbWOvi6tCRsaKyXz95Zrp
+R+l9oXGlO0I8Lb488apY9yjwlu8+I3NhFcbyehwLbMHAQoy+Re9vbBxVHXwbfqi
7B8u167uPb6OQhT2v4bcs0RK2tuFqngEtJFYwQSOkLeCso75eoUTxLYNDZaW6FV1
ZDcPz6xXGXOoNwdNi3wash4PjMGBR6BL6LJllQx9yD3lh+DwvEYW44JvqExZBmQR
G+Tb7UhC+8Ix4whpumfGHU/ytVPnL28/dpEZUdVT6DrzFT/5DF76YBZGBxQYUyv4
re9SsEdysyjuItCRqFhz5aKvoOj9UWkBc0PqDiAGc3U=
`protect END_PROTECTED
