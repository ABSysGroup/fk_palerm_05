`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lqV73DYzxTfPMGQOr7aabbESEDkP4qWrBpTqEXSv1HxFXEnBGaAanSskJp3vA+yz
FunrEl6yRm38Fy5McUbZJpVvBxFFtnle++DJ14YWr4vKIzDk9ZYshOC5oLQJZf8b
r32z0ebwAW1t9aEnYiswdCN/r8bs/pwnWfAbvm088+q+aGOCqvkaoB0GAyT5TkO9
TDLLabzyDZ3+bVlSDYh+CQD+OD71OB/seKZgHac9Mk514IUylQzHr9adxjnjvtQU
`protect END_PROTECTED
