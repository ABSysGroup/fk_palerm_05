`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xAJpGtlu0JEfyV+Iz8vNktrlTQhnVH8xIGBMW9gWuKwQWhR3PAHxZBPVFg9WdaYy
8uinUPY16QvGoPjdGp93zZfxfGzLE0HKIzpXM/UnQtAclMzCftshum6texMa30pX
XzDZzYBW+cgvnE0vG/wiDj3+8DgJL8eZZByWsN3v+m8hwlW8kxCFVWRWxMySOXz5
3QbXJl9TljzVr0H9kMwDVg88B13392DfRsW3LF/WcQoATpd/pvD7LReRnUe/Tonl
ikw9gM109Gw8RJQy6RdlGSdYLWoIrjHcDYjJNYT8e30IPHl/B+QSMm5qTSATEGuY
hNC3k2n++aFoI/g/LCiOsARmiqc4saJSqq2uDzCMQ+OCnL5TnsMF9F+cJoawQYdX
Kx0O3Ss86tGXeGeINCKQDNPUtqrMZ2x9QEkWz2mN0oPPE+6zXLEsPAbApQeQ54Zj
Qc5fO9+ewpgY8tIaVLvqj2R5HVIgpdSnjvY3A4pU4EZSEuEZJNuB2TPmK1ExRKfp
1/0ou54JsHjUh64msU3Q5fexyGQUd1TgwW2bUpoxkzFEOdBPIb0ksfVEdqMwYdnx
HAU40KcEAikCrqqX4CewNKv+f8U4+UAeimeUYhcfipbeesHYMa3Ehmmy1fBa+pDu
g3v4vUBEihVFTbukJoCJyMJG4YV3CyLZZTgwJzkmBAHDMFMndl7/bS3j6Ln4Sbby
RUsmXm4YtTp1wN7kFQNyeJsMgyuyyDEHWyQB7slYT9jLP00Z7JqV9fJzn/cwupto
cFOoTqh170yiJuxGHey4/FxUwbrkjUEMFH/G2jFL0ojJifMiFFZVTnJHhLN1La91
GLd7Pe6CUFE/jIdlyu0/KgvlYzgTrAIwwxmWwaHFuVD/RVvsLXMXe4SpFlys+cU3
8f3yjy4xvlBgRDHgQVs8HxDbFDjtQlAsmLfrTK7psQKN+RTLwM4JTGPBz2yq4+3s
`protect END_PROTECTED
