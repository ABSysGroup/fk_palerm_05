`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VmFEP6ky5q68DQAVoeFuYB0gLigY7DwmXoBT/GdYOZFHmQacmU2Co1coUhCOWC4q
s9NtPM74p3ziYlCi7mY6OTDWS0p8AvDev07S18/Dizw1V+QsLaLKQZOW8fszL2+C
YLrcRjmumXIcmzY2i53HzsQErdH8D5bFhh7HEnWqThmP5JdaM5zaWTe+5+/mPPnY
aK9jg48Xso2kBD5HbP36KD5OSDpkce+leePB2Gh4WHWFBNlWCMoGVpUAOFhju5tP
nVwpP0stitdl1FXsTrePVk+qnMKvZaMmYWwWHSGSs2DJaPC5cWB/XWOav89peg4R
1MxzTEW3+Zn+xQNJMavSLB6P3rPwY4qx/xAcRztBCPmT8APl86v+huqMU6NRRxu7
xD3NVzj4rhFhgrF6cirna+mS7gI3K2wCW9LxosGFy3UT9Owp8U9REt8vcMd3iAog
cv+XTHvYKIWNM454mH9bP+RlqlqhgEpgNpCk6zEMy1WLXo2qnqb2u/JCPOpAZ8y/
NtvpDvaq/StTOnlitUewkKuG1aCNfbEio4mHtNt8BCu3vzylJN8wKeI06RM16FQf
l9kt9YMF8OTYaFuZXF77W/8ZusuZ0WwNuEIcS+be8E2v6HWspLorEjAEI6HOEpN6
fUql8jS5Y0PSvd51Lgt48nsBQ2VaII4yAVb3Vj4d6k9Y27ARsh9ekggt4NC1SgbF
o1JHM8OaK6obx47I6/MH3i4oGY0DX6qzMnJQZF5g/AeoRSi5MUDWSS71/nKLJA9B
+FMW4tH9/NhHHg7lxN3bHxoODmKL6zBAwtm4PSR2z92BqXpoz7zLtxKGI4oiPp7k
LaXfgtNy5aiZ79CwNlOJNBQz04jrdcVSDBJDfEtUfhbnqFGUlsAD6DvjRixYfblz
oxovKizr1dsnnE3q8Eg0p68aYAxxVxAb9GcPLLA5o64O7z+01SilYHPF/t4S+n+t
enZ7kMipg15BllHUfz9ICbJPE3uY7DiI2bhcpeFtvnNj25NP3ZgthempRIZ4JhPI
a/sR7h1iytLqXUokKUSCTjsxM42cPbF3pYlMI2ZEKrSy0/u2CNVThveOCxiSm2Kb
YriOov27kdIUrHfAN+KmhAO+u8htvu/xzDGZMiBbKxV8xgTy3HSUky0PlZyGsQ80
qwjCy1QYFhVQM1JAlr/LnJWQvB2mvXZVhUmx4alHYVcxaZ58TB/wUP3jFL6ZmGn6
p1lMehuxdncwRZHb9Dt0HmPp+rA3iZEPo/nu4fgTfpFCwLJv0v3gaqHDl6vcq92O
uCRO6vpsLK9HVDVseLRUTio8IxeEe3ZsyWkMJY4Zb3T0ZVFPVqp1UcXn59T6uQ+q
Nq9fFGxgw4nxxyb1X3JUgHE2LESxolyRBxjeJLaDgnxnhnDW3I7VkzCCvS7O+L15
Krc2mEiNwU/60FwafqxjopPt9/jDoSU1pS7AoJ+Ur/9gHN0cVusYyTIqOFK+Iq72
xlhxZ5eGmb4xmwxlRHuIGN1pBi618j4IJJx5zv6j+mRjZELq6vsfA9yBpZSkUuHV
sDRHSfXkgFhdgQo+95/4HOvTYujqz0U4CHWOb+rMSdu5t4jest3GwydETClXXwa7
X4zstmloMOhRhDM5g68Ofi6ptMNyTA+wMAxrMNXf7gVVrFhaxjD4uQ01ATWb4Ugm
0sCzRxoT9I9ZjLaUiwWhKDoohTzlfYWsR8MrkoIDzLPpsbd1suurFJLqbXwJLutI
LgNBuFiYMn1vDzkqArJk2t4XhGi13Ozn0y18RUcadRHMjt5vo4IJN3PVwDUaE5Ve
YyU4GIuFWw4Gb3fIN4RVEdrNMpFd7JMCrTKN5lyHUeVHrydZdH9qibmIb/P7JVuR
NNzuR6d8uBvkn+xUC4T0lPIo8knASOfSP872q0VjXhE2SGKy9EHxQAm+msxCnJg6
9R3s/tvKaddPqRyJaEQTXT6o0cCSVJcbb64GD2lBAfX45xnrryuxXi1BGASelfqn
neeZC9PBiuwIfXw4kqLftF/wz3WSj5rO3+/x+d2vty00kyTlfHsL1E/t5QXLrAWF
goG8Z8EBJnG1jngSAnpb+50nayZn8L66eQP9ahfLPa/3Cw9PWSVK7MOQXCwabMAy
eMA1KoeY/c9mGsREsFpKgPjSX8uZuBmBAIJVwIXH53QzuKfXvH9Lfcgqay8EE09w
vNFkpdXOqLJSTA1xRb1oi9tm+Jh1IiGZ0Bur+7S2S8fUUrEqHBWwBUE8x2qrI+hX
J+KggtyTGBJnNISmtSsr3pSllFdMn4jLU9DlTzVsqImK1Jfx7DW2Pml4Zaqw6HnU
yBWrd981WKioQDMBMX3oeUgWy1/WSW+Pf0nZJIq11VfJX10HuEOPTzpceVK9MS7Q
XC6kCcTeeuat8IH+Ia8vQSR3jq512HaHOivypIjcosNztwx/45/Vw0BzoSQlZos/
ZkGOFPnTk8BpiOqenhEKpn8dhFTx3/69CCD8nCpzRuoxWxZ5DmBFrdyNOYhLDL8s
LgL/vzo2CgDIKxjO+n7lgGcEviXaWUUg9kejpGtANOnnzFXjxbu8V7+8sHCnEe6w
Zl+5xsOjoZD3NXN7sLdHbk+7w/4I90s1fDhKGQiW9gnGBAndv80XUy/uIY5im1CK
7LXg3n09msWL1jNyR/hH+Xh3RosP50QfSIWuITGFruxevekKqLrwF1GetmKTy8tI
GtTyo0NcpI4e83iA7o0X6xuT0Zr3iL7OO6+sbYv1vgWu6R2jo9j5wjQcGRENpReH
K1QdRluxABpKLxeiyCQ8coE9rgjzJKlwFSlYSwbPsPppJko7FbabqVvdekBABMJZ
UVOhqRB3uHFVG93xVlE3Wt/roWdW/EjYf6jXSzcwf1PIPVlR9Yjtn7OgD5eM1rcW
wRU4W2p+ZMHcGVDgrlw+eDkrOh4iC/Y4emzS6XTwP4mimVnQUJHW+HLKJQYinyl+
2+eCb1KhDrX3LVU3Wc0MMG/XxKAn7btEw/s/eAgJ/eVsAnIZC9+RKgpOig5p0X9u
QhmYI86ueMK0gAk6MjDsQUuw1m+R35/an/UWiIwFSwwQcvo85vfRvGmZL9LhlEaL
RyJB7W3rWZxWcCANjQlerJLuS/rP6IrWX0opSqRlBoY5yYwM6X9uSv9FNMYERjVW
viYRscLHmu+9eajqahHIEn1JD1l7xGjwiDwHmDxXq5L00AZ+9VQOsQaqtHbGgOae
DQYsmJKgj3fZQlXzjqaDkr7IGfFA6TTjEh9iCdsdAx4fDRILjhz69/K1TSafdHfA
6usnzudfz44AOYiDIXW/e5WGO/4uDEYgkqmrhQjtuAb+EBU+RVBUuDRt9MrPtH+0
53L62eiuJbPQ8C3OBPnpXZn5K7ySMZWflXZgwLlovaMmoVBhn3zkAQ6h9+XhVyKW
sp7SPArhosvQVYC78o9mCsdakfQXGaTGH4kZHZJeZWc=
`protect END_PROTECTED
