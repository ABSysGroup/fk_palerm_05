`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gPSJx6Urp/trM6SatNqy9d0+Zm0zlRpRpWNiYRSkQU4iHl5Mep9vOsDMBHmFyCIG
Pt/Qeubk2JihBaGki3LLJ2htu2PHrcaCa9hAGxT6+zwNOn49vR2G6kOZXAK/H0u4
hvOfz1jKFXoVgmIYfMEuDlkhk5NZcu0DexZtuqSUl4P8kI1hQJdT3AykzyCwQ5OY
4STsyBk7MURkzKGU4vK6HNFxqDyMatvYyLHF3M2xB+Hn27DVeMCIBBOjeeaqFa4R
9CMlBdjd7OaIGIZKRuz2C/GCfT+8CYbgzhaSRJtBJOloyG6KpKkpFtVdK4Q7okXY
Kgkt5jk2ZgLBFawIzmSphrOQ4WKonXx+O2oc+d66wHHdI8aF0xMsp48A5t9E8KP/
PyywrQaF918dbq6j5fyTNpxkkT55bCz73ZjNDCH7YyNKMYG8pLeE8En7iftH+Kst
ZG38BbfnfhTwmgmKB7j7/fiuzOINnTnmQ9XuxJaj22hTFEzac1HPzErqg5y2wYt/
ZhP2DrXjYLi0L7xJXAmh4V+fLtv752lo3LMv/sL19M7L8nyPZiTdSHY805sLe2FH
DMRo33Q2b6O2oF4IMhonVXYiplSPxcmj3ML4CGSTrAWwjXts7B054yatEDCLk70b
RlrcgtHWTB2MI35Yv7IPGw==
`protect END_PROTECTED
