`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EYvcXUVhci0w4LHw6fEePWQmAcSb/uDgs5YpItljy/sE6q9rjKFZcMw/rr+5Dq3r
bWIgs+KdmrAyGTRMOBg9wVd7nnvGZ7i90lBTDJwT3dl15c/yuVTF1o55lC0GUP6R
BhPvWTh383iPnBaMC+mBvZzR9ljHrSB03NDMTwSWkhb+2GUseTGk6m3lTDhWOOAt
AfOtqU2mER/IIjAwhJSCHlUpezYQc62U5+rUa8Tt9oOy2d2fT+k/KddIz2RcpKQ7
CO2lPGDnvINlbGKld8967zrvLuZ3T2ds68DHmn7p9WnyKPNZZEOOSDZr9mayAI8E
qitJQqGVusjOXz2qCIFixbW04Ca1KBIotK19aPuu1UftRpdlaByfvgauS9GY79Mn
0jVguZ6hT2PCZC1tJCnGYXv6OCaHuYiXQRljTONsMfnDdu/1NL9XcNGkqKLB0ip8
hietU5nbdfOwXB1tlq4FOAo7S9kkDXEUPur2+XKLJr0=
`protect END_PROTECTED
