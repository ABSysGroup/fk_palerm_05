`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yu2Tv6W3NZB220NdspAF69qLc2pzDBmHLT/Wd1rRCy7VFAr3zQWa5r6tLbO7EOeO
NEcidtPZbUu20et7F3xqu3b8XjCN0x0S9zdBYZAhRHQNOfKlS3EfAG38JNrbrqy1
fb1xfAf0ZBPQFDvz1/SzaCpe+WvqfGWtKWgZB2jJ/a9mXMZE/FiqqeNgXq7yW+ZE
K8wlIJFdNbc6rRCyQ+06tfemR4fvu2NzJn+syajX3h841I2LV+Ahds5qErTJZcHX
jFtzzCOXytWrg4JEKaVx9CF+P2g/07n2G9GQ+O7+Aefdc34BafMXNvGu5pDIFEmW
emknL9zB2WuIDq0MBdJKdO0ocWvZUNTGig99kxZ5RPFFBX/gxv+XEwjoV7hGkfIZ
Zr5X6mc7UWLbRx21S8mO1z8QDiSW5UMGCHbQeBXT9FSwVrV3moF2IB/rqL23iyB8
wC6cjBfn/TakhUxeFrYgLqQeEj0U47Dlh6y0w3wAupTvSzj2hzuHAHZyykQ6dLEE
`protect END_PROTECTED
