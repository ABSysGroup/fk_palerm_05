`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
voYM7nZ2E0myeskXYDDNJpYDiXI5g6vUdJ7qULLsVMWBn4Tcx2PLgqHfAqLeyCqw
3LAftk1OObnJbsAdQp6QIh1OR45z+KoTtyQ83gml6l5h2VWsIiC5Ijsb/8oCy7fc
jcni4VqucC2m1p1cGx1R+EVdokXzYXQFaKifyliUAw1NyEUzwUWZau34gZ5k81mk
/0MMHwRlyjIzaJWLBitc3OzMoEzPc+CQkOXM33Wb2iO+xQco79ErIuWa+7frL/S8
tE/EiFbZ9hzQydiS3PcQt5IwVH5l2dOYgchXnngvhuNqoRBeyigF6wLb3ryWT/ZZ
t7Y22e3aKSulYNsVpdNX+wjaIGUkdFOj5cyLD/1EAc4W27XFHXa6AOOIDR5zGAOt
x1cB6uS0vz9W9yKzPFgHKd7YOg3ondDtg5q7KJrCAsM50dgIkt+MUoQkeU/SfeVT
vT1hJXE4trDOxy32DQ/rwODX7qUySLC6w/JltVTl9xyE/PaaVQgVvGj+pbKHi0iD
1PtK1ocNgTrlLxudtP7PHwDKyqnWw6j0g2dKGiszWiZOl1ZAZ3QVSAcjlG+IQVAq
8RMWI7cj3mPlQ0Cjey2IZR6N9SGk/xTSXooUtdYigmKOHEMUDMrRgeULJ5pOAkqL
wdGzbTuitqSgtIlootJMIIlAkBVLVTWOLXH4Y5269up/aHNbbrF1Z4owILvP168v
mVrNz83fpejHg6HUDKYRxXP2OuyF86DNipIVEQOELoonVd7aVwCRY6dxK1GbmQLq
gptmW39Z/Yb3XVIb9n09ihWuhY6Th5gPsxrirwVlq0hqJigZZVf+zPN8bwzxVmTH
pUAalKsIUOPMI68+zYAWDcmWnCzwD79//2cRxiaa2NkXKIseWoSnAB3X/1mfamMV
0PKHeTboJblmLh8Fw4Rg+3iGrZVHO/8goIQGzasHzCJabullWLoY77vLbASogalT
VqyUPkJjkoH2rUg/mBQjX8IyBNQ/QAyHi2FdcdCn6mR6bGzcbkuFwjYVvfqVqF5d
toeb8C/qpzhoVynymBUbaWGJ+YNEAi97L/B846eKO1jQ9PJRtdaihcl8ei2aVFiO
h3jTOIC34LA1JYU3ANt546rN5AUDV3M9Jx9RcA/dqXdj1GkKa9/qvGoUnTkfOQCu
z6rt1WysVLQMOmsU31mc2QyIg1Kf8VDZA1OVxOm4VpWpl0TRanOnOeT4/dR/0Eyo
arQs/i6HbrEW93hvxy2tZYotyW9hnOaoUDK0+W5hVKH83yHuL3xDv2QRcF8ngVp9
pJ9DFw18r0azIM+jALt1nWsMrTqhhfzfqCW1wIrSw/Gdf+6ZSGVvyyYZBE8C4iZd
YoOqJ8e6D7Q9y97NdKtEdxnJD+wpQRI5gHTAa5Ai4Tgru+sIvFCkOMdpzS0BTyXb
r2HvRs2wvBxZv/wgVcTP9JNQSlqAsDOOabQBF1ErFtBqnVoB3vlGbVWmGP+PpgDU
3w7bUgKx8s3oBoShJB0r+feYUlsuWSwQ8tcIFV1/wP5PlVgA2xvmO+pEQ8UBOwIY
TBNXuk5RZOOFLSsFCIIqEb0CSJUZ1lllfJ30RszpkkYy8IiKrFXdPdxDAszI+P4H
5O23L5aKUn5WbqTd9Js43aUN+tpZX9/F+A0NcpB3i7rRG3l1ii7GcOAihm/CEHCB
eNCjyTU6eLgvRrqF7YXcbdZhoZNVZX9s4iAhyTjCczM+6zZP2UglWTgUfbIc+fBE
hIo00UEitxs7ogbJcBmX+t+TZ2V4z+T5au7i6HjfixI19WIhrUGCPy+pbj2FnQ5k
9E1wZOEGZpryPiKIQ0yU/9FOo5D9e417SPZTmxX2YHeEm5fv7FF35sBxEklBWYZs
hxxKSz7p0sHTV/WQQ25sgKYsMUHTdkqiphjUZ2KMPGlUFWdfeGbaHz9f3pQYRT1A
WL/dh/tQB8km38155VQHFV7hzATMMDD1Tagta60UIy+k9bUFqzjhktM8A03uHCEz
qyILVAdSfgpmwQWPxI+DUh0NIAzuLVFYTC315HBImTpjqg/leJ0OuBEUMzUuz0bs
OeKZo9vFfHhAXXAoQa/AHGdR5u6HTW5kCLCHzgJjQ0Uc9Ri5qQT+X97Y86TnGu/F
RqU2FpAVw44Wdj8AuqgdK7UNrinbJXcljdGlK0RPvr2SdKQkgPhi30rLvfUxXjbr
gKBMOzDoDZ7LMdJdiz6Mv0CGPy+8Hd50LFXGlSVTopLOgaVJPUChtPmiAnGW0oOC
KuzVKAbjnIa0IxElRBWXhitsJJqc6R6d+aDG3d/M0hMJiTl/9XkqY3Dn6U0NjoO6
HW/TDNVnJzxO7lXDoINllTCaweFAkrR9BeHzm+eg2MBU8QIvgUBbgDpxJstDtDWD
aKFo5/XZWmtuSZ6u849fjhNaQI4NKRugSTkzMJpDjNKps4+QP4svqqZCaPdwirqC
1s32faC6/sAPzVlelxI4iw82MIw5aWIteA/fe1Hvp73iE7WNo9fdQjYVtsMmtQvT
FCP7ty446kmbfW1xAoQtCqNHSLvkuT7FAafArRC9rZoBPJuc0/+T9klv/NoHbA5o
R2J0Xb/RpbP5wkPS4iX4RhkTOO91UWpnAReCAe0+JVG2xgIyhSCxoBeInF2Rz+2H
eiK1YCSLWS0rxizpZOhF7/jFyzjWnumMVN4gasGcvRRih49/z1o1EVz1u8HqgHob
HBR/e4uI8vC+OJ2wpaiwZ7/l7Cm3mbEGf6OCgkxwZBeie/5RbnfLQAc5X6QGLOQv
2Y8dNUpku7sARzxNijqLseciF8y9QNVUjHLaNMRIO1fUgVt1BDseVagGS8PGM1W8
DSOFriYNAR1XaHEk5ArnCopvrmVdhh52wqKXYEUqB637bApAiG/6h6i1E59BzA8y
OKUq/xVg4KtG0T1ONkHBfU2GHDxYCUHfGMtn2h6cvYt07IqfsS63YpCU1MRNAonS
k/ViBCzImKEqXv8vK2v5aQBVbDJeAs3/JV7w30x2v/Bs920QXUa/rl9WqBrAq8sa
kpfUnxKwFR3HDK5aem0J8gqhyJk4VSdhka4xk914Rx+wMlRJqpQbqW4lx4sp1y8M
`protect END_PROTECTED
