`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5DOsr3XZrQk741FQjpY7PTN/PbBBrMPN3l4K7Sp5Ng1X7bzDsip6oVfvYbvmQnEB
mBOvoo+z5vWYSp24jm+sAkT6UnsVZswUdDZWTKU44hEsBNV5v3e+eUZf+mExc7r6
cw1O/epQSXt/Ohwphso5JpT1RxKpEbARg8fT5roSOFRiLcelS4i8+mGsvL0Cv2HD
9KJDeAeDjks2kqvdkE0Wi5bArSfH/lfnM8odzCx6wr9sLO8TsFlokd3xAkbbktl0
VjyNbzFAUBJ4J8f1dpAUemJGX0UZ3pQs1AKaAUSvhCuHhvOyjbwfBd9fK/ny0k5h
mxL+Iuut3fKFvh5EtWSO9xP6n+XQmBAQq7oK+xfe5nAsinng9a8lZ/7z8e74XUUI
`protect END_PROTECTED
