`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JsVKqCyc1c0Ygnpf3imVp7W+HMynCLqssk6ancMNUulp4vv62aENgeIIdFauZQfp
ED6M1Ryikr6k7dSCI5pIhEpD6NLdcy4XOMjvYJF9MKHZeYh26MuAxx6wBzQCUnXy
jf3Zb98VO7AI9gJwifOP1gh7JC66MfrhLUZLE/okZETH4QA2c/XuW0IFUck+LF+/
4WTsUF+3Y8l6qn5NvcU7gu2P5YBbqEsyJethWiR11tjKxVnJQ/nbowpD8aCykcp1
QHj6AHnlweCxe6kBVOR6SWVAfLqvMK2x9fnDafK34xvokAVPmQ36JtgbyN6rpoUD
1mPgeYcQnYkWeiuV+l9xcFhf2CaDYkHYUYC+NNgqVQabPQj7udFQxXgXZ3o+9bQO
rSQHh7H4O1ZWTeYkA9F34KiUzQ2Fh0xJOKvVl4EzGfs=
`protect END_PROTECTED
