`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GQsEskRp9phZZS9TCplCMoiN2+yTqIgY7rpfqOL5k2Uy4PsT+RjTuOTHEzfN9xJE
2HG3VEqRH/q099bXXtrhYDXD38AW1b7Cpb/YwXE9RkQPg4RNbUhc/C3qL8kYdtby
LIsOEK+2rkbrmxHUpunZTvNCi69Alm61YzGvijh5vmAry3+mbFvhy0IRCH+Mkd8d
b9RtARaviJXctxxWZWCmEogGnWamZveyeL3Go4iw2Q1V2MdEcLCE0CpTCYcU0Hme
6jI9KdhddBSLJl5otxi0lftMMMcksYeQAjVkLCa/rcJO6MeZkte1FC5y+kMvoUMR
/151eWDkEcKyTUos8QVTQ2JbL0MifugZ1BZWSSyeqTxTAXWVR+x5vRZueYAjP59N
ZYPvoYhdiQZDyEYdZaT+9O+Jl43oXc/ZvFySKNEv0gUl5+JOX/DCIEg8Xi6l9JXP
ot87etP5rR8w0Wi2/KYT2i83JAh8pP592EDe4TH6flpDv4h2VWmQMg6XkJuELIWl
BwExKT0qd8w7+QVxVWsSharM9dsYWrcxxrGSVwKnMEUDm368uuqqZG5DHdM2Z8um
ckagtB7ajUsOXOOiW9GabEYlcBwRd5bBcqBT6tAioQ+uZfTTPr81Pek3iA4iUlGQ
d/PfMaFuSNdnYDgcoG3bNCVp09lpW+2PdJnhuEEJwzLUZVDvSSJ7B9Z+OMFFU5ME
HOtDz7/Ul1ybQ+vs4ZEM466Efj32UXwX2R8c86YdJbc=
`protect END_PROTECTED
