`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fvt3Z0wWTb9u72PtvNy8Ft1jItUQFOYGsT2lEWFZzw6Eb9lCOb1v4T56BlPeohgZ
/VNs9DTf9WS4MKyeWCwQj4yTb8ilra21SGVS8QsIXaX0lCql8dMJVVQGUXoLjC77
yx+HulY3NAXffBjVN7CnzfZuLrBP6z1i5FfHASBKL1kXRZOwht4zEhDRFTGeGGrq
CIis0sXgc/Bp/3aMKJiZcKwOl8eZnWn6wuo1VnLDXFUCODwjUhLN7cbhEngb8X1M
Zts8dwEnBR7/JxpS3kNUdUcGwVQEvUbaZcuYs0K6ohAXoF911lRUXD3OnWw0sNLp
HrpaDKj/uJgWX1gLWTdd/cN1WXscxDQord1shPMoSoOH3HqVfYzmwW/FRzOAJGVF
N9k7xgNjwoaPXW4HnB7w8a9RSSU225Kd5cDA5c9q/lfnnS+jDkaa965TiiTDRoo3
yBjj2qvLlDBqYPx/6IjzzIs4S1QcdBtchghEk0DfI3LVN9+4ABurzx3z0q3612Ud
`protect END_PROTECTED
