`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ETzAzHEBniqRXlAqXfaqTh1MU/+LY4ghRAp1W4AR4ZaSi2DezskdGWrCMGUQyXUH
8bxYGg+nArYq08E/NrYO+gIgooGPy5hPw+ClTnw/01z723qDRbbU81ZU2n2Vha9d
AN+gDJRKIqgqGtSa/BJg737h1RSk0966xF+4tjNj1tZRP3eyZGIUs6Sl3NRMN7Z9
UliLf+LAtceHKCBBcvlbSJBievh7Qplaii4JpllSlPwWGu979h4eWBB+JAHR2LaE
18QCYUQV+9l30bYs5VTxv0V2SdF12cpcw5s16Q4v3b7L7AR53+n5L6czHZrMXNI+
aPfB/d227NU7XhnPqWvaioZ22ITOt3rvpElwHY1sXge+ddOFXfRPD+77gFJKWtO8
UKjlIHfMi0O0NeO9wCuI9cWHOobwNgtNKopIPvmJzI6xiVBLoK5XUglGNQYxvJFA
qgTqWuKVqvtHs2uTK82kmulZhjVIG542KTxX+BiF6LnVOkthpq1OD2ib+kmgsYbR
HJvNy6JT9AEEJwS02kh3IATZDMzsYBfxPHMgt3xbI/p88AJ5/hzi2mkwue6TEF+J
5vowoo5R3k8sq8cNmvyNlP8PSA3oqpI3GLtDhb+nOTsMIZlR9aTp6A5myPdHoq73
WKy/32CP4NKXY/dUYx4yDTEaS2uWow0vdSw9mbfSdvhH93kLMZCQi10nKNIMYZ1X
MtumldGSJmBjcAoOh2XkJKeByDkhsBBzn/AWnR6uowx2Oci+LX0rGc9Tod1gUG4T
BtCmpElFS5WdDZZMmVhGIQ9YywgmeXF5FyH+thKrqjvKWE8ku/jKwEHtZU1bFs23
LCYPDIBgWLGe1fHSfkCFPywwRjPYaK9fvmRJb7TUocvVM8BC16kCS1d1huxip7xN
KgPC03WIcCtom6IBs73I8gXiBzrktrfqYO/MssZhhWRJcavWNdmEB18ujEuskvxT
H5rqeOlaBKYD3UZox3+X91hEixhMPmdDamGcvp9f9aJNq+bAuNWWgBdQtGMyk4B/
kAVavGggmCJsP/e8XeHDxhnpodXMk6PkiuSSkAYQDdHhdbUlUmAb7VUwc5RG+oxS
PS7LuHgv4CWOU1w9XudbOa0Lygu1ASLwHKo7c3fCYSjIEVs9rdN5xctfi/l8FvI+
Ev0hf/5N3/HqWH0UPGDU3rFTv++KfFaeDk9tR8qMJ1l/cb/0rVPIx7AC2QpvmiKN
+E5lNhagaqCfe/8eHJzn5BOIPwoAeT8cNsstDFlJTFW2D5OnEoDaJOhXe2KOMYSd
GXaeSYHpC99WeVLXX5zXcRXCzFKhTtdNlXTJtNEtAKduBgrRjOMlphCjCaIc+83q
ItJWIfupK1/PO8lzpvJAPoz+4XMUNFc1SjFQC8SYneMLr3Vg1XPllG9D3POSvV8i
UDJrT5GGVJ2R6cV3yjjXFjOWhDEsGK6BjtRY0GAzmKrQaWVin/cPWefJ5n8Qy4jx
xj0di2dN5mVWQdvoB/5slC1KyDJ7986TiH7vZv7zJHpVJdBkQTqMztKBYOuXPc5e
8s9K4qpApUBZAI0a8WbzfTLC9jWuUqrTO/wKqwQSXSwOKw5NhQR+AXY/wd7Rlx5i
okO5Ys0a3TKMsoCDddkC8LTRa+23Pysk9zrxBWZJwbRy8UCWmNxhujNlEeIIQ/IX
hdybrz7niGApZ6w2AJSpdojFkPotdFeFVu3yPoxoWqzTfKbpDt4ALYWQG1QmLh8G
Fta3TS6MaMe1tNuQy7kN7ka7Ja3BcwjUc1zP8v0D+v+5ZnbojKZcxqTXM82cMyWs
2PVHBrToLPZWhttNtVMI9pE4H8DBCfJ4Tm+4tA4qP5651EP9RfqHZDq7Z6fQ/mUv
UXHflJBDtiR5WeRWhO7F8+E6NAbXtg0FavwPyVp6y/O9G8Fg+m1IDuLLS6CZgBp3
Pw6jc1f8mM5pluY2tknLUhHiufDBx+znAcBkNLlQGMtOK6oEhtZY6MFVIh12a75Q
Vy41h57czJIHL34tRD5+okG5dUSQJIOMg5ve5JgqDUOfL76VufucrbhCU+9JGJ1A
jFjvyFZ/v+0u8aR4qrTmg3EqWTPjOPZD40FqAh20u18/HW2MMMs1kR/EDz9//cSx
x7Ul7PdU9kG0ewc1hARKsS5I4WpWEJJs7FUpeM+oXU5Z7L3oaJbWcD9B92cKC30C
xeSut/kD2OpAaHlRwLSQKFkUA2301nsdH/S8fE54FPedrYn6JKg+THQjHF16zjTh
djx9S8ogFZpLok9CdasNNUe5kRrzjhN1WC1VherhWFICrhriCM1Y5v+JcDFzuBJe
v4l5sYtrgcKZWWuFWykpY+fwjDM8tq1oVJ3nXGjn7/Hmm3SIOEwiCEE1GXhmwAv9
M4RGGXgH5wDGzrhRNvFQipS6qrGDt7Xh0iAjUumSYokZ56H3pAD9FF/bU/DBAXjT
reAh0mMEPa5UrfQyRzEbOib33djhERRbC9zwEu/yQE6TDLfUv63CkGsZuSYNFhfi
542yiMUYciir1oYc7V5keeeQq8MqHt8CFaVV15Bstutxm7f1rLxRT0KHZWAZbIIn
uHxjQs7hMnuBwblnUPbpyFP+hh/TG6fz/C4IsLd7BHiW54vR/SFveaLFDw7eRK6E
dZuZdF3CzigdXhV7KDFFdcCsgQB3+dG4OEZXiM13JkfphwUDxQmYdEJAEOLRRlEi
qG+tEkpKel9wuiWbh7oqamGXAHo6ura/oeZHYkBmwacdPccwREpaxVuDAJBEtSPj
XfLfua7THJEAnJr4BjYpSdvo/QEvnFI41xcO1391DdRdjDWE+FTIFDkKeDBb6Cf0
lbtJDvg0yl6AaKRlZTCc8sUBlhC5MNZpKPwJON2uw33AA0DZGURPTsPwe0HvGmUo
2ropVk63IsIiLmPjcgkHop7Cem/+rSP30KqY9J4rm9pHDHTHRLZj6Vz3HPEOhX0F
QdCyg2QdjcZJuf6TQJQppZkZnYacV6rMQT9NliErtR8VLFXGmKu6qNGeVJXC3ymX
GsSDns8oLjmLKgeyveE3NZEPoXzrkDMyeGkJWdCcS17kUHV3ieYKBFcgj+WINYji
TFks4nMiDX52APlYlx0SA9SAhkFxqrQKtQE/4JeVmxfupVP7pt0uNxb55WB4UaJ3
4ps9By54UO6m8hNRfsYqbX6umvQJjElLE9lWrLsjVHtKgMNxZHuPvtRq/3YxEpe0
bmObYBbYoz7SydCwKsvJ+faIrqYj7q98THr0fTDmNSgXNzn69e1gERqExu4bn/Ci
O1Oz2RtsZ867Wtya+voRYHXhWKy8fBzaXDNZqIKJryVcb59OrTckFe7y0YFj5rJ6
Qtv1t4CzXmq2Sccz3cxrV0pZ5uDDFLAzo2440E0o4enzcH1I16+hJ0Ub9AlMhem6
xYfbb4t/6BFvTUvzf0Q300rgR3lUhe2OCI+fQhRUtVd0RRfSTpGxMnUC8mJ9Pdk+
HgqBPVDDQ0zHGRSsvgsPg6Iiv2lVFEYzKqaFLnLx0/Nn7VlFQVvEH48YRwWfS67M
yFFJNYp5PcRlbIyPMRI19+SP+4FuneXYibeGI/yGulRqp9+16SFKe4dt/w4chQSr
T2wtysBmnq6BfrOl8MzGSjw4kfFQ+ZFib63yhe7KX/fiZhRH15m5efQaqNzoPfPB
o1w3p7P5huI7Mp7a6XHha1aMHLB43u6wACVaoteM5kO2DuqeXdke16JiKiMlLTPe
eVrhDw6wbKsL/zloWuW4BnvW31NKZtkMHKqa6zjTI99VsoloORWwhgEhR/3p88nF
ssy25svyltgDUhoxFeaa0uEkQu40UhMG7226uJMko2xcv6ryH6JnJkeISpWIT9Y7
GgAUTJ9zU6n/t8y1ilLi+NQ9v5gDWqp2mFmPubcI77sxpUngsv1yPIXStx3qYIsa
LcjCtXBUO1u8CENaZAqk/Kefp7FEHT8sqov8PBpLVj3Km+kZnH6rfAtYuRCthFMH
4iDHzTlMzGCzt0j4UTMFgDVK9KTTIeUQIBnjiDwR2DaUUuetdeJpQC0e7qtCsgoH
m9e9Ie3NTM5Rnmlh1F5nQ4UNMAOrhx6kzrt+ayIJTJon/bhWl+j+q14ZZQ0YdzdQ
Glmxjxhg6kdKvxpz9gM+U05XFcFJe4O2UG5AnO013RG1E8I6RDSJmq8TFaoE/k6E
dVfXXpj2ZFkcpxOrvi1+9M84NmDiupSEvk7hekbc1zLe4YVGAcnVatU5kQbGLEa9
8QFRDmwUVeEXcCYoiJdXpUcMdX8D0d7IPTCkulv9nDc+WqY14uvan4uh6z3qnvsO
guhUhdAIj4wmxjGmembf5pQn0Obs2qdSvMVgO31UMk1SxGdiaUmNvREovidKUcKQ
jUbWI+U7GuXHOTW8DXkrOymTjYZKlX1ygWxUZRWHUcKwx8Z4PwFc5PccCtsmxvtY
6uWF20+LaOS2g80bAwIU7yjl2f/A8ANyrd0mtbUuIwuQURkpY7GXOlZLYDecWt2c
YIjhbYsUOGkOzeKHv+XQyWAhXOhtmht8pxOT4ibBZQgu1hlhP/gjbh3qZksK+Ayd
ceLRwCM4Ve/amgpj8y9Dni5KXMfEOid7dkkc7qcqE1oQOBolnY4ClZehJfUkWbRf
tTJLTdw26IUmxVpF0CyowqQ3jDKDpfPRcapBKnCZvzSKKcAyDZk7X0HXJJTf4p52
mDNU+LMC+u3oDGwd1GbT+e1zP9e0V2P/CsnscAeqDvA2BRnayi1v4Tr6uErQGgyF
iblusSd+OeIHbizprodviVqMrPlhtDu2SiWPRxoVjLo6cEYjXGt8oG3W71ccPKnr
VvPkSEKo+1vbXkLk5kn7CJhL94erp+671V8MPBLLwC75nw3KWQvDnlqr3HAqybmB
fYiCLx2wHVLtHUAY09SvjBEe1xwpQtIQsxVYEo2V5gDQGEbdxQxlYXvxw/6AYMZv
aBCwlwvAOwGTIWh0GsihfIRUcjEHC7NjAZYik/4KR+u+pK/3fQleUapZBJyhi9ZW
yjih77rWLWRgQlWq+7Cw3WI7t0d0EL2id4SV7AQOLOjv+RzGt+Ay6EI8Moql7agl
VuxMZZdh5h0b6TOKxhQ5GQoTQJmj+FGwgLw96QYsiXorNCffI6w6bfbZ64T7fnuU
fLw1mcvV4ujiTO8i/CCn5RxWg5vHT2MO7droXNSGQPN8/Epp/9viPzsG4skO94kt
frU5J20QH2WBp8LZGtWHNk1vCmFELYhNVBx25Kw6EBAKGcLu9U7+esgAaovqVco8
j1QnyJmY6igI40MwjXv8zvFErKIuqBtNvpJrQE1kP4yluAIFvbkLQUQ68QlV7gp/
Spp1PgA/e2H4nQUokUCXH8jgTst65tar1oHUPr9JJbDCFXrUK8TYcnIT6p+oydrp
zAC9N95QRFFVPrHI2cUhjn7ayCAMIfar/mSthleFdNUjhjYHkAWYYxXCH91dsRpG
yGsYznmZtL1uB9YMvaomkTAC1edKybZ4Z5zdHEjtErY8MkXoKOejaIOl4QYb3dVQ
cLTCl2z6it2H3T62B8vE6Q==
`protect END_PROTECTED
