`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wVHmnBPEoP2j13jaOastaaTddYGKWjVCJt2XK+nkVg0wPZZ9+GlQmOcNyAwGuG27
4TqKvEicUp5JfN2bKGzeMXAo4kZGVLPLgpLHlJ+3exqXz2gSZtQP/gW6G0qt2r1I
GcLB/cjUjomJsunzNx5AuJ0M2YCHvG8i9QvUfiLYCy0=
`protect END_PROTECTED
