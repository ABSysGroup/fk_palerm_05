`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6IVdSkqnVqTZxQ0evksnkV3tLdefmE9uAhHSsPMROTsDwwh1lgYGwg1IXMptBUmk
N7OICw/Op0TKYAm3pxxT7AAB9fsluZE2d5tSN3xzL0TV12ErrI0GyU1gp0f21gGC
wYak6H9f/RcIUs8lNBY0eLlQiGD7R7KBo4znbi/cVaNmtj0pqHV27FRm3z3+wadX
TtBDjcMIPvypIhKTeDiWX6H6qbQvvx89nH2XCw3DdKi27yLI27+87KTLDjdpOgwL
P1tSVJOqrJNPevQ0WP40hQ9MEUvOt5feEOXilRq0zJ5aUhD5eaTN/BfP76k528ZV
ysQgyLfTaT/75kUkRk0fYaihV7+bnZK8mQA6Q+xlsuAxKy3f5xKX++NApTZpYyAI
JNvlPH/t0GAKroP16PsbNBC4E+x52DuXVzp5KGN3jOHlcjdk9pGDwDST0rW0P3gQ
WqY1iLh3pPYQ4EHCyxUAlJdVaDQHOZKzRgG+pdW9lo/8OHdOmOWEVejIp4auxpY8
q40T/ZMOz4zhDSnUKpzzxDdECd1PZbgwe8QMYFEWu/M=
`protect END_PROTECTED
