`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aIqUD7vYjKGPdjcKg8+HdVUoUuUj7EtmRrFeYwLU5b/arLhidUrg/kNW7v6aBILL
5A9BpKjRESdrNI/iIFxXP/qJi0DGm79GApOZv7XCdHTLqGgEHyaozcHrTNGXDDzq
83PBkVKu78odbpKxGI8rGb3BGBhfEdQYQOgBCGLKVooBqTG1+hw8ppkpOYkXw1E2
gm5NOkaA41NwyARMGxQcPhqMTSscyNDR1bxyrdJlGYicLxV5CRR0S4IoHiZFptdv
pY6KsJ/i2979CZ0I7eb95o2qJ7CgojILJGFYih5FhNcjmYWk/e26rxGE1yCH32rF
MUUbG53rHquKahqly2zUS6FNM1AeMewo1/mtQ1UYImtKW8ISwpwyVq9dtnOCp000
54PP+/GWhmGy5cPIwK+LyfbzkW5Ew3vX/HQeU2fOWgjUnJ2vMSCqcFtxVHYw/tRb
JPgfgYxjNq3igq+SoLlXQQD5aC0Pny7iS6bEznxWLu1/98tdM8fVbzkQb8yRMD0k
zURb/NY6VOWWEEhflTS/pvQTgCfhvX2ENgIy16lVudnqr9hVxvyyGhF8BGbAGgiu
ylozFq5VgG6FYUXrpdvTAHoo4t++WZXNp8jGt+gHZ8kkdzLGAgUm/h5qg7pTy0Lj
UznXQot2Hu5Qa10h6X/w44uoZ1ywweACNqt6cNdr2H0=
`protect END_PROTECTED
