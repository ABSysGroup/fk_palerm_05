`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o+czmf0ZdwlW34yjEvOcXdrXPQ3qlDnHc4jFEUcBenthDtdPw+RMJF/RQ3HK+hvS
B92hsxRQeCugoReoi17hvG5zZ1z5OvKaP0/4EYyimdT9h2ZEXX5cOXzJB/3+9K2q
uE8a9+Gj+wXag0ZgwSYQu06+Sv/CDVytt9h/QtJ7CvL+H/wokdu1wQ7SkbO+ibE5
7vgQxbWp9CIO0ysA3+DKFIIMSxx91RdBqUCuQDhXaRnQqReVMFDh/wy0fxJIp8oA
OihGf8wr+Kq8mHG+R5ZpayPRVTepnWW6bUrrzdjcfnXp4ohoNcfqCOYqllJrMGVF
gwn6Lg3hAe7Uhc7ZGKLhpBbHWsKY74OtBIyKeW0YLzu5331B0PdKgpgvAqpmHPpQ
h8ypFPBYLG2tCJrOZO95EhvA/I17JkZa2bg4C/e1Pii02stKcuGogWJUu+6aYmuV
jNpM57fsF64gdlu3uKDdxWJhMDq1XesyhqkTJ5oHyc85Hyn+KwFgezi6CE8GOYOe
Y8qPiHEt92QKmy5fVE0zPs4/Ar6gmtjJGxIrVNY1q/jOv8dXZRMuUb7MpJ4tSkMT
JRU0+tpacCAe59EiEwlqGEHdp9r0IqKa2KaszibwRUTjCk9+NS9UmvCKhWqFRW+9
dO/F1jPKUWNvk+6WIDKxZS6lsCxhJ5tvSQ/njDXRkFEVb5yGylIUQYuMOUzRfXG9
0F8ZOeeohD0gZ3rvQp2NMbl9/7PO+dqgd/wicpfqL//CtMs6aWy+SnQcPMUV6Xom
NTZqPace7VD/hWdt0M6Z6oiMRo212N/32tUhTppUHmZHtFYENfX8+AIYkil3/TZX
`protect END_PROTECTED
