`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iGiD8DrBhILbRBqrsq7DI67mCcKnZfyDFWCm2JR9qXFRdzlehe3JsnX8V9XOA1ua
gmnsJ4GLBfdgph3hWT84z8Z4LHuFsiiI6YhWoEh+JWV2EaoLe2ONA1f5yiE/nyyk
2QFsWCmYyBzpowjZG76QZe4XH9oSBDDphsN/1+vMNrqHi2NJdezGWSXldNlrAlab
CStTsqh8n4swLbhpqP06JHIEi3h+iX5ijWpM6elyyCgqplMrJM/p7ceb1pa5mvG3
ePHzCAmke5GcvriJw+Z/7sgpdZZz0u9ZoXSQIgAxi4fCTMNoRCMZxq0708z4Ww2+
5RYbgryrnIq1CCf6TMD3zOtC9Fitj5UZVRt4MZ1e2IVfDrvXfykMQkWm/3OdSPcy
K64OkCWaM/LPsg+GbVnKiV8cGrRn+hyWLXE4CUxKQ7sNlGaTsgfQ9JY8qAVXGHhA
Zncf5sdCakmbltkBMEVca5Uj9I7VOu/a3z7FQYik1+3ZMFPutQ6AQBzfuztPgo2e
9DiV52u2F3zY3alDBjCPOsSFtPBRtf1MUDX/gj3kH9/Vk5/PEcK3pAbzdAtSYtil
XdUgv0mTx2zF0q6pMp2y0Em2RfWu0bHWrD0MSsQVFY7fjeYpd5s9eGax5M38hiPv
1GeN5SGPkFkK+t/TXvLDrC9Dbkp+OKFoEd9TxHqCD1I=
`protect END_PROTECTED
