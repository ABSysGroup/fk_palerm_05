`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/G7gO0sdMXS+QnJHxBT3cGdxwBZfEbmAmeW9SX0iyopM7EsJQmfzZ/ZnnAgbB583
GGlriFI7Xq+N0OXM+OVtj5vQ9S4qOaN6yiIGtTDQE6vd3A0SnwY8caId7vUCH7Wc
tO5DezNi0Kma+ddN0g2Y749pB1DQTRdEMrwrkUa7wPlaW6jm+hNkYYLNFgZACwXh
faWaSapKJxT14E8czw4rHl0ZFvRyEHRgaV66vT1obPdY5ZWst6QFFO6RGMLamYQW
GfVT/FuxuOibdLiH9mw33UqKHMbzW6WAjfZTQ0FUwZFLz3q1OchznQroad5zTkiZ
tD5eB4a3XVBE5fvnIZwo889FCJbbGffyMedtWjewVUVuJl1ZwEsDKd3wkLIl2TXI
e9DSNp82qhMToCgFljJMBwcJDVhInnK5xuuEAxocy3HLa1CT0w8SQSzj1KUsJokB
1EIxt9TExiYVMMnxdvbP6q4NHMIavsmkBXSG/OtwbEptX3C4kBZDWOp2onJ7Nkvk
`protect END_PROTECTED
