`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uPGuZT+gzei0lYChZ+epmzSBx00Q3QYCv5NY4xTmQCRq3ki9+omZTnozha2xlWhT
mIl3Qf+kjDVi8VBX+ynTYFg8aXmiAcd0amfyKEdgNFHdDOtbLIuqmPnectVjvx7s
0yvSfDoX848CD/37AGGmSxT9Z+WHJ2nfJuqEMmENzkHhrkocycUAtXKIUtumNHNY
yNs1j2McecXSzOIszvwl4CW3kwScZnq/lChIG6xHTkaclJrLhEB0uGzMTGyvxe9m
ijZ+p4tCXPvSZiUufNsnwRw1cEWQyygu+o4AKiOyJFZH85xobOSspdwiFA4tzT57
AfmeY2EXkuIUpOespcwzNg==
`protect END_PROTECTED
