`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NWnVWw3edRZHKsHeN6rDngIZq+BghtidJAY1GKYGiZJL+XUV//iGA8eilUMlYDhM
0+an2sj6m68rFUaKyN4J6Z95Ntcn4OkIDQiF/ryL2Txzl9m0p7IB1XOzqaxuIJpY
J9EtDs6sM+mrAF/PyBj94xiuvR/3ld6VLHcnD87R8sdbB4siuo+Xm7p5ZwIo+1vi
hPKcBlgR8SwfNq5aGzAKCAZOi6AM7YPh/ZOw2i4FcUp83lZo6F3knUNr0UGBEL1X
gqb1NuC3zkzNbR/aESfZUA==
`protect END_PROTECTED
