`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x53KXHB6V0gnZYajaumW2t8OUZHfQ2P+ZKuVagTPfOwsiJIl6PF98AE1BmpaYEPO
K5qIM/m/9ArwGUld8H10SwOROT6XTRWHV6kyWhqT69AYQbIfSg5oTNy5nS9l1FI/
ZExGkoroEck7JC5ZJj68jV86t95rfjKIGehd0hNN0oxWWkna/xw7RXgIg6vML8Or
wZ/ID+0is2Y3kiJlXipEvAH88FiCVUcG0KTmyYj8oyPorQvLp3WFlJ18E0WktTMF
jxynx+91NMqGBJ1h3zubm8r6PSHZDW434K09A3PUEgpF6rTaUrVJ9SssxDFNPIjH
zPwF4++YwA8SrIIqgfyqZnkHc+ynrlh4QM2F3im74I5WL2xZGazGvCxKNxWpfDIK
9dS0vJlfbMFHFDwuiV09pj/+nHHUI2PxCArIEueiv9el3O3wrQpFZQukXxSZKwI4
fP/iDCKvFFeO0/IV+MnYj0lZp+2lkNsft11SUho8Vz6wmX5bFFbcXiJae33+2izT
Q/7V6lv1xsIdjvQ8ULtgo8JkKr5+fOGF0dJCLeCMnT1YimVjcr+4MubP9Z20P0l7
aQmbYoIHiAXBbIa/v0lI5IObbURbWMsK4OCe/vuYNdM4OfpjrANgSDjI/Ml6QwRZ
sto+HVuEbLpMSfB3u1Y6oPMF2q4Y1m03U9BiKq5z2F+2yaJ69t5Osd/0kE3THqs0
4DHes2mCIGHNy7k0elOcPX8hJiZSpwyqbyiK4ytUIhchXJpj6t99mffv1ffQjovj
e+eFwwP6S1RIWoaNQwE9eXFTRxea2eKZq1IJjqUtoqsrGlF5d96DW5siBf3neoF9
WadRSGSz00l+thOqbCcciciSe4FJlhgiCBtB7aQ5O0LCAzmd6Ap6NVJ/0SUzMeGP
CVYFRzqmcO/IqCX0DVPGlWMBTs64Pjz4IbIjdJU1UkH+k78Y08J/w3NHaRcbixvj
U2LfC+Y7I6pBnt0zmTjS/CGvX/sjlIldnAvj/Er6AMYMpmiMruu8bIF2xcDL0xdp
lbb0W50jXp36/xTnDa/2ypSWpNMZKKHCmW+pFgApDPbDox2fHYOkfBDXmkmU596Z
ttzcxonx8nvLgvlNf7E/lR6+FquH3LXUZTVxKbdpeufEd8hppBMQXxMmphJikchX
Mn9J5A8blBR85p+XzIMJmhNeGMfEWyk7iG84z2L1LYZ/8hWjWFP7Yw7X/JuQDJyz
J7cvUChAeixB5KLDgRKTHDzvJ5oEXGRoRcl6IFdH09KA+LwglcUMFZNqUrcdbFzb
IFrD8bbozWIc4vrKlmMRf7IUn2EPwGo2LTv7yJd49ofLvtDZncFwiVVyTf5bftT4
Y4Q1bxf8c5ZSefqncjuqTnQLrn3DZTDWaOVhMC1uHw+7jNFLG56e6Y/vD7tc5v3g
ZrdvYTK9+JYpYx9sBjwqftiKjKIas7XtLtu8JJ8JgFVn5yynwB0i7X4ctXI1WWvr
e+On/v1hcMXsyViOiDRD/mzdUSV++s8D6pd7aPj75Qhs4pUYXpt/+THYj1tjFcAX
Ndki05bHA9rLwLzC3PFidoiF0uA07PaXNrH4kC3TcE+Iw2aLBYG9qFi5+7SQVi+c
VIw88pyUp8KaI7n1UG5LeOoYoNamj297Nz0H1Qi2dt/iaXWghS6fXkr/MmXozgOY
B2RSQjzTdY9Y+5DXZcmsswl0uluvOY3ArMrEGp0qvnx2HLwhEsO6lSYRA1qZ2sbb
PlLhOeG4dZ4QaKpZ3kANHO3OBdq6k3tD+bGT5Bg0zb+J0xds4SupSCbJdLggFV4e
f9yihDwFtz3yLZHkD7sySR35xyLAthh483+pQgG+T4TjmVk0egL0QorSyw8OCPMz
1GcPX8CSS0KO5sCmAvHzDXrKefyqKNwUR/bCGwVTOHzYnJDriQuHQ9mLW2A2z/Nq
N4Rg6rsUtowlpaRsqYiD87PE3/WLr8hHy9gf7NxBJT9glUXCzD6C7vA+2EQgDu0d
z8GqmfZG0L4UC+GSODdYEbStCcY9gMOxht+YDY6802ivYReCvHPho0BWdTJ4ETU8
E7OEnkDPVx3ggrJ46nS/hp/kijN7P5hACGEw+xs1eMdT+jRyxbjkGAiJnwXDiOc/
I0YMMuZp3kcGshCkn25YqkBTUce4Riq/rEU3CKjBQCyDeMj+yzDtAf2+X2Ok+wy/
cJ9MGOiw8LjD7xacGkJF+i4KsH8Y2Eo5IvvbigDDUkq7uLSUBt85FTgWVsuRqg8w
pm2YP2GaE8JRiFHAUH8jgt/WP5neX7L0ezrz+6AZyL/DQ2obODQsjo7N0UPjmhQQ
eCe+JLFIZ4EYFDTnfHmaJpUTlpLydgx45exjOzrQvo+ZKIcJokZ1UunIK6ikCVJx
YMZC9RFCCwDojJ6DyEY0CkOnZ908+qL4JOs8zyB2oyUpQTXHCi4YbTDJ2fMHf4o0
IqhVj3Ta+HpoXwZIcNmzRdQ3H9mkOnB6luzsHR70pFqKiLP87DIkW3x+4KlGQc+V
6bnSwdU4vOJcd4MFF1AjiclX/+9y1hc1T8rorfWRvcZxQHLaZDtdb+NTHXxprDJ4
wtXWV+FlUxsSVV7qcq7Q/jAildHPOjXPsMlk68lkdW3I+dxyXHgAN7FV+o+KgcZT
R3+mBq7NSq563NqsKAqvS8T/Iv6IXeD9TpPdVMJBGO7nTJy7jipJvYdAU19zeh6o
XILV43CXWprovA4vCQzzOkSf6johcwpaxHrQJ9SOAC7yJ+p7JjfWb5YMvBuz6ZWk
8omLP9QIeAecxKzxi5lXPlEJ3AqFs7PGI0fzqBSYFCLYw1CouuvglHc1sBSovk6I
s4biPXAm5ijza9WNrv0o84fvDq9LB91xsSE9qGvkInaXHLimqWpOAvYahzN7JLhI
XemCv1Ggu5Sl5ASYp187GBj65KJ7rarC4VnNP2l58NCkGfI9OrJ8KLoL8WHTI63h
BGzCR4Owa4knmjonJgAphBlfWSXMxWegZGq6cy1BnYARUOmN6rDt3FRtq6CyUlYR
OtpFRgH8/uHQY3M7vgEJiitn6QN0GM8E72TrcLKXgMNhvIq7oxPGOpfAYs0A0Cef
cfhlIxrJ7nRQN5+lIX6/NWAyepCNO15Iu+71DSxXbOMQzMoIXOKUUCvj/7gSzjsS
kDevN1JB77FS7HFVJajAdSLaEtTsCcFPoi+2DyCYaPnp4zlAfsDgp5WitX5UiQ2W
63Ib8UU2qDAcDMv8IJyGs1o8cseQmwOp8c/iTU8J2x9v4Zz7p//jNbHKQMOWqOL8
NpqBTQFTFhSgPxgWaX9Kf61p5sVZTcvKjb2pf1FkQkcZ4o8DFHk27ciwiUa1N2br
702POHAO7l1kU/2FJn+sOozUkUwWzhZBs8pvi8w9zJao//Wbx5BuOuVXyzEPhXHE
VLBCiVYJGRNlVXHgY6foa9ewyB0dBl4vilMjQ6gOs5fSlC61XbbjRbz9whLqNKQ8
9pEMqptAyHpAAz/NMBVPeWXRKlb0ErVzk1EYMnRrnwUTtHqC9RdT9E8piIYFX5pa
ahfXInGvtI5835ElIjqu23c4e22tygYV2JBt9IT1QTfByw6dVf5Pe8FW6VpqcB3Y
/XA7IYbolP5ORq1lMh5RXQN9XxnANIvth1uz4cd37hOcM/v0jKpiQAQd/dOSaF4v
0ChiGE23pfiMX8/+UtZ7wWhAPou8MtHbmfEhfFbUnEFhiI8WQ6aWmqUFOMt23bZi
0cT1BBjb3EvZCxVsnKLOOcC4QJMeaJZOhbvNw0zor1hkHKrvJaluf7qgeWxYNn2B
mimG/nRWjvoZefFab46kIJ0N3PeMsX+D+93oesmZ8zIXCJzFqQRCQ8IpIBOTH8JJ
TR8XX0pI95N3slj4wi5P0iMbDJfVOFL7nj59j2MQkVUfWxb7kdnEzQYmIHC4K7H/
1f5UnUrEQVNmKnwHHqoy8TW0g0WrE1rccRBxEmk9vxJ3v9yVuYqU5jq20iVjK+qP
cObSThanuHwldmKk0Xscr9yGzECs0AmgfRqY7ECKdPtergjQ0T1xNIMZkhJr9aZ2
RMDSrxPopYMKNxMLVmRxi9pvYbROtMwmHGIvOJ8dbKNmszrK9GK9rf1j7S4wK70P
UsVJ3ARBBkKf23qF/Oy5jtyUJt6CO4frfydX9/zsTTI3oPXqri56NP3jZFP2YClq
VnDG6bueZC1UXZ11FDc58mjFxOQEdUvu5l8GhM1CxSeAZqc0jZ/PfIJuR1Gk/6hF
XxReWah7uF/R9fxlCw9dK65A2rEf+KJVcWQ7I92nHtv26DBVWTS6jUy4w2C2L8E7
XIWxDmHP5PKViNTDpNJ+u1pmNnTvfE8s9Xu6CZt+yG96pKfMTXTibBXn9TtH0j0v
lVGVcjuQjohFTl3RbRyyTti9eqUsmQDeNv2YcIG6cCBRdNJujXPNi4ACNj4yAyIS
l2jdWRw2emhOa53o4rKveeQMWeLS6TzGCWWbz+z73OdueKN1hRLAjrpUYoX5TGez
BtZBZqzeRT/VQrkE+tzqIAbSBmC5jFs12pAN/OGiLzuT3bjECUv1QXZ24YNHohiQ
PaM3bvo9DoFJfR3Xts8BXKqFriKDE3452uDtQ3QQ6+j5n1B+etKX3RLurfAvrmdr
n/pTqeteyBslEtlGWqfCSHf+OulxWYWcYsPbVGGXIapaHHVlbyx4XO8G47nxk6sn
200nVBuxKPcmoGoCjWDSjN1dxRbOhkq1JW4/TRD5VP8c1F3DHFECybTdKzytk9qQ
2IFgYIi546DmWqOjgN3A/qprwICJ6uwfx5vb8dJHgj6EE1DwhKDNQB46z95zdU8Q
Yt1QxyrkKIdRELh2jJxzJrIM4Mpu5EE8b22BWoB7rHZnKOsXNAuTPtS5Ien1Bq/s
TBDu3M8anSlCTFwYnmz/siib83VgwINZzyDfOQH0pjbC4r94/u4QLTCKwFKhPKJa
rHwW2wU4DzcQqg2e+37L/Z2DXr3cgsQsGjRS1XupkixH/rR2nh2B1e39ek9hdjcu
hkUpMv8WsUHHuUknYeCc6eLN/NmS0LDr6hS3yVMnh3tl4PfPMKD7IrXJWiE7S5Nj
FKlUnqRm0PwWE11K9qUaDB0P08nMZE72f/mPLMVLhrxpUf9bY07AyMGRuTkQFJmS
ijaPhlOZT9r2wjX4LdhX5aN6g//T8777hQb7ROESXApuJ2TeKv08Oh8MWztTDg+V
xzzRNUas/y7HIY6l8MrsFFmAfldbdf6aJe6g5QS8MtFRtpEzR8b2QYzU/N4s+bnb
xX0yqYwMKfc5X+4+th84IHrbStYbgFSIivZbil0TDmSbPmPyPs7XDrsA+MCo9Pur
/k73w4ZCkF5mnAS96naY9KCFSK9JnVXPzJcRKLnqUJ4GF3IeuwauOu6/rAFmhSXZ
sHk8gua6KB3ImNG7I7931r4v+ilAfXzKyQI6Yz1vO5YqL24v7zEMkLPEvMoOzdzP
OYeTHKILwamsDVSR652UVqsbm7ayUc8mPcKsAhYyLQoA83lkOA0wAwvgu7unEmxp
fUyJp5KKPiIR9GlnzvKZF4N0Pk7VjdGErxPWIpqIYD7bJSJFXZhQs6kxn8YilsWi
BCQFf2qY+xowSsQEDScqcJuALzpDIjG3BBpNn4ZcAvOoRpJaXCNMfyn/BL9YwsCY
OyY/Wn01ovvWMkS3XRxYisl3xZPjec2C29dhVrxaboVFCQ6+fuMqF6pdcIkKTXyo
vYHkjsDWYaWP0xfAnACiSpeHywpmKAA3Pj9seoBrQOaDENBTIxmmmPqUmezGV+Vi
WEDRN/gX690yNw81mBNHuoBDATLJCGInESTZXj+RRElZoF0Y/LBCOy/IPqFM1+xy
zvvh+ApjT/6iJy96JE3ya3+qaRBTPvcqe4dShVlzVX/9ZLtYofbSdu/aALj9KMpl
zPWj5yftVc/ij10rDotODM420+SOxmXZjCP/lO6/5Vh4lSI7rtfMpUBTB+5EtJAd
TdFyf4AmGHl/usnN/HR8g4D4ccf4H6jHt4hlX9vax5/0VUrUqR+F+N1tK2JtAQDk
tEkgZAHqSY5XqD5yG43BFaFNjx6FHThFYRy6uQ03cOnYcHh9tnpYXxmOyQUf1wTM
oNYuKh3kiquOjYytDEIuqKzOMjXDpQirq7mJxl1W7OFC3UvdBjiSuLFMuqYq3mir
0L+wnBXKOY7gUJRZOv9wQg1UgnmJJtD1C2Hb4SUHqZhexrpE9YmnK3kvyr///nXI
LrF3Hyy1Wj0zCCxQvBezJ9b9kmz0hor49Joqsv6U0aEKCldzMKt0hUANO++FbbQ8
tf0D7eQXJsJOPTANpS7vYwWrvnObgeZFdMXE2bpF1NzV2y+e/6Res3RUllKLLoRe
Sa1qB0yWacjFYhMGA3oa+Twv9ypeeN1wpJzHfbA7scqDeterLE2HXzpZ99mqZ5vW
l2HS9FZokOmtUjrKmhZBn6DCtf/U96jQXFQJ1Y2YYmn+zCRNSOcHnsMgT/Tq0Qpu
80p9ufWsQWHsHDfXNFMh0KU6w095zQl/BVNKX0AJKohsY6AmsZhD1tksihg7wMS+
aQmBBYzlbr8ypk1zmVB6aNWv8eWnFvwvarQ1YpTbD6AXdiPtnu4SFRYkU+9gxmye
707dNZR9Cy6TRVliE7lS+ahDwNjfz3nlEsUQfMrxGRwzU8VIGLSdzaF66WCLNbMW
3syGKx/op51xsSBXcnD8/P4JElQjKt0UJuAyYwomLFraQUPlW78LKrq7X9c2bqFH
ymM1wgTPUIvpPHFeq5wOqIC7awv1KAw5YFE/zUmimDp0lop0qD9Pofi81euLJxN7
sAMN+Q2myM+2c1luO9EhoVBoN9NQ7Z2AiCdc8U3z5xKiihXj5yeC7fYykkD7rfE2
oKoovjwp4gnnBNttFyi4f78Zf8uNnOqvHuw8sCcfQdAAEYx1KfVl9rPHgN1yMfWE
nrlKknRTa4qfGbTShEpvwnmlkfs5QcuiCQ3i+Fw2V2bMHIVaDcAqyX8GgajVHLo9
tn7rbAb9h3XKL2O5jRA63ljXRj0Xhd6WIN02nRgf7kKR7ZOEDcpL7u87ZuovI2Tp
nvP6TjpV5BZczUWg5zdbvCe1CAMKoPlN64FVQc/xWrZPYxqwK3AoI6MN40f8PZ/i
S2uQVQm0rptXMTDSUJa5ntg36z/pIYBMwnyVvAiTEwNpd7otz+klcUgv/fO3GUZF
ILzhJPFnbjOHGTGSQdacHvjptC2rN9+6irmqnGIlqabwuFC0vCEOCX5DW8QJOIjb
PZN8vnLqABW2KRWxzr7zNcg2GTCDrVxe0E3PLyG0EAx9r7OTdigHIUjBUpufl9lH
pRS60m1a+fBtxJWvHOXK3UaEfhW2BoAtCQ8hiwVnnw56d7wjMpHhuLiUdSGDv8p3
mXZQ2Qf41pGxKVACAEC2I+KnL0L+MHBCDGIUuHR+gwXi020LB05M5ZHiptO4TovC
9rc3F5obGzVdSUwu0vpTxhClWEnTnfttpemGXLZHyrLHXE18Rs/+ueVYWi6ossFL
6CtXQUrJqQHQiE/iWPGRJSEs4QiscJ7s3CFRLz+mkQMsVS55algJkKAqLKqOS4AT
GcTexW4Z1/4jEE6q28j8/TZsM4Suc2cfE1boLk70ikcSsNhJAHhfCCMd8Rk/xHU3
ZQto9w7jqlF/ms1PojDMeehwOU/U4ky64aanVnkqlsk9LerswS5wVZcJqThZ1HB7
WMHmntlvg+jlOLuomuDPdXAxp3eH1KXTOdreAsnkntUiPZMJGoJD6E6MR0pA1Fm8
x8emaGmqKaa2buAqx2lbBmGpAdTPkuyTzo69hIu7c2Gh1zkzFr7ARah1AUl5DbKw
tFiHVRawnK5VtDeD2wcs5j/TXzaeX/5ZWs1a1uQtHIPtMNchCilwVAHbWFDw2Ouh
ZM61h4EFTZRYES7Rt1nLtn2WiYx+4rkdzezxgn+BdKIg9KhIhow0CSr4A0NEdPgk
1cy99yIFhyIY7mtJ/rt+ke9FyaQvPvCkRpAQ1xGOyueoV4OBhZjbqqvlE9Fv1x1w
7o1RryK/aMB/Mn9+jfLEcfSXEvKz6RMADaUspvhuR1jAHEwsN/7rDPdq6Ex8Ikqt
E543pdoKH+7yosObkzfx7LW4vUsYYUyzahe3VxyAxSPvVejO2dqdP6NPZm6+3XuF
WwT19qnZtTVT2tAqDATJe3weP/VUnx28Ql6uwS1l8V2FRrKp20GmamtHw7AepAsN
UakcJFj3E3Lnj2NCSnK1OOEXPokzIsC5bfr2rrH69AJSncGD6Ok8+KxFOBFFj8sx
N6Kx2G5YMbsSkYEgU+bIWem/3iZv1OLFl4b3jtBIdOEhezPAIQzVp7cSAmXYW2c6
UCK0MEV/d0X8NTrQjy6efWBt047r4gJmz5aCt/ggj4askWuJcOgaiXUWGv0MIIR6
CvtUnXCzsUQ80BxNprB7Y0q2qfvy+bDGKm0cf11rhjztD4STEbL/mgUKaZIt32io
pgRa306z5qKQAGvg/rKSyNU2VGf983YRswcdcWye89uxTQLvw44qzbY1AjQSgvbp
dhJHK5sdWOWSdwEZ/ZIuZ3tcB8P/3Ok2f72VpxZ7f3zsjU6Xe4X9SHD9vDPW017E
wGDBssJRNGknOHSDwRIs9Sh0FrEotZGquxUsqYHbxEXcgWsmZWjpNHEW/I1eyRSg
RdWmAjNn8np5T8vqTz9PRlAaGi2OazMF3TNOp1s47J3T79HA68BtUY6yvluS8ppe
OhOtbc11vdDfaK19HqL+nu5FYcnuGcHfePGxuFNrPRWkXUbircx0YH4R72+ks9vV
oZ5oVB1YUOEb/E/7ahR/uLbWGBlsAvo/RFwtNK1onz6GGipMN5tjOWj+S13Z56qx
h5ewueiYPLSFTOgIpC4MqPwzNxpqacxhZa/M9Nl8oyjXd92392fsUUSqjjSLV/62
kIptsyhFkntc9OGyjwiAdDxaBagWl/2ID2lSQkMC+1Q/siyGXfiOYqrYdZJL2k0c
CJ9C+FBg0E40lOPlTS3I+UkMocYi50pjjtoyH4P7XE0UnvDsX142Qud7iI/jpKEL
CpAp0J5omWWOycanAAtuhX9zk31vYhnmPETKCEQQts8HBOqFPs6M9E1fiJ+8VRi7
IqNh+1KqyrYQEEBGr3Fh+bsskFoQcRV+1qgie411stF7aQQMEXrd24ZzkID3n8tt
vjwwsanR0Am/022f6NHzFMPdT9XDZE5vkv1AvCixav3uzjYRIGGrQNhGaspSAE87
wxBoqNve06pqC9eEJpdYlZvaGQHqlYzx17iuC1wyoueuiALMOyr8u5JkBFJLVPRq
f2cZIkNQuMRPFRB1ysDQmnChPYetY0ZNfPiVCxY4QM1JqOOFavex2QAZSrCop5v+
XDDSHjM3qq8e1AeRXufnfHh2eCvM0yC3rK7Kc1gH74pjQZULu1fRNbvahGZUlH46
hYipbeeeQxjwBeprvwOTHgF77IEapTgmTf9Fd9ZUEk8laQPOisbotQKbuZk+3zqM
IyG9zGFRtcvtRsfrg65imUCiM9zrv4pqNn+A3NIG30n153csFeUXTVQ3TWMmM6tI
ewyIq3llymBE86ClDSaReTLfXH55cj896T0xOTAlV1bRuHLF5/7clGzkj9hxGDPQ
erT0DxhqHSS1CbcZEFjIs2dWfzxE3fbkClKxNULof4jcOOiHgjXbyrER0Hh3fraR
2ITGZl07MUMWJ47ynVJ/0SQocMhEDOz0ay0dwqCheRptApyS20FjRmTwYx4329/h
5KSEiAFN6rCTE0OnuWbzbkhnfbmmWUeH9JVHCcsfqEk3+NjiZOCIE8sVhtky7Izs
D9HqfZRjgfrbzEeK4hnwXn+pnselOsC2lefkwNOcrxC7MJsj/7YD3T9EoTftW21F
66dSZa+E6mblOWgnNZKDLRCfvisYV11G60kBMGI1mFwO0j+paWVC3RH8AwHcjSJF
7FnMhaiQxT/aliLcRb7ZpJg1LISSZkEDSECvV0EcdfOUjXplt/TDw/92By6+iSWt
bMvc4c1aYUFQtbK7buAc2PQZP/J0GL6kvIqCuWOxzuMSaD1p5hJj6a1z/QksuzUz
0eYm42ENa7lLfcP4KDiXAFOb9fmM8byjMJAeJ34uRyjGUnqSLtzVOFJNRvFV/jtw
ByZk1RQ6G4AgS796SpRUx/wGQr4n8IjJbM3hvXnFfcQv7ms8LkPt2G8NAl+xPUj4
xDkL27VNKwre1VfvCtfYc0NDDzUZIrOLVzQSzks6nK5bmv9cdquGYqUUy5m6O+Rh
9gfr+W59Ug1y5LMynM2Ti6Y7neklcJGNqTDxZlmxPneqJ2cdXNJRcrrtrtv3nlAd
jsTZK7lKmP9BROvrenR9wi4pb44TlXOQI3LPQuMzosMzTB1hnZ3TBaWarQ6lKZuM
MTulhGmQVtAqWqukEl8v3Zdlz5UPIvnYa00be/qNWa3KXVgny0nUD5Jo5w+g/oG4
a4YSq/HySGbPEu7ABkkQsHmaR4XMVEK3JJ1/nU/Y/8tKPR/QmFL9o2N/I7lAbY+0
ZxPcRUppKnlUQcw24DOLK+vjQz3Wf19NUcw5vSOIshZTThgaJQZzOdFyNEGORkxu
Aj6lL4DtxeZ0jqZ9sNxIq2nKUblEtfFS5bZr4yGufpYHMjQv4mmjGy5WXxgU7Yen
vRKxo6wKCrWP1o0HGSQjOeQ9l8LqQHWdWbnqcaRaJcqxBe6pkUhd5QKHED2pw4Wm
+abGoB4C6wlt5pxPSRc5Kg8CiIXo++IwuMLu/g3tOnL8dALL8l18Wtj6CGOmXfY0
5xCemWHHigfN5eoHgsyQ3cLCiTcIQv70eS3+2a1BFNdve/1gt3lTaDx2jXrmUHNF
sYl7VtrWCIY1/6UmIljKVnNuNLeSCmBhhG6giTC64RtnQwMi1o4eVsSIfcBMeZkp
Gv5PapfzOE7MA9TZ9nMx45o93AAVCp30ONFWUZB9F/GRh7NTAyKnmNYBlYGkQdEy
kFs2Y6IvBJhDlMaxi/xzZ8sXxZDjHz5xXH6eM/WbzHv8muMIcpP0R18knKogjiNG
a/y1v6ODxg97SWo0o4FvWkRgb5MX5ZMCCmU8bn/A2GhZLhDZRUswB7V97Ur9ZAdR
/fOso/dEhliUTH0/2PO433Kz37iH3bLiWLtN5EfJyn3jA5Gl0QHJugqvs9TBHmX1
gx+VH1VNn7Y3y6u5HgiXea3sTVevCbycVrNg9COr8cMMvAY9cJgtcRk+i8N77lL6
IC7FCTV2xdyu74m/2n7JvTRJRpuBqbNVWgFUWLIQ+saBbJ9eCtMJ7PSPR0eRELQY
xW1HXd+5kmMsvWqVchLbXzdP7C8sX/IHM4aKhZNZOG6qFZ2X1yPDLHi36fLwTvhR
EnSRvl4N7fVMLTd4H++bOMYPlSm+hZHRIR/WCcg6Lg79o/z3MuOn7aXSmcHyLKd6
hNGkNXqR+2AEq+aogDaKetZEh1NFV3yuEd87untporDoj5gzkokqb5WBUa8YXW5h
OYqPN4RvbjDnwIWZwcrhfWpPJ2s0mJNz2McOmD68nq3dJyWjOwGDXfFfnkecbguJ
CJqlK+67RV0YGLXYsulSWD78OgYJL35UANm5jVEU4gIMSeoRIvI9O09C1GjVlEEt
85ur2oq0ADa3Obe3FBHgWyeDU7obyYPEmP7s3kCEcZ+Yq5tuLdZVDpexcXR7YSR2
BPlQ1hDu18xJBJimRSviSWph5MelXKno0wm57ycfvzMo1UmOz/PhdtRjEyQ8q/j0
1hFlihk4ZeIzDGeDMY+RMogqxx8ttG8CAJczkmkfKSGwIbn0H2/d7zyrnIavGx/5
DuzP1GDelC8wIiE6cJePm0bO1a1fD0fZuE8ExwJaRlcbC4KG2rnMTqUJFIAU4Vk6
AAtuCacc4uNNsP9rEGoc8Fr2AE+0k6BDmnCl/KcNvN76WQ5E44iQHg62w+oVbWEJ
QJMBp3+EuO47JAUhWOoMvYYWcD2pxkm9pRZWBtZIr5q0K0TpfxwKBzOVyIt5ObZG
DOfTT9OiaAAYMZnh0iFvF66ULAaj1jTP8Ux737JlHmOxQS4Bqi+bpc5deDOMC4w7
r/NzGWGBBIUYMRgIO39VlEWlmLxz7aKSgiFDeOhiMxwdXczz9pKFz8HhT+aUzvBm
L8Ebx952pKjMA0f1YctD4Pw9Uc0s27SWhMJ49kXcAAIQVJqychhqIb3g+/CYm361
ggG6yS17sU8W2KcWsvmOMLk5lOmvc3Ms9Kjk3tExSKAw81kfk2W50jNusHyumlfX
M0T56gIPmDY8S/lmvcnAumtYzHPYrKch4m6flxcujjeIU3RHwWtmHR699GKDl3ha
eY+Z3pQF2+08YOT//92GgAdmQErreAIMLIKpJQH1PtebfnKY4WLuJYJ0dAYfUq5d
m+5DKv0dx7NUVdkGZGdbYl4KSJW9nl/DK5PLP4q77E12JLU4ZMDH17ApL5zqFUMM
c8TSfNL1z9YRS6tmea6VLEU6MB2z9WdB5zophxPIktUO6+0wlzFdeau0gnjwqr0e
GWO6/Sy2Q9xWWSeoXskZ5rHNbF3vjDo67SmzTCjXO7avt5bEq8o1uo+VCo/sLEbS
FPr16nTuYfGHn25a3sfyJaBmtjmmNqt1TljtCKpn9B6VVHE3toIEQqP7E98QVTnr
3AS/k+Np8pUCe0Z0bKfSwox341+20h09gaXmUKX/0RHV+jA5rRdL1AJfRgFd7cft
Zmuj2jcp+vydnnGqTkYb8MReSo+bYILP3oknZx9Ehi1jajuuYY57n2M5EDGYl/50
sDE1VUbqUO7EqNiyHXRNnPTVTVMWEDTgt4Xiqxxmock87DT0n7VHBIrNgWRoY7Bk
mRJhKN9uckSCeqiqbq52SzqFLNVCcv+JW4n4/FeK7OPr4Ws8h9rw0PDiTf55hoF2
jXHqewlO2ohMhm+5QFe7MNRhO3RNEMGTaU/8PWroj1rfOkgISB2xQH1UftEe0YN2
VBrCIv1Y8fe4QNQ4kQVhm9VmPyu3RWrbFDlrACwoh301d9rnvCSfISZ2UStiGL83
gGKEk/QOeWDethVxRfEJP568vfG9yZjNiRHerNlEYoE+sb27Mj+og/g1I72OQZyQ
ha0C/+UiPuYTt+m77qO4+x0d+3BRQM+dJ97cWfKKexpn0DVSoPQv/GSGmDH8uGhJ
dE5FaG/3gwIGH1m4pfgUX337s6E9AMluCyvFgv6dL7uep8o2VRJShR7EVyX2hIWJ
SZjAKfoYrX2Xy1R9J/X5mNvwNGKxG9SpSwztw2DkHakuM8UsUa/XhNhmXowqllwa
+PtsM1n7faxNHAm545PmX8i9egyHFZAeQ9+GDGaIHb2ZS7zTE0rO6q5G3ZIBRtre
Sf1PNXo2j/F4UwFPSJ4h+GnkpG/aYc0bENnlyikHnG8=
`protect END_PROTECTED
