`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iGSiAGWZZHI0nLhTR6tmjBs4UCo1IQzbGb6EbUrqr2DrdD3C47WNg9VLYT8KlQd8
nLIxp/o0Wgb62+MkJJ9H5U1rD3l1rD8Yix0f8D5QMQilb1vx4cJyLqX4gt+IlwOY
erP6wt4OZDRQYqaDhHrUGnTCXlQBUlXshx600w7AwTV83G35K8L5nIV6a/NqzVDb
lYVJxyW/6r4fJl/DTNWB/cW9nNQ/UMhXU4/yOBhbUij/7H0lE+k8KgPGvalJA2az
h2IL3tjVSj5635qWlZ6DTLLLpt/JOJSEm1hUtjh0G6t5MJwOCLJs/NZSd5/hENmO
q0Mhd2CDcjIO80F17TybNRB+g6LPvH4hJdEeJtGXjTXxyfyNnE5NT+UnZ8gwUIGd
Ry8ctL83R6avyb73lXBk2GjU/eUb8G9fZB3y3Hv5/uJB7vONyoBKTt7lxjg5KzDP
Klh7V58rzMji7+h+7PeQrU9LK58glTjPwZ2wVSOQNVuFTaMvniZ8qt1PkAP2Inv7
dOLLguN+feJaeUCPGChBduXUjyZYVz2yi1WG0gmgcl4NV8JRYnM1cjYWcbWv5jCK
1jjgaumNVSWOfnH3MKgBEdbTaAaoO4lI2Q/JTFvLIacnFb5dCknpbPNeKqD1gqmV
N4cBkBX1Ih9vUy/pMK1w3g==
`protect END_PROTECTED
