`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nh+M/up7fBE7oDJfAlzKPRZcFxm9iSGFWMPCuH5Z0JgYe+zZosJ/fKgFKPZizD1A
tAV2GK3tSM+vivZYXPtFx8sbHur4u6OwAJkuG5numKhzQ6knov8PCMlUxPgkled2
kdAxZ78Rb0JdgidRiVhxYmtYlcegnUhF9Awai9dUduuPP3WgbvrHyVh/co+Jp/C4
pF7IbBB1rq7Qy8N80HnxRzWL+goACKD0WzTTJ+ZjyWkWUMXIx1R3jjy+Bp1nPq0G
BmN76FltB9AmdwzXY2jsmB2THu+qyL9H+4FXv3Xj7EvQprs9Ph+3i2i9txylyFhh
ErfhkB98l/swNH62eK/MIQ==
`protect END_PROTECTED
