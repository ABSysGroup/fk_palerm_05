`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gWjoHG2nTyLAzEKbKUDGbckZeTx9M5jFYgR8YCwjZJuxZwzzveYy9LB9ZiQm9IL8
oon3oyE8AwHyLKBfNYiurqbo+nA/TSb5LBzBp17w3E9PswaE75/kzUp116UzFKwl
bolxnQYy5ZlGu3gqJehGVAkc0u0OHy2GWqyGW42n63D7+2JGkmAqVwbSJu/cOIu3
mQcYT4vfRwiOoN905DDOJgZUus2gs/cgzIBZGTnfAvWIGXCg2hXNPfLd8QztHrIa
FtUp8bbj4fouXtWgsDgJbE1IyIikJyXda46X0+/1dvCUarFFB4YewN6ouFednU42
fSURw4KegUHucSDevE0xkVJZp1DfHSa2BnznBx/0bt+hBAPWqsWwwsT270n8tVE4
e5xfTjk0Ql/gRYFDl7elG8JBOWkLY8s0nJBqyUADkyzjhNH8uAOML0M897bYAK/i
ctG6clxpNkrTbw9T1ZyoD9Fp4yy2IJ7Fz5nIndgOCk0VPf9prObklwUsPE12UARZ
Ro3xYXURc3+QzAlBrmqE13eI3Wh3ZWGKS1GOdHxbIH8m2GOX4Iyc+vcbwk/eLFdF
b/FfmKZPAcxnpOHkdvA8Or7S45TguLYUyHCA+NxJImqJJm/Y83w8k7zD+64u20ht
NITs6tYC97C/I4SVrZy1vVIGkICgsiAwjby1Mi7a6rc=
`protect END_PROTECTED
