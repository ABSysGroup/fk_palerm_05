`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7r/EVrK2JFevqa1Evntbk8SrN1DqH3mwza+7eJN9Xy/aDvftpDidpXyyvPm/LP/S
kMn+YEZ6vCFbg43x96kWMLSRzc9QM4eAI0SIlxWy/VzUjen+0j+xIfWXXcUr2TRd
UDrXblD8gc7XwATOmcXCq2ExvkDBEKu78wQyVGWz1/kmF+TuXX3ZkZClOl4RIUx7
BC90wsGj5LSiQSf+NBYKTKSc76/T/w/a3t/h29aB4LUpg2TRuCM+h2Hxkjr/2kmF
vjZoVw+lRsG5VegAB98gcSiHk71w9RrIDPTzHHQhSvWVvD9PQvZFmDr+mzLmXXec
1isTKywdY4VmRBhQOoDY7rGOS53uaMNiWp75jiSe1k6BcuD9kIZAvuRmc0XprHcd
lSa0vitiS+5F15jEnpcb+a8Bv0kzlLNIsrvut5QmVXn3opIscKRuhfopwnLWJcrW
0/N1/pPN8GjYVF84br59GkNYtNpZ12TRv8pBv7lJbY5BOpIggUm/QgqFMthJ37M+
AaWX1ULkGRbne/fmqhpf4RzYu6CrcWNZeVG0b0x3q/xW74SQb/zKJrJ7heogItzZ
5Tk8XhX79iIrXTI2kDAXcl19dk9NNYGSKv62MDx75N8GM5nFQDeO7tkqA80T8zHK
cu7Iy78kD2GiM+WnktpBp0pEC7F9H2vO7qY6MAQSAVfG7vxAFY8SKvDQencqkDzC
vcqWp+/FVGkwl/qGxppQqymK9T7iHIBE0uPrMUpeWflEl2TogUM+epEnXLHKGZxL
r0DLjT3DNtLepPOZpN0/ja80/KU+EM0r4jJqSdlwGAh0JPDupsGNafMxkNyhYj/V
crgNsYzYGC2TNvNffnqsvndj8BqlhDPP+AIKZqEu1s5LxNe59c0WOIymMy62UnuF
bhoU0lAsw5JQEZBh+44L5uDat6jT8ncAol0m1k/KWyVp90da3Z/R0Y16eq0FKexu
ZERpG3qMjjwWhfjqX5Me3ag/+bQeVZHyP5fdHO73qRFZFSV/XqPNX8++RQSCm/kK
4xliseu9In2wJCw6kyLJ5VfMtqZet0wpYdGp9w6G5RLNafUISg6dydy/jhsoclwz
ZJsS4TOmtfvENh5W65jQjjk12gEU3idxc3fzV6tqKFjCaDpd0UCHLocrAYUNrhLa
reLsNJZYRtWsn5QbyKUiIjMT9SgZ/ZzzbMjjAPjLpPCr19tH2trUz0p7yEagJObO
tC4a0EncleqXB9qbS9160qSymCEns2quHfrk9kDzDR071cObLnqwFr7pFdP7u5rF
R5jMl6Yg+yUgVr6eoiEglkNDE5jasx9/RxlWMGimPTQ2siHUm2sCljyZigjCbC3K
CA45lnFJAU2iZe0bTzoBWGITEKdeCR+TGCG7ChJifzJoToQ6js2Y6TE6pg+wZ6XL
9ckHRs3e3nGY1/bVoavSXXYJzrWQC/Ydp8P5tV4G3lwDmkfjemY1gH6Y+VdWMQJo
vkX/mcaCQlDP/aSiwrykwNBqrNMHQwaJv/FwAWL8bm4wO4sN9I7RnDF5LPa58h63
QF2t77Vqf2t0qZNdht8Gou3CPXlS14tBpjOszIxaOm046AcHLAkBq1t2m3MutsE5
Xr00yZB7ZFujErU4CUksW25HQYA8XfpPN9iGmyy1ksvt1JKcGssUDF25ECsbQIbQ
QDoMmnMn/LdYfyAVyGjGxgcngTpafL8AWPOrDS0VTBoM/7o5anMrnHb0Z4I3kgY6
FPL6ZVBE5FQyl2tBJBFjtbGh7FeRKimuSA92YboduAPP3qQhYxK4eqfyRN7ez0MD
CsVVQNczRgR6/KqF1o9TQSheE5Yg3PgpHaUTMJT4cL0TGvDMSTmxEJPr7NXF+h8D
ngowCD3fYYWDRBEzCr2hzELwvLdMttbtDMdNpVMULD1h9lgx3rxgl8rW+l8kG3TM
HVuMBoH4KsowR7e+TyHQOBFCZQ78Z2uPqbQIgJV9taSdRz7tdWCp+KDoOGNRK93G
skhH8YaQ5azzSyf202pLl4RyehNr06+FAGCMgIKr+WpBVVojs56JZm1W8Zb69qTa
9VHNujrvvD3/jLiJaSOT9whLs5Hn22irKPWreOLIfY6CNjdUf3J3ylWupn+SDoec
y8gtBv3s5EDsmtacxn1bFcQ3T9doucD4wCS/gHfCWT82YAhnbfqId9eHs30v7Uhy
gSzrkoaryz1yTGOxyKXeO/oikcUaaUwDv8qptbj+NgjuzqKzkN3yk/MMgFyPRCO7
Gk0VQFvZh2Gf9gEjwKIBbgQdY/AvtlYw0YQFWcMk0vCVYDj8nKOS5S6sidQ2vbRO
w/bJTd7fCmVkUGsQpkoj4Xrf+6y8aTA9AHt3Y6PEiBxiFdNkUW6HMMzpK8k2Y3hh
1Jbh51fWlK9w3nVQPVZ8ZxzAtYuCtp9VvrWPLh4oBd16xyGfyJk9k2VQgAKekaHf
FL1+6IjR+p0QR88iMSi0jB0707D96QXiq8Ae4+p2dIcenwmX9FCIezMkrbQt2emc
1WcD7LgT7PePn5kV9Q55lo/+v9EWCRjiyAdovgI8JyriGSn2jGlHI8haYCTMmgnx
mU1xIBq4Rjmrni9MKoqI94o4se34NLqy/l0fKR5CBvPFEFbceTXG0gszTEhzRbzY
3rO4aV/5zkYAx36EbZV9Y4jZH4+rXsuPS/HGA8y8NT90apilB5Hw9DpFLV1lce8H
GgxXSdfMFqJSI6zmTgjmMpYR7WgCO9nX2Ka3Ac7ZGPe4a3Kvz3b5dfHNSeNuuVos
Zmk6RBYUFgyhTH9VN6BCi7x949s4qJSclPccmPUB9DcVbVK/1iQ4jlM8F1TttwZC
PkyQFHcC452EaZSOGG5yOLds0+u73R3hquzoTTFWrgMqQQYVdLH2DSiHI5nhnWr5
Va0bxXNRt/Eh45N9uAx0BSzqbLt2QQC1p2cz7Y/Vp8HXgYJpPs4wwFpDVm9DBbBN
mqFY4dOP8lhnaUpZQuCaOyvrdKA32RakvNqPTe6yN/wFlGTOjnMWjGBgZvS+xHKi
blxxgdgGu51LVGWEFYhJIaUuX/W2RkrZ2FBamYWxuGyAsqY9Ack5/knOBWNYELgL
NTCgJmo5VJ5qOWEQAA6ZQRF87v1SWSQhhrf/x8v+Ws7CWmxsmZAlNa+L9huTYaQ6
dX5iwOvVF9g3XxPqQek1irsFnff8sG4j/CBkL/AKApNI/u1Goa8hzrNmmhHfofS5
ddGzmiN9HUKs0b+XtsZhMY5uoXKvmshMbEPKziEXIYBukMS8inHhWHx4I3hjJMAB
N1vcHWlSf5jZefAwK+rruecK7lbLQCkV8c82DeDeZNEKo90LplBqAeM3iS4G23Co
xOU3hV/2/9bb2MxE0NMdHwqY5GjA14IurmHD8cRY2DmJv3RT4uhvnEneiiFYW/t9
7Hc3tngLUMsALsxtLjDgPIoGU3aWxujyKnPGIPks8h3xwkuJhOkrEcsD76/WFlRJ
NuDulWHJcW5VZWgUmfSeieqUYwgPYd4WhW9lRfMzwFx0Lo0jzQSOWa+Gh4zrA3Ed
rD+teUNLx9M5etZWpKKm5WVe2orHnZpeNUpowAdAtULicuFW8Rx36y3kLQDmEc9R
4MRiE8UFj9/M7GCtvrwRILJmu4KeNXRbEiVn7HRFakalKizRmTejbfigzAXxAAXT
dHIhMrKrZxN2QRDZGhVplc7TwsKkSNvk62DZuVvkTX9zk9eCOXLDaWzk/1ZeMS87
58/dlms9noyFdRZYT1oknRVhvzA6YnX7henhVtTZEauV6n1J20OfEstuTR0rPiil
ZvzqapFCjXkH117qMdhKuzvg5+sdojkYUoR7P2AjMncriTtSGClULu97XC+95tjj
pWf1LRWQllyvzDjpYhFjfUV8SiGgBHA5QJvyocdkV80sZR5TxQ7C/yOC/vnFztl+
06N1PkLQtd93/Qyx16XUWV0lmKDLIwvOiE8CBR278iNyOrbitb+HaVOgd0l0A73Y
xadnTZImecfkba5Z4WShvYDjyt9i/TVIc0JCLGFLM5FDGw5cWCvI5j+Rb3GMphC4
FiJeTAqRocn5c8UzVXlwjaUBPguGMpooDFwLUfXoUTmocSC3/MFZlzBIRjysgCe+
6RIuGXsn2OSCr+5K2jkN4w9T0MsX71RFqZTXkPr/IH5CVHKZz9aZyCzHviA/Y+cy
PAA1IRuHUxtrjaC94c4ZrT73t5+WUsmwBGQ36yQuH55wCe8RGIeLlrI4r7rznjzF
2Rkyp3HuZps7/sPVoLZXvWQ4b/qGqipV8AGq7mfDiRaykPUk3/HEmU08COYiEup+
jW9vBFvPkxTZ7iMwG+cyIb4Ww6jaFI4lJL9ZQzNpaP9F83U0+89jxvM4Pu92bHnL
BsVfxErUXKUec0Wgz1hnVjOqbrPzKtz39cqtPueHTaUMYXwzCSvfNOdBuu9j8XO2
3y2SQyaJLsPEHlj1WILmMHRKLjRXLzyJI38/+Eoh+94va/X7QUUISKmuGzLNtnXx
1+QYY0AiFB/y+6M8gCv+dQ4UoPAW/IOdCzt+Sizn6c1dbspjKplWoEDDkFzadwCt
MnxXt6yPAbzzXiVmVj9SWzzp5SHx5lZpKMftbMMjxpkvhLF8LWuxSWYGRF9FUKYt
9Rgkg3ZF5rFhoQFq36+ddUvgymLqPCb9TtXc3O28Gfbh1cyQeWOcKmk5+2DxwMsx
vlxL/WDenCCv/faI4fA20Ck6xKuzKcuizxOSyQVywQE3hoxpzN9TdPRB57Vm4wu8
f75eJcpt5Y1N/YrVmX79707Mpj7Hc6M/mD7ea0oi6YwQAGpMn3hDbeiCS/SA0zMZ
R59klom77bLeDie8Oz+WkWFZ/38SGtLW9+1yJ5uBergW+Xu6SB3mM3n0I6HOOKyu
MpOv5SLjmMaAh9CNGWKYw+uTvgkyhspvHVwNEFNNIKm4pZlrMtZhVniOGukrCL+P
FRdknt6fmgxdEUC6rBH+cpSWWD7JouTuTqj9ejQ0dkEbZb3irEW0tigfxOH6AZAa
4/q41IFbPApvBaJCmSoWkPMwl3IoQllawYQrbUJGA4u8IVOk/EjLykiq2+zp//2Q
bhipYS+rLNL7SkQkcGzBgJD7a8Yiowt6TVY16nXKDuYByviCTj1BALH7DS7/t9rL
QmgE2jm8zAjt+qfbLlMpla6MLlCtpdd0G7r31i+Q/PTaQqUGvrfcnwye3WpIsXiU
v36pqYP29eGtrIuskuCyGcY4veLkvNE1hE4oKB7gSU6ShkTHbrBPNSi174u7RGNv
xKTdwiJR4dCLEZvg+pTcy1LFK/CCP9yUpUGWX+bYwuPmNX7JgYbye9TRJxyjgGac
gv2rapqUvYAfI18WOjCCMj62+eJX+1NhQgSp9xwLfGbXv0Peemv1B3QcPeT4Dj34
jWX/bExDWdTDGAwmebfaqQ3IcNFmCAdywh8jQ4xr1biZXZFp4LDz6/p3QDMhDQHc
jcPBlGuFcXhdoY8n4HnzbU5IWOkhSxKH/fHzwqOoD3P4P6drk8+bHddF/YYm4t+e
KUIvDaDCL3LRXIswsB+CqJcvV+whSEpSjwpgHQOCMpVCl447rGle8iCgpuOHpsIp
dvwv8XFQbtvf13MJkgf9gPXZwIdD7T9Xq7WxMkUI/24pWty36csQA73eHJfdcIcc
Dp266BbCQRgBrusrKkBVRGa4mKdUGTqtPYa+wbj8qIymbMfLREqadOzexQFz3q8F
sJ2Qe7ETSIU/tUngkMM7mkI9WqbYRrszGabpZUd1SAQW/VKa2zLnqBYIPp1xZhOd
JCE2TldqqTFD8b8YJLgkcxyq5f96twGm88DeDvNQDaUDAttrgbroxXUEV1kuZmnY
ubzKODN211MbnXimtP5KqIPKS6IgU5mcUoRwvGL6kPjUbYlb67JYPKxvUE+L0LK6
37vxSLuqk5F+WS7ejI8azQ8zund3fhsjW8V0dyFrDWAG4mD9Tllt10M/MQZW2y+7
w6WZ6HWtsrS4zqcFLdqChnaWFGDBkUOuL3rXqGfzNPXAzH+qedRsXMQDGteirez7
gI5Jqfkql8vmNqFm2nSLQKh3fDra6b0F6c3mJoVMqrBMI1VuLRgyjZ7vAscAH8SU
13+SiRxsRpHuG9fGFh+gOQ1bRCBzW877oGyg6bfH//Ep1bmZzl2zzXUHgkZwvnWh
hDibWMLeU23ro4q1VDtIDkdKQXimgU9dar/2O57aaMFhj6G853Z799O5xjTb2sQe
Afw6/9i/2S0e3AWT5Tt6EZOXsGPLsklklecpvGGp/7TH9ejyPoaA6ScAe7ncBOve
dchPBS0Adu5mu3cTXAyqH4oC5fnTwVbsK40h7c4W0PzolbXKj5ZXvrpQOpm1Wvyt
SmNkhjUppiGCPLVyS2sIDIEhr3Aph1arRdosQPqa3VHWsWhQBEFpcNvEQ4Zu3DnU
uYv14ucMA9vTSqqPNLXgeXVRbRn3C/9uGVdeiwy6CtxC+vKwXs5Fx50r0mEi7g8+
FB9bAQU3r5+aQTXn6RFdHFFzAwLr46X4Mx34N4R/0vt2Gl8hXGzz4RNbQ4caeb0K
wy4Ng2zCA87a9SRw6mW3uokNfXnC0YUbGMHbHRih2vvimCE7IbU9E235Nlc744AO
LWgqPw3ZmxCzP5tHqhjc2+mynkmZgQp+ki4FByZpRr0EnU2RsDr+ojd7JVhNzDeY
2l1AcwUSAwv96+qslZE4mXJzPM3TFi71u6ukfczKGynO6ygOIu6lh1542dhK68bc
2yPdbaMsLw5CibbYBuVzefYOHNyY388tkRJKXW+OV1Kx/7gIGLki46SEKcdo5bGx
br5Ees9KT8UD2shyAEVaFw/MfWOy4BKSb6WHBr5MMvMZB+1b5bFn6Qx1mddKpsu3
u/rla8arkkYuRh99gTJG/upBj+5s+NkByt6UsvTEpnxtS3zw/OQd+Rmhk3VpEhSS
fxdUhDT2MdnukYGCWF8vppRkhj/5Dn5KZscEzwCJ7G2vcnk6byT3LsVxxfMeiAhy
diaA5Gd5KT+Vrjs0fX9uoHcrZQUg/7V5F4eCNSlQj3PoNE6Wv+ZjW+xOiJYv7JwZ
wr4x8QmJ1S3vfuokJCJKdpzFoYZwZp0i0TqgWfb9BELBTA7AUhDCcHjJstt9HmVJ
KdpVMdUcRba04eHIJyypqhI+0oFJ2B21Mx+d5+A+1xBk9NPW+p8eV8L6VuF73Sjw
v6A17mNzCF9NlKmeHpcrJ3ZQUk5Q/e491XYojgGfgqh2WLa74Dff/E7tZO3zkVYb
JdId+6kNRTv84q7Og7JFWuSyupAsMt/RMTEtNmZsw2pLS+G2x3nPCjQlBUi4BVMp
YfowWc0DiRVgsQXivwAFWLEKWJtdi69nhVAn2ct7EwRfrk3kdZqdfIzo+qciwoFB
1KTt7jqDn97q9VOtWb/Qem6JLxoPSxi5gBWCUSVj2UWSOe8yl7a+r+rs4IteBJP9
3bWewZxuIdiY0V4qTW9WRaE4RXKjlfMcjkANLRj9ltUeA4nVsnosr2Nb8KicxqSH
sy40oOq0/tOFG1ni1maQyMEdT03KG/Qovj++CSyJ9BKXh6TqgAg2WuY0B4VsSruZ
fTHKqHDnawCfjXQVq0XvhacfA4Fjao8bej2MVm0IhT8YqUtAtJaBNZv2hRlI0W//
Dzpe9JILnZTfWX0xwfKT66Yn8l/90Z+5syVeNbuj0xUJM8KPFLRtKPIdm+CptWfw
qcxQ4LZmRsGdk6EyM38rXOXWNjShLsO1AytR/PHXPHVhg0XFXQjgDuoSI9F5ZrG6
jOSX7ogFkabYiOge3WZ48wZoXOzRzwn9DrIFqT9JAYQm0Y0xZY6LRUqLijp/huRs
WPhHodOBdHHcC+wbFCX0HDsXEdaEvPxu6M24OwfCn9+y03v1m8LR9BdN9xHpIoVL
fT83JSGFwtUO5i0cq/zNdtLDPCRwO61hLxxcr/MOuLUuCODoNyunRSlOrLjpOO8Q
w/NTp5yWaB/r5nX6l0GziRKP1d6DN7Osx8K6nWMiGxezg/ZFikmt3m2m5tzka5J3
71GI1w4UIcoJcIaAxCrq//2TjTdVbv5uGFKBb5eAYLXopOzis2RsS79mQcnK4WrP
8UUR7jSElayeqFVurAdM9HSthB7ZGwn0AN8Jvh1qFEAQaHZgO+pjMLiAzyY1ndwA
SkMBLBbuQUcvhcb73IxwMtZU7lVa0+0rx4xNUV3MkwMnGFjYYdxE/C4tWbKuHSSh
GUu3X6KKLq3IbpJ45NZdtB3xtSL4CHj7O2KYGkxhyI4XIo9iC93gtX52C4WRvW5J
fkPhnG0gEvpr7zUUrTMhtChHMHhCGcQu5OA7Yf3lwtadVeQM1nQi1GfcpidTwCZk
2A0h7vWHIPYz0QkZTmkWeBS56bjW/CYuPrFj8KD5yF352k8GxkPT4GCjI7wppYFX
26G3Sm75Niv316qRsUzrwYf562C+9D8tgcEPfnqkTmCYMDfRsNy6wY11xxyPlUsm
G0CENEjWxm6pqBsnTsXuILHkWJDOUZUImAT6Q8De37mr/e0jCddS7vZVmrV6FgjY
0XsMwMyItyp7Z2+baO3kI89KjzVwzImuW9GRiSytclkdcdakgPGw/eXJQGx8hEDE
WGqDvdyzfTkTCiLU6NRNBl49rHA7TUzw2cGuoC2mZvclWqJ5j2966GRwKfMt8DvW
mUC7/Bg0kxRP+Vp5WFwH+U6j+V4Msh3xuMZPRv8tj6OnKLN7sPWN9gmEXFxAOyXW
tS4y5im8wFromcSJlCK2b5hP01gcQAbgLT4q0+DFfrDtCL+Ze13uEm6eC2/0eKFA
Ya6FVC+lUsdYKWyz7V/kOEFvUjTHRW5ZfAjFFNtgch2OJmWVSwDvODeoxQndCtJ4
LXNpSD5Y3Rtr98uE5bKJNyVZ5iID1tISTGixVDqf7Y/NJ8YdnYwUWVJeooJ8xY0/
53p/phTEpgnFq1wexHYT4jLmcPaizSf2xuPbX9EOmuqp4KKCcKguQm7bnAw/xd/Y
eBGhtZEYPGYF6DKYXw4VGTGLu/jm2txmyh8Zw5XY++iowUKKNctBh2JxZRvuvJb/
auQc781wUCj462d1tYvDmUUKKsu4JxNp1gGe+s6yPcnx3CXvmOitB/U5H8UB+YhY
fW+QMt758EsQ8HaHAVPphZ2Fiup/U7iJb4eo3H53NH/j8tJHFrnJuaXQKJJbHBa4
xMTRh/vREkNg8OA4QuNtS/8MvxLI3Kivxpb9kKv95fOFk8il+Z3LiMS7WSJhGOYk
DnMM4Ios4yJ3dziK3ysA7mqoepFFwgQKMBlOXDA2Z0F7dzAgZVaYB9X+UycUBojZ
QxV5OEemdd61G7+uE/yDx+tMRCKPebcuH/7HCaQAHogGdfF6np8ypB8y5vEAS42+
IRTooSbPJyTx+Je62Yz37XTd9GtlM+zpoqpUIkqecDGt8KEzZwM/8NKYMmfGI9JB
FiKSRrZuVlDqoieNXmXZfya1o1xbELlQq+ZmBqz03ORzR0Ak3bwB9+0wsZ9xlBXw
/esyt9syEV6hK5GajcUW+Zm5sxzJOaOadkPDWaWEznt2CFteMRdgGr8fNJw3cfri
e8S0Pk+gPpeFqgHMiHAYg6OFIgePV0Z4eM6/r6m90UEVTrW8vt1t5eTB0jyFMgs4
O3/i0uwCtltupv0a9r90Dbc0LpD3Zf4exSFEe6DoAKGsDj7MA++QNZ5tu39hx/vu
+O53BPbLP77puzWOz64Q+O+6/Okia5jcm7JMBVlwhlOXMkFx96aOSsmU8NQ6ki2L
srBoroKZ+pfC+2slfR+z/squifJrq48mI1MycElepa53+IWIygH5PsLpMvLawJ0W
9utAPRosjLqwgUslckdT9yN7RNVtFxe+QvCJeLcoqJ+HxsZccq8/pCnT77Mq8u3W
kSXvQGU8nv0sKGXKhTei8DWIa6v4oj5EwQjGYOvtBYfeJ36lu7HUIUjXBGfYARJa
8JNIf8SDymCI0J86b90pO58x1EYGsVrmCRBS9LuBsUKLS1/+hku1nfD9sw666yFk
r7aY24N4yepUQmxUgc3N5xiV1jWXHZO8i3u3WQgihMZSBGV+rOigGA/awFBJUKP3
vaqBZd4Wv5fWwuuhQ0RXGAvd3UsPUAP586Gnky9kw6q2CeLOtDVVHR6x/eSpCT0q
vya5WkTJcCq0HETHcyzfKKiwu4Mu/fGfQ5H7wkPgjSPmrMkyJWjXCNrh6Jd38H2X
KnD22QVT+tCJL4NUchvR4Zr4on0301BCNUsxvrKEAmfGBZs+L6SUWImXvphZHh39
ibam1qqgk5gN7XYSMjqxISJAGyiSfZFRu0hdUbSvdHBH7S6vI5nNgdsbctnvGn1M
Z0RdGdudcSnXKd1zeYCCT6o32ZNieNutNtq0l+WBJN4JvNbY4QDGlDw70mlmYgRm
tNq+O7k9Rw6Jg3VGn/xBU93+vekOlICPVxV9sJUDG8SCVdjasfGgZPH+uYUObAPw
KbKVWsGyZ4Porj09M5oRMSFmNQfLPHxJwzdpb8GgrhMmyXAcQ238f/nGDwPuk1a+
6yFXAZTb46eo0/1zNqwMFK8wPeA7NVPPWCCgPddgs8t+0NDZtoAThYIHGWbhhrQx
myLhMchhiJ4B3Q2xKxPlFiwUk766TIv1Iyf+rW3KS/TCAgMc1AlWg3pxHmxvwtZG
0K2E4Q79WdTDpVtDVhbiqzj5hh3JO0m8LdHyJl1QpCcmT/nD0ybAWSTAY3eCjXAK
p9W5Qct3GY4PJ2+pUJnlwDioEATRfKFR/ZyFKPJrkak+G/pkYftj9Mm0qswZDJpn
yp0HrluGmGfOcTLH7DROjZuphId8904ywjXyk1eJ6Bel1qRvTZpreCNcjxgISyZ+
QZmRy5BvLBvwvPnnbPNCBwViZ6KaUvTwHRQJFDG4jk1KKw2YcXUo3WgfEq3aK6uz
NQbT76kuSTmK1dnfsJ/VQtHRW0S4BWVmuQCcDH97FquH4UZmiVrwd4dx6bWWh7gz
57LNf+AQy99uKIwy+jgyIxvqDrPCU5zQcrRNBAUX/3GnDxvxAXD+JtqCTnh27Qr9
mCjLtSlH0R+REtnebcun+oNvAHbGC9VU+kQWtFKrUXgwzvdXg/dvLhBPWIHXhre6
zO7SXZ40Y1Ucpfbx2qFAEjsMV8qRkHp1Cw0PODBILQQ6EkdqXF06ViL3xkKmuCUr
/9XAtA8jV3YntX4yNzlooCbV5ft/G28kV9MGUxG5zJVw/74EcHxS03hYl7sDspmw
BUodDEe1znSJ0hdlZns1IniEQ3DJQYb9jOTGzmheyWKfd6ev2IYiyZh1G00QBLTe
5PyAcuOTmjTGHnaQY2nequ5+/tYm7RHI/5n2P6bmGplIv0k/nCY+mHJUiaCWlQNY
CBqYX+WF9+5n5Kkli1cpLzt3IfLDkqMBgpiHoUi7R4fK4H1bRTo6YLeKuRopASEf
PxCCDYd0kaxl48pFjvk2cAW9Hyn+axUpGwr1WtmOdbJSwiutBUfLMhb5D5rUegAu
IhmGW6Idq5amSdiHOshaL8rGBRsNHfGcg+sVFL47x0ZS9eo9+lHjxBpLQcUuqkO9
CdEqPQMtg9pa2S26rWObD63zlQ+DC1+BatrBkxeYD1FoiDi3GUe/YxFhRc1WY102
kA1DiY+Xs2XTOjaD6AYg0YhbcnbYy5kqtfD4HajM20OM3A/DkHQKipoAqZt5CtPY
/KvvyAa1XAopxZlJVBuE7151z4UfYe3kpTgAJprfI+8UqeQGrhjwMYz6EFggalG8
tXDiz6lyNL60hAfMu8NWpANl5gYHjRXVgrMbf4X65o3j6upJbuEzDgbx9oSjreE0
Ie3LkMIQe5Cqf9+S5IBhJdqCwE/B2CsIJ5FbZf5gW65y44fRxVtPoPY9K9R7uiW+
/zFbq+9pciepA+735oWVjmsYj+la796L7eoXehZfQTuEtZqM/88DqPVs4MZawnrc
74ro7brAf/eDqvwhNMJmkXzFnY9rX2pxzdv/lghQHIpK24oslwRuQBKb14+6Ea54
bY8M80+tQBcr3YAadNi9i9NSpgKEG+1vXgGCFyxyvL8i8Rm9gHVnXErPUsHfdEf7
QpdDEIBSXBL5Pu+ZDjh8jWXCyrj3vBBQtK54WBd9IdVD5ltXGFLODkDAflJfsvmF
vQcnLA3X9JgnFj8I5smBTb/xC57V6R3XXZJWdb8+lYC7qz2G8RRv3ic66XCDpPis
J1soOAewSA4+wFDWYTdn8ubMDJLh15bht8Nkp33rKLvdbvLrxjR2iWbn+Q5jw6qL
5+XfnVU8pYNzVt4s3TgW9x+ahisgPaK1YvHYdoF0VfbkqT1jSD9xGvXM/H6KfB6h
dvbJI+hjNkdxtlVeESWZ5yQCL0Tr1Ew8Fg8WAsq/D5Wtk6OFAcc0vrYcg2yskOjo
LZ+NFNhi3Etcrbsf0CBW8+XiLHcQO1nyxkHVme0dIDqsS2bG/hoxwaH+CC5fc3xS
8bjZqBqtagI3jzCwg6jvhFWP2aTN9xoTkynVcGEVVpCvYDGTQVwp16f9TmDY1Hbc
kQcMn4D6BgzlGUYYw/tJ3LJIgWsQ1iPfDIi07qXhwl0vISImMwdI4cp7SBQPJMc1
Xcq7GGphzQYDK9QVazZo3mZOT6+2NnRBeg5DJyCEpQeiszAWEpzp0Vz0p9sAxeip
ixfWONpazS5GshUioXhZraQ/jh9AHwzsclFZNVw4t9FAgyiMXPIV8bFNAcBC3mpr
2Si+vJsemMxPWiMbG2+mzRfTOi7S3gOjK98+cVTtP2rM+5hdar2V0dEDp6JQv7Yf
mCWWEaFTaafrcfn9tMfFQm1AbCyrFyWoCXapwcGIUVavZzg0BatIqe0N4BZulrT7
bqAsTwW0x8Hc/QxkZNjOUt3ur1Wjr65SLIXJnO4D0drE24Ch6/2sNhM/JaAhE6wm
8kNoMvGUhGjuhb7ND6dzToPK479TFQqT+aCz+Lh2lT11FjOWtqSxjsJeG/YNHunD
xk+RG9jGw6w9mOGC3gr3N+MYL7eiiEmGsLVvP2ZHFgn+E6/gzk6itOqTb95cqrp/
T5o+oaA+dT2Ms0qAajzOr5PoxRwVaBHVOZ6jJb7xBa0TyI/EIlb1mfBLSyFuUfj2
M7tThfMDYeoS30VNmsZ7GwG7wQpev15b8daREOM5sGO5kv8JA8Ogq162r35xqIi8
7W/rM98Bi8d8dIS5SJRwrAxPNGEHkeBh8svR0CJO6TOvKrvAmNe+yHQsfdfAa7Eg
tPp1/1clpEy6WXQWcaw3M8ipJDBJCFlUGS9hXWoLwrMk6S6o8m9pBK+jr+kUDI8y
ggyYljdAYHU66hbUOyY00HGCd2NFmSzZ212Lipm1m4s7HBZ4IekAovL9xWO5UgY8
moly78TOhRhVE54v6FZaaAnChCRHRoT+g8JMazu9lPaRQugaNPFSyYoniwBPkKSh
8ynCTf2szY27bGPn8mGdiqmfLeb8yEDdf8GhGr6xvcvu2y5mKyWKn6XkWNCfSpNR
3+pDyONKaUxf/3D2OZ8xGc/gik7TICWeJt7cEMzVYKBQbpTS2d8sbEOsjNJB9XNm
wDV2ye2rnzqsuuX7H0ZnTg/aeFf6+8JGNZBCrPnP+WPuDXSkimpsNlF7GOYTesGH
T6wKxwBB8B773Mld0Xv7FZUeduPCnMm4+d8/MFJUlVCDwF9/pkUG87Ap9nw9PKV0
JJP8TJfqrKYbJOwPAjR9/ogX9sX9T/YEM7Ql5iDq/bZMF+2N9V6YAZP/a+ZpeMmd
E5yCUUNUy2XOBcML0q9zWzzYw4+3yTVOBBEnowJ13pM4QbjGhCiX5M9nitBhI+7o
kAanIz0C3CntVJITw/oixgclNA9p6UJ1d1s4gHrino4EqaXqZGH64hBkPCrXi+6R
rbrjkGeY5rqE1zRjtPd/ETAbna0tP4dfC+42eNJZoftEsx3dSw6JkP6y90PoS48Z
/2D0726DDzcERuNjsuCLyxLeC2H4jEVuk+Nj7PP6vtovRZoTui1I7rGGZkQbLZjY
UTYBtkq2LbEUvSbYWxmCuELWp7XEbdsmpp/DbBFL1ipWC+uvNKIA4YwVsyydnkj1
2McZ8VW8dpYg+puGkTnbt3EbdCFMzuK/GuBgOuQ9Mkg540r+hQxnH+4myKq97Axw
HSLwCl3Lvd650JjW/wzgrtBbHEKF4eOhX+a/3b9iKndDPCu1si+qEzgS1gf26+/1
HCp1ycP0t1x9btGlRgx0W/w2KdNfEsDJv22K/PzMAgQQdO4wBcaFY6NWgrSva+bI
DpZqZ3ywptHcqn8adjonNBbpapQ9rgjBhnJi2/Xc50tJmw5GCv5MHI49PkliUzep
MP7Y/yR/UWe51Kktzx7IUDgaS5bELUJDT2eIU3SeDmv1XyYm3fKmjnYncW6QVFuI
HCggXEDcYoc7oUvsmuZD3x81l3L0d8LuMeZWgxu/fui9KEg1BRxnT8tzA7vJgbq0
BQ46LsPdcAPrEPTVDZo3vZiZmIm3k0Re4RVFHPwvAK36PQs1O2moLiV/DNVkkeu/
lrzazurlEpJLUAZOgqus9FseI81OO9bQZi3Skh1q9XXZPPAuIbK5SykEFYSwTON8
u9CT4j045vvF1LGvou3SGVpVTOtIufOITbk2Fnfxy9da26AEZq5EgRAm7fgz/hfr
K6HUFo8b028L9xraw83bps7q1El5ItK6AuF3si6FISGoNFIgZbHrOrmk2Ad5TZmf
7kWazjMbfhhwGorimT/4uHJOxQzesp4BWCdI3gnbwsOZ8ZlSis5LL0BgLPsKEPGw
6ahucx4p/MmzJhSAIzWXArZjvwHvokQlJ4RCLPmeO4iFnbujICMsrjI+hUF7n98+
sQ4WKHe2b6obJXUTSMeE+vhX54xe6NCHQpnv+7Dh0fh3l+CC2QSXquJ50wvqJZSI
TBvgQ0TSpAkokT8LS5ObQCNhjsfRG9NKbmD/bXDtNc/2EsQpHDWuY5fkPSsdbY8Z
kahuxFtrovF5Qmrz+GBq88Q00fWUsZ6SvdXdsq8P8emw0OQokhltIurx93XI0H/w
0zSOtP1xaAgPRIkK8P3C0ARzJ4s3KV5oU1OXwcDT8Bmf098qdu4JwF51YzDciMtE
/cyLOwrl1ByV00k7rUZtnWwZ9udjiO20nhq8iYEjy9yGytjd2edqDVm7EDLm//63
/SuJiZkMByosNIEAxqqmKaTHQGVxIuLH8u1gvrZ94tEsfG0mQsW2emjhnD3+69/X
7go9VpPIrf3DdpAEgS1qml4ha2P1UyCcZH+HECdUOEBRUWoUSfmZ8DE99AfXjvAL
VtHv086wEupJq5vYOmCQ/nfqxxbeHZ8mZmrM7qrPufsDt6KLkf9SmGV6ZDaRwXud
ji8xuU/2VXj2cUaOdnIDP87HKqyPbqvafwa7bvqDV7XSelUb0v9npZsLlT4lhIrV
1LrphpRon2UST0zxg7AOzKszirtAVFn/ZWqFdG2mpIMsYyyIGthFdKcpb0ffceZn
Y2ADK0OtJemwyXaQHQLLwkja9+8nLpwLRWlRdxhTo3AKetjkeB5PSJyzDBLIpICk
ol7Ao8OcGub73KNZg8ukfBuPOlZnaDk7HQ/3PQvSIPVaAZH+RmrRCM/2r/uooj7c
txliJnv6CXVV94SVbJCJ0j0pUH6mZISW2ne8DDR1/KaAr/JNsvW2HMP4dJdASylu
1i0vvQm6bOAQlIf2deMoA9B5n1WQ8gVtCMR/Z2mGo7OtsQyW17owS5eqavLuJC0y
ToRC5zWQanQlPcBb9E2pIcxLO0baGci7Cw7LefkQzQl40IEmgs2nAJoTMvmwCCBe
EF7P2Nrn7qv/cL8+kGZq8hEYF2xzSR+LHM+GYMbijlI3WfAqX5nygpIqTmo50O81
mkX8TqbSVz9cMTUg5Oh+heQBRX6nyX7SElCAA03R85hqeVokkkT5egvAqYOykWvi
r3X5q6wOlZkSkwSwfZJfInAgsDx+yl87eGBPBUHcYQLivyESszb3ST1XHFS/j7K8
GSh64V7im9m8kocA5u+R4BlmMN5/K3ceQpwGN0vGpVxbi+OjmJMRUFbL+dJrH8Di
ml9uYi3inGIolvWRPYcVplF3GiCeUntARvt/hyzdg20WGJMHHWpqyKyl4O0bDGCB
gDg5kKqCJ3N03QJe40ZQUCeBq298czeOJxA5aqZGWwn/ghOSYQV4oopLF9AJKVJh
BflqbXLcDOmZV11trecu+/89d1GNqUaDX021/E4mEPO2I2x5JADMOiAu9qRrHC92
geIl3Ew2Vlc5dcRb46Xafo+P+5tgLmGE230ODtTN93XHebW4Vg8pvTy6Zat1IAEc
jO2PpQHPZRzin8sH1KroH4EFpHtbF8dEvAX79HPRAS6IMkb5YU6u2J7pXczO7ZAR
OCSoo1aJlfH+UmoPHIiDBDNR+tZaRbkgpnlDdBJPnEqlFrgDpcF5jOkeagkfy4wV
2b8E4rgp6Vzv6s+UyjTl0YG7eeXPEHav8ktAgVaw5HIjmnicssdgQ56LPNCVvqHF
T1o5Ek+O3V+U4elstQADcWtmXpdKXkqV8Ad1u0zn2lBYh+c8WjASglsIZe2e//Y8
JA++EnooiKBVYGGas21ksNOdI5cnjXqK6RM7F26J5a3DI2OAZTvxIW+lrDvyay7G
aAHjH1Ugz8lRcMrHF79J/1xDzXGQEGUxFX22CKlobzYbosfgaZQ0vG1xEfao5mlU
ygfV/YoMV+BSQzAUicuB8/KLn8BCS3IbZYIlK1Wp+fDnccecAVCITWFg7SU08bFD
lUisFnAtC/YkB6Vxxu3ZkbVJCgXG018cZH3fKX37j7HIPR4HzQmrGhQvVRDXOdid
kIGlruPeAXavm837DqD9b43DpADK3dH9yDLohkSsWGRB5VOGAj9i7A1ZCuH7Lafh
Ul4DlCTPPMjWFs9edLoNtqth+fcd3aGDzwuia9d4eOZIs1iXXedX+yA/zUJAwqmD
eud6MDXCYpntcYwEEDRX8QOoQBj2QWR3bcdH4Y8ejUIvyz2sBE4kxBnPHtcGyC8Q
qg8xkJMl9Pdnjl4vbB9TH4xTiKv9eYOz9HrE2hS5iyPnuYF609IhNYpOW+0MkPGj
e/pM+7Vdv8zFwPglYU/qeqJLwme/RGjBpxCjs09eqDYIgcLD4D5do+914RSmKj5M
8c5HVENavh7oQvRqvDEn6tuj1c1POTc56eEHGSOesa+Gob+O6X5A20WxQqlrBqZj
wiAEHAMAX0FVOpe3lNaeuvSXlH36XCAEM7HJLwqMNB/IrEvbtmtXDxykdIup4jlv
FdEulnuU5q0hppdtrM5uiG5XuyH0YCC0JbSpYyPhOA9KP0uBD29sWCecZuZNvT/C
1+7qbIP+hrs1TS+EnaagtCX7AC7KBz0oWdDXWs/jNKbgPvrBpm8EIfDwNizPzYwL
bHEdWSAoKJmpTUz/OAksNdpnwxfrbcdqiDPYkoQKlz9m6RGP5QjQNlRNQQsu91tx
yIOe0IIiZrPIQuIwQqPNbCT8RREoqk/ziUd+uUr3oXA5+LNdg2ljbhBaF3Wrbp9P
K/LlkPHWNv8jqx794DbQBC7vf9BbWTuaVkbVYYjXe3FJ58gNMjmhdeKlx6XtGgcI
rs17T+ahiwgrM1p7yplk0cml0yvfYvO6vXsWbKHR2GZOnqsC03hyxRmZGhV/Fke9
OSXg1UEDCngCJmzC+EJlC+bitL9P3Z3sglioN32ezWR1PU8cnQyeNC2/zYQl7Ehv
DclPVuLZoaaByHc1hZiupL/LYYJEM6XTkH1LyzbLNRQ7CcN8dQUyg6o8JtMmjd5t
ABC09UjbVFNxjRDyy4yduB5S30ihfMpRckRjzOJSP7z6N4q2h1GNnrGHkhhBOSb0
qZq4hiaVcVwxeYyQX8z66QiwUE8rm2AaURph86eB1rB/Wz69+TLP/qQSaH3P69f0
wgGAqoS8FGSn3l63oXhv6s26heN5qwh1aF4dFe2+AkyjLKdmoPOjXNLxgOKiFMbl
yKjV4te+0QQ/PHn3dxHW6R5hg3qzgTFuwX5xVT14o6nu74+niwh8nWkWwr5koQQF
0dxE/Oc0f9o+BCY7pwZc6ng7W1Wg4xNxEW0ys9ttncP5YHilvPQEROC8xIJtkez3
ni3l98mqXRvvDwSIk2ccQcUdY3Swg6JbNi+mDUvhCzglUVT8QYOq67OhQ6NSpLgq
sXnwzNX+DpXwmZ2rzQDs3R/Xm8y3hgJCVCrZFexjWOYMJCjZX46KRNTeG0fB2sAB
yic7e/+zR4/+ojf25PFsfcNw4kYohZE/vIafoI40qyFfCoCxrvq+LrO1GoG/BxnJ
G6dd5oHQ9b/r1WADXhruTGrr6uTBhCWoxY57yD6V/mAXEztgkIkGzqiWOebWs2nC
3vwreN3MhOEKk8hhuqKei08gg1vdCU3fH18u/pKvDZUOHSOBOTJZ8SdonHj5Z92i
SD5jVaBibiRttwKjRk8nJ7jflohBhMUrqO5JtGIlgat8zeaqdAKbus3irlfvueiM
MDCmv3k+nT1VcpOR9lG5nyxfM2b9n+t1ivb8P4hihTPhyEneLOoqYxD1filAQEJj
KSIXE/RVX1W9K/xsA+ndpF1bQdMsA/CJnReJt+BByZpJmfpKPpYbrmnjWX1/hrLv
tyCVHSK4fD8R0cwI2ADT/TO/J5wRR04hdYoMLhSTUt2vBw/1AWCN0w5oIL0aAG5c
Fqi29HF5Tneeiqa5Q/LZbOhVZbBvBNGbgLaC+P4dSzeh34hQjccijjkf3WlUvhOT
Gq8YRHG94tBOAVJx+wgIZjWGUGHHmHhkC1fvjj6ZKP5qanHc0QxCgPfJWemko1sR
fqsQUSm913LQy0WIDDcsjSn0JsVc+Y+zdYCLLNfNswgFZW0Y1jpLsCl/V2mJTnwj
M36prasg0km2FjFHmWNArBKRorQXeL0gB5tnNNqStGkdEslc1jQBqgIS9KD5obGe
I8Y+rlIYZO8eQbYwugiSguYlZJQjZLJcVYwMnrKw3+S1BERkhpwfdtEEk0ugEz9+
+xH3Rw6XecBbvy2ZTpoDSr4iFXgzgezXXO6w7UHGyBuH6kebd1XBSnXPJ7WTqTkC
NtbwdhMD5z59icOBv8Jqd6/m2QbJJmwjtfYIed5oIme3MoXGlgl7HgqZTTG3KJm/
xzLzBc1FEsU4D4p7JPSZzqPXezT+9gkEVesd+AAQCn3nuhz9UbdSLL5AZhv2Nu17
CXtsY4neFKUUPZUYRnT+Ll7ydhy7/JaimovUS1D2fT9f+NXl5R2Pjm6efVUy+4FC
BRT8jveAU2lGN6j11DguNq3aEGHvzDLgIV5gJ81A0bY=
`protect END_PROTECTED
