`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
znhG3oZqyKyqrwVrtI/h5JppEHsCwbV5Y8SvMwca9XJreveUJ63dZEFGEspp9Vit
Er79doJYX3FiWRQ4LpDItPDg5SUiL/Ttu/Z+0QOtJHn+5UX5Cx5akHG9yu+pDSwv
5BPmRvyVnogFi8oNTP3M4ygrh4Sqfs1STsjD7WQPToelhhihvSxXbIT32pjXG+sO
GYcp+mrI3+R3XE8BHdXXnky7Tu69FJ82PDZRnTNvQNQnce5Y4DWkC0m0xyUYzSfp
QyC+MzANcVMT1PzLXBOmmsKWBQUBi8lky3POChm/ILJgTzucZhUKyrfyd0+R237n
7zAa277O23SXOizbZkXd6Lix6OfpdztUTk5j+BHco3kMZa5ufYoKWPXhMGlxV1My
oj7vTFgl4FTonIfXV3YXRSzXmw2ZxligBdosT0UtAWRIHh6oYVjPCptigSsE4JKG
Pdfmusu4+cBR4OjICiR54Lix3VaPEDNdsMRyYZG3Wh2hYOLJ7jerEXZVLGn1Txj1
1NllvQO93uE1U4tKYr1Pp5go7DJeMA1naxxVuRELzc9hi1Ii5XFuaVL/sxZS59SU
GPav11LL/Un+u1HnMD8biGD0wLwOgmqfAgd6C0EF9MB9Pn5+FY6XEn37ySAGOtJ4
4kKJ6fGz3g4v1O3jxV+aGg==
`protect END_PROTECTED
