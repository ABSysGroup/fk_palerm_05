`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BQfUcHBNZ5n3giaXIV1bSHa0p2H61dU+zEP2bNvEVsp3Qj9oGfzyALWd2kPlC3+I
jC8AIPnWrhMVmQeRfHg2RuwznjZML1pf9R4557ktpBt16c1jEbz5M5y1KwjXGbmQ
F+g2X9KntQ3rm+xszFNF1M7KdbRaW+QDyk0olBZN6F6g4tO7SOwqNKy94REgXuCu
8sBWoFoWBsFdIXKqKb4LBG3L0Lw/foQDO3whmaWxpLtzgxA7UN3jjM0+7N4TWP58
U5kV1aCjOVTmRJRW+XsJoqLR8Ybm1Inge8cyBX7Ua1t8aNZ+48+asfTEYYnuv8q1
V/8k7oMcTdbxmHVx+poe/MI+8CWpwZtUWEwapTdZqUAqxG7t/kNc+kV85pPJ+rZ1
VbDL8WQGglKkbFJt2Mxtc1gpH7E+GFnaCUJU0D79c5I9lLq5+xoXqNCh5OcbaE88
rcu5oEVY1gwkqhaKB2jDKD5ZIMi4Y+WC2cnZ9PI2nEqXr36UmjyKG6nu7OLC78ry
ck0VURvCqjpRFxOr/+NEGV16hITlyFdEXsSu+iTFybNRcG/lDoN1JojMSMi0ZrYq
0R6QjSyTOSDUsx6u1/qxrhrenRBifzpo8vZqTy9tUpEGFgt3rdBRHdwOU5BDOgWy
EiuYvoX7XrKPLTrlKu9au8cVQ3AeYRgEohFa47eW/ZI=
`protect END_PROTECTED
