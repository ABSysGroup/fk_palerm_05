`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oHQwCyykS8h/7A1WXjaZq/g/8N2osM7R2R7GP+7H6/xMEdeKlFXFDsiP2SfNSpE/
42/9cA14Y6kvURIwhutEESUzbJi/tCAOOXmpvwCdAIxHAKuN2youQO+xLPRRV9ox
Im9Tc6eMxX2+6+uJHIdCbgkPVY/PGqBuj64LK1gBgmKwZ+6DNbUwrUev55LPQu5d
eS5el+Kz5rvRmbEyba+QhcoOXI1T3D/W8ZkSBzYeAlwLsHA2UFdjaLm05HLxcz3M
BTESIlLuGqtp6GM3yhklhi17R7OfsjoJwt4Muv9D03SzXnxab1pw9QINqSSPKrBn
P9kx7FXsm3aSvaV9JoSY1oXVhHeAOMhg3hE2BE3M6nVbo5IUYBhvKaSqvaSe7hEU
`protect END_PROTECTED
