`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yXHw8CN4FqJzadM1ViMMdUrR1HXt2eD3szXmUNsUNSpUDNoxxCJV67SWgTiO5k8O
m2z97G+6CPieTCg/cIO4zMGolLSGVkkDju6pU5pfjCJVnRTbsW03pnkikojp9hbq
ygw1NwuPL7b6XwojGSMaYpKHZzIfxrJbCKirEbR9+UvEs9MDDmRyNMxKExCDbtlw
ppAn3ni+a88xbE+Te93c2WPK4o4m28ybxDYplRlinGO2ZIjdCt6AhfZzus9pr4sE
BxbHa/kNFHdTSfF+2snHqUN2QwNGx7/dw1mk9/kzxuMbr+sqa3+98UhUrn7soB3a
PaC300KT5+HM9nCgIVF0/V9vz0GyFzPVil/V8X06DQAxu2wCKBu0Xd4frSiX8FHg
UCbiSav6Mz3aCtiV2IvDs6+BWqHUryTJfb0OYWFN26II3olPeGx7/7Pz/1LZ3FFn
AtIzjUjYxwm4f2UNfKMuCA==
`protect END_PROTECTED
