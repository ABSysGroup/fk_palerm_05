`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gai2fbkp1BJTjHdhIQxezEPCG95vboR//wtVsaymG7yRb62H6/aEHXnXf7KSzI1o
wxtyUMyUVac8/5eys4MXWlX/BX9asZy8TZyYkEz9eH22l2U0jj7LwfLSVNfiirCD
e3XM9DyWnDaOhuvMr08UTRbBFD5LGNkIidI5HkYVOPr1n1xKuQq+5qGMM7NSeogI
/6u8UTvbDFJWek7ANaQ1qfiE3iztOnina1jXQbQQSsA8SHrG6voHURSOvbVLWHnj
xTtBifMcDXCLl6JjGD467DpOubVDOVYpDl5Jaw7gtYergAC7t/cX3vLkjWh+GNza
4q1gmqwAQ7D8RbHiS34azCZ5TTmiGc7taBfCu5W8pbjR3xpR0AcFZ6YgdjUC74R8
9c0RiwWV0NYn+QJ/V2/vdzWkaYPiB18zqyYqlcUVEqjQzNo7W9tS6UjFTqOFvkeN
z6wxyklkl01b6UT6vNeCw4zdy8D81NO1Cd6UWY+FOA+BmbVTYm6rnZGtsJIhJVra
GLEAz/vN/SpeGw3imyq7sNbpTRR7jujqHXs78HlT61AejgY7wNMvQRlidI1npHRo
vRqN/hKlyUQZLigzbiqi+MNPnlSB4+GeJxof15C+uEjEqf+LzvM2Hv7jxeoCkPAs
r34FisvTLLUoXbITGbTkke7QK5he7qwJES2QXpRU4eJjM/nt3bP07Idu237/4Zr9
iGyjSzvyiRNQFsIIsrzUgM9dxCaKXLAL/X7QM1qsy86/yZlLO3I7lMwt4cHarb9o
acOG+h1u/QS4QKqJo2kuuKdkn5CFw0ymgTttJIX3u10GTi4uXjovg2pgdhy+3OI5
PPChy1Ihst1LkONEIVTXcGv3Vr0Vu5T+UMjCZkY0hlmauDHU8qGmwN0ZzHLnqYOJ
Ce85HhqsZ4GxGlnULpU3lajT1RwJtFe8/ksMoxm4L2JMReC09J7iDi5/kq6HJ6B8
ym9KIMlJsbfWyBMJ51gjzYSpwQVCMXTzwsG7UjS6tacJSvk0W2g6Heu2iO4vCrEi
h5eerMC2M2aG/lv1BX9qhLoUhlR1TThyH4xu9jzbuI60w+TE3iCwlkFjwusDutHW
cjPbxPAkurojEvFc0oR79ej6hZ21YipFQ+TiikwZWPG0RIQRw7k38jHrum1fiQIG
3My9jS+wh5Mad9MTI80yJS5K4XabWzq7X1tnGDjku4kZUL3Fxxx0ZXXoq7OuVA8I
qgTuFOAj9P7pAAQVyqsYM0hmLG7vss0xE2EKmeTJyZh71ARrPZQatQouq2/Hur2r
8kCfzS1jNZAuiX4yl8AHQNmb0tAMQW6iBeHwXeeC7xDrW0BnzxXNWrM18k89Q9Zs
UArqNMaIkUX5wFnjx0iZ2NNxj38nglQhgwhaY31TuQHhxRc5iTEYbULcgWvJlZrA
PjO/s3F2gy+Gf3ALyKq21HsSdllhNhT1/pMY0/qPFblneOZoPs7Z0A/EcLI5jtiD
Gr6DcyZ849rWtkKP2oJelsW3BWwy5vT3xnEpim/vqKQQFU4Qq2sEvwzF0E3tfx6k
G9EDFD7P6P8Jy6tytHA/gMqafrhDZPRGmTnE93Vkjf2MP//0G/Wmrq6LHs26m3Rb
kFN3gVZQzj6QUmR92sVCSWRWU7m1e4KUjZAB+3f5N5HYvpOkiCcZ6lWkul9ey3In
/jO6+xvqv3vG0cq7X3MbMeMYXwFbHXusr6+5Vzxh1ITEZQ9zU+K6lJP64WHL5Cng
nvPYuhCKfDUt4envURm7n0o17M3wxMzvhFdh4MsmH3TqT56U4RrnLOfvd1AJr8JJ
Ctesc7nqYTvAJbjCzISvTuIhv0dy7ftLbbYrmEqVgCMCWStevlsF5NRajLw5lmmH
RORCQJBBpWbINLRNkWEHdpdXlfsV/4XzxF7QW5mURLMxQqQ0yI2+jFcPq7ToScj6
0kDsCYm/fEKMbBsGAJJs7NrTXjhaY7M/6+AqFDsEiL2r006xg0HsscGSJdKuGzPO
2mpM4WWYc9U4/XYLTlf1pSsEgy7YcRWIelak1sisF2s8N4FeHCvPZSqjGHq/yQFk
fStDpZl8BVMfJStT2SWKJ3gtKvCqemW4yAtWbHY3Zd3gAKA0PwE4YcsKCnTdPTIt
at3TY0MYP392a14E8E+AwusOrs+mLhL1hSySYC2o28ab1kRQ5vaIt2vr6jdbxLQ0
jXWqbfFc7DzuvATdiOshCjFcvnxpv7tbWlkpdOrNilgt0qLwd4iVJw7J0g+yX5kw
krPSZNH2IqQEV11dnrcKiIrHm40BxuvjybdK+gcSTu1zs6kLMTe2GGZ73RQ1t3Xl
jZR4qxBTb8wi/zb4LdPTCUos+apsJo3DIk3e9GAFWgO5BXKI43G2pIi4ZhrOa55y
s1iYCdDgC0QAiW6MKcSn2M+TwRsw8YXYlwykfcb1Vcy3OUiwATXVFRDMIZeV7LBo
79MdESihut+7/abtG7BkOFBOlWHt+AAHmSomShJv5S+AJ/5hiCsrPyaR5fRUxdbo
`protect END_PROTECTED
