`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pcheJsX+nUDRrbA/qfbpjMhXIjejXuLyNSFfEAz19G35c1gQFvteiggmOYZnF6/i
OQrWQj+ldiHFyhzmyOpzBJ8Zzm4lvPC3ZdAAxeRs4rlvbDkiJSQBhXVO3hOIq2DC
/TKqM7EjxamZapNYljIyfSlSSKPo+QPcf7r68Q/IOCvTo7BPUruLWDKZ/AKFu0RP
ZTrMjqhkD9PL7DFP5RyFDTqbll5elov1lEflpBS6xzmpLpR6qOPRJaCkgdYHBjTP
po4643C61ogLMIteU/iSC5/NtEnbtzafYRsgch/lSYL18wZxrbrt4P9Wb6Et4CtP
WPJS1dl3mpS2J3UdSp2KCbo+wQKoUUSjvBzskaEPNniEYxKp/rzvy/wuECM4DLfs
xU0ND3pjJvaBgkkKwC8VrK6BAbwKjOOw2jDOiSVdCBujoe3VeNAUf2hlbVeUUzli
p62I03KRJHcYWFOYFSSj65cqsGu2NzpHpektrHSzl8ajDn49GT51DBuXTQtqLobT
GFKlqDsv/xhPrL6w0JCvek74kEJbzRJ4QQOJ2t652bM+AWy52Ip8lBsXJdMFqTD5
dsW3h04boapnL2h2slaV2HF/4Z4oBtNQdQACchaNZOUcbD65ke3UX15yYEmUz3UR
bFwtz1vZvpg6U81TnHkN7pjrCQxuNc4beyQ4/ZiAbeNVbVbl0hGLMKRJQ3u/kbeJ
tXdrXPTWUhnmeEIaqztOHlHoMMmlsA6nVjaB3cq5F4d3ht6W80qdwa6HKvyVPBfh
8SXOeRRB941jcz6BahhaaVXuQETZrjVFQ5uHm7ql/i6yNfRqKMLE/+zT7jqSf9DO
eTuP29qdpCFitm7N2SABxe7mwj2NLChLJVnypgjN5t8ONiZYQ9PoNxGHar4YofHl
T5zjQHoO9VcRQv0H6M8T1idLV/whXhIBNzynB5wgZQ/TYjhNQeNxYQTXiGmqK3xx
dTzGDP6M7VfemRRuGvLwhY+ZU4AHkmkuY1AQ8nKaSaL/e2bZQdUxrgMPHQirC3yq
C0ppDOSHYRDP/rvzZMlsDspNA7rA0uwo6qRllKBu6wljxM1XaZiQzvaeV16cgrEt
eHcrkW2Ug75C3Kcyos+kAs1dgHrgFwKT3FWDo4OEwS13uGFu9Nwu1k65Nd0FJcm/
LKrjxFz/Fy50PdGD+GCY67VdPDPejkfbmRlk4mYhueXgw5aWV49mgJ5zNCi4lEiv
+kAczGZh+6Ie1cl3rReLay2r8KCBnQOlOKZHG+7qhGm3HregGiuY6o25rLbjlLlR
1gqUapHO7iCd1tBnQAph3FX4wDANyhX1sgn7p7TDf7svuiRmtDrcO044TWdTvoFu
VRJZAhAG9hOqdC8nSC23NtPEUuHnE9PM7GQBhzdLvWTA5hD5ReA/uQT1qJ9tz5x5
X0JeyJQqltxLJ4YerHxQnZ+ywuvLIO5949zPyKMW7f5R1aOeBAkK05VBBF4EXku3
3FC5i1AlfFGHPUOSn7k5TWmN6+q7PLgZNzKnAPv8elxmjyJjE1KgIwbOnyqYT20w
OCq1HuhBLiU50e+jLZPvyX8vuMQq2rcxEI10pyWz5gw4gN5XyrY32zqoUXg1rhoP
CEphXYtCha2dndGlldXZ625aXZhBWmPw+4Qq8H+PvzgXJF+455pcwslZ/7GHq/jE
F2h8YQdOvOvgc2Bwy8v6xwpqAvGDv3YweBPvEwsHFD77bcyi+O4NidyqeJ/os4IE
wT9NUbrI7XK8tnBbhJELzR7nW2YoGQWJCYY+KH82d3fdCXbka6cvdk8l7OwJg0Y7
XlNd5byLrGRHlCouYBQj2nfqxbMQqqAhfQ3WyEQoaMtxhTxBnIpufCJEzGOT8oKM
GGCt9uWHDKdN+vrI1CmYQHXAE9w+E6iSdCBPLn20lcvXRuDU/wa2sD6Bnyy54BZS
9CXXPTWEl2JeMpn2SCf9k+8/vnwHMwEaF2FRmTsUBdBjuX8tXJaPJMJnRrcxV/V0
CGkMIosRMgp+K+DXkOMnik4HwVirA7WhmQaYu0Pxv8hXRhH6WioLl5Xs0kiJIf+k
57pz14GMYSjPrV318DOGFfGE4/jhbbcbk983rsthyypK6YbglzLZuDdFt7uwYiQ+
WVhsYYSooDsg5XO53RIjPAGMIAdDSSucSEVmf8ZoXDr5ibRj26P2V41bDd+iZy4B
k7lPqPLaxP/14yh2ky5p5XA6joBQvWfS/ntMvQIbws4fDij724+K2mMLRu6lr53O
IPv/P/EXTzulB2X5Els2el8WHmxdqjXaal1PB+Gnmnz/TubB1LaDiHlj/shyD1ue
EsjdXCCNGbQ41qga6VEdFarTHAaW91qKPOtn8z7UshhXKHgpXEJeRHy6C3ECaojc
ayxWmfhxJ1MJNhTbAchKJZHTIXbwKbWTgXzaf4YQN/nBhenYsVg3vF/5P5+olnMc
qyFvvWvA0EC7buhs6JDmfI7kVt9OBnFzftoJOASZ8DBAmC8q66uH2LL/QBJrIVFb
7QuHsSK3RBijsHpZNqBA+GRY/R2qxvoWSYCjhkKcYSAWjGOdEZ6yCjIwIURQKyhi
2tSmSzzgkt+WnYPkpMfnuAQUv1D0mQzA/r2ocSKEqYbgUleUccTNDnuEAmjbYdxy
BtPIN+at+iKQLFeuundau8kJEZ+JdFt/LrQPw4PoqDehNCXKH2PqGiw28h9Ei6hq
9Xlc9/Xae/wCoSf3V25yZO9Tjn9EAmM4kJxPilUOFj6kXTkfPkbJCZ9ghxT9EvyA
O5ATqiPqr2XstZ2DRKwrYLeifwVwXneJ2ZmorW98ts8wgJc5SS1YB6KskTJCbfpy
4CCHjgciylTSCvQ7MxLqnEg+45VRi73bjWwci4J4RdMdYm+Adp1OPwXSOf/y8lpD
OiuTjyb7LGG46AVjFZ2YaF36YnLbrhhdwxPTcv4wghXaGlRwtsHghubyyFYF947B
OfcUCNtY/T7LxAyNw2k4ZLIgt0DvPu1K+uodN1/P/79KYvb6vSrXEEmy4g7CTDMK
ZldWFW1bbaTpZswZhihFFOXREKJqFdiUnCl2GVrVZ6vKbOlbEevUHsUIFH1kKucB
XZ+zsOkPIEf7LtgBmoUU0LGgnGKnUFg/WVKpiCS5Cc6d1WJOa8FSagE3DEQPvJx0
FAMoM+I8p3e4NwSL3Up2SeCxrOI13TB6u7r6jk+WaOU8Fs66xgzN4jV8CgbLN1+n
fmp/wOzSkls/J1/a+GC/jcUksR6dVUAQMqtgQFs8lKskJbAR9fp8E8BMGRB9PWXf
V7U6o8MklaVH6koTGCcWqu0X701u/vFU6wFUarsYy1kSk6fE1/jHX1WNIzktg3QF
lARaXrPqeXXO3xFyar4iyfuSmeYnD+c2137OWc8v9HSfLRP9kC+eWSo6lRzYdhy3
9PFvXhd6touDS+a5XEESIioFgJWrhZ4S5l6pX02pLDOiBaMKhpoNkG/Fab96WgHd
vIxs2OlduQWt+z3UnnLYLon3zwpJC+lxBVYG5ox04C6cm8+G4eQ0zKE3I1bnaCOt
LPDq/4qRY/9I67RZw415SLWN4qfi1M794y2On0ng4pl+A0QjCgBmVMPUB6LyFU0l
FqIVHeIpIWHXLeJPR1GNIZElyQfWiWBgekLcfhiTzG6f2GJ/nHZBc0O1KbGcwz44
0iFT20SvCQzD7Edmw16a7KoWTUnGfTEcAZqhfHmJ+pWteoxIVs87JWCesymw418N
TD711mz9WpJB6d31lqxfxgTLrtPEIFDwyW5sly150mtMyeLDONUyT2VJ8xtMv7RR
9pfjU3imbaVVzvIVpp7wUF0VQR4wKHdy9PGpmO8LC+4dkq5J60PH2au94nhNUpJZ
W5rucOJgQU+614NWReSUKZCviM2F0uM4980QpUdf5dlVNeKTS6WMaOZ4cxbksEcY
J5q6ruqGiHQnhwTB89Dr+Pk6tRLFHVTHZU2EOqtnXth3cvBynufmjhe73IAx7xs1
hbAdE3KVGi8IyiTlwi+Thv9iuZtLdFFfj0KQ0YApJOGEmUKbKp0rTwDSGX8Aqd/I
Etk8Q40o6yq0lyofHTqzwEieA/XtbMYX0YuXpZ3/pVFhQ7xtqTQGSmy9+S9UfZMJ
/qLbH1poqKXLZZYoyO4a/mtWyvwuNVSmvgcZH5BPqmBLDkb2pJ0KdhMDdORtR1u/
rsCh0JwH07Yx8iIxl1UXOF8l2UJp6X3OW3cA3fn5Ws9md2m3vJgPBLyhHP0Qfnvc
pDx9n1t60mq/tdBW+GEu+BrqMyY1Jd8bOWcbLbDN0oxXO0Xvm51liQLfsKHoDZWV
l/4SgTc/Lkgguc+a7g+uBl+nqXoxketWsUDg0Tue61oJ04LZtcWcbTeeCzQOXwWP
6GNUa9fZbGvE1ZbIiQT0XGC9hYXnA8IiWhH+6SPdHDHNwAlmzBLt8I/PkpbSEgNB
DS09yOCKnj4byx7XXJHh2nlGJpD4kxGpro16fX22Q3UnpZSpOyPvJ4Q3gcjDSfaG
gzUuYFA5rbdsbE02yMsF5Gdy3NCiUwjGEMnEBhi+iNEk0dp2AtvcVqOz/RttBFK8
aX+cztqqFxfP+Qa0ZAFs/ld22EZOedn7uw8Pd7MMcMT/TEzpNmHOUNCu261LuMd8
neUacmdkDPSjpH5+j5xkqKHuuYVGqrtbLDEtIDVvLY5d1UwvLCMkQ1AspPGR1QaO
WzG4a5NYdzeMh0TBNXV2sMpb3X5cZjHIYX/+Gedg+mNZXSWh2MMptooDwObhCx0M
KQRW55aTodbf1h3/2Zv4fMXC8oskKZBuyQtnhPPYncvB3PXihv8qSLhw9Akh+HuH
PaxvCHACmUzBkLJBYPyODuzKm5I5aAEOpulUgEVtuS2JXNt/CMI7nzjQA9fe0AWY
KAkD4tPcv9CWFzjCN3UTTculYFPYsN+bbnRylQ7Ce2rMDzp0rQdKRT4eCcQjs7Q4
EhW52duR0WrNTbJMyqG3QbueSpwGYlx8nt4TrZ1iJz9qy0qI5+PVvge61+1Dw+5m
mPz+FTH1OR+D3HvPQwUGTTqKYc2QgBYBsFhWctvU6zZ+UT9/qLIRloAm9sUjTR4g
LV9t6KVylE8osme0M9Dar0dKWMmAJ+XOIkAWuA+5ZCdTcKY0Q1pzpaDPhUsE1SwT
tiPFyPyhQ0Ytbkc2cumSius4mEfULF4v7WOk70zLz4g0kisG242kY8fD1+hVCKwl
lsaMkqsjQAoOuy8EFfD6CIL2jvFIpT6prqrA4K3mElbo/JX7wSaE5ijANK4nxRdH
VzbhGfbt1SwfBLy7q95/lDRggSjYNKRiK1W2FEr0tVGOcwXkpGlkcQnjQPY3hXbB
V3lny+xMeqO/PmahsBwwEv0BPwhUI0mkoPNqAnOkaDyEK7vt/l9mBpp6Gjr1B3aD
wL1TNH3n0Rl5HjAEzf2te41W6WQmDKGLXD8icPPlh1tmnzg7+vYunZxrz9VtULOi
7+nogUf3vAFtBIhfCulfsZDizuUdPelEP5EuC+oIERaN+Q2bMWTrX+p6dp9VDiHr
6/Ni0UV3dzw7VnpgTuUz+z8aIlPexlQUIIQJ26D5/3LQ7SlxqkspjqCog0Q0a6U8
TueHpgOB9auY6M31KroQYOxhHtK+JUNsmdpKz54NrqlgnUa/p4rgfKl+827OJrMV
SZROoww/gow4228B9uZmoPYhe6DVusjNLnSzXbskUROOe04zhoYwDx0yy1TrsENb
5s2m9zlPIB4/58jbBJDVJRAJzPJa8oEEdtc5A9FfLg64/ibc+evOq/IKz1v61ebt
1ebuE3nDqxtJVcsXJTRsJLJeCEwRb9tbS2IkVS/M6a4nTbrLmTPrCHjkaAeGMUuy
R9UNYlG5rfa3EGfICg7C8yZdponT56zXEyhX129GdOFzRRTukJj/Bhp+Gwn3u0H8
q9A4K60El6vgaoUTJYn5hVvr68pEROLME5fCHNBpML1QBaumeesQNvvRy7rLq4Nx
f0I6/eBizkpT6gWo1rJzDF4mVJpUWpI8p4wMkjilxOisE9IE4OIOHlN93Gf6mSaD
ELiT6Ge3mpm89b3Zqai8W6ZjusHOMZVH/+3oaN5mO9XxHtl2lkqcRYhRnahyDvOW
ITQmFlgMi279aNf16/GsQTflKCINI45qJYn2eBYnWzt9n/exXJc16t3AnKojq1Fi
`protect END_PROTECTED
