`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rlG2tFDkIehIWaZQvIejw3Tt0xxdZSI9omuojLHdPg1cDVLaWkE1SfV+9Ad2LBMW
tNvawmR40PHGBy2fxE76Jq1pBY9S/nHWZBLnFM71EpuEN1jPgkorGdGS53xZkq5B
Cgh8du0Fhb2yJEQeIVVMdzin9OSq2lvLAse7HdsIK6+LvA1Bpqlj6YkWEjTyNNlh
8bH8YV9BCB47zFXo2P6U/qZcwloLQkJKBlw/+BS/c11PQbj+EMktVuj/RoMsxvJQ
HIVO7wwWsI2PzaHZCx/oE3vwph/XinrW6MQXhv+Z+EVc9RfTnP96xn1PFH9FqYvi
sQ7lffB3/7dn2PNf+8qoNb7ojlQVnr1KHhkcvY5IxbVouUJjly3PouKDObFYpsD4
HQ8K+0gYlp08NAHCgPmWTsaFLzil2zpHFGxFf3/M3VmAYpNEcjwv7h0quZxBBkBd
hoRpaJOuqQlNKzx6p7EGDboTUKBjQSQvN2YxvlvNe8joYmUWoXOYA3Q6e+SC05I8
l8fCAx6I0ktGmtJaMclF8rI4on+kLNOvkhrhSbeGsNZd4AoWLgV1p88txK5WdkCP
+7TkiRpPRlNc3Pdj5wV8GebB8PNt7i+HvtQAZbO3qow=
`protect END_PROTECTED
