`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eXUV+AjECyVYTS6lO0FnTF+AEnyaewrHGhlW2oZ3/YrvWC9+AEBDGDKv6zobEobt
1Jh90s2gpCXuxFM6DCXssgDAjek7OVGI8JwpkhCB7r3CGTVwVoJYFunulcEIx31r
tH/jKL33ceMHNQhAWDeDFS8Hjnc35G31+SERA2A/sw+dH98d7miR8y6bF9Z1mmC3
+1UViHX98piVh5IllCt6LPuEfC02Ca4DTXzTPCKLEXkr7LFLCOh8yuMxLVb+xF9A
0nkEDQzUBBqwqmPT5A+vHorhgXfZIZftnjUqu9GEqfP+cmH4LO1Bw3QMi90vVTog
daVHU7FPaxhFRownGyxDkbp9t3SnDgeOFwFl90Xfpdk=
`protect END_PROTECTED
