`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KuE+y12Gq2B8dlhxYJSFSUq57a0vJE24YOMQFZXOOBTmPc5OJzyy77uwf1DHZkSg
0CWb9irwk6E7TkRyNmTVzxAEAEYHX/sz75ZFe4YIr3V5RCQNjK+xuh5IIqz5ODGv
IhbIbjAIUtbpaTwJEV26boyncWTjB50A9TnhKbkPw9Z2lvjnbmYzQ9HS46QvzPI1
Kzqo8AKvjumZCsB+ryB2ChHpcJR594PImJLqn6wMTiUyFVI1SJjP+iG+MNZ8Q+TA
wZBAA2vIAJIV8RkcIGKi3qaYefAFMXIhN0Os4HgerGNRNt0v0h2nS6O+NawRzXpN
M5qPGcW3a0g9ZrG5Xwn4Abx03I2Y0oslrDZ2IOBaLEJ/51UwU2LNqMTx2GQb3YIg
2Jiu4GAIWvlcYrN9nDea6SKEgxHNhZgrjEk+vxkFQMIWbNV2xl/TvI8c9YFuOaqR
AMsdrew8E7k8cpOtm0v9RHIO8hg+9oKGYn1JxdRErLyREqgIZWOfwcVL/J6CV4iZ
n3jqOpVJI1rUex3TrXgiIUoDgA2AqkznZjsSi3v0vFrrzQw0fXciRg1DXGp03Dod
HSixNN4CNldkZyLsrzjwuMgv5FVlr7YCQrLzVQTmre1c0hJgxY7A287jjisQj5tx
McmYtcb0G66/FsFzG5q8EvRi/yxK/7lDlHeP5basTYyN5WZX1muv27tsTmZTNCdr
6BJ+9fv7UlMPrFqN+3BlTjI7Jb5760ag+qigFsraooUPwyKzwHSD2bqzcbj16n91
8TQNdl/KkL3FAEMVlwFYwPkOy7Xjeoh7ty4omaI1UUQvbBJGW0B3y+ItVGfDn4V/
ONKI/ThjApEfmoOavkbWzfQiqcmeJZwCfGlSsHhRCWPRDtNyeqzqXcqNzj0R0h9I
m0kRcHYwpFvTSgFrhEGScmgtHHOTVGUM9jGo/Mg5cWRMnI53I45JeuPL/YZU+Afb
wDj98tRTgQ35UTlkZwNQK27KjQmHylAGYHhDZyrDNxsGFoAkpVdt5VbCr6DHsvx9
1tycfa7vkklqmPDcGnS+Q24VDfLBPcj5WG6jMgZ7kpnhaVDQKKH54rdBZiJfP8A0
7VpwzQsjXcFP5BxB41a97b6J07uX+LqgMkBqQFeu/0u+XBm8gdpvxx4qL4vqJDdm
wwWVb3LdxyKlirvZ1eikyhobAR88hsgX8nDuVBNtpdGMRLKQbNuDp2xZZKHPqWiH
rCgqqx/VZmjhhJ/1FeZn7UG8CT4CUj7MZ4WpXdDh/eLNlla+sKGL0Vp47f6gsrWq
dNTcRrJLxvhPzpIoP4/mtcByUYZ+H4bfFDX6HdmNVKfC6zRhS5s6wRUDwMsNRPUm
WVOPl8k6oh+djbXX1K+W0f1YJNq82Dr7FIxFw56yIw8ZmOtAhAUWpFQiWdSPQmnA
TwVy1+A9elt35XIdClm0w2yviWFUX4ogV4liqhIcfxQrIvgymIk61rOvbWEdeXOW
vKOFGsJl2bjzn22dsMDAJBIq8jPv37KnZsSj7gpZ+d2FFEhL2QUmX5ylZhU/RfCp
zMdP6eBKZnQlzyB6sAYcMi/KXoJHyM9l+V28Fl1jFzFbKi2RMx+JhRISQmsfz3QN
t53l6u8vmuqfgeQ3NINtguBMPEi2qvbRTIooAXpQUzmeGBU50n86Pyc1cStXH9p3
i/8M53SJKd3EMSUhnyUOAiDQV+GVRG/j5ZifyDSlmlISb3YgJh2/KHsCQkYeUH7B
1U/6f3EK3jMU+3wH6hMSBmMEg4etkAyX474/1OV9NVqG9uSy5NDxi3Ymx+CJpPSX
yrMzIWao8duevmz32q7PABq6HiIl3czNADEPFnM8muGOU2IIujnE2750sHpXHkh3
DHvP/pQdiy3U9C+bXebttHl1olTQBuDHjWIUsnziyAjJpfqVOa24PZVHOMIququd
mysaa/dplXj4m0AZ/IUEmRQlvT5vYtyoxB9TCyNwfkuvOuTf9clreqfz6x5X0X98
6I0fZjS0F6yemlgJITGHpISRfAooNRBmxOH8Ji/LH7wm0FSuSkpULCF89aD3sWQb
5ORQ4d2Agcs6jiarhZWK22qtPOcf1BORry1hw0zvtaoXTzh/gPqXXq6TTbH7uzmB
7Hno+3ZCIHLMzZ9DpjQZtfDL7WtaU5c6+UG3bh0f+ZU1FFHbBRwdBTmrogGqgwfF
uY5KaqL/TzPEfCrtdu2HF4jYeDMy7eMV8FWQ6Kd/LKF6kVHoorHeQ3kZgEgjHB+/
F6OtH5MhY9QiSyDr4pVFQ8TU0LmcvjcWjNPgqsqODxRaxW1JgNsCavfAdch005U6
ifP8HQAxLaoUa3XtkKQGewZHcvramhKpAJ27SHYoSkkg5aXAXCtOGpe+nLEVWvd3
NkXNuPaa4TGMS/R4s8Cb3AkZkaGdLnCJwJF+oPb9hZIGNNYz7Ly7+WKIf8IYrFUg
ehRR1Rsm6yNV2HWDBU5eTtUk3MZEB8ZpfJ8b5YOJSt459BhIWSNjCNWL3Y0o6GQJ
s7EaZ7vpLKUGdAwjLwylYZiUhR9jtvCNbprQrEhDlQ4lSAqX7Y88khlDi/ZLmqVt
IkunWxDod2SWK7QoOvgc2mYYgABosud+O4zQnRKjCCGUGUO/uYB3nWoiZvQxuoPE
ftTB6jOEctDDVN4Gk+wiJJu4vscyXw4BUKUJeB7u+tuKk6NTUOZsRdSdTfx+ysDV
Vz/meXHjrZwjdAaVwVA/5uzAxbGp8bs3UZXyDhk+LEUwfEDyokEEkzIVOWWFYDW6
lCUIFrMAbkpIohQn1+gipA==
`protect END_PROTECTED
