`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jXAq927dnAqmfK0UJOXgiHsYZ8MhyG0BsJ52lG+9upWD9R/rF0CgOvl7trXtqm+g
UqB6RwN2koI3Tan+b4o5ll0guP2Wtg2tClZckvHlC18m6PtLfWQZoooE96/3gfeJ
zvdFemysRIyhTpF0nDpHCn1KYXYWf7bEIaPKDzmXDMSd4f4rOiSMA78PujOyv3Bk
2TVcYxLErYOVsCtFaG1v25ldvZYzd7RS8bgXead+b58mzmPdyMoUTu2ZA3k8bNkH
A/2gx4GTCMDsatLgxGhRmXSsh0ii1jzgAdSaCSikQY4gY6Zx7xntyYYDKTi2ZBsh
JCiXN9jDw6L1HdbRuAFKWzUEzWg7n3KvuFoVsVDhvWnncToOBGyOjNALA0atspKW
P2H5/UN2epgopSsOhVpmAowUsuQ+LknFFHoXkxQO8IUEgS3LluT6QX4J14Mq5WKv
n6W733C+lkIfmNC2/gw0ANBvYCjTPkY7+xIOhBRD4U7XPOW3vpqBM7pnoegZxRA0
DNV94Y2HOg8H2O3Fe+wbSdt0nAWF9TIGz1a0UUJlDubzHThg5x0QEXkJOKUmyxzB
GCEBfPsDWe1+mfD04k5tZLEaeBPiBOzuIZwxUzukVTOgMxFSLbntxTbF8UjSoUyR
cwvUNBEz2yd1pR6+1RqYFbhYFiRxZkZPXKV3GxgtCcAYobwex7+TeVC7T6gsTpd+
PnedTI7aPgWjALrxmtNqLivOL8u0KPqHizYISrpaiEBHkeWsuoJKvgxUP8l/5mWH
OouaGxo9LzMP3/d/P2u2JXNTfSLzuPcaB+pUqLSa7+j3uAKu7CGN0ubqoVdwc7xd
IhWtx30PJnL+g58PW8T3jY3sNrkkdU7M+xghtBybR/Njpfl5ZSm/DY/0Y5cTNlDx
8U3NtkG/jtaMPSOQw2CR35fRATATiw7M66UmtKCOvfZlDFpP3Ix+04eHDLO3CNe6
Wl9m9GcXfcofCZDr3Vd5VBTw3mmt7bkhctyHRRZaanHFA/5BpuJGOcGaMvYil1XJ
A/yX2wpQ7iNqHSuQuTV1heS7+cAwph0XNPegliGUNESWq3eGl+nCj9fOvwG9fh7p
PBKFft+Dtb8gSVvdYfI9eBYchfOcWDidTACdvmxx9YnkyciNKpD3pc1L+Y2rOt5n
W4Gwt4Ys68M11/F+5+X8Ua4fwPJ1SxLoiTYi3NgLNWf3rYRy6VW5Yl2G7tL7/XkH
X8N9eYFbUiDSyUi8wiVmfty4rZtQRT/dBNQ03TvZ7mWuHDd6V79VSCV69gFHIdjr
x46nrsu4lL2Uq13ZrLHsw2srbY+mJu0CvashLl/9mRDZ8kSMd3SOX21iinprD4PM
/Kk0Yr/F2u2hDlSo9WSb0s2H8EwS3DLMWgikA36tqSvHnnHkr4T6KUX17TFTbYPu
5nuSUDxI4VLj2GxuKmFetmN99yyfO/ez+LujKkq5d/F2qlmEmiiN0pm4KJmhJHhB
91FGo+zCvWuAld5+QwRCCBnj3VSlX4YOCzUAlPkF3ppoq8AExqWf9Vsifgqdu+ZC
szgRtP56Pr0w0eUwRHxqNAKbrPeyXPftVzJbp8nluLPIXV3zftFgk2+YS/0Zqw/7
ylFqmSEPvjlEbNC3aa67nLh0RBNMuTPxXQfIJnl4nCoTUTdt1l/MKuxky48w2wi+
/VsXl/ks2MGamDtdrVzUwWveuC/sHlG4Fn6QYzy/1jUsrL3Thf54RBpWaHGWWfzs
0CuX5jCGCLdwhj2uv7L/OcQz/qbl6njO3LHvTsksbsn7yVmO+u+NLIKEKPEy1bGl
YYT810DerKqaSoFgCwxaSep0ivO8h+DBdASt8YLndC500T5hbwo32M3ss6QEwBY/
dqRvbm53hN6FBZISQScYeVQVDzWF3SaaeZGh7vuNprE6P4pExHo56CysvmeNKGvn
EkR4c4olrz3md344MBIqBiaqY54l/KNMUvmWB6Euo/M0aRBNOWWMniZSz4zF5q7q
smL1uMKg/DklLc2ja4nnXdiBRYx4q/x3txYzfJrvb/ZY/TdeDvyl1ycBQLMWofXQ
PNAXEBFtFz28j4wNQuD74vxeY63z6n8o0rglVGeWOT0=
`protect END_PROTECTED
