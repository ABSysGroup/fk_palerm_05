`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5H/GLhaTlksgrBtPPd6jqR6M7K1tragmh47vbs1GLymHSyU1WlFzF+lu5IB5unj9
igvFil4djCXzS7I7Ppp93OZdgHZMq24w6aFPu7OBuwLJ40IieDSvuoh3dUXcutIx
1THgU7n/twxLuoD0gOqt4SzHkIpDiOOmqbd8t1/DhUiGEbawZBe8m2Am5grKddmi
LFYmeLLIg8hSRFmQrsLf1ivDtGcB2wzLGGfQbXMI6fjzSoun13mtqy2QUivf/oik
ynfGG+FWvAjYQI3/uVQ58aU4l0+9LCFxZpGBnLMjvZygm28fqdy++S5/pKIaeqqN
Hy5CfwCqlWBBjYI9gRN9h3w/Yvo+PvXJroCSJ1gvH9P5JovufHfZkzwrLxGHMD2D
2YARBZsXX2otTbj1/+XAxMf6bKGvy/zz7W89HafAGH9x7hpv1ea7uYBI9CXuZcho
qpfu49I5v377BhsGgnx3nEwGZT9KO4oDKtlj3mnf3Pq8iQpc9yzrSlpChVRaHVPw
mlKzcfLpexqq+gD32xGLyea+hBQmSqqox392jX8Vnspf8GjQSQk2my+CYqak6aTi
wjuG+x21qktA8LVD5zZBtSGLFTJFg0rJRf2xWLgJOWRUnj2u+WJu9swFbguC2pC3
disqvb5apLfqYL7xPiTU6SULNa5HXkQk/6DaKuE8r3o2Wk2jECvbCfjprfkTgS7D
ZOmTWj9V89UqxbpThylOfcttADvgvE+JbUs9SpBDnDd1B7Zon9XcKZLOvgQEl1qP
7xqgs6zn6jOHDIOtTjN1i1KYaZ7SyqM4MMhFPqCrKa571i7l4uLvVZYMwBLOn95c
vx9ZI51IKBbj1duDA2z4LOELG0F3OuJ9qhNPAuDCkRqjjB8t3NbbeixWiu60dLPm
QxumZ0D7a4+TbLZyW8P4zhgLXC17JgBhX5XgqgyirmMBlwVTJ3Rvas75c0ezvOGy
uY9JW3mejt20Tb3T8okIm0w2PmTj0dEbHDHaZAQ2inIrjqda1RAlqPcQcEQK7FkD
tsS2BrdWGaT9oxQIr0Cw0eRmFbvRWp10lNL04dpdxGugDvBCD1wcqL1CcWEEm+kX
YL0srbqW7s3sjGrzo+RdcQ==
`protect END_PROTECTED
