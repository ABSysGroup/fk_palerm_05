`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q3uJodjsyXk8tX6Pgj0EG/EaYVe1qJgNvgLM5jzz/XSU1o9Be9ErrmZxfjV3Nfva
Rhvsvm9k/WEcYmWU9odcpsPoJQ/OPVEAj4bkZ0fng3ox0LqLbE85ADNqaGvGcpaG
Q1Ya+VF+z+otlSp0b0NihaM4Ma/inqZx5dKRSJNBbigo6I/h3AtV4Ipqt6nm70PT
ZHb/lH+Wx3YaLqc1Mt1ri3ksowb3V129en73zSpP+u7g2uEwc3ztzqadZoLrY9W9
b7JEUwvE/BpuVzLE/7kQLRtyhcVtvNe0GtPlOIXGhBhWshGvZ7HiY+duT4SRUoGY
mUvo2wqqHXOIIkQogonPB19EtJiw4pogSek9HIu8M8n2KGs7JUV/SePKDJbokUUF
RlmXOx2W38RfVdxgPr5Ui4QXksY58Aiy6dcnyN0vvP3hwk4LOdBctmGYjZEX6ohK
j1kK1SFBZB4rE+/wdQqJLWIphExeDM/Hiv0wb/t2DbXc4yaKUTmn+tLrmKSlZgLJ
UP/skEraFst2iR40K5Ubjge0HMhfS35uXf9e9snxRHsjupLreGml0K8Jp0nIqayp
uxlozk9Itks35o9F2QfENytGm+RApM4Ya21DHV6mIUgrl4YLBcy9mtiUzCBEcj4X
vS7x8KeHRVep6QYrymLSiddkk9cZhD6j9VMsvH31Bv3QT0c3F8gxgJCFOjK8XNP/
iyZv4lJPF1eY2OcTe60V8fX543lPeG+SxhCk+SNV5RmSpSms1yOG+qJ+ntneaHRB
V1Syz6YsiA4KyPrhLxCpsmqrOY2szfF32byORJ/tl8G1keKRY+6xCEzi8l30iOeW
1WmVrPor13q/nvYmiwuXO6ZsvbzBZ7RP/NrrKaZc9B7uVNSzUOZz7y1tANCX6wMg
t5zPP9YFEuzp+RYT3Kj3daKoKk3r52fa8o2aQr8gRyiP3DiBYILaPkNJqgfM41hx
`protect END_PROTECTED
