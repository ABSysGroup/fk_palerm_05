`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oPy3EiXPfNAS/a65dOc740cf36x042i7fDhOg+l7MPQQ1V7XTBeeYh3uPOuCSHX0
kCsKndj5UoNEfnK7bPAhtlJRLWlOd8ySZHcROyEOrBrfgIHuvc8jZuRQ16LRXBIk
OWjgMFPLMKO4ow/I59y/82DT5STdIyikz61BY/AetiqXXurYm+k81BVRuxPo6IyI
JU5hyvfMoe+S4Hkh5C/Id5sii2t0HfG7nGmn8YaqItTM2TKeOid9/vUvmZtfEGNv
76VZEhzcQu6/3e//qrHciPetwhIGdWtrQVdoshFWz7LjZfcvgCLGCr7Dv30c5xK3
piCOwAqrxZbEV/lZS17TbPWwMUd9IzryKeeuSO2ml/c4GVui5w2f2mfc1UA1zz4b
mOq55ZhBkshus26p0Z/pfOqF7/0E25YpnPZ1MuqXynNNVPxxURvpYGCMOQdWOrac
3RL260iX8b9kAUIpniiQq758JVG5BeH1D1OzfuUf1Abmsq4UA9/Rxj9jMxW8Le4E
2YrDsg3hQ8wcE90CKGLHM5ORafdn+xMc7oholT8fmg71dO0+CHOe4630LJG0prxy
64GJWIV0qK9YRdholufpdLulnAYPzN8StbaiSGw0POEB4m9kYmMb+dWuy2Elpa5E
FFYHA5BiVCugEouR7MzEt7U3v6W5LmdBj0X9V9EGrg3trjO6adt5ZaFYBkXKV8mH
7laDJdrouQJjn75vVAGCNe2mP6vylWjYmXFuwme3q1J+UCtbD7jS8H1sEjJU4gag
t59pRTxS4MZdvOIaK1/QyIoNYIKn34z019tiNOIEMFTw5LmDUa/hwA2sM6vmzSjl
`protect END_PROTECTED
