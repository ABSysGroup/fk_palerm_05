`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J0qhJJxk7JKkX5fU6zMQo6Cvqs3rLvpR4C3Z7I1FErVpywPVcU5tyoEKZQ3PNwCY
fawaeeHc9PmIBqimJznu7RZmYO/sv0CyLBbaMMAg8Gc9yrZ8EtxMomdztrwxP/5X
8EAv60vB14m0S08+mY5tl7rWDCbQHgntLQ7kNGVrvvm6v2M0LDuca7pCKV++h09w
/MLy39/Mp8q10BxTl1WBMrNlTsDUW9BZdfUoF9vTk1ufxIKiO9tNeHc8ghXq64BT
yTPUMK6FyhVSbIehhkU7WPzQ4VZZg3iGsPj1b2nvUT/XDTpkNwve0OyXsGWiFcW6
VOyal7OqDqxNJFKiqR3Jw1/hKBMRrfcDK2ymu1yQki/BPnO2WbZ2Mzl5dS/iXW/l
mYPasfRd4D6exSxK1V1tlU3WETR542eTLKCSYV2/DgDaAVf28UQOJxIU1RgN12gp
1WfJj9KxSXD658VH4w0t3aPJcLTXfurNmzGwriDADyBcMqeTDqLY0HYgfEJqKyhW
YyeC+LZStyjcziErhGPcrceI504E8D50LPQeuM/CcyM8a47Mo+Rk5W23Z5crVkdJ
SgVTNHMIOzDa7VYG32nDUsMlkQE3XjLZA5FaBJ7lFjEiNOySMh/5Z2HoJEQhaCua
uteBbLgunTEjH7CfA4et4HLbwirIdHF5+wdbZLqBMGI=
`protect END_PROTECTED
