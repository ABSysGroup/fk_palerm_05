`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
efmdjDHNigiWuW6acwRSBXOa9mlSH4rg6Dd2iB8FkufMjBTLTw6dr0aob7F4XqKi
35rvmk41pNYXwo6hn5CJJco5Eapdtpay0nIKuaGuB8UQPi2ASlGhYCbarApimPNF
HAV9MUPiVQTcAxGoiv7LRvy3gtvag32dLJsUUIt6HQz+qh67DdU1jgDTUr/N7yve
v54wBXtxJmCXmsU2AwQbMSYzg5Kit0tMOA0Dy9htb1rlruF4evkh95rChzn6D8kY
XtHJv80G9tjTc/7SZcFBOvXk1hK/KSZSanL9qgPhNIAK4uCRP4vpNkEeG/qJUCDz
uWM5xCIvW6IqOu7dXy6vwHMNbmLTqVpe6aDRmN19L2cXQrzgOzq1qPz7+jLrTadk
o6+cXLtfIzUeZl60WeERg/FxtBaN2JS83Myt61Brr/HpbhfPK9BJVz215vGqmKCS
Wa4XgY1D7r2tH2+7MR0dbVscaptHd9HWzHxrSfFRmqbBY3Zf/9pHDqrUrn6aHjgY
5dRt9NQ8A4cS6tcZWkFzCMJdSQsEdk6qUtXA11MBeV8r+g8dgsC1hoFgTyd0HWRY
qYkw1sePf3V//v2DyjtMqXcXxJeAiC668LmBmYVvsRv5H3vjj4W3286WAXlgAUt/
cysFFV2YeFus08TOweKnT4LfnTLek/BPqM5OHT6ePAG15KaYG7R1FM1qghGZZWpe
2frRPbmeLyId9kKxGezeQKCvzIo3OzOIf9eMRe26fWxAvQsPT8t1W4tPlJ1bT8ii
KHzGErwYHemVQ1rWTg2xJjGE3DVH5qzHZyqgu3AYebp5tXeGf7krd7aY1xSQl7tf
ULR0PnQKqvpuQXv9geiXwHCOGBTSmQLvCGVK2Vb1C86mQXlYyPhiX/FY8I8h3zhQ
xeRuHiA4M5PSlfVeMcFbtXetobaViUOUWgusdtZ5CWJENXKLatO51MBST9dZ1T7w
y1zCmW2UxHG1hI4wjBUhMRP1D1KRbmowlf0FmiOqrsntcs0Tq6DY5zLN55XvfHf1
mqUlrflaLdtpUnN8TYOXuiWjtYoAhuHm/CmOOOxYYDkcjEei5eak/mTUjp9VXWTc
5s4UAEBR81/gEA5kMwaXHxvwahdNXRTuS/pTH8IUMkye3FkGJ+yYVf30rPe25XCX
CurGvHz0ChX/OO+gVSQSbQebeCQ2K2o4O5NjGD7s0VPNYxWcWU/K4ldy7eQL3+E0
0JFOsEU0qOQwXomSF9Bt64aUn28g0AvVkQr/zT4IoqW06vmzPCH8hweC5vrLJv1l
qRDwIRrlXrNxkRCQxMw4/XW3aWi4vz/MRviEKgF/6PBso9emdi0tFgHDP3Oe1ZZh
qdekNWb6sek40UAHVo0SIGWkT7qETZKtjKeOJDbqgkR2egs9L2NtYwgBWHCh+DVL
0+UDs/IT6b5xJD4s6IuD9RJQtbGq3cHnOEuvrqE/IhOxxzENWsQeDjnq3AHSB6s8
1uSqQCGXgKfUqhUkrTUi2/cwt4JTUBzNZ9ctmQkiXawqP77sWPLARRVXweCJvePK
0nKotmKzS6FBQZcR/fVj0XFMPzk6KGSeqNy51IFzpX8fWQCZatVPmb6xFGT4Hj65
Nv/8auHn1w3Qd9O3PCqUWzoObmx/HVCTKb/ZE9xwmWRiYW1XueLlStrhbLaVeSnO
bgRhVu1PSE6gpoUkdaP4DmqDHNkJeHEQR3LICvw+W/R5IDFX49EUes5TMemYd1fS
gq9W0t0/L9pCjYggJHxvnvtEZ2BF8E+ErACqhIBZXA1EP8yseR5nt2QxiWq83TjH
TUV3+jJmeBzKNLdTZzlutXDN858BJgb8oynlazz3Y65C2dagJCyt/OVxyiwA/GR4
SwelseL6b2hrWiGKa/OGEI5hjYtNzC938TD6H9jzliB9RdADqvI4IPPnXmdhY8gV
eRvMgBMPyp3obQ4i188+x6eRcVJA+RndSkD3eKEGbx6kNhfx3qShbxJDBCubiZJv
Dh9D6uzp7vDM+NK+4TgUymvg8UT92Ekeu7eVFIahxojebt98/QyWxFLD6J2KgLle
mipc+dgqVFYf6gVwweHY214iWU4hNeYFrn0z7LPOs0FFlyk7p0MUZd1LjOLI/J2k
zCapHqJN6/qEBmpoZ0eQ2gA1JNPmvWn6/jXzFpdC6+q4wCpMvqXT1sZPvR6RDDOW
4Rk8NGnJCFfY8JgSnffrZ6AKLoSTvzqJkWrFj6B9ew1+NSMPzl3rzdCJc3Ogf1ke
KqfGeFWDjUr97iG0nHBP75MlZ02VUxT78lYyvQCrFq+czgZWJ1dHbrbLFc7ZxlKN
7vRHjClQEyisYs9KCtOXR+E5XswRezN6EGzyQCGc/zVBRrt4EVEbxNRVNojh03dC
U1O0j5baEluSNgEYdNXjnDxdohsqnUKXkZQtWtRNbkQfm4Vg72M9qqDfs1Tt4Lqb
mav/4L7ELJescTVO1CNoIrhbYkw+rgBLkAuaTNAM6Mu0igU/WQe9oJpsgVrAPrNf
6v/gXP9O+J0V8mpsMVoydDi8R3IaoTaSopt2O/N2VKGM2AUJzVGrxh1WoC4DtsYo
6rOtCsUy5cts6CLKkgulPuXE9IF8jDJySkWtD/5w3odBUT9cLuUd0i/NJaBjEiQX
T8PQvXWjC8WLrULO+5nClkD4k1smJu6vgbwT/cryqlctGvX8V1cwcnk1oWTt9lAi
CrAfG00gm6EbzWUSITrmCOlEG4ndzBYBPoyhWg5Fd5yyW6wmaGr82KVB2AvcqNsu
Y+4JRJEQ7rR4fv6/2C8m3jVGJqu2d4z6ujqM98NBDujvo1eTSwrCiq4eXzXhDj7h
2KmFFxyir9A54jQxtwbCxhgUdBOsjNUk+0ul/hbuwNeW0p5xDKbqx4bobV0kiEST
uSc4H4hB8AvcHPYpFd+Ea6VtVWKBDBGBLiEJvGs9i0xtjeI66s3ySAw9CXGsD7t9
8p72R/qrC+dj4G78J2pN5uFWaXRItWJWolIeS80wkoFRAzWzdbFS3U9jsKGWWUyt
6LER0K9x5Zioo6jdT551Wl4i5cR8QtERZ46+OgDziMXui8w4CS7Z82xkytJhAzBe
dEBeupWiqrho2/u0Zg+xRXVmMd7tx0EyCQHpJjLvc3oerf9y2BQPYK5TuA+nw0bq
Gv7doA0VRZO2aCXwHx9s8ZFRBqzFF+j9mtVg6AM3EQfcmIBgJFpdp9biy1p0lKZG
8Sd/RUHMrLImb84BOzvdrGRQOqwBWrSlNcp5HeRoxPH/nsV65ZTgUg2Q9LXyrtkc
K/fBuL0cWv8IZJgJ76a+92+Q7n7L0UolNnibrQxQdxJ4JpT0KQ7bJDv/JJFAWU7O
iKMp/0RX5tgaT7pVpP34QxMsHLEiboTbBk6O5Kskvht3jrXd1L3W61WtKkVil8cC
Qr/qPAE0mM5PIkkcfefWF8kYcoFEVp3hElO+2C2x3aOxB4HyThGgtnzMiMy9FAqG
p6qKphr/Aav9nerBC6/GiNQopwqkDAVe3P9n0ey+TURXr5/WuTrFW1HPfpFeI7NB
64oXRrDOtL4T5VVAJchmCFE8conTMbFG8BErvKdgXiKFfU657vGmWXHTRQH7RsMS
qt7UsKjRte3QfNsUTHNfyOOukgH8hsDsx6L7ZdAyrsWXGegEoYDAh5nQ8S+U7ZIg
mMyfpSq+jnMRwIkvHA2ai8wnL+gcEiykybkAYTyQGqnl8fSJAzHAhkW72EoNPTIW
P3RPBSq9KQ6lPiU3ZEx7F2NMbGlsx8x+F1/2uVsFM2sSpdUHq44RgxqUuWGqbpXR
EA/TmyxjQeS8KhcMN1JI9qyXKRqDaRNPXCqkQ5K32LFqLGzrD2p7bOPYynUvq/mC
ywQ2huzzQJ9fkhw/P47ffILPp7+tR6W4NEAgrWtFdkeVi3VdSTdDpPx4LZq7UgpB
9TQraJ59v6h3mb9PkgdEYJiVjdDuTmrVAI8cfEMEsheexW7I9VoUZKWveIproiiU
REJBUn96R2xzUWyL6Z8fmJlZW/Fp3k1Z92+iXVqW2mfankUH2Lss4H+zkIBmQXKw
REtNeRwLIlnn5lBQs/Cyvqk2FaXOAJzxQ6v/j54JQC4AUESUPvm6zHs68ApxDLoh
pQFak4vlESy33kfKG4nJUQhmq9dWll1c8cWL8b4L1m6QQjK5TEASqRt8QNQIXVxF
6p4jnPd5VISKRwpgXFdnr8Qrwlw9k9258fzkLtIJ2pKVcgwyte+IIWkZJMjZ6wxN
jt1MXrE0CyRZ7Xga+MMaiY1RToIAap29Z+vFSZKfHPhCJ4wac1Hu2tT4KE7Js2PR
I7a1ro3OAeXKj7wOVlloZBivcU7vLgM4l76lIhtB9uHn8+O+VZTftwsEiW+CqS7Y
WOMgVfoB9soCZLbOY+L2eKTvSmPgHbxueUPHa51Jk/4wmK6JUu9lXOSDSJvUaBs/
vx0wu3X3nSE8h3tb4EOowB7ExRdOuYgX/B7RwbMQL+2mM7Df4TrZY1hFLhX3bEit
LkJSeJ4pMgCvwB6LkshiRxFzQazVqg/oisssMKw3LS8HQlGd/TeeMCEcmHPP+7aN
T4aBe3GS1xJpPdfljmi/9BEuwGUQXcfGHLwuBt8QfNXAj6r1ld+ZX+quMKmY67Cb
J+El8PhJljaxQZjT91LJ4MLBOnl2ii32tdDVqdjFRzoOESbkya+goHs7Um6c9obY
xWvLcq9EhQnmaQz6YYIvH0xoHGc3wBoioGmD01gp0vgfkD3s5zuv6xms3Pv1ck8S
M4UA+HW18MGfNpdeC5pA2N13GP3YJ7rW8huGZQIpg0KOulhWiXdhGu+PJ/NgDrAt
Mf/L+vioVJCLFPH+koQ1//hpju7fDzkJiKgFfFryflTkL63Lg1C07dVP3iWP3p45
HogBjM75jJflU18GyHG1eHCppVX0z1woDDAk2xD24Qa0oYB9AEX5V78b86kaTP7g
TSO8EQqAt4Co14PztG9fcXSDMGpV2UkVG+tnG3fpY74Yp600/FvZamIWB3u1ruYG
tFvVPgsGhtGfGmygNnXaTv4EKmdGtP1K41UpzYwWDY4XVuv/umUv1SV5NhyBVxfA
0JPHQ+5XGS0ST0rpXF0O85ws3abllIjuP58ePI6NS6VEMnJ8W+z3POdd3ozdxAco
X4BuTS2ZdToolpCERNab07CAS8PXeWz2qjMkqh/DopZG3oBZ/abHR86yvKKbDiu/
PrIMnE8lGgdBFtPM3BFpFUYXTihiVbaOtk4yAO6J8VHc4iW9d5xxDYYo7/BG9pZ7
2zhu//7W2R6JAVlKpp9duUyyIUsE47YlS5BCswyIgG632+FAjEG6Km4DZoC8UqOm
GbXza248mXcYBixebnbij0I7maixvYK0ylVCRG5oY7yzcuyIDMJMkDDpizdDopcS
ewHy9LzhjWQ08qLonQtik6TPBxYCHvg4VMhus57Qg2PDrR8PuQhaScruIsRkweYb
4mPmQaxUFuBwbOsqpDUUadcf/04MYebeeMvSHhrls4ezZGPoXq6zKDRBk4wymW2x
6IEIdpmdBZoFagxS5JKl5MTwDppxbqpP4SBpBOcDUZUEbuQR/cYoZjqTkoayVD09
3MJqW9+yFyU6FCEeoDxpHUQ4inK/m6u4GOpRWqgHq3/BbV3cnIVZGCYC3trvOCg9
ZqISZELUDIDoMnv/Gt6nTT64PdQiInE+UwFwdUrNhpIrWxvudcRKX7dx2O1ZQF1q
XqxaXB6eBCTPXzZQiclFBc4HiQQvhiOBmB8bMZuzhKDAtZPaSmIcq0H/TuBgEqX2
qT5PV/30a37BS3Y6VVAxe8NGJLajRFqd/B0sBwuTaySzYjIKGw+zZzNI6O9b0UK3
QOD4IVlVJGmj7o0YgI0c40I/IZzqOn9nEu5ncn3ytaJWq0ZAVgwWT8Ld06Wp5G3P
fKrP1fa6ZYM+22NIhAWSUzWvZhfQu7c4R/CM23xwa0XztodtorMkyHhSfb+pdYhf
6IKLVIF8kXJaqZx0qHCGdpjM/5jxFyzTxxAjRsELMyripOd1uAV9nI5jQrIOjfwt
T2bHzL0FkY5PxT+qUSjqBCPokDtZeZFOo1nf789Zxb3p/QPX8AxhFtouo6G+9r/v
AKktyBz4IXYsLfRY2Ts0qXFOUXx7Cj/wC7J8xPnoO3aMo63V3mFvw7dbka9WcWD/
Aa2cOMmoIT7JJMZJMsRxONodgpH5ZHpCo7X6+LK2alSDYn7SKtqedQRlVWE4KkdQ
`protect END_PROTECTED
