`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GEX0fgOsJ8cnWbe8x9p+Y/Ufwx2pEu4d7fQzRn5IvJZKnAV1C3efsH7wpcuyJaCU
+ZQ2alDDj5K6WZawf5xc8jXolzjIjCZ5ZJiDJyI6jPL4dlY7wdg0mXTYio8akxjA
KXzSVJMic7ZZC/8oAyx3Lku20NTZxxVK0pUI7JA8uk+NPNRllGXQCPO5W9aaec6o
vrfW6u6jnZ6uySi2o1LK32axGOSd5+DhQzALiVI2QuhOT+/KX41npvsepH1O8Ygf
V+MNDHCagLicRg2OcFNUb3UIGqblj4HbrxyO9S7NDYmAWfWEhnG/rYT/Z1cnvgPm
3WihXVF3g2CjwO8Zyd59LE3OtMb0H99tiDjX0TY6HaFhO+CWBLKhJNk4oNwfAKex
8MckWcybEHrdbGdYDBAVkJ9sHdXnB/WNIX09o+tLOhaW5s4mSSCIa+GhMZSBsnRO
AD9Yad1B3H7ZpEamVUMCBFiaFlHVawvjQJaUq4kp0vemY5KLnsf5z1V0DuwV30eT
OhyBlGhJs1WIvx4gODvaEOhuZKFmttV5OMJIMjDCcCyQ2EuuJOgvlmF5x3231lnx
DE+Q9rOtvX2fx4yuPQbOFpZepwMkycxoNE8SypUp15+5/QubdUlMLXU0CgNINs3a
TwFnQ1CAtjIMqEhrIx0Njw==
`protect END_PROTECTED
