`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LoVnX0pqMFxhUukPQss9+h2O7+YBdhPQBkk4MQL/Pt7FnnbSLji1Op3pyydai7RJ
dwKERAfn3SucNtoDaoLb38OVF5pw2Sm/g6Vr1ofTgQvfhLsRXxWTDpsZyenAh7py
VVq06Ku6A9X9MKtUw9agwgu2jyprNnWCriCNc5OzK71ktX1magiBwjWIosU1HlvP
r9KJD3c+l+hY4K2K4pZjihJnGFrRhqvLrsiuAWw3VOn9vg5b/2rVz9JcOwKrfKWL
uLOsA726nRKsV0mF8utKIwWVVc8NuhWGKvhHHyRDrZSiQmynJDVx1NmTp93GYMkC
S232DnMXiPFjrPk70F84Pw==
`protect END_PROTECTED
