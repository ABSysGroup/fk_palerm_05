`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1bUjEvKfeRKLysLXkmuurVK+GKRSIEgIiZFSShoXohMLdbXp7fgjoxOkmAGLZDDF
//JimW68Y3WbN6P5DJSUJ3tmlW4Fr5uyDCwFRvftaJkz3U8uUgxxynCOIZfKfQjd
GSq/0idpv5SpDRDdlAKmuBNjMkxf+Y+56qI7MNz9vGjOfOL30zIDiA2kxLWXCgbd
cq+2D4Wmf+fZg1DgcW1emBZNr7MoZ4oFt2qEcvSwI5L0vvmHNAYbqYkL4fQxIdh5
TZ3LHqg0cJjsxg3lnIYu8Qv7LK6xcYtCQMHLxzI0uTVWZbIG4EW80IrL77jG8b34
CJf0qMAd0GymMd3nxI3dixnnJZE2bKKn8IcAaTQ/mRcH2p9GkmhUFtqeCGmpdWIh
brR+kYFObSAAtuAgaH1mCfVfYWwB43Cwehf1fw9JWZlWUnMzwuV7jcOuiHa4w/k1
jLSv1bdZ+M+/h1WVYtXxiZx9yI+5u4YnjALO1BWUHdTvB+wLMOjjBoeAHN0cBvWT
`protect END_PROTECTED
