`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ONzZL3p5FuR/wP3RH531HVAqfcHsdiGqzam8DU9iR0p6y4nSJNfyFdknmvIn+NcI
2C5NISNxCSbUThMUcqfeRiEnpEtEzpB8usfxupGTWmgRxMpzgk4dqw18iQP4GZ27
WS2i5ILat0v0EXNI7/qSaos9OGUWElC61MvcFO9ErzEA24bcmavR6d3ZXutH5V3+
trbt3UP4fp4Py2tbrNsWZ4vo3AZ/yg0fpjZ99cNxd2Pzhb/TrHniNqUwZKiEF0eD
CRIpHpW9NNk6Z53jW1QdIRNPsjt+nQ/VZ5AmO5m94YfAmPDMjOBywuB6SI76AMHg
+rMaB/VWGZxI2K95XPrUbESF/jyhSmT3qNBsVB455WiZJpKquR8RovB6XvPiCfOh
ZsSiypqzltEA0zFzKJAQzdwN+S+MgZZoRL4RpXCyNRN3dbHGA3Grg4Re6ohKJPOm
3U7ET4eSphXuJftUvpt6yOfa982Ln0gCKDGY39slEyIKc7lo4SbrAdrVfcLBovrt
gOnS/I7lyCc18zmBPoI8+tbgdCezdhfqx74P2Ggb37URtKoy8gHt+fJJIWnooboK
o4vi3M9kHP3ygJmiLdBxET9XhV/z3sD03KduC9vQE+LjeoNNDBejBdx/a1GZQw5d
ImZVaCimaMK6UiVMaSAY76JHweqBVQdsInGZLo2KIwXPUsGBMka6RWEl0KForLy8
skxvnvXywMk+Vl2y18tZT1qIAofC5Sc9Gl/0AxG7sYlr/c8jXebnQu9Sqi1jAGIk
xQjsumZ7l9CcBJAa6EroIUUGjZMA4QK+EpFD1W+eMpbSjyFOLRQIIBpBTLoUaANv
l6lezmnqybKRwdb9ONzdeJmkk6qERm/yvKOSbCew95X40+sIBTgf0MDsFtb8UJ98
yj4g0XKZTr6sifoBoA+9mzHzGIPEjROQu1trz3q0l2g1fQqZSR24Pc1bhfPHPo4g
tkcauwGR1GUaFYYeWjiwpyaBo8Jzhz5B+L5wZYyMTjT9Shx6lMSwQvAx4rP+cfo6
3FT7ImeaIuK+iCNp7EPw5Ug1UG7jY41ZviZKKajKjGYJ2UGkIvH5B0rZP/jHHLZF
fqjS7FLQkgpB1ldRTX2Rfs4kdRawbTamISJHPmIrmW2u4aGYZ6woI/v/vT4gI89Q
WWHpPyfOjhgzT1Iasfc54p1gkJ+K329Z1L6mA3aXHUi/czGvo6Txp1Khh2DXh165
LayNr9CPIdUtIIYb8p2rJeUstpL0BTbnoMrRSUoHmTWgPuY4qi3+TIvyp8Y1SNbi
53URrNZHj/78ebGwEAUDYY8ek4c5WSkUokcJjbrI8Zq56YthdEV/nkkx18ai8C22
DaeXMnZ7JyAxycKU4jv91XD0+uL70KK8qah18TsDcesNt+dKPpvw/i1yJzOK2nJ/
NDz8expUJQGDwH0z8kh0/tYBzncGXeiVL3AdJ1kzPPBcIQBlBPMtwIsQMKmEqhX9
FKp/sSO4hh6lCJ5oJmKT3yf6vWzrjH/yG8Q/LTGcyATViVhPub8l6r0dFBk51JTz
qzc3FYIZd9cLmgaCM7TH1YgZwWPPY0YSN8P193ed6hHmIPJ5ptzkoloWjJ0SXj0l
n20mKysYGupOnW9fKCpo6zzcIzypCMDtpfUVZ+stTH8iYBmBx3Gb7rPF5/mbusiT
LAsahpInfBtAJ2gx9HlQnhaMh7rQqFPPDUyRhGKJBMH6j64RLdTYIONSFPoKITRU
J074UbalKVejDoQsmhMqxmpnQSMTu1RSyoXx4E16CmrLkv/Cyo4M5DMKEpn7c4di
LVtKCBQ5bPreSuyhfDi4XdEuAcror558rr/fYCFyTkWKteBsaTegTasU/d1sEXUn
v4F7K8IiBwZBFf625vxwEaF3uXwkmGbiE0Oq0l+0JWwigj+vRLwnbqimX7rDLZeg
45llFNFhd6ImwZYMSQqaIgYMDlpf7h0352DtZJQX0Rv2WBlTJmUFmGS/6Ngt8oRo
yLsaVNegeoYm4in4tptP59kRlaI1sYcgaXaJKeScHRymNqU4ubN77cb6bMQizgZT
gKRxLNSwQ4BIaVuxPCDSydA0Ra6Fya84HsemHWLopn4fjCk42JvvH2Kn8zViCnbq
tEA0EoDt43jh37MVo2AAlPus8pyJH+e9ZrL8hbMkM+TqE4sT1AvIJBmAVgX539Xp
LOc9YjKpJ56gvbszZuOaU1o66HAjVjGR0gIV1T00XvQ0tHJjtbIGPC4N1ML1+wtO
duLymAHF1ANXXaEk/AJ5REq9YrnHghTqTek7u1ljxkrHt3s4JjofJiy43P8CvxAB
KGp5ZcuW8qvFIINkvVCUE8jR7R2c9Pidvcth2S3tREGxh68dym2+5ba1ezQ4TctG
0KeopdKYb6TcG61Ef91WRNKq0badBh8dHCdnHoxMYHv0xkNNEF4p1VyxKaBbgDze
8pMdn7dyBxNMO+vBEBoAw/pENcog3XLTnuA3Idcfs/gjMcpKkDa49CqpmA3p/0Dw
0D+1BGH+Y3otORcUOV2ksI/tCnTfwaERz6eJD258qsK020jw7DY7BXfvIu8hVwzz
0e7v8l019r08P/0+0pRYClbzSY65kZnpIoP43LJ5Y/hc4dagKgcggpIFdzUe06Wd
izHLy0POIjcjusWPVT0lpxpQ3bYtxMajuFs421IptFFUoOEOyIGlgqyQnOkfDiNN
EhaRUGNQVgSZHv+jsCi2ra3CSRL+7t25syN22r7+BED3lSMf54WYpzEQITCv/XgW
qQfRd10qMfhZRyFoUsv0yksgKcVYCbu7wmsyahs61oAcbohGD86DAku3g9l5pqm0
7UGfug4XOLNY79RnD87YDFcygHHq+RGk8MPbwdX6LbyQliekjXKksBq70sOiP9z8
uSt/pKtN4xI7WpaRaxuzymym0V2nt1ShIRtUeJXHbW1rHW7X/oA+Rncwenc+wmP8
NTDqQnpGDd///eqO+JRyE/Xc7MwrD5ajvsOodx9DGgY+nCQ2705dbovgeZuSpia7
1oAII/XiNw1Z8LOSZ9XE7wdnEJ3pzAw18fXzVSdONRCegm3bLOPbgv43NNofqGjT
prnJ/0HNXCLx3LeIM9ejd9CyFD3GFX02VO7AWUz46iq8IYORYrR8ayX6Cwu+w5Y8
tJ29iEbS2WLHa5aZANbdDPS0KEtS++D2Lv6Fhi4C/yISYYU9f1+TY0ec8yDOr8I5
BLfJla8/EX7EMmjmaLLxk7PuBnhZHD+wwg6XA4hOR+u/jqdwlxn8AjQIRGgSX5cx
ywfMZvjNTDozsWig/qigO/Bcyj8FCaDKSI/Bo8YEuO3awV7nbIM8Fm6riRyBfZ/3
IlhlTWFcDUaCPB6I2cj6PcC5weUHHNxig6Gg+seKypM=
`protect END_PROTECTED
