`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VWX27Y++XbzY1P0B7+rBAF81Mi2SD/gfrVBSMXjAjL5ELqQwZxtSeO2TuhmMDqNv
ma6Mp590K1l5lM2PaxdusmPXnKLUepLvTaUqAJiizis4JiJZMqdAvMH3Uj6MCD3O
s0rkI2CiYvACXqATxFAPA/SVZIJx9Yvs4clIu8VN0/o1aZsw1VG7sjPTDW2a98EY
QVsAXW1KADwQCYwIh1HhDlWQyB6Eib6D1wRP7Vy+MBOues5B/gvVYNeKtQUQB96h
4Hs4xFxpkmGACR22A1U9CrY2RHvvWQJZvNFeEyxIf2k=
`protect END_PROTECTED
