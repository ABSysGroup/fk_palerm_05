`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ScEDx+dibgnWMFcIy2BpvgRllSXI/CRKj+q4T52sNUJ8fSjxMaBMOfwrtOD0LjJA
1vjgYjoyWBFkxZ0ZXipBxbx1lc6A1w9MYRaMcMKsrisShI1P7tjptfBCBjPtzgxQ
R5km05AnHJyVQhN5GxUbRt5KdJI/uTkQuRdllUNBvjbvehN+v5p+KR1o24flvOCw
6f5oEw1zjujuwTY1aX+YFdR8IAfcIePb6GTLixM/TkyXMgoXTKNsCdy+vtoTUUsX
6g1buCRrqlHp5hnUHR3KCCjIurzIt3ddESLqUW+wZ3VaIvTVOOb18qejtSjHhulk
49GVx6WCfk+m+u03zvktMWSOAdLetUzEhUN+i8HPQuctx5v8CUecjREM6hPcCqVP
faMA6aP15PasDJ3fyp96Jl9eYZ16E/98DwWPCJOnOXSrscZmskRx/LrH2fr/sz44
yCSAxhs9EksUK125v3GHDGo6pMTCjBJkvFtViKpLnNs=
`protect END_PROTECTED
