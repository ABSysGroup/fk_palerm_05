`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x7JJ/a20q5pFxQkX00g5JGMgjByv4IP/b+P8USSUq4LJ6V8YbTB2xf/U1Prbtrxu
omqIoC0vttySBtIRVLrb8Oe+4DnMwjKxj9gE37az5vTxUqhWz9cP7qUQ633rQ8bG
Djdx8t9pAJS4VMTxsQWzZ7Bt7qUlKsCSxGTU23MYUt3dm5BHWl1NC/z7mOh6uRVl
TJg4SqfQZAnJYV+wmg/i258KfutFQI8M+cchJXPanHnB0ZbUFArZ6lyvYIZ4vebh
VqNG3z56OkQzjbmzKSQ4WMTbri57+N6sY3THRbEic+MyOhMBckWcWe2E92X3BOOv
kXTezQamJUHEUO90gWlZZLPYaNgLbnjMyUmN83/IfxrX1gH+kjBbj11wd07jo1K4
gQ5/Q242QOsDn0i9r+vP6w==
`protect END_PROTECTED
