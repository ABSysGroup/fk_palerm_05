`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E5oYtI0vb7HZlD4z99GyHeisB0xeqfN3eBd7PLP5U0bm9m2iSr9uTE9MN4Xqg4yT
0PGKfx7m0t2Ns2keJILH6tPlPHI4TSE6YFPcXyVhkSt3X15yUoyJ0gq84UlXRjiS
7cQZuC9Kks2kETiHfP1MVI5o8rGnHT2/EKI6a78pZdfnF3NfEjSX1vt+VpxWmvSM
p48thHErj8SWSfQ9aZf7gIzr9MCg3IAADmq7LMqP3+HBihb/biwU+MpgaqMV0Nyq
LpaJCgiWWNGOPtXTI549dOar7d0Jp1kFyxRi8NKIA0WtsGPxkTxmW84F8LQRXtfJ
zaCL7mq4+ayrc1ivPV1ifDpZN6eGd1wnDnIsT7V8q/xdaQBzDVQTCJXuMdgilYm1
+KR0WrJaMGSYRh80QuxE4xCmYp3tGBi0jBRTMKN54paUDHX3VIf0cwwpBSrZorpO
`protect END_PROTECTED
