`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CMAE3TLHbf8EebBuBBM7nlCwrwQWfKb1SGcJR+UFKQ6svhpP55Q1e8m2UEa5MgSe
sPclACStsWGJ0/NRb51ilDjOyNrZs0dTHvxWMMisOffiXt1FBL7KGATUNvDq4A9J
2N0wLWPCx9J6Qs9JMdbK+AEsGnPDhDdt9mTyHSTMheHiq4+2wbJQ2S3i29wnsRJ3
aTsssz9Z+au/u4V5O1XytA==
`protect END_PROTECTED
