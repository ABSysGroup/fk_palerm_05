`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gUzyLa8IBmx8asc7VTzX/+sH2uAFrjHT6I3YRw+NDXgyVog7VZ2/teicIgR+d84s
/XN9XUPft89553x/lcE+l/0FpJekYQdTmVS0KEZ+JcMkgcCYlVVwjYEYpAXQgPVd
yx9W3RfUe6d2mM/d2bLtWIStjoniJ6o9KplX8EBZh0g3A1jSBZ+KvEXyeitKiSci
5K8MzmLCQc2zm6tRzyWDijgVbO6d7XjATE0bYH4g2uXWbW24/5iNNm3rewdIoDLn
hwHc+1OAT7cyo1bOR/yQYHWDmyDbpAd4NyVZCAu3OBREfZ89paBxcUrSGVjulbPJ
iTA0YjPAc82nwYXyljW+0axOgg2ejyl5O4j5P3oPr9igL/Y1VIyIZTVfLv2Ig2Zw
m1WmCwyXBWNMABK7XeXbQR1IdWpEDkvm4shY7jAxOgFeO0H5Mi38YKELykDYfCw9
3B5OVpUSV68s++qENoG5gw==
`protect END_PROTECTED
