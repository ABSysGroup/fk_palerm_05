`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l8woLV4apTX9nSRrVZcVd78lcViaRXVrmYJdbtF160mFIyWbkJm061VgWGfsGyWG
xZOZu4kUDWC+1ItCtU8Ayi25veJ3Lz41ldLkIGhWuPAQR9jUlRd9KKSx0StdbDUd
goEknILTCu43Bh5VP5L7llZ7lIf0GjbwqcXP8K1vFCAVM4bQO4C8l145jcbHw/LY
nEQTKDNHnUxm+/6tcn9zznQcd3ob+7zGRjkVacmiTaNPvVj7Tiev09cEjOSsSsgN
o8W++Qm3oS9p8/ceDIjpY8Yx6emj64+NsvV1KWw1/82URqVPJWHm5vYXubW1B2XH
PpJEUjDoJGsWWOBZrVgo8oLSwI6yZZkeTI4TQ1c5WYJt2sWbuvzfJewlGJjXbOk5
+uNPtCoAmrveXx4W7cGuYWVvSiiQd2p9bGgmlZsNGTb8/fEWu2hb3piv8nQwt3pd
JFzgwVzlqmWo69hWvMqn2ORVIbWNShJkx7DWQY/wVVDLAzwCVjo8ZTLkKfvR0J70
GPBbc8EWU4VmeoOOhURiFAbZlGYk/2rx2/4J92c45RA0qaxtHMKllfp+xEu6RQZr
ElLV/IoPX9U6aJ/5NeDx73mdSIxfrpsER1kcy9knkEAp+OgedwgbdFfFeQzvdUk0
qhjQI1aWLsYNMHmt5pA0dCLd1IkvIZM4R6AELTVBOZLXalb5g/K7kuVFCgZGa40e
3KfKtOp7vrJfP/r80jHeaP+ije7iIXJoNxnR7ZY3rOJgER0tCqIsEvvCZ95Ji7cN
o0Ou2wycDWXwmF59FCaDTQ==
`protect END_PROTECTED
