`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ddq1HsdwjSdEyymBqN6a5+F0lW/5fHkj/MtZ7RGRgemuZWrxnM20NRKRQblZheBP
cYeiX+9mPBZ0b5WYKpuOSpGG0GA9PJUt8t6KbliNg3YSarpgy266by7Su07VyCrk
a6RkuNBmm2Cv3dKqZ7iZrKjb0toqRbQjKwHe0JmefUe997OPQtt/QJGcTtJE0Rrs
XN2yvF5gplO8jjdRFmfvziB+23lwm8bB1v2GCUzk4ZZzwDKyVxrVJUWnanYI9jUD
3zo5DJQR+Pc37J6klvGc5sTPGwJQbnEHDGa+TsaGuO6Frx2gHsx5C+BuTy2z0P8o
7Vy8QYlb0ih7ErGD0MHSSSU9K+pyOsfW3qABu9b8lp+piJ7t8d1ollBfMT0ABUO4
a1/dg8mJY0Ge7FlQOUU08u4ecBr4UA7rALm1WnynBt2oB03Zlrxkb324JEbgozqq
WU7mw/Wvq5LCaXgr5cTT3shQrneJ4nIxTAsJ1dXX77oy/oLiq45SSkXdaJ28P5RB
n4VM11vIHilFoqW1qmLZpubUJ41clLjHLdqhX6bobqhtnSXo0RnVf4vwN0D8yAx3
XacIQA5b3Lry+8+b7ZP4tsBkEW0UBJ32bUxTyuoN4Sz0iHzC1T0v4501gMT4+AFB
AFCpzlYpeH0nU5LZI5hNaFYjF2Fe0zq2qlEo1Xf/g8j7WYetQJT/d6xqmX5RFaOj
GCNgZZcIjgZTM/oIxQue0GFBNPDzC8DSYP8bqbQq2ddJf6KhH0F/1Qn3ctavw0EQ
4jcW6Re3zffMNEGbX46Izww8BIxGY1YsO2mi4nYdkCwSmX41Crqq2R40DNqTy/0K
2XvEZzfTXXwHWY088fOa+S/HPcD6i98Nw9ZASHIibvidXX/XsKNtq6KpzxPnqKQy
dRXH6F2+Rwp7AdtwfZic9Q4j68BZlhLu24YMAF93q6oLz+GKxUj6PPJfSeuEGPpL
d79rIPcCzbz9S2hmBGpcc+KmeKmwLMgsV64N/3AYfBPl6HVbMLHgsJvKMTsGy/1F
Ad4kies+NDTb+z8AX/u6YwiZPyo+t44lBqMmVYPbnUyQtc2f7neRqmlDWMxkk3cP
RgXzES7IOOaC4SFZXa4gHbJgNusyHCob3TaF3JcWzeQ9yqB8RW1Ghz+6jFDlyV5M
WRl9kimQbAplpVad5c0cUzvdNSMEFhcdKX3J4qJ3cAI9cFuw9AMkUXA269boRPP3
wNlx74SdcwF+QNGRs3qSFE0WWb+hdvmNtyp4JOMckJ6XlHS5CmfxnIrAo6QvjP2L
ENSZW0a6E1G4b6i6ljzK9JPFwtrffhEs6ewWtqg3sjaBbwvLdGHjboprL/gmY2xK
Ncrk7mXQqrXHCllUShDJk7db9vFOx2pb/u2GE/AmfxowucbDydr4KdY6CazXksEI
4A1WDuRHJxGI7MznVJd9SYatep6x13RshY7qF0fYafhfstL/PdeEhxODuueXXiZ6
vt9gOw+3GzMheqS4/t5JirgsZOBfQq3nBBEfjqFqDIyn15m3akkcxCmSIzzRygL3
aFUM5vf6RiSnLY5wzO5Fng95eB7fKcrGc0tEj5cw/vmmC76ndAe89LxD9tisGKVR
ksS8ftaPfWM1RM0KeWkKeJ4plmfcXFqQ5wpwRTR++cgiTrujwZpgQmQDT5/2B/Mu
1Izbqb3tRIo5U9ydk48KM9RZ0q1PFp4Ihs2xuiGvw54vdZ6snE0yA3htKuAw2jtc
nle9mkL0Vz4X2wyvP37tGNN9BSD6Hq1fQArnXahFhic3TETbNL3QW4eXDnUzErys
bEuMikrGR1Rnos+5nI1dXWhJrGr7onOCeKk8sAtp3vbkVxR87Ttl1V+yg9InDCsX
fr70j1gV1Fk4sa928UGk9X/18KRutWg8xcqoewBVJ7A0k4hIRGsuiKEl585WABjM
VU1e5/Ix0CZEXnfwjaeHbFk6jBcTTs2nFf2pfC4uqAb8Ot4UcyTeEJfdmMKtedi/
muW+8LGn0jP6nqOxkj3rlQ204+IdtLp5iZTqDLVOnAP2dxeAGnapGmEK6E169s04
gjTsRp/ET7FEImI5ODgtazvDU5vhXvqAYB3t4natUmONAagA97Ioch3nWIhGG+X3
Hb7VUXMVYPsh2YT2QtwVKzGJwFwuUxP3raPa8/a4VjU+Vi33xJ6aBYI5zXqH3kuC
kq2i5FWueaNFmiuNwWRLknchjd0QE92/BYYmxa7z2AsL4r74gn5DxwTxN+S59+lu
UDsRWJAeHRv6DOQn/IdstqksXx972CEGvMGM2oOg73mu3BjS/jyKj95rs9zppIlz
7TpWajofd7lwHGHxgYy8FAo0LIyjEg+tyzWdmT707bzchEtvh+xZzGaHIQ/HLHr5
yxVusBy5PwVnl8JHuOjlWlITkOp6mL/pzQ44CX9NHxBYFfRVNORhHReG/u/6FR9b
`protect END_PROTECTED
