`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aCbzlc0YvOLvT5lLe2ChcBEzXDaB/FJeOIxv13RFBn1edeIiMTKPThSxnYhVM8TJ
U+i6UHrBG3c1U8FH7Hzj9Qu614MT3n8BFysL1F0uWCjXRjO8Qjkite5FlOqZnnwF
JB6tswa+7Tq8jiJxIK+RvRkFigFyLBw9h3PIN2/HGmRfVSH7CIz7l18Jr3TiHtmb
8hQNpQ042VGw3MZCWY+XF4RCBKXG5laeHkiOVK0zPzansxZ51iE1L9N7U3Bg9vtX
0/3T+HkWG/Lk1Wl6qJZeP7qCqbdoaj0Ia62SW1lSHk/8kmw/gw5m848KZyl02Smz
9BYcwLWqW+R8CLhSvfq5j+Xssk1fz3Ssk1K7g91GPMPtcyybs6QfGSSm521Y7a7L
4L9y/6M0knmJu9BI+jtcbyXD3U3J8KejqwStDxcRo6ReH8fESNKBN88pxiIpD0RW
h5zFR1JsxC574ta33OP++w==
`protect END_PROTECTED
