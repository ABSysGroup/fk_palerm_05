`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yfMbSqhLVr0V2aKOA/4UDfOo9hA77/m9H6DhDf64px/elhtOXtnPWShJFx6MaIBJ
FECCp8he15xtIrVKNKKxhJ7YEfCqv3AI+oiTn1rM50LegbCNEjZ4a044t0yLCoRv
xxr4sVRQZ0+vDBkFmYi6dB0fH5zEFufTCTYkpFHlpnkVEDF+kasj40fpAvI3mvhB
UvFgyBic2AC6jGoLvLWWfhCiz5q1npsYI3AYpH3bddlWC+XoWq+OxRW0rPuzmVKk
DeLlkK+6CEDYDetClS1kMg9YU4Y5R7HTgpft7A50lPtZ2mLhCz1hOxgzmP3+MHXh
Tb9Aqse604+ONNsTFxjQxYIXstdxpPwps99QXmIQIYe+fzxEq5vLLfg17pFe/gIg
eF48Z/7Pp+6sC+FcA1H13XCQz/u6NTSFhuGU7/AoV5RZyVEZVxkg4cXPfn4hKwWu
zWGtNLXHKuhloZ4ZGGa/aOwwomlf6vaW9EcU5THukHzRpqLm/7Hjs+s/cld+QBtW
iqCA/RekkTeLCHqx47OnXhFpSWuS0tJr5pzEwioLctx8+zlbxPGaRGpmKs3+fIlA
1NJYwGWleXfk9t5Qwk+QM81kJbIArHDIPmfcN6m6dWJrMrmiGOZStzn/srejRII3
7jDM3iTe8bQuyAJN4AfALoPeqexr9T4pSANKM1+oLgw=
`protect END_PROTECTED
