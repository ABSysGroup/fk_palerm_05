`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JFx/0gZVQpSHtiWn03OE66Jo31zqqt20+ocvfNf5OwFfTfHD/ALpuCpEfd8sB6TP
iKv0cUspqMPLBhAWSHkvHcjldf4bLIlW3j/b0GVwZYNN68RONHNpRPG+I5gqlJo9
KLhciFFSgq1fd8wvU6OlTTleRCiP59Qfj8o6zh89slcUHDkM610SbT5eRymNahDt
COjJBP3wPW9axwv7j+LIr/IgkTBmNLYtB2jDlJiZ2+yieVocvrwx7cz1xxoJ1F7T
8bRqUWx/mVu3DpsZToMoo0/cJhNHKjVGrxymYU8nSo0W9nFSWXurznOURAQWGnPG
9q0FvM4uJ0/oJ7AhOxew4g==
`protect END_PROTECTED
