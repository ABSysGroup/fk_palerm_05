`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Vi9OkFPSUAsxhvuGcN3Ur2VMFNGmxMk6IWEVgB94KIKZbjtW6AQYHnJTA4AyhSI
jXfLIKkX5gnLvNusSCcwquOyF+GSQpYQUkxCuim9qAJOko5N7aLg/rgT+fOthY0Z
jXIVEy101cTEhw12M80AzDjQgdTYOInjaj4qhJKKJhFeTgeUdQB79guampyOUZ8I
rDVrOdi8XJHAwoLtC2EA81prVI3XJ/fozaBygp/L74/V9W2k7Yvmt8uRnRpr2DxZ
QzkoZcq+C0ah6EL/ZY87/ey4QdzBAQm8S4ZGh3Y9SZtb8ssrsHqLZHillzw1xG+8
0Enwnv4dXgDDqJzRR60g89js47EWvtk+nKwp8rQ2VbyfRCkyByU/x3hjUoGwhEvu
RQcUSLTqhDpN4QYx05TY9V8NwMNmijLNJTbmQMrIv84sNJnRCC9IipVIwFFn8wSU
CodUUnbfk79D/jQiYWs2qn0o4yt5VMrSOBMUljWYRBBtBrhobcpZZCl2XRI6Uc7a
rNh9+gQzLYIKSV8ETX7pHHoVWQYW2ysgKvYPykNH7PlrNw/2NgsJzS9cGWQDJfbM
fyMkcoaQszxSOzF2eKf+QNPJpP5NPSBsz/6ChRRQnyDQ1+K3d4qCcr4n0QQ6ty1y
pMRogwS9NYSANRsONw2TQQHyMKAzoZk9L042QAOf41roiYdhYMNI5DNiHnYKsB54
GskZwa8Dn2SgcLPtR9H1+dCc6f9Z9n28cBmJVRVuvacQzxQceThbuz0H9LgYEbMQ
MI0Y8XdxMOiyHAxZAzDdLyK4l1AOgWvWyQrp/WzukMnfeht+7djOfeJgjnV3rx2H
FT02XM8i/YCajOgIvyWaoA5hjwpF3+hBitqWH9wgu5kvIVrPHC1tB+v2fnCUGBIk
Bzb+3Xt6k/wm7WEP+DN0N42YFDKFq5aJLeKZXibGcEFCflo4ilDOIcP0OQJODMPm
JNEWIZRHekAvFftWnG3TmGx//fcw6jQVxZJmDMhtigN5KXP+UdDc8Duh5qX9NUfB
DPhoW6/zue7nujY+0Wpt9xyeP6HJ3hJXMPg4r1f21kbse5bKmdigglIpoRQq5stH
viCM/b/65O5ikpuRX52/qayJ+ZziR88WWeNZVE+UPQSsf8ofaKoAX+sgIPWg8Ll1
9RoyVVrKRkHqizqJvAVE6IXSuTV9ePHhsdk8liXVTloMtMAKcNaFG8t8KiHKy61P
eXUSk4c+pbF+Ts0JrOMo+pbfc/Wx9WzWuB+1QvJK3K/JoWrVpylVd1iuwqaJlbgv
2Jk8XExXE0rJPZzNlS9/TLbuNcYyoHzUaWjhPzpagenR4pqfe8ij8M91EppRz5Hw
mkM15yexLUNJRvS/t7m9XRbwRxu6ybheE41UO2FUlqj1vi3S5SwS8/P8U8y/DPvh
e4f5uHS0ZFNLFcKah7FjyzilGWo9r5FEMZATIsYixh81yA/S/r4EkORwbEtYAlW+
/6rD/9Qfc6A8dHBM/wlrJLW8AccH7BZ9GGVI9hXrV7GbR3crahSCbH+rA8/7kNtC
53ewzXn3y9fTbxCzfuPbXD1VSkx3ls3g8WKIWc5avCibD68fURWLsNabBQx0mAgr
+xANQl0R2CuWPm6FC7Q+wiL+1XkhPiyq0cwTRFlU/54ToetwCSrlfo6gzOCSwZ2g
RkC2/PnWOe8WmSiKleHL4X2dGTI93RA2+m2p6g31v9uTCbSzRL/aPBhtASWedQKa
xJunvj2343dfZLsX6ibobej4peokiBgAZrMurGP27us3t+yAcms3RUyvPNbw48Mt
ec1tdyUdSZXqgdg41Y23EJRnwwtt0JUeuJgpGAJZPnS7CqulZUeV0e593zzSau/T
2s3K3OIhowfVpu3SDhao4LlYmQQq1oRhwefnVfpkkGonqxwHMbQ+efPZWK+MD/N7
gtiCp734/xRqSPwcmii2Svj5CkoVVyIA+JZ6dygklNuP7M6b4LMIeabqn/Fia+x7
udlMnnZyapEZV3+rzsRovg==
`protect END_PROTECTED
