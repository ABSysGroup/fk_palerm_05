`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ih3FoRWoWwLha7CJ1vBII7pQ46zzB8FGY8YrSCRIt4cf5eb9+J1/kHN6/bLnnc+i
8gZO2nwtQA1m768vQMnll7mUlHJp3QgiimRqO4BLlklrWPpsC5/JRukpS0Nkdk6t
IiICGFR3ats9H17/ArUsnzcnzjzAj/nhVQ2RnD6zjXeZz0j671H3399dCI45GHf9
KaN4CRXR5W7mG3HIbvd0CIv5x51MEIzHeL1DNRi3oFof1Z976XRERoPdkJzmpC53
FGg5P8n6PaR9bp/7LuZ2DCsewonCWajHCrEEvbc8Ge82LrR9btD/zMXjwBwSAJzm
UaD/CxhFgXCfkZlVM8SZavZBg/sK6bM0xKhO9OMbRjPInY/AskvuxXM73ElKMWAK
px409eUtxa4bB7cwThPfo4Sg0fteCtZBgVRUKHKgtukrQ4nwtSk4Vuq7ES/Venir
KJ89FCCU1RBIV4V5oomzHDflUwchcJ1g4gVS+oS8KcTgn4ovTR1hxPXA3o4/fyNC
ALMLm/d9b/C3d/Y3i/7wIVD2X+tbUDeA6Q5HMQFqYpYt7eLWrcc2utZnCyMR2PPc
/xK9JIT5B8A83YrfiupNMX9E1pz/q6vvt2t5PDMuUC3HRCDi12wjsnXZ2Pf9199S
57IOpZzcoJeYXT9yrx7FPz80y2/jPHZsP+g0yMYSdO+zsOff2XA4zbDVbDgm+tta
BXa3IMWLeoOyFt9uT/kNISK42e/mBy5kiRAz9BCpoXL/OvtX7j3fz4NHIAwGKcN5
cDgevvjYoq0Q1/tucVJkRjKbbJyu3FbhjC5V+5zFjjUs2Po1gs2g8ecYpY2BLdTi
Hyvt66oBihiE0RlxyjtN5dUxuGXzS3x2udD1A1cU0OCDQYMlD5uQdQeg5wzMFJtn
JynLsMtJy/KzO40TkwIlfF9gcc9OzopWKTjd8H2E0JHlosR8ck2Z/Ic7HuKl9nha
CiiCRJhwp0l+WyL5RJ/7S60RVkJo+W0SNQyytBxFYihVnTJfZvGrlJQYt34qdY0L
YCsJtCf+a7OkRjpLEN4/joNT7xDWmeu4cYvMFA6tWWft6pqKqxapnPItRWGnzZ5b
jSS8TfXbxizZlGgGe7gJ9uiSMzGcc4RtnllvhB4fLeo4OSnvgjFZ7vOg8QBigyM5
6isASs7lj+lv5dfjKlW2AVbv8EmwitWkdY2r4o77nqKQDiGaOgf4aKUhR9jlOsCy
073njNZQXkP0xEyI5X2ldMG8AqkWQrA4G4+0/oMtxTfFvGgQ1MasA28zueSuyumk
7yst5PFzYP9gOBEsh1coDAG7wEY1nIFoxRXp8WHqTxPqNEVVAbyi8QxGjKvpNsIE
ggPnqGOvDx/QDk96MfcDz+CbAQEQfxh9OXzKripHfwGUbLpwAH682kBfdaXsEXWm
+saJxXm6pkfGe+0xz5RHof2o4lNqK9ot9UigXEUV1QSk/b7fLuJYUTdktGTzIXeT
d1xZGJMGvG229dlIDknjAVk42+NBpdrbGL454TrCibJXrUgcfsO2EdKBjTWNdUKt
b8DIReILE1F5JVGg14H4M3HDhXuN0gKgUQxyD+UQjtmmn7vn7voHJkC9qzqNBQMo
fn6pWX1GLVYc8b/7RiHsTmStYsx5VvGp6qT9OAJbRyaR4syK5BSaSB6TPwYZziyi
fZ+6VN6033Yc8gWO4/aDWqhOa/hWd921CZ15eVtsbqTwCFpp7X4j0i7BEeAYnMHB
G9ylVsFLhiKe34mMOANfjmLZCuJJWJ0Egid7/PLhyb39rzVF/qVv9gSLt1LiiYeH
XZWYqUb697N4boRzfCHbflDwiVBUM73zsDbwhjxCzZ42guI1zFYU55cifh9sVbgp
lFP9ushtBtXaaYvJ1zCQz+B/S0jeLGApaTLOqhUX5AMp2j+hsSEBIN8bQ3/BPrYK
NT1oplig9EN3GPdH7o1RFiRVRbcDGE/tSmFjZP0Y8SS31d8QPXH/d5YUkXNoiUqj
Q/kgjQ8Tt1O4feA/CV0kxw5Bm9tzXipPfYWvzh+xQZjHcK/QK1e4PBFRhIw02gbt
828jae7LvuOakG/s1u0KnsutkItj79YoO+LwXZO//GPtdIts8XGQJ17xBzF4w1Yi
V7ykKWwK7bQ/4XdosJKLhyJnsAxnK6FflIlGV6SwAOzys/qbEHwdt9Vo5AGbrDhf
uRb53cUBVf1sdemnWi0mnM19JmcoTrc/Qrdg4dbou25w8jJYIn6/C6QNuz4alCjL
Y03qvqavrHy9Uouyf3aDBi7dInwfzFyXqwOEvuarnfikSITN5qchBF+QGRfJDmN2
xUgQIc/cHNSKnltcs0npB+knSPJJdsFp5+ADsLrcGv+8YfhEpQXBuxyKG1q04+Ps
lZDN8l2/2hj+2UQ6/KZ0w6+kIe0awRyVo1pFsmqhexd5mMwq7MfT2+fOlXssV0IX
ic1IpFvAIhctgm8DJxK1J2logD4aJDy7+U/MypTjsFMnVjJOmZGP3iVYKjX/c2+e
3hfoFSBz7JkiEPx7v1kl3dbH6ai9Q9zgB4PiX2RgY/kEICUOdSDv2ZA6MFJI+btv
rTP72U9Ogi20HAAL1zQVFZ/xlHrmSZOy8hBxgFW4Emvrou8XFslS+Hk1TfEz7hXN
/ezxsEIx6l+0/4f5S7mn7c5rTPpTNkEee6QCyVpVLccXv7uVmhXMNb1DxuS1degn
CkS4/DYmgK+VIpXpUbI0ivhq0DR61aW/WkKQAmIqx3A2iqZLAXbiMmqa+rpulU6N
sqO+9+G93isAHKV0ePUWo0LyS8kF8NPQ+1KFeesfVePI/AkmTh2I5We6hv1durK5
5471yQ6PGbXBfljOoSJwEIXjML2VBdeuZcyerx8XzZ3FLKpLaY1bGiiqLwjCzubU
fr40zAYVCI1FE/v8s2KZQq8mktpj22drFLpEjIqvGvJdiFwtFKKGlZDPQGFjfMbj
l9WpVQuuKxEmNZIkJtZ74/AZj5F9pj9Io7haeMJkyXnzWKdZpdhXZJyqF8vkkxqs
OTQJRY+puAxmOXzroNqMr8qT07cWKXQ3Waf+PH0WzXITcLnuIYSr/bWCtIoQbwY0
bt7FsYOrrmpI3IlXFJ+S9AjDEyfmsJyVieN5O0go8fqJ1sCfEUBAhdzu4SGssc04
KueBF1KA+FWvJPZfPXQbS1vBhwvLrj5SKS4aVW68llX4wf4pa2t7IMJ30If6YBCx
5vBKBtr32gog9Xtnc7si3kJhlSBM5BmJzttcxQ4gyGiLgeQagJGbP1FiVqR7O9G7
LqEyjO/qwqnKa32Nky7EAcJv6Td/RuKlJQTXTJzQ5MOsKuTfSPu3G3g7Xiigw4mL
zkOhyycQPCDDd7vx5CuEn4JjlVqa/edD3UNPDPZyu/KOQkRkx3FZ5vTeBSZRRFuL
lLzy6Vi4bIvExrO6pMXFD/QMRd5qrqNbz+K+mDGS0jcvZOYyjVM54/zUG6Z83Q5L
qkY/xiz5yxo2FOBs48N6uScKb7tR04g2DPvxZ2+Qz0A3xYlKTjARBkT2RK2Stmvu
ByOG/AV1QbC6sOiV3CKGP7qcN9FDkqNOLONBOOwPdBVSWJRKJdZVFFARZCIjUV4K
LdzEwPvtudM7pyJUvaQSgAA4xP1hrPkD/c/t6r1tLgCDhth42CCeDy5++PBIJ6xA
u8sc39N1B13ubI3qayod1Ewgz95iKsbMY98aA7mTc9n37O2qiXnxP+DTcdhpx2iS
PfeE9SEfiuFy4zJ22hetfUsyPNFZEZM8BNR4+lW86lRTXmKNxkQpaLFVAPmKqrKY
vywolESomqIu5Qdt+Ula+veDE8eq8eoWdx1Hr08E9XYf4sWi56rMlkWmJjIHNO4B
C13khMkH5Vkfva5KajTcyguP1uzvXcmCph00xtJheu6hvoD/KirULlZr5Ox22YTO
pEk+85mTWX4R/koUlNKBy5x2b1doBqtpk/N9K8AeQQa4khDzQa+dSqrhytIRPKFF
6MnxD9L/iQmN6T6S33qPcH37RQRSsdKxfp1MQ+5f91ZjkkJxGVN0GaGTaErxucYa
H5USQ/UuZGTKu/q06vwj8DHVh/XufY36trgrce5Ao7R2aV9lFAYGoPA1l6EF3okr
YpVhrHKQVJ4HFG/BRNbvjJEvWrhm1NibNhfqJRwbzsdfUHXK7IgdHBtZLLlZ6JLL
Sgt2rzwL91rBzqruaKmFjrGPGoZt1bbtoVG1XQS0lEhMc3LYXenb5kxwVh9bopaK
GwUb5O7nnIgu7/tXazBhAaCQNJV2YtiGJme0wOpkujRz0JdG3rCz0XVCu95MKlcy
Jv+6xbWK8li88pt/1QNhZfmd/oqzwxXkGiMUIuMdvUr1N6RTVXd8MtG8ArN0YoKF
WzU7GJKrGWzrV6mNKf6u33UeU7iD1ee4/gZJSfRRGSm6lG2Q2+xbpGbyTSIogZaN
xB79xsmwO4/elXFJcRqE7oUe55UHc7wXwxBHEqc8zW7GQZIS9joJyF07Duno3857
/dYko5O3LCLZ+LNAe5XeDN+ybU9g45+PQVewnfwuMZxFm45L9gOAkzkjbte7rQPH
gbobYibiNDiyCQNjhmu29xCYuxe8E9bl5IvhQONLFgBW8PvXQAPbxjFVg1BbJr6t
5wZpoCejQkzyHeI/0kt1/hjy0N7bYWruVTDxh3dXXtEZvokscuYaLCwUsZLlRNWZ
uUqppdWAFZk1pKHYt9gMcoLBmYaVnB95/Nf0jEjigobyXe9EUBk5rw5TD2b1Erbf
yYyxaqe1T92a4LUPaG1MJCg0Dy45EqjPZJqTgxeJYEnCvRIuqzFgouYJy/vqfM2r
cvKu1qSvukmIxN6xhP0vHrtjiPQHTaZhb290S8M5xUfy6LZ4ud6oiCLfE1dx9Qjv
P3ooGdYKX4KlhnicXIc7VXQjWiu0CmuV4PaGMV639RTLb30hCJ2SCUVia08eIerk
aEGIcM+eplnlZRPn215HKPM51rgGprAa0TXoQkpsLCStra6TFdet7HgjyJYiFTGK
2X4kKmSekhRvHair08mUO3aUOpS3+OgtdJp58fKK4yi6fg30/1WOXCuu/DOPhaDA
Wn5RvLWYCewboz59aDayuB9uC+jvnLmNMLVey/vcSGSq+XjhSNhrWPsrx0xpskZV
s4fcs7JZEGs8wcL62zI9hnBYKC2TutDVqmm4zMxKrk+iGAHZqFU9+MFZ3TK2YdkS
Jcdg+6akyQxsIYeuzcJDLKFM9+iaaGoQdDKku+Kq+gIGKCyc7Jzz4OIBNdr/w/AO
kjxUL1FN8yybrTiNZeVllTibhYDFbU8NMlzgBFmr5UGrrwH/Fo1k3tF0ZP++ik65
yGGlmi4X++9G4JYOGftple6n5G2jjkoBdcfAxE+6BmRepN5FMCm1+ur5Yl8UGPm9
t0iptK/zOT2UjB6r8pO73MMNQiFrHyyWvxSh/cXZRiFRW1cKWYCPtJlSQluUIY3T
sK7/Wdem4/vSulm2DpjBSoGrWFQZO001OsCcOh2Q1foOmsMqouA4Hit9Ou3WBi71
2lsgmbwz5sv6C7HEdQMoLdnPtzeanDW3p2M+/peg5PnLB5RQKHqjvsjav4iiWrvg
CYHwbPlEi4Z9ip9HGv0BGngfuElFNQED7QzhrzbUQdSj7Oz14mLl00Ey0NcwZ74r
589MXbAgeAir4oHUcP6cJykY4wdMv7dXn+LBbSm82OhJFAUhzMvrLHipDxNUSvgw
ULVnpDaQVCQuPApQNpBsv1udNsMD136FS6E8q0/oFyXGrotnXsYRGu0iEMeVW+Mo
AJSmHhTdyVlyU7Mlzr7RWKsCKmaULI65lkbJ7IQ+cB3piqJ1ToqxbbibQmgp6T3s
PANZ2FhG2cEVxwgjH/d1gT+JW/rkNFGTM8LdR2DvZbi+45LVD91GDMJKo4qAtzDg
C3tk/vYoMFHEVnZGG6dScDMu0Vthv1Oe72ZehBqZv5nDgc/HsmW9iwJ9eSWe8qqa
3RDvdqIjgKV/D6eQaBsWSYO6tC8ZN/LkkEHxcPdirnjuBLQnS4iaaabtYifVwqLg
E53b/AP3nWoJ4DUq53mHsFjcxbootistWxbhJIMCUHAvrl/XxTh8NcKjN+hZyeO3
X7pLZ6w8xjU5TxJUoABlBcz9+un7Sbyq6h2jlEqjwvWLygZMGx5WBp96SoCpVjrr
Ga1tmR6+Adc/XrL/uhx9cMgudBNH8qi/gw44nEpxmyM9VRom3zR69dAXS9N1z7oD
H6pJM6CJeT3hTZS6BBWftgUYVb7jpoX8ft4S6UVtOLwMOPSwdkZcTwr9VxUbTMp9
Z4yUZ2UquWFPehhHGhl8m5GiWG7J4BJQIKMT0AYTGI0B9fgBbzOFvOl18XRSs6Tm
oy/byEM8yQ3lA9Lgf2G40QPvFk0Gqc2O3gCPEqyaMM9sG6pjxyr0QBnCIsXt3MkN
WjQAUOL3jxXKqIErLylqumM27a+YKjLYVt2F/WNGFamrFNF1C71+lG5sRTd1pluT
fKBMViHVjiXXi3pWLeX7S9e1hV06VX8puFy98fqgtjfA7OG2zxh7Sd3uDiIcqEUZ
tzmDrFt6scCHnMb2SO8HmMSxMB7qDVprcEMA286qtHy3jMAu7fhZo4x1hX1z26qO
yAb0kg6THXKyTC3+4eYwTviUtfQdNhIt1Q/kZAyzS6pXQQba7g0H8B56LjvtgDha
KJ43ryWtLBBOEgn+XW2Lcw7/o1NzNSA2iHqE7s2u5EZJComdEztNLUB0wQx377D2
oYh2+L7OnjznQ2X39Fh6+dLqit121LycnzXqVPDMkvUkUFe5JzGY3/yKAb5tmsLS
sW+Ts9ppTa6e0ds8dEKCErycDmW4DhKUagvc2J91p9XGD+qyIhC1vKYsYWQ7/lKS
ODbGUWYfUoOohnJQKd0lv/4DaOJ5P01SEonlRO5AQ1hYRuj/+Nga5iR8KUIK+F+r
PJkRwPA6M4B9e1GURAZsfAmXzDJgfyPnXtdT5qiKiYrhKPL5nSgnHzi6ID4NvFuk
+J1h6pW2EKxF76kSkSGSaAmy0cl+uura6bh7qIJJnNYm3GYMPobuXwj8otuHLn0Y
6zSRcG8v4rbucN/lR8KNmbijZk/7Mxwu1dtSB8n5Rf2J44xiNw/Ww5JrvI38TqH8
La1Zwdo3EvHU8NWbjhr+GVegxhEIxZdfQgA9jLplxM++mIdEI/UD+6LrFSTHbw9Y
mZ0/Z5nZm3aGsiixmwnFkd+YVkri2WjGYSY7alcxIiwCXDP7DB/rr2DkG7QYbTq2
WvJWffBms4SZsEBQ26IlGooyRNqej2YpbmOYURWOsRVBAzctkrNcI25rXtrTdHp/
Go7aSr9UOJdfH/Blm25RIVmFLS3AwpEnlb/wOb33zWliTCiRDso+u80odNU4N8py
YW5X3upfTKCakEBxzf1Gy1MyOd+772zdJo98JPVxQLn30f1BRdEu+bgjiFuecOX3
W8Jhz67TN7Ao8J9HyzdCsA/1XjeG+Nv9mVo1MvTHdHceAAWEckDx2L9AmvwM7qf2
WX1RfoxhT8Pd4DPP6/I3H9iBM51m/m0U0pBzNn9jOQ+GhM8gBbKM+SMRjH5M028Y
dI3ul/nUkvXY4vEGG0xE/kQJ12uiUB5Qsvr8PLormmsHKpQnVn2YEtqcTsajTDUk
nt2VwYs+nQGmNyUTYqBefaBeFJ3TQ546FAFz/fBeKeAfs4kxCkZTKs5kOdxnGTtD
Fb9bvF4XBxBNgY3lwR8uoPif9gCiIWHqtxzu+eXFBQDs8Z2ePkAckHIPr53Hkvmg
6Ie8nMWRwBZhtvUNirsZsrm5GlHut5I+JJEKJReBP2KFRfuFSlbWdHejhwNt/BhI
zyN6ydmk1T7S6NHO3vw8hAKojceik9Zj/sEZ6vajYAG2tb+dJ5KymwxhyIavx/bi
NBa+tuRdc+uN5zw/Eb/qkMc7VZd0A40XIy1EEIZDFrhnzFO0sFiZ1sMBttsf/Yht
6rvy2xq8vZwzoTnV9fl5ATcMbQARrnz6iRCV2QiYvBmTOL07FVHkeVWUQq+PlQYj
emhLn9/71S7vKiWN8VmPPKDcK40oOAJy8N0CpFUnZQScsb/cz/5Y+CzxOns+GXS9
4jwYZXDDqgP2j/zBvtibhUY41/2+NN/bkeS1J1Bfk8bZolE9CAOOpazltrRPAooc
fuU1jxnv4DMYVCAlVOY+RH8whGFHMxcI+i5tKmyRD4vIY1vcVX4HYX9IvpsqUaDD
28GwrDcM1WMitMzkFS3XVI++EGVH4AQjXl6Ziux+8RSwzrRRTEELAyDAcDG6gdNs
bNWNzqq1eKSiZVKtXJBhSXwYiJkAf7hjr9C8UC02xLLqygHoPdoMd9EhAuk3CL4H
2Bwn0CtdlNqXhKFccjqUgMtUaAd+hGPeOAJ+cFOubKgHBs/9h4WIvWqWjBe5PeMy
DgT8HlO1IRbGj1wZcoyBYckjqDFFmqm1szqbdlT8XlBv/4WeUPV015kKrLcPFUAp
ZV2zbhuffH62y1HGzZWw342W/80NNuqqCSj9UsgRDVuPlg5jiP5AMAsmpKoJciwc
jwOzMwqrpNxRgEmHDIUADXd9J2PQxm6jFdM/B++EolfdX+4ZEbeoC7yEIWe4CLt+
GSERQzVK+0gukQ007wyKNKCFVWERTpM6+x/n360CnhmGt/jVjW7DiWDAEj8d4mwK
6KDxekAD7DurN9vBSGCFOPK/S9JO7qLfkdBkw4yrlW2MRmFRf6VUrzNiZ3fuUL5V
IoyXJWp4CzA9mAGAgBhCXNxgkfEfsDkGBQ9Wkk7yS77LUSEPSW0LnDQmx3xzTDDD
GF18MDVcqKRM7aZhAAhdJUYxgn466Sk/+Tio/iyENAos4Gxb5B+eel7E6yE9V/lD
iPHAa1U6whucefu1PonMgWpkFdIqE31E8hDVzR0lgAEvrpTgMWu7oYwDxFdYrBwU
LEcxqDaJv3YAtG1PrM1A409oU+UBVUTLIQrv7utHLkzndhtOCe4Pw/hhuAEztoOV
j1KFyCHpjYu64KBJrculgV+yTyFlZysjNv1Aa1iTMkqyI1bsMYi53/Hr97bh3+vZ
c0EVomWU71369sFaY4Mm78XhI7Z7R3xMJw+hQ+7hsS0BAimAMeBsmgh6c45een+V
zj2yhnGVXxF87yflWW2XzFbR1rl/Es/ddB+Cd05UlvSWm78vscu3Amfg2voo1+oJ
5r/53qUyjBEQCq5RGuJJubUnMAp2DdFPRTf+OjQirHQZK/Zo5Ac/X6dmrIH0FHew
3xs3rVZbvdRMUvyDuV4J/FPx4TNuWFofcaVXkefEGdM9et6VLGis/uUubkYz5Zci
weVrh6SjWMUyjM/6DzThWjBvsbscHEoDD56sdKdwo3KebUvsyizCRkclQ9nLHAKf
/McXIiHT0gUJQTDeBI1plblSzaUoRzVWUdenYqvBjQMcLU1u04jCYH1aR/7BejhQ
90CddUsXPJG1IpneBTrC101dgji786z7Hb/QH3xvkuDzwz0XFfDt/PR2TIlYD+52
nveqJin/bwAMuLCnZXbXSRpeA0UdUDGx/NudSWzz9f1i1bIW8j+EnhDSP/jvv1Pw
G7dRls0LmZAv63kNimiSwWgODU1PbXrCGTAGOl1NvTJ/0TKUpJbq4ErKr5I00t3n
lAbVIdE205PKKKc9hRMoPMc2bW2lqAvcgewIv3qFgmalqF37r6PaSkEA1vx8r2FD
0yYVczCExFcBpmw3eU6QMDlEnQck2a4TKv0/aK5dnY4bEW28LJH/1rbOC6B2vcpw
SUmN+AmLbcEODdHHKkt+l5CaqvQagARX/GdYciBD+kBy4H7sIK8OeHsbQE1DYXPF
y8RMMNDzq9oKaPoKvEpZEha8IyuKQAPxukF7rWD5wqwdIryJy1u3P3Shi9cO39iS
Hn8A3Jo2r7A76ryRbTDS/q/pDBwG13R4dAUO6yqHsQqsC34RMavo3eJ/ZLoexUF5
zFBF95C+6ZWerUCZWclCLZVeOYJP5HdMBpvsBS4HJPuQr1ZMGHwgvhg2gW2fz3cI
vkEGjisQ/C1TUWFDy/a/ceHVO5YiP0Rpm/LnykRfI1a827R896YgvFzqEArlwYDz
Wka6KivImZVhNIybYdEi5MwXgI8Y1eF2BN8uCiut2RYNVm58wUaXr5Ij+omLQkPl
jGDvo3ISMMTZl5YOTeR/rTO+Z1do+VJsA3WRlGHgQrpq7LPkp4m5KIeYP/31MJd2
znZ8k2QcupWIvS51A+YJY8eDQPGcHd7DBhT/9TSTdUwXElxfiOHeASZr6Hy/xPfh
KgmIZVLXQDRp2mIMPmw2JJNBr8P2SXF9ODNgZUiTDQJZexdZAtcuxWFWf6ceCFXa
TXua1SGaGsqsiqoGjGPH3+AjWkNia5a7piTWAQ5O3bgpujkHIT8bJUXJsTuUGjgK
oQp5bqLpAZw8cSOcfrsuc3Wogk/Szr31BG5wG3DrGGHmCiTjk/386NX38HT05LHt
1CQGvZsede8kotCRMOSgK/Y+Lyn9FwuJIxce/tVj2IpvukoHKWE9fQBY926Chq0K
rNA0hMD2i6rBGF1EmhgIjETGB/NRSB3g/f5xCJmsDqrtvzSWp/Y3celG23u0QL2P
f8hGGyj62HBqOGV2Z7D9VUPWBTkrAg8GyQyNmQUUlsQceAIp2hGD+U4+O+pJfmzC
afwacWNOI5dDOucu4DvzlQKZASlFmOkQdeKuDTZdoozzjLXrHc142eUVBlHkbdxT
XKpsNDpsCs3x1b6/oIxQy9n7SWNSlSeK70aQfupESARKgoxtHrlD5EyNUnZIgZAs
wvgZX8vciZE7wuFAOWezdCBXXbXWfWL9kivOFIRZK2XcsM2kGhqxGxjM8szlXsVi
iiVYDy+CKlXhQPpK75JHzJt0gdRC44aIr0ePgG4A7w1cBe5hKHjqb4rpN+cmFJKQ
fjDj2EsatO7wjEpW8WPRJ63v74/MaAfbwMPwwpE5GEUMudu2DyVfxTXDzzYx6tni
Z71wNIY3GHXy+PSOjS0IvYWvBpFdIEzj1IbN0K7t6RlBGBRnuZgTxb9r919z2ah+
Df+JBD9hM3gl4LFq87bnqu4Cl9Fb7f/FW9DQ8N6JjOXMyR0kajXXwAuzDxFocWq4
gLQUnMEMuLZ3qrI99C8M5isnAAJyVk29CEDdvB6Rc1o1SD6drizUiDdas6TpLzRJ
mjTF6USN13R9wV3ppTtA1c4cThjZLYvPYoBxlC5vTsuWflSR1c2Onsm00K3Cgej7
3KMrwrNahEW7tmDKRqstxZ/15qDhcsNzcdvaqrfCc1rmifodvW/GvIDfkKhqW2jX
EpXpGw62WUzKIKEXiz/hv/zXzSugQXUy/IWS3IFfUyL4TzXoBw7FHlCxfY4Hf838
A6sZ6KIAWeTR2GYAFKUQ9ybN3KQmtG483ui/T97x7OEI7yhyEfegPOl8EslVZzYu
/gaGoWXPBhGllrrV/GVy8RlB4ZJGxwm1Girg/QDLm9QhOexooAhx4JEIAwdLDZow
R9Hm43xRAf34P4v3JUNL+8nc1FSUhI+9lrHIt1FF+C1TUaLhhW+gA24P8aSWRowV
Iyj4pYE3Vjv++wHf6JSv9p8u/di99HDONT2PWyhHM3K4wVAeiN4MYbQtbT4VfSak
xQAbDEvCLTFnjhpFavimIbJudkUUWWaV+kE3p7E9JC+QPzSQKNW73xe0mI+XZ+OV
vGb6NOW95Pb4TC3fGhZDuCi42y0uyWHlGungGYqOgcP63oO8s8EpAMIoFZCGu/tc
Q1AU7DWRxJJ15H/vrGsW+24rlCgE7Q9VxSU4dc/JmKjNJiNztLPbMUjoxcKYa3S+
VbdHw83xAguQsUA+dEXvl3n2Hgh88Jmlp1c/umx4sGc7qgGhyvBjv5ZeTruPtsny
2yudey6BHLTWKQLjANkvunNEiFjSMcTm69r+lMG2ck7dzmcK7uRqG3CeGDcVwFxB
XvP3xUk+FAN/DsNyYnllmt0BMysS2cZln7nuROBqbtsBGzvcmqGyewQ5jAvWV5V4
YlTETf5DMZjpfmY+Px/zSpXSs/LyFeW3IDygbyCz+G729k90VcbzkmKW7fhn8bec
IPEn9XFOi5jeebjbKh2gMnB5EfIoOkmhtol+0AwBZ4bbjJ9a3/iCAnv2O7YVRnRX
wWgF2a/1K8k+b9AViVwSs+Yq8sKbqCDaMnMava0M5h2BRnIVzontIS+D525UbWS5
jx8qM2yKXeo3Ej+4sJO1JY5C6wvjq2oMNiqfNOSHdFRDnGjYg2l1F3d7uqyTaYX6
4mJ+YMiZLNdnS/DsYOg+M/2/NlCnewG7GbtjCSy07ln4O+6b7bYpsiYp9t/+eiZ4
0+eTAtZ/nj/URLaWNLlJ+UnxUvF2V3SoD9KHZ+HK9d5466WaoEpZqjPYg5W7z1zE
Co5hlUmJehhKSiWozYomHDi0+bqrTi631eIXflRKda3psfWomLC7rsL+NIU7kEBz
gSkoQ8WXjyldaVmoI3+ZVNQxJGIq5kc5Y3G5NCsEcIF++VQBvELcm1mUuU7i2TsB
GqCIYZuzv08P67Mt4ujGTG9MA5xBQbku8/CUTNwac/KH6wrMjNYc9hZTlPvxsZI1
uhGwXGqxwRlKCUYmEALMqYeCTrKTGlXJe+3MPIoP94onlBV5DvXVRpfcEZsWaxEn
pgWrGRHBrjYCpMBZGGBxIGjEgDOOLj5wP+hcxgaklmYYKRlHj1PNs7cMWaq5DrBd
1OZlrW4jVXwPC/E3Xwkas6qukwP2kshVV3THOmTkA4hvqM3R+zYEvCrOxd9KVt9N
NnoiKwdf+K3aVD8BENZ2I7fKXVSy59VLu/REctkE/hJVs1qfCL+EV2XBARpaz004
ksvqXI+fCjZIxEzb6Faa0Gqafjcf/R34A3EGLu+/P72rzaz1G0T6csxisoeJR+o3
NqA11yuyd2TfjZqfR5SjvGWfcr/VZe9olRqfIEDNsn8ggUbTFUEoDan+UH4I8Kao
MdGlOq7OzDm+lDjGhfoEwzh6+WHUkvtfnc0kwN95EIh415s0MLdqURSrY3DQdx7h
baQEybsoP6q7OCGfdWZlvaMjkk7ZnAx4B5GqF2faWEgKkaJAcrOto/O4ONcDi239
ka0F5K/yofQkeQG6VsH71mXk2V/2iAFzezU0wtrCMMK1J8Bn+zvovU+i7kInqDto
T315xgAqcrEWWayOhefI6TI3esAcb4xm41FoQzhOeXUwg3oj0aJHMGOdH10+FrZN
tdS7SXKBRr3c7j2xtXRLMUK4Wzri+c0IkSlJ1cSc+ilxrPf99LfLLhiijApwRqr3
FrGaMjkdvtaG6XWJdapccFyvaoBTfyDPjKbFf4fbJnCreMu/4kMMqhqTu/cPN9ED
JhPtklIxSS5SpHS+OPL4sFFGC6HaZC0k3Q+rfL/WYqDRjyMnW/EFVw6vnYiUG0gL
DLPj3g5wh6xaB4gqRET+earkAvMdXIlEY6EoVxG3OivChGdfkPrWUUn9CTUxhf6Q
KYkWHYL+Er05Y24DgAKP13Fuz7696/btux4KXuEgYKy6M2MEOm7lB3v2D4UYxEoU
PPc9jBNXeWYbBdYzWTIupcQl3VShs9RE3Pva8LmoFfdw8Xw34zAK2q7cKi4e+3ay
58+40F/MsYnpep0I94iJzwowEtDhy15E4QFgpPQKyfJKgGLUs7/luOKJMg/kG6Aj
l9JeRw1NA6opzG6+UPjbMhK9EQZJ8juT/3tnO2EmYJVufcbCASESXRy6xo6w++n1
YXawpuxKbTe7t7zEF7x0vR1k9bt5RYFxhlfFp6xWq2mEpdz/79zueCdI8clroZYI
zh6LU00TYwUvVGu80evy/lVGQ8sEUEqlI5Yz5nxZN9CGZxd+5jzGHBdrBTZVtcVf
bpv7OzeJwB5u+uiuO24oaSUWuPpHH4cnxpmaNWlOr/S8F5GD1omkWr1L20iv31MC
yQ2X7s4GeH0aPXFBnzoDr8xVoJrHuG0aD/WKBQ25NpIMJqz8KVT9U5mVHLF3OwzO
tsnzmoUFZy3K+aCobsYJCQFFbbVnVIyKAoasBE7j7vonTGN2r5t4+xrmT36LnDPm
24v8MwDg2LtNj6veZsdTU2WrR4RakV1stSBRLU4Sztlb55BPqfg8ELVUXjGdqbCU
dY1ixCsngN9lFKySnvQLWh9AN7Pj9r17XqFII7+48lfuhISLI9JyV8ypPhHChKqd
NUwBf+wE47OfHFQmivQlYVh7hpiOutlAA4qu5ewdomJLnspOp8tjPvrh9E/4j+sJ
4nNSqCmf3rls6WNCzUNXb5fAcGeNOKT/SNsSvjrJEB++UZh2TPH5SYYe0tPiiWl6
z9W6LQV16VBSKKP6SIc5QkUvBf76Otd03Vj6dy4rNOA1MhHsQu2qVnVCohv4Dyak
dBog0VxieE7PjOKV5OcvI6T2GjFUU5v/y42k7GaswTQdffODPtxKqdjKPEDr0RCH
BBLI1tRQs63OsXXUA4DvK89mKJH78uAZwMJwqQBNgDYpFylpkysLAJ8AsWbQoBAf
5m7BqHkhUxadAShCmIUJdkPHGEDjaHHwMJG5U7UNfdKtOuTiT+Y725HYJtePcJM6
MFjxGpulJGjA0OPpba+oNn6D82RcVHwTJUCTHDZqHy21Cjqz6NBmtvTkGhrc8ydc
DdnJDXocEPpmFcTlikmhlo7hc0rNlziOQVsn24EHPAI/PgIdea++zBvxkzjXjff2
zM8TF8+tfOt2xJVNyGeiOqnpWwt1AcGRjJ72NCWHcNnvXXB8Wn1x0YJud7WoSF/N
10rcK0V0UyqnXjQws/XN1aXluzVwUFnQvt7jmVmWyXnMsrNJCuWnB2jCgzj/df/6
CtrcbKFLHTVMTssUKF93Jw0dGNbpckfpVezIcRWVuwZKf3J8ygkGaDMRtX7eA9DO
4U8BtZtffnpICKWoOGDdvY7czQVSej2kibKpIAZOGoNXhgQzAJGR9dvFNNiUODUL
dP6VhbxSpq6eniDkLpx5aU2ImROurifmQrNJliUp1iJQ3LgUxJpYkKHK9hjAPvjM
jMuyDkg7pE47CYjjBx3mSpC3y/iX71offbCr4b/v0EqnFp9KveOxzJpl8elpg50g
XWgS+cDARHi+b/eu+PU2ynZCBWuw/05wS6uipPrXtcpwh7duY94iEnzt142DexMf
ZPEBbN+Wg9vdS+3cv14qfS1M2f1ixADipv+S0Wy00TtUQOzU1K5audv0GDYSVV85
PASBxpF/J8Ee/Ud1m6Nk9NlVhVIGTZptSurFYvUPEPE2KwVCZ9xo0E1ZjsS+yQyb
nFJ+Nn7/hnzClgjJMgvl0QvGWqwGmoMCLaj6CPHw3xOGeD5YaSRqiJJXi+N22/Cs
FnbYqwxy50i9FpizNvBNk8T91bThTEW9Xi0QljGduSq0ngwr2/xeRr4jutVce3pR
gWYu+ATReugGlkd1ub/snOGj24tfxvhqPFu8cDI6WM7RO3l44v6Pzbc/genfr1mV
qYyumGqX6jUX0FCzr/rLWTi72/lParEpCJoOOmaoIT7q4nfd7w+aww4z+k5uf+Ag
mumIx0TZ7CVtuaxaWv8uav2PSwwE6DjG7Sg4iXwINZnDoVvol1PLef52vYMQV+o7
o5R0hwm+dV077ivh4B7y7Je5SN0qG0D/9eV5QkDr80OcyIYm31HyCJH43B4mSph+
pEBkkbYVz63l1seR1yUTIwzazbs7VCvYbRtxNByRypXj3lWqrMmWsWFN0X6jVwOs
ZzgeSCImJ2LAhhwBsQCgYYPqVPM5Db1/y9KlLAq4adi59RLShc51BfbT6Cc6qHfJ
AO/cntW7TmHubQA6QiN5dg5liIGnEcR3LQwDCRuuUxso3t99MLTZfzRWVrn9Z6xP
TexD0UFe4mlnTaW/pQI3ai1S8zSRGhskYMCXq4GhX5EV3WEA7FAz49FFvNQf7paS
cPLVvlkgHs5KmtENsawKEABxXtM2th/1cYQiWvfWwedR0rwDViM9ra0fEimGh97R
6noOyq2zVNf5dbkzJYCVxG9VCREcySEFnrdacrq8f4D13/N15M6KHweVdDVpAFYT
Veo7cDzeBrJhg5mdqA0DJJv1Rklz2e+rzUY/64Uy1DkrkCQ2IOkLZAhfJ1fDODjz
qsvgLhYeoOmj9SKfEpNGMMxtr7LJNeZrt/3A8rXMufDgQ6e8KVhOKdcZrBvIv7E6
p1Ar14WTI5hRjth0k6v3vL78uh9ML/tFlhhQEHnUpNYAu5Pewija1jfkcYX8khhJ
uLP+e/0DPy0eqMIsBpiaMj1q0YxI+pYWN33XI9stvbq4DCjcsxggtJXFEdNvs6JS
DfL3bpgCCXq0epoWN6nK5oouPYhg8sM2Srw9Rbf74WmTPAQrE/KMHU7X/SrxmZY/
J2ArN8RH7zWLQTwC01tXzJJG44ily1uFsAmhxH39FA3QFq16TU0B2GSGE+50fG5a
hHV9lokWkcXIohbyXEAUik5MlUjM3pLwBXFkfF+iY4WcZRWab03GJ4CvlmBznEIl
OkyVRWSQHeWzSQuIpMs8qBLyyOHTrICJTyujMBptcNS7b1Usqj8s4kvYKF5nKwzx
rVeAoYsSI9xx5f/1jiTl3Ww+oofLuDvQ/Iki0RsG8h8GoIX5mdaB9DmlEievL1gk
jnP3Rfmg6vnzjFWdQPBn5dQxog+bv/Kltx7LyiR3w7/Sy4/nHeOxqQPsKr0NIfPl
5zMPQptBL8UY/IcTrzZQfRrhr3dAs2cWHs3Zk6Iz0QghpcQy//Y6vBMfetDJLyd8
TL9xoXrOJing4I981E1jaA7rFWMGMX5/mgFlPO95a6dThzHqivCnj5wknTZ7RR1m
B/MhydLa5+V/qyguXsr3tA4XoobTBSiIYuZl7uBa1Q6kvhN9b8XBjHPAyUc44RNm
iv6YrISTgzZbKlLPlHv7Qt9PBE/d77QP/hSZkNz77cFeCzAuN/970FGns+Mgn9cb
qGH8KMDiDrJ1GTP17VBLsBu/kX0auN/lyFQ1d5lVo7Nxia52v8chBWviZC3hXx0S
+HJ65pm1zQpTa9jdw7OUjjTzceK1m1r/7WWyyCXSGDRdyMuaLQ/J5DmmngrSo7vn
7ey22H8pIxvfv3EeimGMVelm/aZWzWS0N/EFIaczg5UdsfRTZxhwXzNE3EDo+Suu
LOlHwLnBeW66jFvbdoiM+BS5fKsNu88v6Lqte9+l6nEziC3/ePT9zymKIAOiV2vn
K6oEIw61XSuT0DuFB0ekON5ukfNj11iXtErZmejOlyf0qF7YEvM8th23vDPjB0t4
W5n3PR34KUGJXJn6yNlJibZmoyZ4TxjYdRjT5O1AS07M+i7W+SnWJlIWD7SHjP5G
rZTi1v39KhBEVDcjY2JpTpvUGR0kVtzKF/szw/OysyFigQfLeO+h+Ito4m+Spz7B
c0OaF6HQGEPc6y3YbHWA0a3TFPoTE19UuICCjOezX30VmIEqKvTj7NKglongz/SQ
98eU9V/1hSWCvVoetpZAdls4JUvMuN1rkDeQZMX8H76P2k8vd1g8Czt2A4l4p5Bb
1Rr1fFb6cXzapabTHyGz0agJITmKKWBCY5LltxF43voDlvTNF52YAMaRjTQncEWd
GlNRlWpEA7q9BpzDNaAXQsNRZpI/J+3xlZgKRhOMp4hVjAOMH5f5/jmXW1hZ3Rgu
tX5rydAwFvxyjIxbu1GFW6Dkam1J32pdMhgzOlJ/fRXsoOpjo2PGrXOIDJTtr4TJ
2Oyp40S+rZzR5AKvZz1uiQ1fdUB3b+MBptOg9Ml1Rt+qYuhZSBt9BJ/IvmbS3/ux
5arxdtfa6OWMJsAgjanCluStm7Jv3SBmgTYKhYnbCPLvqvZhbQGQQQfM3RFIMdfy
cd9xL5nknGY24aSpnIqvMmoNtCE0R6f9+3QuQvGkCkudzLNJBJC439MCAiOXo+F/
EzZda8AuRavx6vBUboCUSZd7p2HFC2twsiz2utu3Dtsm28QOLFHUhTEyGjgCm1AN
1vVJ0cWcSfzjm5sIppg7P1xK1/HN5+zdw2rLV56A3rYmFv27nTk37fDXRZydx9VV
ECoQSo0C5oDGTM2QbOxoJ+8ZiVwrb3+eDQkhnQf5Ddy3j3zJyLymJprpyn0UF4zG
fY93otRs6e5I/i3hBMFh4nbVMxK+t3Jp2FvBtyFKqEBxnHKUN1TF6za+cUF9/3I0
8bL9rITtMVy7CpDSc/z4fHJBnBk72XMXqGrYogWZZM4I60wvRgdmSAOv9/cMbiKP
bPB0b8GZMLe852RTFhtuPz37APRMDPcGH2zEJ+lDPFgQLjp6+sf1nn6uheFFQSSH
PCzztgwD2HwimVSwln9+92RZxWy11jvbbMocYNP3P0s=
`protect END_PROTECTED
