`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5iduiJafcNvGy0rYm1PCLBD3mDA6f0ShFCaVsH0gZFEgkR4wgAh4a5d8A17hGOKi
3XMZdfbnCJBaHNgHYDLnHjufU5ezCWmF2ikxtrpwtV3GWJlGm8QtR0DF5d2NY4rd
rD2HYXd3ZtplgRCs7gKGiHLuV/FVr37Rb7+Re4/R5QtMLHNcoyho3BxArYeVn+rh
d04Z2onuq6J+iBs4o/H+Fzxjy/6YDjsnndNs3/RXmmT+geRTFG/wtJAyhFWeyrIJ
7sdO2BzjuBc7cUXWDe38jnTD5Z6QIKGVA/Aoer6sbVrnbEAADMlCcE0igOkRuHHn
7n4nrJBPlHFfR4uGLLb8XueKWyL2Jq08H3knQp/8bYqd3CCbWn7iChFrZI2pk0LS
rxHBPeMLihbipGRmzLD67Aq1BdQ5RA8+DqmEDTK7TqiV+HGGFpxUvTxGVuCVY5db
XHPvglX8X3KDVN9DcbCzhgE2lf8Hx7vVhKkzsMAON90=
`protect END_PROTECTED
