`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+5XiJO0Uh+tMJMN8xMuoTDqpdtuws0938giqE3y2ldssIlb4c5Wz+suDoGkKYIL2
Qh2O98mIQo83MGt8i6RNdT/TJTosi5hnKCWBT4fiRM6RCHrusjzGNLmhWp9mo/ZC
YMIUsUVTlJcEk0J09kwbFn8pfLDnP8LTqMLpMmgJ+adSlhUL9AJVj2zEL+85PuCR
M159n4FJRr9SZG71Jd2YLcv+G7bu6kqRIMWod+YWuhjYgKnxEkN7hzw9mEEawcQD
J8mO0XG8s5963CLUsffZSrlL7e4K90gLW9t8gqV28zjQHbzu1U+P1KDAfYn3TGab
7RyDo9qFgsNtYRt9qJYnLKAurVF1yvd+wSTu7ve5pWiAC60OeHadKbGUNubFQfl+
5IzLGywBxwaGNMFWzonTrYQXqTFDHb4yzsZFKHJCJGi1DyIiWFwPAhg/PZayea29
XMepmptOeyvDSL/pBfjYRa4r75nZDc3bKLopDcdTFUVUN+eNGmzuaRNpbw3CdQU0
TAHfbpxjauD4ifYTSLAkx3ZjXV7DlnJmfQK8pc/xqDMuOtpg1pA5XAWsHNB+c6/w
5bgn62OJ15K1dgUBAhXUMy2hhtZ5jQt6oABxf47JZoH646+9VBQofWs/5kZJK6/t
uDuWHsk0vwbciISjdcgNJX0OSsDaaEmWfW+C+sXeL1X/fTwz6f+wEV2KCtSoOjir
T6Zr0PmPJAPmB4os0Suultyr25Sk4Yd6TFEk+xwOiDJyCCnKmRtHPwwAh36Hzs3l
lSpg8NQtHD+GRBwKrivi5/CzMRaEmg4iNsbn2nYdW4XW5y8NH7DZML6ma2ksiYBF
U2NyqA/BRTlVffSgXINW6t2R6ShMJpvpQfqQTqzTflsDnDXby3Ed1bUGtGXJFrsi
jcf88swkDynLXXLRxufthqHtfOvE6k53zF83G19E6Ix/wMZRdMC1YPBkR2i++oux
X3y9Y49DXykILUppXWoPehizbL6gi3JAmEWE7W757Ei3EKyFSRgVysUqMXB/vE8X
EdNsLSL9YB3Ekupq8Ywj517MgY6i65dbiXXwn/RNhXjvVEKimxJhMv+3uWhq9Q6Z
UlvSCsb+BW36nByHey+Z2YsXdaYODBR65nh1MjuOiv5v534qHguB8beyZleu6kSW
vzBYocyYCeyS7gkEMAYU9uQgysAmPQC0eT2cpd7fXHeK8YuTqVxNYlICNRqxQJdS
xNYlArKDeonGeZIui9ZFgqA1WQw9GPeVit64CyVRIf5CE/sR1byeigPZX/Fh1MWE
70ceVmbqW8PhnC/YaC8UMeGUVjqC+c6SXfuZ50lMW91o1fJCg38uQftM/RdFMuMz
rTHVaZbaHc971mfjghOqIg54Zhn0Fssq6lwAPA591lLfZYNoc5HLXwhzeSeQw/Xn
WueP0PBwhN/mZLRx8DwAaHF7ef3ADpyN9DQXxL+7j0UWoikRLV0zaMTZ1r0j8VSv
j4/VkPPYNVPKv02WEAY6PXmcHVtKCEiZhNw3phtkwgg=
`protect END_PROTECTED
