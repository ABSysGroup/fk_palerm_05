`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Py27/4cb6nQTr5uQYgCQiSgPomSSYRw1tXpIlXoGKa9bQAtpC0LY33UcFsTLSid3
niimYT22nPhUIb7da6J9meTkzQqfE0IML/RJMqzOS7WtTT946/5A8sd4C4GkZnje
ZOjzvOYg5BXBVlYedesCF5WBKTT444jg9XHieML4C1DUGXNi65qQgxS3Rp0aHnGG
kzrPG1spJTPMuyFH7AxOnmqlf6z3EXinuyib2ukXg8umKxxJgSurGB/QyPIMJlwk
NuQDQNUeGArkNkquG1P32cF3JdDtRHmVpxPpMUWZNBRYf3AUQE8KuJcsHwUpf3xr
889v2DkMYTaXnz5hGDy6+ka2+IzHl9ecqBRakGaTOrNqtsO/qey4kQn6Cf9w8SGM
I8HMajE+7JIkNiHWQSIU+ZlxuTh8mRHbOEssGYOIpqpXcPbQaNxunYsdGUtnvpx2
ZkQDJoiH9iIwjX0qShVXYR/e7JHNu2MRH/UCUu2Fbi5RkGQ2vIC2db2eE91Ehfwr
inkmTUuN2z/YCW2zQj1iKs+iTMii6yAOslgStUPYDPZM7MidulJXLvkCp1V+xhcN
`protect END_PROTECTED
