`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8zwTX/9CCaJxqqrcX6hZcOIEbbhaHN5gkf5E1qpy4C/KCgKadJxjB6/TC+BPfHFc
6HkoQBsoucdgYwpufz6FYX+MZPnMYfvl7GRW1New4uanowhaL7/sYR4fooybqjpm
z/iyvx/RSxiQMnR+gw5+r1C6RUo1XIXotzKqbTtPxbRRAy2YJ9XiIoJLccObU4WL
Vkl4AQgXR3YsfqR7b8XVIw9mfSVLROGKut5j9TdC7Y17zC2fQiNwMBRq1UnWLnh0
E5Uwc9/39b2880jDdljBc8h4wxWQhzQ9YELdAl40BAagXMZteHSgUI2q8FaS1M19
NuTb7VpLP0gvxifbxu8C4KC8fT1U5GxuR6lDSoP3J0q6Ek3hGcmKsJfNhaltw0r+
aGO3QTT4ChUaSOC1A8eDtRI8hQFX7UZJ+GrFcCRxDQK7UkIGuZWyAil/b1SYUS1W
5X/7l+iRhtsTVAd3Vcy1ckEgJ5On7/XHM2i5QuysDy+7iZFtUu/6sXG/nzhyY1x+
X7GtxHJFz4+DcacxsK7wGYxxDJsMJKx9R4lVHy3aG3BX6tg4YsQ25K2o5Y8lSfLL
zBD/QA38iQjyI/ibC53W5GUvoqF2Nv+DcbWU5Z48bYoUcrNDg07AWjdqXRiKRjC1
xoHk/87fccAFYHPwC/GIwS6QS+aH9VGPTSBJp1kjT+60LmWbgbxSzhbvk3b7yEcR
a9gYHPL+KHWZSvXz2BbmeWgm3MWCe7qfpIUjbuBZfwcjRVAsz46fnAATFGS71d/o
rlcFXeDJR1aHienhDpMhwmox4GGnGbrb5pIGt+hhI6JVAhOwTG5JmaQBpneDzWJP
YWi1/W52M5z1gQ+gbHEd2CTDYhbXQZ6v7UBq7vnUuly3w3e3Y4KcPQ8PnjYgIl+x
VxrKz8aRON2fpSYpV+5QMyuFiGoaANeYqt7vMNXf3kVMqhvRiJxInIPnie3cvmWA
tLNINS55ZdhdmXr0p1Ij0s9wIvfpbKO54CkfSlj1spY3DPXe/tySimnqA3PtVbnz
kDnHuZXdbR5e4CD0PK3qYO5AAN0zZ9oqFAx4OqqVQvQ45iKDZswuvICGz6VjtuwG
EuykhN1ch+JnRNrUYDss4VKSf8e+AsWp/FgYTG/5fTduPYpquGLyLmjSyx1MOMIE
dPWf1SgpkXGqiKdCefO31CJJxrzidsu/WBRsJtGFCgHDNesP+txrwSSmYkVH/vHM
r2KCtg4DAY6L11U0y2h7qhEIMMS9XF5HTdDnNFHPrwAOdd8/rR+lzx3v7fbHGfuT
RcWpCpAzNMz9pJmv68FlE8hzEKyxnbqbaBwVibo5XH1aLG79J/3LAZHq+I7hkbjE
bFc9d+AkudskXPYKsI2zQkl5ZmW1jn4/UsZI7NjGaMeG9/p+GMJQ4f7X1lNFV7eq
PFkhpo7nJdJUc82k2YgHcTjjKUKJ7k3tg29CrbhYyx6kDDEtREhpgKoG/fY4tkYG
JXuqfPC5PS5l2w9E9oYNLizKT5+m21Fv1/jWnSdOA7A+qbNA2suH4gXdsyfX3nut
GeE8I0Xj0usePSVwp7vBjfIyv3VklhCimCdPhHH0zms95jDnFMVDv+DI7pslDaWC
hlu98Dp2+9qB1hkdKS0CwxHrdAqM9+veyX6WkoUfBbxtf1OQL5ZwUFU7NglWzCM+
PMjV64WtvEYO7YxuXTFCaCZbPI5mhHD+3UFKgnKAHTfnXSMvDF8kD7thgV3DaFie
zXv2FqnGUsebqzMN/qa+wikk9Ump7XYe5gapND1j6UmMmio7Gzp5IW8x6lfSsJzN
lghR+DqEkJlqbPB3NqsdPNooItayZY2g+I6FNAdIteZaksN+1CkJYomowXWKFcx7
wV1nQGAR567scOqu5+SAmMzEjl4rHnOtykesxYzlptmnL80QLXDBeFDSgaVEa1lP
n3oG5b2YQ0nuaILAzoPPvU1SnAOHcrqWIc5huO7yAB+O+wYlAbXZpZ0icg9PvKoP
Lu2xGUlbcfZf9EiY2e/TBgM+guPDRYw6hb5r4zZUftlqq4cxv/iTLFEwpOomC7u4
rBe88sJW7PEAH3Hx82vJ+Rl+mCjEW2YsGLiX3wNYELA5DuJPJeTYNPRawpfkEZoD
ztxEMjWCzYpGhrt/6sYWt+87qkF+SijKqg9M1ExLrIn4+RCWx/GC1Su5mzztDoqf
aIM14L+MITH8uA2oBnyc9lvkJ8D8DIDyaA6TI6s/7V7xsr4KUWHm+RcLTQgjUJfo
o2jinEx9/4zkNsefBKTQn2ioRkS+QLRw2ShkCYJYWepdsQsv70V5VBYmbUpqiIe2
bXP9yR2wME10SdQSDeQ7cTZBe4VgP8tmzHjmuxVxAPPJjF8+nrHtq6tHQV5azj8e
H3kCXpF9bwerk/q5GFEJ+JYTZfcC6Sx6sYKZPnF/LrtbXWeninePQk7oaTOD4nSS
GDhrghqSRZsXFfjpy+fdzfCbdFcOTK5eTWT/2dUJDaV4nw/oM3sjt0o2LE0Z7U/P
gGkqRPLcYLAOekicpvCkoTEQU2dwnke1NBImsVh8mAdXN8/40GF1ubDnt6XI1wH7
vMtNBQufxYNdeCjbEyJH6jq7lhqU8oj7qtiLtrF9ZKO7Az7yZFdM7f27eMG2DaN0
mSE8kIUTSo0VC6/yMwCLuVIMV2C3ELsHLYwUgeJACQ/aW1sdO6Jn/5lQfJVW6jZQ
Nr0PNj/cjRO4p69welbq8Fterby/X4gTLFgJPb9TOE9SN79/bAa9w5G3GTIm4K0i
lcJNYxP2dxMpm/2gikkcM5tJx+KKmuCdFacw7p9Zagc0Oj73UwWCKdMoNUyWaFgs
SqWxFFQnHNbM4xu9kQd10ECD0pEq7//T8cRqGtKAnDH5qxHPALudgj8h46ECAjbQ
3mGsxcOgOnkJI0uotF2qAjGwwGiEjT3mCxmbakqdopBAGUgEjI418Qz3O8BUW3+2
UEVcE+vHEocs+dp++3f+WHYcI4uK7Ok7SDZCdqggLvtdMp/Z8qGt+JfneM/ADe+O
Kgxn5sxdf5iXNWRsfJj/UWJgUSTr9RUbimjCupRONkanJHR9jem0IY1GyxghAgVK
O322xS0cEJeA2fgiuHcW0P7RBR65S7WU3Nbq09CA1LE+5pIY/j4sG3LlvKVJp6r2
vJdKtGhjVpE3pyXrW2xuwb1j/E/bvIAyyEG7XNXMT/u40RdJa5TBfbWJgtM9EQ+h
aZFrD16zzrcRupaDbGkkBTdh2K8efmKkHDhUN3GcjVcwRMayJFUWfFKRD62I8sQc
vdLXOoGBc4eCaoDeamySNovnfScaFoqtbwq/RHGJRALYZTCSpCKXoP/3E+48U66o
2itMit4Miog4UX0rZ7rJ+CoMNXoC4sK5IJKXCJAM/Bm9RnG4skjHj8fZ3j6UWkGF
sV8iXcIEvpG5S4LreCqsVxLD7tE5zSbeF2G08LS8svKpWCYMuZB9B7KteOIN6AB7
z8/jmJrRO14IJAfnBvgwyjrCG0gwFqV7lalkR+BIGAU874A6T7E1Og6IVOWiK3gk
hT1BJ1UIHwZA43m1A+sA20i6A7zdRyx40i+V7D5JASekwoEqmig5K3a5z+QazL74
FlTkEy14ZwqRyPu/mxP4+hpq2NBhEGLOabTGFZOnq6HCG2gIJzr8ZKZzNBg6khZV
YMmUngoqWATWtt4hp6rcXPs2wsk460X8MAlHzeosPoyp5DuJ0/jpxSNXcYtJnaAi
lzeOd1RqXEAHqLmdiyhfsUAaQtEPkKUyUrt9uzUxc+82GefQ9mN7gSmXSWL7MIlc
DNMoU6GUKiYuAD0TwvUaN4DGVKMDRd6PyDoo9LiCFoMCDx94HkRhk1r8rmhBm46R
3W76clxCVG/hk3cSndA1IBgpMbpZRhJANFM6NmPKpUThzMvuHgu1DCGs6e8vsBzZ
Dhl7WpN0ZLktsGODU56TNGKUkgo1l6jR1SWBR2s/anNGO2KsYimJiFq1py9kqmQW
sJ52VQcgOMqyngsX5GPcUR9n6mJHN/qwXEcuckFmynGNeCj6/F2hIfJ+ceNN+4IZ
znZUeCEGLEqwgQ4vThLgTkywlCpDAu0nI9wL8qyZ1meUOMKoNWpYNuiI1bkkWzf5
80+pTNXlwZ8O1PkQhJbFTYYazAOvAK3fPuwkjNMTXp1rVnFA0R6tTDzOy87bSZcS
EwC6pflCIxxWtq6h3yLjWH3Ep28qa20DMulP6FS92wtXYNT2NZy7VO40VSApox5r
U5wBKu7PW2992KUCqLitsJ8z3c+l9qAqKPBSqYAr7/s1uQcyG6n/luopZY2gP6qt
yG2E/QaDfyF37P6znkCuMNex04FfeRRogkECKXObnfuMGbChHm/Ayac8t4qpal8n
NVF4L743r06Mrwq7DP9GoNPSG04SbYbK+i839LwXkcWb5dSH3+3caUY6/qC0WXAX
SSUxbkRcBLa7bXp46nJUhK5o7Q9LEHbYYYy6fqxFFFaK6MoqwVpX6vs8Mn6TKNOX
TtFSIX/SDUxSzyNzO40PO96qH5trLjdTaTPe0+3/7WZbQfRMTXpp+GPKU0+d4UBs
OByfdWwhwnZNlJoFAs8KjMdnJep6QbM3gcpGyZeEz1YQa9/1ddOyaCJpTqTAavf8
sIhEcfGeW9UwhWKWRKIxIDaamVLLxqgsGnaaKcj+AEJ28dHcc0Oqi+pWalZFm++O
RRFbujGEDwMhGQXViYjnlsavS4dYDhh/AszwRiQ32NeruI5wDDKpt95cbu/ESV+8
pafARz/YpHnzZU33Tke6ETWiasFKjZ2HIaSwX+IiZ8X0fLnH94kVVaNCsZnxLrYB
1RV5gy0dTmfod4V3h7ash1FVKHn55xKR1l1k+EOc0nt87b4ENQ5gU7HnbHIZfkxz
4jzCdEwkrWmMegHJFbtnzgdmmLiALw4+p/2JvcmLVs5Goiar1wgegWc8zU6rNBKO
K8o9I5NGSdBy1mU52Dze+DMkZlMTA+XWm3r6Fjsqpv61XzcqM7brbLv6bfckDByH
K3+1vvqgpY5VOu1TZyDzmN8eQTVOxVNz3wDxywhiXj19xmm7E/JPrGL0spjxoRtX
MwNVNQIWgscOafzp/Rwg3cfv1L6bckroG8MrJdSn8568rfz3RTjOjdqX8kqIVpaM
6n8TLyXN+/nwp0V9zBrP/+p5vthsd1DyJkH3D985UapBJf/3B1eepgKmSOCQ9j3o
k22RnjgqygMIEaprdMqHAA+hWo5adqfNqdA3cZ7epcGGBJycuHxgCXNzAuPZG2w9
dAprIT41ZZ0ciV/4QPjODqrdJAWOqdXQWFKTztBlhDIIeXu24dpF4XBikjI5oXEe
ICDJU2hOXuyHNS8efymuEGdKMHquvT8IBB2/aYxYmPbXGQM4MMnHAoy4qBg5fw7F
HS1PHXEDBw6HawaTU/Wt2wDCOh6MITtWMMY0dZEulOFC4UsT27BQ4X5LXrIkzGmR
GEMZNXaRK7Skaao2rc8r7vU8vvUyosNPyJXK9XXbsiT4mGB5N6pIKYCOUqS8vVyo
gwH+mWQLiPELv0G2bcslrjGyL/sJAg01wrZX0Z3zQ5L3QXra0CQzX8pvqT5cyAli
RFg5J70nQWDie7Y7SC7RTZT0s6gePG7YBNd63Qw+jmwQKRMBkMSSdbahREtfAi2S
9FGdYtTa62Q5pW6KYuBTAvLUaWkdOKrqz+nG//TGvqwaVVSzo6mraWTbB7kfJJIZ
5FxqJldOfwjqG4QFF4rWDe/KGqXM3DvqW+2Qm9M8F64YnmZNWXwZPmW9rxaGqlIO
FuoL667dcpWu0Y4Ih14Fd4X8wKRdpszClg4DHmr0aorbEq7A9U3YtlZPtTXvk6wX
C/jpwQvvxASYResLPaAxUMkhxD5VYmim1pDMrVuc3y4JEFm8Xt3STSW+KCdhET3Y
Z1Tqs6up1J1gVPpLp7g+MWGAQDvNN0JHY3Du4w7C1uDhk/a0OSwoBUafudhDLAnT
JI7/QCW74WifYPAetWFgQSElbhwWTed8athMVxF4bG+xSQ/m5K365fQPKeCFmFkZ
/Pfjk/GQuzGXC/GDOuFRIIIVcgyvitDfHXF89mIuy3J7DsF0vaua4FSRG5ycE6Ny
4AUJ4x812w7K8xuw2gM03SD0dMhvG2UJv4N5fxOQzX/5QNZ7j+ObTKKNuNfFVjtV
6E4C2A6zhGnzOPVnwA92x9cxfbzHxvyrLB2znndfnnFLt4z7WSaHXzLk5VByU/J4
jEfnnuNh5VzDGsTpxkEJ9v9BVY0vhVuhWk36ElaaT/u1s70QLvPFMImsWC8yRk0D
wzk9WfV8urKpBat5zMoy7n6wUzWW1qR4JfgZeyOmj/L8QEG+ZVbbofciUN4qYPiZ
je5TiyLI6Sb3bJYjPlUe1UKnsuYfEcPXTMDxMMuYITJdE2jPnH6rU0vdWvtF+2FK
LrYAROPz/Wd5TTih6z2H+Sb4rU2I6/odMyqvB7lnFnnDVCmo2dc0RLc9r3iaCNbT
P8MgyFljUPr7ne67glLku7a3mxsJKwCWqVKP2FI1A2cey+ER8kM6Ks9Q7Soy/96c
cM+KxZ2Gn753tTOSqojPqWWw1dXQUxSoNHJU5rzN8IXE8kSqMCQEC3PKx6t1LWPc
Ir2bkBIkNzaNNTMEWE2M8LbRgrx2zfzPpBh8KGMb5wGXM/nZtrLvo3xEw8jcGZS8
MdBX+n9TlfMhvfM8tGJzxPRa7eiPp/+cXNCp7/4evK3fVlj78xWijkbe7T02qriy
IlSuQparJpGzFPukeOV7QkFk9ZEu+lMFEz2nC3ky2ARyN0WkSFzZBsQKWwPS35ia
zqmW5Z4nPQhpdmply75WOm11N/P7MdHJhB+pRScUUf3LQlMVn+FglLpnY6cdHR4o
Y0RiYD/qpUarJ/Enx3esr1ASD6ZufQvQVpZa+iMF1KbH1Vz33+xzDTmqhTRECuZi
/tv1rlIgsMDNTGbCd9/3e0PbKu85X9FWkgQalo/ggCKX0cVpsr9tKu+sp4g+kfpQ
3B4Nb0RIOZ1kZbs7jiK/kodc3tIICVtH8ggtBQOwOT4bgqVt8JUQQaNhuFk3JIfX
juiQtc3RNcunBvgNco+tN6w9U6Nfzayyx5XcrCLbjgzVITNM46W6GsXa3jwEhn3F
gJwZa/bqPRZOyGb7YGGHbQoh7Oznm98JxHedkrmOgFetngRr3Zf7IOwnkUjZZebz
5DzYVbQGtCBQhzk75hbN+aP1hDTWCf8EJkZ8tD8jqKLzczUqEE384AJUnvM7dqki
7IXExVMJ6zYr1bqU+T4vZLWWNMZmHwc1CsB0obhorOtfly5P3D/YvXQ1ak5wwN2E
AxpDOnn7B+200UX1gXQ2HmC+e4HLZQVlpYeZRIWco9O3yOnGgyO+d0k8hQWg4CQ8
xlpMp7zN+9nuFxK7WDFsU6yzKtO2MO32AELYQ9sa9A7ogFQxEShneOS+9qgseY/q
S7hiIYt6xJB3lDaJ3LGifxLm+LjAyialOJR7zm7bb4EM9ar8TrD7otjiHFrKaWXe
qEeBnNryQ3G60akd8dtER0qovgWSW4fDKt1nI2R0uShIbkuFJuz1Prner6f1bdBU
b1NKJo+Ri6zUeOO0Z1fPddv3vL40jWAC+82Ic91C1y24caSGGLZ+7udpP7JM7P+l
Nl7NPyBpCiS9sUADq/YirEkl64HxweIKYE3zB+1dM3IiA2FMJ2UjK2o38BturlT1
ym1IxyPwe0eNw/czf3RiWGm8kZn2Qyrt8Osv7utkcMfg0Hc/5J7vEGyfSvo8TLaa
ndv/xkkybaQBxjCBq9dNqPEkp1OHZCb/VsMxlU/5zhW3YuClDKYCgKR8NCSMsNAE
F1yWFXgOXBFGJseEsEcuePHkpl5HKrC9jYZd55lRp6yWGRVGn593hlZ3VFNnX5lc
dA0hsy/6ZkjEPCd3SUDnJZU6qvUckp+MbPmA1nEdrN5VvqGes1M0sKE52xBxWkvx
Fg5f3oavR3HP5Kxq+CQUWTT8De9JdXrJNKtuhRAf+pQeaToASMgDmYYfTAnL/l4b
a0CfPIXwDDqqCZKcP7RV1PPRv9vz50qWwzAwFYuormZkUhw/PHdIaqiw5/gU+4cS
NT7ZmWQXRt1nkRYydAjuIZ+pXeo/aU8W1bdlThwfxSnvVTGk5sqa1XBSs9oZFfzH
YepkmRbN8+2hIOXLtIgSg4XoPyP1ijmLihQL7dii472rkZGMj41LMZ6lWNi1wsEg
lH+qIkps5oGOg8lfp/TI8bLxm9yUBWilyELPGozEhj8v3Giq36/taNp6Gr20wIRh
EOH2UrPjp9+7sAH5dxDWw/vVGV3Z0kFfqWV8Cw/9jK7zLkM8pSIs6WQc4qslbokV
eIr57mf0RrmFbo06OWKjR7gVwhagwBD7RDXYp8g21q1k6KOWVpQ1Nvl48xr64u6P
hfA9A0VrcSUZcEXNleh3EmaTJr20Eoy0Gh8sBR5d520bXrbdNDwqnvB7AojSCLEA
3QR6LylrcxyyKOx1/uf3CLKMD+nJCsHK3TqYm6882MK/D2TD9aEVSTV6h86ETEiV
+hxnC3D1221YV8vGZl6O4zEdt2XKV5/4egyIl8Dded9Vqru2swSuVaU6aXdvyT9+
E2/X86crr/ZFf+hoph7OtlpWA1n5i8l9i1qVkjdJ3l9t4pyHTyZ+jbii43uOSNeu
9It/bkogGxGyI51xQ+w4yVuqWey3SW2nRiSjhtI0ye9637bQ7frHK8mBqI2DNcts
xxb0n7gZo/IMnHjHr/auIM9t+xoFFDc2mk6/ZK+nRzWri+zxy34N5+LmjV3N0XPA
VX+/XBh4AQErRwaN7E8kGLOYtasHQXfp+9oDBn7Wvr43HSPshDZVJcd9fMqAeaLV
R2+vV982TIfom44NHZfCWtNh9Imov2XOPP5a1/Ya1ig8T1uvXpWvC8xSJX1wQJ2r
5Ma07hGOOtf2awLWRQY4TlZzzHMerSxAyng5EGMiALIcPHXvzXUJatTNVnxgvCiX
7hzxwZbquGJ5jQnv/K5BfofvBX2QXnxEQe6nSv4nxGylxMnTV46GAgw2e4PhTjST
YWYZw3GtctDbNlduDfl7h0X/ci4YZDV0Kc5SIn+KvKLjg0HLUHc3x2NQ2AT+yHk7
lA01T5MPqZmsYzbkusBa6fiPuuUz8BMH+9KDM1JkCQmfEGeN0KZVRbTEgwDDQeix
sOawyg5d5+Ns7EJw27iJxs1DzR07kG47u8fp65w/PwG5CocJqUu0UKlFkdJW68U7
3tq2ND+KTYaPqdeCA6bDNVorJ18IRXfgwU+kYNGvluGtBJQ4Pjs/ps0ncxgFiZgu
Z9vRzCgNBJ47OWb0OovH1NFjTlBgTFKHw9+UiCsnPAZeNCLmnhDoBaoCvO37TgB4
Em0WF7MTc14cL/v6gs/yzgrOAS2CoRg4//slVCAtNeeqR+N+Tcn1v8bHGhzCA1XM
Nzrn07jwzf1ZHUrLzz6TrFQzdFeRoEcOlFhhFELrtfO2MuvBg3ekoYloWBa4lK2M
ZAmUoocmEn1jm23N6jVZHRb3/GFwhCDAWrYJ1APC4/YT8Eyqk17O9xNC/RwQszGM
QhgmhAiyNEmXRfn2uEwS6j8OFfvFPHMjYDs5JRovDNEswipcFtVMPokjCcqO5Rin
p+FgRm+T5i8/5GxMUfAnFFfJo82wlYB5VSic+LFzROY8o2aQzkDZGK6HoRpZedET
6+VKQMCQvDMOH0lFlqBgrdKqXKoB7sIbC9fTzlDxDTAVU/D9ttu88xx2rsVxwXiv
U5+kVvcwDwVlry5YaG5M/xkVViiOQmKuoCx9yl4+eRnDtZwd4OrovK9b4MoRXC5y
hBjpwQLI4N04uwrYPYllSHsfA7xlEBDJ4H4xDo+ZQZMNbNy48GE9iTCg25zxEWM9
4vUAxIGuD2GlkjBs6cOsGLbmMlpohdAVEAkXVfHcvYt5P+ky64+xHe720B4Eq7j3
r139owEvllZlNWSdWSsaLXtjXIrMYpoCrZr84s8PZQSiYF9EcbSETnUQOhz0aqlc
MAFNVltTetcKS6dZWfOzZGWKkiVQ4ERfFE+Dv/i48cCueEXl/4oHIpeIpvQy5DNx
o9ofhbw69q11eG03q4XVwUYPqkgf4N0aTCXKWHPsdJ284p5p7/yrnE2PPttPSqlH
XAPtd2KjmEEDIcHnP6bM9Q==
`protect END_PROTECTED
