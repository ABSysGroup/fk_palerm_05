`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mlnEiGozCdjvmxnC9erXGv+2LHqspPwjQHicmEv3nU3naIC2IW+KuyXBa1Uj/i2o
gEJ3p0MBKed5uxPDtJcfYuRnkXNYQt+9UH/UdnyVZTaF74KQOgs47KUPacpL92fW
1tORPaIYPwSfnOzaryuuxSfMU6mjmWPPdnz1Off86shJLMW5AddXyDhH9X9+Ntlu
cN4Bezx3Xb2PneHnfjn4/5Y1/fl5QwQePYXbQAgjXD8EezPKL5EoqVQmITGLAFyi
oAYqVtdAYaydexcyTIcFof7TbfYy5KpCZEI9LXPUoiopmcamr0kL59M6KLRTydvg
Wtjl5R4SD0PKg4n2SBqXn8mqyHZCb0ZV7OkEJTTUljuJ53thcZS6E5yXWmO0Ychq
J5bhsfTmSwNeSwhKXGVtPqT0CAxoMrDhKB5+AqKMW5C29WNwP5/L9K3cwDdzFpzw
lq14FgXguS812+EO/M1jCwxxkN/AmZoYA4g4L/tCxOvVJPZkMO0rN1iLW3spUg2B
CgGrPp3V8Dh66j/NqRTlRssesdlrW09eZ0w2WNyVtpg=
`protect END_PROTECTED
