`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Orl7YVKpSwG5Q8LgWAqCeZclsaz9rLE3eHlzhK6aTA897CQpzVqPk697917+GdCx
8HRzTBa/YcpCMxRIiD/WR/fzwNVTEFnvLPM9qJ4pJq9HxMrSu6H7AGoYupJNPoyN
rWiQWRKGJ+fyK8sM0ktrj1XR2of2WIyDBoP5rGEgIker9fLnWaOTgDnZxP43/YNB
Sv2GXhxNfxmlnOAgFW7wjH5ZE7BRCkS6jO2Mb61bVKbQXWgMHrPseVsdcybjJqji
FKJMrAtGEtuFAvSuzfTzp6utxyZr0g6zvnShw+uKW/lZwASz0wt3K1aRFzLz6rZH
1GkJET/7zrJ/pxWj0YhmAeJXGt+MGtrv6lB3dTBNUqC4t2XtOpn3lFEU8H/mmlL6
A7LlZMfL+b3ei4ILSp7H1rNeS12j7KHnITDfWiIxLO33vePMs3B282NGDyc6IHjn
KFmwRSS3C6SzIpq9ZUXRR+mp99V3ezZJYv1q/l3Eu7V4DBfAoIIQUPm0m4a2uWjm
xZFZqpoUXzQ8SzwaZnhZ9rgg8keV1x2Lu5y9ekDlPBmeoAatNaYXDQctkPh24RL5
OiY15qEYijK+wFJ2+ShOAQ==
`protect END_PROTECTED
