`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fp670sV499dKIb7aXNvCFeg0MQn8woZZXXeE6uh6uS/g+4Dcv+NYYDgw7F7Ujg/S
ueG+J8OQl6hvg9/QgCIrK/gu0/KYSLjjpXkBi9VuS6d7iFtmGmQ5joMK1ef6mctr
Gt5fu4XR/7Xgi8JIbQf4FDHG23MGorf63uTPtQFR2ZEZDcJs/iqMJ2l4BccHZT5c
4FPVNj+LbITMjBskndUKfcvAj2M/5J8ixrT/24WOCWebLcYA+NoJchU33GjnsOpt
Wr61xWDwUaC7s86ZS/OApKOSdmkqqZFHPlSz4NUxA/KRd+R7ueRnNhEOqFxvnt2I
ZGQ/3mA2uPfwpuixvu1ADjZGrt/OQ2P5AGV62/jfYASEw66kcDB8KETsz5oV38AM
p1VCCEQKo/NM3pi68pGzqR1cUeLJX51unhxYowRSk3ifrfSsri1T1Qri/XZzhUZd
5ccg9mXrPhGXbktdXnFk8XEqapzGtL88sUe1CXO6w8NqyWLgq5HaPypuhSqZqGgo
datJOCt+JTyau9Kfnaqke++8wg/SvoD9VJEfenLvrFdX9gDWjyS6viSo5VIK9ArK
ubX3IIUq/5lFkBcAGS1fzqbbgUZYqg8HC6p1Tw4YNeuOclPRfs0UaSwEv3Z00y1W
7qinfoq7si3KppvJCf3/VPmDeXNv+6ZYeN1TtLAQ9jnIHZIQPRp3WZijxhNQLyW4
cKtlRe1B8Ab3GjhuPBgN5AvCCaNxGsG1g3O1pKcwkDh1hEytfjAV5vgwaXmWAVPF
vC9EIfc/Y2dtgXnp3/palIl89Jnev0qIh7zO6NyoKNNbv2t20/EBiVm2NftWEkMc
g5RwOjcPMLPl8eRmoJRGMC1rnOdF8/YM5T8kUf2/vrlhzx7nlBIdZi0t5V60tIPw
Iq/17yl8bsKiX/rMqQccn75BA8kpAWxrOgnU3mroSGyt62ZLCgGbw0ecA3XZIFAL
mRwSyOGRgtzytgCSwYb/BVs2dZqne00TZxXKx+vXSl3ucbh2K32CRcvVdeO86g8o
xychra7FW+k2CHrwxQFYd2nsGJ8MjJE3F3mfvG+GCQAO6IKnuguJ3kNmuDjy61uX
DJQzOWFPvPbyhHVEByt34aMeSyFIeIydZFhvhV5wyAwo9bUe3x9Mm9onKfmHxyfS
0bAYqbCyWwXkgZgFcAdMUe2dWHGeYcXrM/yXVEJycVl4mQ/DcNjobiZU3scjiuJI
wA64TCnKsKRjOV/Ye7amtnlPXqHEgBIstBNSe8QUbFn0U4S2dehIqE0x6OMooISj
oOYjMnAs9rYyiAvQmcG60uc1T4hHNbCrwtdvIomqd856DwLblDTb6nMrqJTpLchz
D4Wp6AYBYoUcN53Rru1FW9JbZB18hoTxgKwsYH58yGPjnJj9cMRvshhQmEfbmH6I
`protect END_PROTECTED
