`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IoFCW8SImOk9GiCDo0OUsA7M9nTjEbvIBhEhlAT7e82cDk6TE7CEjeYURYo9Oo2A
ebsyLRUKT7e265n0q1cVD9SWXwOyVfpWrZsdgeLIuUxR+kTuDlfSvFmqZjTCnhJW
zCK46+/EPdy0Bzk6QNRQbsODbHGH7WfDptsSOccpKvLobUyvt7IpUaRHBKWja6l4
Gjsw2sSGBr1/hL4XKXS96oo12D2WvMRjK5Q3TIEihGuD/23bCTRZw+FVbNd6qZuP
vq+uYrjc5UNU5Gt0qMj0BD+syppLF7KH7BcYrQrzRAz4nmPBqqfgHfrUCgzAycnk
V3VVWNLvYGIpWdsb7vYOiB99Aaebr29YMh+HQ3cxv2JY3pExX8w2U4Baeq6G+2rB
Yyei4SdsCzOiexYlgjKYmI5j4FBDZJSO8kmwLrqo19PTDkwzGb8k435FHd4sZPkM
WWF2jjwi8mKeMtcphGA1uMJV8mfaiFCleNTRCDJ067twroYwEL1TIyNeeRM2lNlh
WJwHcgrNmT6pCqvQbzdDstyB11fMeVcnHHaaUYAM/5kqw5wt4zguuuDmpdSNRvil
6YEa/O+3tdUeUZUKgSxBMMmbNI6NHsUR5/e5ECVxfjfY7TxbCvtclwjzsfFlSCS3
S3+0e6Ovk/4L7KS40UOLrg==
`protect END_PROTECTED
