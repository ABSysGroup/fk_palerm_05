`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7tfpHyC2TvwgiKWjYTo6lz/yedenhbIS3PiX/7Fu39hzpNB48nm6WYlRNlmIyR3H
+m/W7AtnI1SRA+K0zDZWnPP7q0P5l+nyRCqZNiDwqbJ1CD0L1a+bT0BWuzgGu7pP
ZNBXn/skDFees5l0ilNP+dIVHPttZexOsKmqE0HhKiE/vdjKqCU2NqXmAx0qOuW9
+2rRjMgU6L0/FyIMzQB2sUKTkRtJZiLAKKsW6Tw0VX1IXS8Xhwcp5HMvTGN1FHZ0
Dr0BzCjo+30EeqVtdTSioaICEixXi6AG6PDzuYCevdZfWXOPcsvrcX95TRCK4z1K
Ud1fZ1Gz2YCpT8boemeiIjzObbylfvm28HVKz3XbklB0FBGzO04ZHrb5vcPwAMHX
I9fAtS5UQDCbkboDZMQhte03r8vQ4f063h8jatlikbDIDJcbGaejy0TjNjJGTPsr
lxkzcRo3Ji62rHuIe70trXVbBTSXINGjd4cKe80rLpc=
`protect END_PROTECTED
