`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4lGuw0KR44o9N+dbGgw858EF9jOupq/r6PjreWWf84UvSNtqLmruHZmCpqFM7f9A
0je9dxgjlCoSrUuqhw+yJsWESomz1h1HjRt5DPDfr9ymWAdO7lEA/HlVaHHgWuWe
7wirHAF6brk0CMShwuoSigoBc5uIex1L56bsyIGT4eUgHvKpQLTW0ApfLorMNstD
V04h0ADa1kYBYfmPHR7G243PfR9uM7ayG2C8FkiRCitUw5qaORhyM1l+SgI1zv1W
H0wCOSSFdDZwWH+IsNW14jChU09lncAA0LwCvhMioDo=
`protect END_PROTECTED
