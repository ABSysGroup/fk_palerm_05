`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PDGVItnKmHhabaDrSx5NU1352236cGkfLoscNLqmHrcI5qjP7GWLhykzE1Hdrd/C
DWY+CkcpQFeodyn1oei6mxlUYt9ye2wo6edlkXU8gKr7GurqgeHWNLKP/vMkYXm9
mBfsaqx9LwlZnHRgJYid4zUOZ1PMWp3LVE7iUgbM7khC7U/DFnrhMLgK6SMiJzJq
y5ZDOTu1B4efHdwcSGAR1ylQN7NqtkaSbn7memVu7WFUBd5hNc+cQlWEa2LrlfFJ
brKrZB64j91hgHQnNBrWeT/hR3UjWeb7OH3onjhuooaQEUOJZZCNnBgamgFz8bsi
qigDF6aX7pz8Jjn2CpaETVL7QgtEmbTCrQCiHLGbhwd0cetUJElG2gUFgIlPjw1G
ZOJibhOxw2j9UGlNivt0T+Zlia6fX1Wx9Yzgu9uQ1wIU4r6ZDV+s63ZuYBYEcAd1
/q8xJGvbcI5/mChq+7KWhGJ9ba5eykM7eghP6LAL6dSfNiwGXmFXsigVmF+1RAvy
Hc3la7wTMBh5Er1AIsVj9zj+q/mdd34uBK02xwXo1VVWOwPoFFXe9v9odVmnjS4H
ZggfNeX1YCQ4DrZZv+ZitcnkM9UVbC2LvZsMpr7kLoBXqePZXG0ndb7miE6PQqY3
g0Z5CQVoEB16E4xJI1bwUO2NLkyZfUOlWl4EauSyesOJDawIwwYQionBqB4kwtFD
WvP+EPWupeZJcXZsoQ5FjFPY9EyF0n7PbWvETc4elsa9TJZTycgKB0vBzMQIt9sa
rxE9ti8fnLS0Uhi8LGuAIQ==
`protect END_PROTECTED
