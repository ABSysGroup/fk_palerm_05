`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C4pqKwUjCY7pM2pP5l3FDt6+IR/cO9KBxKPpn1kh2kJ8ytIVnv82ssVerDa5OQIh
V25T+xZ9/u37L7MCD/esj+bu0PFRVg0ALRkewx5JY/JWNp1J4SCqRvTMeBbh6SzA
BX2h5hlyqVRM7WIHuhBTWdbzgcQhBi1zgKkAbkxOmy7+iOWHMBDJRqNxU/AFnKf4
zhToG1nP9Rz/Qqd1z1kaX3z9rbXoWhYr1p2h52LdlvKeCqrWa6ShXyRxnfl91tOW
bn6nz59BrRianADPvMpoZw==
`protect END_PROTECTED
