`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KyLZydVZfcnBsI+Qto7ZGAx1FL8fi74L+X0J2wJLZZNxUVnfjWvvyiVEhgFJFEmG
NuUU4OcGa9D2W2E8lHaLsJef321SuGa/C/Za6Mz+GJjhT57kwtp4Dq64Gcq3p9IT
yNdaroPJExSPJnKQc8yoa+X2ErF1JnosyLEkXJO0s/DcFr+vasKKCsmnpWZEg48w
onUne995coqGt8s+uNMFWrVzb5r1Wte4VfvLT+X58Hb5vvR9nT6Siv56T7KJW5Qu
QIccaW4b6EMPl2oVdy7+Dm5SzzAyy8NTdmCGl9GYuGn0DTy932SU0B6WqswhxLgA
dRHyzQbBH54HsYaqaAedYfeHgNuPblmWGZAQZ9numlgQiwFzaSMdaauQnU92oMzi
/E87lg69RZAu4v8Ykfvrh34RGLZt0i9fC6CwBxrLmn8=
`protect END_PROTECTED
