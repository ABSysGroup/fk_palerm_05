`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
53OxBs6JuYYdYolKeGKKyFLvRnGm+aEnp7SkHwxbI7lQJc9l61Z2S5ky+Mapw71O
JOYOz5o1fKeOwFrdbvYU2VEXGbaec0M0uNmwbiPVooBvde6zvx7et0jsoIEKGWnj
8qqKnfuEFj97EMSa1GJMXDDGDvegmz3tbiYWjO4/EzJFJQozdUTW9gKmqMKizvi4
k4UhC/+Dc2/sK/F2NnIT2JNHH1ezSiSQZiF0N9juyu/W6HV5O/izHiTV7RdOl2HH
+C48w0fEm7iU4gLoJT+kVoavpgmWj4R3imYi6G4umZcuIV9Cvoi1dpfph2jFI0sF
9ae5NgHPfNEstvuddPPQ6PbQoLEYiW/I+OPV1CZrXt6zccxrmegiU6tsGzUnHHjG
L6UI/ngxSxHPWeG0RyKuMCBBaM//UEtGnwshtF3EtzB2F5zg7+OO0dOjnQ0HGA9B
3QRsIVdw3tjoliIuShtqxw==
`protect END_PROTECTED
