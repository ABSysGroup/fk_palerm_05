`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/lOUYCU/eGFwQUgtZj/w1J6fBA03Orzi6hoaxsA7ZDXCP+YrZv3qlCt8LnmybrvK
szjqFmFQsgdC/Cyqr8vDoaVoGHBI7s7J3C3xxRu0ScWkIMP1useIq4kqmdyfaqgv
o7Ig2GdU1edTrq9keEmvfY77q3K2TwP9MjU4oRuAfwMKpl07nRghn6IrBfzKTux5
+wCVBu+7wb9zuGxLXTVyjppEKTYW9H73daF9k05Q0rC/3/lupWE9FZhquN2X/nvE
nfG7Vc+ZK2j5yuBJWr44DbrpbwCLvY2fhZ/MPk49KVG42H7RnI7av7zZ/mjQN40k
ATWD8jenE7BwTmPLwpWlyJ2pQKkCf5BaJKtj5iCGyfccrwYsL5cUozPMfAqm6sOI
3b6MGDfmRZ9yh9pjr15NvgKM8e+tbcfxLRd5kNHWHwC78aK6qsIwo1/x/h8UBlVN
vcGAuBJLAy5mDuMxIS+7F7XTpEcozGKFNNAX9Jwjgcp8X7MTvhs+LWGZdKL2Erin
UR8JBlyFLZbez0PhLr18EhM+jK8hBfqh877heVR1TqDrFJCkOS3hX9KeVPigsmlc
2scIk+bhfx0Zcxrujy8mpnmfLZSaLKBjJbJezeNTPB8=
`protect END_PROTECTED
