`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DzXgcnPHHepi7ykPc/Llo23OkXNqzyS7wGoewjkJILnIH2LnMSScaM6X5eIJ13an
jnfRHGLioBsgjK7YzvKC3ZqlYB8u75otYjBXHtBe9dWk9HrFH42kw+CWlawLxWt/
7cYjiWnJ+LkNqhzIlIemjLhZrwI/Wf42N8QvzJKfIGXiXr5Ai5jGGrs/kPKN6i+j
TrRPgYHGNS29vgCjF1nQr6yGanJ73GRonPEBMCYVZed42btGJA7mEPjy7Sw/ttBg
O6HLH18G6nSxYdq7TwSinhKBfIrWueFMzV6Zu3/NZCnmt2LV5VSJby5WdXn/BrpV
FbCuX7xIgVxHXbK1UKmZqlpnXIkgpRe+Qarn0jjV2r4JgR0QloQwjXkoAnmXbD+q
IgbB1uks/qjE6V5pkwC6vm4HTVNEr8rtnfGFCRVPBTfNWf766KWKPsVGPq735bmT
VvdDhlUnptGLTxLREST9M5gGg0AwStJBNHjE/xtkRJY=
`protect END_PROTECTED
