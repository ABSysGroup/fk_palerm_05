`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hrejUcMryq/3cw1uCcWMxS/P27S+4PDu4+O6/+2BKolowJYqSRENEaUf7DmY+Wq8
Bu7JClX1ivFuW+qCKZSa8RU5kXwWX7ByWwD84btUGfJh/8gOV3Y14m7W1gxJ9/bV
B5uTtJV3YPQWBD63oMm5j2F0yho7xXnGJ7uG6opVhJjQxh6f3383dDlSI4INyRCl
tuo4eEhEeMRX3BlBQ7PXumRV66paynbPcGsTN+1nIGCpsYEJv8/+QlvOE1sTawlX
9Yh+O0878dne5snPrqMy0tjTOF3ZPT9+rH+4ynBXM/U1Lukvn6BfYe/s7nRE8L/+
sXcmsfWbqRg1YEA7UTOiRDUklyhd8IkFPLMJy1RlO2A=
`protect END_PROTECTED
