`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ms7w7RKaP+6o2xDzbzkLjTp0ZfR9zzCxC5CgVUO73Li+2wdua50rJ26LEKpc3/Tg
AURta90Q6WfE622MdW7HvLunowMZqlycSSmxr5UOzhgjbOrGZzoL/LWREes16krE
CZmrGtq/SHmcGda8Gdk71uMvZ7d94QofEP8LQe+wjJP17aUx0BoztvRDS2FkwvqR
WI6QZ8fyzSBlqbLWVimtXeI9THiTodP3inQ0PGgQznoAlqbDcjB7402N2bPPlS0E
W7/mCTNLTG/V8bfaNjRgqcQXGy5e7cEKNv9spfycMyWXMUaEbx1n0db8PpKOnxZf
TsaDssR3ZGbw17HfeA26IQ==
`protect END_PROTECTED
