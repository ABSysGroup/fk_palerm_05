`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EvPi+znkqCV1z8XT8hL8kT/j3zMjl2EgBg6u+PjZq+zaNyLJnG8mYlUirVY1cDtJ
PrBvrK3ngTPrSKnvfgPpxOsdEB4OxFgn91OE1ofxsKXrK6qCpb9Lh52AIX74Gsdt
juYy/Gb0T3DrB/DszvUTMnJqZfCtedLcXc1Q4BA9Wchr9c+Q0IE03cYeiapOcVBz
dTyVP+4Xl4MJAo1LJt5MBnbdncbU8rg/465iVmTzQ33T4c0vK8WDV30ZUPdkj2yy
zFU+Usd/+ll5M7ty/Jztl3agu/lqxxajTGrARjCFSK2siNFPgTdV0C1MC3QccBQS
SqXNXtyqa1dc3UNY8wusNFZftvvaQ7WJ5E3nXWf5/Nj3TlWNAwkRj1tJmbO5qzAp
uWUdC/rwX21jq167e21d77Hz5c3k2vEzPDtmw0df9X/cprT65N2R/WDa5a4zT1VN
Vf3oZrX1ialgVAYqedBfrs2n2LxshgtMv7OTzVzSskSYY01U+6g8Kw4tzyhCcs6Y
xO3JrNHE5u2HiIK6B9GlSZLoD8OOMulE8omUD3EAnkzSKxhd9wCC9+3fkanmJSew
TP9vNEPeVsO/rnFv7noDrqG/16vG1RKCw2H4m4CZUDW7fLsH0UxdtkDyKknXIFDv
Ld+IYInz85SVsL0nDDm5GcM2ClKbhy+TrMKG6jJXhvT1QlRcwpoREw/wf2m1nfMz
0C/LDevP1hJga5BVgHbdoig0yEHgextj0LbykTY/4kvebJQdLitViBoKFfciaypD
ACZvIPn0e3Hft1nt2EYgluwkUFJWJEaJwL+z+cj3DtKOvRPFnL5T0HIFfBuDarXW
9aqiLQqvNtpnphpE74vrBtxY5Z89S1n3WcqlV3HLmJ1aVMyTX6ZuFayJlCOH7zqd
4HkUItDFEDS4SwZRAw7zW4xYneGVE160A4yJiG1kNcKBYQeMMkpiaDS01ox0vxax
GwgCmu3osaOjiKWhCftd5s8t7y7rfEwFZQy+gZfi2+7swlmnpM0sOJ4ZB+P/WvBh
SHajBEgjUAVGUXMn4GyQFHYdZOqtR6VUT222DSLfbhdlrcCvfz87EpCGGeu694vN
JXcQZpBxYpP71GYiaspHvQQ4ixdgl2OhM2HMD0J+oTU5CGV81vUkW0u1yN2SHkuW
69H9ablzr6xPOEeSLMYakG7TOkv7YKi8dvkTU1A/3rDhRiCs2N7vRu6Nb3/kdZeZ
IY4OeD5M2/sUQMaL+BQGKyB1CxV2CgGA/P3dGCV6MK3GTfby03squPWuDEkQ4mmo
wU5HJls/rAb+C9lmcWMz28CuqJKxpDZKEPrFXWWQV9DZPai6Zo2QGkKxiJjFXixY
iGmThzR+Zv7bffPuaN952TaI/6ed1l8piJNTRxhbpTx6074qv0vHLvNpR9WPinmw
VZBFNzJTmy+Oa6w25sFJ/4ACuuqDuYyWA1wiuhzUsHG6/DoWiWfrfRKs28CzSBOe
A9uKfa9tLC79loWqtGuhfE3lKPHvOpaPrk6a9eYv2AauZoS48arIMfBZd8BIQ0yK
Q6hdnq065gLK1ZfiMBZfJJPdGzee+xA56/40l5TFQRd15E0iBHeeoVa5DE8p5zse
DjIYCGjCV/AV3TjgN3c18gj/R0k7CcM1WDY7mKvkJ16lnzU9VARMAgVaELZv1ooJ
PQuEWT3hmMIknR7caHRnFCcZPiG9qP/Cbog6ygfP3xItJZ/bZYlbQsL16JvA3eKJ
cTQZ19SB3LOBiUjmTw5x8qGOyLuXCTYon8xaqGqYg8PfdTEvkJmspNzA+uj84fb/
MDGR1Ep5HoBs4VWZE5GIf+qr6V6eAFjjrMuk8G/NBDroDMX5f7KcDg5jL79AqoY8
YsQEoJCTJFhNQz2FYN0C3qAa1apYqXXWCBBH1vONARSfm9noSWteTq2UX+/dYoI1
+M+KqrRuaFXexlPGq27dTgyBHq1Q2XrUf/lzrTlQCDAwek9C2KWq5tI5Du0e9pqt
+bIEMUR7stvj+k2P3P4WoZ9GkI+m+umDdmmp+YNhbRC3CgD3d2tgZCfdFP28PTUI
VvYsbXbqBPmVAu3PzX88DPqZOH9UPw1rnhPMtHEnl9AtZOjldv3uKxnu9chJB9zC
1b8Wc+jY7iFwMTDyBfaHb4MDrLqCjPf9XlRmsnsbah0xRyUJXMHmoQ28vq22cyNs
zRfc0mIvDm/CS97//33JIzPLs7LFYzaEMdWOvAfgcijEGhlcZZMBXJP7/CUy82+6
TNzvXhPuTUYpGinO2LXhmA4IORH0UY0h1N6mH3aqPZTddABi/k33O6vGkTtcOePt
gh1S08V50aZS7tnN4X1FNP20WxFlcODzeu6q2pxfXbE9eMqvsWhznFvbSSuy1PLO
7D62Cd9mmSGRd85obRwzHpqSupgcF5cb5X2SGPd9MHbi0bhpwoPVugBN3X/WcCCm
cXmgyw729tVLdFo7kDvhgNoLF/eN3rCCRnBxPCpe0OCMGMXVnan9U1POQdzTJL+8
0VzGoduWWMFWKKmsRYVFbxXgtLdutib8y6JUixKVyKf6Tthazf6DLtg7I1MekXpW
493hPvpmq59xsuX6RPncWw5EhJTKdk3Jl/Udzxb7t4f4gYCDOzULimNDQeKwqiLh
18FaWoo65Gl4kfVvaAaDrL3UUJFt1K3OXUNEKvuL4OMkpyiXq28MpDakhNn93K2r
vtwSVIwxXFydji7Pe6f8uzg0eyCKUtsXZkeRWaaaBDEVfdr4u/tOKCyQmjBu8TEp
DYyoDd8+JX6A3ri90EBvM3GcaPcy9vWCQmzpUIwqy1aPJn/7xnbWfrxuHFD1444g
cxsmF8fTbKs2kWR8nTdf7Lt+MZz3DYnAyan3nsKEq2TnECFPFRtaiwkg8WNiP34G
R9mVDRupOGDfuLmNT1MsvzEvX6P5AcUoMgHnqKVAHgppUuNFpFkrWNYyTwFqo1um
CCzL4+DV8fzbl7tBFW6Mb4KjUzXkl/fTsm2Jiwakuy9lSKBnaQdlct07UB28uT//
xqHYQugPFcVzBCjQ4ecreH9Rib0mtLY+qHTrNsAqQNl4ya4ey5rQMZnXSle+OfZ8
fx3EO4xi507Pfw3GLeVqLdxa3C5xDOXEDqnftMA8WRwxrjMiKmSTgJtRwduoJvKc
Oa656lt+23oCnqSfQkSiaMfe0VCPbfxeiRsfA0qfQD2bqv9nl3whUNh4pkjPS3c2
QkdGiyb6MTJSOOifox7g52Vm/OcRo1/XoUcGUptOwS9Zbw81ie7u7HKG8jhs2kfS
PmyOhntkCSMgy6D9Atn0aXuiMB4/j9R2WTFl58w4ubLNVY7LaQ2Eqzmhw9bp+ahH
862p03JaiUE9GHKRDchkT6fMY0fNCjxYuy20etFQkpirGDr9lRrK5US2ATtLAdmX
GuSixjVT1hNelqv7Xho5m/dv7S7FDAZdvU3+84edz3R191op5svW7WEkHlzxz0at
wclqSKo5W10Pv7ChIkEKVaiuF+bUxmq9UA2vmcCGhKEG7hxcZIYGQgMNzoZSqPxO
KlrVnTcWUK9/OHaaEoNrOvH5hKyikVQYgxgpdyWUG3ztByjt9IculYKF/ibs/Lss
YmwaEt+hDua/cMqhVVDt/U4fBT89N5EJ1VF4n6PuFfA+YyCOjcskHeUUmijf/s7V
1JL/PDTN4H10aYv8wiILRZdKi9JILyW32DENZMH+OsPhhIct1pO6W7wr5pFBCLOq
e9ReGaB0QKhxQbMpT9h4NrzldTI0ZGjJuL+1t+VdqO9ec0CMn4aGWj13Z8afaew/
LTiKSIZG864LwqSwoO3wY1PUg1h3tUj/f+3D68muNSK+4RMqQw6ebYkcL8woOZ8e
iM5ZcabJlQS0B2wi8MFJbWyF0cKo+TAXRHejTbOabP7LgenTbdXPwtQTutpIVHaZ
DseiE2kBt3PzigdSWL3f12H6rHVHMOt3qQdlI4CdMzXFbqyTrnZsdy7dIkwOiIzg
5cxeMf23a+Lr3qltI0sdKKxdhUIIjdNxIguqtgQYAyjCgHYU7FkcRz3OB0ZE+4wl
8cFfEv4CGiqrTYo9s2hYmuIzZTmV3U+5V6X48Qy4mg92Kq+Z2gbObkU8/7VYIjSz
PcxleOrdWaVDp0dlSMtF9xvH8hjhQLkjlGfAw0J26pa+Bb7/AxC7qQ/nydrPehoR
EQE58AmJ/mxJAL8qJ9k5B1yMabLZnPJPokAJncPogXXr1O8CmvpLhbnOugzA4zzV
wnWgW7yWn9venaNFud5itCMMj3SDpoOLXcZMVgmAZP8J494cbl6zM2I3/kfY/GB1
KZDoh0ToZz12bOQ+bljSVHP2lj7BlFfaMshss6njQTzcMiM5AcE2q0QDmRL0zeot
9+1ngM8ipvL19cUZSvmXW478OFM80/gnb29n5rTnoP2+izwc8+m+Yu3938lVhv+B
Za7x8Mk3KmWCUyQ3pPs/Bdvt5/3EulU+xFZOMb2rRVHxc6yN2hpLTe+RIuLBQZ8C
76TOP3sfpnvvXkiOL96ZmXrjvcs7tzRVx1SRrxa8pDVE2WNNNoxXwe6KhvlfKHDr
8RXOZL5FpByFUqgPFzG6PU2t32Fx7datOBqQpV4JzJNL9feIVEUQPWFWJud+5ftK
JayGztRKjAWeGbbdNx0DFzPCYBP2SXfivLhzTA9zDwkAQMwo+oS8+orhdMlorZ2W
HLsYf0j7nyajqlo9Fmr+N7w3MymEB6N+a17iuybiWdEucFcS1+giFucRJKbsVNk0
oXfBnKVjNSU/Fnfh164tkHxVa2q2YUnljmzsgWYoGLmxKrdfSnKhaGEoYcqD3gO4
ofh6y/rt/+j2DNEynKwUbwOEU4hY0S4pkqkAhZsZAcbJYdj6USncYSbVbg8TJlx7
bouMF6CCROpd1yPwprx9DHbfcn4GiwFj6RnToDVMmfUh5vpIxjMZCpnIRUHs+f+3
zja9+MXQQXcZ7TktmPZYgcuuVtrLVkCq9Ij0g3JlLac1jlrRzwREv6FOVFL316y7
oVv0WoZ/4yCe94raie5fW91GRl0/YMi4oXUTepU0OOBpCYBKi4JKzyWZCNCQrgZp
1eyWIUtVfXp7jBjMjz2Ss45xyf4AxF+10OMopkhyiFyyJ4jp526k0uHN4X03qbWA
SIJ8CWDDGPvC4uLOPOSvWBVKjIZaT7+Mrelt2QNuRjHZ5VnoIfVEL76y8hGuZvMK
FMYV8Cz3LTcsxph1s+s2nHDRY2VYrNSYU36s6geFLS2EZ9295JXhfxg2pTvADnOw
eNqK0wM5F0c4HUyKdVhkP/8CP4/uZCKa7u3vqnr+fWLJP36SRlEO+4Zt445scDxB
rPwA1gJMo3ULm5N4fJa2hpeAF0OqyeP8HgYGtANHSvhq9X+geyZSgDc8QhFE0w6V
h/qTZ5h60gy2RWktOcW9UVmCHkmMN8SqP7OJfRezJhqqMfiu9oNtvD+wNrOFCVq0
QdLdp2aLmXU8+XKXYeELWv+SmwnjmS0cvQfbIW4OR51Vrt2cCsW64dHGdB/W461S
ANk43xVZ7CbYd5ZcJV8n6KewOu/Kb5YLFs8DoVzYOXuGoR8qsyWzpitGQghHGihP
IFZBDhTyKsZvCdAb+2eKGwrADLA7Xb5wU1ddMyiWWJEL8CXMOX4mJK0jHC6p0S76
Ih9OVDK+hkpu5CFiE9YrFcZOjYTSL60whSRNx0WEuGV1a57LCBxvjuVLAZVk9mql
7V8LnwLQ2Q4XsU3CBbiJtYwRIOUuTDB7wKLAJTExttLrrhr9EZnlr1znZG8+QeVb
JexjhT0/BXsFjPx2KlsAajG7sqJsBMhNaOpFMPU/oQe/cBi9vReEEgAnm5VPtcXv
DbrwhU5BKm5KxIpvHxa7eRFUIRs+TrgLkH4v8PlxuyHWp9MywPbjfi2W/tZXmAk0
wBPbMIvNShV9mxLRpJbpONPq6iU3IpfPV/0N5DKbUNPJB9CHHigDGy/B6Q3lQbBt
xbqMNqTXHlbK0W6gU5oHKziXFZOtVSRgxMYO/c00chlIxL4MclOUhtjcoT6VphXI
UGFs00iL8loy0fxywBVE2rWSwumS0JUBm3Fzh4fe+aiNOowWLlTaAa5D+BxXAZKR
M42rHq7mVMSiJMrqmZAsBE8oAt2ANiarRvsA8UoJAQzaKbvm1qiV0Y1u9dfRUINI
FPBMT9jRSaOxuCVw1qOFBI+41qf/yyygSqdif/MW1xmti/X8ViFz9ZLHOg4nVq40
7peTp6YIkBmFkdTHktRFPWlMjAOON6aGfNCTKtG5LNtKB8tZeviARo/kIRqd0j07
AxZZqAUHJ5vyLGxe4vs2n968qC+WcTcu9GZPsqMkHBGH7tnOjxUJFViicDI/G/9Y
5UqVG1vIns3ip8UA9IT9XlQGukJKn/qPp2dhN8jk1lbz66Sg2YqbMWvt1ISTNrc4
D1x/A/ddlF7NweZejtRfMNavm4wRpCl7RSfmnTEakfGPo4aeguPOxTPZYnPCG71k
HtL+3O3769OK0BcYJHc68B1YueAyMhNlMazzSG7QsqgnFFyMgKWrWfe/PWuS+RNq
6Dzqlk+lOJFQ+k1Q8uUIEl1xv1mWwHHTbpqCKhFA8plIDsTPj6I5egy6lxgTmZKT
2vvMF03qK4adQvsy7VbpR/yGwtieLsA+StvNYi/zVvz5Rau26XZubrNH+DimdcM9
HnhcPgWr/AVbubPppIC1xcE+IQBBcnifM3J0of4NGVPNOnXltsQR15jwcUtEtIk8
Tjd2XPeTG1CJhXOcEVu1w7qv28dfl9tPqkbmZH4PD9xjPgR/FGJvAXwa6OFXzJCm
NjfAO7PcYbYAGC7kWLcgVuMib76Pbo6UxNyA5PeGKSuQ4oBdd5Yz3sK73SiiGGbf
XykU8MeI/Fh1hM2j/PHyKQ9xeyBgHtubj/AU+2NIBRFWDSRxFpxv80sBxwJgXeTE
zs0VI85TV9+LRVXRoCkiqCXQ3IsObjBWfLP6yXs+SZMxzMdwTJX1/EPJNuSmNbKG
vYMW9Bu/YwlQXzQvIor1d7UvxP8ABkji6OxsY6v/QlOi8qJ2WkObMkkdWUIQ78EG
q6XOgTZISH6H76LfzP6PTf+0ioWnpu3405BrwS4XJwAhfqKRgY8hLUlmciEJe/Cx
abwybcS39cX8wma1nDhFmEkFrPn5/kBAqy84nQ1ZWdnOo3WkCGGFp9F5fbDcrTvO
jYE7vnau1W30Uwa//pCqfj/ZvJbtM0TifeVdXiYAw/dW/7fvg0d6/62lzwf0u2Zq
+W5ZSH8TESw0zWz6myrdZJBGuK8VkX2oeJ8+aNdw5xxixmBG78jlo6+1n5g+ys0Z
Fuu86F2PLwughxu1xKT4P6ui/dyaspyya7VQsqftVqlCJlVoIw6daMMij0ciCwSD
q9C21R3BRpVnAbO+e37w06G12OH+s+eY4LSdmZBr9pkaVqvhSadUvnmLc52kW1pd
9HzQdidq/GOxtadnK6XpszaH/XLG0vLJHMIZTY0Yu5RXKhkJgTKLBLycBLcHFfKM
rDUCpQ7amFleppb5ykMeDKAcawBIe3MWIAACTopwDRR9Bbtsj4Fs2ywbSwfkjFvA
pybfPh75yHu5wq5KgnSOObnSLtchN1eny///eIqWnYVY70VbkpZ569x4F1atLz3J
V8l9k49TIYVjxkHV7N4OZHUUb1y0B7uf+AiDMHnLGsFKXubyHYrVoeMlCYkjUc5J
GXNXHF12hcb5ZlgMr9yMKmyEnNuhm6/lfxmcGOlh2zdGhMwHWnMhTgm3nKpforDB
qfvxxPRIXZ7s1hxjMukD/+eKy05T8c+WGZbZw2kaxvlyXr60AcrThpqm1zb5Z2np
z362r6p9mOh5mLAFvu93GvKzF9tCbEHQ+/B059muwBxu129bm2b8AfyaYnC89yfn
6qQRfkH1fWKmcg/QCT4hdNTy+th7REwd4uwhTo0rLsqpX9jJwRbN0FoBXc3WB9ku
fmtjJEVVyzAikbpTKoKh6cQuo/hM++NELHC00CT6JSgevipvzikbBq8C6iKzzi6f
UDfUX30fSGOeeepUb0hMIyV3VSaNs+3QHI6FPh2NyqVYqGb7viIFzbQbhaSyHkLJ
xviaEWldfvEhP2w00GHgz0GDLENLNMoRdMyf6dgdw/q8MNBddLO9Q75G/rWBqxyK
HMgZAm+cyfj4n6RhGm0tfR7g8AiyZCuPfNM49ouAL0yVpIrGDa7hpyiNuvxhku1t
i2FslsqGDcZX8+9nufeOd5UdwJV6kZse8mAKAAU4BXBCuGt/3pI+NiZt7C/BaEU+
+pnVSOBg4RtUpIy3SLkiW6/P04lnMaeLhMhSurerRzP8SBRX37b58ig58G9Wxcta
KgQAv8t1jEvNtsSJjQq4TlqTSpXINarWNmeNRY5dJC+a0Xl5DgYLp/9VZHOzd89G
g6JwM14/cOY7TsJT0aoxn3pnt8ZbwlsaX7V/eB21gyGzoIjZhjjCddstpb5ke02r
f3NJt+sXLwGvlPzrbxEu+uW0NI5NQ99gets2z4KLbIB8cmqaYmfWXbe6IhHemKQ9
nrEms1IDXecg/P1+1zTovWoZfbdmsiGr8syb8cBhfFnReqV5gLekKstgK1NiOSNP
CfLSO2ohL9X4tCak4lsjy6b3tBkO37XKnfJV9ERLXL97C1yzzbaj2Hrpqy+bFk5s
b7N/HoRJxXtoFjVg25vk87mb+SRjjmtttnop50Ctvo0ZwdvxD+7RIv1PtC1nLhX0
s9+T9kXG0f8NCyQZWNAPt9/uz64J/1sHqSuOt5yP7MXgoGjnbNPdkmzOpw7nX7R3
D8JYMRTjk6wiw7B3T6quWUEc0Xc1avRFn6DkaT8WbSYnq+a2BZjGjchC/pxSstzl
jFRJLWZIcu2vnvoLePHsfmhd+TCLiw07inX2DzIEQnLRXs96K7i2jfh61yG1mHHr
tcBgxv3f9yF+00GdgXa9/m4KG412vjZAaNPAUhkftDdFVrFJjI0/eBJZBFSyeBnx
nka64XRDev0JpClfaY6J/5ohZbAs/L4RaqWh2piqWJXrVdBoIqonLb4tTX8qR/Pf
I/Zrb03O5dTLSh6XlyLIATKLtKW+kMbv1yiGUDDtuscqLMgT01ZQa5NpPefzp3aO
1DnjzYtzcqn7Bl57wAt8a7OMnYUn8Dh3V23rBPucs/6JMwrvGIzsfdLTxfviIlWs
v7jCqYEF+3lq9KrSf6m4ev8w+GHyaG6jgl2mccfuaBHQWcAw5F5StSG4lcncxDbM
AQrE6U8lRlNoqROPpDhCbPA2Dwf5kax6MjIFHh5HtM4HW0k6hATYgPt8neZxT7F6
SYjY7xa648gtxdEGR1ztXGWOOUeNeGKQ6hWrUSZ/jLmg1fPIsO9qta69vYEKPn26
lJ80cZRFWIJxq0M6AqY8z9hxRQL66i5EggluGdymTwX/UjTqsMcBlZY9OS7TbO21
Jkskuy6VVBTNEv8wAgJgPgcI2GxZ2U84TNg6z7yjEUPCvQ64E1IUWZt1/AhZiUYq
DEFCi4pOaJqfBnLGYr+FJg==
`protect END_PROTECTED
