`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Co5HeOUtiIBMpExYXmsQr0Ydtu/f4fFh/N/XN00mkiYTiRSdE0Er8E+of4DD6RZ6
53Sck3VFJCRdvzV4IvWxEWPZn7JX9KTFmDG39kABla8YV+iJgvTuGEyBDoI3IyJU
wdEXSoDCyxgT9vzGfyiXUbXlH46RhSS6wpR5Um5ZFUeT0m/DjJoTsHySYSIyyPUA
RatoLRjZ9/sCQRHTVbF7Tn/1wXrwRxBXAQCUXVHTYB5RDqrZNSSL8i8Ou8fpKYMN
OCvgJ2AeME+cF5RuF2PCo7OBWljt4WSGfXSNNuEGj8JqPofNYXL9nmxFU6ji51TJ
bFDMfhtMZQ7ixRfD2T0LYeF/Uan1Kle/087yNY/14UuFhYGSl6sokGJOuCuaeAuD
JxvkC97Z+tZvavMdUPZSulO2/Zh/PEO9A8TYBn+3nRULt+/+07LX//u9wPq2fokA
uic7tU8JDIiLXAMKSuSxurVkPHrfEX8MhgCyAEFmpNRtof3JMj5fai5DaMfRzAqs
vHIMfTNcrrH36QzVjGgfHd6taPqozmOYwVQS6sHjsltjNs2mxr41QugQcQFUkKKZ
sy6rfzFA/u+LS1KkEN91w144EyJYmpNPmuL1xtKRxrVRyRmr+7TpQoyEo25LwNBd
/IeMZhXTJMEzap0Qo0pMDQ==
`protect END_PROTECTED
