`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oLFygTHDrTSzXKxNqiaJv/1zgJzNj4ZwikORUiWUsLyPYcEWUwXJYuJJkw2PNCl3
CNvEiBsPBOy0Hl5my7cnEAmP5V5McE3cFVyi7PRlyKidi4Y//ojzzjDIm8oglyLy
ZQTxEVRX14EvT4xyTaQm5wrRzNORJ7xn9Szhx9t6Oy6TskTNK22EbXnHDhO1v0qI
L0iARapK+9gWU5FyxCZkOJEJQX71iAJJGw3/iiuqF68kTgBsEEj04Ph1gJYKL1Q8
S7v0gdzy2eTDrxSOU6FiOA+Hv4s0YoQN57M/V6nFJiTjLbodAuOdBkFxng/ZQJaO
+iYrZNGlrT79J+SH55pSp8pO1w4FTfeJljtdT2mmCPLsgl/bgN1/njpL9v495d4S
tG/RlGPHAU/I6Pg0ueqOKw==
`protect END_PROTECTED
