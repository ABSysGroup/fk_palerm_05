`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qDUXMNlqjKDBzgKvHvs2PF58Ljraowt+4vIT4KlOuh4mp5qbYEi3cJuEaC2hAX4H
e7JxFZcxE4Ii2u5jkugxAwDcZDgospNyTKCdOu3jqHyGqIkNWapgOdmi/y9S8frz
5DAs3pKKlN1ZOr2ogKiatQZff4nTKVTKVyD0XhjfmPowdGjQNL0uMAIavtoHShpP
QmErBSyzAVQr1CF5sCiJZXJxADg/5yLYHKxpIOMGme9pB9hF30sGTYFG1kUbfdYr
iVupf3IZzn6AwRysdc/I+Xq7BXhd/HM0rrVcoRG3Kvp2MnLSML8bYYUeuMVsaIOu
h873oJO2nd/A5KtV4UW+1/MXJl4AvqBjCc7w3rCPQ1GV7bbqixr7ykeL/86MUxY/
lLjKo5HAPoVI2tvh+T85k77blq12jMM82/cR6H8uts3JuY3mrx8LLEYz9BzUMRkU
fGefZLdkIh2BMr6Q39s1B06ZAUNVAoMwo3bXkXgzkaiuJ91NieLBujfL7j2yKU+e
MzEDIt+IbDUUrUD7uGNr3Iml3C6pDWZcB9p5+92uQ4g=
`protect END_PROTECTED
