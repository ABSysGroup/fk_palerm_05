`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hZZUwoCkXUmjaEgBJAaRrLIsiIb43EVZqzNdszIRQN3IvTvMhBWnCkBg3FWQM2gE
zV413M5mOjmQg3sJQ7XB35q5Y1pG22k2QITP8HcelZKqyeakDUaxsrCfOUhsmZ3H
IcVwAmvnYjKdT+K0CzZY6Z04YuAYIZ4tjmPDjZehYCBymqvDHZxVR2yLrVSgwpCL
E3NIYH5puzuSTiF1Lq68EVIiN6P0ihP2KBbnaIlogHkZE13zLqeN6IDpQa7gLrbg
1lNqCTASiEQeP5zcSG5h3eOyk+6ycZ0zSZrNvUM28I4ZKL704C66U+vVgqixnboY
FYCYw+ChQNz4THP5KF9eKQaBpMG5OZUBKkQ0/ER9NjXNkiNhp6HGihAVCou1DkTE
Kj0Nkt4INXc+WEUvmEYZaoEWI12UXazCaQMrBXX/f929CX+94NbSce56k+J+ywNv
7NYDvO/i3XvWqkAPv4ZCL18vmn86z25gymk9NbbE3CDfd3ugfIUT8UysKe2upmLg
YhoLczqzoAzYQ1yNJwxP5Enn6rgP5bTOXdKPXYsY2XT3hf5porbjiAkKZsEaRgRv
qwkjhANXe6YFkxTQC2AX2Aac5RzvNN3RrL5DKNaKcYuiQGA5a+tcfgZPPxiVbJ1k
0CifzB7UQu2GZVlSafWw+rPeyD71YMH6VV+9LDOSx1V/KCDpILr41CXMjW3tS1S5
O0If5Y3KmOBK/visnNMyNbrkvpKlagslIvvL88wX3c8wNKPGnJMskx+as2On+NSh
J9palduQYo559wJdCgX81A==
`protect END_PROTECTED
