`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j9/jrRH+VCCqjhQpka5YYAxT7ww0V97GbQVbxYvk0W+zXXubIUE8BS0Cn5mqm3Ap
oTaLEMFtYSNP6PWPFB6IBI+2ICKnfnKCTI659JOFcn1dRkSpscmsJs8evVrZzS94
YupzuSvSUJwFbkvLbne2MgGeer/UuCBYCOJE88oVgGbP3G9FQHkPYKdCv1TZnfzf
vjmx3T3R+biI1UG0dE1xWWRtjFzwbFD0XbLqoQzpeAPQtIv27rMREasXjXHw01Ie
8gdwT2Puc+8TkAW2IA+soTldmlhHur/l+WsvumyZFSHyfCG9eGY0YlR7A5HB+HCj
TEE4jGipBY3MvK7LbN1FnSEFf4BS68yk0sjcAUMYNVRJfCmYcK7tD7ufAC/JZ6Hh
nnEY8ukc/RoSp2WbXedXoevNZcxFpzBpa4reOfJ4hOqCdlQoIj8p3jz5dijltqZp
0hOFqE433/kzoAQM9WrQrlxQhVOSy/4b8Y6ksui6M8afchfATRMGRMDjj6R6xPr5
kP54JAmcivFCJLv0wkVvdEAzDyPzyOIpOMum7T9LNG4HALvtnjd/7TvyRgSy1fk8
NcXGSMbsDv1CBj/YcNlKNdALyq85sn8TklrAqTLtjBPVVfn07NnuTWIvFXQy2jfp
kACaY1Jm7ntWfOetxaDYurTK9LeFpK2wpF7kKVDGGLv7+JDTq2uyoV8j2nJ8BBSu
0B2wmtU1d/U3XxIWo2xIJbWLH8Y0HH+IhgT+ie6FGnvow3w+w6UjEjdyhuKnfQNs
Sv1PGjVSi7mugo3q9yzIGpNsx8vE+aIQs0ZUhmnuBMb7d3S55NvyeCi/ciknvNdH
hn+fh2Bfez+WQMJWIQnBF1CMt4EwaX6826+WkXD8X6+GtBq05u/658K7yLUSao7O
rVcrKZ/tlfPTWCbv1ccm6w65L43mL7tPNbbDRUMdhuuaEpYrTqoKfT1gtgh1B5MS
3PT16I+Ex8cxBYbOjHNPv/9JZ0ITBOtSQrdQEF77KaCjdZvOFEdWvG5w9hjOeVPd
qvDq1PApHWpyMjQsm9wAqeW4jWTbr7WeUz/67z99HVvbBkZsTDVdxdaAObX3ysZN
yNmyeJgzgbddv5NACj7Zm5x1b+YHz/vLPwTd5ZaQyGGe3brrW6Otlsyr1rqAhchR
YX9sc1+M59ROhjTTl1wqLbXpg0d3KjA0O4sLeucbxs1PTj+TuaUEtW1Pe6Agie9I
w1KcQB93cQx58wwdUpIsayPwivmbPDDau7cm622nQs9d4gAwQQMQqkZF/pNdjZVq
GUYlGRSOGicoxoiIcTfP2DWu8lHJSFBcQof+Ov80Zd+VGY7KCfSKdHBmkAMvciHA
s1LngQbFALgeLMKmlEDkQp1vZ/onXpt3kBnEgurXPk0AA3MkAP9VjbGM9seFZlES
q3/2cVwDeaDkRPRHFZWc1g==
`protect END_PROTECTED
