`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/d9QzEel3hRL+fgJTLjSDRqf0vEM40KaQgwAmSXz85HMP+1tdIPHfnrmnY4WqLjh
CK6I7RDHQZhclVybdc//7avKlQStiZ9+tQg3SO14c4t9t396NamVkzR6GQwOToTU
GoKaeSw4BDuApbDJ81iWO+05zzft6WQepC8W0XjRpO+jD768dfvWAOiloExV2BDT
21qsgzUg517CQgvEMgn+AzHIlmab3ybuZWEuv/9rGL2uW4qG71fDmJLqRTAtii6w
U4ilNowBrd6FaCaoqcsJJ6qTBgYLI7MFME6j5yk7ZGmkaBsrsxN1bSbKC5PFEGy7
2ZaQczkCQVHg11Ygis/RBCTmNJpOSejdx0lcIUgpsqyWsG5VgHjFLSttcYTHmPtA
ruZVYKgYpMVwSz382uwsc9piQRFN2JVfhUaGCrIlZU37aOBBH1bjvp/lUhFrRQrn
six8uZIlelcDq/v/2v4KqdxOGxbyi0Sc4hZY9iLvpPVIui6de2h09Dqsy+PmjAgT
n0/3VAN2m1TIDVFndSE0EjLL5kVJMHfHPQfarQYWmdUuD8xWDSIiMP7yJHTjZxak
r5/d6VeaxjFyc0MVQ5/QXqWtYanWP4kwMJN8ICnJKksvucmlb+UkWrDZ9/Ko9iD5
lXiYmDnF6zAZX43+SJu+kVbitKEc52/+CXV1yMwB26mXF2lRk3pQf+yTUWCgS97Y
`protect END_PROTECTED
