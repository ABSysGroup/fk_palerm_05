`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h+XIV4Y3ZhFr4XqWSrNwIAu+rG162VuBtjdJFyNSPoJ/D53gAX3ammdCFPLjq0Ub
6s30Y5GO5BF3GekaAg9xO/3IP1BMIrsMa4UB/GNceCXLYIcTj6iXGXOr4cVn9Btb
7v4x5L51wENHVGwRlBrL4QDDwGv4D+twwPZ4OsxTwXWT/HfGKF5PXrynmamCB0UA
FbxYb/EVXGTOKirdA3hSwLDW+bMiSuHk5Z//DnTBM/j+04qH9sezi3IPFtmDMEGi
YlYm3+ArhHAZqUWJs8FHLA==
`protect END_PROTECTED
