`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TtZ8ll489pY3lJmFNEQdj+KD8WAvNmz/7ZUhEotAiEsoQhX2DENwVEDsulxxW5Q9
8MMnXTnBCNDoQI+AOqybaKnOqfbs6ZPxDZ4FbGzuzYwbkiOgtD1CJqbm3Yrop65n
WlVKnUkkFIteXKlEBvJVlwsnmVVjjQwiPSe5ZZu4qCJlowt47AJbbXMSpY1JNY3i
pWczj7y7c937l9uhPf7z9oTLSDGVprjFxVpr6PZ56Ix1hK46C1WMVnCA1PbV+BHk
asS7SAOccIT37ynXm1YO8f4qJlpzsPkS8ZHzO00fuXlmhXXIOfPP7PTiuuqtqZIs
rzXUgBclUWiXgN7Uam8LcQpLLpv9A5YwK30IER14liIwyvpwTp/ViWZW+IxswR/3
tPOpnGyRbiJBoiqITXNYDdao9gbS2Pjj/wKOaGxRinS1NeSiDj9kutTveQAqfdyx
`protect END_PROTECTED
