`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jG5rvqAF4crdtt36FiOaFGN4izAOTneLHO/Roia5I8vjUiAsalQYe+6gTPFLBm4u
7Tl9zThx+W31Z439hy3o4LrVTK02UTKVp7njxjUm+AXKb4pN2FQEQS0GscJ3onsR
6oatWe/DF0KGYebs+lSl0Q9ZONxrnKDbuq0SHutcg+4RFk5dgnOJR6ahJmaIY5S/
J2J+3JUWJVteRdQ3huUpcRzM1YXo6TrzNngnoT7+pnQR6glQlkEu+AftDEN5YyMX
QeJ6mcwk+2saF/GzZRStWclWuLwY01r8+kGpUREijHgqX/BYEvfTtnPQIo6wveNT
ztLXuOSSN8uc6bAbQFWfZWOQstam1Ic7os+W6M8BHxE4AAAC+dh0GEGsQ5bQ9EBg
liOdvaIM72ySDCOKbBjjgyi/E6V5HNw5hZE88iWyclg/cz+JsWPBhs0uELq9rzSv
`protect END_PROTECTED
