`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RCXKM85lbcWtXae3/iqd6Culur55+Vz6O+eydCxtNo4U0QShjOWqW3j8V8x+sjTB
2zq8hfnuNxFz7b6vgh8gL0JTULcxsGG6iR8eHo8l6l/rz2X+vyAmRSrKp3t92qvH
Bo9vwVX8SjjWStD2dOd+PuSa4JdsCBuhK+19yN/MSww8b6h3NGPU+5RQrSzAOr9x
nzeQ+j4XV/sjE7H2z7zvdBfj+NUNnqYVejDU523kIhhIutBlI36YqZBnh+gTmhx6
0MIF8b/W0auf1zv1WjkHSMWvqd1TrZWM6BsFFEQVQLdQ13M+uPNLiB0VqmbFJYER
l1eYaH8TYTwBOIwSHbiEt2CF8HfqKMll8c/HjBvyTfavzgUbMqhaLlRmLRyIqLAN
wCS0eok1KK4TQQwpWidtHqc+eKnqzL6lCh8jBqSi0oW7Qjrtp7eZ2RaXfs9EuvTx
`protect END_PROTECTED
