`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kaWXRcdgVgg17df+tDgDVaN0PV8kr7/v+iuloHFnBGd/nz7PLHUiQSTt5Z6MhT4S
uIz9MIKgBx5GKQEWiBtc/K/vjRGeq6k/5At7gEHyic4vsd3xwXWz1hWtKznElh/0
Gg5pWvOUyXy0i7Pa5evqyqDNIBeq9xGQcEcclv/A3pgCy3qkzLubQEqvtjtPVO/9
ktFgoxAZYMkT+Gt9whcHALpBn7PCOE/90BKqCqK1SuiYkzSi5XBYab9HuWeRs3Oh
hBCIOD5h18BEmLDHw8kw+F8L5yYXQx5lypjrFUeoC/FZt8EsYM93Zk3wG69gn6Z9
C6AfkRp/OmiQBW+9uba0MJCkDXN9SlHLsyRoNPXOLaNdCySNkMBgsKJhrJ352RiO
82UzI5ersDlOdWw+Gpu/k2jXJPUcTqiutIM+8nngdn0=
`protect END_PROTECTED
