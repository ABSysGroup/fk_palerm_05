`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ypuS4+h1GPh03WPT6d9ygBNN1myTtT4mqTZXn/lJd6DWlORjXfoheArT9MdYQBcs
5aP3cKRuDlnXR72bo3agDFokqH60YMdVzRPXpoc19oh2AZ/LpiAnLJ+JSXq3RbCy
Y4V3riIEptA42EMu9756q8Rqd5bxcy+OKAktNPeTO1PJaM9srFhVNfxAoS2uNWtj
TRZRWxad9kO7PjRzWAV4BgWfVWP0kZSvR8OYfoTSYvjuRfvOEx9wJqXaJhPrvkW2
kGsYfzr8YN5WPlBk5Dh5UMEtwrcEbb/AauJ5xxAEZR2p3J3jRXzBmMeVMoQTYmal
o0HJQjoN4CWPcBqE9s3gV3bIIorzFJI+6vOuKWY34qSRrEHv3L6cPpUt90a2yfDh
BhRm9eZ9EdjTJmBdY/Rxmh7nf1ZqBs5zc3nOsWs2jA8HLMoNeO/2WxqwXSdQwS8U
vEomS9EXw25EWHMbYeXagk2dgdhZrEZCFm+A9ytVoPF+4EHT2sQVe7nq64K7U408
e6HjIBUINNd5ZhQEJfvZNzAIDdIw0UhpY4N+3/iwhIlfAf+vG0UjX2MMdgpWzl2i
YDrYAvQb9izSh8B7jRvmpCDyXGbUm0xc4SafWBOQPW8fWpWbB6j8BGzZdOnfR40N
kJSJDT5K6yJsU6xt6qIty4bHG/TuL/LgqoaKr00WxVgZ/HSCB9wGah9LXaEKaAsW
IvQ2Ome7qkpbuWy/8rj/W69W4tFG4JVS1XgSd6d0AdPwdDxWHlnShM0/RFeJ4jC/
/DPzzOc8oWiLKNInZCbBWhmnuUGj6lohGUztFcxsef2XJCU/cmwVSILR1D+AMbh0
D+XoAq334vgrnz7El6ZklU9+CwjPx4NjTnl+6/CvFF+GAWx+jN626JAsVTtHy9bA
HShyjcpo0eMxJhwm+35ngymjVnUbiwcnoad70D42M6HQ+OsoXcRIWiF0odKIogpo
I+BXmO+shV00uZfDYaZTAwhhtuk0/1qDGDceoh691VV5wBu5XnoSs1X7qwvZhxhH
sI8hHfb4RkhG+RzsyxXly4ekm2/LUZkMZapvvj/fqwG2FV/BPMRgj2Yl1mZDULBm
/YiQfES+/alB/phH0MWAkWm4Oi5TjRtSOVgIEB0SPKoH/lQnv6SYQvkELDemeQRY
v85WKq2qg1PPamICJeMTm8ZSpmNxW+6m13oTMTskJ95LacNpWzRWCZWR4jN0Np2W
ICHb2P5vnnMK+K5BGtmTCF1AjNWZpDABaCmpZA3DniN3gUXWl3uEZSKvhg1RjhZs
5J3M0Lks/XSqtTCxWyG3JigVWi2zz3VBJIb8xXnlGGyODe+SatUolHs+yOtd9Gc+
bXB2mUa4byTHCvpox0rLBK/zTKnZFqGzzraU2jJ15a3A30k8xoYjj0SR5ukMfZJM
1CINX6AmR9lYZT5ShmVOkb4WF1ecQUmDRv1qzQhyOU+xeLxe/BAPIlnpGqKzTiM3
fh+OzX3ndLePB4PfXOAyOuuYfEj8PAay/lAQ2nLjntFSNh04EvcgELtx2EGn/cTQ
tykLum4eeofHnKsy2ezMpMPED8csOVISPBtjAO/FMTqFlC2vzx53uD9U3ZnLtBzr
Dz5Nzg6U8cWm2UWvJqAlGmBlwynSXJB5AdAdc47w0l32ta27ie4IcV/AxPwtr0cJ
1tkIaqybtmCi9alfYBwY9y57OLNENP4jZFik34a/vD8NZerwv3c97ntzh1Eroh2m
AHjflZu/D1UkD4xzmmmXY4645+aECz5wEkav6Rl2K9FmeVEPXMOZ9wUnx1jXui2e
jlX6twbPdNM8avpPeoW7nU/J3JXKKF1Fr8tzO3jVbuTd++vtisPcude/AOnM7hZ/
nrQy+4NJpogDQXA/P+sdHA1dG29U2CuBbwGbNiJ5Cfe95FUEZ1luuHpjPt2SBEbZ
xCEYmB0RoNZU97H5h2lBBtRVwn1IIhRprkiy916ZzJLc41LEvjet0opbOxdtfth0
gn5e6bIrYCBXuRDbZ5xavd65HopBVqlL9iI5FxFk8z5Ypgf6TJXVXfm9xXPTedkL
QJPfEsvBNkRvY0xwlRkAow==
`protect END_PROTECTED
