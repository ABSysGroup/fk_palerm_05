`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zJUuoM+AGnUrEUVZkzrE12G+AOPFoh/KXIZaCKA5Z61D1Z8tcGyp4G5P/HJx52B0
t9gmE0nj+TuuUbDLNjhv3x2416V+iv1weJedh0B0cHJ5smG8YRHQPzq189c+G4NV
1gkVQU+aZoNLbg23jIEOgD7ASAhHYsjm/L38+bFky1X9gPHeDN7Ba/JiZ5S8ObZD
wwYJtOgzfrr4zk4XyXCXFVez+8ivhj9IqfVZS3e9R+JTaaiWMmnYSB5GukxWhpbt
n4lrjsptIaHdfcPASg3T3FAAGgu7o+7OOiGNdcVtg21DAKc41DKx+zsD0hLObtgc
/783o3XpUXnMzxGS5qHOthHeQbxK61TluO3b8jqngEA38RXGUswZ3VXd8pbUTE98
n+XEGYxkzqyTE1YM3W1de6aIk7JZXf0ZeQnNoNAIbwrsOH9k8SF1cNYVeQA/tjVy
Tz6o8MwP9tciHkptdcSUVxNR2TdbLXn5Cw22tjoFUap+XROj6VNmYyZPAvzso4CY
WinMzvQaURChlVqGdEcn8J4BmFar7b1DEswOrNWTNz5yflBcqBI64kIguooysmh0
n2CQlHyx2T8brXjIgEyWmUHWTkx2/ljJ35RAUvWQFYduontXOgaNJevCcRwClOhB
qF9lyGgF65yqcFtRQ/pyE8UIbGAD2ys9Ua/+G0HNC/a+xkT7vbRdVJg1OMqNWjyM
`protect END_PROTECTED
