`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WD3c1SKU7RhnvxXsTo+lNn8xUuWHEDNCVBwX4waD7NQVNyTU5rw/pTQ2gyb4zE4r
qxyvIJFmve9CSQJa08rtFTQw5ZZkPq2/o7pnqWyZHJQpqWec7Ohxxc3eFeoEzmDM
JNxnX5zSXwt/gw801uxGhL5w7RxRcqwEyfNwOQJPRBvzF85BGXjvlj/tVUKR+/o/
bKwX5iplAzXOxbxlf0ynUN/LfaUq3+4LIkfLsyVPgOIH/ylBqbJVlpqHyOH8USF7
5bLwTqBnTiibl55c5+hy+jylG1aBhTM2oguL2zdjD4pVwl1d+NlDcVZyyPS0tpSc
SDlqVc0zoZeuem2i4UeL3w==
`protect END_PROTECTED
