`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M4S8eCwsNKvI0F4QU11rdVlUtN8r04n6lS5HE0LTQ6jAlDhfNBdT4FySwn0EV8Ea
sj742Q7r7KjOdBDChzD630TjJD/V6Yx3dcO0C90uYd5T5PNIZGOPKCETrXBwXnnn
tqIFu3r67e/OYMoEXswR/PkO0YI63ocAxZt+xf3pHSQ3CLF01R4WrwIlbFd/HXvj
1Jd/mOJQoMQQfEvVdcArWKVP3nIup9Tbs9triZqBaIlqUxqbdZ0jN3VViYWuOdPQ
S+g+hOPH6vVHxjbj159ctN2D1FVA2p0Q+UAfr0u2a/R3aINgPx5ngXorJ3kQbEoj
QhN0by0bdX3oyMxUmCDabmy/9P7G4iMldD092+ONUmpeoTSZqEqgG77sWDmfO9Lt
QmfMkP7MC0ztslRSXUievMcf+BcZj/Hq7q8cH6eop+zpoMwLlsZKmDOQj1BIrBbU
iQIY6u0OgOdmnZLTVVWo/pZq2oUHihVMBXr8nvJpDwix/qZXgMD/JFvNODEYY6W7
0wQtkTg3cU0TPIBpfgH7UBZIvIlwUjJ9Gu1mldrK330=
`protect END_PROTECTED
