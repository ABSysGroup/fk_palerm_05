`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
41VJtF54gKuflNNnrC8cXGv77uT5caHIMwy3BRv7+kgCAmePRhnkk6vjVBY9gzps
y+5Sd3Sw1UwUpYhZ/fMpxafMkHeVEZaAZGh+SM34N71Jw57p8KFnxjh5Es6XfGMa
GK/CCLpBXc0gf6p/F+AxEdmS+z8avvo3U3U/QF2Q1Cgf/ijRAXJ+LeeHlRSNX1CN
aifI+aemSitixG9/MRbN3PnJQN9kLrkpQWiP97kspIFGkPFSWQvvECD8xj4z4Ocr
Ykc7GB2OIL5PwhSulymdpzUlBK8G693TrQDL74wOSLapFGCwQipS4pZNftfqIGS3
acMlHze8Gn+ZCoiJyNvq+k6w6YLc4lxkRtZqT7IXGwtL3OsccMmbqcZZtOGSNMKY
KfKQl14d6zV6ZOIkUwAuyga21Zs0CtnfbX4J1D9Ry/A=
`protect END_PROTECTED
