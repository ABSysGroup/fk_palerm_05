`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dZdUOwXiKJ05nHXffEcDIxMPz73FIHCN+Fi16GzCYA2T4Ws5/93d/WrfH8aWaBSr
Rj+12Zs1QxpgiImGA5z1K/8zxFGoi09bqhqIW8O6V/ij/SM+fdTlpduwVQ8KALQA
MQuCqr+PJfg899OxSimowD/aJHG9ttIB5yDzcfWvxKOp4vJwypKbjezLXH+uok5s
euR8V6c+YMYNF4wX3bgUYkI0itrQEtNOeGnQVmfd0xPB79zxk24bx7YQzpNnwgKG
TzOrobeb+yxQ17T4a+aqog7O+RVrXSoG6JTL+dI46qtEzg3I8aLLLG8X0tNc5Q0A
4oGK/+ATb+rW6YI16pjMjzxrLFXiVxGezMLHGKZHtNEpIgTUpExOjKhjAZVdjX6d
`protect END_PROTECTED
