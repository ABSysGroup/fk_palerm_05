`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lySMcePop4z+1GBH8bqedQZtMGuBr7bF8Ftd8OlpCh3P5+XXGehfwdQYwW0f6+5Y
0QktF4/L+kUi9D/2R/LQlBeK8MbNF9eZzG/9QwO4ZoMKJPWcjTas0K1n3ByxYOHz
FfS6GTx5/+wyotjw7zLPpNpdMp41zrqWrUVF80316s8t8aR2twp4QDxuWC8gy4aZ
zz2X5V4kg0AX3auLrCupkB8dgUeL/IKFpTExTLIh0A/U6yUMLTihie8V6RHxZxeo
bsjgiUMW0jx+++7ESpvIPDCScmDkQRtM9xdUwKlxG0uYR3wLMKheFOT56N/LRmtV
SuOJa2vV7/AOcyAhOy1S2RfBaCiHk6ZgIFDjHefHfYaQMlV4JXldWrS2qDBvGe94
`protect END_PROTECTED
