`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aAS9O/eoC3A+LlBcQWl8Ck5DiF0+LtCKyBRDuVG45GWOJYROA7g0BvS3AFnTZLzY
R5ef2BLt/IzX5S2VkuKQT/FbSzua3ip/NmTAAmA1WIE6J0yG8hSuIoHK/DIV9RDT
I5Kvz8/B5b2vZ+S1/H97CwNLfE+7SHFDOoNa/uPmQFbJc8mbAJJYMeuYQ4m4sKAP
HmBqPB0VMisDuEO/dk+Xh490lAXRSGlcG6iKWcge4ifVJjKvJk8V54wjVOsyu8XZ
JQQP+KJ2RU79V8GUhIrXx3rMYVyWXVT4SjTREI/PR0MlrDlC/7WOh3cXcEjMTjb1
iZ2AFsDbrVGsjng3+8y6AdK0rb71j3OV/vnfC9GZnWDZ/v6TIAZQNPI/K7zQZFX4
fwkl9zdw2FL69ko9WX8HHSqhXuFJY6Z00AaF1c4HUp0Lbq8Qxh1xpZ+EN6Lz48Ke
y0xBJQ5CsyZKC9IFekYz6JvE0kzwfCX+4Qs0wmpo7na4xnB7sYrQeCeq7GJIoca/
olPpukszzYk4x8K5pR0YC5gPgw7mDbEj0Fd5+aikooMCW3RIX7dNuTA/fSNk8u2P
AhKt5vI1WA78niUXUjjiBWCENqgMXKdWI6F7dX8Plf7hKh0d424Ur2ZBKs9PWcCI
f0nvtg6ieZk/++oUdnI3Yw==
`protect END_PROTECTED
