`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PMPOHbZ2R2sgxhTT0wV7d4p/Zjrg4cP1Hq3rpF92RotUq6fimZVoloFtc6MboRRb
e1580bHOFfH/5O7TgiZ/dNCzvi/zjHDUmHGZNpUacT8GbQQbN3p6sSeR902vE3bX
+kjBqSir0fr2XlAVbfECUExyoxUYjInScDalhIncoIO8h1zKGJenU3rTokdPPVf+
hr2G2ZtUp6FbNMz+loCVGVEo9CJ5Ldx2FVsVLestfmqopZ0NOvsNvnwicJXDJ61R
T9KqNWZSCmla8X2cVHkZ9J4JLVvIM98ZMQTRVswYj2L96xGXHRANErsbICEcGRbd
C1SYD8UGCN7/LTnjYD631dxHyxZsRr+Ldl811u7g0QjyXwqp0MEcADWqw3QcLF6k
StLZh8EsLbuSOFsE0UrHVqgxvQMKOBcHBemnbH5nIvveg5RrQ+Whj1hnCA0YugDl
aZufD+1/tqxmPsoXIpldcMoraogmzT9fxe2UGyArBJFNBIHl3OwaOyCscjtEZkMD
8OAgjNpchZavlikWLDj/y4bXMoh6ajE1cktT5/GLfDlVPEDcEKF/lLUJ6nnpREOl
6xGSTWjdA4WRWSJdzF5tTDTrCnTs6e0CjmbOz+L/bPxrLJ3AzDvq4WrEAnrE+H9g
wi4i4o/g4hKyUwYmuqUdA0LhgkUHfUwHL9jXi5OEIJwJroJKSKHlUpyPWLmgCyYv
iTJeXcUrAfgIZztb9qmztOVbNTehNWm2hYdEXy+JW3sdE4lkRG7nxZiwJv7KEmH8
PFEb94JyeLGfCXRT/YQnT5Bphfz8pzXMbg9G7awp2saW4K0f1HDDmGng++xbm7tD
GrgFOt5eYK8SYIMYZdORn3AIQNJn+3kvqiTb/V6acJwe2TeK2s5Wwn3nQ8EL2HKw
una36TVB3XmSIjFsyqgRju/LHIRItJavPEMDaz23YbGSU+5C7bBGzUAA7u5Uz9Ir
NbWCTIflTBD8hR8wIp6po3PfUuvmWz2naR1/kNPFVqET89kEoe7T1IDZ6iz06dF9
+m3NM8pq3QiUqNMblEoheDMEe1dwJbsEqhUEHm4eQj8cYUpHjZxttGqgE0008/zg
K/+q9OsUffjRqWUkqvyRBdT022NeOU1rYMdkHbsq212B5+v9229Q/003Rb9sqORy
uWfP6p4JccEtIy3itSMwMSDOBVIA0PD96NCT8V7vrYtIdqBbNlKH4HH31bfH+Uto
a9TtcYVbXEHPirzdNPmvQbFTdKcyJaa5V22vaqfJmRUtZvYLZnjvp9LUv0JWQtbW
gP4cQuGczFW0kp+0z3kBM4YOcdM6N6ifxIOKFc2o0HoNd69Tc+aKiLVp9t66ONjy
QzESufMtHMiB8ooezHGHw05pLtZVyZw6fKJUS7iDe2r5jVK/ur4r2fLEPQ0RDCF6
I8yZ3zaPN3Uz3YtJ4Ab/fHA4LpTJOkkWU7dUxbg2iPNRj2ETFGZSskZvul+U5rcm
gOQ/XSboWr5f+AmJxrX9S4ZFxORd/5FRdrjC3I3yYvcXr6jJ6ujsK/wZObpP6ygF
koesjSYRQLsCLhbb7FNKKkMtd2+GYYKBtn/7ieNhjdaD69OjKHgiijvnXnlQG1Ot
f64P7FaRrNHeHVBRAuIwOcIu0r+I9tcoB/SJI+8dRaa/AufEUFZq55O5aWn0Fu1S
ukok5jLyG/jLixIx9n/wjopJ+qO+WTgdV9asSHn+QeEeKj8hmHvOleRnCEhV2yzf
aGjBq1gANJHJ9TsApQLXy9C580NTqDlY7emScB5GYsBAtygQziZJSlU37GYdEU0j
HquMuVVnpgQ1jtBiYEjdMSAUPvD/JEWYouAWNHhZu6N9ko8o1zRauQMYjfVEAVtP
PqoVl9nfi/4iOEdZKXju7GhiaN/70EoJk4FYYT0ctQPGtZyIzMgr/3Q4Gu82+jJN
ONdKJK4jZ06/RRgHzc4W5C7PYyg2xwGltwBn/WxFysC/MZFPg4fPXXQyNhiDnxji
hSYR66Vyx5WsnfAzPEdROJne3dwK8peinu3x3/Lh7igR6vD1mk741AwT6c5dGXrz
Ta9XgLFVvmMpFrdSBxnePFfQ7kgDtIX7HpHq/guVKTSl7ydxcc23KqcAUV6yHZ4y
m/zjhy9M4o95gcvkR1Ca2vlelhj5sCNTnZv/4njUPKfmTXlSg8+TVun3l8i+LQKr
CYdT/P0aha3tGa/kv+Gew/0X8zZ1SFbFxi7BVvhV90JiL7y1cy8lRpd/X72mP1Zv
y/16AzlLolM54MiHTiFmWj67aTQ0pSpbcgK8Vde4eE/rt8RsBh4UtGPHeZgdUAb3
HFlGcAWF7nVVUpjd9NaYjTh5d6soykLHSW/tDmIeMt09agsDUM1JJz0hZ1GrMMeN
KpjiJ4CgS4SDU6aRKe2xj1+TOJA8U8dDWPDDS1LXQg8N1W1qaRTPHpxEZnRt1zZt
2LUPzNCeetx80TPWUHSrV8P/XiDTrrQvcvffkKqbR1IKZtE9gVOkgbq3wTL+8OL3
CcXJdI7fQ3CORuh45WuW0V+8NyUA4tgepXRxzmNZPm/EiQDm4+49IZUB9UeR2Z46
0j6vLLaAIon9fGzIFy1iiebZj/5hW9RxdhrKbc/w1Lu+u3pgIQlho/C6cDoaQhWf
GufLT7RSRKxbx0/uMf3YRZaw+P+sfXB8IX1biJKoiuJ2xiYXB3a6djAt+JZMmdRq
kTS8VIdiWVUz2xCdAgJWIbYr+lyaYdLtePk3b7YNjRXT0NOHFt9wnTuGeHbjMe1f
IuiCFB4XrzFkZ9m09BqVSmgewcekD1qJLwwgffw0eMk91O+gCqEUr5BIKSPljWVv
/IIJIycTvi0P5235+Me5Ve/Z6b+qWP+4I670ut/9FA6shhnLEldYlVqNfl6v2+E4
t1pnkIQFsMQ/XY/vmTzJGOnFJTTAkB1F6O5s2G/eAJRyI9fVo20uu3Vjm6bPxV8I
HdZb4tlfXVXQtWzWhD5z/i1fll37rTy2PhzSxTylZdr0M2wigvcQs2mZjR/Flijz
jl09VaPCs+wCcKwI1qxhhhDztuwbkuHShi4UJefxcKRzhAkYY4PfifQURCMDxrLj
biYW6ihDm9KDv7/326LTrkgyyx9EfcOGs3nMi8oi4ZyonUUekdb34tHTOpbYVUWu
pqxKAg2hTcQ9MpRAXXOq6myEpR12mLqnLb0wGE/Jky/mpEXJAi+eqflEEMvvfysJ
oSreKGok872jOYYlrH6jGdG20U0YsaMt3e/ZJGeG1SeTKZZVSWJHBjgGeypNyd2e
pPW9xLpC3Uw03dh8PmXF8Uqb+khQ5V8RNYOF/SDeVU/uZnNUv0PGSOZ4p9a4iQe/
hycu1xhK9OXwn4LC4uw0crfnqm8y+CTMxFQ+7rY3t72Vl9AtNXUcphA2vzn1yLed
JtSyJfgLKrmzv+/kpDM7QRCgEwGNzwb8NHJW4EUdRFOLdNrRtITBKKNfRUk+6mqA
CZemwKH6ioiovX1h4stIxTNZdd1DuZdg5tIqCtB7HTAmx6ylmsHBIxxBPxu6wdOV
MOu9nA0Wzh4d7VZqrWRVG4a5J8cDsz8ousMFfxA9VB0JJObPrd9GycI8iBWtFvfn
PIm0xd1RMgcYFHqJXKQIyKs3bQZiGLW8ZTyLTuBt3FwBqnbPs+PUFYYH6EoEt9uF
16iLVzvOubDhIui2OEkaPxKdh2CD+wcBCgIf5RZZEkwXj2If8rOsPVhM3bGb7pO3
z2wr/FH4w0debn/VhUqHm4vEADYxt1C8Gq0BrzKh9EieLio5qlEtLej6fiR4GRHc
lpVcZKwlzpU1yrosj2CfMm/pxOY6/BplCvcnlicFrR5SSe8qecnJSU7eQ7QC2jEm
rn6DdXEBokGWsILXrtKQSlTy1w/jo6VcK2935B/VHKORYPMiuTg3jD9RulDDMvTk
tFtDRp97LSZbE9SZGg6dKV0u+HaHmyd0qOMFa5P4vWqHpdMZzRFlCGkw9xKmmOnL
hYEY5O4nofLGBPRHjaSgS/xF2l3ux9RD5NZ9i5nkFEcvz8gdA7Sa5I38RSPVC247
rwA7e04WtINUZ6e95nTuiu9f1jHybDakl3Z99XkXraWvLNiDkOkSSy5OMiw8b+p5
kdZrsxDb9z5VjB6PeAD9o3C/CQhOIvC/LZ69v+DXzCIlkGR/uMJlmYTpOcrnZXuC
fD72A6hobPM7/wdB+SFqSgV7jN6cELXJIGMwOpfm1xOnOzKcY9HPqYkSepesSM0h
Pdk3uxFpVt7uNRV4ONuCatbmaMOX36JHZd9+uQ9WkPXnRQKA6wngmlIR57E4T/D6
50iT544NZbOwkzb/ItH/HP66fhWSMc/+3W3LR0XW2EO1qLJ6Wpd8jgad8NqC1MlZ
qwICKEVfJit29S9hHKt3/72I3YIJVme/w3vrZRuJMzu/tVMhZIJseQi9CPrq+ScW
EJRkMD8w8csV86s0GAUaEXg4gZQaBqz2fxIM5/W/ONkHopfpwjBtDvBTSA4S4fXj
aFBadBNfM4R2u6nye5/yLcJPysccsnND7G5ZruPdVLc1cT5gYcyLasBmOT3IiM7o
oQv6oWHc/nZIsN0twYp8wvFLhOoOQs1xVwxM9ZMnvNdKqw39tGPirEGgk2i/Jr5r
zFwxVnbu5NJ5u2tVw5rcywB1xoTfKyyR6t+961YMBTldLF+BY5XNE0RN3Fw/waIJ
pooVZFs2pxHIT4HPcJI/r0qiyu7WiQl4ceebkgJnVCADrf/grPfj4DnIcDUrAPXh
3n2GWO7HMm9W7bcou3AWqKsc2bvoO78CRSRxTFTVR7eSCmwTNQC3HHeZbEi4cYZ3
esGU4hvSMILCOeNj95ER3s9IaX3QwjuM/+Re7Noj31czzeAzniIwvcRoAcEndUT4
9XfRayykZg7SPrHAz6dor9SlgqIvbhPjlunfJ/Ny2xLhwGRca7O8br1FU1GEMDaW
EcTEsOxYDvXqXLu6+OXFTBjWkXqmmIu9yzkFSQiB/5xkbnB7A41REN0Y5Vn0D/J+
khNmmZZ4Hc+c7BID6l8GC0iYAYSrXfdzjWQG+Ae6CwYv+H7Ijz53ZMByuPbYgv6O
ZTNve0l230BQEiyyqiy2Tv+qJXT64xjLAqE6JnbYyVeGJiNjMBJCLN9Wb+aBV71E
xV78ioVsNn2VvWtcJvvzhiytAWYJQtq4nlm1AByI9hcKCC13vDMGRffwAn/Z7F/7
isdrOO9FJSRTLpwZ5HIZJwsujnmW3ekejlQPvHFpm8yvhazc6pEDLUedTAOVU55b
hlsGEHuPESLc/C/uy90k4T6mHdMZ1LEbuzCuJu6Z5OrNL7SxAOahqvyufafbxIm1
EsDfTLXj4G6EeSRPVaipEvOzfqPR6ShrSMKVHj+5HrI4kyvyqUempcG9IhasyxH9
tVEDfYJGuTr4VAkOzKXaybnGqy/jnx/Ff4C05DsD64qZo3H2OKN1pbukRkaZ8ECx
5noBrUMNTcDep5qzyYlDP4GQ3LCGbK3Zr6Hx9iTKswn71TT7arxTb4wLyWU5f1Eg
sIrJZ028OVSzIx1v776u8vReBzmnb7hricUYUbm37opPcQWIzr7iFUnbSuBbeWm+
vmC2O2Giek2Fyrm29D/5k58A9uAGqS5KqBdmA5xs9wIxhop0XyUAwGEsgpWIRIwS
jOgCM1377MvVkXAeGB2didA2kDzYB67aBA/Jgm9vScjUWmwtnYtAIDpsKVFjy3xq
wjSLWlbOtuNaoomZWIt0NV03HfuGUyuhB7KEtuzOtxME5Qx5+Q0TbHI5531ReA+5
Gd9Uk1yyKBALKQpmEXYI0Wa0Tpri66/WlHriAURhnuvxt34aOYdqJGSeTpVC49Mj
fvv45W+Q6fwaDNo0nQVqBBek4vo2+81Ix/C+jbLm/cNukiWDj5pxM6LeOQD+ihx2
eYfoI4oSdOUp5o3lRsUg7WTAU03V1UT7zz/gZ+YtiHVvdl2/zlK+npfvD9pBNjs5
8pD3O/k7bJ/84bX9d2BLZS0YW0DZM5H9fTe/OKD/r4v4rUQ95bDqWi2qn5xIMRxn
A7Gq1zfxInjAlehiKdFDHDe8cxw/FPgxLnuBL4R5uwqWmvGWum5uBDAWm+hYCQEd
EHQtisQEeGsuhIlEATSQPzwxhSF/PhBfr8RkVD68x6SB4FMJMbYwmkxkzc8tFnN9
uxyLtHEpqiNsZJVIh+0QI902khyNJaW02z63F1evM2kXlqBGwFyqPTVrp2g1CG0g
jlBu5165D6T7VsTzmORjQVbf3xaD6fLdao4Dd/PB1Ktj1CtcLAwFEy5sAwcByEw7
tpNW7Gwkp5477bD3opGJiTnhJUrx/tGmalDZrbZVJS7e4pBtYS22xzW2FKwNUCa6
151TZ8Mx5A4meXwjHmiJt7b6KuuqSwzSX2jSmC9lty844i/rL5/mXjhvj39bIn0F
mEK0kuQ1pd5pzlkRgABAfVObu5+JOSefqQTX8X+68E76wOTeKaY+ntZv4j8BhyPH
M5eFsxbZyRJUzHNVY3SfnYVu+RBgkc504+Hiuw/A6HAjVXZ8Q0iMVzyuc0DkwK+8
jjocJ4BWCtLr7YioL17dTlkoE4xzkRByycO+zDENo2dq/vuxw4qMEjVxYRPcswky
werJcAZlkguWI+2H+3goqOmZ0XTVkbwd0gw9a5Wr6ksBZlF7xOrTZXIiyq8+UmSD
Xd7ntQS67xcdZ8N4VHsNLzeccWHhYmFpnkMDaPbFucFFWehD6OdPVDF6AP6euL/q
y8CPohO8EnZBEncLdF4y8hh4a3Z5b44EGRq2SHJUcp/R+FmcnGdKH6mGAzDTyi4P
b7G1z02LfPzoZDumfdqPJTNI7t+wvV8lBKFN3QYWTjn1me/UDIImfy2myrklvx/Q
ONRFKUrOHxIFw/VHWonQE2SX5w0JYFxTp9pkKOL+eXa35p8W4s1sbZP2z7jPkStT
on4c3Utlfocys1qshd5nde+ellLJf0NVT86wQYvjPJXKCU1P62fJCAAGdL2rIIek
Wrf4t832tOpjdLuYGMdTANnkq2Ya2RaiSGDlsJ033TGfThnJ68kP2eKsGzwggSdV
sapVlH0iBdnInYeLRFtJ7SXuwJxRv+NGJIF2Bm/binumK50KR4/Ohz8BIkklHUmZ
XkHhlUUQp6tBr0EtpPxlINrLq/B7DwmGVWoMmPQZDinsFzUABjLGjJuGmE5ZJ0Ry
+dO8mNd34AQIuaMb/C4xf4xY9JYu8X3/lBgUyEV9aEimOwJ/v2eXq2QZpEJZoy6E
YbUJNOjWwKlNQG7Vz7+Cn19k7AjW5Q1Ce9j9Fo20ITiUSdfQUeTk3tFDuWvsOnki
WbWJYUm7ktZOqiZoqkkz94Difb6VAk394vhE+E8ej3cDUjyud2AwAupJmPTgZCBo
IpSTL3cgRDFGFwasw8kYTSCXUUOG4sSpUG0uQLajJG0lVZ1x3md4fJAC1IVpQrz5
VqQ0L9ZSEWh8irolRDOuYWBoSerhjmgnuDYlUzQSKv5ebginvYgOulxEELZ1lZmK
Tc09DNFonkQnb7VcMwZt1uq6a47mE2Aox+4zzcDdkJMPU8oT+GcUp3uIPvLahpMC
3phZqcTq6Yq4f3JbQ0xcJwzp+TF7kaeCN8tcDjybk/+B0vIwdEm0ruDe2WLYf5yD
O85XO8/ocMTIMrwUrlnxQZZgYSSKdCbWxPCW0RgGSsWd2W/lVnxCq4MHPyBdkhYw
AiOzN83XjBDr7vTGxNxHVzSPqGTX3jhspsSvpMCAYkR3hAcAD5IIUC/+YjBy/PAz
nO/0Vy14PULfRVKqG+sHw6RpdIerNmvtiUBwvdLUwDMNUJllMKb+6tcURSCulMuM
8JExzXXtJMFQo5gCgXMDUF+x3rnKocYdrxO03TztUOmZdKbpJq+0D9+QvxRmUujJ
Pdo6IIjnXigIw51jG10luA+wrmP1DxnpCMcyG+zfGOEHV02TulIpVPeDlStITMHc
PmfTkP3Le0NBHF5sd4Gu557LC2tdvVPNvwcOXD62KF5Au85M4awSdq6xcWj7g72X
Mif8GRcVi4tp/NHttvH4SYSEE+RyN3JgYRMA9AchPeukYfm+tyCF3CiE/7trZj1z
A7UTfdxNSO3hD9nsV67HqbYvUgGq5t6Qz5tqxnABamnQ5Kj0fuh2hfVsug02IcBw
lDLELwjws+tNwZ+Pw5KpuxAOe7y+70rPSFYq3ocYX8qjvws8g1noeUskYrMw+epA
4xDtUktjWuxPD4tntHq1IuH2MvEQRAvOhiOS2WRNJox59FBv7XI+iyyc/en8FL0V
PUxA3o8KZiDItb3WxTYMH1lTwUbTIyF1amhsDPaL9XycCdnI+Zv4Hk3wDWBumqQg
cmYroDPmyTH7sBPdZR3oy7UsiRePxPVleM5H1iUUS3cqmaREuas+1Y4sni0699Az
D+pBp8ACdYFFCdJprSxYy8a70v7Gmd0S32znPfkzFM+WadCXT3v25WN58hHv+y+n
qdqC3x5v9HUUBVsCvYiY6e5Qp8sLp1bhvT0yIejY8EW63HguB6yVi5YBmiOPFRt+
P/1ZJSeA8F8EQKtsKtyfPuD41sa7N3AEsh5+6sCvHy5h5+tWHwppWyTJTqONj491
DTM1QIR86qECVDDRFlRYxRropDS/nSq/4rUBTrpBvBKwm5AqohUP3V/XogVG43h2
CEjZBm0h0Gaarxm6xWB+O9fo1jju9nG7aQTLfy5Z+jX3eCs+JZTybdEymPVZhbN+
MkCxxVAoF1pyDt9XcvkxJnAU0gBpf7QGBkau1wKs3dIlUjvu4Ba7s5gijDb3leqU
h9ef29gI1CmJJxDSqwtflcPa9KavY/nmo1iYiGiz/incpy5FmkVOWMLEJkNbI4Bw
5DKLo4kgTc71/Rw2lDYkWAdbJ2Op5auYVPyccNmXVPIr21cudJ5fvsaU6vzyKGKD
eaTfeqNg0pQTX18qfEOlEJgyXImGX6dY15L8obAfBK4xvjKNevBC0gyvR5iURlpQ
KJ7/E5Ao8e60b5ves8s0nulhiSuwz0IUFqzhohoqehm+VMmyGIXAEHru6r/8f3fU
Ddul/H3XDFIi85FkY7QucTUV8QGyYbR1CN4+4jMogotBRv25Fyctd6bZJvwOYI5c
edLPRIRJ2C+v9ukZnzC8truQ3QHzctFeb+VEMUy5/wslzBByIMUBdWmOthAiZETZ
etlDVjq+mCfByuHLvdGe6stllnyqa1IcrjL7HF1Bh6KH+/lGgx9OdIM5pntBwYOV
kpYCt3RSjKMO8UB+8NawowNRa4zNry7Qm7Raj1vyetHlczNmS3BevqSLTsbgFZK3
v0U6F3b5XapLFNoVjt8edOvlZIKisaiL8sxczoSaeCd1Xh7cQxrdZHbjJt5D4ikn
KqNAmiwebwwcvW5wiMvGCY69Z63TnqTMQK6maF/1Z0iP94uRO8lewuN3WyYMJYDu
3K8AJgGKblpXwfLgR3X2vqofgzFYk9o9XBPez411JjByWCWktLc1zyGdfsZag7iJ
z55pD0IJMJ3sEGKm+mQx084/YluPcS+RnJjGxdBYUnUTO8ijk3ZQy+ynHLEA+V/w
3pCA7/A86N75AzM3u9Nh8TFB2xH4FeRIH0Sx7sSTVDCZm7d5ssQetXezpwZE0ESt
IASe9IY5TdcWo5aAUaBK9JYf1WKYgzmM3NYFSI2Rc22396uH9tdaK83hhXl0aZrn
lKfGEWe66unVecYEhXdl7SRc5qtNgf+vyZmcsBZpOaHsWBhcrP47xd/uLresyIam
Nf4tt3GuwtTHc+YP9aMMWeep3lldNCDznEx510lxd0cornCCSsB0n1VIbPp9bAmz
HNacmFKNAUvx2y6rEaZ8NJRfuGTryPB6OYYeSO+rhdvDhhDO0DX8Y4O0wTRvc37+
VjseQfDS0Rz5Ep9iN4NJuYWtX2Z24bRaZoXUTZJFGmgz82vM/ysGwkmdfmlN7gn+
+BVFHs8cUGShMHh1JEZcQ1PlJEvpj1lkOD4NaCI6vkjqKFD4mwuYEgV/byisy7tZ
2sGiU4ponN5SXcNwJySyuERfgRlLa24Cix2FfApbbvc74Fuf9CbhJBFuTOiHujGt
kxFoZjIbprkISaFLd3uNUNkF9oOHJQAetXh13UuEGTg8d0rFRgrRQHOTp99ibS01
a8obSgHikSdGIMgRJfbdeq+QUjrmEJYbX7wYt1KSuX91k5xx2ydqfnvH0ae32MzE
xb2tPHzZ5XziaGmRiEfns1TEzAsFQ+l5T7FevRK9yh9xSR72dLKRLXN2WuNgRcF2
7X7ediMpSUnA/iutbeI4SDhfTTi2lfaRO72eo3vRvi/nd4kGBG3gTeTJ4a8Wx2Ky
27idgKzOV4vBB/3oweglNOHnVAdoAvs5CwELNrI06dKIe6t5T+L+Upt/cDdpNpMq
89tN8tuCPcD6xQzEqkW7Qng7KWOv2R6aH/UlDDP4iCWLk1w3lx5tAhcps3mi/zCk
8Y97Sx7wFQxsRzQJONn1gWgi1tIg85qm8ecTZZDF6va3gvxtPkeDeYeegj+Yda+h
aOaaFQC9wJpCOydWCcMkD2BxyYhyB98hERyoLY9qup5XQIkR0qPRctnIUTKErdgy
mkg7P8IR8scRv1ST7+Pkx9UrSQ6FOSfgLkHBz18ReV/59O+oLSS/fKSjo39vTd1V
++4KuDfP3i+/wOORA1nv28IfYwaZNEo7sUk4YPf2Ky5ZHhaTOBndjFbcLTtZS0SI
qn/v77onlM1c9KlG3QX+mk3PswbdpcasHIDDnOU/TFGpP1X0yGI7zUIxemuXN+z9
ulofoRaY52jTjw6Yqz2SM4UKp9esz7NT6GFF8VzRzwuKuad/7eD93YZZVM2ZAIkb
UR+W3CIm9VH7kLd2rk0acj77eMpb0cNbLkJMF5md3LrmcV8A0Cs0ORfuxpebvtX0
29hduMRbpho3xOSxqr5irmJdYMYM8DkVOvPTiyDmtIALqI0c20QrQ2x6qzzvyeIy
6jzJHYBII1gHzKp8xkzUcWUXqgaNIcQF2cvKaaKgV6PUan61xXJM3GqH0g1NSpDp
fbrjKIZja/kCVCzZC6arC/yvpaI3VVlFD+WBJE9c16wax/o+O9GwR/tbAqFfpi2U
9TDk69tCJXxeV4/BDyIximZjdDNg5eEYMEGv0E1RodbTqUkd7EAtvTUuaDjoWe3Q
YteJTzAPMBuT2e9jnsMZlOSCbphIgFdbc/G1zJuBRav/O2fo7+VDGBCZFriGOG1J
GKlJaX5+AtACcM0BS7FzFXLXejz6eGU8b7kTtEb1GgLlj42ZFyax9XUPgAou0YDK
QWBhs80IV6ouroQL2BGCad9IVFXzMgM4S1DVsiqvQkbj5wmcomsVzieoHAlq6wRO
AezghQazr6Y5NR3sR6bHE9JQPWQ/TbMzHJI19o9Q7669olDZhC46/CHwFuvXZtic
hhNVfHgv+l4JROjy8bF1O1xLhICjhGBXf4PtG6ms9rF3vfjFDu0z2wtCNQ2BHb6O
7Zc00v7CyrlAX/eVS6kGZdi4xpgexRqfNQ2DH3PhSe/pZZ2C69iMTAp9n80BRfcp
82LDPQOmI8cvuMjarPI4Wp6Ojzr3EpVqrRgTuACsLxIO1FhI3m+1d8EYHAXtGc0f
c+fARcCQWp5yfVGrNwPrS9ztCEGjPmyUHFDkDwFdy2G0sIcinakCkqJCbUs3ST4S
i4ibE53uRpb/ThtebIkihx5Dz97E2CB/OOb04j900182eSXPv3IhVpuYCuTHWorv
ZsghHtS8r8A4mVn3CaRjYwvfMpqp2krAKnw77OyzpUONQUzJPfIpsfGPT9bygWFm
Gr5ACiE9j91p+ATx+gwB/cetRXMHqxBea+LTfTRb71/jK6PTB3bz0kSl7UVRQzGT
ZryeKdazdrvCgt67nQKdwYKCturMp2ZCoRuGssoIohzeRd8BP2yEIPJ+KhHHtQIZ
eMizn3/3PlAzmdMMEo8qlIWLPZGtsrJIGpspoLnGYoyDC6i1QH8GmpjiumxpjK7G
bRbpwyFBNrUYgFGH4I3MdYLyj1tI16+IHjQkeVqaIBeEB8E43zoDQCRQavf/NKtH
CT0lCs4ETBhTdi9lPPid2GMnM6jm3OPSKEM/ktnQD7WF55VkXlqO3ba+rZSkkpzS
6s3NsWER+txlDQFvaLjjrDVuDSu7NOA0xDy4wyVZggQC22SvlQIdX7zEtVg7pBMc
k1uzzp+m9RKK7RiFPfewgm2WlRjcF5fO1FVrv6UrAghZHpLPpjtghjjVe2Q4gByM
M9Zq5FiyDOV71cPp5nB9jnjdSgLSejr97+C0Ya8EQUcLtYw42Ij14g5RApqbF277
N/ea0/mpQ3pAYw5SbR3HH48+fvYZmIkvxrxjJPlxLXfkR+Hg6LB3DRoMTYdSzF8U
3wZHRhfC1AUHHTHrRWjpDJUt3GRguId/K/F8EJtgi/80e20JXab+uE+DiYdzpaul
4trDTL7sSpZUsibUwQCxuouHrhAoWnW+oDLGMb+JZ7h+iy6BOIyeCJAimjE9m43J
7fEV3a0nxYjslYVL08KVoliMw+QYiJSYCp8PxNaUy6tu+MuY4NkXOPwHpPYHmTO+
kl7HH8yCmL15J4I1ADS4kGJrbsUwlLbVKChrR6AdUwoiGCDcUtRa69uPevP1KKTr
6hBCBUvVrSwxnC215TZ39qXRUu/hmWABXIbeY9kv42rhZrBqhPHnBa5+QVnKNTfR
geyY6LWmdOcleYKD3hIga0CrDNwvixrC8zAS0wNS9GZwY0uVwSzN4EGWvmNFjU8M
yh1alzTWr0wN7SocZ+1O2Q==
`protect END_PROTECTED
