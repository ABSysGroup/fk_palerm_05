`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D5i/u5vW5sjwcDQjM1HeioaNBno2YUkGvCB3LsyADZ8B+z2Algni3qASsRa7FZXM
fGmfGFwpKHxKiJyGJh6sRQ1gDFY8ELhPRxzIZjN6h0GremBwjLTvg7v/SVY0asjg
iQWGjDBDedLgfvgNsILX2Fr3TEnI4tSbuHEdba1zOx2C0sKF9lJWIGI+pdFJRWDy
3rheR3ll7b/v/Vr3pBHCy40vWuttQ4Es6akfRnoxB3/7qlg/8c7uGM2UpTTyOyXs
bOGzx4fCtMosuGjvBBbSx4/mXGvQtMuKv0aFrdK5Bq8bw6x4Mjc+4uXTkZHXgJFf
jNX884JlNQfG+JQIbIWySpWEdok1oEydulzc3v3Zzq6mgu9xRlS22IkgtwZkDx1t
1tp9gTtt0mC45gp8hn1IqPkHTwK+WCetJOxA0NGkvcKA1WA17XJp/LcMpdsoBpO3
/T5rFUhZRcg1AQuhzkpw9j3oD5h595QXEzOss+/jKIdLT8A+Iqmp3pzwZpVmUJl1
eKuQLus0HWqD7kQfVPHgqF/AGvedQgkSo5g9wG+iJIXvQM0X/gaG81jeMbS47wtI
CedvGHjSCtb455dyAIspjZxrAlJW3667lLdC7umClIU30PEAwqXX7B6w16X0mqOw
Yz7pd/lsE0+RCFCcK5e/C5d0KeH6fUlJRSic/e1NU1kIlWfq/iQ4LZNlueA2Tx/f
fhvh17h5j+zJSoL87kkB6p2y6146518RGY9OCJAG10Siq+XCdf++qLIleajv3oXZ
6+tUJTVLkVVt20Mp1cfybObd2MnDcT16J2W8lW4v8wqenv47LxKFeDMsXI+SfmG7
X4hp/3dF6EnsiHDdupQIdTZT4lzlY2TzLjYV/G/JN19dzxB/u3RatlztG9y0EgD/
61tnG96K3Xz0WasPxr4XggOyRwT3sB5M1wS+MJ2mziGwAvog6O+Syzrig+CT8bmh
W8gEKmQ3UbBtTMx3bTwmSQ==
`protect END_PROTECTED
