`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bi6VPa+rR3hUI29UTlq/XnXb9onY1rChfnHFDeuSNeuuLYjHwA0U2ph9UGYNAu8R
WuiP+pNJ33FHGmQhwG9n1izyNNaY1GvW+Eu8Ai5XACHwHauFNFIW+I4vBrgU4q9n
U0jmxSigRpQ13tSnIOucLKEPpM8XkGe74a0u4ep1RMeZVkT0zWrnMNf3Vr8kh8Yk
A+W0i/291w77j/fGllXJ0mTmkDdIhjNvE/WbSiXMz/58lLYZQYIzsR6rozxZrhFX
hdwKfbqSVdCjvC10o5z1y9wxpzpF5tL+JeGsodqyWEB6JTm4f7mpPn/TVn+bcdfI
P5wH0SWJdD/L5pGnakvmUoxsAuNsJ3UIL/1x4NyVAcjTOvyyuqCxfc0+4eqFIRls
5+Yvtc/2+/QFw6jN+KNC5s7p14mQwl86f2tEuZ8GGcQ=
`protect END_PROTECTED
