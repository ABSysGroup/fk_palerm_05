`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
epWNaOsor3k5VssZenUXBAhAqXSOiIB8KppIOENwJYCE4wC+Nhz4cMO1hHNr9A/E
ZWrGYv9fQh8EF9j0zJxAD0j0g13vuU2kuAP5VU1s+Zjr6h2jmHoyWe3EhqwYdbLV
XqCAwNNa9GqbocRG4pM163poOo6E93yd3lqaKExT+y0ICjIlQXEIS2Cogx4vgcAI
1c5Qm2aZYJ6Copp8PpcE26FEooDpnxoLVBV5sFBj8C9S3ea2Q4LxhlduI3KXluD8
7d7f5FMdX1yM1/IAmYxVGGg12NjWgNxPf+BfkCWymt/O5Z+g/kgjhWrVgVmCBufT
wA9V8/b6ok3TobKqd45uqaERi5DB1L/I02HYzkTjq3u6ATcSmX952kbZjsEfG5ND
LnGkdJrzz1MN0tsxfVy9NBitbdEsa35JZc7aoLejOwtf1LXNKoIH/ITeyJm+HBeo
Rwk6QdF8kmRoQy4hys8PfLGxoDuxxprXiGotLTgOwPI+70h1xVa3aDRChgNyXZs6
HSCtTKMTMm7sbABcrUI4h6dm42yTFqctcxNLMwfVmgG7cdr/8FsrdwZjxdL3Wqgk
0tRbV4DfQQxQx3H57D/v3Y4wP+03lOEjhlm0UpovcwhProtCgAtzGjTTUODqY41o
t+lsb19QWnUIhLe6SOL1UeNekiJk29L0yQsUORJbxjdGg5Yw9m9+vFwLd3b+t6Wt
qG5Aw1e2ARERzaLAf4OcJ/Y0TdkwFTTJ8D3oAmQWTneEDjOX5tCNq1EiM+msAIpE
NuIvUsN5q1OhfLJmW+CfBMwevO2fp19sw8/9v9tey5EWYyUwLL+HfimyFCo43D6N
qtLjUPTanVm2Un1BxtnwmR9Qy3ECg7e76FMwlVevXwI3LGnZDthH/KqgT9qYUDLt
tkKcmlJ+KKPFqJUzYFCUt8SIWcnf3d6VJl6o4xpJDncYofI3jonUn/hEDVN+Nbhh
WPnCHp/Hs12mbgw+FL5nHvkrx8nxjQHgdJDpxytvnbxGoMX5+VJw1UXqVgntb6ch
/TGiqZvCd+3cQEAz1v63kCyDWXr1IeUkvgLV6eDlKfc=
`protect END_PROTECTED
