`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZXEc1JC5xACFpQVaRqrOYjIqmtOkTFMsgi5NSBOsBDflBwGdXD1Ifb+EYFOFqQ2n
15qwbNrQxWf5FKvpcrg+X4O1J6gy5Ho5pwFJVCjzOI6SKFXx9jym3BlSHpDFjIBz
notpawgV8hp2SuhmWEXUVXVYeQAvAYHrTXlUHRc193Q+IVQTo0I5wrbqXj3CoLjc
KdilF66WJyyOp3rO9gQIVXWJAROaUnrdKtRJ/4hRdkRMRdXPIGJnapiPwsktw3Ir
9ANRvDTk32Be6Y/mzM7fUfRjqS6tReSjLrAF7h0dLDUsSgvHTd1yVvR3IYON/Szj
lKWHTSIgO5rSig6bpSMzh5KlCwo34V5alVCe+ia/yNuxZ0OmSqcZlSgKxhzsIMm3
MyDLSxhyND2e6luIjiL8kZ/v5yeKVT1IhNqNk4vSQP0zm4UCq54EC/e5HBM8EEdg
BgDyEjUDCLbxWP7dLqw/GrVZ20hejp9XPKc0RpBNgFwPO3Zpz/ZzTbXQ0/1Nwhlm
Cnr+xs0JnjhTgDwL1ODdL/G8NTYaUe/3GC1IdRX5rqhRlajhLOuawTtppwgB8Pbg
xGfV59IlaGK8fBh1inmtT3diljXPx8ds2vb9J6f29FeK0oHuauPlTXdeWDe88VFi
w3QMe8KzLtP3dg7XsNsU1j64qgwRa2J3TSsOo/jMZAMjnlqfvQjcanEdya3MGjEV
V4Ms72N2QO9H/PzTXmhsu1e0ui5NL7pZtFmm/Y3X4Y22cub9sUJCDNp0fUNVBFz9
jnzQd3b3jxG4HsU+ykSVTE6+C7/ju+Tuz/FIKvC/e0ZdS1+CUNWEyA2h2hCdTwAx
NDVSeVBmCTYpeDV3DukGyjLwE+X6PWpJMdP2bY8rhuSODpZXvasikKwenIKbN8Dh
8qcwMXhAp6nvdi2zPwTSED9/HIRyfZvvetukuUcbTNQLF7+gptXPXmyYHjD9U6C9
UzmtDG/oQ5yO8FfucxqKXHVpFfxh3s8gnGsY6AWbKaJy8+Am6fSRCcEntxqtxFH+
4vLPbrIM3IlkdxUM28lSeTYVBcBXUNIJeO5CX8GVIIR1Oipsqw7NqiupaWv12ZgU
OQukLmNqyYUZD9pb3L1GRujpa5h0uzDYkGM4Udl6ZVTphgD77YGYzGHwIvXEWxcc
Jd3lv9vzQXbJ+meAkIQFnx9CnU/bH5bgW/h+wnDxA6/jCV9uyjZmGHs2SeyPDDP+
xVO81SvHZ6xDtiEXwoYyYLUWfc0QOdvtDK2+ncHMVf+M9/4fKAMvcYc8IjRMDGH/
spRKU/Hz3UqNMmM81EzPLEkCcaTGzjF2/3VbOYFvI3DuS2MtqnK62rKHB71dWDzH
hwB4Uyw+pbJwHQDhmYcI5LwQrRaB2PitpO5YoGPtJPUIeVQtrhpCPgK49RRzALAS
muRKPhmq9NpzE305Zkm50PSqo2kfAV9nNccPGIS8V7Pe3hBlM3YVveIxpZMAdneh
t09SJq7ISFqBQwT7w6U7+10BXE25q+2yjhzj/VcSvDTJz7J/Dgq2HSsun1BzXYRU
GRnq/i2c+Nk4Pxz60OIE1gcxPcSxnkSJVnephD4YqzYKt3HTC8tWfdEwY9uUdE7m
s07IKsFarBpIjiDIK5qn4VFI8spBwmkX9Dk7YEB9CbBGSlLD1DmZ731KWefTbzcm
a1QL/06boR0UOl4kHT6dq6ZK7bVdrucUTY8HKVstSUG/fAJq2bTln0LA4bokQrih
/4F4VnFY4NSSctx2bu8EKfHEZENoO4o8TB18uciSNf3uwgl2N2bT3r8enqd+mwdz
OUuHb/XUqtLXf6KXiwGSdEn4l61Z8zWFGKhQVQod4cOINKAcUp1I06g1izG3RHdA
JNP5kRpM/oPK0DAnm9EBsJj5Fm6FmX7IBZq/fVwXrPUDWNo4wEzj5eI5WB42JFVC
xw2xY/YwBxm33GawfRNF0pOYlfXIzsdlKR4ext1HqHRGNkybCwHLfn9OJFr0Anjp
aAkf8i5SKew+5xnq3ULsaZSi+8lyAwBv75nPu70+nVJ1AIL6HdXXLZqJUWFGiYoi
xIjqAupMVA/BDrlfl3MUBso6ayMrNSpgpjjzs31+xOQuV0LZ2KCs3sCXZgGxmvpQ
sQrLWW076WDO0ScGu7WUbMAi5SR/GVnr7yJjEI27VSn6wUNtSYjUEQ2IU8FZimwB
d/WKFXNKNLZnJ+sFQCrd7tqZaFxsRVvxKZ83uhvIFPFhzeekwE9Nc7zSdK5RoknR
rksPUoqRt9l+tpbr0uZtZM2jq9PfjFoBebwPsEoAkoxqLhlIvuVFNF7rmzN34mwW
yKF/+f8TIcdTGvpjnh5iAtAocKM4nQGfy1VARO5erFbT8Lv3bYRx7RoQ26FRiRfu
fkjXR7bfhryA/l0vxVtAjP8kmmpcjJHlktjwYt4tQng52C0QhGAAfbZM8PwRJRTu
Qey56wVOjeZc6l4umYebhNz5VWemR8RCYhZyLufy8SQuHFgmz6kskZqGfetWrIXA
9QWPRb18lvZCr72NEw5Fu+thxFKWcp34yZarq9UUcDBamowVGzHyFs+B/FSEAdFX
ykrwxOC7zznSGSV+80QTjRmSkBR7HaoNpByxa+UETt6VtiVM2OR1+J6Q+nvMnADc
TnhSfcxHssKOBqwCmHbktY+xiwISXUsgiTfrEOGXcSiLgSUWIHYcGX6HgvTGeg2w
ZXTCNtmWisI4qjpxqf7QzU8Mt+/rkomlFtWHfEt1c6hVk+H4aHzMTrkdhguVNyVF
glgtLeYHMrauDF/BEDsCajrVPtGtPBpb16f4du9Pdha8rTjQuNiH/pCfnWMT2ta2
2SrqaitsOfgsxpP+TS3sCIcv8PiG3ybWR0xEKyRCtxjlFluUAXDD+5dIIB9GI7yq
VOMipHakuR1vhn2nAdiBa7ZrCmsm6otTuM1TZuYnCo6LIUnYQNCGY6+Y5jCYysjH
mfZwOB2optAIwFLa0FT+E091u2zuy3DqiT1guaAzm65zhLwxJkjImD/GpGkm7KZJ
cTobpcA0VXlmu2evi5QoaVQ6/DgQ1ECxhVATw9zQA6Xd02w+R16AoCLTBneKBeDM
PRn8Ijt407T0GwrojcINazKQhj28RFsGg0tEjoEvW1ynYTAXhPSDI5uRB3kZXrRP
NfJbu9W7tAcHZGuxlB1lACoQvR1WDKTEV0gqeWuUOQC6hX+kQ9GvJfCudxxRQaP3
nZZ9Hf253e0fJRWkVY0+MKJhnRfZVwhYmEoPYmsQlg9UX00y92Y33qYViTt9z36q
N6VHM/k3fqmiXDO+yIFWW5LAH6KKzxSveCU4RncPaaLkGkWGPl89Jxz6ZMpviiKm
5I4REWfqKLkYTOFHsFBO5cLWxvXBReySGFjGZH5E+uxJbPTkJ8g9EuqAv7HmRGXS
UgB8v5McPGTkdiTQsdPuxh4hNnZCDVfUq92QJ8wHGFhBQ4YHinlbhutO8GpyNtkb
us1unhPb2BoXpZ1QnieK8UmTLryBVppNVKBLemdLxVmH0PmRl3Crojz1ibe362uI
yZz1HFtSiV3sLYNhs4KFZP+8S48B0WUNqzIY5gv5y3IAjdYfY8VNVVZyzVumfQ5k
Vb3VQRq1dlUkgEa2vmbs+sS7Phn+qj5cbU0pPEeC8sMerqt8m/ckNJQ6VJlXgZpO
mvo5ev9bWCOMMGdhyVwR599ioVYxRiPXBIr0YcEb7/25NjYv+CZox91aiDP+O8f1
jrJa/rIG36dE81rhbRVxpxSk6nEbWCaSkh5cPVlFBh1+3OwZuSc0poisinjQKEEU
QgbCYq+HC0atFgLrE0Gh/vvzsWwH0cZ2IVo/43LZaOC+8JvHPdNvIZ8K+DLS+yfR
hPrY9TXp8zsL/9yctevbxnXXIs7fUoqGt3ogWYYTccudJPVDYFyJNN09w5Wlt0gC
K6vGeBc8mWiTpduAFymJYv1Z9UwmD7wpTspYu/0aayudwkkoxDRlJR2niL1m+mTw
AWNvKv8HB80DhzrqNLijCih4XoBrRkTR4IMHlpbPllCYtnROD90UgyARHScHgO90
x20tQa/Abvr76xMOhov4xlqdW+0RNNAhpOyGl9W8Xx348cfIjUXRd3NlgRbrSGAL
KKfIuoIYHTb0TpXFmmzxQRFatzkGF0gBX20H573m0Ne9sCM8hZOXfIqPEgUQK33B
f3EQMQze6inyeLxkrv4SurXf2V7svWn5YwL+U7TsUmAsKps0NY8gst+SI2zSFiU6
Y2dVH5shPI55OSspGSv5hE214fujWHNeZIid4qcevWlDo8iTDUMPfSEi211DmiqO
dkR6z4urqWJFWUx4DyZYHhVuOSuGkkenmyAahGHvQH4EyIygMgMlA6voSY0bk9Er
m5u5BMQI3gVz4xVhuS4fXxQjrcEQwH0BsO12wUosddV0fHDoBRrBAdTlyZIv1ox5
hc3e8XEHFieMnqgDVYtYk+o7s3JA7NHhGO1yoLxe9AOZN/4pZ7YeMzA0wPXISHia
jiCJ2lZdwyIzVeKqRbn158mPUg2XQPYCu/DqbRxersh2ZkKexCN6IZc439vndcYz
FIUpy+sWmvkED3ZUeV0vTY1zxAMtcKWyENMXlaxr4llKGEzqZ1dgjlinYL6PsXQZ
P2ERVi9JaBY6VyDfor90PyDSkVve29Ddn4BY/5cd2WDfnRJvQu700je5CWytb7Wk
gubqQh7rurkyOlPmNmz3eHaoYVcHOFZTjy4ihI3ubxxRfiXdnAjulrAhA8S9wHKg
5nQVv8eQtMZYaKnjo7orotbjheWliJXf/Do1v387oZIp9tSubzQ8UotgoiMM2NU1
9lSarv2qz8n9f1J6bp5YXpVhlGq9VIWOSvg/uiswau7C13e5g46BIuj37R9AStwE
3L1Gi61249xeWzGhhn5ECr6gFGiIwNQkPq8CS5gWEq7wYn8HS8tIw8WxlH8XGyqU
BQZKessy+KOZhsdKpBYwyrKv9aF04alLmSJKbIqrscC7V44WdCanrcsi3AdfLXTU
mCFFg9l5yOi4VJAYbxS7y44FTVpqb3EGF3GkXDRosRUeTU6kSOMvbEK8LebF8yIP
87ggDugeSn/yGYEcWBim9yWiQsyOLUD0dZkjKxAFuYA5Th7AZJZbb3n5oFgXw/uM
Mk16Gh3Ko6dwPPXdjIYngxX1unwLQGzjVJlwFILX6vjml2XeNbOuVVJfTAh61IRm
MKOb76MAxokLsyWpkFV7MgAs68NyU7j3MADyL9t4OrpIwnFlv21CNO3wGUDzQoUN
NP7YwHSHHQzOjDqHal0xi/hO54IMp+4+6zpT7mNfaYqElPHZdpBw76bn9qJJ809N
T6kYMClMNwtwK+ZayssVabDuNJz4BVNKZMAcA/b1YXYAcct3OaLjuqU88D6MOLXC
Due4kQ7aoSXcrzfddNoldBrwEAZT4UWXf8ShSgBGL5L82zCFdLCzNevRkZJI4T3m
spB6/QVekrKxTeBmes9sHTqV8GABrsr84ZK/hHwWkxFfy4xvlowRaFYykZBQhs30
40DvCEAIoJFc+j0WAPlrsMF2Shl7Peq0cJ5haovf5KVxsRTBDNrsp3lvxWsV6uv2
KmfdpcS8Nf6ouQThvvKs4v5rsEwXM7zGYKH7v2I+jfrPyX2CgBq3Gz1gtBEepkgn
B+NIX1RpvzTSZlaK8MLlAd0/80RE9UV+a0YDlRaTGddOwJj0l8lDrpKU3SpXtnNy
Yd+UtYb6e3e8FlQfTlCswfQGhvgL3UF29TnAhBVZ7Lx7EL7ajXhli4ueI3gzucGC
VbY5YEyuEHGvrgkIFrcg3hrVWvBBCOD8popfYohkvuUn4iaeYKh/nXJ0GeLIupDJ
Nv7G1Ta6L233wVuU30wQIB2c2mVm786GvTxNIBqIjWQSyE1ZnZ8SeAUnXOKdVAKr
ZpjqHgXWlpCVDVHW2eq0iCPIo7FAQwrdV1l4pGeKDrUR6R5TNccDiLy9sbNLroVZ
XSL0ydbfGvWNb7wgznqzf9f9vL/m6bKH6Uk+X+CvYtkpEw/qBd4tMM90Ua2/JQBT
ABEQgfhQ0TulU17BNHQL+/U6A9V++u0fIhHt+/nJkdCkNqx9JA7yFS0W/6rtl1dN
PXwwSaxOmmdx6AQoRleIJJvRvalep2vK/frXy5BNX15TOToAjt+0ZvWeZmoLrwjY
CG5oZOlPBIGNcCZjUrwTWZKx7hO1T6HQVlGGMNSVuK1MQ3S0D2i0h8Hjjn0ytm1O
kKG+oXJKcTFDSlYlnF8YhwofdiSe6RjmlcONOsvorH+vw1I2ONjplxDuyUE3xaZc
xv+5sLVgRIX9xSPLkb266xP9iFb7sTJ/fZFt8oV8tsOyh/kbZNYN2l/aMrtZ1BWC
m1y/toqFPoZvzA4X7FQDeAhY8kryGCma2X8YYBRW8/aSmzhgXc6TWAuyrK+42e8n
yMptMaqZi0Qp44p2NnKpaKDIY5UW4QSqAJboTGy3AiuuBTqkqOFtXcM570qP4NnS
+baBfTLuEhd4xznGYyo6qTVfLJk3/KF8JVFx0JXxnBOMM2zg8/dpCRRXsjnWVmCi
DZfzw8zq9JokhRNJILREghZpkUT+HTp2tY2gqooqQQXR16mw2DqvZdSBLa84Feq6
YKjvRtjzTdVcT5b3/7Fk7Ol2Z3sjPpgBMe/Cez3xOInJ6871xDcozT7ztjSEOL+C
ey5fC76uQuIdsPdtZzAGvz3FZPLc2j8cYCifqQLoEJ55bYn0PxBIIFheHyQQKkCf
T2ZpRQWn8OTIAl5Bhq/uBGaTml4G+Kt2lR5zgBkixG1J7Z9Z6msmM4TgThV7dsg1
Bp/VgIRegkVbW/XXYM9Og3n4iOK8H4We/DQ6WJExk7ky/+WBdOF8Aslo4o29eFU2
CJVIVSAEWpYFmkiyZBfC5zxZI6/+0DYNn6RPIN2aA8SNiy2K0CfO0q2noswmNbQ2
99I7qPxKpr3zUaKDesmJeqrmvggUpSR4DUL90/hIz2ISdhxbmsmFrzb18257Ak63
turoXfrvYXaoygQQZv+ozSZXkn2gWZhC/qmY3KrkVe4CoH0AbSDgw7Nj0bXFRhaY
HEWxd8w0AH2YYrzdE+GEq2KshRy383ZBjs5qKXUEbfbWQEG3QvnX7eGgXSluohtw
hB8lMc44osaRUfETdyUrauPbUpaSWJ4fPl/h/fFmsDxwxt5+rD9dv4tduS4DtpVN
6nBJqhVPRnrKqIXeRF7zackE5hTP9MsSZAtv8Lac1IuUMA4ByFArHeoG00vruQuG
KwYWzgFnPNPjZ6FH3uih4/DZIKM5qbuwrNsoUB7wtf9W9GJfJV7f6OgRi3pfZVvj
yGwfbQqYuhj0tIIjd/ubBhcl/it3jNgaOklfEVXI046bs5i4Db76KL7CbH5eAR+a
ENmSv4Q+/zROTRPBARCxkg/yPi8Ivvb6qcy9IUxJzo415r5CCLPJlJr2ZKAnLvUB
TNSAgnjId5baoez+B7IihneK11+jnAVHM5eIP5tTnVV/TnCy6SQBcD0piT7onWKW
JHl9nyTDBKhhy0w6UppwlI0yotN6XTM5sm4jyvuO/Bj3gbLzxkC1hT8N4i/lqrW2
Fu8+xeY11QVLeIsHEkemClnGkl2v3qTjE1RiEKSVG7jx5bdc63h5i6bUWgiP2EPH
+ltrUO1VmhJ57ICMsOwzueA/bjwo2wdVXqUVWCCbl41WD+NHLMKhZ0MXeooydbHG
sD+rGQ5I5kfnEI0P0LyqZfubN6c85J56a4JBfN1FezPSavoWeqgtuAyqBHLYxewS
INS1I7asjjpaqUDRDVSFutk2VvytXCgc/opW0hwENLfOvpOJpkfZe5w66DjeGiHH
Nxv8b1KJu/kJiwU0UHs2Tvot4t4SNWCKX1jI6oESnQ7kCPrIzR2ywaFki/qiwoRr
uSleqk4wYyiMJ+4uLkoKpkANcBJQnCYFLFpP7w2UmEUJQvDUiy0Urijm6pP+orsT
Gh96xrlW1kmIRwZ1hzxV80SgActWYXMdpn/9etebkhjC9ZPyCUoore0zxwd9xAcO
UVaJ4lZkgmq2xgfyyvgirqJ4h/ix82KrN6pDu84GxnijkQy/FKXygFJK7A6BTGmU
LmHuc0RylJ7aQUU9qAtE9uvEcnGUVaxqNbk1gjB4MJI8vaL1phqKdkjf1sC46kph
MnID723HStYgQbBRxZdCyBFUJFU3Zb4NotdUECyVUOhUUfZrIsHyG05xGmdJFLS1
6wd1ixl6u7e922R79rwsKIf6K+6g06S0V4MeCiD/I3+5w7AEaKYpXvPqgqsmVy/H
kTiZ6IekAo06JEW0GY0b33mbBW5eSxky6K72iTU3RudDPkRCAOGTBU0EshTE2cot
O9GFzJ5uHFfejMw/OpxEo3VGjuXOe/UBta5b2rxdt+TMRTV8cmrUP5ioLC8bNCx0
RPESrYHI9SVqSn4S9bNLceNfR+7vl57xRW1me5AbR4xi2UDwbX+sYi7uD7aGfDvR
jz+27+r17jc7v0o7kVsbi01I8hK60dnOBa2ttnEidbpMpYjYJDzJeYNhLw5D7oCL
6ushQPP1sIe/22HpZnfrRWXnSpNLkG7m1qlYLOL9OOqYTNoYy7NmUqq+7zwFE7hO
7R4lGRJ/+ZPBM428hXLyLeVskP5yG//IOrcuvcd66DrNZzw0zOsSUErwb3d/9Ivu
FAERXkB4gawBeeq3wrLRkwBOxi/0pDZ6T3IFjEweysVgebmR5qFRdg75M7o/XLcG
d8bSv8Zh5qO674FH55owZ+AMx3NtHYa4HVo17t70X+0Ops3CUGJYUZAmytB4MHU0
WAqwk5OOU92RTfBeON1+u6f9x5KrDZVgdu7L5T/DsDt9e8lkxWdm0aAP0lnPlHTI
2DpbnxiZG1VGxkGufNxRKWdBfJ8YAYkbO+k6Z1nHtuDIUfBUh+CQns3AYMW2L5wY
sgcQIhtC9ODwDAynNdELiXUbu++04Ljm/BXDB2gqPjgDguBCMAob3Piy6DtAMZoH
fSWQRncrS4O1gcbvbqo9atx4pQeP+m/XyBckH58gHTS651X6peoBDu/Br/4KV/29
S9jf3aLrEbs19NW4nmtzn2/1JhGSFARBK5G4GnLjo4KsSzrFJfh8ZcsNmxgUvfGZ
zQj6WDG4q2/1Vt8GafuhYw8IKzVA3mo/PSr+XiUPc9lybtGzKxuCrsKtikYNJVIq
QAqPUJuisFtm82vlpsPes6ieAodVpWkxfxVKgdfr/Ft90JjYq2eTR8LLqgIiBbOW
ypaCwfLs7sJy83GfsyAkVe5HLujCe4QlDR6YvBxO+f2MMLuLWg8K5bpD73jAQRUD
Flf9mAX2u/AicEB3zJP6LejsVeeQtTCoKH02hZsG6h75VordjYhR8BARXwUaCkKK
Xuti6k1UWWUciGrCFqW9EwA2FEq/OX+pKwoHQmW2qLItn6CUAN/E22zSk8dO0178
6XP7NrX65639Spdl05+dRLUcIh8A7SRX8w0w5H0dtsTd5vMEvWn82tA3MW2i/h0X
gmGL8hRSKWHF5PLYuh+HyPXDb46wkv6vyp/jpa32JwL/BgwX8FFEe+02taX6+kGW
X86Ms5ICMOGoZ1tMWTy5D4xTIXmtgXzz2/Hk9ReLxTYYx0i/8K9RKaqBA+9A0Lfd
tENRkVAQ5Dc0vl1U+XNwAqA15JIoNtROv3juVYBL0hhvHxUvO1GJUlS+HEyzdK1F
noalhtJgxtN/79v9sSEmJRC2fFzQ22fY+dh7xORwt+jyxwTAm5oQ9D27IULvUrFL
QhbmEcqLQbtCiaOiC0HEkQFF1QRYtWABeHFwjJiC1UCpILwgD/H1WHqlqcs2eJMs
BWyZnHHA9mOW5STW/AIVz9gmcvum/yauu8nQUxoJ87hzwDZYhTScL6rBb3WGPu8R
CtqdsKu5Nzt3h06ZbaB/9mh10MhjwCmu1KCx0T/5MGNNZAXfP0S3HRJPiMwInwnC
fsuUMEvzEfgP98Tozm/XFzZEDC2WoIOKkodCWtU/urnEPoTzf4/dFtfnQAjaelkq
0dxJtro4qYJGlSPSQ8Cgs1N244hCqC/AddpjkRLRMhXnZ42M5Nf1JF83Pa02uC8K
3apLWQ/Cu9oCH1bu9svz0DsV7ovRbnbv92+SjdIZHw3regd2NSc2YpIwbG5Y+63E
OrcZFca7Zki5lXwuNUIYbEc1AN5slKSVaLMziJtHU6fBtRCRkPO91nYbXmak8ZWw
/2V9dHP3Gn64hUQhb18DM6arbiFCwDywm8Sdy2tjQStvASu8w3giveIMj+/UAqDh
d8UWJaL5pVfJ09UyjT52gQ==
`protect END_PROTECTED
