`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wiJZEhiA0xfdHMgkONz/H/5z2i18g7cd5WWKyfMkxvmBjSCvYw7dZ4VnCXVvgm9A
i8ouaNdHA5FCJ/umbifBnGxG+jp+6u7SuRCTHqz9Kst9W0M/gljyWr1WgYfQfyhZ
qRMB8n0TtS+pmI6zvHT5uNioSVZD0g7CCVjBjYQyaRSAFywSTD8fpLDwQ3P4aYGl
fNgd5SIXu4MnRJWQ/B8r4gl6DsJIWvR+2R0eMRQkl/19og1MUTKZWq+1zmkxrQMD
jirKA5iOvcLshGpQX+8/N6MUVJnCp5yn0y7heDjj73HmzSanqF+MRtruRY4KwOSz
YRuDdD9XZYHJxK3VKVGJrP0TTZ1wIjGAkgDIKOJXEcWMAfE8QBud9RiOBxl68Qyx
IhQPHYgyJpOf7YtyU1/msFkI5ebIjfcSQw/mMIxOq5TUuKuToh+99Ls+O7vAFWun
oTP5/QcippmR5pq+Bl5p7TWyAqKFOTjYiK6NHTtg6Wr09BrhzErV5ExW9IaPFQEZ
268mJ+QHeO9WOOWcItBSRNDpy0QUPJ+Y6JrL+vDCNoN47HpV1HuoqZ/jZwpfDlZ5
9QXcRBQDLZ6ZclxiodBIZt/ZxVDRTnpf4OW11q86CNl0yCG35aI4E/5HU27FHufA
koJAII4VqFnxikE0EgbOSA3iiqIptIqQnb92lIL+Ydgqodu/J/iuC8E29Fmmn3cR
IHNw193+0zCMMPTzgLR5A0nBlxJuhb3ZXXn/izBMrp9fcsHJFz1lAiv50QRKsTSc
OXOck128vF0n4x+Cc3/c980XPRwWfge3SScQ2nlsFU+HLPi/lyspjx2WWj00ZUEm
TxToSqol1Npixmocx82MyZu2v7XUvg5/4HIuLmIp3juZoRxWS+/3VkjFuoSKOK37
Fnbz7QkOuioc5OvW4Q4PqRquX2oYCz01GLO5FBxWoscdkTiMszBms9TdydgoCLpq
/l3Pz6/pFtlQuWx3QWDWRg==
`protect END_PROTECTED
