`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uc9HMahHBfKh3H388Krfb2PraLMrtaOKRW4jqE0w5GQ8/qUYrLDIHe5edryaZ2Nz
4+ZWyR6prxJ55D2zSTDWX+VVchYrt07M0qVefKaAnKfOaJw5fYTtSQYWceuXuDnK
BhdNArXrZMUwwa578xklDd6a+7fqEC6csGAOQgmAw1KKMYJgft6FgOsoykRdmoJN
qjzO2gi4zN51l58FzKl1qLTgzeIUc2OA9YFRnfv+zwgOfPcIs7/VILdSw7QCuJh3
HXMq3RNSyzCRp8CzulBWfPgG+SfhnnJVHEpVt2eXpjE2BAwIE0O6GSeYEpJCvct4
EsAXpGN07FU5XlhhrRq4yoDYh/0+VnBrn2LJ3hGxk5/50OysdZqGK0KrYdc4VLeQ
roMGC8W80jUbUqyRSKlGUvXjOK17HlvSp2EqKGGRZQ8GCmGcQ5ylSnY9ZDAWukQc
s7d9Q6MPMR8hO2AVPbFsFfeC7ZMP5WD22Vpx0PI1+wLxMF+olo1h1NsAZr74I4zc
g26LFQWD0nT+qqGYEteEepas0X7U8U3Nodpje0cqMEceUfpEo92GhW+wSLKDxnDd
cIS2l/8iHWByyyjL8lyXGVqwVgIMfFIuuR0UmLbOQsgljO16EEAIWYQ42v5DTU+d
23Je/cnO0tRowJrZmm+WULPei4EeAXqOL05hwBOzLczO0GqSXOmqu46fuNJYe7SN
pgGxYgtfnUBd7rOkrIDryOPsApv8QNP/9UqIOTkC3fGMwNEvY46tFOquujtMFk6a
wEif0oaNbkkwX8PPuJ5Ljw==
`protect END_PROTECTED
