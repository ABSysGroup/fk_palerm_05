`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r9QUUAm+D+oGFQ2taZlpnHZv7iJcOiXXjRg3C8ElLi+qen/dEtZQcGJfhfMUEvPg
SZVafhSUo3K/e8vVblYW0IFgCSbhlew2gpPTEsdKlbyUK5T8r+48yrjCSq58y2PV
uCPC3eMVP2E4nCr8TzFbB1RtUEbDWoQJ1gvgX/hJMwwhK8b28XPRLR5v6Y02H471
wm2HTBm/Fu3UzsP0KrMzzKAIfrDegUXNJt5vSZ05zKJioIwY5GwEIlq1d13Qs+hc
jjuIjqirpGZkvv+RQarC1V5vi/BFi2Zmisrmc/ZaKeimWI2a/84rHFLGxoyfBkNG
uv0EXsCQrUsugAweh0bmt2yGWGDWihZd77Qlp6ihm/YM5eMQoS9uVtqQ7xOF/z4A
kq35Ojf9VcUdgoJ2C3mgD7gp6Drq71AnqxyRbvNTs4hLe1+Ka1uSAnd6eokHCXGi
7jlywcRFF2mqiGysrxzXYwy4wcI2cbOwrhH+arOqgYWjtWCcd/tJs1kdmxptrPQH
x4hya1k0+X6+B2Suj1v+Yv9wP5GagtUBQp0p9iFcr9LOrr0QX/BGT8Xk9n15pVVj
PAMqQyj3oPEBFm+YbNQGlgdSk4PWGt0ud+BL167jxcAO2udsOpwAoZ54D/NPnJdi
OPxa/sEcw0PUEB+8bOP3B4409X8/XZJbMMl2Ha78pq10innAZVS2lQVmKwGodxU2
LAC3552E4jJu18N0aXQuzGyks1mm6/3lBmo27bODgulu7irjbWfDqiRpYYPJstcu
arV7IE0OVSXKrU5m2v6uXzZ3TZFy9ThAXcSWte6HKOV2Ktu3QV2g7YqR8aDb7lJU
yllWGL8TwKK1BxjxSBEQeJN/04PBwD9mo9Dis5iVbkSJvmR0ooTKRdX0EgIsN0j9
pqQTONN28hXfU22CMUsp6RCt6McaGRxgiPqk6gArBYgNMG31dbCq5aSUI4uAyGGm
ObEFfFoNw+hi2eeT20b0QIo4CUWbJrY8CtMCfUXsnMDdYXdoM9g8ngcBGBO5w2zz
ZMZDW1XrMCWLa5S4HK4T2ZphyfMm/EzCJ15aMQ5DGb8=
`protect END_PROTECTED
