`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jRR5OkWp5r8WqUjdYv6wuSwJrfxDUXq7+OmJXIN92uNT1KNZn7UHY3QA3HlcYTBX
CBozUzowR5zLGxB3H0JMfclDFqXjyPU9f5gSsRZjdMPN3BSU96Ubb3LdP47tT5Nd
0B7mVF98hKXa9i7/6MnLm/hd0d6wfrUXJVjYZ/Kbn+PFjZemAZftqBpnALT7gT3X
njO7MNXkzbnvbB6enrdMFUk4wxYlBPsbNU6mbMaIdSje59Bvf8ncnP/ZxSViquSc
UU6t7wS0ocjD7LYijchLLz6USj2rtLGK4wD/4I2dQslsmeciL8qohxztcUOMFqrr
WyGy0Ebj53iI9iePHTdboRMU8/g7KVIfe0z6x8SwXjE=
`protect END_PROTECTED
