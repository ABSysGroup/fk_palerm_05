`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cgqsygDSw35+Qbe8777J4e2q9+XsWeTSk322gOqwoFtLszaCczrlQVdO3rxJ0qzv
ysiU0XDDsWNrqLkG8i05e907Rn42hLufKIHeXI5c2zne05Vc5WfvHR0MQHxxj+Ud
Gz7GLau2l0HfkVf9HD2ZFa5ek07b8u9IRdG+RpyPF89HExZ3xBZySCJhCMhCgz2/
8+tjWASmObVe9KMnJX6WBEObYKcIKfp25ksdrsCmCiKZwbaGQjM0q468Cmz45ayH
R/xD/Jrh+sh+7qeIKUvV3UE2FUsYlq4LiU9WeyCURwcwHW2k7UmlZdhKjtFyy8fd
r8rbilWTaRT0jOyk7PuAseINwAKP2RATAi+0aNIt0vtmQzfg27y34SxLEjs/mXnW
`protect END_PROTECTED
