`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I6qGb5vf1hn6Srf0m18hKhPKSO7Ubmxp6RQHG72ogpHieG4eIpHyjzZTvsabMrCn
AaQ6RUybtuLdbSEyD0T5/Qxecd2c4XguW2WueKtCEOjQQuDsrFbro6p9OSkEFLPt
1vCUtyhQBiAqunbUt0pWA6RIj/eXcJVuzxEZQ3ulOf+XCux4mwRZjBsKolybuImu
PNrPQFv6WYkWJj4zQ05aSsRIH2F+gG2RGYgE0eMIJPSwV1pYdZZO/EScXGfBM3Ci
In5EI4L0mSBdiNSmwbfeRUxS3/DfIHhkxCk8T59h2+CUFfeHfgCFJy8KNWN5850j
hJXSmVGM9/Nvb5LzHwwxTnblu9TIS8nGgW9DlU+YI76qsnKrJQJpNFFXfRxwxoAm
hhZsAxvK6Bd1HrrjagBU/K0PoMyn9HwFbAJFA00fLsGL9C7YuKSQYKSbSbIfdc55
FPxseAXDzCYmivxVA4wpl5ZYalJYqkZMQDsa4pWw+IGli4Oy3IRfaDjikw6FSGWN
damRY0qT+PQpGDtqvDwE2prUgK+jPddwR5XBl9zC4fnkMCJT9KjBH8D/pwoOPOvo
CjyC2Q91el3LkwG0W8qCDc6rtTFRzQgX5XfRfD/9MvvIqIAQ/DmtPrm0h+xMYBWB
kFUfUlYN5VWP8TF5NOKuoQ==
`protect END_PROTECTED
