`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OBefTAezgcbSHgE0VAvLjizxZ1woVH82Bb4zZhnEqzeAF5JRLFDrILmqc2XA6qvN
+mCBtvnKo2mRKVJKZJYRDYjxrujqrNHXmp1GU+fbL/As2Fl4KgNYVMQjeKxlxy+f
nnIW0CEpPv8HUH3rRD3kGyHCTmNMfNH5mRw16S+Gu28TVnyeJ6tT9y0YS2bKNiH9
PV5/EFsQYSFq38H9fFpP6R1dv0kE1YHVKmw2jUUnakqEynAh0ex4O0W1qJqPi9RW
r//mDG4hnIZMw+ETdI0Mhb7LMhUMViK+PGyh+TwKtbuvsXA6dboSlM6p/cEYP2MS
tnvBJMzygn6ruZ3p3T5mEgNx/KvutDtZKknaa3dgGrjqFfeiq7oaRo9fU56VzAyc
PJV0Qq/Y9lcEj5C9uPgVq4buXRty+t7LajfFyyjF5uPzQJ2ZstPtRqca9KR+pR/Y
y6sUBlYvez1DjM/PzaLiXA==
`protect END_PROTECTED
