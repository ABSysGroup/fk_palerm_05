`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fdkmP3+tYuBYaSFFi1GyDIConHaTAXGhmY1KPrfPtKnJmCwzgeWW36HJeq6kcLne
D3bjW97zduFytcbIeK1QwgyBRQ/jol/zWCGv0jxz9StCM3SrM06nxnvBiZoBGPiI
jSV+5OBx1K/0xCA3Eww+XxOf5J/vTm1sgSXKYvQMI0QaRm/m3EB8CYraSq0UFfRP
evVZRXsxXQReTzXEWyC13zLEBNVHuC48sG7ehjw+clGC9WxGOcMT23xJc/+cmaF8
xEC+oyHO+F0bE9LzIVGY/UFvYXiSeTS0ZNq1iWN+Amycdd6JAe1HIkCMx+pn3Pps
OJwMa0TIgtyY/3igXyWMf63N2rb7ampO8crDah0xA4YUzfV+EqaVRs6KHLorJIGb
oNkSBu/5W1Rgb/VP8mha9Obt0Onzbnqd7F+OvMrw559rbQqgBRy56lTm6ckTCEPV
lBznBJw28IfdQrOBxv2OLel6E/yeyoZfoEscDSnstBkpw8QasmxqNNtAlQ9iMjJn
o5MG8W87BAiw/hFOy8fEtLxuOcaSB6ZV+RTCDGJ06bgwNtMTwhCTBGWCIYEOg9sx
`protect END_PROTECTED
