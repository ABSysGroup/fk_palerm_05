`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0RlzBW2IyaKqDmv1nSY1sxW+xLNS9aAoV9c5UX065wnYMOI0ODYvBaDiKVc1DDEg
80sIWntvC5801mjIGvZsGjM24W10INRbsM2Qn3dWWiPpLJvdCaAxR8YEh3/eoXmF
GYTCiPWnygyjakuir9k/dkPmn9fWTbGrlh2u3FeNyvkbS5bOO1nCp4zTpFSgCXJT
7dZwj4FqpfmlpqIf85a5J9Cnr3Bl7oTIYGRC2B6zOT3v9KtFqGMFM7zXFHavUfnM
3sc39mW61bT7RuHDjf/ZDs2EVzBOBcfUJtVUoMseibeLdLfH7WUmKe4E3jY0S9dh
zMLij/XMMNIepD4oeNlVVhSOPp7InBHqcspwLMwwBuZQ3UVhG3cOvgqtZFhFrTKz
WiTLkhN6zRwEcN3EBBvm9KVdtkyVyebBZTAu1q8XbLY9uBhi0lW1VePNTK2YZo1+
kh37gmAEI1j+lh+18fFMQg==
`protect END_PROTECTED
