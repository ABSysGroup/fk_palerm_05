`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Paf6uo4xE+3T6Nf6H9WQvjwSC636n4zSfHuptQBPGNvQL7jQ47pRFnfzmg0Ic8T
v/rtqmhlpkzyZae+S2E/vUnmNriZq4YeDXo3SE2oSmh2Ss7L5l/1XTWX2z6F+VSh
27snUHxBttEuO0HrK8M/ZVjfG2bVNzm3tk5y0q5RSjNktqmstZbBIe7jVTOWPTSx
0FzUqYOLJkPcD21MGfKVcZBNibycIXpGlMP5/nCMLma18RskCYFzamY3vCJ/Wwe0
a/jvOLBqfBsv+tY+4WQydUiFK6JcRtZi+/mf7vPAvr3aN08iagDQ/o2Wd8rMmBX2
ZeRgxowHowpQhWU+A4wlww9amS4NRYosR87E/zRHm1flv6ljLXS277RXLc56mVvr
ksCHQ6iV2MK2luD2DH5jJr1FxWO01DXVj128Mnji/mfsqXSFeuOydCiSVKWJyktM
JAGBYqqoZxA0fvYUE6iuzhaFT7rhgEyKV7+pjHxr7FhTZntnnv+itQ9QeYBNWxP5
p1t7uoyP84OL/93B1kda7WpTE4O92NJ2pvUsxE2wqsmW5Q9oX4KoTTWonuAeOxh2
un/3g0HAsK1zgMAze4cqRPSS3BADR7SgBQmYuh3LgXJjMyeWOQK28ccrP20wcA8e
96Lz4gOQl7yXIvjL3JCxARyQwv6BsILGezj3nEepLcBhA4/DsjYryDTLOu3r5Mpy
ocLV7oUWrnoFnPvS+xoOrbw6t5Q0ZQlFvIcA8rxvNtaFzsD72BRzrfJhy3a3kFd9
uOov7fBcSd7FYSrCFqvpebPz5dTRKnWARiQMF930bZvlehoIYYk3K2w3jJlxld0r
98vOMG2lz1E7ji+Bs2ChRcY6OV95U8Okq8Ql4+DD14A=
`protect END_PROTECTED
