`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7a4maTiBjaBrZ83HuKTFiFLRYMHUceCQIiiBoKEUcdoQuFrcdUl5Yd1v15SfxFvx
jZ8QzuPtlalrL06wlEuRaAIVYU+W+QYG6pe0OscSigDUOitfviWRisOa2ntJY8uv
XUN1jrmf1ntXlHg4gj2TB0sNm+CZD8srSx3bcxy8Pcf1Mq6kgK4CfsmB0ocT7zdN
cHGHtPq50KPemjjNotZkRmgikUM/7jjHvju9lpNoujvnx5SOFJDF7kqdzwRsm1vJ
aBgH+GXns3eCmIKDGtjNrQtAOYaJgcK9pVTMsIhzMFjcM+pDAX1nbHYB1hnnYh9d
C/ysvGIz9vgZbTEFukGo3ppGfwYg6ushOGqyXra3DbfKDCdQ/pn7so8GfXKHRRN7
`protect END_PROTECTED
