`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3C1QANZKfRy4NBaL7ErMEZle555dGDGWf2EAZ1byB7f/u4ewUJm+V/pWE7VtiFiK
NFpWskCSNXduNMEhwJDBpvJO3HtTr9+jDA/xDtzU39sinuXTRG6s0HdDj6pxAkBg
wrMuVT4zb1MrCG7R43MjCJJPify/AnRiORFMpLFv8TGlW5f2A90smF8awtPQyGE0
xaaHghlwVILJjvx5QD4NZ9Qhgd/aawxyODMrpLZ6UR1Oacs15C5yv9AU91x/hP4t
PvMEjtcBoupk6a50pzonqc8AEcmg5L/+0DybmfhWe6vtrsmaTVBjGfu8qLbkM3fr
QMRW7pWetJZeaONoQivdwV7OzAObmErFJ0y8YEKPkGUKxKAIJz0UDiL21C6osRwQ
JuN8FhJ2b3gAcqbCl8g8fB+IwL/T31Ve6i0UanRHFrwrGX83xb0XP85t5hWvAMb2
FH11FDtJnvI020U/04+L9Rij0pV2nxkhRAQTHlX3UecAGIpBzj3IvHuI6IaJTiVa
3fReYKx1J0RJu8gCjb/SFJq1NL81bYwbeUvfFlqlMxX/jt5UAKqOR7pvps/ii14x
N2lCUAYgOsFJlnUaW0F7r6GCcK/5WpWt+ZjAOZkQnOmr3H5lVw6xZE2Cpp58djs+
ntvSQBUptMWeHpO9FvLK3bTNEAD7ipC7P+a1YgbGN0U=
`protect END_PROTECTED
