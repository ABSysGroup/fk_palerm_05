`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wgu6NswjtPli1utzyM468bY0Q06mmxzcZotKfb/0OUn+yojE+9dlIduZUCvuK8Ox
Va7OkJSZUp8osSK/FqeenPqjP2Q5p5q4K1TsJ5qtDRGQvEPHPmJQERE7V/ZSYjpY
uzpMNG6MCkO7PfnvQIDrKtgRXdh2z8p4hOOPJkDibvWQ3SXouw6pERhoTw9E/Zq1
zuLzCriuT4F9hfBWm45kCDY7yGkjkMaC2Wzf59GeWJWH+Xg3/YSw1UdvlUqo/Kvp
cqIW5RY1DD1jMLodLQEMvEymfKWMQe/wMX2R4GdZOt8d8HQwsc4Us4OQlj+RKBWK
pEAWsNdvLqoGtPabAQABcLfxD4eHkoJ7/Drr7Yz8LMJkSOOWPO6VXSHxFRUfBXml
csdBgh3+h9aCNcRB8To42coxwIVRmLdmsA5+fuX0dzecQAtKcm6O20AYBVwVrJIv
SyfZnZretgQSiTZWt7X5Tr2StwxRODczRiiiMCYqr/eBnC6e521cALlfj8KA1OWZ
JgS2tt8ndAyWe6odJ0K21qCs6uPpz41arCIB5/wbMTHGMHVD8XD+7hsR0+Cq1q8D
`protect END_PROTECTED
