`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+uEOl/kHV5w3CHpMaQR5FJXjelp7YtUmnx1vjLUBj/6XUGI9XVY+W7s0d7hYn2IS
4fHMNVrm5hc3H63dNNECoJMWDRPA4ZenR/8+AtoUG4Esoo8G6hwohMJYb7rFY2pn
anhEGVx3A9CIR8cLg7IfrIsozM6muFu8ADGb/ZqBR2qxmgr9/Ip8+7nqu9QnzwlL
R+i7VUur08RDjIF0ZMCi/7fIrWzoJ8zn42Tu15TlyYg20JhWzqU5TcL29PQUwMoi
cmobi/MnegSl6KMY3WcHFjEJhFqD5olyTFUcwVsseJpli27g4YrThMz+JgTiRHt0
erKOLTcixcC7E+OK4kFMPQgQvN9YaTqc1SihUUacHaf1iQvUSywRJjc/EvlkXaQ2
l18T8fGBY8OD98/Fd9bxycLjpnkkETxxg6Fw2p4rIKKw0CiqkqDHWK+cWie0GH0f
fG2Z5JMC1onXfDuRV/WTH6Yp5N2iSJvNVLNZJ0J+C9hLlhA9KciEXwRn9Lpz78u9
xn/MpzetkvnW+20HlyeTLx7lRTd+84UZP8a8Rn+1UdX+4ANZGZR+o5tLSUMLRqym
tAtisaFM0DDzsB23hSXeqqN/bd6FIY6La1JBg9aetRGTjQRIyX8avCM8K+pXM80R
wlJPI8BsE+V/sA8kGzIfMg==
`protect END_PROTECTED
