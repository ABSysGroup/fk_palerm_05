`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FIIcsZ5BY0r23kvVALwIoYQTL5j6JbHjys73kgX8L3Yrs431XoPl67YCyBq5Pt1O
3/YahxsCMtNn8US8hDvx47BKYXF5BoWJckbVRd/clZfeUuaBM7iM1NPFQdaVg89a
VHpsTR2FaE2ErcnknLKpdJ0S0lwspmeA3pG7XKU34XkLqXVA479jpI/pbOHsZvSD
wYf9ySKCW8n6tFyHbnU89rUjOHnta1AzJPVk2un/sKVY8LB7Wx6TwS8+zvRJu6l2
fCSPtrSghNPMThs5bIX+TPbFCaVdaGwjz3MV9M0VuGS6LHUm/BrK0wzFHuN9SjkX
r5FsLxjX+hrdw1yGwSt9hqDeWk40tL5A8fXmk0xatQxJvdpEpuZIjpWrzO1J6K3E
wpjPt15RPDRnK3X42btATF+OuBTFs54tm7zE6yzd1I/QDA0DTCp4HxUsSyl/gFrQ
7eMDxfUVpQspFbk11BhuDpUq+jNXBOOzMLTFtEC0s3a+4Ncp4rKRWUMAhCNNRnWg
DDwjhGARG5E5zZu08E2Y/gmDh0whNmxJ1FmpRj104hAIgVUS3mfE1lNP+ODs/Z7n
bLpgBHNM3joWenw2+9p1u9l2DOEY2d02gLtFfj2mpGmPm3rahxyikWesLmlM6vPw
tT31iYH9AdTCBro/zyf+pNGYpqrapF7MNNXCNrmgg2o/3mZ1Ayh/Ebf+Z2Y8AQqW
Uxhxfds9vxKBcirtziQE4HvF27jH8QNbn1mc6aMy3MBrhHh4rayRdRmE/kkS1amJ
c/ld4LzcXfbb/6K1b7RMtVAeGvnZpOt5qVqNV9Fd5+fw0u/rJrZTn5zFduk+++G7
`protect END_PROTECTED
