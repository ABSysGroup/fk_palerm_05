`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NXiXejGxiS0FBZOZUkWJr4DgrKhIiGyaiPREpQUHWQaeLZkcs3TmFIW/K9gGMzov
ti67zJUKy9Zl98AwUG0+5DxC18+SJj/YSDiC9tle1LyT8HqDM+iw33iFfNw0W1Pz
SvExrF8zzAt/dLcBZLNcHYEaK9le3mV9QiTyWb7bRI6pKd4PXFf0T2Ux7k4e1Gm4
SfuiOY+ZZv6hfySOfKhaK7dVR8X4R6RysbT/DSDJHjANSUK1+YwUb3HF+RRptlaV
Ygb5Ym5DrIVguC+rRK48/cwExjHJ7Od0MLFGhauhxJghWgZLp0kwvqxluX+e7zNU
SgpVdIgn8A8EG2om6bbb0cAxXzP+t7AIYeypJwq8H5lRiFXp519faZgQvsj7kyma
ntYRbumdKVxJN7No7G7EDxc92bW2bcZJoBs96FdFGIKGXaOe9AriSxi5uJNG83DV
HuC1fMbWxdj8ki4YwYjyfBBgE95HTVXQ5CtYoRuYVQW0aVKxk8GuWsiWdNC691wD
LdQ73+4gkK2SVwLQOQ3Nvu0g608sq9m8ykaweJro7wqDl67qEHlVHU6rRngtzYgh
BjZ9oxreP+XtIklzIl3laQ624WSmKjvu2y4e+ybI5m3+LBBgsvbcertyi3q2A/vn
KNLxccxYm66KhE9ePdWhNU/Dork1nJEF3JoG8B8/z/d3OWq4+iol9VYJukUKjUoQ
LW9VVYe4N1tB3+cCZ2WcHKZX7M7SJwfcVJ181jTtH0YLRvuRSGOsSVhdAPVfxeAC
tuXNqd1QOH+fcwMsGP4591zLRcB49fXoFVQEs0xZuBGTPHICoW+7Da8/i2yPiy/H
LFtOI7VsQ5Z0LIVL2nAUXZ8bimao6vaobP3mPfYns7dtaICsb7ifuXmLDD3HuIp9
zNc4ooBsQB45husxmmGZBS6hhWETbLl1qNK1Y+1nNIdeENzx66R8jcM4TrfA/zSp
MJjUihaohxCgdsLU+TwvaMBuyuOQgtVuUicDKBoxNWoqUYXkz9v9Mh+ygJMDY4Hh
uDxI/Su4/Q5xWtae+smtn6IEyjltrryPwXdLYbSQkMrxj6r/cB4eFAkAz2agdtET
C1VPhwiIE5nDNuBA5ILTHN8dF2V2a+Sf7kGaDrHmF45Rsybsi8KDFeTdreMsRw8r
IT/R6/05FZm9XGX6k2blNDl9REeJ/8igXH9dVHtnk6dGTD14yR2cch/UlBa8YprK
TsCTUg/itC2B/EYECCk9sSAN+TwkUShoiNsZK2VA8+5GhNsx2pBdSzEMlTf5i0c1
Tk09aKaeZyJzLQhpc1O8aEf7zxfTr6/TGwTkA++BKvos2XPVZbWNpraGbKUvTTkV
e9SX0BdAeApqFEEvWdvG3dOFWTY6PeIkEVpD6A+pq/8Llsx0dz02nFk3WsCPjOY7
`protect END_PROTECTED
