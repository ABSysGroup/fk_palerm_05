`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r+VbS7NVfPwVqsHhT9kM+lIHsiPhvsbuI1CgQ0ijf6kSjX4QSLNDYVQ1fkY8grrs
w/szK7l18s+t3ZTji7MfeMgcTiF3bzBZBoqrM6uYS3/4Wyj1YIo/gcqnHvIHYXZk
rf1Jfs25P542l2ppVob35/BzIZZfPShB94G3ZE1Ew4LT5PoUaYnswQsl+HQfFoXt
oVPyV2FPspr7LAUkCtnzU9+t4KgB33Sg8JWOU2R6fQQLHCp+NtX7bUOKF9pjOiq5
Qnc3Nqq66mC4U0N2NL4DmKyZ7u6UcCp9CeAjn/F4qYJG/TSA2wV4HZcVRSyK6YMx
AaoWx1eGHgdanTCuaDYJyQtl6btHyezlKSrgBhAk49H5QYviGwVnQJF2EsYXHwDx
7ifegj747VAlJwhB/fZvHpAu0ibhujZ/ACf5fBWN/rzDsJwo48ms6pM/fkJWERUY
i3pc4wIig8RpaoN/OunLnWUHHn+yc5sKmEIgEss0ImzKw/3PA3yuhrqemSum5ziT
KMzoKx3rBQJEClBEELJ/ulioTwL5mQ2o74y5vKgI18IEPKDnfD2D9auMZF/MqHL1
CdndEA8AgsORWNPXSTARuoSmCl8hMzZY1KCzuo3ZSsWopYzdgAm4RdnskOwqXzXo
TFND/atwAiBk5zs6Nlt49sxUXYTprvSG+HbfRk0H7HGc8QSblhNVsITNhrF1dH1n
yp9JeYw7UGWg5A8rarwaXR0eomReLcuuYLwlxf8zSr+APMP9Zsf3sHFeZvE9Q69s
gX7rUKpEtWQT2dz3XyjusIyQtUy/5NhJKAV902Is6gD1Bt2yvjI1U/1thIj7huUA
jqI6tfM8U0hD/Fsv+1zGlsxR4kNjy6IrypItQOWoeTCd/j9wM8tzIzcmbwJe1Bdp
7I3qR0k9WJt9bos6ZcqGmu12sAxP48PVqYc63oBVeKa7MscpWc7t0xK6yxKVChWg
`protect END_PROTECTED
