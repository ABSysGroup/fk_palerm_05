`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2kyD6rYoV6h5xbv5ZnzJZO4vNkATwelMJIAOEjoKaEvzim6ypZh7Rd4/V8w+U9xv
R8LKqkaTAYOpDXpSxJAy3Za75lbRBpAJOkUep1zOPToLoUQXhqyl0prFaCfhO+kO
Elv96mErwd6EgS/c0MPl9qUAaSzO4mSLtyp/MAhYJPpQYH2XDy2Y6a3yVF6EOVNA
YCWrl8+RQZ71rli5qYsHjqJV9LAUckgwA8dce7WER6L2J8ISJvAZVda0y26ADYTz
jKmBgiY6D6hBwKvnrWnbqpLAPsBmrb1liFSXCulEvt/yaaonBjxWBA8RPnloPhw7
6aJ47hsKx9lYy5d+prrCqw==
`protect END_PROTECTED
