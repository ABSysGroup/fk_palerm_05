`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WIpka9Nu1gkFS9cm2T8iXSrlSGdRiZP8GGcU5seiW9/jzYjQdPDT3rrxH44htUuy
KvBaUEA/x1c6p+EFTMlKMFltYMykSEG6sZkGaVEPnL9/i9HWstXWX60MwXZiBJNF
q9Dq2u9c/6NDVqHK60ryiIYTz8ehAyG1QmFBbvkyQDtPgzonGw4RMEfZRDqcw5tw
GUSyOL2uywUCXR+ONUJcBecxbRR61Zry135g9VSlPeBnchYGvRcKSJZwnvW7ISr0
OuhWWSh1GtP1K799RHPjN6rLk5qqeUAwlKr4UNtBhig=
`protect END_PROTECTED
