`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U1vIv/JrMcvRc3f3y6/eBfT2h70QLhWT5mz3r/XhFAyTy59+wNGE27AY3Alv2biT
eZxltshx5l3SW1dSVx1T2wwyK3TNzPT8f0QQ6x8nBF3BmM4/koqXWwmswz1zLXtU
yo9UVtm+RdCz/YghqesJe9fXv0OF1Bfi2iD7PhSI0WrRsrUpzK6z53vx7AFZ0oir
xZjK9t1K00kJaANBTt8h3Q==
`protect END_PROTECTED
