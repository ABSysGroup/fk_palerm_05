`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dbepgGz9CrMr6RMke9h/tX/gpHnyryCNfee60Jr9VBWJ6Om0NMMKJVKu8Tl2hlIk
fWKw1Qa3Q6Ea/Zn+w3wRM2yEEn5D2eflJTeHUoQXtYlGvFb7r9soyTusQRkoFhKv
Di/yIC9IrgT0J6opeMN/GwZOTvPgWKJnFsrabNlgUheiqlTxdOl3ovjFqcxbfcx9
P4fE0moC+gvpXND/AK4ISek2LViyexMxxzCTqCNFGVrIHF5ftSNIMJZ6cidx3l2h
t3y4u9whylWOT881nCugXhwP22wk0917IPMcQtEL08+x3mM4LlGexqoA51huYuzJ
`protect END_PROTECTED
