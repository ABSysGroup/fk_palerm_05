`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fro0S5hyTEKa6uzmdVfUsS1E//yTLI7ygw89opqJw32+DsKVqPAyrB0lMza6v5XF
5aqso4bIo+TqUjPXY8Dy2yysZ3pO7FjZ2h3ty9TxXuBnqnAvlaoJsKIxHZOBfjYg
bOkaDqGcwOThrhk5z5dqK0oeoVbfcqiY5bbGaJMFQlQJmjKfc0QWbXLsh3GAjSGc
p45gszDxWKn7jGogcLcYK4UhvSWLHewgYLTWdg4Y/Z/8oRamaB/vSQ5wIkoHopFH
gSpUPiFv5vRjJBFmcd3LaZJzd293IFVs1OSyWB+tZhysgWeWhXO9lfgW/5Ip6PJd
9c2nkq0y/8T+nuuQai8cTlo4P1g5TZt76izfke6cckYbFkdzNnZi9l2pI8X9n/M4
eAiuF/OO6Yojbnk6nQNOcPSUuf2bn4A/qN9xXQ1ws9lsfdQ087wqyQYU59qXuGYW
fmqbj2rMpKn1WlyrsKgVdNckonWmnmaVzLnWF+s5gXpSi6lpgH6AM5VNS4WvrhJn
3fbPFKDvco3piYWq2b6NpMivGXbIKNQ9Htlob6bqeAK6OxHNFcMiFXVYytsvCYd2
0XDCkKHRkzf5fKgvKzY70N9E5Pn90rNv13xHAo/Qwul6Zp2wbgbo6zPUpuhNxvBB
9ljZZ6bBo7+8L/HIOdiRR2tqU0NOB0DlniNvTgsYDjKF+Ex2mAo+EM1EBG3h4Ik9
QWN9YauSxjaZFaD2xYO/R2j2Cd/Zg/GUSpetSDi+jar5aiKAKHE60MD9ELPSoXLU
uBsYiJKWRN0nzb/YbdkoTVLPVX6WlPB35lYxIeiiir8NcGnAAOx/JjmrzdUHVQrY
mi4DL456GWM7tsar4kV+GA1KhqWIQoUDeHQp5hgmmXbsGxGqoS3/mF8+IrNvf7hu
g65+4XYS0uKc6DHgD/D3sxRXibpBM2F7d5ITt7XzRctcTN2KARlrCuXvDzNksc5q
69jXlpKACOLSRHrdjWRIPFU3I/rDpF1D4DDqOdm4ViCZBH2+WD6065knbJxgYLbg
Rbi7be3l4ljhl197pAQiuKg6kzTX3LqsPB4ZgO0J/zCSgfA1fnWqWHG2FsnAYCeh
mb7A1n+iA2Qsuoy4KJIaknqKupqfVwmq1oXHnng5A6go7Bbo/GyWPdhiUXhYw45w
YWO7kZFMQ5YYQ4CqM/HkEdnCb7NxvnuyymoJRdAm6Ezc8lhEIMBsMF4YOOWjC3ka
OgrtfhQ9j2SdF2vDkt5J+0WTq1LIHXShp6sf7JoAc60x36wK4+frVSTbJd5ohxAl
PtJqbWtCuiy+kDFqbAIIVcuwa/yVhwjYz8XYveL2MA03EdrH3S9X442bHLdX26Go
kFImOVHvYPmzIfFBhvJ3IqXsCERQr+0tpsyTCH8vi5+hp7VPY5FFpjrhJwjtgKuG
quKJrXrmJor/Yv41TgfUxRdLVvXG5klnJ3anP6m4WGfUdF1eCBn0Wqrgyct6GynU
lyvoyQ+5G5fXHgnrHWYC+pKEbixtEkR004J2MW6oSIO2Lzg3/moNbkcsuki80Uqo
qHe19NCHJlDaE0F+26lZ3axSCd+Aq0Viv7XBu9XRdT+2vd9pQGYIR1alQ1g+IlTD
loI/+Mo1t82pxun1zemTTyQR4gJQJgA6/GBE8WariG/WHwBqGJ25s1ODKw6aDcgr
zu/hXut9kX8+/FQkjLG6SkIQknXgekjmFIZQvIazQ1iFwonDkr0bhWYBii3HCPwG
VKzxTDUHv9p+0U0SvfNmOMgGrdFtmcvUmaRhDeDeFdHobyLgl4DC9g4DKGrPlGec
T4sERvxWtzYsyATU+R38i0lZoBC7MWtylZPS+YMexRP757gZ9UZYUSOPNhVcOoDw
T+VA7qkAXCV9P1wk4QguFzVCLfHzLrdtzC0UVQ61QMWRVij0U6tj7TDsI1YbXyED
RH1aEhd3jc1Y/h+gnvjDPEWACfMC9/otaSq2/uhA4Iu/Qu94qzlOY1IM4bKfomZU
ru7jXWnNevPlbc+bS7DXHEHfpUqVIkSL+OJnLSqnetn/WBsXdU2Hv+4X7FvXo5QV
/mXNZqqXFOWNuLjYNVBe2VlMLS3l4OHZSahLBvhL8+9QlNrpM8Oq5z/Mz/rAvaRB
uGy9oWlReWrAy9cEHol1TtQUGhMxfssFFZ+tGaZ+IvYJdsJTwjNqr1HACOEixp7I
6MqzIU+/clNzcf7LaJwqcagXzZR9sPZC3kfHBeGr6iy0cl8rxwdkj/PaQFgKrshy
5r8MwB3Ea0wIQEAHMVFaEJDiXrW/POiptJLZxzpQ6GOYQgVkE1lTrE9/yvqkjob8
3/K2Jm0CKfCynvhahx3866h6Sm47Cw27f3kDjxEijImEcDB29fLBMIZOurXjZZjF
1vUCgOrMvD25ujRfZwa0o1XdZaiTJJZkvhL9AHTUZ/avMcxjT5X+a3hljablAs3O
2Jre99p8FnaOS8bZcffmwfgmHsRVEH0mhDQ63jd3VfCIpIs0eq8GVPm6y1BeCbII
RFE5/ivoR9bWczJNU4czOYdDhtU3+HvHlk3ypY/e0xjuutQAIquOrpqBhmdhWOs1
t7FBQFC3ShMAJbENcMM/1o7Af/y/yLr4GXd4ief/GPGesW0hW/x2YA1mL+vr/7fD
lKf4XcG8+G15v5kuG9qGdDhU/6jEAHcTE5K798fbMo7EIYg2UPYEMQAkkipU9uph
2g2gqDb7ul1hseB5jgdQz/epfuw8iQ3EXkP3jfSxOqo5+BGdzYtnpPKAhJYyNZqt
lHHygv8ceTt7eohGJHgCQiIWHxeRM5F8fDhPCYyWBoydMFNb6mOstSJx9lVb/gTL
rNkkOWyt4ItH+F83oy1KlJMKNg/PlfWsjQ0VmA/jPOLLCSPI4EGYnFcdf/jfQ8fa
5r2Vqc4GR45sDCkBFf9qePBERGMYDLyv3xD1Er/Uu7nvhAWIQu4H/EdsVNnWtQ05
IOWWSoUjRXEsKboCIqYKI0F75fJKBvswABb72VwUIHw6Zmbd7Q0wtX9QbsjdNhTH
GLwHnUMSTb4yg44mLQxENwi/Z/x1Zc7ZgMW/U3QiVQLDuyeQhw7DfNwHoHcwgQk4
eDQQ0Fva8uDPDzGWm4SsTzlbS8bt0vWs0BTjsr5ZC1VInic4LiRGrAbAniQmMokS
LFFCweFdUY5AKtjozFElWKAk5kSl5H+c8hnk90hwdTWc4xZPP+e5PFQ/4ijOvV+J
jgBUegS2jiJ4qr4cdSYKZUz+XeYqdi4uPcs8PPCtOkvhMl4JORETX8pkqmbRycEl
5i6KcxHLsRdTUq8Cfpm9WwTynZrUd6vgZcgBnEe/R38RslcTa9rYpnYw2sbtbvXE
ryk1BGN64UjY+pH6jzFUNPWJK9bzDynlalXY+mEGZ9mHejNz3quC3ZYTskWMveML
OwFbVwgIfrjP0joeIhdons9mhVTNnb+wyQTYLPZTzEeI4db1dXpaiKLuOg48urAB
Li13cC99WcKQGJeDAzcm0kimQNSl5lhVkwlRWYk90+u4SvTd0SmFOdXCX1N+Si+O
iqgYm7VOD8wRgPSOW6kjIrNv5LdTGfV1lcuqX1OgtzReJFRXQCOhsIgxl7OJLqKh
LCm2LVOh+Rnvjy7LdGl9JicWHbWOg1ytfrWZhdRAjExQvqZ/ZR0kZclwfTONnnJ0
esIS4qQ/Hu8yd/Lg+f6FsU/PHKTgCDT6EBMR/1U3vZfikuzHeb8CUgQGZCRTI6AF
0pO/Ja+y02FIPZG3tjTP9Z7q8nCi5+S/hP0fW8m/jJ1PHMGsuisz2OXl3DUMCErX
wHw4y1gVCHgF7TxG5SemF6o4RTHZ3kwcnXuJ8qoqpQYkLWl3AYoPr15V/fzYMQbL
1jwaXtprd40LT522uOkmMiN0k/ZfEt7Bu0txGYxRD55FG3i4z0E1RqagNiCSDdpO
DRO0+6k/ecUkHbFl4gfMDFdKWdbVT7mD/uyX+Nb0gx+8es8sElT9PGAglf3dfdEF
R8Wdj0RDaTno1vxOKD4WTVcFE/pMXBfcIcGjVSnf5au1Kw6NMlPTlmbR8G4va41z
5BHIeW0UYrcNqNGs3TLw13WZ88tP4/RyFNlRcAoxOeB8JeElkIts3Ls1a8Fj6Luc
YYeDafYiyeN2Jtq2ZfbcnrhIaG2r/NiY/JJI+4HaVe2FDVZXl7qCvAegzwWmtLSD
G0l2D4uTk1Arqr1nW0RC8USkCUc/aFLh04rJjlP9lPafZlymv8liLaXq0U+8B3xY
qjm0x1l9Pf5fYdnqFAKEtjxImN0W2M4owSibjPZkr1wU3EdQKNnS/PS8Ozk2S1QW
qKuMSx7NGmgTBZwz46c6jE1k1SN2vWYca7vQTsPT/KY+3XO29LJ04aLWp7U7bl7W
5bwaXtqVLau+Ui4uKP0zhW3GfnhPu+gXxPm2ZnCiAVeqon3fUkv87hWnaEw1FTBk
H3W6q1Jf6WG8QFbaY4E4hNKCyLOKKYzlt3xRGNFb2DiblnTgNCxi4LSCbFVJM47S
D5TnIDUFnpyQ8qbx2Hq8HIe4cqlZZJGo3WXVdASy0GeWRsuOoCzP8Qc3aHBIVK0O
tWP7Lt/HtQDDiiRi1+M9vMuQgM6KUBnA+TKIXb7lPIJxPHPbjoV9A25nj9F31khl
TD3FE9MU0J0MW/lvsZQD4zpEbIFflYOFt5GjRmixZm71/TOSsj34CYZ1Je4AoLs3
eH5NYs6ycFwFVZ5ik8oVLUtygiZqgZyPJjpC7r3+TCZGWyWm75rqdJu3sx4G53j1
lKpeKsfg4MX8LwHNwNGPl8rvBtcBCwl884QZ5ETHHkMzVA+PaILb2LqGtv1wokca
HRJLNSlcboJRjRyJe73RHEkDRm5YK+JwI3bA3TAwLk8CpuR9iMp8XyOzDr7+IzSW
zO+fhX4gksS4vxgROG5RQDh8Yxbe4UXPDrhXdOUUGpsIOT/nLK+LSTnPIJ2jgn2Q
EVreI14Nr4gr/tjN/kakfv1nusaIUvODDPQVq7fJ+ZH0ZVsOdpmrGRu6LO/iljtG
lP/phQPBxJSdLcv6z4UWIWzWHnG5tQx/MnjcUI6UMyAiyc0IDVgia6rwQ2J3MiQX
KVBuxhczLOlK5/3FPqvMAAS2OcHc3H7jUnE/jBXH2KKCr/lbjP8k+wxG42ArM7rU
Jm+XhupE/jBe6Gj+3/CDom1kNYP2IK6L68Wan/MCRVUy3yN1hf4TOXlPah0GltFU
SwVU2j0RBaZxZAwtoOLEp8tqnKILOXnbY00GXEO45oN3aOgREg6UB3Oky7tSzjUI
r5ad3JBgDCAA1gU98QHq9a2RjiKzDznX5HExKVHQzomY/WOISz9BSuTELbf7N2+j
vOpfcZwrRDBF1mwxxbfHZigSkvXmhktL7c/FDSnZagNgJ37lOFtyoN1TUjcLtlRJ
vR31dyrlnapYzmWfKQRNum9Mkxlb05/grwbonkLqHqW5acW5h9In9xA1oi2G7S3T
fcGynYRbg4d+bzme7MnMkRASLGQ4l+jVL5qcbwmQQM/zumD1rGBOC7gGSxWPEt8l
U5Y7tgwFZYjWg79BP8MBTBj4X8djotY6widk3qW5l4yatlOJmm41QIUV1qvMZuy+
Y7Va93yUBXCvZCjEt44XdW6Ow6RP3FAYWDhAoiRnOFeZSAQgquPxp8hRkf7qSfDU
FVpOOAXaXXSyw4QaYvDqzxRACgOBbjAW8p6k4nwvkF+Wsu9GfSJMSeWKryGHpjd/
Xvj25/+ifyiGL3DTNlse5sGUXijbOniYRgDfDae5UHH8oua1D82Ry2abHtcwt1Ky
B7q8hPcFSrnA4FGqse6pfWg6+NPeC9zQMRe9a/70WlnbFCF79XSvB/+AsF+ht0jI
tit1qVJr5R2UlCoKvDV1m9h7jvQpihWlpWSmaInZWIzvTAc6MaqPP59s7Je2311i
8zHKBmlFfhhAPTa+MqwMrhOZ+qrdGR8rFLiuqxo/RsNPccytUmimyFIExuKo/VU5
T0EQs9FBtScZCG3RXtxnLy3bPkmLQ1q0e7Fch3l3YGsI9e+/6aLURKcxtNV4rBkN
Eu5r4u36VULj1UXWhvcSKIozHp4WELCAfTpvRaEF8NPs8gAR1UMlQHV85nT53TcZ
g+nHms9rmDBy1wI0unz5iX8RS7PbJPGXjwq+MWzTyLvJFx6e++tak1h3F/zw15b9
u1WxmWTXcrxCdq/Ms1bTNsVfBEMxOI+4MA7GqHtAZgFgRJTOomo7muDa0zyTCjAI
gqsEutfK0PVNU04HqrLquFpIWhltDzMXfkvqI5X0K5u9yxGkFz61/9lvt81Jk+DB
R8OAuF8I1AdQHTQqW4aO7hxBjkIFrUdZx+z61XM8xQEole+c7dAd7PzLscGqjM/U
cyDTF+pILCv5bpUGts7P/nICPfqnEMaNkyGijvqyAeaZZ/nS1giZZBdEKiRCjB2d
3hG3a9qdpm9vb02loXdVxOnvBUP8QUCDpMK3SNx5AYxWBxtKrDdOCRPkYK7jsfcG
Ltq9IRAp7MEGMNxBTsG/pfkZ0OM8I517BgQxi/fktBTOJMIWrFBMFZ4OyyJblWEb
nMGrlb8p3SpzXWc9mZJ2rn2fC/lXz1Dkk9TZKClHlh3bRJoEyeaQfTHfGnSNRun7
dhuqOQkG/pwg5B1kSj0NZjZWEJDkQDoFU3WWs7ZdhsHNT3FwDkRwygFNdZIOy97/
ZEIUVCyJWUGYScHlKe2ivGZtCDB0oeTvBeNM49hCqb+4PPEsvbh4e51hid1HBzin
qTPWBQg1nxNRSzj/uU8n1RSBwSIb/MjgeraWG0HaC2Om3YTwU9BjUqlXMsTGLl3l
n2nkPYf+ZjpGISZ5qNl3dYI2n7YBwdd2w95Wxhm//ZZeFKo1bvQjW8Jpz8grq7PU
QYY3srHE+R+bNBKrgKQqAMiIblQSLYKhCHojr5+opHb58dGTTu5mhz7fd0YQybag
m4zaitFXpU5ZzzkqqE13bNVTdrBSBBHQNondIUOTSbsrj+a7fEITCY4cnoX5h7QK
t4JaGm1a++a04KxONQpRePhu6+cH+HrXhc3yNpJ/8u0tqgWDCGWvAvVk4SHQAH3D
sta7KP/lmNvODNuiunDOnHUYtNUazFYcvoDmmAt8afb7WOCvI3Gyg8Ms2Llm2VAr
LsbMmKkiJVWosJohxlEwFaC/IWHJvKKIu1WKUqMjzq3if80aW6xrf5QOyPBgwN+/
JvqhVl3z8JIMBHaO6tTTwlej8w8PQEluGup75uXDMkfLOd/kVHMdJmTEtWdnSPev
1Z9BfJzbg278QG3xjJ7OI5TFNhhOCXImTgYr3Df2HK2GkgF9MFLeAxpB8gNEpYHZ
jsNBP+C1mj3IvbFDopVXsU6VcQQj+vgdNytUFtZHhZ6/kdoe6eYq1HvmtsALLvZX
Y2UvBp5pMS+1fYtm/8l5DLaWg5SzLA86FbBkq1DcqFgiGQ2V0ryCwSO4jwDXgzon
dOr8RTFdcgpOMQuhHjwcB9raBQF14xxbgMRxgEzbRoRCcNaV01DS80X/cfrE516f
+mcgOEZ62AlALrM1CrtpUbX2kCA3eyBdbTpeknW+AsBfCVJDOit8gttRUBee2Veo
yav7IVgqae7vkVAJPN9qZS3JMj7scmQBa4nBk8TQTPEgG0Hx90KsOpaaMawORrST
O0YOdeRu104l9yQb2lh2r6nODpswo48kBv9xure9rPbFJBPiwrxl3V0RL+Pxf7Tm
PABOs7/lI4VawTyOwkkNwO0+h+5XgzEFugQ1US1q0VZCOzXWDzc/S3rWrsax9rTX
+kS5H13yXywaiLuQAv/XH9ejFtYCuQD/6VhlSt1YK3AxyZu37CqW60TsBWs0ychy
9DmwnP9cfHOhDkN/iU0t2fr1z4jvnuBul6QiFX2vj1S+fg302CJvB5dcLSkADh1g
CmzKCLn3kGvaAE6Y4oZ9OXoNTRZBA/5IjpGHEq6qCj2O3j8ndZww0QYNmd+6PZ0t
PxKsKzkESsGe4H69TdQeCE/gto+YT3OYGBohtqTDK068MgZOPhXJCPJ3bVInj3RN
JKgjTizSgEiOcFj5KskFs3XDpwEHeNzwj7wPBhPb6EZr8dNCvu5oL6eb57ZngJin
qiw6ocZ+75SKIf8WUJku0Un39hRL/7AsHWKkS3jikv0y0WYc3t40s98G+lAtSO5G
dLzbmytukZzFNBa3ZrsCV/egdrz6Zh0yj2iUN80S+bHjjzAWQEkSLzCMcnO+1PG9
069NFZbKdRXrWwK0LOS/zPXZWR1mkwbrz+oZenH6wIYNZfgZn7ojZsMjEIyDCB50
Rs1rKKGJ6HE72INuBWLeNeagMV0cGa0Bmj9Ve/LgBoBM0WmZxhIwbJkce/fSYSzv
GgIAnUay+EFFE6eR10mR1Tgc4M/Zep124tq2yyvGY5bG8vMyqsM16o7MnjENWCeR
FsOZomBotCWWJexll/TJTr9rjD/XDmBIz+eqYHbOmVnMW2Akfvf/Y0C3IC4q5uBW
gEf/OPH5sdLCdsM6vMGgOefllcfk/CZ6FsR00AdAzkp0MHtIzHeF+iHV3ifL9NuE
FLF1y++GL/RpLW3I11roUJv5uoaXj3Dg3GcDECXNqEb7UXnHFiS9doN8dmky9KjW
QX+x9ZLsUNq25OsutX/wkWK2xMdFCFR4RS38bgi3eF/jC5G3QPpAbUq1THfqUNtd
Du9JC2I9DfNYbE2CSOwgVDYBPverWz/1NrVHZs722tivkRIBW4nYIHCU/+E499rS
93VFwAWGNu+n4zYcM2Z6rB2/S3NBMuDK54kA1uadoOqSamOXJ6QCwips6IjeyMkf
9k5Gs+n+3//a1KFddiJQ6XhE0GAZhHuPm8/qo0RaZS+H2Z1Vb4fff2WhDbpHxtjn
S+wsgms80E30qmt7Nn7LBx+1SMgNUBFvR387pqvGmMowdUGnfV/jj4kKH3rUWwbU
ZVp/5rCXlyJdfbqAEqIcPhJMFTNwSnPGqQLJTZGnxNhHJ2Cin2fum76rA9WxGZLG
gZbivq/hjpf9ajytXpf02iQyhem/g3h67fmwBsf3c/qHZUeh18WD6Hd9dxmghhxk
xo1i616yP27UDh5Kuck2rwfU3R782xqUd2NlvfCkBDUVDqpPl9Qwhc0xCeTMbGYQ
Orh8edLYZqeQOQAGhPopRBUmfkt4Zbh548SHw6GRcVhJyfXyMa0Vi31QksScFuDA
24MhFYDHHAGGYJue3Afs8gaV6yz5axIvtTGWl2bATUjCNIKeruZmjRw9BPvA7gWi
JCxd8KJT+t+zwFzh4lsvQC/kZUeoUos2wpCfXQ0jAIcqdeJHMmAmxb8q0Sl4jGJZ
0bP+hZtjpNYyGH3D4czZ8/JRqQ6b6AOc0eSjwCS6FcZ90aZ8d7go7myI3A7cR0Jj
vQdbu/LmQcqkTPuiKgzTfisc9QRm8Fd7luW84zQu7DjNx/l61501nogW4gQ05LWl
lwGuAc0nkoTPJR+rNSxScpdgKHhD1U5f7UUicGZxmKA+UXXu1DSlQMd2BXjLIiB6
5/WLkWdMnCA7UhD44k+xafGDeKtQffuN2FNvibmDKvugHMpidzr/0XFr12DxWbma
jxk3kATRnpDGX7V1/cu7GKNVsC/Bg9f4TzGzdOyCMonBkpZdIfrNAnJ0iTYIxTei
j59A3GNuVox0G+LfgcAXttnsSM0xQg6SDi0WiwqI3jUrxw/jIR/AtqZXtaL9TlLG
HPYObdnCjDgmPgeDe31kO6XhJlaiIvMuPIA/G910Vg9t622mV/11eYY807NpATGK
HVflxJTkDSecmOqTIglHgBZJomfwFEw0e32FP/mcRSMA5XuXrUtXufAofTflDmO7
9ZwawSRAclxOD5QwhxbNFUOpUkpd2pTN0tkLOKfdrOedVAOiQI9vm+x6K4eyDi2S
hlBqeGAaI+U9A9YnTeiGbBQyb0k/GPRmveToc/IbM0eZoQGPBVBPb72N/oLRdb/Y
xge4Cr7lI/5npbljVR0X0Q13QgDEadsq5aBsMK4t1ziJvT0SwLi5TxRAxYHg4lH8
+Tyt7ZlIePM6kuuD6mm1LV8BMh78ljdDHogGtMVxbZlMX4NTwXDN1zRKJKYCsQvN
9BCNz4rplTR9x2DNJNjMRBMipCiDWyirlvMwkNuth0VB5iXe68zAwM9qjKhkyYQr
VLr/XC701D5iqrR4nubhdYrRkQHSwa8mVb88MI1FAR42uiQX2KsnaaQX0QLioAxB
bnkBCGdJKAw7DNJV5u8Sjc/Dk2433T+b8XeMQeWu2ijoba6a47wqOToUri7SEoZT
+u6DzAjSMio2rpcwFQ648+RVwWb6bREhLfNzFnVDJt8I4t8iUFKnjAnP8JxMxm+H
g3lSI3GVFkaDnbZ0R/qWvb/VsGtvCDaZ5V47ZgnTVPra8tIkSuCxwoT50jNfaUCj
b7G2ZWBBKdUJAawjhVyc4JYYU6KcBX/Xvemwj4cSySupT1LZ0cG5lPLsGibR982A
2TGWNNxHaJvYIFbKF4d2aH1YiW/0JaAFsssCLP4hoDxoVOvpd86LQz+99mVVWM4M
XE9oceL7gsKv5oPlTKjF0sTMO3oImeI+pGeYXq6WU9y9j5x8iJ4gry0th3ujz4Q+
ke81hfyD30R+B+Otcdu2CygiP4YpBdRpO+WkfbPQUXFoJYBXk4qA8Z6LSFUPt+Ax
SZqq3W2z9SW0g9hu1pRnYN41F4f2mt1mPwuDHwQRb5rh791Acf2o+fR+iHmKs4Ga
KyxG3iRW7OrMbejPWO3+z4s68C3KT6K66uGdP7GZ3DhJ+QYMhVgCshOHN60qxIRH
DZy1fzObvCwo+Lmjqiyl4epD3k3Eyi/Q/cFPud7W9faGGkn5JiyDiskWV6cy0MNl
VJ7LW7KH6KDTGSmfeMkElQzy/XZYpoC+N6+KvS/C24WUog/TU6TM61N54sVEGjoH
Uqvh2ZGqoauedLRjF2rTJKWV1QQQ+N3Nr8+lE3ljlaAFhR92PwmTr0vdofyAOFP+
tDMoe/y3joHXbUaofe/V58EkV4bUZ56pVcD2YnPCO8nzFkcE0jh7IBPbI1hlAg3B
2p1x6f0extUDsdtjXBfgY2Oc0WoMfOieNlIHUT5yzmsFKeAQilNfRAEWiDEYX9f4
6LecsrkDC2Vqltx1aeh/q+qIy0mv2wlK5scpT61Cr6FC9xOHm4N8Z03CddKH1/9S
zPEW5rWnV9iLVlndhoNT/0sVwxKHC8+BC+quS5S9REu34RO+JczqVS5uthO+aDK2
wTJy3A+YQjkanHQaaKp9Cb8NpR8hgrqPWQIFS3Cz1/kZpzZRbp5MK/KlMANfc2lU
DOdz8AJefFTY3ulf0v//ti1gNB9wY4qB4en0wpc4XiXdS+F7lX1e/4YIGlgwYk66
1OTI7/w8OswTEONtWzWZRiA6yYzAOOAZJqwvr78Zf4gxhV7jufB2Gnxfp1sWiMpw
Thngl7Du/Iyl7VVYnwl1JF82EhITRcpVWqQePT8zfgUP2lCRDo2VE/sL+/64bPEL
P+rz3mzq6QyfaHGNsy7lRASwjCjZ8Zz3QtdVN8yiWEBLmHdoFnMsdSJi1GWJSHLM
zmrnT7AIud0sLEl7LQshxCkbZuJeumsKpZIuyNTYk36C0G3c6Wg+h56QSwZAkQux
uUv4UzhhQrE1uCmLwqhTb3/CRjXbQyuMOfDEU7+WCFe1ON82Dbc/ZR8Bmb1/irRD
gqwJ62Yk0xY8RTvbmBEr0TvzynGS0vu/pHRNC+7eH9x3kYPMb9fwVQ3JDwTMB8yt
tw9YxRJhVKlMzJGFL5hb94pcvAZs3ooJYZtEqanpd1401OU7DJmqE7aMeNFmTyGl
YmoUrdhkNYN08xnmQACNnaHYGNUmv3z7vtSIE+RYiq3Y56IsfFWXTwVPj36Prb3I
dwA91HphnZ30ZQZC4dgEgABe3EKdwW93ASeIT1P11Ecp8Bwq/516WAAa41EXQ8J7
d23yknOaV/aSx2VuxysU1qys6o4RrtaNWXuDdTM+90MOpJCgYSJ9kt+WydRC4FKd
3sgK5qJatH8b/mS8frPVsV+am6eIdTacqlvijjSYe70mD83Ro89igN784+DhsjqJ
/Ogx5d5MSJLxlwp8+i9ut7GJy2h+KSOgImpBOGq/KpeNISCHbmVCB1K8QE4h53KE
HeE+b6GDH5srZ1mOQ85yzbI7xVkXjZOdoJH7tTjByJooKdB246you4RkUrsovQVm
01sZ7cFKT+FFzx+fs+FsYFvtHQIB0dxwGwDy9HV37QNJhbagss3Ll1XNs+7Yx6V7
5UdOy1g2rly8/ghZjDfNBq9+JnLin0b/fR7wgnTapufm5Cuuj1sEsJYA5/5gwgsd
Z+0m9JLDQUs74FUFO028ysjCopldS4+yuemo0scDu0tQFh1Efxh/Xx9x4HDCjqZS
eEpkeFJEkh6eudYWE0UsI/IAO9FzWZJCK0/mf3ylxa+QKsMQGyGNFbJAUSTqFY+d
posC/P9NquHhb9+TQbtp40cAwoN2mttNx6conqzs0N4gCYIrkzXTTobwXuyjiFqO
GbrCVtT0uu6EGysxEjBWWn4g5bfkKeHNIREghTJVd8xxBfUo8YExPA7A864BeFbN
gf1QW5HgrEL/J+SACip4KH0MjhAfXKyeiFe+wygqTkdFAQHyND2U+a00QcBn0lfr
lwgJBatJPEVsj868XPbq6geGtemUMyKLWCrMnrVsYEaPvhRRh606OPzc8rruPOrg
pay3SG00e5fYhX7nvIbMKTf/PvfvoIY00cspPk0Gi77h+JrlD6grY1fEWS7Mr7xN
1tGWxErbbwTeSmLyRQhYRQheWUbgCiTBKequuHrAhzLpFsHxkcL+64TujjjAIUQF
xxDb2nZvzkj3bxBUqaPvzo6QCBlWspy2SgqzbQlk5gSOrOBZylPrahk0JGpxelUi
5nhOINE09+ScTu/+rKqk8ahWBfJVi+hC3EIP/VI1qz1V1Cnq7ojBozJhB9b8vqRN
tjy2Rw0mDaRyuW05/E0msRPSBtDnMKWeTovdYJFDQyd/M7pHrzLTvjJ7gXkWhjIO
0XdlMZMyaQLLI1naHrU6R8eJ9n5d2hPnGrkWXXSaM70F8DHVf8O+4ACDVk2To3xt
dDzb0NOmr/lagVnMTr2bbNs5ET/bfZVnYvb8iLmcWsHIRapDQhjhWutRzFULPqjq
JJhjTLW509xse17zoj/I2TUcMWSFVEesqq7y4v+TOSoizyubzJ+RnM4h6MVNSXJ0
OIFhlur+x4dUecLdg1nBQ47kkXKndDAzEhIehBHE1fEXEyvHLJ+x8BzrcAdD2/uv
ULRbltaLkn0wHPqPT21BdRNJ80soOarSzSyhrlK+QwQpu7SP9qb+sHV+S+hmggWn
ryR1m/NfspOOLqUAU6t88RjvYxRZIc0SdtLjyX1rXs/Ve3giVk1htHoVSM2uoXoe
L639rhXsi0sPKViacp+WQcFM2DBe/lPdq+1HxafRaLnyMOMVzEHBH0jlVCoHb7bw
Kpg1iObjTd1wzr9B9oz0LraVocTae0RKyPjG0CA7v6Ww08kI9+6OVG63kbGXWMR6
Dc+jUNyVb531oNsH2HIaCQccmWvSvN4c+JU8WiyyxcikqqBa/7Uvy3rY4CoBAOSk
KNwYPyzxEf8W8r9VvYzHzqoAgr3+mslo4xApBFHi6tkrIMPg7/nyDvT5wiymYIEA
SZpEyD+0uZzZe5HMw9OulCbnxfB5dMbzgvZYsYq+lPbJ81oaOqX+0RXTAzWoYt6N
HajLULeueHNFYaQsYOLPOqlbsGSH3ViCUH1ZOt+48L1EXeqKrCkfJAuuWl5F8k3T
zwL9N7QwNxP6t8o4Iw4meLQjdzEIbQZesNFvo0fDiUNlV9L0COq0oQEyW+JXAXfP
R3+ecH5AesUk63HQjNvqNGjZmyIbV9hL8zwpy21JtI3rD7ZV0GYcaiJV6bIZyG0e
SQJOElHd+v79jssF1rZAk+thCbOutUrylgKjNrOmHZHXap3lOBXZEhEO6TDkBo97
kcl24yjqt8D0C+JLoEujJeiZ3U0+tpBmA4aZi8YDe/qZn8XgafSPw3ynBqv2OePB
i2Q7R1rILHhI3qjSf3A9GSY2HUbYOz2OlwzK+swdZhsS9rHaNak29qrCSaLxFWDk
XWAg7TmR+pniqdLmBYeUMqw8WLzGHADgMzGxERl50AO9gTHf2aX1mtkmgeG7U/HR
2K9ex4Sc6ekS1ZMN8tID8ks0w69Btb74l6i6LW6Bpwc1KOlEVyMNs9vCwfWe01H4
T/P0oscDu7umfz01edEFDQ3xYfwaRWy0+u5KWTk4EqHDuCLPQHAl3GSyt9y8xn88
xu8pU/rspI/nUNGTLF2yQx6L/TlQDYrGZgz1o1uYXJoHTUc/DTPjWSYdaJ1E4Vgq
4L3oB0/x87Z+BNlCVruytFGNi+DnOmKjmaLnO+33IXqmznB5qzfF9FLUMAlBlEWt
xjddkWTrAUU7X5lg1OAnB8zOlXS5HFUGY+XsgFgIoUPaLUI39ZV5FMiMSl92F+YZ
Nrn8zWNBvfCLcJh2drkuWkN5lgKM7EEq6qVQIYsTrImsD5JI1EIVvv/4MCBHGID+
5Ll7SKj3/Utlybt5seQImVGGtQGTBwqzLsIeOuXCoaU7IJzzQ8vSYmgoYHUcMC48
WMEJT4SAuJfrRJy+uLiTBF2xymLd2kxwuXwioTy4tAdHX3FovwdpRmK6SWjd6ri5
8g5M8KYc4/UAqe6yd72Jtfoys1uBaYqhw//GoQ0kWoIxENcOzjtIZeE6adZVS16I
7fjHqcU93ggvascPfTLP5lzNUt4Ttex8Zhfi0qeVv1tikVDdX+Hv4h96oP8oA6MR
WSXd+1yvXbCF1pmo/yx37HAX6nlE2aDnqwucDEDQ2efYZ2+KWbITHQE8YcsKmD5l
zk6h1ogclV93fOrO5CUmH5+Z6vP7mdFGhj88Yzsfgr4e0xtIwk2kPevGsd//Dz48
vGKdrEXU+xSOjS3HDpclW7QNpF2z6uFtxoznC6NeVXevU6Bj5CFLxwfxgVNAR/Kt
qv2cAeBjND0yHJBMsyW8R4Fs7ZejOhIzeYZUDNQlRtOBuNGU8qp00NoCBo6AqJA9
oaDCC8b6GP5JCphabEYG2rd1imUvVMliRMOsrB0bhP4c4qzJKw8IxC6vysV4G1Lo
VTlmiLtWc94AyHZ48bc4YrqQgRSuNL6H563c1Lfosbq3Fcewx89i1tk6jkcJ+rC3
XHEJ/OG03rtZH+gZPt04qF7/RTu7P/45/5eXr1cMX0yTVtWvG6/RHZtN06nxAHFm
9njfMnBLMJy5tZetTEgH3O/O0SkqPbOV27lOB+P+cNdDMNeuCyphaCxwVZqcKfFZ
0Siul2+nUNaQeVZqxxGvojYYg362N9swSr1K8xI/4oFc0+YOBgx57lgwkDMW9hyT
NM17L9jBEzXm9eoYRQg+wUVitKBCid9cTHz9nDPGhV0p9etKVgsEX+oYgk0u9nyu
tirxy3oRPCzMoZS+Pjs7hZnuh0mEohQ4uaahYSxjfyrX8lYwY9XjSVXT+17COvXm
7+6zHwG9trND5CVxuSA3eV7skjrS9sbzr2bh/gKfSJcfQ6kSczm5UNiSsyw+biKb
8+Ycipk9g32rqe+3Co9Pm4kZ//u0ujuWsYLromIKRqAS88l5eLEGeWdTSmxeZ82j
jvKmbkVyzv5gYxrDF2Qx827hrg2zHhfSyZtWSZYZqw67wE3au8xx++Sm876/Dqfn
VLMmvG9peKIWfTV8tJGGG2VzlBn+hnDzWz+iueYOXBqqr6fM6ZFnuekZi+BsR/Qs
shF2YceQ9/iETV31FYRXgFz7abCXgCRyNSJt1l/YuxLCS46jBfjcyK2gH9PlYZzT
NJRC3ZU7G3jWyKmd7WzJb9nR17GJVKoKed83g3Awz02BFdykS4nGi/A8yerhx0m7
xG+eMu7z1GPbWtYsRSBNFmYuYQKB+26yYQgR1+PP5auP0QGmz2kMOTqBV+tDww/E
u9hbWpmskG47dK7IW06kLp+Q/6SbfroxB5JiGlRq18INVCqi98e4vtIRMt1OI/fv
VPmISFCJPF4qEobN5fa4PQ44MKkIJeb9HhdtRfLoR9vedtIEs8rQs22UhXG5/t4d
UZ+7UiU4W0+tGIwJCvirAIQzZTqTQtM5nE7JionKf0kie6lPWqz+daiy+Rwf5TjY
+bDZ2EmnX8YQ/oq4WNymKFcPU5Kgtgpo2kBo13qSIB1XX7q+MiyiF9pYh50ZJ2rm
bMv0f8/3fThJENoSG9HGRJElYf0TzocpO1IA9RLRXp1679ZqUK7NIgSbR8rWn54+
39YUaFYPYVI9Aum/+cSdGZTJqDk/xS0q6s9kw51mptiRe1daQgTkRi8uFFx2gmD7
M2QfUO0p87ZilfmgTW8zQT2gaYwZSdrUTtolw5uLLDiB0BpPkVdyZWDRy0esCx4J
a0jONBVtaIBWBfpwwvoCJLvyqnBvgOlWFw2LOmFGCQYXPLIKqrbf91P4fVAAmRpX
cw2C7N8PPnTgbH3AIphzOh5G3XN6KRdInZqh5lG+GFwHG1i283lz9PdXAo3nS9Ze
q/b14xTrqnyOW90WPiJ6dJZzxzT8TYVVknNARKQkrBlNAz174R0lDjo0px1XQOzb
AHAAZUtnT543ogG/ZJ8rwQya69Rc6JV3r4GDMqpSDHdZ/+StPlhTI0SbDxkpD8GP
M39KvRICfu6NCYxvGe2NF/ssIRUOKEMgch0JssgFtEQE9S+ifYUZFIR2DiAvlgBs
XM+qDS0oYZCpEDcBQfQrQG5vBCo+OMPWkBj9OFxlaC3EP2wGNryPNRAOyvph7hA4
lVvjmS44CdndcisFuLCkWpsGKBdm0t0FBk6voizYLGW3r46UkIc4kfPcZJe/l9dx
dreaBCltM7nBUNK++knOLWfXtHeNXOzuGS3cuWs+/3gNSVe4JCRVxdBR+Dsl6Lr0
yEBsFN1Ce5T6W8k7NkBuQQalHCuXpq3jO5Ss2E5EVn6cbjPbd0ZT0dr2RwNCPsiL
V3vyNKrzKmLkb4mj9gkoq74D5RmEoLJpUXwbxCIJIQRaJDiTfG0iiettGl/2TMgA
k7MfVXCuYXUx1oJh3IFPl8kMgJ8TPIkrGsmJghWPa8uu4wXGw39pvGVga9gJGYoN
6n05pBByOZzF1oeo790+RsSA3qoEZXevSs9l6UIHODSpCzKYtVNT5Cbls76WUr1g
Xm1XYxZNKkL73lzuNO7NNiI3ZYmH8B2RlusifKkOK/0d5fixsQQsC3Im/5B7IGIm
b1QDjFZOfmHja4JGKHb+5lJkWlK6r29Xd7eOZvdby+jYi5l5EefdNf4hoV3jpSYE
5ywvPHuh6Uic0E5HH+jb1cGm9TReJIMhE47t7xuaW7LXKMwkTG5VpViNMfJVQw1y
5VvrHOA0/ZaO4yosYlbmVmgmSRLwo/kpvf4lEw68H6FmOOnR7t9bPYnPvtASUWSw
LND872VnW0K6NP2nBNdxAx22OaBo9RyLT+/p6fUbY4ODrGcurBd6d69YeTP3JwUy
ry/Bsptj+90lKBDor6gpJCmG1u0yv7BgRXFFbNEB6322CMGpKZT4xFbc8Wf/9GyS
0CBN/hbpXd3x3Xh7krJtnsj0IGiZ5b82XByIFBcaAriEanRifCr9QdY53gVlnc+6
vFuugZwkln39CulWOb0mVKJRfiEpoY8wNvcCIDb7gTVx9uBQmomcM07GCUC20Fwc
FkjPY/XBJKLk3wQKgDnG4PuwiBQOM55S0IwTeTZDvtKDsUDUYWae5mcNi22YGFLD
yOXuPrIV1jWyb6ZxAR1/Jg2Tq5DgrKxLj6JahCs39X9j2bAneXRdc8DLSFdT4Tjk
COWL/DHq5QehdVNkoXSKoJtD4hKl6xgN/5gZFSLl1WlsULEr/F2D2QhK4NDOnW0a
/rGKfExpBHomw7zzz+cWkqy903fC6IcZkdHhfSjo6Pr1qtjj6VqceVtmMCAJuJvu
HdtYiMOBvInnGAfguWJ9UxUq2LuXmwhDgm6n56iKs+DP2FF8b9q7Lp0PK0CKtJzO
V6Q2KMKS8ib3FFq0hAlmcOUoSwyQJO08A+qr7ybHpVyqvTCQPAWDszoC68nt64hn
6T9n5zXi8+bt1ig629R1EHuko3hwobwDKMsvYY07QC2rh5DeSxSZA6Y0PosXDOEd
nImV9++hbGhCKfAF3Au/QXGED01uUJCQEMosJdHyzwLC2D+N8SUFZgB4v2UORV2m
Jg7u1mNguY7/VtmCrEJ8jTvTCTm/KDApe5qt3XVfBxuFJUZXeD9/KIQPZU3CtDPW
KJPYLG9e/akrE1Po6b2BmslWbO9N0EWdEkRjUTODCkk0urXe1avSkj5dEJt/th9e
SbzoeGZVy94kd5YCIwkwHqiUoPAbENpsdjGPt/+Obucoxr52FHaed7pZzxsOCilm
z5l6GlDxSpU1mzQQCp94bVsdm9OIyc1H1qyQx70ol+Imdqu2pIMLDAwA0iCRszWV
lTaPCb1JfO4VSGlHCAb0awoGpN3uly80eUnQVAYyy3n/LxRZ0q0dclKmd58/xp2H
dDWSKdiTVpUoiY10eDjXQl7hIPhnGnqUpQ/I5LsOqmVLPoB/tOsq129aGwpQpolZ
wYi9sOAkuzjQYbfdsyTmcWTw9/bHWdzdpSiOTB93Y07YLgsOM0oHaRXutRs3LYoK
wBFrFVc0A4LY1Q6YwW2rkCEnEurQu5aIt5aHZj/EsIBtiQdefS+O5J88d3iFk7H8
kxZDGXgZ3eBAiBDe2CHXA1a4FZMI4LBce9xHbGLfv1+Jj7O+y2j+D6XFj/Pjqcb4
ezk7TwrxCAzOd3FR/rqCCalLxcC4Pn1BLPpohq6vex3+6NqhV0QIq1Q1sk+omKkp
8clnrZbcZ2sv0WuYhJeCtkm2hZcswnK/jXk6T8zxDwkVhpAHFm5RbIBxD/yWsyXA
SvtR2odwxdrwnp+u9ASbwdNgSq4EeJsUBmqJqXB3kagqt9ifWZa0zl9AkMrrO644
tDDqzLiCkYSQSxnBl5uaSzj4f+r6cLztWa0DhEAN66lgwhSAUHITeKV+CEtXhPtO
bLQxn/9uOFlSMqY6kM344iYlmuPYETZzKj98HzZQCk3YJFSW7hYqwI71KhUfXacp
Q/a+YCQT0kiBdmvt27sDU9wv0lYSpil1zyG5Rl00pjBaFPSOYKB2jr7mKmr2NrxA
sgkAD1fHs8zefKT7jb3vwdBB634cBSxAUQsN1wU7IiA7ICyi+riDFuls7qzHriq1
nEHbDg1JIkCnyvPahJH07/ZWJbNKprDxqefex9ccdG0rdXHR6SVRGpyGrNWbfk8l
EwYCm+dTeiAr+exlojTTvCpzxdQL1X+Vmm8yja+RoGBECUryLbwyDYdf3KudqosD
OR9mwjdnnSrbJVGgEKoRcyFATFYYcsM7xFncRInCxUsextMpwkwdvAxVuDo+wf9H
sGe99R7C33GO7IgDW5vVkEAi8kIJ3wU/nabsdRokrp3hlzKG7FvyBS5idNRyhVUg
D55gitx85m/gUT1PhTlUPzfcQ4ilsbLQ1ECu6An0oFGBvRpv5xn4BgtLQ9oTmJ4O
VRs1z4m90D/hUWnM9CysGmNM2TzOtjAWBJ9m0AUDiV4CGocslsl2accUrE7pZIpj
eonk6AsZir7/Yo948l9csPdXmnNQzDnU7UTjo/hiX2WRnFzNWXqoT0sHSIjbphOQ
Xoi3jrQrQDBXLNHHwaHzYw==
`protect END_PROTECTED
