`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yrGpUSjrdJkmarDQmCctWq35QwXU9vNiHVyCaqUyUENYwJvfd48eWM6icicMe/OM
MiCEbXeK+g5ht4S+Cg1yL0D68RF3pndGi0W7WKf41p4ohayAFLZA2g65L0NHQHOU
0fv/RhphDUG6L6Wl0DASVNHP0FbL+PkwFnOweHC7JHZulpk2iWHqh+FwdLn4qJeb
Wf+ppMLmGKQ5gh1FN/01EJe2Ewk935vxG8movvRvLLImmA6jKSegwHcH5zXm524W
vQaOceVgnsuzc0tJSbRANdk424EYB3cAFKwxDZfev7pElZau6m5D1HH2ZBLl1/MA
gbpTqJoGdNdBmg6W4Zcbe7fV96utlVKYzfM8qF+ahfPtrtSpaZHQnp/ljInNakhy
iDOxh+ruowL+fyiJdUWVU+3ACxF5fQbxlCLX12/oO9pLLjxXs7FJ3y3dcMhv66TO
9OalT4Dr6goGiIPJkzJEWgCgAMXqVHQsycBZePvzHFMZYydw7OL/AK6h+xXO5tiA
AXEOvT/WcvN0qIMCaGoQ5GbAsAZTy6g3oC84Cb3YnFETac8ONW7ZJ6ryzNsP9OwS
p5t5PR7VuB3Q5a5HVMG9YcI8s9hcCS+9NpgIA/nR5MIRGKGNEUQ5lh3qdWdRXxVX
`protect END_PROTECTED
