`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ML7HRZeSU7Kxb8HjjpDXgC219XVO9H8L3HH5iLIwIIrlJInCyVqPkkfHWykWP7zM
8UeKxrsJ29Caf8+tTHEKqccaZDLgiURnVgshpWgln2AMML8sx3nFJAZ4aksPQpLU
IMoaorVwJS+p37OjiUuyE/R5sGxyOmBigkYSWuyzv9+rPLWxC9dGPcorQmPUL6Ce
lfl5qLrN0rMew2VeyaLmDaSuw3oGDaEuFTg5BPjxCreeg/ovNXHaYnOwHSPNDto+
q/lqVKMCavekNAArvdlOQoIYEfZthAwxf4UVJ0HB2qX9MjwA8ejR0aR1nbWzsvow
cVHqp9bWo12sClxLpL5WJ6GNzEq1hAjiyB5J66lyS9BCmBNKcif3hRzFLAfrihU3
q8//P9KF9d5kBUXBug7dC4nEnM3xdsz2OAXGtKeP2GxwZkvFQSrA9oNDxpJOcAR9
zKUVVAR63wVcqizUfHwh0ytwdHCnqKnA84KU4Hn1TXzydTsk+5avVjqOmfPlGFSh
eVto9Dbk0KM+GFNQiUr0n9m414q4mKv5pOyU+AWHVpVVmTAUZYyf6bRKFbWXvibb
7otzkRo6VQbo6QoauJU4FONu17rwu61aUugkJDsjVlblRgOmvBzhQzC7roEordoN
ovmISA1ZfRAtyuORBhkao5Zsgo4B51GWSY0rg3HmAWRyDKnXDw3y41ZkfiCSQKtI
1J9xjX6o1TDzEQ/l43DTNNiszzT+z64W+Sk++K72oYrUi8I1Zu5DM4l6wOGm9m1j
HDVW5vhhWegisUAT4yt16Q==
`protect END_PROTECTED
