`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
86cc4j5DcSjil+C89T/7DrjUpBdCseEDVCe1rJ4LcJV18Pbc+scwxVX8gIuY+9p6
KngoSmGFyXsOPBaJzabjcMt+9ZqyTGNJsRSIK7ETmoqyRCupi4505tWZUOHDDUnV
GOkKa1Mfiekzj4g+8lV2V+LAoAh78CIUi7vSrrMEkAKzTDiHf+wj4ZiKJL+A75FE
pjMZ9fXxRPMnbq/Dr/77TojWQLZgp14sw09XkShtUoDSMBQNXnOyTNPeuWJ1jdSn
AUsupYWKKkW6X68sC65ka0X1n2l2ve+kYKcI04dlLqAOb0PJ9rsYGNdt1Uru1ok7
CdAmcWhM5ODQtOzWurhzd9s/8NJZp3GGX7Q/eronhXSqky2TwechM8MlkIiYrnZr
C4NdBzuMSPu8SkFb2b/0sr+JJeNtF9CAyvkBtyKaY7Qc6KuKBE/J1/rn3x8bS/6B
jUKtWVUeg/Y0nggvr6RKra7xH5baGXEYLnTXzcNtN2XuvocKzh4FriE7HbvD9s3y
hqJnWPrn3gvHiJNhUGPBO2xzcj8iPh2LBo+Ye2elg7BywAFtMbejrn0Vv+ckRpeD
6RSNTQ3owEJbqKePqImsHdqGm+xi8L5CGpolm/AfPEIUMvcXnmZHhXOTYjwgVerW
SIEIuvKe3uyZESPjPGuhXg==
`protect END_PROTECTED
