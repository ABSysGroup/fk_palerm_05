`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5dy33ofNLJXVHg3aFwce19zwUfIgJr4gUJIpItAfLxyBpTeuDoO/8YhJC1quI/Ws
pUm9lZGAotnSl/uoVqZeDapEfrW4roLq/uAsSm+bLXDJdzQjb0KEOhoD3RLjJpwS
VfdID4tn7EonYV1UUT1WnCrUoj7ep9i9zTAykCng+fbo2gkbjA4nWKzYP3XzQIYI
ioXg07OWqn56ySuEpbG1xnnLnwMIpAB3P4z2MX453PN/4GT5w8Va60IuV+th7aYV
LQ/BhvrZjOe/V4Ws9ucgDcKTqmayJ78BNTYu4HCt7NjqY/za0OyTOnevc9N/VJ5u
xfuiYXbEsrNYP/WMuKT3+21zQNO9OiGXPPHS/DQuuAPVJMqX8h8EgARf89S5Gm3H
QclYS1HS7v/Gth6yTJeGtMzJ6X3ReCRe7MvgtAGihVKfghzGxJwuGyfekhlBzNEM
51DLq4+Jouj8w9y79J+faSHFSqYMseL5V2uuTCn390+Ji2pneWWjYzONQekMuESi
he5u8M4T0ZXX44PrP/e4REwvOBnaYvIVqgnPe/GUftMY20ESXEH0f2hJZ28dQBTt
PiDxaw2eRF2KAkxc9gEeNkbaZ+N8EU0RBhWBYu8Fs9TP245uC8LSii5RZdghXbTy
Z3AskWVyGHCa8rsSK++V7jfYd68kb9dO8j6YU1yBXTlg3sH1wOl4V7koajT8P26q
2qQfIwVMUKTRWpGhFw1TyOxJvFMMMXRgYooYgaicOGU2Yc3eh4ZkaDy2JlQgq4Cj
z5L0+sAxtn/BxDXq2pg3i1IrsoMgRTbeQV2n24KRKT3S8ODprt2XYZX95z0EQRl1
+QToR6UiWIljchgRaD9Fqn1JmED/b2A3OIgcWiQ+Xe4mwlXucwaBa4NxY+d7gKZK
gNbaKZFvPE4cg8piqiB977d++fUcwmSbAm47DcLRqftmhPS1RwqLPgXfzuM3uPoS
50lwGsEXt2ZbVg9QRVePkUO+th3oETpClkbq+F1Hr3deixd3cFXYIxOy/sOTscy0
Zr7wq+lk0mbRkOOPSBzW9kVQacFCjBWkQcrpHPz1uh3Ou89TQrMUbzel0BXWnPnV
lKGFlc72cgvr9U09uKxq8IovE6+VUdUMjjqYdSQtYaBiyl49xVP6ag6gEr2uFky1
6gqDHirPLTCLdUYY4+CGZC2FpFo2egPMElqmYexrTob2L85t6OZ2Q3EydU9PNnKi
EU7U2pMqovuWqrwluARMOklS606l2ZK2dEne1xWUMsqRXVr2xhOdSbpkz1ljahqW
xwn6c1AENkS2UGcZBEa3RCc/ayMmEinhKH3YSNDPeIyk6NanbcBaST8nvvG+TILh
Xoma8DGENiMNL2VsoEuv3lpceFo581dcxM9DD4C0CS0rqWbng58sc6EWuBI0avW4
PSCm11STEC+X34CW5pppCQCA+LZAsgdO00xwq/YNkXVh+uPm2svBvedPGPzC3Ucm
i9dpvJdVGpbzBsEWXcAfTuXFzZqx8bnXsgGHNQESIZ40e1QAtr5UKf6zasFfegAX
IoguEyROVywO+wYPNOhe664dyrFWnc+3HELP8IrDbfu/Zi5uMzNRsW+HVcjCNPUS
g6xiThxxluGQuJaJ564WPXoKc9j+/UyZLspFn7ivDk95JVi+zvGQf/onH6ZNH7a5
kF9nzqCiEYvNRjSS2idGlLxOq8JPLPxgObmcEJJ78oa2GtOn8Ft+BDaLWGnhwM0H
k9yF6GuOLHcGibFUmSUzdqpjPPBd+YbtEzkJ6EPkecMejdgJ9+tNHeL/ZghiK3ja
l+OhLZq2N9nJKYVDNmd0vN74HI5Qj3WDSliHK4KDJTfHImm+f7rQWyGDepAWFQHh
BMBaMv3O3zvLiSpvKnFshp7c/Ht78LQ5x5ADq462qpROERjOkZdhS5qoU/42WarJ
04uL8khr/+dupz4foZlSATrIaz90aDc5wtUeFJFaw3yeQhVzKYQ3muhwXsGG2T7N
mzx6ETYOY2AIShpDH3RyfyZ9NMUEg93maacmF640nJ10Rr/tn55hkVEeU3kYtLhs
4SPPWvVvRb9QeZAnx0iAf8qWoX31+7ayLjFU5qXm/sd0tg6A4KUSA2oHaNdgx1B4
zLs1XxGzrbtwXrjbTw7XZ9OXE0f5I7iwjNbIPnFnIzhd9iBOw5h6nLX8oHgQRGOC
Al0EKHSSNLjW5EgFyB/AqFgWL6VC7WHcq2cXbEXR7YLs7Qnd7iOCEktqCi/06K2C
nK4XMdOMoM2BSvY8VMIrGQ/gNIGHMYq1WMbXKS9BVz8dnUHw1n6uLado0QHDuL93
5lOY8tbS044QZBdGujj20O73YoZjsBBb0IjBmxMAWLxkUC/hSr8Jj6o1Kx7XQSsk
kdXqjG2Qy/FLeoexJuA95rUARLrFpdDa+QRXhquTohE3Rqe6iG6XCkf1frh7To7H
kHgAFM4cnpM2U999lXKO66ZoTrnm+bvF1iRVEifbAtcpNG7P+VuFH92GFwiu191L
PE5GVdtg7uwtCXWC3BUr5kr7D2fU0njgjovBB/ROmBM4QjhlhMcYR2mSmYUzZrvk
0f4KWJlnkYMkadicN86Sq7a943n4nnBxlaK9DZ7w7qeUoNsq/OmCiVJEbImgkhiB
tB+TXzQqkaSLlYEDMulEstbDI1PYo6Hun6MGl2X3HpjUYxVdaY9Q8bodYeBAjKyt
CNNHfjwgDNiCea2ej7ClDOICpFeYrGiajPPS1yIc0Sd5EABrgVlo6+UujQJ7a4+X
ZG5Hz5HVfGH9MZgh7F88Io+Xzk2AwYxVo/LuMNikZ1Mfn7ZeXF37uWtaBF27iBiS
fBWiHvd96G7KDqY7zi/mA5FR/146eRhdx/3uMoDIOP/85maiqVbDyCqElEXXZTmE
SGXss8b/re22KzaZPLSB/+Cs1nKgiUoj78ZH5dvxktthnKaWSXEoFrC6rArL04M1
lUL7m7Q8oPEZmKAj1kDrAX9I820WDa01FMkpTlCsbPGXPMI9fl1ZQ3snUr9qeq2K
mrGN11E2YbM3kkB4l/SmaNCV7im4MSkBhG6afv9Q38y1v1VgusvgDDoV1xmhdNIf
0PxujwIuViC1rP0je/RmDtscS2QxCSFX+3e9pK6IImVGCD7ODQzxKFtovP3QiCwj
R+QWxyt57eHawmvnTWir0RMRP0IFRoo3ewDPNnoEcmfTxNQKnQfO1O2mwY9WkyQq
92wKBeFe4maNzqBsh0IP/itKmhBGJQl76bXjixMZw/x2o5IWObV2S/ugHmWH7hoG
LX0UnLUbMtzpltzY5B6IS3VB1OCuKhQOw4hoi1pV7dN9KRFdQkX3hJxqsMqknQq9
ioNJZHrrXQDzCMpkUz2ntnE8Cg7ZSg3Nq574WYtIORUZ2XCZ7Iit9V9L3mlXBiFa
QomgA9xQfLcH1g+DtI7yoLeXgfAhQW6k74YQ1fZJ/hcF1U4PBr5q5mKpndocUNoz
+wgOgto6GQWs+GZV0gecdCVUlRp/o/OXy7kTPsrs50ChntJeFRdOxyTi/q+obkYF
kQnNWCtPGuheMZqVArkikAsFqcmfreGzQ4ILeQ3v970iAiGSOTtGggGH6zD4+eYO
V3LGlZPx7dDbLuRtEtL3Z2mqB4AvUm7mrpdwG01TBjV3/s3x5Te4uRfiorUChN5l
25Ws1J3lQYlO3vN+Gx0LdfQ8l8/+kB/f6hHOoXl4lzk1eEu8kfYMM4xyiO+Y1IMs
KV4ZegiLoK7AtVcNmQaoLuEIXPW+e4M73s8YYtbMkB3lKJBUnB+4urUdLaWkc4if
1kttu4r4eejnYQ1f+7Wgb40bEkRY9yqqMKpXPwdOZPMrC740lTfH9yyqYKgG9ub5
uIU/Q3MqrEKPHnfluQMIAUkJ/oyTp8olmtKb0km7ShutN3INAcLI/kR9aD0V7Qw0
L6Anf01IjX6t7vPhMr9RSk9E2R8WQ3IQTBazA/piNBTW+MZ1PmKyMbd4CDDjJRf1
VTPo+UobgBN62N7tMnqFzAxniY1nvcYAcHI9wE5kkq8pdA+mcVzjS7RH28F4J8nX
ja9RoBfuWvRbw7/QC7jYRE7LcPJfnyj+IHaJNi5G+iEXAlfCzd9SOKvAFw+LirdN
RbXQ4r+w2vVONBjMhn5qKzeSfNphLZNcQtWIfT5kxok5tXVjOe7kydf2dIFOQvtz
1Av/jaqPc0N8ZEogxNmDVoOzZ+mEVApcLwI5B4i612VagW7jPo4X23y4bEK91Ubr
KzwRtL1d5SAdqyuTXgvV+TEGLULzTAQc1W8o92ZDau895HvVCxByvDkqkoa/185U
uNXoCPtYPHytGscrTJyXrWQ0OvdWTaIfmT+rYLqDyidl9s6UyDu6KRG0+eMMkvWd
sBCbNbfqOMIadR+JdcRCX6wnXBdNn70l46fMwLOQeyl549Dq+UBiFicmk36qXOyX
Uf+JRe0fgAFgu2wI6s70TTXQlwNT9S4Cd8WX7uWOFitGPRKIixT/OQ3fWj0oEV+W
rgyXxl88fF8LMCl/13kolTvIw6Bj2hSVowBUBRbMgk4poVzzYToATon8J1Xipcgg
EFz5OQMGQ3d6ZOhNpqdalbpJCw7IKMXFz7Ag+bpTlzBubOB2FlJw3XvvMr0GLH5p
PMFyZsNSPqj8uAQkr/4btEbiiVWhDa+g2qP/Q0JCAEaLiychECRbdQTOPHmWSV8+
2snqf7mXPKI4rWL+1WTHCtDzsDBZeEcK1Wo++EmoTK2qolEQ5DbIAmlp3QqWnDlH
Azryr60wQB7dPrYMBvJiKvZLLI083hi4Xx7WTB/0n4P+6nq2rd9PdmxsHWWYOmDf
9COZp7YJd+eqd0sZ8CKtJn2mWhTnjal2mz2ZMiosqWIws3B/FuUDg+OtNSmq7lz1
iDd8GdwX/PgHe0bBd3tW9ananjC2R6YiqZCpJU1rQ4pZHBa8YkCu9E4+Rz44bDLd
HB01/k703oXIw6W2NioUNPvss38Ak9SF4TXjSxM3dDUTmSFAAjRycnaLHu/RNfkj
o1XZDfVlnZ2Rs/oDxML/qOibVutIYnyDNzoq0m0W/A71WnunAzadBKGWHK7fBEu4
9YVdPhqoz9jV+e90Jw/8ESfRpwYpOINPGUTXaO+cB/6NPT5M/bZMtwTiElp5S2K/
/BT3h3N+jB+zuXReqNneBsPMbhAy7luFQD538ONScdY0eQkocyCHdxtj/AXTKuTX
D9tXS7Xv+CnbWeM0Bl0d4VQlK3tD0YrYyHcwPfMQWk/AyBYiUNzs9mjx8c9a7sBh
2lWNyfyymAdwIhgVUIuVMGdgfCaIfHKsYbzxg/d9ojgsNgb1xC8l2TvL44Ni9Kzq
v4UlSyooaKsK9Gj0gVAxAkwJi+IZiM6FtQ2yrUr2+XUq0hJEiB4e7BMTG8+aYu6a
4Z2hmX6LISoZ+t7vxf0rZvZuQ/CV/TwTxzOEyvN31JAeH1B65OEKC8+zJ2BSSc1E
3UklZ0ac/iD6wtPKlWHh2HvUpF9rseU0ttMGIYk3tfigUQzqgCfuDMb3vckwZSyP
h8N+hIyvK0RECgsJZCAlyOz2kSx7eh3KyY09RbYJrnI6kAvj5xxHG/Zr1qg45J9M
LqP5Um0mlje2Qx3j252n5+HuU8Hdh7bjAiFrxcBjpQuSuO1ZkoOTD4JGhX7gj2JS
2hf/RVI6QPMd+p6buJPVA1H1jNwvzeaePzcDFv5fHML/Vzcu6twYucVO39N2NVM/
tbbCZTpYNzOEAL43JZBVdNqTS7Y3WYaeOBp4YaxtLPQNtLab0lASd1O4LLCnPYxv
bMnWUHQ+1v3fOXU966bMo2+E2280JVqpKWKPAw+VAjdO8fC6eY8Yy4ev6QXveg5q
bd4mosRQxEQT7kMLbznMoNCNiQdLKyg4y7xr/QgcviGCR4evcOCpzdwqiINTG/D0
mwbkr9XjQwasJ0STfsYiGS2J//vDhCMrA4TNd4OMJfKjqpYecbSH7r7Seem0ajbR
LoNm4TNFhJUZgWcl4eAOoK5BSQJZCN2tOMUr2EDLFYdSKZ4lu+VhUw0fjFvc2NI6
agiCnxRlvidEb7kyImqBShTWW0bU+hBWCTaq64U/Wq9BDa12URARkRooJN9MV6lP
5Siq6qhNYhVDwpmEp11sVsWdrC3FfeXPaG3NBaozjBXRrYk9TL9/2dHFH9p6xoy8
W3qVBdmTMXDp9MNI9rEcE2iKhfp6/60KTiQwGwn++Ge4L5bO0Uwv2yq4C6WajEkR
9HiFDiXueoZcBv01XbloxXsnkSX8Qk8zJHxMgNUrmEYLSbiCGo/Rgh4ymmAs4ICK
hCWWfQ8Q+OsgRrw6Xa6u0G5W20HAVJpda348CGnZzyyCx/QLokGKBqJ5I8GSCS+W
Uk8T6YbOOdKxuz8qr7wj2A+SK7USU1MAGeKx4ArSHmlb9FU7J7XGX6DQvv9R5alN
PRZSICZyZjK4HtPDpZvZNxI4ChlwqIVAi5reglQ0kDh7eCE0OQfnQQRyYycbrpwK
Gb7R/m4hWJZOF0bD/zmLf3y1T3OGrK746T8gt/ETbIIm3JUvZ4LsO1zZ/f4gqpvq
ok/jH7ABTJPmtMSYT1wIbCakuFQF95xdWaUAzNzWF4Vk8QPe9PPcAn6gHFMaNuHC
A69ErfK968dYOtTr6EFHQnuEHO1tIqfwz50HybH8BbhUjP+lXtvfJtkfEm8hRJ/n
tqQyiYMmaYgpToVjw+87AVwo9GJPdioKj2GL0/1NHUB11odZZRppYgRlG6xIvbo6
HNy3BdxlcucXX7aCq2kwS7fI+NYOEfLpxhQqNGiNGDSIqKGYLPYEEAS0b6nkRJyo
FEvL6wDk/dF26DEojRCahehNjli3HU/ajRXOrtJFjCV1impUqU57xxvjVW7rKLDw
lbqAMbQ2UOepop7Hz8NrwdDUO5qRLfOSXLrZOeyfu5x59lBU8wd0aLveGmQPa7d2
AkoiyuGg/i6zpMNpGlk3Mqi3+93RrdY3dZ3cd1Dj6hZCt3NI8/qr7e2Wv9rEIt1F
8WMHF/dUQ0aG/5zP6R3gZ9wtzMPwnj0tpwKUIyYdWaw+JNmMjXfX7wOZWXQEd1Ho
3jH58SAs+u+SE9q5IOOnkMRjTUId2JPegLaihvL6mbmtl/bw7pu8CemcL3/cEStL
O7Fqip+YANoNjsiB7AuVpEwthfng1Y2JbAn2gheYkgwLli3PPLEZ2Huer/FNWfvM
hi4c0qDHlAdQV72EbMwrEuRjWkIZApyCwLRLDE5kWGCZKZ51SosWJmLoqMQYSYlv
lHpgS9cPpzRoUYz13onzcV6NnDmqV4VqwL4McO5TMcLtwTHgM9btPva7oEwzcqBE
358hewQyIw6hDdNP/j54woPFGkdLcS8lGdJ3eFMq6TCjImHrZKGD6WdzXFqa+Be3
EffR7RsOrU3m0do8Kr56Q85cHVOsJ4+pAsckSgeGYij1UnUptepFg/S+7ODjBI1N
o6WREArj01yctsUkvxAb1aR80U3JFIROArOu+VXY8trrQcPO78o7XkpPyAE2CNnu
x+DX7cuHNuYei4pf6GOb3mEfa0oLdyJ4rstAbVR/o67nDp2d0e2N3tr7+WwLES4+
FCXl0/8HVxy8PiJtKdub6UXPwMQxhMtscq0vttrpYlQk43h3JWnL4JMEmiUJ4OHU
Xcw6o0P3JcB9N06f0/Cx1avEJADOfCUTnpOH+ep/h0PzsylX1rSncFJQw2YwNT//
SaEB5rYDsWdTM3XFq8UzVfbBp6ngV5JCGTwcLW8hjjS6PhYA/1Deng1LJ6T6HS/L
0eYUr7/VzCEV1IR9KtiKi7AJ7hNF0Hp3zm23Tw6t5sezgJoArhgFlsGOV+6Qt83w
gmEZjB+0xcQm6FIRQ296RKXsSnhEt7ELtaCOlKt2lKOCkHoLvchhZ823bzIDqwt9
Cr9jTwekd//nZMUFzaXffpbt5P0DGJCecjr4pxp6mTjwTNz1jAOYnrmEmO+weee9
e1gh9Oa9ETvbiGRilydXxpMibTGeT9prY9tU6hEVHc4bSRA39Tnk4l8gO4d65UqW
xBxQP/6E6rMsW8Ck/jOAYeSNw+z0ukzm43T6UFqGR9q/G5FORTY7fIp++yeOsSxY
r5QWUIicmwAo8Gp5fXX8SNFzE/CpYjebDNuRCIs5snQTTHXW5LItoerZybI2beZd
/swiwjXVb233FILZAcqpkwhL3CwH96RG5p/ztFcx+jiVqL2x/a+9oWu6TOfnqjac
kl0YbVqDIqK8IEkFD1mbKgVh/cWCrLMV/rPVKpJxWWVuMEHf9zxYj17OhOfFlGEC
QeyKqAGD/QF76xEo7fI2qqyhJE3aijbEaDJ/WvZ51c0M7Ze8Ic1NBWwcIu1FGhv5
WCUP7ZAlBULsoeZGpWErDNv5fD3u+TH5KAT0xBdGn695T2h9o5R3bvnITQeBKmi1
9G+nLKh3SvW7NpAyGUv62R4IOFByY5F4Yt2iXGRKkcMjUxe6NOiQTj87urjaHE+H
evXeQQybcV4v+g3LW6ChDHriLLzu2l7MGLJc6RcjbH5DsZrTnr940mXNJT8xfRSY
hzDfF0lT7wpXVOIRnGMfN5olW4hWnRTU3FhYCfFB4Fqd6F1UKRHTVvfua34hdal4
+AJcf3EPZ/PpbpCQ9yA1QDh9yP+AGtyjo3RgFKbLSr+8nRTJH2Kz0Or4Nj65UAD2
Q6cv/nie7reIf0M7cCFvTEYQmoh/S33Z0YOJhiPfbLKgNrYngCQJ5O3TnQ4kTarH
AIPw7DGRoapgkDvJOmcSgv9Ihmn3J+28SjKmB2Z1wA+VpeJZ2eaWZE2weGpIyDwP
9H5CLemt/LFchrLKNhn3E+y3ZU16B19gpWm5xXEhZrUtVq10MHsiBbk8InkAdP3i
fDdKKjUvXef7F6dXQPsHVGCNGsnHHeI2OkDNiKvU8FdpTGiqIe4vnae+zXHskcvK
2t8hdomqGqXa+bn7c0kDVjQlojxsUpcyXnPTQZCCyQXG5q/jZyQgc7AvdilteM/W
YWPycAo4flGwhhdBlKgQ2tCR7TpdzOnfQ/Wv5OweRuSkPgVBrvX06ewDxZ3Lf78e
Aqp6NrCtlz2rj3ksvyGD+vjFWWTzlinPgC0UIMUoZvwKzFkYPW5sqF5w+cpIsvBJ
zk8i24wMsoDx16KJXPMYS0STciDBB8o5BObpNurrtqx9tJ1lhJ1MUgSHpyWIb7Tm
JQ8wIp4QxyWZT7T+Z4EdQGaQyXpmrRPHwarNfIsjETW13wouNa6BL5KrpIg6BSr0
c4uVuM8A5n3w3pNfPnbyDmCcPXkP7cP9BXeIeTGS+0IOq0/th8asg/O8U3ULDHrU
kaDxx2pjYvvQvn0Dp6kYMuOkGOhUGtLkQhAWAT1TCIXDC1vFadH1WGn1lTOGYcni
HcOFoTs94GedbTfGBrTi4840r3m271PMHO7NdJLkl9NSIWoyQ81NAyXVViIpoVrn
In/BbPHAQbSAATMFItPq/pgR9kiqhtaPHoDG9QTJE3IKBABBwpBhlaJqCSPgIZMT
Ux40VDMnOEajlD3OJpX1CwbN05rB7x3q4S/tPWRRz8wfnTyiZULPiu+6bhbV/w5E
7dTVP/APsVFqGTNhPQxuUqTXclo2IDhq9JXsFW17M2af5Y/dNw6yI1KA/zuMfYwq
3KXAwWCi4yMuALpYHai9hHbfKS85A6NGePrAHlP3nCeJh+YhDJCEVCO3S/39v6Lt
3b+Lq72coixWWjNBS0mNP844wnq3ePb+9gflkE42EvFD5u0l1uFkZUqm0EtJNgE5
W6xjU5lMjPP57g+P64sCpvBY7ZEozi0hYenOlBmJ5ZRcO2GroJJumu5SaiCKojHT
xQ8gFECX2PAVct92X07kHH8QY0BjIyKwW4V0tZQW8Xfl8qJylTH/sksJEibZUCLQ
DNR6xOypvxOmI+cQYO1xZ8VR7aMMLc1OfI6PrI579rO4t8PFHPFoJinARNAsEOCN
qhptsg6CitjEkzkRhOlWMId7nEnKelLCVoJjV/71jc+oyZ7pBew0CS2fPaBSLrp0
oZG5/am8CtOmq/dKkyV1iEJswyAiA5fLBO7wQfKud+WuxaXoZgow7ZnUsi+shJF+
DdeoQUAU5gxsk70eYA5ms9bFLhzCu7rltcXAsZvzBBaWu/rERqAmkduiVGsHOqYZ
8xHhbRaOHiue2KmnN/vWGudx0H+zyo51U8O++B/KPcMeb8zCrI2VlZ6C/1lp1lzt
0AVEIstix8euSYXy0NsyOx/cHUsxDY2Nsm6iTytSa4YfOw6ORBHWaeAnfBMCViVr
+3nJI1HVeSmP7B+frKyUhp4BCvnOxyTeHeJQSkZkvMvKL8HyPo3H08WFFb9oQlEa
+9vtZQRBYQszyQKDRVg/uMYoRvRkhLqOi86YHHAk1eiW+FxKm+4QuvPAS8waDmeE
rxZpPc2gJOiwhW26kMVe7/TQWeTA3wA5lqHHZeERgqnRxnuXz/uoZ9A91AlgEvhz
SqR4ZZtZZ6qSeuTpzwWhufcKoksHwOwnJN89egFDs5Uj3fBihL67mR5jQxgMcTR+
/piOIalHDDgQPXEEbKeSvZfVcl+qPSvzWpwp4zGk3+LRf3mTW8cYt1Gxxg5dK8rY
Bwv129iOWhm8YjMDX0XaQ77LJzwk2cJ17sma8LSMsyy6pE1X862qMA6ABz5QDlLo
97jB3W5BD9TVVC60RKZvIdMsLyjIVZwXDEdNlR4AeCjjU5DErk4/5XYSjq6+ceTV
ZcPMWitjo+TN/GaZp1dKfE8ahIcgaacnEbexYtWaXlWeA08bdRc6gzHqIC5yus0s
WERQW9cp5/3gWsyIQQddw6LcDRGQ72GRsYpeyCFbp/tu0UjhJnnhkyE/vVkq++bo
D2+cuR55UQHaJrZkgW44TZnyvUzF0/vhAB5j1hBXjAXoZK3qpDl3C0D5lQUyw2QG
+jqCOBtAj+O+BCQB3Ha6vuqrcMzD1aIJHh6qGEDAxewPepMiSd4lekRgPaz+9Vl2
PvCFIYtAEPr1DGPLmuQrvDoKQWfzKpRmg73pVaBcONiQeiO4ID3oxSEmtEnAxtp6
K12EWWFo1gTpK/nbmjInOG0ONFoFuNj9K2t97+7mBgA33v6wre+C3PcWvkI9mf46
aBAw7Raq+4bZtfSEM00Mu1WuZsfyh6RNFBilSkdp7aOYxEXCIg8jV9dn2oYmaA+O
fIzdwO9V7Ouzt1aSSBPOMLrpaMzu7ytHveIQs8O9K3mo6ffOUzGlxU9TmQlNpYjw
1EXebDERRzibCf9vgpmNqr1EQ3EnLNaaNXLpkpmfNWPqX7mKKhNOkuTDIbRyaexe
n6r6Pj8kRsw00r4P2veSXITWeWDQl/II32h+axfF9N+LWkmew0xTwvm0lMSDp6sS
KEY5nYL4lfunyXPyNrL237qCogWWFdDtYuMBXJdxd3byeU7OjUa6NhszAZgX5d3n
t1iyLhwENat337MuyKvHmNwBVW5MjkirKP/wOAD7cSqCf4r13vxrxvjFXyVyrsbK
fWjTsJ+OKA1/RgwX+drLeQPJyJCZAloXHbO2bjjM7+O+uu0M91pz3fIVON95lYOW
GFFLfUcPZqXPTLw3rzn8ygqOUegXDM1ysUOPrRgTgAIem3wCRvVJ8pHgbC0DjdOM
2vANX6hEdQ/MpECj+8cydNZefWHPONtMYe45G4UIZBDUjPMJsss7nWqr2m/DRP85
gdoUYZsAsC+HRI7Kx0nWxJ5vapwjjMzsfiO4RbZhkuEaoT53TmDMwzwcQZf8TiuL
+fIO4VKTKJX/1EFjQy0d2Y0Edz1qOIGDq9FcHnFnFWMB1q9ylIU9RxtEMhzlDlMH
/fios3pYJ8Osv3glgYjJUoRroPJwGSKHb0k2megVMIN3It5pIqMYLAyAqPqZ+NY4
yOGUSotSOCLZSu2DqNJ5b4x3PgumxrR4UnKNGYgRF7HqcreOhMr+T8Gi6wnRPYCl
qTshcEDgjOREVB8kJpetmqAxoIJnBa/DOtamUCAgfQ8y05pjeBEGq9jnDTDws/5B
8VOnvU1tBEdVnMfxVy27k6Csi5F/R5OiT0B9+LuhBnpEqXOgvBnK/ZClvUuNS+DL
DuaRG+DUqjITNl8mD5z00qSk6vRiciKm6JPHIsZbTtUMur95CvG8PBMypGE74hED
J5P7JOP1rsHqLl44sBu/HwLmK6zJCm4eQUSnzwXOHAbYAUP9iWGxu6/6X6+PuNZb
gc5FAoM2lBkU1fPGg6Xb1h4Se+htOT+5vgMAkuCUfImQPWTD8vCavoxrnkHyuarZ
b7PDOZXyi2CnXyiH8CBZSfEqS5fRzHBMUkPc21YP9m17nUHejiZOUXQI0BRjT3Dr
hXEptneY+g98og1KiCRI5FuQjMwCgfBELnbglffe9Q2WQjJf3W+JRO0BsuQQxQ42
W8nvk+wMJ31EL9Z+hXt00ehHO0zEQybCKx8tu0LaGXoIPQn6jP2XlQlVog8AIvbO
regc5gl6KBoz6w7BsPrPDjmqkqcJU3siW1gF36sQtQvG37XMnO280wUZpnIBwJfk
Yt4cRuEvprcosmUyiumE57QzIaigZ6JxAsGhHi2F5QId++2X97uvFG+R2PumUfOW
BkEIsC18AUpHSeMso0JF2wQEDEsWYZU9/sF9JhaFxVUg9xDUjb14+wqyT+MW3KQJ
yIH48JQFQPugaTPDOKwbySWJ+ICS4xXPI9TYyoqRHgBnc/ld/lt4S7pPbl1xgBQG
FNQKHRuCzesQ5rq5WjI67C6iORfQSqAEl67yFQxy2w2XfiuPSS2z2mZhTCNaI8VC
9RWYPcXBn05JTknolSqqd63lFILElFO0n0bi5drD9Y45nMemz6yciexgqixZA6Mc
FcPhVjsYZE5qmgmVsEgd66wGPF+Nu8SXQyGg5ZEYEtRTRUeELK4eDVv/6kW2bwTV
Sud3eYkMxhUVHdBLHjCFoWByhgvDp1Ann4smP5lyKIorc5PGudSns5znXyR0oioa
htOdn2ZvQ10buDOatS2PvC56bphkBlloKvtU1rzkNtT+JxvVZooiXsm136s7u0ZY
aWFdB9cLt6aWGJqzZ7U07vOGAjVdXq5YEehPLi9q585n7O0ArJOgehxbz5UKDKzc
1D/9PVJbxr6nCjrr8WS9tgJL833ER3KkiG4s3H2MriZrGPUwvt2D0NVBVVvoPeKH
ohDDSnjyeCVAKK5DGaKQuqDQn8JNzRVIDzQmGJXnQdK2cnlFQnIPftqel2a17+la
sjZqYV+qn4LB8dGwKW7UBoXU1pHmFY8aklEsWFPpXPolp1Oqn1/MoP0ERNmW8ofF
JgWdh1WLmy0o5fMcE397oSt7FW6iAhlS4caYuajVQt4HZ3aO0inFmkRkn2WNf0Ck
2cfFPkBf6GQtN2TolPkbigSOyOPno00jqmmmuvJuJxBM/3vg7GOPV6VLMEnI1OF3
hDEYtgfIDrtkndhwq5uiDP8o/83j4+g0dKGsq/8pTVuQKB58eAFXyYdQ78VRjEiv
PIhVAf4PZNLdDU4W+UCZYJoQHI4NQ8H00lzJNANuSZMbVpAGofHv4oJ7nBTSKeRM
YqTUfvShvjkRK1b6i92X1fRTgFZWjfJMZl5VPQoKhTgFCwjTqtcYHrbr49kQ4pDl
lwo3MGJTJ13ovtiZ+9r++lhPuTZ9UxsGm3e1khoQaNVRmevp8MLhQnA05MQdTv5n
s88Y+iSezVM52oqGhW9iW95VJG5t5gIWr6jH/++Vwyqoi+paNlznaptestDzpG/p
C99HMnjnKK7KO78JJi1dSEnKdmsVxv+7JJ8FajSP9OJ6WUEqtWAD1fyrnLSXssHO
9b5Hy1k3FYgmVb29cNevaDfKyJs2hthxc2rkhwmrxdYY74azsnd7Ls64lZ49D7Z8
34Si/Fgkak9iixJZjNlpufYbkM5oiJaJD/A856I7JNEq6BBtKvy3DPxrrjPMbuiH
u/89dZV4vFAXK6GNq4UV4A7CPfdsd73r2TUSmNa/J8KugLDhcgp/IZQT1It+PGt+
UBDrnQfewtWq3XpLfGueB1NZfdjCTppXjLo7vYBDgPiCRzWkw/ww6RLzmXfwiEOU
byiA8orygxtnBSSjexcBDJxXsT7gvc+vpPtmVc20oRKwQz77VIA8mVsWYxPv5sLb
ThYOV/ZRTvqd4GoXnsQXatpJ70GEKOxTH0l1gjidWFInOPi3iinYrkezqNkMOIno
KmPtsuXN9mTbut9fkzfGAH+e2BlCgZAw+HtXzOsqxv+1xgbF2HoBA9Ux7jqoqvKt
nNTfjOWOKwQrskKHeNM3TkJpLMdTwtpEkidFE0m5jaJiq/cCl8BdtUR8yG8d9Cz+
+i6/k0mPQ+wflfP8/fTmWN/obJhPOEYEEYd7nzp9EOiAhfkql1qgowAGudcS1HdR
HvdCrj7ldcu5q6ZBc5OSWMA4TL+TEItLYIk1ni/VtoTR8EC3FDvr/mSsynvbvGMs
+iAslKqxN+QWnl6DvVryqx5w5y+SsqZ+SMolBkrozNfeSjSboaz4nEqhL3u0k00j
zDqBA7sRGLx5tbHaHoLEYbheAGY6cBU3E8lCEYxYFXT5yJt7IYcAN1B9INYDzvFU
hvkJzS17T27FaKuH56dsy22SNpspZLYARUCsKZ8bBApcJAeYD0P9PFYdp6reSlVI
cvDUOklRsfHkehM7VcTaJ16HUF/Ko/UA6ORSWeccOW9IJwGNEI+HzkL1wuwu+K0C
s2WJgCp5W27rY+CbqNvQS42r4PqCCBsfxc661yxnN+RlyQ7bNuYvwRwn6/T/ugr7
0+RQtVxX+a3A0wuGYnccUeeS8bM5jZHkk82XK+i8pAmhUsSAu43TGm2Sqjz9vx3I
HeVi53yGSZsHcRqG8BlX5tAwz7WCBUK2rPu6pnw6Ye4HuK8XTqHfAoZ6jK9Zql+U
NAms1njik5WPUYQzN6hxioIRGetIxxu9rVsaWeKZvJcUnC3qig4lItT7asT1UB6B
kYQgwoDmfR4Ltqj1YmJJtEbP0tWyKJNiNNk9SOZeduBOj+tUVrPnLuNkVdL6w/W1
+RxXF0HOdL+YYZFsnFI65xxcYKdcp0y9dM3Fv1nRenlzfd42IuLkttHR2jHGuvHF
BWlQeuiz/AifxrzcKcnP51mWmohQiPWvVfmxyEjSAucCCJVmgAjRP4sV9WuoDsUH
0gamzij1CuW8Q1ycivcXh1xcbjgZCHC7jLFtQJ2ly3mkG1M+HMjF4XEWdO8IIeME
Zt3NTq9CpFHtJ+SjmYWCiv7lls39RnwQrTUtDiZW7JTO6N8eIgWDjnrskdB/vnJw
Nl4j6D/1qM+9iwieMfjJ2gYrXfR66bwBcJHsT3JSHQesTMJacdUKNdFpvg7hX+JM
v2iF0stXlKlReKZ/FPHA0oJ9szsDX02Y5jOLFhirNeWMpdmof9o7Qlp4kUeTf0By
OXMgAQVeVpMRdlCJO+a/yQnhPwpMGoyyeuW4IqfYcF3kpK8vskGHDnmQfurNp9Vy
cdaH9Usduu8umBtoB4U2ttYugHf1qYwc8vnzM7XQEj9s/twsbaH6grq1w6nCoUxf
V4ZkiqGW3BlEWBP15L76mSZv05/n4eUqPK8AkXY+eFV/olj9TapcYDi7N9/Hvwdl
4cZ6e7Z8oMsse4dQfj8WHsoig5t+And1xgnF/B4EzKtUoLjnNCMMclU/kg3e5K23
ATnaa/gThMU5BqmeoRxCi663NjuFvIPF1ZyFS9FGHWr6YvqkNPtmA4k9WJ4fSZmf
22VRrxcZihO9yDeyJt4t3NcuIyu/5uSGgHkFIvxPV7vblG+soCs6iP3+REW56udk
GkrXs/AJQdXs/ws0LkWhPKaJcdnLyk26FbHb2KQ7ZxBAhR9KZFQNSNs3QgW7WyHy
ab/SIB0S6qQDOOal72CcvHPMoKmCGNnfFRdgSZ9N2FaT5uYCbLuqgHMXcABdlIvN
pFSu4YEyWpT6SClvvlQN86mH4W0I+NOJHENjDI+dUV07ZjCkuDBvtkv4sz66hjiw
mvBFU1SB8bAChjOHLmpoIJMRImP7k+Brkx+k2HNK2mT5ZzOlIJxlfrAFWAokfq18
POSF/DNj+UpCVc4EJ1tu94gLFmc89N5n7vZ3yu4FhhTqy50s+Ydb3QmBLGLDqazY
Dg8oBFkhlQs0yFXQweBA7iS1CDki4ODIE7lOad312krtctdnkJPKS2+ffZf/9b3E
PqGSgee0lsTayj+J7CRJMc7DlQjHuE0n9Aofezzwjmpry6/uElmIN9Mp+foBtCL8
ctcx55T0+IYhbvUqKoQmdMo10gS5wbVVwUyOJxSkyO3mjuWjmjP6KBug9zdyeDAv
eDKAYQ34rwixtqs2DmvVVCcv6OtTnHggOVG0cfX7H+RoUj7E6mtADizCVt1nxjL7
4vWM1Hkz2qRzErnYpgU4ShcIvSIK9Ksl11lqIaDqkLW1lYtcXl8h+Yx9SPe8/VHN
igKXBXXeXQrqeOuSdUyGM2uGlDqk+FgBw1wFpwXOgGGugHZau8i///fW1c39+5pE
6O3wM/BsyrmgCWdz6XcL7V+Qt2IbglU8ZFtpP4cONx/XoQ9XkuA4SwwG+/5RKBos
+Ek7pyEmJmiGeknQoOBr9Dsz3KIdOUDCgexxOHUudxJOI/XRwCea6GQIAapogM3z
KplClegStSwDkztrkFBrsju2LQjq/K1siCJjgf6uvS/pATSZb1yBREPRU08BUsXi
F7OKoTR7LM8TphO5A4nd9Eq/PwyXZE9LP75EVqJk9OygmYdSlzm3xLhBHb1SKftZ
dldCMWGgWz3r/09Y1/4foaNshCSSQnbkMBdHVrkR3SOWvUwoYeJ6nTtw0jxGgr1O
A6ZXvUh/uGeAm//k54i1+5hlODGqkzLkDoX9i30LL8Ct6vJrzQlp5KiajWSefLjp
Ju1+QEQp/0FQudpOX0eV0XhGt7Cf7UX3jIelUfhaL5AbO5MaXetlDeXd6qJLPHWT
RLNZgyxy/DQm0U50z/i1azGYJoufBKsny5lfyHCaazHIduEZlCtRPQ4za4kabxN5
YezXA2x0U4C9+B1Pqzy4/vP9RsqRKwCGrRw6G4a8JIv+9Ey3eKgrl+83loILo7o1
FZjn7qmOfimoGm9OcK8LdUt7WrSOEiYywEwLt++bLyGVx5oelnHrDg//6qIgG772
3D5/QEh4+zin8BLyU0V0GijRguGYAjbf2UnI5Y71xTzVw2NxU6eSuRw4h01h8Yo2
O2mkZ6C1FpNFKeCzhG3Re5cD27hu2Po6kKnjwAmHBpjGt9dlzUau5i2G1v6bpNkX
VWOVxCKLFEnl1GeJV9nXZyPmUE7X+H/9hbT0RlmFc+2yFUBpCuPSJzmuUmFXcpog
DFnO0QBsgPK+FcXhFND+x1DUg9yEXNG6eXULhHwOKsUvKMnlbC367Tlz0Y+cZp5x
XqePgs2QgeCpoTDxm2yrazQx4e1H3NOyBGDfheb0TTCSdVrA8EZg7DJ/vPorPEKU
DSu07LeacfKnQTNSwvnugX+rRzldtDsL6WNQvryrSNcNxz3YIhfnvSutLOe86oH7
kmGPffU9XfKCLUMT5MXA3uZ/ybqZlYO85jwu6wXufdawj59yomdr7L8EsDStgS39
wcXivU+jlRfs0RI05fi8juNpBjdnIf9nbqHfVgnOuW4Yd2mp675sa5Oq+vEq/d3P
OZ4XkcoHZryD33WuwKHMWUH9cMcWaF+PgNt87FNjIKT7inDvLjvg1X1XdP+goY4P
sOekberKh5Nb2houn8YvpY/T+Lp7zjQ4vg2BC4XW+i5T0d/vqvtbaI7Z8U0H1MGq
4e+MD1vMSDeOnEKsZx1Ny96ENZPRAfYyHK/lLYikLUgMBZtyC4Fxbg8vo3sxcoQa
DgUUXiaK6fB21rE6QgidEk5LG4Gcs3AjSiGZgVzz3BHnQJj2ePgOTfrykCwA2MgQ
R7URgd3lhuYa32tFW1GUme4D19ok+JpFPlirxeh6LArdGB2Q3EQ1jCC+mzmXIOhH
Qowt5gUvsF0VnEOM8Pgp6XM67o026WICYCpFjAhta4oUWUTaqCHI2pYeAbaNmoRH
wp4H122KAUOD23GoRK7AA9aT1XdZzC92aqyoDH8NPimPnDoy4Vb2wxs3skLlygfi
0dMVg5zhe7PCN0YaFQnzEVAM238zj7mzc252YUys9m5xitJ9rKEM/YZYWbNZf2TS
ZK7APTopCFlDp9LZMG9/XGqmpJ1SYnxSzSQ4hcFSk0CM0T9LZ+9Detp56UUactTk
BPqd1xzvfvt+s5ApIvlOCIjDWiVYtZBbl4Sa7GqNfnXRgeiCqflhl3+o9i+jDzQy
nq9yGVilNrVq1UXlD6H1EEpxbB8/eiYazlRZ4VvtdVWjvtoeRyY0jjqMTNWmYxtr
0ouqjXQygRtDCcFES+XTikIDN/G/BYl4Im5iNXnLMI8r3iQ6nHoEOSTXMxmfstiU
A8CZJn3REcn1qhR4Yl+CsP2a12jMA2dWhzQfFpnJJ6UbqUBqb3BZNIpny3e1zCJF
Eic1jKhxV2Dc9fGNrBny9ZgvqDc4P8hzy1tSGYAU9mVtdr8QIgph+/NudGJEQ96W
zCRbe8kxmNFsevLK0uUzYexwPZyaxCRNkrjuAXMazL7nfNtZuuF1bJVVaTM3jux7
ocxR5MAochlPxDQGk/67pXVgLeOMaz8kjwKWHnPS5KBydDVjoT8Qr4o3XQFuh/ey
NwfeQ9HFBFp6HWhUXU2R6b2B6fBg22HyqyYMvMS0cyaorqSEriQk/8p514L698HP
EWk9aRKz6Nw4MdOg9lfMLcYcg8jQru6di6hLW1ZbATcivG9DVriZ+MA0cPVJeovd
BTX6eAwom1zDK/7hA63dFj4scSRsBobFb3oQ3M/1pqI0GhKqSl4PnK6BnPMlzmZF
sJRjOYBIJCah8ek6ndDBZtUIC/2eyrhxbPA8MbvL4YPL+bXjFjnLCP0hAkoHUr+v
xS4rcByPY4Gt+Xbva7Rapb9ql2w9X7rhguG/Zbr+kuBq52+RjM389LjcWyXW8VdQ
KY+YY509bH8HsEus2F7goS8nYJgjb3kYCK5IzLDgp6nsAphIh2tdRHU5JaQtcdUv
ox/yLlVeguiDLkzzO+/sIoKngXLh0pS7ofnjN0d2ImJWQx/O2CdFbOHE7C/Iy+dg
4jrmexiPDs1c1fJBt2lQe1SytT1IJOV2596b2iwqjFEg6qlaZ2ViL8lxhiLT7iGk
J3Ch2UAIMxXXi4IAr0lzj6iiDjtwKrKNAR+VkrNHrTksztm1tWP1kUQfLf3+Ecct
3P9UFoosLz6j0u7rFD7xZsfKVXi2OtXrcyf4TJM4677dtHOsiKTOEJtJDOePUPp/
Vxf00B6y3+kYaavtNGHquDmB9Bbdfg3yVhVV04wEQ5kUaVJDrg74w4KFOEScAR2K
8flIzauf2C0D4/D9pLg2bqP9j7R0O9Hm3/P9gSjnEC9AQH8ns+IAWOisidHWsPZs
ZG0O25BoPWcIvvy3qctLLMWHkd47pA7uvxIYV/maQ/nBYu3zA2HFwZl8KRw9vLh0
WaI7dIj9v23E4aWRvGeD8X03rUWbwaxfz/WfBnRe178tL96LBKwvuffWcptC9VJU
1D9vDiAJBxTnqV9TO4dnw9PGL9Uhi1SQwCiyurm15sdvNKHA9BpFHCWzF4nPMGHl
IZm9XWR/9vtsgy7fcIj2ciC9fWpuEXvFt6bU+rkgY0ouqkThYraAGutZ+G8xEoig
tWRmx6GrEeP1Q7xEbXfoq2sMiWpnua9kslrL/7OVkFYOYA6yR85Cs2ksMaYuIMaF
`protect END_PROTECTED
