`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kmJ/ZpcFotfliyuTzhA84P/jhuYTSksoKhnr+0QOO1kDwAAc9yetSxlFmHy8qbnD
bW9NBtXBbrBkW24iXeyKT7qq/5SDkeptvQMoJ97QOQlDhykWH9DiQ2Q9ZtAV3thI
gTg+578dkqGzM9YIiWEKmJFq8c/6FCGQdh1Uq0umZhBKQxu1fXz3dlrjMsrwAUf1
MzMu4mtwT/E6xj5L1ZKLz/kZ4RpowOYK3hGOq09/tXwuTy158EVL02PojTFT4PVl
eE2SY+PZAtRIAuoowbPcqA==
`protect END_PROTECTED
