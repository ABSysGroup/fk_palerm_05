`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iGjaPgD+w7cKEzKttK7hVndPBFsDhtzu8+lhzwCsVUdKX68SeAy4wdM/oS4Iwmr/
vx3XS1F/aiuAVUwSErgUZwkfoJlKRJ+WxT4DR+NUsarS8H59uaPwwHnBfXp6h3Ob
O8o6b5fuk0NJBylJChZjLEU7hazPcrOQEBXKEvTMEvXAARHrO8LEGrwCxltklu6s
ICBFITdd9+aICvPPGNgtwRFjkKrT5KgbdBQLXwHwE05io49TKc6txraXJyYGAr49
4QYDpJMGJ6Ta3th2+jiJ3c/x4l3djVGPwNdO/XjQP4IYKAj3nkTlS7BqKgL8JWnA
`protect END_PROTECTED
