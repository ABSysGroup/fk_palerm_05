`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0jie5W/JGQPQK3TrkUPSopv7jDqwi0qA5iWhPbHE3dcQ12P9kxjex87WuoDCLt/D
VX3jvc7LNHic/lsTRmiYiUuC99ozf+0tu7h88P7mP64IoYGkuUMnp8vHFQNBQ+ch
48ofYMqbkQoGZVf2fKK7a9XMQGWpEY/3W6H9Ay2spNc3kNs7gGKNjLd55KkU7evk
VyZYJ+pYXOgGsLYDB+Ta0XQa9K4v2KyoXNlBWrt5BLBvxLYV6Cin5vUcey8jRNIj
t2j9kCzFVUMj3Be70XANKzTylqUD/VyRpS/hEPSKiSYMbVbDzWhREnxRn8EpdxPy
+c+6x8eSfB6nNuJMaB3cLJDxtrQEbXOVwzRXHNV13u3jTfEnR6Dlh9FsmHqvuzKF
ekGhbz9qAbvHfS9OCD8GD7a/1+VuRgwedyB71wySzkOISNXs1IPdZrC1vcC2E3r8
hmGuMAKSunZkPlDCFRZ43f+u0fA0NL0XY49MxBn03fPdydtwebLwVqhQOZyLL+X2
bFs/29Cd4icFt8kEC87NxpnBeZQQss06VVlCOg0jJex4gntc3dSMGqManxL9Iv+5
hQ/Ld7eye+N8CbwwQ1QTCMNTBohnaCPxtpsfeJTobLL4kQ9d4MAf7Oj5wWk4RD16
0KYDTnnoPu0ZpiDtfSZVefgPh2blbQqvFiRY3qyCdgE5XH9VoZRVqityUcvD7iW2
3+wQuvWxAa/BWEsgXghLHoKqpzcmf2ZAWzOExUdqlRZ88eAEHUHn5PJub4tpE3pc
yHVEKZOAP2RD4EIRC/zcse4zIaI+YgfxsD6jrNppKFMy9DLp+Je1H5gzFybHKMQY
3M/b+CKfwMMUV8f2JRkNzL6Dx/j5K/28FqILjH95xVUlDvmHTsKCrjl5i7jfpDlg
qniz1/K3czefAlCDgurEGo+aMkXP3qJOo6N8v9LWKGUN2EjC0PBz11njr8kTXJMn
iMnJwUZolQtOnQzqnSCzuBJlsV6rnDVgdj0wtAKTg18B0Azp69gAJb2J+VsMzCOV
`protect END_PROTECTED
