`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fFdxkryvMr3EKnBWfl2vWm3NhRQwQSJYGx7v1REfFp8ioLJDAPmjkd6p+4RVQpkv
WgwkWh3GvzWQeI2F1vLe+LFZAuBBC8r8nZvQ+ncC2FF1m+NzgzVRFmxNc2TxzVR9
Bjysmr+zG+//vqDiSnWhsCGrWs55muHOQ7xQWxBrLap/k6Sefn73aqFjT5sNyLuq
TRx5yK8aUA2yoBJumjpborjTfCfhNXdHbaI0TorKZw/KcuvH5RzXLe2ZoXYk9N3F
rlC9foaLX3HOPGIBEDvixm8PEGE4D8ajJGF9WjNPexn2Nr8H8OEkUPLPfBkTvbW9
LDn6C4uH6E/v8qf8NLkxgPJ1In2NVigdnacWaq62S6BR1Lo3DGa1u75DrIg8h4zV
B9blwyFD2BJxHHrXztohllpA3WMDe/GP6sIx/zWdFqrMWs6FPC4enDtwTv4apqZB
BRnmdHIqsNnS4HakSnnwoQ8/lc9RNVNmYJbyhi358Tf8DZb21hIysA2RxOFKXpT3
7ORsMSZqVvJ+wYky3ObIuVL9t0jP9IoscEh5yu6jbQM6H28C8HLc85ptCu64i05a
vYeFJcgsB+gpItqOSsOCD8WqwyVmM7vKCqaVHUioetX2EEf4ybkNXQ7DEA/IMFM3
MSOfh8CFICJs8NX9gK7rsznvR0ZzIAhT8JuWyqy+WEgFS9JQGOEipeIbgGgV8nRR
nHx45QGfAGNRY94TFj/oM1nuTwiixex7FP1r3TgXA6y8bzGC1ah6fLA/wR+yVHR8
IoHy/fvEZKfqAI7a2amEVdMuXkeLNl1B21pZqvPze/J3vURyveVDZmdBzvmKxxm2
eU6P1jO7ej2AHqerJBHEAdPBWf/dBy3lDGkXB9ZOEArs2yn0PvTpNq2bbU3nu3rG
zJKwiWvZuw5K7PHcZwANnxWkpyZJlRyRhWGMSx9ZMuYn388rWZL9zQA2wh4iI1bw
`protect END_PROTECTED
