`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D81rGYbnN79wHaq43+RulS8PT2jvGtOtkPaCZOsmqwnzpJbFC3Ab5j8F00l+TjSh
XbkNrdhkDZaubU38SLxmI67Ardl9XeEkWn8NYGFqZy9wwvohcbL88TKeFiBofhA1
9H/gBK48k3Z2dBdaD/PZAbvjx2tbYDlojqEVVCwE56iJT92DO0JrtXsR3PhPTiyG
Ay1C+aCFzdlihZ0XNvDw/XQQ52qTb6Zas2Ya67lkEIFzuAocf9040+sz1k6IAu0N
FoMe9DkLRErjzCavMDVeag==
`protect END_PROTECTED
