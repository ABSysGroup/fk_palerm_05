`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4y9Vd8P+MNi5MsVhsylltC+NPxlThG/lWrgVtMc2ovxruopeDhGSuFTaFTXvRxup
ntakWsIN0acEn7v1LflcVTIeXGF5NEcLaw7oA1O6nfRR8HuxCMkTjqMqdKkXuKSf
dEx/YeHkyEyeodtUaPSx+dO1NpyVvuGvfIIYbIxfAMCdeMl0GD6d/S4YDzQmCX9y
0KBgsBBrlDS2ZfwF+OuN/1rbAUcyrZTeRkzw2GcvrqMyEf39oIN+Z6HQApcj2tWo
F54241YCNXGTTC1kzYhpljS47Rx3YZpNuJxVHQrNl7sjaWtWobiZjPJsxuJDu9as
YjgsDJd/WlUB7MRVoZWvfNdgGdPWHpgPxvpr6YruQGJvqW88R2kcfgWhoGq/9hK/
bkXFL0SCxKB1UFhdTpYwC6Q/Ssi39Z/6mpGSWjm5sYkJh5JPktG2rFXdXQbpDALz
qVjfAlKM1cUXB1zA+009Yct2Et0IVdhwDybnZ0VYx/lYG1Oi+umJ7zbOpSI9Pmmy
5IxgRO9c47FFJl1VElyqP8XzNPKQILA77EzdtEe4mRIUU8S3j8719Yozy8cI1jtP
PhqhJleBcd5hOhAkCLzZ78McT4I91T1scX8zdo92PP9JU3imflCoBzKcD7kVrFAl
GZHqjJhtdxjsLka49jeOFhGQlj2lk9brZplQ/ODilHZQk9NWouSfhBwr9eIvEGbF
RYurcxu+jrvAmLTIEPw+A9F7l/coWChe2g1YBQkrY9Vz9mCYrH/RMJl8t8ysAqbz
s9yYSR/Keegt2J2ai7qWObbsKZFKwvwrU2hCWkfQ0xv/Uurxayh6gxGpaWYGJEYI
zWNX3e4nrSFq/RRJQ7IGWpUGn6To/yK2SsNWcRnG8K1B/62SGseh95nSeyoCsLU3
gGXj+irKlleQER30cAHCJh8m62oyvrZmm4ygj5AprrbY178uHI4qE4zNh2qAe4vh
jA9xoQKlx3EmXlc9Wb2LcI1einMRCBSGPmMl832UFNqvsNDSNEcPQ9nxlxM89r6t
9bKfZ4QUQF0XjYCRKubBQKJqbNqnuPLtVwNeQcz9YqgasDq7fSEpEbdCRm5mUHGf
LgSmQW8SDWOpR8gaJ1bigzHsydNmIB76crNerERD63nuxZCE43Ww64qStkUF5smh
ecELaM63eqnQ9UZHTGqgSlKltg+xnhmZAgy8NrrHHRSqxY6pmrreu1FD/p+XPZV3
VBZQxni6caDsAHr4Z/5zZwMNv1JHWRZjecargPnre3232kSUCqLU/BhiMmSkgsXV
IJf9j9bto6xW1iVEOhnW922AscC/JcYhY6FmNllUWhnG1sjfuLZvi806bm7FWb3R
4dL1DhI0zKJLblYMEqsNOWgT4Gj4Bzbul0hMHqx4v+tBxItY3iveyghA7fnV55q4
pAgXabqfdLDie6DWUxPcg+mnCJykQLOUz+lqWyloVdA8WB/Jp/V9rqwnBUvtfhGh
rFMtwqY/JirN2lPHKAniHhr7rYJ2xtO8T0snDcI8Du9J5vv1CrW3C1430WbymhwH
oYD0oB+Y2ZiOXaJ1o83XFeVb/M6w8c64+yil58y8ykXbsIh4B7lofBzPWfuN38lA
V7k3ePZqOmGZpl5w+lff7JNOnw1GaaGYbev90S+yREroJBB1iJsvW4XLgCeJ11LO
EFtZ+lMwXgafUBMNStFeXmn94aDkm4FN5nF1hEG2O1ELTzNp4lYl4HmfPnuJBSQE
VWnSt0i2K4oQqovlGpQNeAJDP6LDnuzjxQ1ySgszZS3DWNhqj1SFI6P8qegvoxWd
Yc3N6lpu38SsMxf285ny3JjlXmthYYtardBP5rcC+K/OBTCqZM1fILFJz1c3xxbm
ggkgT8Rbciu/7lN+WIP9hcICDnkHs7qiiDs5ylOuW/vHDUQbzW/PjAe3Na2P05UK
4StGZFZ256wncThiwjNxyWciS2ZRrMLbUk1FLD+pBMwdZKJrY73DjurBVwBQLbwD
i03Nc02JZUACQ92OMYHjv7DWRxLfwahzz9ZbogknTrRC7sO32nCnnPox9/EidlVT
krBJTT0n2f4LS7Y91M7p2ayoLw8V0QuqoHwqMfyBk7k7LoWwAX5CGvD1aApy5gBk
+pEx1Bc2CWaCVD/8+P61NJS95dvr/ho/TNLDOPUhgLD2odzmcDuP+ZhfS+B8wIwj
B3Kkl63EVbAROurOgJmeMnN4VNDXGhBlcRgekRtTCccjiT+YjTqtzuGeqhnDCmjp
2/6Sx3QM8DQf3mCkgJDiqSMSw9jw6Yj4KmHUk2NLc5902RUjHdOA+HcszgSyRpY9
`protect END_PROTECTED
