`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o3bVWT9U1+R/Yntutx9fGyFB1k2d3jiEPq05Edlk7u6K5Agj0tmrQAvvyECdekum
cxmHNpDH33edOS7FqXHJTawMasPYSb7RXkQzHBbUi+JGVk7DoQQR11842V4nbRBa
rCYhztaNSQTvk7hGZJw88vcd8qLxO8feeiUR22GKPwpsrFp0i0eu502wWc2gbvMu
+zetx/omyBfIOIBdX6YrvWf5LfTJyQFZk2/OC7Ej/pt65mdq2IwlzeyPokfKnwts
gUQEN/h+6MdQDW/LK1ZHmKRePnNKooOTtMgORFrJrRoDj68ar0df6ij9kjNWMB/F
LSEVSggoas9U3umIPlD4ZoQDw+NxJj1paCw08Jfbp5/uRO4Obv15QVzZOfTP0WED
HtPIbiIyGetp3H/mgomTvlXjAyaLl6giBTIvZjs6uqh0T+Hi+0M9fB3kwS37ihfT
bHxA0u2mGPE/lw6Sh0qFxv1GaJ10T3DP2Sw7mlw/p9oD+a1jiXyA+zzmZkceEh2R
hM1kaBDlPYls8ULJTABqhZV7/SQmqK7LZMiIPwjCWd5gvBzioIopnYDmnF/OsgzY
`protect END_PROTECTED
