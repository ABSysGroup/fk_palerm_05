`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AmmyNM1n+gP8E62xRou9s82QEJbdk3JdlnZXmemZs4i4fPgKrySY7K8bxU4Lc+0j
I6XxroQ4Lf5pw/avLpifNgVq0Y7yeXSyFMrBCbFgE35WdlEqHSHAMGmmqChkM9pj
Hc8xd5VuH2kFRATmTIfb35o9ueQKSALuy8fk2NX1VaNeWJg3I0+6QtbrZRHY5gOX
XMS7IWDWdYKIa0xf2GIp41tXrH1qHzZ6nA0H3bKamAhbPOijZDWJ5GiMp41FA4fi
lH/JrBO6l5T2lZyTWOM3e+LJqJ5j0UiAJv/dzmCo6hX9ihHIJNjQr8otbpGBERti
xVmLySleyFY2rGot7Pt1hSgKvlJHOPt0wBaKPn9wkTmf9VdpfG5Nddga6YHLwLHd
GpHf8RS++7YEPAhFt9KlJm8G84HjaVl2kl/MSPvwVhDdj9luDmBfYm48iqclxRpW
Kxtms/C02XTDF+SqVU7a5s2a3vr353hGaKPvPYi3UlXOT5h/So3CNNcE6Z+MYydq
boSRGTQnnbM+ZBW6klgT8kH4aoq2wgAXubj4nu/p8up5Mpwtop7+seruQElS2kbZ
ddHbSGisTbeIm6xW6jv4z7t2azZIHgPcVtXQYzE3cnibF0o/KDS/xWF3BaoWM/5J
cNz1p9YVF+q3h+ZoarLIGg==
`protect END_PROTECTED
