`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/XTkNQ6wcdlrmvhHwANJFwCDkst1kLGythkxwz8RPQ0UW6Vadcm3Z3cwLFOqgaE7
hWlPP7jjUya1DQJsYXHI8jN+/S0SYkW9z7FwR+QbW4bHZG9bOq51wQc3tq6PBDDI
scfU9PjImqRSiSUGyAYoiY7lFNMF4tKNHnr5xhXr/tacWCXp1AM8cDfzkhygw/eS
SzCdUCK2XhGP91UB4Yt+/15/0mNfVxGGL7g2Vt4raGiDtfVrQrZKGQG9268Q0Mkm
bc3HYSwu/rmGnwGvS/8dAGEhjNOdEoTDC0GFg+rm0EQWNi0cjyPEQ8sNw7kFGpa8
KN3vUIUrPn1xAHgI8tBSXarAiVPmozj71bFQowUKcY76BaGasSjrVocrQmeczgd0
KT+d7EiiAGV71yb1H3TlIhOQ5lronE4B4zSf6XOALVxL/AGA7Oeqs1KIWwNhmc7X
aVZh+jVwr9sY2EreGFTl0U5it5Q8gvM140jpCxe1ksEFfETFcXdxoJr9SjbOy51y
fmc9eCRgeLA0Y2LhRCfn0h3Uvvwbq+vcDmR7vP6mRsuUT2Qm/tXVy3uvFX9PvLig
EVa8cqXGyHFtFDX+NlLRh5hsJZhx1d+IpjcfDagvZq1J3GHiPilIaLB6Wqx4KTuQ
OoAtMxl8a7rQQNsmt6z6YisOX0RSUYrZzodMdD7nPDQm3eIRSKDgUVuOFyS+bxNf
bgG12wTSCo+52PAqTymO3jpgYya1fWUOTDJfpcR3sP81tWojTqplqpL74JmP/NMt
olu+TrsirJ5FLC+aEGscANepbs3sMReKMB+6dZMuOKrfcFWcFTq8A/cnqRweqv5y
xoaq5N5Kt85Llt4BOP3o9gwoPC95NZh2fipdjaHzA+cEirZKp96+qlHrqvY5z2rb
`protect END_PROTECTED
