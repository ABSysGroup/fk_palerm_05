`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BMDCjrB+CTyiDHb6USRbfJH1FGCmyXrWYDv2UL+QZK/kxk8UQ55ChFWVDDd495ly
UOADZze5leE6aEf/6lku+NPst8G4qwCHbQT2t2vQ6yhsgaPbk5tvgZoaLMPBWJ6O
f3xTm0hinz7vnlp3BjM64x8OPSCGD93dbS+Mp12j4H2EXPsVmD3jsKFljURYLwEZ
2wMQgY3nAFlx3+24sk9ZPgL4OpFom0HVrsXMrXbfF9oS+eOmQjeeW0ulKHoAv9k9
8tTGiFs1whqCJvMeqU4XQuy0YzSFcy/hbjeN/IIMGUnaxbPiWwEGE+qvEuL//ZP2
96UG88cDRLihCMD3+AfVZXX5w+i1Pe1XlEF7aeXUXBOy9HTSeoUPu7PcXCnawiH0
yyEgWKo4YehqFuwYTiY8uQGUQ5V4Jbjx+6/2DdLOzJvtOYkP+7UOk/yH7SirRS55
Znrey3YFqcGLvVCHXyW3KQ==
`protect END_PROTECTED
