`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bCiSpXtQdxl2RDotBrYGxRgvlM0eGWNeZKYkAkUPE1YAWmX8tk3Sk1Csw9DUC0p6
ibHz9dNLIUmubf2PG8MKrQqvLMdGSZSOy6ekMqm10QjjxwfDhEBs1rAWKeg+C/02
wKJcWN0uB9FwdLVgaXD3DPr5SsefEclHunxE87/Bzl4PyfpSwKgbgxSmMZUJWHcj
J7r91TGHRPDQPgprQNq5ffR2dDE2K1b+YWvqY24ytHeGXgpF6dcpKb4RSkwrgKV3
`protect END_PROTECTED
