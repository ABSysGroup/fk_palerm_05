`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aT82F+0k08tBVXMkF3bsLXJjuVmakNgYUhsXmstf4+vAfQLxJt5AKpA4l6nWv+yq
0qsp/Vbk1b4D4wqN5T7dNsUwZTC75Rd6RrZhN9VPnjt2BbdWPam6aLHM+0EubJq9
ZJAZhDmnxPcJWIq32jQCGZEtEbFF7EOokP7SIUwyS3sTQ/dbYUZsfomL0H4MWnog
80uXymMlXUtDWc8ppLNf8Wu3IZH6K3q6Xr9GjgHYpW9Hj2/Z3SvkzFSTsTpvtXXY
SNprzDwnnkHPaHFymFBC+a0p0NyPWGv8NJwlih8LpYgO9UFlrVmwbVHXdHLLoUEG
mt8Pqpq8nhEz26QbvLAmteWPHOmgiKl85M0IBMjdz4dPRi7pKkuv/h4SRnHqBOK5
RVwaSOe61OMgNnZ2lDZoReQ5XcbUiHw3601JGNYBvupTSB3/tr3rR1z8J+ztLnjh
JypQE5yQt2j5VaH8vJCWibQXOqNYv99+q2Os/ooIM2I6Vd/x2aoOS/Zo1U1Oq3iK
H0BA0VwO9GD8r5Ud67z5axNM2nQDzyXOaSFmLnae+xQ5F8QU7C2Rn40uWx2AOrMa
sYefgXBIe6As5CpRLCn24FY+C3VJYdzkTDm0d00kgVbTF2Xkc4exU4OphQqgfuMJ
WQEGKpK6gQj5EPJK8uaPXaEEadQQVK7yy8cokGYw5fkgaRNMb6V9Ou+CGMUcRWCU
7kCkauZAZnIofO7Tucj43w==
`protect END_PROTECTED
