`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nnE+FSpP/qz5g13RCPnd2vX2v9dc9OTHVe1P3B3lEz1YI1QiIHBpu7B2oJ8wJdrE
/xIM5ivzNqXywWnz8rsrcNfgsOEicHS4F+m/X3C4t9aqS6yRiqpyb6OOtcGAz0Dx
0bTRM0lyACGN6ieE7bDEh2GO3yS/AJMo8uh3wnJtNzarIv13V6kPXwYnNpSlpojk
z/fh978ajSJG4NNL3Z1YEdp2WC7pe0KD9RP/6mIxMwhA6dZ34IPXCH7A0ydfi8TK
KZKHqrFvHKeMRwRJnWFIXOYez9f1AW4894bbJEfGuCUanyuc2J+/EdnGcNmba46u
UfxlV6oWeXSjdgON0xKxRQ==
`protect END_PROTECTED
