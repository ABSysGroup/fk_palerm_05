`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xT1fCNWgCYTwthBwYyHr+Gxr3aLa0V1XSqWCbnVRJbPqUGDJIJcr2m2qYARNk6kh
AhEWZOs/5GihA/URwDTHMOaDSfv35Gt8DKzKhu+2hB4qJTWhT3XTDYFywm4gWGdM
ZVEkMJpQ1gw5bQQyUYe9X2atS3azX22BbjqEexwvXibX7wFLyy4hIhFbupQHgggK
5HOCQQ7xLBwQaCKDEgvtvF3ziTXBLLBFfhMSAZS9vT4nC1EV/NClYSpIPVfgi8s4
z5fy01T+33PXHNhdO8yCV4YMhPPC+5TqpsurcK8pp5iWsR6zm4HJyVJ0oqc4pNhh
4vrnoNcs0Ktjod7FDHJ2XaydtIFdtppxeCU8XPUsyQAe6NQ7qCEzSVvV3pf4aYAS
uVyJsWOv2JTf5rOEVawvyad/XUwTp2Dz4LbGHZg9AXCxEmmYrcxVn/X0Wk8eFKxX
mG13Z06XQXcpQES9HKoxCmkWffO50L7B42c1mfX5NKj4qQ3equGtglHj6GPJmBcu
xcoL/ChM0KuNz15AzvGbWelUm54WHENh1BjwLdoXljVVlmE5+xAHMiFMk0xydF/A
N++ifeOzzCviNcxpqdGuVhaCUEWdTlJOlKEAvMvjQv1yJBrzuv1D8HCJC/jlboxy
ctv5rd7Zc82Ja40fp8lrHiLSenophmqce9yQzJst8TU=
`protect END_PROTECTED
