`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uYPX79ZjlWLS8goLRzeGK8Rl+Eqkc88JvYeT48MRPOiUU7yESsYTSBTGErhc90qE
1Kv1FMry25NbaCdfd7BXnUnqmkIuu73vemHoETganD6Uv7KNYre7g+mAS2qkBVqT
4wJdDryH0GD5wCGWn0ozEXUgdN19J1T+13i3gp/phOAeJ3e+mTchM4a3ZfOQMCFk
3invOA3L5Qz2UHTvrvNO6QdgJ7WWYf/ECpPd4CY7HvK8+X4MhjlkkJWzjhENROI7
JJX8S1H4wxmlzPulRHsFrYxaMZTaRfyI2OmZ+XIkgd97y+gdWfcV01vWgzC0Svu/
hBKYu/YgovJSc0vMSCTM4w==
`protect END_PROTECTED
