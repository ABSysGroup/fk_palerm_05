`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MbrBbc5PMOxCEewO8rlMnWAy98eMfqc+Ig2cQo5pAX71xsS9zRV3tBmM+C/JKa6H
xaM8Vz3CYBOlwPDX1szuOLkeQD+h3S2MxlZQvnGX9sgVmwM1tAd4u2MByXYnJENg
PyGNxAIepMNOiAx51eSO6l4OQH5hXnXZXEl6SUPg0UNKkYp91VHkkC1RE3UlbzE5
2IpGH1zvCV9oGLt0ovrFbjklTfX0ThFCTcJ2L/WcymasWgmy6RyKaxqRQj7oXHcL
61jfRKlp8+SJMIj3W9GXFZs7zqySOC2cvfESY4AxFje4KVFh+PNUYp6Jo1ZsbkUf
wrsLs+vXBjSzxy2f2eyManGTRVffZxKY9/Vjd6oVJb0laA2EQsh1cgMtJjrz1T0X
q80mag0FgshmjFB5bDn+bIzuIX2pvVs2Tiy4K/tmEfGeJn16pwUV/Manf9iMMsyH
Aqd7hVr5SEU2lGaQztSGzpMOheyIxbE7oH0Ma1+cxKth33RKunArQ7NuXOi5lz/m
qpLJ6Bu4uK/F2VNFelddZ9X00LdxncJ1rwhnKnTMDD9KmeWkK8sosR6acdIRlj4j
FJbkHTtrZks5OPAE9Kl6L7K4YCIxXZVyeHNPKiCyCEwW381SE4kxSHO8CUB32r0h
naokUhCOT7/1l5vCQ2fAphWYmZp+nr6tjiSOlGvKCZ4=
`protect END_PROTECTED
