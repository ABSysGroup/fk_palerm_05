`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EHNriPjYGJ+jldtCvFj3KZmV4NQiPykrNXLsfIFYcjU1MOQUJTU9o6JiWJ3MmQSW
YgoEwDMhk5AVhnhTnzC2mSfiYa3ORey06RYXMGREhXOmmx5Nh2rLXgpPJ+NMo3NN
d06qsmaRcEk2u9mnEozreU61WHGNALj9fZcEQGjFZfe0V2wK/S4p8qicmY7nA4Oc
aOkdHHagE1Q6RW0rz2W1jopu8Nr/rLsG+W9592ij5EuDMspBqxu9Xhdp3Qxak/gw
eHmdQNsWMmErvI+M7T1uK53k8aNCsT3BtBnzI7Irvfdhr40PSJJd2/o4FSszaMmc
9K37mBYq6gRyt0kn9f0bp/mgnNzE8iWxgcDM3vhiyjgVrEq67zwdfJE+MIE//rWx
g7lbinXvKKo9/eJgJ057ngtOEB1PX6cJFpaCjyKHOpC7LnM0K18b0yO856fH7VZA
r3TU8cL68AHUF53ZcH8FT6Jv7hiqq6f5epwxaVINuprFU9HpLxXaOfZVEiA5lDNe
FMjU10VF2E43AxAyFtea5jG+NArEJ5CDnup+bvXuSATxREsnLF4tKiTojxOufRf7
w7Z9KzLqqI1bac20PiCtY/YjB7vsHjhh7dLJg+uLi/i4ghrmchtaq0LIvCwZDVEn
bembo2jMZow9+SzPd28gzQJNHf2At8VHu6XtprEvKWULSPL2Ge/w6Z37oK5u8lz5
OEHdb580oZWFu+flo5eft5n7mBgJ+x2Eijz3wuTfKg3roO4omIKXBp5xb4/sy1cC
k4tuGGQEXCdd83Zp+ADNdf/KEPUc2eDhvKwzDNLqjSELGzjT3MSHMj5zwuLBAPRh
z1yTxDlj9kWOZR+7sPiXBbE2hGZCqyqi6qWPbgV8VNFu+sGgITHqw7O1BvQIHRWV
x62crojXnNu7NlNtwta3Clv58wJOj+sL5t36G7vLMhBzbHPosWheRlFoaf/OoLqS
`protect END_PROTECTED
