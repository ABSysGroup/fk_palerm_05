`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AaolS7N1JtIY/TukVPJoQXT30JfZPG8KBzcbPay65muMF8VNNVl98annIiQlKP9y
vfVE24Fi2AQVen76p4tOnmuPHP58UyXwOZky0ufIru8qaXOvPcmfduNYxGjLy7Ug
l9ebSN9E9LBug8kwm+WAPYGT7T6O3kLWyWphgIgp/xavPR/ApzSnqp90e9vOiqy2
ZMEkCTYJSBymB0ibY38vhti+raJ6KDSv4C8hmp9bniHN9YPzjAc/LRrW9XK/m7oy
/3jdASMdbWHkhCHZIQiTdNU+Pkyq3x/R/fZLJ07gRD3bX3jY+36E6v2Mhv6oJtqk
+wf/jihoMjQ1P61hdS/hC9eqbCoankSjjHBwTMlNzTY0PEMr/okWmaqP0rAm6JQe
PIL4w24C9ZS8xpm85OW4RJ9VTZLBuBeXqlgjIHoYzY/d7A1EBksO45ulMkUCkAbG
OST1PT3VYkhr+6eyXcT+TlwpjcYO4z9NWsRT/c7AMit6Gc4YKqVvnKiHlIRl+6BL
o4euoD+Hcu7JKDKosWfhJSNc9I2wBuPu8nH48HcL4H2BjS6VImqBtzgYAr4qcLvi
cmCZGWJ5+K7g5+g+xDJM1j8dV66LmkFeBhAzQBSndYTN4omKW34WIHRsbz4ySEjQ
b6CjMZjGfQsJNb9btOJCCxuOvjYSVYrFh6GW4dOJciXsnjb3SwBVH1w0sFmakQX5
vRogS7EG4oe//7Q1Fk4Hj0Q5teSLbcuNDaz+2BeQUT5dXZg3P8KCGltr613STigS
NQel+BCWUauCJRMQ4L6N+A==
`protect END_PROTECTED
