`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i+3TKnL0MMOWgm549MvhWTCuvJZTnXs/BGGtPeSRXdM4ekpPnVKBW48VjNKz0qo2
XhIjnvbw1PSGwIVobsYSfypu92iL/uc2l1Hn3TlUg0IedT5tbRkGPKd4Dkk1SKhq
5bLxH9gO4ieZ3MJr4F0sRpIcpl/s4nD955xURC+E/6QBPRqyRLSVntYTMtAK1018
CZt8L2/oW1TJ7rWpLbaEywt60pq9AVWOU+1U6/tVm1SGFZ7yDbh3/grcdMM07XmW
mc6gHTTksIjBJTwQORjcHnXn9cByzBfEjNI9+GJHm7lm9Llmpt1pDONhy56275V6
HukX/HWsQ1YHlYg1+n7sK+VDFNpOrYDV53NH8jvwxOMHKMNjVXKjkEs8UFHfXE3V
N2Gw/MVOLdTQaQKmcd3K0M0pOoJzTUX6fHJn9rCRPskMWQVk7J6BUUDG6LOjyhIh
RSQR8Evi8tvVAkZ1+1MMGTGgdep9niAuegE3rbxkkaQkXsWRGU4H46AFN14paLCi
kwgF2eQQS7T+ev1YhT9pt+UjwKsSzlIyzlqKypMyao2/PeTUc+4h4WGkC43Mi6c1
cbDoxcmDRB2ElpZ1zIOF5kUbDUunVx5aA7DVmzfH2istmGGlmzQz0Cc9OkOoCvWq
7QMzPGyhQ6J1/pJG+Zq990cB9fFKdrQdVlrMVFD8tzifVd9hyC3i1QMU1g6dMjQz
GrCzqkqAqYsatfbnksc8YWrZUhmE8VqRyTsyESkSyfw=
`protect END_PROTECTED
