`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5pS/sWJLjMvanneSgKFx+bbAm4s/MpKUEFki5hyjhwcIhnI/YaEVPfha91EEV0tM
9/sCbzR6ZfUYc+A+xCo2FTWTIM1itKaRr7DiIUER/n1puxW68IDAn7zUUUfmzLE8
edWHf4mlf8OZz+Dely6oqhRafORQJVKzH5E5et8KCZbJYxdgkDKNDPMa9MYfGOyl
uBUuPoXIE62NP2XPbNqD0CWErASOg6+0RpXLEr/aBp2psd8rOVO9OWTmdOgin51x
M7AGHy37ZN7QImqjrlpkpUY6NmwtFgTWH/Ut7J733dBQCIfBgk1Za06+FqcyZ8HD
xdxDbU6p5hQtecD001jYXKB+tE+Cc0wNKt7b0kHbHef0VCtJog6i+59Y4mwOzbhk
SRFYgUFv/ZdPfV2b61XIzwPQ1+X+iX2QgcVI50hdb5Ej7dJRoWCJn2HlESju5FiU
4Er4GeMubf5H93m0x11WJ3qBU5lyQWfyDhC6Q3b331o6lEZulcML7Zbtkn9M40uU
`protect END_PROTECTED
