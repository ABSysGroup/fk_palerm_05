`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AKnsgzrobwWI+r8+QbgYqlL8tc78oGiPJYmWTEpc74vG79hRqBMNabWHRu+GreCC
EUHZiC0IUGZ4bY5uNF4ELrOgjJ9/ORt+QWO/0a7Uzi+32Zg9eGhIHPyaLWzpbIFZ
sVwbdzFPZ77rm0OumhmO0nB5XMU9HngikhSU4h5ZRXq1UaRLGHLiUleWw2yzPL1V
Wkdp+CoZ2CEj5pKIphvs75XdNJrycgvVQHqzOCqNZky4TRfS68aTW0kgMIDd+4LL
dIiAHAuc+oQCIhYGdrLe9M2ZDri11Jl/v6QGXCNwhlF6eNYub5r+tH1D7roKrYYb
zCAXgAb8Q3YmMrcIpgyGR9ljq765p/DnehQuCQI4P5TqTQRFNT0F796GnZzvogsF
mDCm1yQXODrwVHv6n3v9wJ+VPOawbe+Odg02+nv+sdPolWtg7KOkQiOnRdIinBmI
`protect END_PROTECTED
