`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NPV3mvpOfD7L5bMCt5kRodvrJ7t4LVk5QwIeLvoZV8XF5GQv5oahz76KzpzK125j
fBusB6o8szxoeI3ujIcVFmVSQs96Ae0psLD58y4Yh2JLALOBplDd6DLOEe46IOlJ
ny8aQvTF5Nh5KBLBQ/TdWW+EMxppLV/GDJmH2CCxvB2LNeI2Se/+ICZDu1IzuCQT
FauPzvcWCTg+Upi2oSQuuZdQmnn02I9NbcNT8vkY+guL8yfOewfhaD3sdGgunO65
KkO5AyYgAgubOAPYakdKOCNtFnenA9itnfgt6i+Oj5/Fy9q74v9QOXtN/QcFPkLs
oKWhUC77xmE7E1cp9m1PFqfWIS7HPl+PUdAISyV9cpB7XqjNuCZ21ztMBjuEmsFe
7ZeCfzQMlTBfUCV0UcJeKja/2NJaOUAAqP7PhvbnGzgrmNeRnIN2k/HAyVDQn3QS
l8Uiomg9e4VUWT+wQYUn4w==
`protect END_PROTECTED
