`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SkurI7O7b9YIpwKzwvBwV29loNaqLsbq9kv6eypoQhhgY1Tb6zF4rY6xU1D4Y1Ni
h80jIuBEk1qHjDf0Cr47mEYALexBo4M509iKErUHHnVfJf0b1baUuBAZ4Ng6cnzL
MViiXDzqtwAq/p9o1DBZA6LBu8rrM3PrTbYh1HASdW701N1j2uZ2jDz17FJrSsDn
zX9tl3t67NMiM9wQowQBAUopM9TXkYC59rvzZSwWR86aAUwkKAgK1aD26chZ0dKx
2uFysKSDexCqcgQdqwIXm5rzP7Ywder42iSP3ECeGEHKIPP5eseF+HQVg7jvmUsc
uucOr+VlQ2maU/J7RrKjZ0JCTG0zHOAq4D1/cse2uqG+Q93La/oagUZfKFcRE2ES
rN1vgjm1tsAjmZXFViL1OLmH0VQG2NCOGZm8O5+c2pVzgamySfq3nAZCcjKThuFm
Hz9vJL2nwy/ZMMhc1ijq1pJrU4XWC16M05na3NQDbjLqdcUDACn+vsYebyLBhEhB
RrMJqy4CfDniFEXDK+uQIV5wzMSrwcOYPoSYBKszpdAUu569dxEfYPALHzqXVQp/
0yLekqERje5XW3FkLFJ5Vj45+bE29iTm+vEAgqZAcyOLzE/EcxZ1R35Bc+E4nQGE
CN1MDaGCv8cwEEFWbMbHctBeZCHodaxEwwQ7Z+hDKoYn3JHBnEYIccH38nShkugp
t4YY6mz2WFv+S7uCbfFc1mrAspx6ECSGqELz4HuQRSzaIaZ0Qf3sKf989NMYaPFU
gKK0cWRVQLCwNPEUfZy/RHUI0p8WdSmRO1qw+GyM1pL9F4iDOGQWtRfOM8GPKgBt
Ac6Fh3mfFb50efLrCHeXuAcR/prVKLEtH/d3U1qmjYMatHEdNSik3bMmYVsOIzhD
W0ks2pWJ7W2fh+1SzrSm1Xyoak6sXV+EPRXazzTx7SlYj2bklFsZwbIEGk5lAKu5
+6mXpGt+c5Aj1KjMo7Dr7Ro52yoRn1jsAMr+SO4wlP1RBmprYGq2nz76+UwVrbdx
5hSFOl9TfBGrdFXlERxGfS8XxBc4MxiA+tiRRJxKT1Uxhor+8pMt9LUFweb8nNx9
hrpGEalS0kG9/L6jBZk0zOsl6u76o7hxAQADHZNHRAxAmHpDBvZkfr4T0zptTzUk
fr1ti3H/eTC7iUxKPnMg+2Meq7Spt0qg8gneq9XZvYOiPh3aHkj5ihSjWJjsj5qR
qVJrWhr8eliBqt5neNQ1u1gmDAXmRDdEujhzT7x4+Ub8ymzVLN2bYC3aUaM/cV2n
mNdedehtz2gaURlriefAPv6dF1Jw31l94/orVrMGjV0d5g4dyFxnni3w8hk1nZEU
fBfsJWbzo+DEQPSobyAjSwnC8+ZjTdfDwlB41xhQ6YhrQwBhVt7VVh53GL/2HE9Q
6qYSEP27kNvWx44e+8mJAHUiYDeUZzkysEIEXk2WFCRxY+67Pykns6xQhW2fHxcb
AMHXj8ZNdAF0zKnhHKard2OVdQsU8URnQXGFWd9AEizuHeAs2s2CK6lB5cc8H7gC
qG2Py096uv7UAeEi9XoHihVDkpGz5AcCVeoJEhN0FUkUA1F89wtQJxGspmB4F35r
5ajDFe+kruSCM+pHNYihalrKPLv47qT3NnxBjq/a9sYpe+gqlPIpq++7XCVut0ep
+CUOcgelG56MIicQ7IUwz5eWALofywYwuU3Y1dX/bpKq+Rh8a0EsE6jLc1qZJEo3
nEskvMUrMBdiL7qASMjXUBIhKN8xmA+xU5pWJ6jYZGIgJwONOCNk7WXh8q5v4P0G
ex+AR69ZTSqKuLv2t8Hc+GbFE9Q/imBpf+NwlsV5CdbuJgE1pyv61Jeg/RKNjuTc
LyawXk1locKVj3bcK6rWFGfuMwOKfHOM7u8HNHN7TrIM2NR5qv6Aw/DnkmkHy7+s
fBy69VPj8QvQOpQkSB5ROUZXCJHTmzXEPu3HjLPzUZ8hXdLtBeMxf1XZswLSSwUc
dyHhQys88mzsEOw+WDodGBWa8shGIT4gmo/F9WoWYgQ221U8mPGrSxalSSq7ln6p
l78GUV9LM58YeIUCBcHBqKvsOH9M/Uc3/nno/EIb9pH7MPeu/dMkoQhFO2XTjjp/
3f71XXgql27JcUS6eUPs56tAIn0oPipWClTxBo163Sstyp110KPeBcCPe2a0dA+n
z5vZp6o/qWqnTcy/H1gedAxyE01+YCRgJFQV0R4MNVQZhAVD0wpamE4QCYubBojS
u7EPfLdDebXu8eO6RNlW7K2dXf4cViVz1EjoEf7Qgnxp46AkNQZIgbgJTtsLtLbV
qVQBlFen2topJ0HwDjFUHHDJembI7/YUV0qff+rzSY0Un8jqAw5fS5+61EQ7hGyU
qke7upW/onKB/Y8O0BFmvkzEc6r5RxZSeH05T2GAAj2khN/KtFcfm++2SUtqgWBx
wSt9pMwpZypYRx0emdk5NRtruB8AMVnBAlxyRVrw33kAq1TOYxxsZK8zmvBGbK3O
WapJL3PohMwCUIBf6G/KK8y7UIxxclfvIi7t3XsulJz9EZVmv5KzNmu1ppIioV3Z
yNOxSpiq+CqGQQ988JtDGE2DD/WWVUxyXz7r2u4E0jnhSPDURkkvgo2m2rfnlo9h
4JiJGJbXvP/llFBnSSIbA4TfYJrJ6SqyGYqtq+k638fOCIR9Yc6NDBNpC/2TdV4F
mCSrEPkryoGubsxUQlfjpgZ+V9OrWUYqvOdylV7TB3oMXME6yYlxte3dtodS1LQT
17hSR9mprEYnB2SWx9TkOJByomw9PEB41ModP7YJZQhQY28fumEjbVSseUqW+Eam
lcycowH9uTEscDe935//sZ3FqI2jk5Rgm17pq374eLBl5f6qdz+jxY0G/qHHeAAA
HWUH6UEyhgbk3ysApisu/UNhXmbqsltEcoh3xbmQMLbPTUZjkQKfewvYIqK7IH2h
fYUGQnNW9i65eowUlDQV22mPRmSjNXohtL4rXBgubyXuC4t2w+DYIho8Z8Npz0tt
tm97mpRh+LT3349czXIlajEYAAof+WJLKtBAFgI1/Y7IUIX9JBM9rJzbWABEdn8U
jfVyw6TEWcBamIrLWLGdJa23XsrjrniaFR/OWSAYAReSeyBfR8kyCLaMn96Lqu7A
Z1T3C/u9c1uKrJO8SxCnlSSFgfmXjEFaQdO+4BLRdQbkJ4vcGZL8Y0ZJo//6JAOm
k0mfoclS3h4SZ0ORbISQj1g2CZ7DXNeGENznTzEQWGEqmcG0XLjiyNWpND8XTmhq
UvqTC3qgRStFMg2li5lPI+4ITM5In7/Gn9tw7NAHcQJktplMi7IzTg4eAY8JlNZJ
AmloNnMKKaXzZDE3y/OMyM5RTAGo+V/VfYhvb/LXwLdfbxXB1yqjYYxHTMkP7xUJ
Xq9qRWeItxCJmmYoiCVe9phOJ2RiZDXSGhU1Ysq0um6ROdjgjquTrWiecYU5Psb8
Gxqxu5zBYmPjWEl79+iywCHunWes3zZJ4jOBGAY23kxgcSNnhZfmlrZiJAnRPQwb
rLfDU/c7XOVyLiDgyO1G3pyexTsjPXgW19OOgzu+423BG8nJ0k3qfvAVYwfSmDCx
AHya7XcUWCMHOZHeKLqNyfQnm7L2py8QJuZAG9k8zKqwsv1IoUBKbHq4YWrTIulF
yKKJt6bc0mz5w+4okTAmA//y07MC6clAz1CTMp/dJUYECjQcUydWsNH1/Hwh8vxV
JnL4g1ytbAkvi8DZGewxnvT3Xyu8UNhRmbpOej8CQjNgFvTNCZlcUSl3C8tIM6/t
7iI5Euy2CbtmgIbyCz6wlc2luJmZP4sDcNLmzc0FSh//XtOweyatpywwQVktL0Jb
GJkxkH20sH9Xk3zlE919Lh6DeYXdCiBZyCoWeGsf4MtTF5paWk0x8t9X/AAoZA4p
OOxM/7hnnrZmrkAaa7HE4xg88K3WZWNZXFkEaAaP6QQiIg6psCFALDjuXz6G/6z7
Q/zo4LiZSoyllxdXptjdGhHVjrw6rRE0NMJKZuyz5OJS5MBgdW6OpiIOhC5fs/la
R6drlnw/9NOcOWLPBsQvAXwDsOApmW9uSZLuJSnZx6KPrVQJ3HzHREBuhS0vLHVf
1u8ifi7iNO1NUXvOcZl13E02xEnOCOh9GfZHLZ1jJcHEjMhWZzzgCthsJdgNEoFD
9YGFpE3tkfwzK8AJS6vNP7VE0qQGtBROFz/JWlt8Cqrw96lQfWn2VJpPTnIrwTjo
snsRaDrguKlhUEYtCVcQwpSmZT8QCWgvTXhViZAOfRZc9YdUX113RRM1PJHgBcU9
Mz5xVkHwgw+fcEk/7Fgb5Nk0GbWCglGXcKHfhCsYdXo7IJ1boGBu1zW5zObxnaG6
h738OO1I2b2W8EvOIWERYvMRPH5PapftwYBlnIXOh7xtDIv1MkNS2ZC0ga9nm82U
uh1Owo5ByMX5i455le0iMVoQO1Vx+xNkLHdAMNw9cVAOP3JQXaBDuBrcDmI1++jk
0QfKTcAfZm+2jSbcoqmLhSVr1itg8JwGbQc/8WKatL6UrKb2z8ZOONE4GV4LroSa
p0u8NzXeXno0WUNvo6VHig7Gaa8GSyX5deir/nF6geyaRqeJ+sfR7OgR1y+FKjE7
Zz48umQmDV9RuXe19nw0R2LtA5phCzpFN9lajNQm57axzy77Hnux0QkE74508XVt
3xdaEjDZQN1qWowd4uxrqr9nxo4o/fNijDpPBF0z7e1Rng12G85nLAoYONxpq7JB
bvq7o2vj2WhUREpeRM5SW63982+FoJslSVejPspjLKLeeSm/9PmPm5wFLRZB5HM8
FV9nk6JpkaX5MA3v3HhquDtCq8PtcLATDeZQT4EqkTHbkReVcjNstJefy1ZAlVI9
5GoV64fRE5ANj4/JwfPLWRJb4AK4uPZzyKF9AEaE6J96VMvmgpz2h4iLP5zluaCx
zqYpwr499/0QSKHkGvMgi8om8oiu9g9JBA2H1B+5xfkXDLo7E+8kbSEob7wytwiF
DqZyRxaNMh1tD4d5akJOWNjeDbzUamCRiLKQxm9yE+gR+ptn31CClGnLb47XSR5u
pehnHnwNZEuw8B+3vcy25XxycQ7GGvZvcLFHgNjQxnJ/D4EyN2X+kny0keriO/+w
6H3SOFdwIplJVZfSPwvz4fNWgLnjs76r9SHXT7CVCJUJtBL/u4ZkuifMzaQpT0eY
2AjJs0BjObZ+f99SPDO32GonUeaIKa/HajgSjNKrKlD5TsPZcwnd/DvpGO3ov0iX
rWnWwv/64eK6kWgXHVVo2qHFx+SOTsNQIJsxVQzrSYCtYapv7a9/uyeZ9EXo0LlL
zBsAdkVHar6rjgajfAkSOm1UFZpO1HipRfw367WulzeG5VuowefUw2+N6D0Bcnsc
tWqbck6HoactndOTeGJrCE8c2pqgAS3hv+nrmFSanBzmJYQxHXazM2jaWnwlPPsy
6Q1NrYK9SxeF7+YDafWmHPfeCKZ3wvQOOojcdYokZOvdtVvQ28+9CnUq5ZDXdJYx
32ArnB1H8e06fiyDSD2nLtwOwOp7exMKyq15trDJaG+VVykSuIrwv/AsInGy37OK
Ho3T8F/TmgP3FnApLmSfebRXUc2CjJrbawh8zqiFLOI71FHRl0Zq33ZkNoEEyipZ
9JL1isFZ7QxVWG2ltIA34ZfoixEDhomPFidvEAz9SY6ubNjoQBBIOdczCD95O4cZ
LZoqc6G6lHZWMboMPSl8opa7WSzyD0GfbSLqIXfOdyWfQAxsqiG2C+Pa4u+ou2Kg
fCQ2HTF6kpeL9XGH4Eonv01Pk1J1uGsEul0Dbq7AxWOESseOjqnmw0YdW/hz+v3v
fu57OtlkVA6ZCAW91YKGdksn5H5mifosAksikM1nI1frKYdi8bbr55TGHK+yNVQT
627hlNsTBc3eLRlDXJ8tIJF1Jmw7puGXbQb00rcBy57hR0sEl0snJeDqdxtd1478
FJN8TsG9cmGyCGc72Hj+s8R257l8uNgl8kyavsPpsMu6BAQbhdgsiU17Gqt6roZm
Q40DqkmubmRLBSw6EPPOVdDEt6/oObyObBTMuhjj4aD3q3rnEfUxEKAZeKpi6kHA
U4VI6+Vg6fEm03oufDvlGg3ZtWWF4OXlIRzmRb5BqPEDvAPQLIFe8gYwKlU7fv5j
Qc5eIlyBwVJGo9EoUQSYcjHQZ+7znGlJfY2stnMLN1dUS489KAdloe/a936Yb+OI
P+UJQt9ceTBatWScK92dTfnjvVGAkN073B2YWn/o/a3NNp2pGj72eElpXh7YKr69
ixt1OrSnblxt1qSphAC3zMeXQZPhf1SajFqyC3WWQt72V/Y4JjcCD444AVIEdSpX
CX44slyMiCPrJHtdEED8Icgsha+tmmOW6mxlY6e7w7pPy7FCu7fBGrIJKDxucZqa
TmlTUFoqeCuLVm+Cbsj3dewWk4chSfEBdMuUZ13Qodca5dSggvXu+f3o48z3SCWC
ituFaKVw8RMpXiHx/zRPXvE6bhmXwub8//YL19VONfrbc0w2oCajbYWH9v2a9PI3
68OUaS0trcZNM2fnKijkofg9lxqbQoblu8wS3G8s9C1fTaVm/ecq2yKv+9sbIpqU
ibxfpRrmLdwmiWqqgQFC+wjbv99tJAgcPigyqd1TU+k8ZUFAbEmsEtlQaRqddR3q
eCEIRcyDk1SDwwibCQzRhuMUR+XuF9RnZmKYBW/l2E4W2N145VFr3Vz6ccSpemgd
xQTHqAswcLx7AgPNIyLcJHxqo+y800QjfSad5ilhRKhb5H9HHlve806b3uSvWETE
f2tduiDDgYkuDQ1EUOk+QWNNTvqd8+V24cQQR8AA5narAYNkS/cPlp3HUXi9e+iZ
jE1vaeTwbVJjGsF0cpRhxzhN/tT1GpPGT1RQchsfW8ROCW97gy9JrbtnU40WS3w+
`protect END_PROTECTED
