`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Os1Ec+cgwSQ8v8AarZZdXhBrFMa9usHD92Y3ZhgnRD3vVGfLEwfaJi4SES4UxHaI
6xpzWMJzqYVSEYwlA4cogZ1qCgvTBA6Uzxr9qV6fKOm3gHqiTpS0Z1+7U0/ShhKc
wzdv+GKlLnZo6G9fnj9YaHhqHSRoCfOa7Jkydp8wkRYRgikoJL/9TJOEVyyxCXnR
HUryo590uWh2dK3pd5egUPX8Zxv4dhZjUlVypMneDLWKJ/xKQaYuwpqxKJT8CwTy
rSsol2gZ5Qwsc5adokWM161xueLRnZ2c/PUQbDUvjp8IXXaZgLnw8Ms1fVKqs26N
brauNo8KbpuWFkodZYf8r+HcS9o5WWxPx6a7eclNc4clbA2TxqkNntMDBt4nBYQM
w+io9m6s6n32z4zrbFWUgogYqjb7+a2LUPV03KjWeo22Z2qi96/A/Ipmmr+lOH3Y
/YJHpb+g7SDsg3ia/dxkYEehORDqCoXNRU0mJ0x3ROSzZBHKejWvZz/VOPA7bYJw
gQ7kmFhT1J6+vs3jdQ1swCG2/LKgeywsSuy6H9CVwev05G6xS7N2kA1Azp3zyHUz
diKXjRLXlDvKLIhGRnuh6tH6E6kMdSw3QCu8UX5oZGCbTQEupqxJD0lSzV6Sywss
4eP1q8x2m+Bg7C6s6XLY6y2tEpzbFQL+9AqVXdiB7gQAp3gXsTVgMiT4NuZ8BBLZ
`protect END_PROTECTED
