`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AlsI1ug/hwE+Qt3weUtP+Mv+BnVm3DKZfhPO/+MBFgq7GSWqdipwySn8G6GQMhlG
6JaUHtRw7EzVL8vBOV/lrMiQl04npMfuLIuWxkAxG61+0hv7f3EXt2LF1LiIbeRx
FqL1yZOWqkUfojPHr0Jjznrb404A1fL63tOcPirQezsHRbKEDY5q/rDemMp8FzhJ
Tbqc7RkMG+4fIF53R9azXU/BTeyRUmMPhQ1EVdm/agRdofXh8HnDtnB8G/UsZQEe
Tlle0gy31LYD4x6TH3oLcQf+tVTAOxwGrBqa+fTGrHYFDMh4Xx9QQCZTFPrwaKbb
/LZjdlj0vVpr15DTBaBKwHYJawjv3Gouvee6o3/KNSZuOrms3kzwVvjKDLq0QQqe
V+szj42HNj+PeuxUvaHLuOB1OKX2jy9lXSvSta664ILITW4FJMDnj6suBPR9LHuY
ZzNFzZuyEom4fL1vvTIFzx6eBOo7GF7jBgKneLRCqEmru4WOZm+F84FUxvJVSVab
4O5azamL7nXh9Wl6wjPFLc2T2DuxA+X1mjmGxHRSCdVMPcAmYTazYXmPmPFw19cN
a/3fe4O3LNLn4wmchTASv0Ykei8QlAogYibQergMUbRQjObiHnJBB3TWVmnxnHCr
xbx7DQqQOE6gdGJrTx5KmP9bGSkeYaPVDQ0H5AE+L75Qz9ks8zNcfIMWzpt30kX9
gBtJHdPHecJpd6YIiTInDYA/KWRBLhuot0eq+QMY/3RhZqYkTFshGkVhy5SmMx7d
u3L8QxJlT6l+DcfeNKFJfIpMQWFVgnkzSTLOgfN1V5akz/VkfgWUqACuEHFxZWU9
vNEI2Y9vM1/HZK0JlEkfKj7RALGALYRLk5xcdVTdTvo7ydE3Lmui1JpDOBvaP7EE
W5xfrw80iekW9P1gqQVd63k9/qXkAP3Wb/+rjW0DqlmO6lD9myFR/A9ywG2URmwi
EeGBmCa/qt7NF+Y94p6+K49MYXuabg5VmeVcT/U73kakXaswE8etxvA8adpYDcGK
S5AWMHFeKaS4SDKjrkbdfpj+ua0D9hN3hJtNknj+8z6NRRIU8Wpguv4SNVBjHPC8
Q4NHiu+r8iD7AMevoUq6Z8BBEfVmooSTSu2q/XGzEynEHJOl5DEjYLJblvHULbAu
yMKGo0yHyDwgSmJ0Q78b0NhA/UN6NMRQNVLZzra70RLYK6pbE3G87T5AgqC9iE9u
U1B77O5/7C+Cez0JmK3zQz1B2KkU+9vcbeq1UZ9HdbzNvgmUULGsplK0AJCNOBu7
9hKFFbtsUv7OI3YX//qe8AY3O8MGn1R2U1Lm7quVX7KoYynXCg5jxHD0PxlSArez
PGr3kwN1PID1XIOAo4EeTHP59NL4UpV6Y+nwuW6i5DSYRCBB/TXRzbEfgEMaKINA
aui6IdtNTV7WgnsSvZjbTHYTWRL8NzUDzIXI3HorK5t6XHcIey1M1d8FH8JSgcOE
gFFirZyv5VCdPcohxZ4vkpy78+9aXA4MQt3cslOHdz2pGU9RPBqXHxgV9Jq3t5q0
+pZOho7C96/CJz3Tn2HEOh+LMvJfqDtB+N64cKgXw9st4q832u+37jjsvTW/zi0G
f9CiEa1L360ALOipd3MdE0dqlg1JZzT4hj623BDo0DSms8uOZJxMhk9jd+LpqSzi
Xh/9sDpZklR/4K2VSjT1drj8JUwj68OZqzwsXTlVT1c2hraJ50ngevZNG0z/QQOJ
WU///ZnlyZMAcUI4Iemzwy52zZpMdY61fC1j5xqUtRj5C4ORwjXMRXQN8E5JL5mN
USD7hyKNLF4hX+TR/7ZL6idXIie/AxBxJ+1XK008uUAvsoRV5tAAq91vg21LdZTT
0tztHkm08BAVFEc3CpbRd0mQRrPKhlvv4kj6mjjrAM7qif4hvwBygRQTxLUdkyB0
VonHIX23IpgE7JzLtgHlH1Eb3Z7QB0e2lUVN56+4FYX4M4lAwEGTLtbsFzdU6w67
Brma4ogij6fT4ZHQ9pqLwPR/0pMIzDXzH6aUCrWNJn9xdDC2qiOL5qxEHGMLiWGR
x8FdBAbElJKyaOVnwdxCUriyUwCfxtH4creXiQAD72hNb6THfL75s5RLNnFwm6BZ
IB6bcS9LqLaeTEoxPISuwWOCIG/8Aflb/Ku4vd2IGNetBdYLwmcSw9TyBkyI41eo
/rL8lggbVuzDqEvmlHfbi+YGwmt3r11DmpSlFEe9xmy2Io1GBJeomYaXMfWO8nkh
VDZoF5v+OtcYtHEao2nSA1K7R+J5AH8iIMT2GPpwnC72v/eKyUg2XX/UJgQDqEry
x4UtWbJfN+tqPreYcS02V7y92nfHF3BnYZErrrBUAl1MA7oPYkrfaMQNDtdvQ321
GWhCc95/OEDS+kCotBa79VSNt/+79+4w8NQfdevrAbf89OKEKmoRQ4vlfRnFYA9d
NDN9OnKhQjLrAm1lRho1YhjO3k+J0DzYxF6QdzlsWhCweN3NwWYk5h/PcH12NS5N
Tb117l/w2G2uoRzl5B4+0uuNupYhgiuFWVZf59ew9JHuI5ObBGhu1Bh5Rc+jNvaz
Fjt31WD5wGpCAmjTyYuXBgj+bE8pCjPGNLXbFBFNDsKymyEzCSJFBuSBPUwvbFoY
sLJgQBy5u6aLCe4Kzkk4jP2kLrQlK5br0sLojjPmmNTxlr8OhDxxUMuRq3om9GH5
GLdTUTjxnx0q8GOdd625upIJT2FhzQaiZF1GYnnMMZ6+jBiI3VdADhS0y+upBD3z
wFr7txsaEKyZLRrAwBhHMG3IHm0faKwGSIR5hEcBeNHYt2Pqt9tWMp6jZAIRy0aG
N98I07kzY6YDqmCbw28cjd3a4deDHI45x7aGqt5N0BVyWbghubYycb7GNHvMZmnd
frNtv7etKzFitc+M/1hXJFKD3xJxa1p8+hMkW61OlbaNCIBYEMaopOJuFoHG5J/P
xjEDcDqnviYFnjaZFlq/OCNsnCICRlnHeylzKu80DnApaT79lJNCfbzM+aGtr8RQ
qC9MzZAoPIAJCnwyXj1WqILJ+SsQqGMy8isOr4/hARwM1Zcb9h99bXmmNDPB8N9z
yZnECeFJpfg0rBS1JYoe4k6pLlqOb0sCfCnad8sw1gf23H9mYhyXPa5X6gY/jjsA
pVDqw5PprMF9K06C79gaB/xR7zhwO167OqDE7p7Qa9YVi7fvU0Pt/oiqRPVt18dp
Z4dLHrtf552KS03mwh0xlkpa1l+H4uJMEjuScAaIwGv/A/J/3AkVfpPIpOMAK3t4
ZIbc4guEJ60vvCRZ2nE45uMusUiUGZHgwQ+DKRJMIwCL7T7DCwIN4Z4Tzzanx+oC
Te14zIsFzOvqlAcUXGt0wn+o7kFIzwSYCaSJM+azNuOppwYIx83XaL+2mknefpaH
ileXlqRl5JUspLJw/G+rXy0T1o1NmBIz9xvPoDGXnl4EsRsWnlGEd356aF5pdhG1
reQSMuvf8Pi3lQ0DI3aZtLh+ba436wwFibPGtWMXybbaKT3kgtkgG9QuSCt9JyP3
U6iFYttbB2aM7oRkNeCjWKWWilbTW3TRoyPAWBR9ePj1B6CFyIQO09JxR16qizdE
rLR4M9vh9p3LFN1XnMSdAfwhUJ4Hic1hEol6IfnCfYPb2hRexk6128kq1mNEBDvP
Yd36KUtkVTlQ4/CapM9R0X2PuU2WxkPx8YwLR/4WEzDcRVcjMLociHYPoYwq9qGv
bF/1Z+tlaWsid0jp/EI23/9QtaRIIhq/saRx/H9yMRP3idKee8be1iEJtCpnlpcq
Z+X51uWDXuL1JFSQX1dNCazOdiLfGXbDvPTZDLZy8rfmwLIScdyjbolkdh4cL8LV
Uwvrzf6YUEQhJ4NpKxY8Nr/2O8/D2tDMoj6PI1j0hk96YoJvaCHjN4EGAEM71NgY
lFl1wrdvPL2OlOtyYU4rRPzohAvf7sFvqSclvRn6xm4miPZKduH+9g+prrZeJzLa
GU5VKpRakC5smLpW/Klww2vnbyynzb1VgZHePK0IBHtmi9nX7iTIiSDErD4KmQj0
BLZJBYYs2F2IN1D64X0+SAp8yhO2cnoN1ZVM0/JyV5G5BAqNit0zc7fypJNEw97l
1Y57LRD18sSHawTzeBzJNwjNLa414dSRLtroDfMFTgeEFLS0c9kDOb3aHm8PSM8r
buw6N6+pWZW5uJtdidh3NcGwWkClKSBPLIwRP/9myt8S2WYf1RK4YPmB1YSIAe+W
/BqN5VXBXSEWLAj57NjXExJprATzMb5rOPrQ2vXvXq7rkuBLlXCF9lZ+TwtRyWKV
xIPw0sbWksvgFbowRhnWuigFSdOU4gLEZtVmvHaKXULX580ooWF1jARSfFBz4AfH
KCjx4JTCmlABU8P3fSXGGv5MwXsp3PjKFYaeBBSM7WmmoJMK/ITN1EhYqfDVIBx4
jO+iTTcN9PF4ofI0iyFJQfa5pLPQoKNPAZ+rf9xT0MEcBOTD3rmnaDNUinUpgGeF
WpcnZayF1aawUBZbBidnYAq0f/zFRuK2excyOurqre3Jqxe+Ol+zAmMkBNi+3v/H
YEZfFMWETcTwQZQjDUSFA9Oeah93JLePjapABL4CvJBduVgVw1+4RaUMy+N+Fjcg
SBRHAHfCQdaN4TNrTm6dDUdzhu7+/L38Ai1aJxIf2TMEjgJuNk+4dfQQF0iO+k0U
tE5oADZfxsEo5eiDVnHkxneXiPtRT1aSyb+IujjyCJyTdl9kyKc39DfZ2LX2Qil8
jIXtngInABOPochLHlAENO1oCjCwWXbLQ1POMMZsNGmi1wi/bN9D1DBxRLtbfx6f
fWO9IDYBjsLMuLHp4/FMFJ56yCJkpJgmql4lCcYarDP3CDa/gKmYLxhURisnq2gB
Pdss99A0iN8euhttC1nAWE+M/63isDJpKZaqh7kcewZ0Qi0SKlES5lN5QQ8dWN1O
RMobVH/EUknkZr1S7DQ0mAmaDp75TCZLCYV8B/xzY2QKdSmAXT3i0MI6v5dzCFrt
HUlTT7Tu2K7J+oK1LiFSf+vEeBYbDWLfe+qEUqUbIcREflEWaSitfRPBxWFzU0fF
hv8OfFQK4BCHYuk/lIw/CdJVefugWtBCoRz11VexeXuXSDpqD2/sC0dGUphdMFD6
bH4hEkBpsKnHh2syCkg8Oec/EKntKy09sqU9BmUUft7S40cxUvwk7ozXo4oAw8sd
rfoFTg9ki41R4ksAe8EhQR/qg69q36LGs3U/UZLpmw7Eaw8rIqPFipari3BQ9v5Q
3CvAvUN7/8hwYE3uM+g+9UNaOicMS0Zw1gsv/IlNmiE=
`protect END_PROTECTED
