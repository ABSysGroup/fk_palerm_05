`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rnl0A0cBzf0yr86TOXRiN/P745SwXF8HBwQSSTMP5VD8mCYYRSHYzAX3txWN6+ps
F7PZq3xCs6bgn32vgKiiCi3F9dkKpDiZrkSeHvZjdfmRyjjH9bcA3MY0o2oneIJM
DxaeyeiMhdx8fAHJyvP5nLoohldGDBzTddHfWM083CcFce9c0kcAdq29CpkpsfbM
7gJUI9BQUM134JgBZsHvl6pZsB/XWE9cMn2GCqYskzjkG4xZAsv1Xt8l2HAMsLDj
dx1OJxCjATcGmL3p33+zCliZqklppY9VLwlA6wkyUEnmzAQK/1zSV1sVDcfEE/88
Lm4JP0nRbJqZwzPYyvAiYEh6CZGLqJNopboc5beMo1YijUQhBre2edFSDQSh0lTR
Q7t54ZT64E2SZY+8zhy0nN4iM5gxy1DLYglfxMXVb/8jip2RrEx0VsExMeVUP7NF
EKbvxH0+lQGLSdwB3OqzgBLkbToQE1sqW4xHJUQ1XHE2tn2uHLKOZ6v+EO4hzmwl
PxOiuXfTN5lM8zX23rsP97M9Bpmjm90DE0zsd89AMqXDyY/LqNzEMnXB5+Jgak/P
U7fdBXKuBTDVqwSBAUYnz5C0mDvat65xJjMdghDJ7Aqy2hKq7B5sN4UclSlhoHtl
QOFj3549Chd4rEnqUwM3TvPSjLgw/Iyr+ierFD21ngIpmRGOKH89b8vz6Cka3plQ
ZeSamZ8yt597oGA3hEUFY0YoT9r4S1QFLGS8kT6gZ6TXdJZXIj05bePGETy7T2en
ECknlj2t7fft8TsW1zEg82jJU4bImTOL9PDiu/x8vh+71PpT5ysN44AhWsmtiv7K
LusZRN+oC6ed22leYq13Lif5lK260px34aqWjhNmGGTeLXjih0hM4PXd5tdb/rPS
mWOw+akU5ZCMcSTOZhmMbmQPDbTxcG50lGm0u6tZ6UvuXy5LQJwyotmmsBXwUYW8
0jbTc8p/to5rOzYQ3jhzrKT5asTG09VGtF+hPW1kuASa3IvTu3oiAe5i4GCFxL7I
jg0pwFeZA2KR+yGAUhXYF+a0hhIgdP+B8OsKI2V/ItA1e7AbdgoRUw4yILZ5gMY8
Gj6B3a3SFcudnTnjXsnSY8QxPEgVcwKZzJxQ/VtcELWLvCX0b5V8rAj3bDee0tST
cO5zP4nvgyY/OvaHKu+eFi3gdWXwIQvnWsorlghizAynfjCQheDXUQ5Uv97Ig0L3
QwGKmussuPtP9dcY5efqoIHzX3mqfvZySV2iB9ntvHEHD5fffH8NtwjJ0PW/8KhG
Glg7QDMJOoR3FpYN67L0uym14OsJFMzBqxNTh6/iJCOrXfPFia9w7V+nfP5RYM7/
6KV+arhUJ3WGqx59r9m/vHdL/zJ8fEpAVAnou2JBirXju4516+MyaoInpBqqE5dl
Cc3FV9ia1yD5GQAo63H8Llyo55J8QHvi+pkpNOVPWaniqztUc1Jbp7lsZiioEyBn
un9y55inmk0SEVH5MiUZpgmWmkcpBoKqjGMLMEEn3q+WmB/A0mWUEvQcqHUJxVXI
mJTTBrwVKs2h+VwXH0uET+EhR3oLQSjLj4+phctp6qmmzwa4+Z97eURwdAs6FOrL
Tul/MpdRR6Rd4CscqPLaWf0Ce9U4eMsYqdIVSPW3aaH+R4xH4dMulpk3ZKsdy5KD
ZmgWv6SkU+JKTR7S5DO/ruLyO7T210cxbzamCrAZ6hxPhyA+bi2GkViVZroTjcvm
O3Fd2c03j4HdFwhyo7TWLbCvHEHN+mGPL75o3NFfH9Szf213A3fJYxMhkZ04dSJP
i5oSMvQhAAiqO3YEr2c73mcszOAVc2OWiTec5lcewHfY4CsanQraE+9vrd+Y7GaT
kTYXF2smzeQdyc/tCJ8Ru+fYX6DslFgFP1uOtw6RMCHthe7SW3+SnnAdmk2dnL5j
qwNC5xqBJkNCyiU/iIQfPFJFexoyAD1xQtgnrnJFGWo20RRP+JPfOw01B+pWB2Gi
WwPXffmF0+AO56OOZBsOrJs7JN1iJDHV2N/wu1cRzmBFoQ7d/pNPnrIqmELryqAz
8xQ0Sl8VzoO5hFiv/dotfwx8mZP944qe+wkKF/QLZ7RHZYkR33gdCKKa881WSmpx
UmEXh0qUu3WQo7Zlnnc3Z8PaFoXPpdA7gDw1I4BP/cxRr495i2zzzC9/7E3enHDa
LXRMdvPa8NwsOH/3Qedm+S+Bp+xmgeMk842NSjhQgyrZyd3Z2LuDdFzoVgY09c7E
iKzQ4VZQXKVqnLZXZ7OZm4REMax8RJ63LTzZInsvoORrHi0vMKySxKY3EpB7w8zP
i7KfM7GcI/6/XY2rAEEN7x11mDrqME3xXorwam1vaOJ18F/bxxf6fa0ss/Um5Wwd
zWFOOXSEGV1WxsR5gOEnuCThyrtgVRFCV9qFLgFQ1MbFurZsg+qu0AmFFSPGTGJQ
QiGRqEYXDcpCJ4ngrJfdJUAI1P2DIt/MdAdW74cCAV/QHgm6fx8JZbyW63k9pC7W
5mOrKkpjMpH5a5+DLsBEVMULVhuHBd6EYjU+vRH4mXPMB8PIi425zK/MhPxvsX1t
clv1mM1T8LAdVMpFXU/G/4vipeg30FDZh4GTyfuaC859/mY7v0oHM5PoIwYFAh5a
KRfRQGcQdJ8Zbi8LjXAns4Vsh2q8MhM4/Fd4ppwdDyuDP8UTUL00D6NWp7N4Looy
c4nqjyWb2LvffhTKXV5sYUwWAv0aqljmFfvWScRwko0aeyLzCGTlcGykNhtD03Cg
OLzWJR8KiieUlW84RK/PFYpTVaFL3I+ItpZfOIZbBMSUbLry1ewmBhAyTUuahcvI
mj3mwNFTkSfZHiYqSq1zjymlbMeVVelaZBbY/VAltpzO5qywxaLSPcdvoSvWToce
MyqVWPPpEoxHASEo2LS1QWxEvjLT0GykOScd2mISaZ7v3UP4LgWIzrilPHKpeR4F
GFxbo2YmkKlHO1q5hZn9nbTy3GeXghX1CcnA7fR1D1kVZMrkb/F+sGMNlKkZzNT8
Gr/cmabjHR327ZPwh7QumELkA6W8zMX1dxr6eR7XiJwVRSqZW6Nvzju24MlRAU2F
rjBARngGofWBenxf5CWKNIUW2dF/FKP7XrRr1Nj17ei0usMUYYtCdp9OEL/I32Q6
FlG/npCHoCshr6XDBCSbEm0N/Q2Eg703eqkursaohIBvdNnC0tq/gEV3SiS3jDBp
QLUfLfl1MYEU9ON80WhRWfpc7FYK6NMHwZXrSL6yuczd2j4evJaQziZjv0rPDLHK
aEf3PPJfRYm6tD66w26qpwaZKFQ4P7eRT8BDeRopiFr6LQpDsnl/nYY1aGtqiZUe
PhmVQX/mhiAGRNHDMCHbe7bmEF2fS90qn+xb+6VUtkKvED2OONAp03hBI3oI6lfF
wvW4BreThtiVKh3iTHIvXDkI96cV74M8tJm8E0vL1z3tQt5lZeaChdWlgbT9hLGV
1EOaSqAGUNVi9mO9uvICLxWuyzcIPrIRemf/2SwRpjqTqDO/woON46zjFFKwjpM4
+JSV28rt1MOxUw1hILi73n6Rao29BEhWZdJM7Kn1OIkV3u6cmuY9HG0wHj1HjlfU
nx3XrMKlOzJYWiuD2sH88kdaJqxJTMNUck3TnOBmz2ZxtIcvKVT1ii0kLj3ZhyuY
Nr7LmrOYkR1r1YtLcZo28Uk8cM4wdzGIJpcpKxKlUWe7rdyQLIhwcQmYbTLxW8qL
fdPpG6RxxRdSULPPfvZdTXZx+BAvDmTurNjFetl74Gc7bmeYSjS3HrM7vZ0v2mvz
MfvfjTZXIhjRhG0x5W7YHVqoOpbQqJs7PvqQugiaf5cvFOAOg2dIazo3p+GCAQzW
Gu7ED+e7uWvvhq2lj6jynB2Skl9nj93Nv01ti+yDN7QOpXL4D3Em328ssG5xfUJG
nrIyIayhoWI37L/UPvHEgl3SUF3ayiZl65t4BnUzuU64hUHtwU4s5+GM0URUvF3C
FZSz82H9H64cQ/D39B7Wdv+jpcyjbw/NZ8WFTmhtYDUxqrsLCdpRwXBhu4mhXsIK
vOuaBqZyf0igoY8iCmPNtipNZD7UUp0jje+hac/4ix9czNZc70NZu8L/jH9YtCIq
RzmL+KSYvOAkTboh7NSLRiR9r+iyytyw3Tfawk7heBjn6M+YCsSVm2P5nKsNE9NJ
wtze+FUl93EYogeA+o6HEWxsAWFJNnvRvS/hZlsAS35qkwiUTysVvwGDBKzTbGm+
HdQro+rSw50T9HtbCX4yBuNS8eVcXNYdcn0wh9tUZOzGAYBvm3sxqzw5+mGX4Ef3
yNhiRJUQbK8mkXvC82mX5JOQ7z6xsR7lu7ceDMGQGo++BpmxCzXM+bX6OB7PpdXZ
H0M45cjnRJ9XVRtGFKBPDVQJTkxnKsKWnkw24j6WhIvh+zLtUDZ5x28m0T6Zgcoc
sbSohC5BVpYv3uA1Sn89GhRYzuKF4JtNmHnFCqnTDhvhDlLnLawYVdLcakJlLYGy
Lj563jC1yMHfCpZ6rX7iqcvZlNf6faWc4dye99PsQPCkA14Ev/PAcOjT1NeP2NAi
Zt4Cu0Nc8WjxtU6+WHI5TRE73piS4RZtQ7h3N795PfKEfgfbWlcfd/FTF7pk03sd
xaMar9D51K5G3gpzLdIdEQzVfyqe6edauxekJzwxXa6xO3Q61O1LmaQCujXxh+Mz
GbTb7p4egHojze5DXiyRbg2+JDLXp+KRCX1CY5jaET3IfYdApM4vXgQjlY1Z8QiL
wpFrlBWrAde2Ru05qjHy5hkkUl50UJCa3uyWGCg/eVK3/XEqskCigIW/3MkRGSn9
oUB0GPvDmNgub94QTSzHzFqesx82A1h5JUUhMMyWkC2GUBrkwss8lYfewcU3AoS7
9cyk+shlOuNRw3mrRWJlUPD0jbLgckigvlDIGTXcSwp9H6PF8W/E1ImIz4nPlnei
Wtha5fSmDjHkeQcmp/Jh2IC31DnhYDpRXHpYTCRdxoVOETXLyiEmTtxHrDBTcR/P
nQalo/vy/Z5Bj++v8oNlheNG9NrgWnL30q0Vu9qVLkQRqIGj+HKZH9OAZdDRAPmz
ixe+I9bomtg3VcEfLoFdtio31vAsK1bT4x4jPaj1K9blDgrwe3CvLkt//wub4oKr
AmtXUUNs/K4PSRnQOa31uobF2nEkXFNR7sSpL0kfKnbcQrpc9hJHXWruMi/BtrfC
FtL7HRyqZMWB3iSn0Levl6ScD6ezZ7DXTEAxIGbKIhIKlMeIyCi8fiyUWmON/V8w
w8tWhAI/bjmWt8t1dSWb4jBcmevXAH3bHhvHhmD3pnW7+/fp0TyOYUDj8vQ765rI
eIh/pnx4Pi28sI45A1jm6PPvbEFlNmsj2kEb0QiqLyPyHQhTwWSdxGnYE9NOe03t
ZGbjJ+NptL7z+qiNTPuJv+nG9Fc8lwgDV/UA7kgOyKgcf+KgyOpg96QFUJi9hQis
TlmHU4TW844H+bN4vRCEc8Csd5vYE9k8Tcsncmrs/YPtPZVKsJaucpNGkgXFnS+V
J0nytc/4a/q8VJMdLt+L5EjGOmoziNDm3Iy+6Ylta+UkA1cJkbe2cgoFfNy5wzbZ
QB1tCkZrb3XpNz0j/MHxkaGt7dZs7VVjEpVEpleILt4i9zRsnlWj9Ussfhiw2HNc
QVElE1VjOq8tWvCUzlQWxiDkrDJd7eFzPF3lJGTkBDWe3q3Zp+AEZJDPe/8o9opI
sddr7dqe0N5lUt8j1r930aZET5QwuyZha16q3sF6zXoa0L6IKFLZdfL/spyGOEfr
P1linVuCrOpON0XF4Iw5KYSgzBMhRw8X7vdbUCVirzvbhejZJmDBww42kmjHCVPl
E+khaSyzj6YZJe2Ii7rIRu753npbPo0zVnA8gqq7nxzwWWml3ul2A6LM6O5OQblu
VKN/Esx6YEbzlgZGYiunsCb8+6LK5oWxiiYGYJ67oAlz4+T6NoSe6avg0IxDAsS0
SxUyMwjTHhxwZn37vqx9GRY01niTSimGNro4FVUXoGByLS/M3vZhppoPVxlnRhu4
z/xsViE1y77PAo8TJYOkdeoFrAj6KIrQxy4GbnzOcpsFLdT6yTFMMN5N7EeEbVZL
+7BtcDO8j2uCIHDlcZVClcd/QDqk4fnhIc6QM+ucTevjwdwbbiubYgDo2ULJWwry
0FsHRkQ77wGA2Y/RRGIMjK6ZsPXoY9eXvnRtV5sR/PJxWCXmXwaACPs16oi8kZpw
0KCX/T2p5aHSeuKArofXlNa9lzZML+Ebqttr307R0O5TeN9FOVykJtuM83ExMt74
+OWQvfeyFcEJKSTxPyQeTsYxcTINn4k33ROm6zw2kpTqN+sLlwHRLmpOBWd082lO
uQ2+C3KKuarls8bNmIPEG1DbLjjqAxnzuYu15jkBTFxvy2GYKRFUqFVO5W3okXFq
eUEkTH9FUJVe13uJlA+rgIDm5+vSTqzPrGSl8qF/WbJwmdXy4SBh+ROPLLlaGesD
ek//el8wE0DGwBzyHNkkCqitXm36GUJZ6oBfl8TYs4oH3e0tx1RspvqGDc15ttU3
hkIp1q2ls/7nLmSTWkn/tjKAh+eJU4leKY+5IR+lakE6iwRRhcJs8KEUY2uhDg/H
QYVp/WgbysFDNrRKoh3bez3DXNOH4c/LohfVr+xI8gymQ+Odr3M+1vihWiOHqsfh
HkDk+xmbBpRX7y+SYucpYRbgQFsdrcmsqQeJeuGpMYwJ5oaQLjrAc2l7gcZoaR+1
uPkKqTPUfEWx/L4eprOCHefm8mRfUDTAxn3sy6stvZ8vhkZJU1pXFRfIqzeOOKKJ
xVahaI1nBF2CTvcjdrEBtUWoaRH5jh1hOV81s7UdsUO9vBC28Nxx1I0lAS0JwJCi
Z7DKpBg2YG6BBNgQw2DKn6/EKWhl1QdzAAzTWIBJauygE+oU1+NTf3AQRtvXWwZ2
h8nuo8HO7wb7jsyyL1VPND1qHFElv7chla8JPaxRmqLqZYpCDP50PQf1Tm4gqIgT
f+3u5udmlEw1m6qK8YdhhrXGexm7QW+j96vXkl64sL5MAzWpB+ATbM+Jn/RIyfMG
8T8BScTeyatCvcpV4/adC/M7HVmHtbYNzjUZ4JCZuT/Mf3+h2hNXIlogIZOy+/h3
0edRIBtUajxj8CUq5FC1LWaTFifIDSxvMFwHOuv+jFUrqP279WqydUwhgBAhrZos
ONlo4EAOB9YCX+6D8Em8coGtHcM4g+tETPGEXxNrfTOTlbZcNOE+eVfLUO7uQLJd
2GrFHHyO3wAp8eRvRTrepJkM/8JYotJOLxxibISuWJ5E62lp54w3OxbgHKZDkp05
BBxXN9xhcRK9Z/Y9OYfCAEQ0qIf+SgmdPBrsjRznMhfBlblpAODgEJSO5kee7iES
Bzf6HB77/3xhYfE33kWVEdFrOpbDj5PPIg4R9YU17kSg8sIcEvLFGFcff3hX+gM5
ZJlit+dHmt/GBl6HDwjoFp3XUihrpUE8E+fQcxDBBI2cjpzPM2ubSB07HxIefu9o
2yVhV6xyOdDze2vNgzYI7AAgAn4dLY/3DbQwFMv8ZCKHfOIC/hk1g1/wU+l+xiJa
c9cYeBmaANSnCIIdXg6EqnupMvQi8xT3GtYZdf5sLFQu2RGECxT8VEK+OnulzNvq
z6ktF9IxB3y//FRQA5Pm5O7gUEOdRQ8SyrpzmFOKMf4P2XAaDuSdSLo7PpScdA9N
SJcAvDj2y9HmX+76gdN6wMMEtx0+0glcB00xf+hWrUnujGHhAONX6D2U7fid1VsF
+3etv1HHIGva9ieUGtoOUcEgSv9oxiOf4oNTtQeulL3eO5OXQrctwSFhPX6mT60u
ASAdGhXAhfhg3oEYIlcMFzFPHG+VkI7/2vbP02z2rvODxOFqLOgDgGJVMVz4vvLz
OymYIrEIsVHcJK3pxSJbTGZjvB+MMmz6S0X6izzNQ48AYE8MimUmkbsxWhdAZUOo
WTxgKPRkip2mTxCZ4uhL6JKUNsmhbCFCU+fWMJm1Cba/gczrPoxgDQKEHYryyxJa
NRB5IQMP61FfR6uMgAdTIFEDz4bpLdurEIVOtyarsIZnBLmpvz/qTYFCHSxYliU9
MrGx0+JVZXFYNmxuewB7fXk6EeE7ElzJJv4Fm7ZVH4F5S4skJkRMh7dDVqQBp8wr
FUfIYaj3sPxjpWoYAIsqDYTniI09JuFwwV2CJjG9HXZuwh8/CpgC9Xwgi9o6eITE
K5bduMzJsEOwljmVgoxe4jaQYMTj9XxgviH9qiObX3KGJabO4NmW0TDhP1GMkq+Q
VALkqyGfm1ndOPcBY2lyg48VoxqmnOLQQWqekAFh5A/lVpv4bp/HqgHBzA8dHHIV
PTTPQyyjAM/vSMladTBWTlfb/KkClOzm5L3vELJvuUDwokO+s4FQA3Ib3IZeJgUG
GktyZEJhkewhEK0Z2S3JsIbILQ10CEnspyCYD797WjucNzeVJ1r99Cw1LYoZ1jIs
0licgsKyZ1pBOW1uZt8Fc6RWy0kY0iaCWbZbVwI2EBu4elFcEczSY/FiSo/D046i
sCnkEDMRu24AbT4CSuG/mGQZ7wLqwlJiHwoDPig5lSa0haYEY42bpp9DI/xCgEOq
xwK2siy7PJcuirs300M+xpFjY96hA4UIHySD+do9/qzsMTRYOP5N4o+fJAd2Ita6
Wpuy9TsX+jqxlxPMbMb7GYcMX+bV0sxeGI8HLGzhIZmjZXnTKBKZOHr4TcwdzUA3
pZZRxbooJKCgFbjYe4Nx3pZ4C7BBycuS5Zn0NZ0DFRpZLrz118ovASIb8YxK9t9J
g3CtSobNeWtmAtKncEjVmvItd69+xw1kbpuvwiGnoSsYEY/Jpfn/B2h3Sygohu2Q
Zs1AkNJfM/KYt1uIWeKcsF7lY6JLsWR2pBLOutCHCYX3vk0T9QxIHDUSe+QiIAwf
Wh7OK1+1mGZ9TvVM/oHGczArs5A2X8sfsyum6FG9l5tX3iYGADczKTWCF7zy02CN
lkf5UySFKJK8/rQxJ07oaunJLkN0f2ZOwS8a0zixDAMgv7dgjkDwk1SKFjG0wGsk
VKWp43kTSsphTBjdC3s7lcp78J45387yDeGtY6/Pq0qCn2aCqmdPeZxHr4ACqLde
18JuC06ozuorTeSXSOJIXtPHS4WOPigHn21N5k8wGGHYsFacqv6pv2UT1gns87dg
nH04h3Fa8pvCTS4TaZiX//ovpBoul71PDchIcPNfjct4SZhMARV4vWO26gx5lz7/
PLc3i6s9imvqht3PeN0YkOXmT7UVA4FzgF0Y+ubuPcZUBLett7SB4yqg6wlqXhWu
ZaUDr+up0ASikKYoZaSnXMNXGO2qKsNztNoPuXwz9o40J2xU8u1zBjbJ3T1pBgA1
ibiX5wXLyJWt+tiVNwJtnjRR5quwRjESHd9OZ6L4F/9uPLETPVHy2ZRV+nL6qaAz
XDsWesNjUu6iIVcIRXntDITHCsWoW69SHfrvga1OOaZYpUVoHTXhc5BDUUWNZB2m
2aocZ9SQFBk6WbgZwmZfToWzfWXvl3a3HYF11dZnDn9BPNDo2mVHZDN9bcfexReS
Us+0T/+cFxXhTSs/VL2T1AYAkL8KzLvcBhjcBQlGgv/8iGYQ5wzf/YaS8wl9rhHl
khqDQsLW4+6zHSNdzgJQ/RlQMQ6EoJqgJkHiNE3n97y+an+1eKhBvFCT1msB5C0G
gv0ccAnPh9i0Sl9TFLhHEg1u98FJVnnvAaqPKOE6PCsQldo3R8x1hd1rjxbHTXI+
lI7N3d1kNlZpdof2tAow6Lwpeh7TaIhI45XiXKKFD3loJljvrBjDkFMer9kjH1SZ
T/MDCz7/VTJ6iQq1MpN8q8M6w1soIhjpWiF3dYqPmSWIl8QORJ/WnJH6KDZQ7Rj1
9sw/CAhE3YGRfIZ/PDBhjDaP+hFmlsae0DpisfvMT7XhvJ4HTAxhFcllszt8MKK7
vjDYknkYNHjJQT8kn6+rlDEMjOb3txcwUsXrxEO4KqvcoiX8+eYvPlYYKECJ+IaR
1xhPx/dBAV+Bw2Yia1o8bbTf68vWcOe/xLzSEIpggKaIhx5ByfwWyaCCNuWrIquM
S6hzU2Txb1TscVQ1G2huXxa81RRc7kzNfj1FTHwu3cx38g+1NvciBGy3VkQjwQ4U
M/H7j16IcLW6pvgBJk2jpH9MpknqhMBdXmT6lpsYfZ0+cbkAOovTLBY6hVdvLYFz
NMzOAlwN4fdrGw3pz28gW8jtjURgr+OENd6LCWcIAvzeru3EkgUdps0H0xdRj1T8
V9tpm1dIjw9virw5kNyR5Q39r5pDv1cYZQGDlezCOtCQ56C6JOeY0pXpZStrddw4
Jv31zPS9g6npyff3nmNy8DCY8JG8rHEtt1pKr83c0QQ0SlUmpPZ3UToO5Cox3WNa
L9b/KUuIu+CRrInN1h+JfOJz+M8SltCbQdpRn5WiV+8tb9oFH/RUnhi3ona7rXag
K9g4VNYYSD1bRbvJUpGQ3ngvdZXbFMIdZuI5sXvd2HogMMO+tRaN2CPYIl+ve3Sx
wOdXZp1QBLIjIWspVLcHFb6cqlONIiH0F6HgzSaacrLa0N+wRB5nwPOtFEJX9h8a
+o2uS3UpR/c5qrxZNswQB+fUyspa1QyZ4Lio3VXfAkS5AU6JB1vQ6q3T/3KbK14A
YqrMOxALgkoJyKI64Qgo7oj1PowJgaG50mKEWVRG04NFmoT52lhzLx/5NGwbPSdt
HygyKDclx0E1ib3I/j8Dd8VGWksbGnex4sxFwXZDYrXbQ43HU0r5iUQoroawRSeU
sQORalPPnye2uHvlASEq8/WNBJozTU+03lyHXFDXIK0+C0hoJKxPzoKACdgRU3p4
sLyh/uVR0rENZPTbwar67IoiHhZFdxAFFNeEhYwmH2zQfrUv1/MgQFPgA2++PBan
4fMh+D6rA4uuXGorM2TRl+wV/srSro6M15E2JjRK8/IEsjnvZdCygYuO6tMNVuhn
RWJFKsb+1ovoU6WRVy4hN5Lq6lgUzt31zwx/xVfPVcRJahoHl1/4arwVi+IWSZ3j
b8qcdu9Bs9WonUdo6AXNtpflmET67SY6a0rHNMigmisLB71BEQkNzerOceOR19VF
JU6i6496XMitXuzYKPSp/0l68TzO53dGYIWkUMcHSPIPbYDsVbxuh5KH27+pSfPe
kLv8YM5sWEeSdkRLdoSrHkQ5pG2NxnPEiIpSbT4WFlkdspDfZ8i3D88s+OIXnO2W
yKgFN8+1AEGoXE/IF7C7Tvm9f54BGbzKY6S8iQrCIznrSkhtboFv4hk/aEs68QKv
zz33wOXTr+xWFpqh8vlzg79mXWLHQcNHQVKFGpbkpTyPeFhOm73nPKCCnN1ksVH7
QUxXC7Ydu9OSmxp+bx5ZGPmTsfvYBtWPu3hM3T0Z//gr11Wbbqyjbe18c1xN0LJU
KlrL1Gv+aFa2Fc9vHMG7llcSms9AqRXomK/c95htJ6tOYWPrE5cnqbI+nGB6EGv6
ZyeXVFfpWz/ChUOBrQiAtzzN/L19tMHBczJ5Ti8HY/v/EPHQiWUzulp1lnM81+w4
wD62U7RW+mpJTeBfPW9F+gBZTZtMa7iP///vFV8JgUWnt9skCgdnVo8TLOSGju+4
uVQXOIOLeAuWICiF+NQlho4EVB9b2rNIw24RwLPCRiimi8MpTMcZ5YSJytbR1Iur
FhAciC0PvM4/pVJnKWQMmHTh3m3FrQ4OcqIWEYBSosqGzTKvj5GeS5Hh5Qcvk98H
dcMZlB08L8AbbM90iM7CZ111rO0zP8Fv6I7Ktukx+2HUFympa7aczttxCF47XS6d
X4WRjk3nPVCEu02TQ0MQ6SEt+gDy6fJ6CxTCMByEaakAezJ/aFbiEZS/3UiU3vRu
+O3XF7M2XZwY/u5PiVCIrLVBfNRIrHUj1Nd3N6DjAa+SIpXQn6Vg5CASnDwwWZGi
B/husF9NdZPVvWS27fzLX3T2giUzA9NB26f1D42U/1Qul/8bbqtxq6LX/BYNByHh
EXciGpB7U1CDl5lyPh8TY1+JJFCzRymk1fpF7abcjVcnpoquAk//Z1osXzZkS4eb
9iJTxVXIidW9fVMvOn2pYBkT9r1neFwxhjK+F7P25dNCxH1EETKdzlmbMbn+02r/
M5/1141D3lPMBTyH9QPiF1Gy5JDnHdVh6xgt3ofCHsD3MfV/rX/IPk2gAUkKKU6u
gKmR5cgu1Awoyvqs6KlyIFpKxNUK5rzkSkm5kpD7ir4oDX07R5l/HgWTSQNL05T4
UCy7DcMC5iV7fRopaCENdtQwp5SWwdP3pJdipSMzXQtEML21/qKK+viltX5w5Yup
MrEtlCmiBv0F93/khV5PQwXxnfSrjQqJtVW5yFyPRLxZfFDxlA1rxr/djiEgdH9H
gvQ8oEdABaZ1uuqP02lzILCtx36+svtcyLKTwNDsCdOBWYp2KtbLKs6UmT9rTXJF
jUhj6n3vAtcd9ionG4sxc4PoZeeVoc7LVgP/TFT9di8TN7SfGHtXrwt1X0+Oco2b
67pdkahF32ZCvjoEFHWhB6Y9urP4aqXwRnUovY7/oapsHu2dsv75R5k8hSzjZCz5
DifWcopFXVUubnwOUlzp/hp8lktc0BthIZKc3FfKbN4/u270B8WzNPzOicVL/jXF
X7srwaTK+Dr7u4RRslqqu+Sm260aLcfGDSN8QM6+iQ2Gw0EfnMLvzYcy5c3LJxiI
jQ1Mb3eFQtd5J2pRR41CqBxqDA3w+/KIoJgRflZlCZmgHb8AYGdFuqNtKcWyIl3M
Ao8Qovrel8FYTne3rvO1kQpCr1Jaad9anuXRZnjhelrA41I41DVgb3sqfIJB7rEX
nZgY+qWrGSw2w5dvnV52Jbmms380FdxmFGLESdZpJlpIM6m/BlJk8RAWO2Wfe0Af
KUfBFBP3B3Kz5Pr/lgCfJZztxcb7WuGlU9pNpKUGOXMt4h99i5IMkFhx9ek6v7eP
st8TMQpDC2UjyM9OLN27ccHSd3vxjMu+cwfPG9nDgQHFMI77d0Q+f8sf5Qu89Fvo
uSq0c/mnlQz2AWcjH/M+guFCt+mhddGMFFMVnrzJHhBrEInan26tbAGb3nYtIbIy
QqPb2vzpuJG8Ow4qrCyjMAX2JMjD4NXoHn0mrMpDRPiNkxwM4PNNFyROA2lWddTv
CUTLEBxWylSRDtQb/EX8hsWu4+PDOaeKsr5BbhyQhZiAtxggfEsGaKN0IEkxMjaU
4Ess+SNfZxDtcvvSkrjphH/glvAUu7yUJAH3h4ixANTyZDTAva+GkwADrClwdJpF
iS6jvZSwJlkBRBrKlfkNKSatfD3KwleYxGMbL2Ks8/FhdLL4SFABl1s1hRaE1D/R
9aRW0/12bXPwssMNr2o5rpA1AqSQPyrwy5iC6KXDDCQcZcDnNCjgL8wRzKYrzVdG
E8aSKbXQKCrtZbXqSQQukCugHeY2oG8Hy0dHWsVOr+R03yF8vwCcmU7MEyaPEgOT
m85lYCkC9za6DhiaJaEgLGnZgxY3KVl+FQdsbEVvInj8nw89vw+dfKSY4iP5ADln
NHyknwpyvdgVVAD5YMD3N2PGgm9saJBJ+uqOVdKV2+/qWGUIAqoUz8ndD3iex1Dq
sdaJH567k3lwBtLskZO5mNFQ6GGvJ105kQfs2z/SH75JUa9SoHZpm7OCAWPcrvH2
P/Uoj0Hm3qKzMHin+mpgSLYag8sg5eSKLLdoyUuNj88lGa+07m8sAwOmAnQgsKvx
CicAi0QkUEEl1bSV/rlPXIMrO9XlOs18865uP4OZPFAlE3K8hYr1lb+ImPuW7wcT
3QQZBrtcccTBDDu3/OBKZBCNUERmuDr3vCJv/V4HGrXh02pNHElMWTFd0/cDybSd
6oi4sX5tzC7yPEqYtQ0zENbboLWD+nVgcsOSOd8Mv7yNxfqEB+xwqzcnsfNcaf3c
1N5/wlJlOYVplJVJEo41kE2mQrf5LAeDO3hUcpYCfTl8iqUEzd8Yy5MGUy9i4ivN
6uqaQJf5KD0+USChZhztvIrvnsTIKxODWOXTqjl6pWW5OIQmTSDrxx4Nk+GgZRDF
Gy3ZsU2YebfNn0FBZ80OiPBW+MZclT9jlVqABvCsJqk5G5iLb1eAdUwsM6RDTzw0
f06J3PswOUCD4jcQeH7Cwobp9DmxE1Or7Z3JWqqT2FnN1aSnLS/wM4e7s86pIoM2
c83Hz6Y2HwmDmjTE8dWy46bir36GPuWXom7NHbk4as35dnGW5B4oZkvDnisgWfxf
BYueSCf4EzG945v+t/Gqdwyq4+H7ZoljLDzIIhlj0JIlVdQRH4VdA1bMWSTXCNta
ybbGsHDZ0Fro8ABvYXVLVLJPpxgO8XskVIfRbhJNwTdUCK3xFsfyHS0fsWmoS94F
IPLk5okR82H8d6pMx9alA+26ngygOIIo4t9wvrNCia3QidY4efTcSSzYR10ctXfL
dEtr+l3j0PQHkLaGz4Qqq7EIoPbk1TYHybcQcTrAnRgyGN7u6LHiFMLmuyybNMVp
SgCBJ10kus7j1HZZtY4oKUD+TsfZxjiloUArRSouK/P28r2U5NxcHIjhubAVIdHK
aMzan2rqK/1mskZpHQC/vnsy9bC0Rpk4XT5vQCI0vIlczDsIgxf1nqtK2ZbZfl+R
/zRWgJqYReLvb3witUtlXCebaKFumW9DdZdSeAvA9/s4Vh0MMQXsaor6cXRxgt8O
dHUUFmKy6459nkQvffCKS/hrl1nXBwkTyYrfimi3Q9e3goFborfHDx0eMmDuFGpn
MnTUKG6iM9OXsAwuTYuOwg27UWGTPeIxa1/vUJCYqPhL/OrZ5Y9ua9GQHHgCL81W
F073c/ZGD2BqghvQUbFAtgaI6GUuwTdnQY+MKKi5XIP3vLyDCXSxcST7hnYY7jgI
OlLkwAvNVDWRkhJew8tGe11iJjzNANUwXzsftOtAoFFfltWEjtxVcdPGgSkuxvCd
hHgnIxXOt2GSEoQypI0+7AVpYuVKTHtc4fyg2/BZ44chEaZ6Q4QhEJuapaYk8T19
6sZvfc1XtA1q3OwswKLGtdJEerleWwiv8s10XKE2EjSmX2ScRh/CKMKo6Z4WtpXX
e3qDEKjgJyksF2xp+2OO8ST/1isPe1v7pibW5Vm/oixiBpxl3ezM6Trh9nuiIryT
EO5l6MUGTPfyKEHnkI0SdSp10LU2okjmO21DPZN77hJHmP/GNriwJ5dhvkyi8UoD
R8e1XKIx0AFORaK54P11eqIQsLJKEH20n04XZ2ZLoLP3KNGevKvmK3YyiotDRnO9
ZJqZHQKjV9efXqRozcMJwlzLkW5oYMZ9wtEYvI5Oq3VD18Ph4CZsqQbt7zIw43ST
gVosKuH9e2tUC79YnKVVNApKcDsV1KwoOm1zlPeohDei+PjGQrnzC32vRPe6Ybml
c0cnD4okqNJj99WttuwBNI+uXOyiUrhE3NpvX7DU772xZnmQoQ4/PwOSulwRvzPj
++5MCRwbY///HR5wf/kTd+0IHxIJ4LjCl6TCUHR0q1yBg6BXBvrGvNtZRbWYDc9c
hHFE3aeN1w3B5iHCH3kN81rFEKfHAB2jhic6mo+UYd2nu32sbfVavOrrAYyYS/OE
XFyCxlJ+m3ZPuenNzSlZhA8mBXv9Aui8qGGJjfSFc2B7uIg8xxli1+gGP2aNdUYo
meSIO0C+Ieb752t5YHe1pxQlwl0AQmhIvI7RDMbJ8h+SffVo9PA+f3LoUHiAw4Lq
ne9vrI9NH4IjwXEd8WPQVqudWeK9gcojQGtPBpCWog8yM3bU4qBOwatJoUWQ4JGL
RAwE813WJAl9+Gts9lWKBIGWDHSKIdpSL18p1eDchhtkTAiWcL2KVhWt+OsF0mC1
0mmnr/XlsSM63yDIxR7YKYVTnygY4t16XH2dVoKpp+34KBIgnWDu/uyueQ3Q4mnI
PW2bTI9bsVRWnrOpew3Qp5E9Xveb1uruCWPAvm0U2A2nd66JNG72ZM7llH8crdsm
RJoSTS6Hmp6xq937hmLRG5DbNayEocRA5tHdRuYjVMItp+Rds/vdb4y4VpJOovrU
IsXKGgbpxJ/pOOldqdRqLxHE6/BMMEhwBVer/BFyp4XvByNYXqvx9ZbEGvMdZzl8
hGR5I84vA9UVxCJ42nDskGNQEwexPplWYf7EKlmSGttTrOpV06gbzqCAVybm4WBS
9n8gW+XIZeRPtOn9rErwyCfyY2xsQk2yknq29jGp12a5gQR7bIQiW0NHVAPXz1zt
IqCv5U462DxO5/EyGr5Ku/XxUy6BDAHLeBZISntSBiG9fW1BVD6cFnFA8Dj6M0ZT
ItTMAqyyd2Uq+6RA559aRwVBPLhtu9HacTydb7eP6D4gbKdRj0ek1jXOEzfOoDUq
YlEP9klGRAMLGN8+feB9jUYRmCO1ZvM+lwqNPhMjZxHYIEgdYx7w4tkEYK5sE981
SvZma3xbFZNbp3tfOXON2TKJWxnmF82pvzCCzEN+ukfZgoWvW/P5i2lQBRvLMNVB
xsb2AfKx6jYVISuxEBYZbcpoCaUfemqoMaa3Zn7vOBAYVPu777dZvdaDD8I/chZ4
sdZJdBQ/ccogAdKlkCA6hkFFcFFch5qeBVo0ZpL1RT17ma3tw+ybjvBy5Vjc3mi/
gySGET66SmhWTSn/RvtqiOkBPEm/gd57QtlVLEIlkbw36UG8/p/nTrtsqdCz6AKV
PSfN63bO1G/VdqA+HftzgLlAUU5CQRmcDNRKP8K9jOOoUmVFpyY/AhDXeo28n7dl
wXNzwJowK5c/tatODkfg1L3G8YbRj/3hkpeuivXvb0VmOt6kdenl0XQKm5+6zLPI
PUeE2hilNUMDqfWcg3Ufw/VfF59ha27PhkSyTDSe+n+HgRPvej40OO0I3nj7avGa
I31zR23LJN5kqb0Snwarw9g6DOViBgjGQ3HJSh+Y7pLO+/Te2ntSDQMkTSe9cDJd
lBSYoyF9YweAPZxNeD8wVIMgmtRHQJv27pLErRZI2BOVk9qTua4ggyAkfFcZ/LuA
zV4METTGQ5WAoQMxljLHlFa6Jh7jczK1Zdav6hyMrmbTtOBtPDMacL78IOMHAcut
X9WQOizX/VZGUdMFYgt4P0n/XUzT/SYDbBEpv8hTm3onl8lVPJN9dP8Ps1cV/MA4
+oHCuXAyYiISPnpHmKuYSMcJYX2gRnx/ZHx1SBmxtcm2ULPlh/Gki6TQFbcBOmuZ
U1PkzOuPXs7K8TWPhhy/DHRzmPny76QlbTlVKLeUnSQP+bh8SRE057v9SO7LCR1/
VtyTyB3hi491/sDKSHpw1tDRFC/nkVQMTmndRollvj6d9w6iztw3f7jh0ZFoeqyV
FvH13by9VqfxfarQfc/oLokxBn25oWF+aEE3TdGpmsmED6Cvr6sGtKPMufG3rvzf
yM1njc2Z8383P8PYHJ5y06gYRghh78ea/RmbMDusUZx7Y0Yqk1hOE82TKIa+eDNx
JjLpCPlDJhL+gAhiSwitMqPYhkhc5wvHtKBYrMKWRRi3YjG+9A580pCDtk0RSCqT
+wyP6ifH1HF31JTtcK0n2qRKcwO+WBarvFnvc8+v7h/XlM5OMoQOo7aG2djkVWWc
jclg2XJH7aZ8Wssa5GzVERtqK0YneLY/BDxNSOkXTsh3F8/lBb6juyKb4F5n4Oxs
PJ8Q81expToq7D47PQjmt4CMX56z+4hRa9qSDDB/gRfYX+aDznae+oEhy4hUlHSe
BaZs1oWdQlouGlyrFnkrqZYlDa2u2Zcu7NFnGcG+lpK/iMzpggMJWCXEbmTtXGL2
j+NL5iRUxVAZ6pzIfVBkQpPg/VB+FaBwp7Cr2JKG5105AaSc0j3adjFT2s4NKdXe
SoG3VvrY+xlVNU2Op3fqGG5wDPNNY/Oqe75shlINtUO86Bk+CmPGtGza2So8Git+
/FETt9U2cOTnXViYb4XIbS4T39GNJIeKyTs7rxAW9gkWHUmSNBoFOO/FJ0JRrN7A
QJPTYaL+KXqVf+7h7pIoMBNdrXUKEXtZX/SFBzFFawOuMrK0TumyGQbpOAmhsRAL
8cyhVFCXum6FR6drrXFkPPumG0a1fxiivGYcoQAZrQX+a0NUcVAkvnYYDy+gg9M3
Bc4v+jbeuLfPoOcvkahakL8A3k/c23RnXS5fKrEXx/mUMg0pBPfvp2komQtBJDWA
G0PLVBXZ0XmPHz4Ai7xJb9yKRJQX5nFwGlNLoMiuzVI7k65iXlvxEd0R33U2oiuY
1YVHxI+8jlhBCvMJDemxtDWlXscNwhAX80jpJBhYDF7ZEu4b3WH0Luwhh6hHdgOZ
/3nYNPj2G+It7UKlyc22h3i9IyZnfVM0zUTTFX3pXxYWKVCD+bo1ojRDOONIYWJT
LERwTE5TAamSsf3mDKdFGpwwFH1WhHRQsLUk5645Sf2mr2BpW9c2SbAb2HmeVKAm
3xuVKPibsQOWXabY7PZD8bJ2/KhVgSz/A6VUSD1B2SBM7PNukziIbmsh5Jly5OKW
yiBCShCwWpStHoTahSrOJF78pREBTpDSE8WtyM3BOuOd6haeYxX4XRqkQmkTVPKH
p8/wQQzNkn9Evz60I451jSybWL+mIvoB7EeTpg0A8tpgGnKR0BA0z3f78b/sPUSp
Zg7hahWzyGMyql8lEU4EqSjyj1GIYReoRBW1gRDp+/e97zs1KCa0pKtktqAu2VIx
LXKBH1XMyQVfyERK1jhPQsCtHMO/eSdQS9XqMRwUgauK3JlgwvdAIzxdj0atDMjw
9gt5AXkFr9ByutsZRtwXirQhafAjGW/uu19W0vRBEeEVnHkT51airYz0feAb8luz
L4RiGHOMH/XG297tU4GyY6Y4KQPmoExR4xOtcJHdlsqCj89JkeWsR5hdYThN7xW4
EmE+NTXWPkSyUUVgVRW5WaT0ib6QuVbeHhPhuSIDgHwslR+XT8tliqc/iizvwS1W
LGJuZ1Kbk9P2sZzt5b2SbWc3MBZGHgMxTaek3OhQILYtoUlnPYzTYD2a7bYB7rFm
zVHQalyLrrayhxjHyMwXgypWR4qv1VsD1EQsMb3t1O7VvILJsBt/87m1DpOI1wfq
gvWMmD8l099wOq8BkmEshguh1H7uG2rOJKBaKrulYqh/ROERNkwRJonTOTlXPPht
yAj1Aje2WSCqO197/ITdozbeR4sg1MrQ1T/9tMX5Tro3IiH8F270P/pgMAu+g1U4
GLBVUIzZihU9fO2dK4gGzriTKF3DKtKx3NXzXCsrs4sjhL+ZivyL5V90RO6JHs7y
d8m9EpsxVp0QWS6Ioi/gqw4C5kZH48a5QEMvDbCxDa/HzVRs3DApkQ3vn5+KJ5iX
ZTYKFNXwxLquOkqwRv2kgrpuVz4ytkc/vmj5+shZ10SWciHCxKMey/TS7oKL1rHb
E0WQrj/OHyKbS4cqe4pRza1Y1mzD2XCvT/m1abLFXhLa2IT/1gCK4cYntwLXaHCn
hcLUhE/dIqkATUhgWcJzEAYVmxV+NMdABiHGBqfAMWOIBdGAYTw+/0toT25wLAaW
FQUQkjoHb1JEoRSMfneEAoerS4bZKwEdCkroQUHJgcTLq2RtNcVcEjoFXYYYFPLa
Bm56mDhIJzaVkdV1tAXmD16iToL66MsYHtb/zE76cUnhfPRpDftkaaXQpMmgyVDF
sJNUrx9Z6btqninJdc7p1ssB4zZZiEr2FPJj32KLt18YVEqmkY9TLy59pkJfHU19
bpOnnM90mMK/8xbfKHdWbVkyTFfbydqd4Epdlq+2/YjsaJyvcZN0FqPZP3Fcqu8x
Wk5ZNhBDRlgen1pv/TrGJGhvgLMxUu9jZg1g/x576pJB0z4IFnHKYsJ5h+fvpwoo
XR/Pr4m3FvrlBdQmSQJ4Vslr8lzu7LCMX+H21skP82eOqRCPiUelfDTAcWS/2pKF
TAqq4L3Z6vNOhzxX7LA/xoJEJ/7mPgP06VCptpxsF2S+yHoAlTcatfIJsIoc9bMv
S0RUgVwd3s51UuIj9uUrhg==
`protect END_PROTECTED
