`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x1XvGN1F2WPevs9EWx3DdZCF5UhUf8pEHDoStPiU4sEL1R+F5zIxhLTW+EjKqokO
i/E90LNYXlUWyqRKg/mMp9MIKnQXuiF2CkOc2z00AKqGJJQaSNQRgCs33WszWP4F
UfGeU2haHXuqRcor1LewTbkKaSmSRWG1vphIICPIxbMEt7NvAhwyAnE4wCts+PjX
Tmsyo2k2V/CAI/mPrNrCVgC3BrYhnfy7As+coV60bijXNs4KUms1J7NmQ+JuIcUj
7TwpCNq1pzVdG3EGBPkTMz0zwLoCLwyS793+2b+TNV5fGctFw/nMVKZ8gN3n92IX
0KIQYX7zPv4iGD2ziizvduRG7XIsDKb9D0WWo3BtX1kHHoBLR8geYBN5lreIdxrf
1WaU7igvc1WPXc6pIU+/gCM7mpt/SL9zomOEEG73OKJvVPdtexLJGbBEWOhXevff
xLn+gnOu7zHNICLyCRfXyb9K/1lbsDB1+d/VvV28VXJ370c15dfxq/gy7AmATRoA
0Iawf1yKXjIH4FAMSvJm4oFSy30HsbzrH8bWFvjwdBAadd+yHmbRDQ+SH3CQIbvG
/p7cGERlIOSDk9yKF3HeeNYMUhxNNlf1BTpEa1Fk4Srz8JNvXY+pOEdyEADpHaVC
UGmWIJrbakqAKrmsubdfqPAXlriCNqHP2rE0fGx+B+VA9+yZmJg5ohsWMcDLl2pF
844m5igHXXznNdrIMbbUvonFreu/nDHiGmMtukRTOUDoaeLf7OhhfCsdo6sHzZyG
ZCtXbYKqGisocLStdGqJKqB1fl7QjOG0KM+gTtJ82qfgSgbB19ReM8bkPEjVtiIM
1R9MYrdwtXUY/s74YlKQP3rqCizhTmLOs2OE/57KFiMhKIA9ulAqe+xqokA9HQa/
05f08nd9uQWrm6nkddv6Uv/jpnVPmmYVNSDFRRBnaLL06RnDXeTb6lrNvdSqGA56
a9FKPMbhxEfZD/15uqsF9g6yzNtR7GKRjtKHKuI8UbR6L1pEf4BF8ah/tcqKrgzZ
WcDlJIZJs1+vqVOa2/hZcZc3xOna58HAcfI+Yn+ELTQcv4EwSnZ0/gG5wFwPdZyh
iflCECNlCom/CFCNdx++1W0gp4XTqCHIFORfrFW5ypkZvGfnLrt242+Wt497G2Js
pz2XeqYkVF1OyK75OmOzyII7mKpFPbGaspPNPBEqDTPJpeDNTJ9kFG6HwzOg4G2E
kqwarK4Q3+4jQp2c5WagtXIKePXkuPGIqeoQ+lsl+un1XedueO7qPpEXgew6/Ztg
g1FWFT5TvsHGsSgw4yrT59JD/cc/jNCKIE8NF0IEF1LXGJg/gCPcwW8TcGWsA57B
MEg+0C/bOE8Nbb6ZQ6bp/xAEkOVo5l+b6MdUzSsOs0ugTXxe/vZHRGLxbDGcES+r
2wgnZSodXwJ9vVQZSNAUGDNob0A9VdEYvxP0weoEMs8qJjFOIZ47RsBogIfcIDpY
/0Nf61ATRfvKJlsiz7LwtniR8nXoFaAGrwSApPBCI3i3i61cfAfUT1JKJUfdK81A
y0WrdqMRH88DQXsHkJn6B8tQorBy23qVPdAp+X6r6P6WZKq4zjlFh+4ppHsnJtfP
p6vB245erEgKRyghEFKfgqn/ptO4mpuuoVTsPqoiDW4oE5Cv1zEPjeIi5lcc5riY
mg3stgnh49l17Iiy2hYqGu5H8STNGojtRvdYkBpP2TFuDZPBfZIZeUjxoZr+iPzH
aVuPp4QIo8A/qdQIRRot7/Z3SYXuYy1vtF2OS/ZuGQWnIwgCmOY2G4A/UiASvFen
JxoDj/+N7Er/kvavH6q+J55ZuA9tpo8Ji6R4vjn7GQi/dCsFU0llQfqpqVfPN6gK
tj7TknTYOLavKockS7AyZA3qHFUpMTqi9gN5iLmbaYXa1ObgF5lgSr1rfPWImFpS
UTB3MfNx20NnXe8FPdeIpfT1fUTO/FpAno1UsA+m7E0he37bXMaU0y6CrjSVUb22
FGTAYckSWJKZpK+5e56dBFE6qEftC503+c9wrrVmCq1nszuv2wtq48r5vJrP422u
P6JU9/eQN5mvKWJPWjDU7UMwXJQMgydg6tnJhnxDI2GSCqzfioMugy2t/ASwdAVQ
YkVgggEzO/cM7v15VGAkxrwDJHcXblRSM7N/xVHtlj/TIs6ywPfEWWXpuJShCSYX
+4oHsc7067pke+29rBKvKYjLC1di3AAocqrD1V6OmbVJS+8EE1TMDoUeOH4XuM/q
ja4Iew0dqHRmwJTE4iNWsyH4Wfu4+olbhwXLI60DRxcGBk/lMA+uVFYoWAlW5ysD
Ds1lAoob5PNuhCqaf+0MZREu2awMVA9UzNP4ua/620F0HoPGcUeUq/O0ssKka52r
raa/iK7HsKJpqCLfZSQ5cwSzocIozfW01Nz2zV8JMzbe2y/JshLMnvJgy+riX8fe
Ymw01sP/yWJi/kDlGhKReIUpd/qz02qpEv1Ye4HWXF4doeAe1/VsLU+lSOHXJN5w
B0j7Klpf9l/raxT9utAP2VP6gQLDKbOQS6CLogqgYlXm5ue82Kuw3MV4eY0W18j5
nsXvbwPAGdApCXEd6bQF7uJnr4N5g2wGyVOdgc8Di/T5EaDgB1/Aty5X8hWaBKn3
SbR+dw5xezOYt0Onu/COzmQMPa34q1xe33VARqz0QRSyr+se9z0rktE4oFKiSF0k
4iAns31rDrGQF//Jx2Pbqdd6FFkqVm5ObMB7GBcQ3rWQ7MHP9EXorejVUX0bQ1D2
+WuXhTMOZnMxWumTMo5M8hcaiQJwLoXioLv1G+TjvFPwKa67yDs5vsrRA2oNUHQe
N9KKzoEwVAhEtrXo/L4/u/EFEMt892ZiICj0flym7RHgVsMGzi7uu606KRCR4BW5
/ZKchH/hTKjkZ2imfv3Ark0RPWAQHjJddC3HRf8IU+0xstWoggAk2qcy1K4QH8bj
VanC9fOKoeZX9qBatGwEY2dQZ6YWuuGGwNWGGtZkH4KTc0AJYT7e4+NtdSl5HPgr
hkiH781+bnUjg7N+fCBzUDQgP/wTWaIKvlc4GnGed0kAUOY7H87R8Q8VQ1U+dsjY
CfATkrBSZNtxxaqKRBBS/Q==
`protect END_PROTECTED
