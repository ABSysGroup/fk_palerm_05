`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6bd0cjW7MYDCcfeo/OT3zX2d9OT/0VGBUsF0XdFZKL5GhBnaMUKP1a3xucebn5nl
reesRwyDknpg6l5nsAVje8pgUbJtWdWxLDdot9rIuWvJoloOgIaIkIHfXJLKxZzi
havY+6LWn+bltJFNDgwIYpLja9/KZ1nMM2ASRuH+QrnCVrDgLf+sSClcB6yGCtW+
4BjcNE+uMGA9oquItu1PyzSfMxLsB+2garOb6Wlonk//QYduNRGRROOpo7feTQOf
B3UJKE9B+H5KjbpUIWhaXoQAP8YxykZ9maT7Sx3q6kZih5OMT1k3C5x6QY4+yphh
g7pjlJvl/7NOQfwz2z3ddBsU6sagGq4fDSDFfGfeiUz4pAn+BRHl2Hs9Yh+A2R62
Z3WVyCgQyxEBuQER5mPc/2RMmq1AbWJ1aZwlSLwLPcabgvAgdxWB3AmYrN02PhxD
csd18Ei1wCmqSwOVRDaZn814zGibmCi6vWPQKZ8yK5nWyk/Uu9DRB8CuvQLI58/d
jTLMKDVCRwQlnhRNfaABA5cBjoXb7xExTCJh80bGEvRZ0hloDMN1GKQawdn2E70v
pGDQL63EA/Tb64Q9LpLTUrESrJVA+lnLfTkS0ezQnOBcFCtS0Y5ka84qNK+FvI/P
a/nS/3oIeFAy8b/FlpFV4yYgQV0G6Y0OJIJVT/ZN/dHuvLeCfpk5YE6jqbFMkrYg
EzN2ezDmlZFHEH9+Ele6GUdsqw2U0OEYLqm7795P5cT1nSt/+47Bw5ruEWn+4mmE
Yqs2sNITJwNrvOMj1i1HEipkfnycJWa6jy450MFGZp+OTZvz+fKKd/Hne0/eqU/8
HDZJDU9DpNefWz/3+7bTlLLgLI3sWDpH6jt8FHc6Y5Y=
`protect END_PROTECTED
