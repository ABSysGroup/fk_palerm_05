`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lPp1e2BBlIC9XXkAshMscHMEE7mxJjGh2EqYBO23/pYefSZB+imskc49IatXSV3a
Ct/ksdlgIfwvLtBogl/SGK5BUfLCriXyh3s44EW5ttPWe+85l0Htv+igXXR+WHiS
1TybKDPBKDHyw+n1vYFrXziKRClLdGZUWNlB/oc25TwBw8yrIIaQ2P2ASOG1FUfP
oZqbWpm9b2+Vo67VFMrrEy7mFIzi32u0h077Le8XI9pddGSr4zH2zaTTgm/P2e1e
J8AqhsPtSwaTfA6xf/wUztxno9pnxxDDljP6SsXceLf10sFKB7xTTGLb3F+Envkp
13vB9rqkLoQscvfqrCMn5D0t8gFylPyofJFI4t6g14lk8fllNyi/cEovsqUDLdz8
3JKJiQuN3PH++HJJOS/vxDSwjXh+a9XHTAjUTukr+A9/FDnB4A03nSweYnIWV3PM
`protect END_PROTECTED
