`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lx56F0j30Sa5pLiA6BwMMF3HbXIzEW15o+DswxwDAHwKIyDeKvaaSrbIiE/HfB4l
hQvtW6E4pgUOAu752+4iUqAsEqmyiezhP+vOvi8W/bWuZmp+d8qwwrWXXn6O0YUm
sG4R4ZpAohjo9/VXt8m/X3bcbsr7EnymR+CJKC/rEUYJwZufgBgYokkq1OlA5s1c
tFww7HqOgkUJDK+hqdA8XYm1Ck9VLWdMUURyNFzJJv70JeySQNNoUgEf4r1wRNOk
lBJ8uM2nC2NC58r8TtxHhbVqf43GWziCYLA7TA5qhJfggYg5gOBHDguFLVc1n2gJ
27+zlQJHd6pKs52e8DxcuVj5kQW/OehqQCGhI8S8uGMemhUAfKBU+O+ebzi12eRb
nJYWgyOmWnOYTfpjHihzP0a+qeP/ss5mFTi24RVRcKbegUHSn02yFaX1/IvrLYZn
1er8JN7aBDYf4Qt8IC0ptFdxhGeERRZu9UEEzSQ6sammqhehjeEqIqPdnU8cxD1D
7q5jElvrO48tsxSo3rlnRiBRXma9/ehU++23Xqi4zMHp7R/RysU155/y0UyFzZD7
nb7KaoUYveaewYfIYxS+mml5NBHkgb4tHJwezKi8tj4hx+UOHOOkGx3wonpa2EFN
OiPLB9x4BMVnJLUHioVN38HHs7NE45LVC11BkO14L/RMlEXVwtxFXKxStTaWuiNA
wyjzTorIrBAy2t5u0q5BKtXWOR86lOMeNNt2GjGRvhL9Kxead7i8hY/9e4UQKp3B
4cTNLQhERllIVSupZw5hxZueqXAo8b6/M2W/kthSG6bcNjm/nMjyBJXyNGOZLsfN
tyvWLALduyqERZy65OUfV+/cqflh0BFm8yBH+++NyCgmxL/axVlGj4piQaHiaHlB
lExu2WRRvfmCA+2EdTNBsLkHNcU9fIc+w6WwXmZf/iF4FgdPW01lr1XceeaSxZyQ
`protect END_PROTECTED
