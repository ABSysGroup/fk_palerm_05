`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
csornZGdyzRFsI0XsYkbZIhokxWWZ0hmPPM0HFLD3TSKXipbqct3ZI4k/dRwvfBV
FIIH+Kal3W7Xj7DQnI0a4DEgSsleMrrzb2hXpry8ndmFdJJzMT2fpO1H6Y3JHESw
MvixQMXdlTYZF61HqZ9amhgu5aVwoTYrFtPYudiD5/jq3eApNiTAsbZvpZpMt0Ta
MbcNMKRWyKGX4G5/xZDK7r4RiRCRs5sSKil78T3GB33RhCsYK3i0Odf37+BSfV3s
hupYCk110KylkfGfSpJp4bJ/FZe2+B9JHwzTT4F9OKc1fPh7ef/YxXNKhOO6TS4y
xswq1EdKhYyasGJEBFoPH0X2HbUP6IE7gxPrfMDADcUvpdgLf20WzSEpwLBQdnJu
j4QbSGmar9j5mx8QpZuAl4HgaJzZuyJxjhd/HUtihr0pmBb8J03+CmuICRNihmko
AaPBgEQJzgHoMTomRMjVTm5B9KPGRTvTjoTDstKqrQjbGedjk0h5y5PEdvCpsew9
g/UEsd9MocJ9geSA54hocuFEx37JH5RSs8VeBWck3mqz01IGDTD28ASOZYX0dX3M
6YMlRffZECZs00RrcSX/+Xhv1qPnqFA2iyj2C3TeDq6DCrX9xHBC6NXALaUpcGdZ
VrZ/lM8ZpdRgZjnhqlPxGaaQtUqDf4c/wwJTvq4WUexD514zp9JP93BnGGnVeYGz
NqhbU6seYdoHCnx+BmQHNydztg2uEHsKTvbg6K2s6bjCE6PMwllgJ30X1Ujw/RuR
E6jdk2UYUMvTDpOCtmGig85PKBsoLenZ9QArulx3EoJX05fMlhRhQQWnsFT82pNX
pjOGjc8O+gfZD9jfgU6+nC9Xit3xClhfyepevrS77Zll3Hlgb3B81Zoh2w82RNHE
b3NlfBFO2tnE91LIXkyo3EafjXbSxxlrKxnp/v0DSZTIWIdShNpHoEwSF8ABqbY2
`protect END_PROTECTED
