`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kAglpnX/ZxKHg5Ut+IfSLcnR1He3hadVtPEkw09VoHIAAOPs8vw0C25eDQgQ23mD
6Sn0776kg2CQOtyxFGQTJ8koTtvfMIxQS0yZSXec9P5nR1ZiH4Id8m2rbIgexbAv
NfERn6gz3oossjsoTY2vkDA51skJ5P7G48GHZGIMLhhTeDFaZJ3kNIM36/XQE7g6
s+UeiEOex5QL5T6vRhPqh/SlFk1zEkkdOzcvUoCJ5Q9ptMFgW2dSP73uTjcOKq0p
kNM7wkxDZCQ1oZKQgjJ0QTvf0ftMXxRMBhl3N1C60WkCKgfRFHI48cPY6sWJKHQE
OEzfwBUGz8uzA6vmgbRV3w==
`protect END_PROTECTED
