`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9aRGH8JnSfR1UH2GVMTKEb6E3UbXoubCZvoQ6XplvaecQUcACBwfRQ49wJ7sukea
wA+L4JH4yKRJ66MgUaNhfjaaawtkbCPTVTChnW7eTaYjt32fFRj7AlvMMIAjRqaM
Xbp6dBZQuwnknPvvh5xBrIrlG8LkMQjLlHZ9PGCsdzmGmJnK3tA9QtYghGthiyY3
IBbA098Q5CXy3x15AJR4u8m2FjN0nKD27sDYdqUUq7kBY5cdmOFMRPWYbqMU6uP+
Z4MqfRpIJuhymUCucFNxWTnrkrtiShhj2M/8rmiOS4K0U9j5785Cr123rG0XKlzi
xTHvIlSFxlM/JM81wJHUqQEitvdvWmpLYVbPeOsgLFmj3jJ6ospnGgF3+NgJgKk0
CxuWaPBPOTwu7GmO9BgQct0aEs4LRCzUD0M+8NAXCTi9cVq5QU5I1T8++WNxIneM
cj+B1QkvZLAsNEoj3SUDRY1MI7J4MGoK1Uvcj7iCC0GNWKaulW+NVgDzHWb1G4VQ
5cQOSwJs1iMli+GVdT5VPAlvu21zXS4CT7QcDF4U9royqAVjJsP2FR2fYcIl7dSa
ZKSswydLX0H0dk8qu970nRho7Np63AO3e9/fxwVI68ciPM9NtrwvdlLi39McBC77
Qvn8l7tc6zRR/1z+436v+HCx5+0EXYJ4mvjTybKKa1hJ5KEnZpo/F+06FXyWq+9E
6sWFCwVujlAoMc17xjKKYyxm69BmAN8lslbXbdCGvJRuSnd33+hHw7oDeqJWe2B8
rtbTnUDiLzEULQN1hRcALDjmQZk6O0mE23G9mzMAP6mw4nanybIdiOohWYrkYrtj
i1fYnCRoooOei2qrofJp2ewQxbjfADIXCTQGHdONcXgsrEu9MSsfjmbNweuXpEto
oNqLfwCBBCj8VQCsHLuUShZI36lMpYszoPtmIvVEV7yuUvOXBapF1ab5woUQBU7V
8RrttKZfYhr4w3iccvyIYn4ElTeCjc2zUnBvOFiqqUsZAzgCc2P1CYWaQG95ZEEZ
Cb0nSNicJM32c2DmnrXn/mtGy1M5XrpwbTgbvFEjBSmwxtoh5mgF7VHfpIftxdTV
IG5ffF6v8/1CkgZRjKNLGOjncyQuqs04l71khO4N6GWUwIP0b7dzpF9Ez15iib03
`protect END_PROTECTED
