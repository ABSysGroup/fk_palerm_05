`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kgd7GYGYXkMf64/ptBu/C0DCVOAMRwOtNp+3ASqbAjV+lLDHxEtdaGSUO4B9DR+w
xIwhI0kH9qnwpa83bLrMJHmBzvAJCxAbATK/7VT/nbgb2yonPxenedfDIHbZVmyW
rWdpIu1On9jA70C7ll7yWKtBW2sWAy1g9ykmFgzmjlMqbYe/uLS4GtOpzYvj0r3g
gYRiuUvFs/gt1TWlRZfFinvO62EszRvhNkZD85/s1lael0Zl9KRSyXxScPOwnOpz
6Uw6bEw06EcFbgGYMP2eZCOfTB4SHbVoSPC0MI4SB15si+afzYr86MegGDAnnzjx
x3nShg43m8ASYex7rFGc7P7RvAYZRbTzL/rgfHfftfo30oYSTTExKpMg+ORJmTvA
ABtMtBtO6e5UacxEOPnxpt+EKZUljzsdcDAdBKwsIow/DJ5KKkOUbXKLgSk9Pmfp
Og4plZTADVnR6BH4tGw9c7DTOD4loFNfOYcRdVINaiLWXGYKQMsxKssHY/ALf4iw
CVGYC0CYNLA+eXOzUJ1W8a4WC7rOQWMA6+C3Ji6oX4Tby6fexfcZOxVxIeC2qHac
lp5rI0B4KfuwBRsDZAbzMpCRj3+QEgXeSIrSB58mR+aPuMdTXmcZuP7Gi+jIAkzq
p0RgkJR5GhIdyOXEP1S4G1FELNjRCWabcLfcHJbNNtPTLRdoD2+msbnkzuw1X1P1
NgNyqReCLPaxt6J1asJ32L7ufnks/X+hnFipAA36cxC1vDF6pdx/ygZwn/Zmx+3o
ueEV1nGBAoSUBwdte2rczLG2OlfZhj4CkyRQb8VxorwnF5qmkT7v0Kj5boB4j3Uc
ogqwpdr8MH+Hs48GLlgjZVrysW5jUmndoKPfDBGYXYdXWaTrNR8lZyAuOljuVmGS
apTDdQml0rantVbsDXOCF9uo7Qd6GOP20f+jn9Emnh9V+ivoyCYaYBBonoICbHKp
Jiu9RhJudB5DJCR8BFM5sP3WppemFDfk51hs1j40NOfimQcd0WYikAYdrBmbMmct
AMzJVfcF+Hs+BEyk8Oza22GJw8C7c4SY9tpz/r8x54aGmKwJwGboAUV+CIJ31RAY
ulH2Y8skpk+ukEW7OGgM8fPK4iu7rC9MOb8c3H9BynbkuRh06Lq2DbbsbAavPWkn
f1gAA9iUm0FaHMaMOD07JDFwqlZITx0M0DFbOxrVoEcfXUJwbmn1z5zEQMweq/Lr
9jKi4IBfAFYRFlV9UXALf/SdoNi5M3FMtZkqsiCEPpW4VqBnMlerQG6kTaPtBZNh
hf9WmK5SZA6nzj1TwzyV5RtWfllsoLeeBkXA/7d4YNTtExD5HI1umnlU5jQY9D89
Dj64scleZmZz1Ee+lv3flHCwS6i/sqUWUJT9kWUP+NJEoZYcwt0Oi/+TN0lYB0o1
bgeCbG0AIfQ77OA1H0Ytl1aY475/eYAHIyAwowZbGVlv3hm/256Fpvxt39N6Fjb/
+zlMT+RI1p2p8mGlVJfMPICdIq/6LJVPyexdKCsGreXgsWnjfKcXbA0ynhR0Ac8N
wRfHhqavAo0ihMfBUtfR4xWRp3AFschLkSkKP3F7kFpNIFA1+Sb+vwUWmP9Efgo9
AHDBAbyGiLVxSh1rygHPP9IzVuAHZb4m8otGfa7bg0Lixa7QPIB4kjQSEmk9K/JH
TKRcHFbYVzt5RC9VODWi2EyGFxapCCND+qFdmdmInk2J7OPXGl50HOzgGwIbhwUu
UuB3Co5YYel8q0yRc2Nmq9nWWr+eaNkHgxhdb0XFj0iUeDIXbQcrx4C9pOuH+hvM
v8rQjgrduDmE/7P8HrQLnEHuSgW/m9Rm/GjJG4exRgKliAJSMKF0g6Tcr40jSUQT
kIQg858o7o+5OV0TQUQxlKVMKQ/Ixml8GHRRpsOTe1hpIUzfji8k4XDOETsCiAkM
MTWB6H78i4u6NwZYuOzmtqxiveyxZXu8fEDlG6EK50oMxTNtgRCNevr0h94Fv4H6
OAYhhdJx0awKAdEO92Q0uh++VibA5US8cr1umXH+3Jl36wtQF9wiDEUMNAkkGKPO
LO2V6SUS+7mQRSJB0QW5akj0nd9Z9sV0tGf/d5Rg/kA9w+sUdy29H1vnKClpniEk
8RhOGEsE928qtZGwp0tpZdt6XBZF3UqijvagmMZT2jP6e6wCtAZamIy4a5Tvk86K
ViTPp9qUQI3sWhAbnJnLROgRQyvfjD1Y77DjLxvaca6VPNqu9WKTo2UbgYOUESJw
8nbfs34lTuuPF3xyrW5NgJwvZThoFs0uHmNoDLCWGhgb7S2Aic2f0x9SRbKTJ9Oi
/7cc8jEuf4eUnirY0U7YhwcZWn4riPzYMnrfURLbixDqn0a6smSBDIaHR8za8gAg
yLbBLT2PzkkZRq6omd+wpTwWAxfWqSzqnPuq252XjoJLvkiyjwoxIa1PLjYn+aeV
4h+VV7r8dwjTMHf4TAUj352GQE1hwHEOB8AbulTrPcs3gPyKRum4C4hsVl9KwWJX
rbGJkmK1dAchu1fS9LHYObIeJUG0JMaN/+jD45LIBSaip+hfB+b4tpTVyALashMG
0ThO9qPl6RoF3op8WdQmJDPcpnmHXzs6NKWFFp2j0Ypgyq6BYYyM8H84KrMt9+Sp
1U/IDxFA3urGZwDg/WAgpd822QRtNnTarggqNrvPPPpk7TG9cmMJwx+hZL8LkXBV
BIOYUvsQ5rSQu0/owgQOtyBIjbYfraCmjNdLsgWhC75FMzfxUEAsgGuNEAlDhoDf
JQzbjQ4m4pu5ZJEnGZfDJkR58TWI3esgkfuLK4xXXXZ+ZkvyRtAL07jiYKifiGr1
5V9bI36GCfVTG09Kog8Q/xYCO4GEXLjQ0IQZdCGaqbn+YpteVaY7XEl6PwKqvq5q
L4ByOv1xaecM2+sKAYZ28w3CGWlhHecrWSi3S8z6pO5it51D8OlO4loJPbcpr3DP
cWr6idPak4yNJxDIkjmQvK023uuJ4lJFbevwKQSm/j0AC9mfdvmWpiaXofvUCyF+
wU1RzdvD4jhL/eBSDGOh77P8U6MmT9PbhjuTohotrbtcz+lpLvgJu+7RClU+WHY3
Zfp8KpGOXOGbtc2ZvA67nBBqrTdHpdmgp12mLIfWrgMfA2pThA51xZALS6LH1CGq
P0J8ZHKcdXckhGQMeEOXY1xb2NreereZoH0XD/Z40hdb6lv/pdbYScjZLABxenz4
bzwzmvTIevC6+SMFNzdUI8SpwrqUxAIAQ2djU0B5+irIPS+8GOAmAL3jwcBlWjNU
nZO20kWLlXLLzl6frz4I7RUzmxtYR/0ADcXjEI4L4HnEq1XLTrRbfCYrh/x5vAJt
9QMHL/fVPYNdJem31W1jlBENJeYvPKTYNPlT9aCgRuG89rJsFwAhgayGyYh0b0yW
57ieEGcLbe4k1D+lJ1ziPLgxw6nEN7TdAIywM5P3WsDdxJ9LsGZEw5Ok6c4XuTcW
TlwP7GzdG4+Vc4MUHPvh5QlUvJH/wBfYEZmI8zGYojRTwuxkWXPYRCCXnRu/XEh1
K1VCAWavCfCVgFf5vCrmj5AGdUaMsYFy4e7ZribFZhMM0glcYjeurn3emRTBor6d
TFVkHytTfkVx2uiPMTT0pUcZLS2ojKFm9sYSqsb5xnYF1PVYQ+2CTVUoFoVvvU+C
6OTfQy8fprV0GU9L9Fw6ZKS/SBGrb+QpYEkS+h5CnJ0=
`protect END_PROTECTED
