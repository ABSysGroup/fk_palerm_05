`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
63jJfjCQNIX55xASRG5jTyfNM8Y9vSBAd+3OPPfjL2wtx+zROWV/CpUm7RAO/u3m
FFnJnXAf2l7LqvMUbMeud8NUavPKSHVhC9p+DorFLeW5I5eFhHf8iKOn1WFzBClH
2UQ0QGCIBkywqekUCuHrY9aYNU9UiJej464/Fvudos1chHs/QxXyWsxc/4Lccc50
uthGgvYvNnV7ZA0nyqUL+jHba+U/21xJp7PzQ8mAzSLYjImBDe5Fkhk69pl9IeOG
xL0anBZ6+c0PGEY8RR60fSGKokiWzFmQFmfXx66JJdlnf6qycapRsl3NFuW15zgQ
6nxXLtMPMg3lIaaoRozDfBL/+NBpItoLH3QB/tMzMglWWzwKseRrkwVCTGyJlsFu
apbeFbJ4gBF3ALZF7fPeZXZRByBwvGNFyxwy+xhdFJgJTZSSSYjpyep6r/g9qmXx
G/w8rpAaYS7LshbRHk2UC8pyJwtzGaWPOpxGYp/0Ttkw7eunSLLrR95QeBYy8mcH
sQUdQtMavf5PwaG+rYFIgpPHzj3xAwKuu4MnNeQ1w6uCDhebM4cix1XYsZPvvZWX
8tD7VjTG4ldXQtGZmr7TYZbHQGXHJ7ZrX9UaR80YAbjwphbpQXlbcMnxxCb9EqUh
rrzTqQB7Pequ5Yx8eF41Q6yUccij7b1jqTj5XGqub7bFg5E1OQmaF3p5chYX1U8I
fqB2+ENU1SM75EMYUAfKddzKmYqdbLyFp9LUx58ODe9dZ6hYdjLFGllsENb9xDKP
wK8LTuVbhW4idvCTojQhQXCTQW5YXp4E3JiPFc2FoI0LqQZmGOdf97PdOk2lO2Qk
3DCY3D9RDgCh0Y+qB273cqSR95EbEZ2IYbOr/gpAF13z1J0xlY+xm4hT8kuhW5tp
IvQqbnIUxBrs5n+UxlhT7E8LOJVW4NXgduLi05Ul8zzM6ag1zINgHx7+ivsCuVlj
`protect END_PROTECTED
