`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Noz+vaHCbJq2MQFSDwRepuL3F3eBLqSTkXkO9mEvqGVjU9ph84ED0kKCyVoBFjWz
GNxfl1UgCdTwQfUNGSMAxhjyd+Y/sXhHybHY39DVxbalSPKGN2hc/gLf22dCNTKG
z4UGQlA42JldeDwPjLeKWRIzoP5OHu+PMLZq8DfkdNdwXCaSunvNiFdoeYLYL145
e9KzZua2gf47bErHdkxJrUZgm5Pw6VeuOHFig1zwNuLGM6hUe+YwAp3i7YBud21N
lcaeQOLTihAzPDwVY5yjV7EvBUDUubYitDyaoOfs6jV7ZfY5quHc7umC2uikGKeO
Do4TEYoYC2RZt7u00GVJOcNiBJz8Dsok4TOpOfpBycynFSsz3YfBI7Z3/nv2MeKZ
OMMBZKlG0MCyw4lbaY12RwTr0ll6VDZB5mKcNDAy2UD3nRKFjhWnofwN6BvVPkXP
XQUmYw6aWGaif1mHFiJ06/+HghuSPY9iEb7qdr8hAhEOuMQJsO3ouFWQfxwwILuY
Hmc8WpyeyvvXh0pnEdLxAOrs9vdSt6aAjNQS3xwU/6ACzS7aNK+wQQS9QJpe+Hyo
VQZwXIWeo1f7K4FvEeY4skXjLcpO6g65RHGe0I++qe+OgjI9yv/rgleomqGkWbzl
e7sB9wStJJQtap7qn0rbQw==
`protect END_PROTECTED
