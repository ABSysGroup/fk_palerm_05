`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PpQ+5jJGkEtKVLDMi+n7Bxs46hSw/ct1U4Izr9UY0EUXWSLl+9aYmi+yx4EwUDvH
2oqPbXVjMA4SBp5pLeFR5ceEKzoPamfwr6MZESX5eN/OMvkrr9798XjKWXPYq9pn
HOrqO6SWB9pcwVRxXahmm/DeuIU6mAXja+V5Z4r/YhlNa6yWFCv6x2u/bvPHqxKv
jW6rdv1NRwruZoix2J+IQOGH89x5xPhrarxM4gWG3gjT8M7RoVQvqOnQd5BsHvm4
X4S2LslqVhmb8J06Ds2SDQVQ+UeI9kbUm7hxc8fYmTUmKZ41Sxf+vl6SOVc7t72S
G2y+uRrxw6PWBrU3pEsZZD0etQ1L7mvZcMCuN9hPCgddOkq7CSrJHSQ7SI5Vc2TC
XPx1Gfyw+HEj7LB1d0U3UDFwuRQzpEJs6Y0XtICC60l+fRkI2q8iZ8B5JoInUGi+
ZD9TRK70JlnhpLvXUm1n+tt9vQoZVsVEqXxckUM2HJY=
`protect END_PROTECTED
