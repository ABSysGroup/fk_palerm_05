`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8gIL9FabLAs6QXdf07kfTt78QyQe+rbJJCP5LPLuLhyNH+SC0qqe4sLDLSvGaFHK
eRMEe+Vidvlb4fDsgDuA6kzRqR+Vn5zkgmzfeRMqQVeA1fU5X+VXg7Bemvo0+URM
uuvCtfpuUsKs2tWUVx5l+9/EqserFIkMA9DAq79o9uHBUuAuVQQwOL/wUwrTbs3X
Shiyi4X62JGN6qpjStVVYfM2ASX+1jquojLgyqko5HvIokDKcoYaeouP/65kmpio
0dPztHgOxX7BJrPJMW4iYDpCJ+PfaHCNPFDcTW/OUxAg27h7FgULYw6gyptcMQDl
M/say7o2Z/NFzIa4ct2NhXfi1FeF86zAA0BB0M3BPf9Z2nrTetdo9kZ7gHOF1Yn0
tKSo17z6+BUt29gnRBRgh+wywaHmkCfv+BqJPai+qymue3TCaLVTweFuEX86eS0B
et0vw5HgAGT8W+gyspNVAWeteR1+HoX9Blou1bBa1G+1S5NXhtjwDog/5x/4Ob+w
thTMRyUoN29yfdlq809Bxi5/B64/MeZ18yZ68shzbhKS9/Uo9OlZYiLjArCJCutf
FIghTGF8AjZv7rMU1BMMVUuBDCahAUitnFRnJ27xM6inuG0Trmnzptw/AXjt6il9
OnhIYDMN0k5CkNfLFXIKu+H4Bm0JLleTTJg+ki7iDujrd4cGaXeTjiGb3n0othuP
tVMUVoAPLpjHlGdbAYs1mpU1QKLm+BXqbRUIKKbs8CMMqaQLW5jrj8nVGSv+5Zst
vKjNRal+2FA2+x1NGxz4X6OQqodE+r/Oi0gTDeNGzI3s1OdyMq0T641uGIz+DWl7
yNH4xJn1L86auhdYsMDtLuWmbO+5cp/bzix5b8op8IQpUUkhw6DjKJGVzqdOrAun
6mqadew4DiD8qKYzXkTNziz0Q8fKKtu6KFiBA3zpYCpKR7H2/6E6wvnNigEkiAVg
`protect END_PROTECTED
