`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XaF0N+2aibVYwHztjrs3vTNnWSjQe5sce2lIg0G+KTo1zx6fNXRMwXkPHVG0Uf44
UNc1I0keNKTQy1UaMmXoQRx3gw418lPtWhOB8KNDh33XeIjo4T76iEzjuDRcj8K9
UeRgCTFLom1wQJqYLHued8EVKeUf3NQhuuNxrxdBWBVHBgjyHD4a9c1+dz2SbR2w
6tqPsMcZgVb4ORNNBD7qggQQA+EH6NV0UUiCNJxWUW5SxfxoqptFrgePWv+jaC/N
YjYa1FrAzCTv6nSwaYvaK+XPz25BWYvjrG1f1CTDBmwqeUrvtQQWLiZx9pPkdzJ4
moOC4BfOImqI9x8JFW+JCfvuOf/pTb5qsfaSmuDT2B4BAXQpLqTgGvr0idJ2NoZm
wDuLqLojjQocENf8XEvfHQnTHx3XVcLqFqKEnnPqFQcfHHzNI58xSa8j+HMgvsNK
80RbR+/ihibQhEMdUmKtWrJhlmTKjztAjflqZ3AZHJm6QKbc1Zqt27DZhNNl/Hop
DPWTgNWRrsQJ3nafiP9tmOvBMx61CWsmiPTfLQ7lz0ZC+iALE2DUGexzyuKHHMPn
`protect END_PROTECTED
