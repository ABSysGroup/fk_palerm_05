`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8hO87Fs6YconyQFzY4A4h1RGh7By7XcUreOBpdLmvDe5057uveK8l34DBN0V+KXp
AdXIsc1wDvDpsPh8kK79MgzuRO7+Q3gnoO9WrYBm1pZBVJZRM5L+tMA8/q51RzY3
6arXZRc0rJvX+uiIq9+obfKAJnU0dWCQNNfoEd38mjpXC7zJh0ghQKtKR5Qqq2gB
g7YvCSqRmvjJPuzA1F52HYhjBz4VKaLW0Yf6cpFxoPff4twPFB0jARK4zFG4NIhc
l/Xz1DusolypPboxEhBS9Lxv/OWuJGKe+KAv5rQNSnGzicNPP8d2oTl0CLpstRQ+
gCYGeyKABbSjmgbMUDqqPIGOyeN5w361oc+oQrtRFrmOwHeC041VqeBKRL9pPmG+
olB4SwkiDMDDSOTI8v01MFGmBCSJ97NbJTjFaJ3Z9ijurx3+9zkpuLVIEqzMfvWk
2eLWrBFMyBvMgo+JokULeUcpZNQhC9PilASeL9+Ee/0UDgHV1UvGnfJB8KGSU3g2
y8URkSmEVg2Zxam8KZoklqBzy7vE2AMrX4yUAkUag3xY4E6qoddTZ1O39RYVZ9oL
7WIdi9azZluUZH8w4ottb06PeXFLzgKWQVAtiFo3EIjRRrqQjclncvFLkT0Dq8R+
JKdfUhnlH/cMupmRrEnMwMKED1aPydc2gfER2bCtMRClp85c1SrGHi2h2MJUQr8a
Ya+4nZMLV9QBVxNZpHzp8CGvWLh+C34kUhT3G/tLNgfgCp+N857jDBpg28i0yYR9
WnHOupY65rB+TvrQ3RmTZMRc9qg47rPSAQj75mG6GuAEtcZtKi4jHsJcGy7eZvgH
v2fp7qK+NKh0eOXIcKNXjJ4vfvbjSFp6d0IV/KCqt4RbG373t3FuutziXjTeMplD
vY67F9Yj2I20jb0uVe7BT5TzaqSNg67KNTnCNoYLxUiVIkFp0QoQ2zhQ+5yiSXXf
lrgCvR74tboCEmpMxx1ZL5eU5aAyhhJLPaFGqLmdhhIid3OIQBRaH4FInAGpWLLR
N1reonSN6ZxSEEmwUwxqBtdBR1zFQJ0GOo3XHhVCCKpLBHNMJXmXbfE574G/aTDU
dcUjz2ynzjQ+DefPuxxtDbD6SC1EjY1imGx/MyDNtGdYjI8HPu3SdgghKxA5bM31
JC87LE0pToBVoqCyLB1l8j0nMM/aof2J7tbU7zjKqLvgnFhKuJ5wtcsURNR3zIiU
M9usyNt+TRSqGWwld/qGOL1DueP7S7WYWBDbKlAtc4oCSZ3CJnsSIPl1Lr+PaFQR
bggK37bWtMT3lfxmDslrqJdAmwandAKRJ2wc+8S9M/DdKcnQVhfexLQbvj6hi2Nd
iCfz3tgLX035qAX2hzC4jGtxCr1Mpsk7OOqo3Zw93N6idIJWrhSXQz/U+8Sh28qh
GBmDiou2L/dbr82UlsYGCgzS9hqsNFiTe8VClpGTA4rjdbQnTOOBVfB827KOD0LB
adwOvH+TGRwzid5wLE19xJiU6Ida6+VGBLfUCqlCcm4VVP3VCIxCmTnknltI8BKJ
cwsIVCsc0dSTqVcp4a0X2juETMxvmYtzINbRi/EOTrRlVa0VCHMB/zivT/WGLmVQ
DZKWsHg9dvO8MtP5W/dA7G6SkpVmpx/wQez2ArYUJH9iHK+9F6fU+PDc0aC65ZaE
trfkPUSpCs4so/TdXeJOBOVf+HFDwX0LjXIfo4FI0hGdiqWDVOl1OPONZB94pJx3
+6FiPXXBMhuzF1hS9NmXlVpdWwoQGPu7z0KY21VvFGELhTw3g6/L53uUgZj98rGX
kw6RZJrX9vD+4Ut6+pk7psDluZvBRg7VN55ze4P8NCTmdua4efPem5HE9/BAviRC
bQsILiBevSPUunzibsHBKnk0Or5JBy2Mr/AP9xFFvK/JLhjyM1GSIUsTo2nfDoXu
wgmKo07l3r957z9prLT0QIYvjpk/gG1EeE7Sy1waHmRUCdcHFrWhKBf0rnE1vOcD
8FBCMYfeAM4eR0biLWL8Fc47VxAFwf9OEtWg83KO/ZbtmcSvjAVwNs+H3AYOsgez
2Pp5rWJEB/MiPSL1ix5fup65tPz9bODZY2CIHFNr266m/8nfk3KFhVjnxMqrmU8f
aqqHAUGE8ivRxZDJNOnvYYP/oFr21yzlFZpfsMVTYZsYWd0ePm5+kXQYPCdoKyaV
7Ouh1a0Hc7yBaNir78MQiTBi8ZOypDXJ5pJFxEqn7sL3Bk8eoepdj3sbYwk6aD8u
NKjePKs30as7M8/DtOPxNsAIht9TMDe2XhHdbmcTZ9iBH73lijRIuo6fp25u1nWD
CV1CIyhfCXOz9zIhZL92VVOa8dVRQGpGKI31LzLqc8REqMVJvQ4sElNfo8BGAXAO
kB0ZETX5wWb2Y64LVxaBC3y9W9BbgR1k4K76DFSBChjaOEIfL6OQvJRKgJCHKYdp
N2vmoFleJ34Pk8oRTe1d7aTVJLNEea4YVE98rPvpCvZAzGCttvlAp/GZPw2MUFuV
uDprpML7wYukbfVbHPVqRv2iOm4fcQsd1Nu6JgDq9dgKdAGutGJez6r+xs5FqLZR
MHWQi1Z9kY3OePzKPhKX8Irfg4oM8ozFoH1iuoBWuK5aaMhLvZWsoLIPDlv7YTCm
d7tjuyhovB1nqQRLagq1QmDcGgZhKw/Z+76o/I7J5bvwZJFXTz9qG7mYihzrQOi4
yWhaJOdVlabiWO7dXy/2lDjAjkdYJKzfLS+jCbbUUTesWhpc48PCN8MCD0ML4rGM
UPlD0nT60AvY0acvFWfwCRwDSUT8ApR8fxleUcbf8ZriGD6R0CpThmAbOjwW4CEN
Gp/V9IZ4SFr9HQDSt6vFi0YzGTLDOimSr/R5rIKfxrMwO5SwV/GhBhTmlXJT7cdf
rz3b6eG7i0dYw7vjDuveGSZORdUMPxvF75mc97tWSF+/bnKlZpsxFPmcJFaznB50
SL8w/QKxVcH0wm/4iDayxrgb6WyMuf2XcXtEFwLimTv+XzamYuyFEY0Z2zCDpBtu
FEQKQBoI4rvLpU/GxSYJ4nCcNwgxm5f74dq7eicWvWGBa4u1HFQcfnpYSk/emGUv
YHcUvC4HjnL5LVhxUeW6mnl5SdnAzX5C9CQl7Pp3O685vgpyvy/0UNgdSj6Rmr/q
nu7SB5hpHfEHNv8Do0zYppVQB2b1NoQhbcppIl1NwTGyzMJbDsfAlfsEZjaGW54m
4Ju/Fw1P8fOeVjF9nScc/i4XD0SqmEHOYQ2zWOJTfU9xquSMT+YhtFwMuSUqIMok
Ce9k1S0CjTuk+0f7T9PYYzzRkdfA2V9O+Ow92APlHKPXkhg3XmxHuhP89ceHb/qa
tvPPmJiYRP3IHSlDXlr9KG6y+OHa3qZogGYd/4CXzhhn32rYTbGcWdWSRcqy6JOC
6UfnVIDmlqHn1dXAZx1PjPrjq8Z4ipqKhyhJzsCemmqgbB2Ho7k7ytVl846usj1g
NFKjDdchWMeIq3ILqmvHdlI0ldlfNsbhXbffeOc7TmFyZctJCSPpImhUwlrV8Ffs
GCxinmqrZuMW22/zfLeC2GuuY5Sb9JfuH2GPg+U3VEsEwqnF0IedSVKpG72vm3gI
CBvcLaXy+pL9XOItoQeWJx6uxfy8QhCpj+Eb/ZvUf9a/h4ergkUpHTuFQZioWKL7
oWEcJJtqG+FY79+4Hsl2uwyE5rDUnNievS0DvCOGAVo2Dxdcfw61fR/SS84sW9Ei
zm+E/vj5uZEUnW+lC/13715EqBU5heoYQgBlT+KSuPgzvqQXJjY9ijrN97MNPJUr
UNDzBe7fsWLKBtVzemDQ/34QNu9rTpAo7far8DJM8wC3xxetjzTT92yzUkiC1TOG
Vocu0bDiSA9EKM5PUXCavPrpBM5EwIyDkL+sCfuKRPmrRnMKCisEpHnFBApUVbuB
AZT/RWMnNOqdkiOOv+crlN5MKREYMMei5sE9V2AWWntI+vy3F7DsVXHPBNnE+aIL
xVbFDyDAMDxeaZ5GUk4m2KZ7LDAFTUOJWyEDQLYn3LiKYfsnqbBHyhqPA6nv5az4
LDtrYV5Z/hDs0wvoPihzYeFmzIlzGQFzxGfRJMtIqy3Ldgz6u89dMOGMteHikbwW
d1hHJQ+OqIp3qtqCRxo8YFw8PabXheYYcpSVfqmgkc2l2FdH4xiIo/GyHsTmTp0Z
qM4LHuY5IAEAvifqHg3ViYN9chzQImYGr6qvyt9nEqS443HspuiDWoVQiu2HdgOg
z/BkQqXBtdwhxLRNIbnTVdrfxzmm9UJvww0tb036UvP9TqRgnwOtloHZ1aKz5Xt5
wQqIV6TRoUhHn1X2BOD3oIDEZb/rsQNIrNdVeekeXAqN/rymD60/P73awZX7zoSb
Ha56DCA7QAfm/5rUhOxnhTqVy6vXDn5l743954/7wPeS7xqYORZiZtShxhSBBHC0
kp2FhPmyTlcMX6BxGoRX8/TxCyph2OFO1S5d+T3thpdcmEqjGy1F9D9E+K0uVVDU
oIPM9kISX+vAnAt/GuoglT3X8m+YkSY8oGZJwNM7jrJGL4rQOPyKkKcJjrW2tkkc
OrUsz9TlB+IO6ryS5JotRZ2El8CiaD8aNFojBfdz6ieDTPp5Rogjgj05z61p0JZN
k3bNHH1WD2ntz88O5HkJ9XaaEPC0p4aAl+d3hzBCeWTdKFeYmdvVPo1ktMkrYxeE
rB2mMu6SHuV6RpUhxGSCrmjkj2OnZuj5X9G1+VXz6rAmZwV2gCJM/joqLkyW29eY
VXFhEeRSkJ3dAPZ1xIiiF5OZJ5kfoBCJWHj+P589mh9n2V6/Dtfj0hoCvffb12dz
p5zHEI0tueFqEUe0MKaXheee0nuNCsAq6GvEWuR8o2q9T65pG8HntQTfgzImvGDm
sH2rP0dIDebpOOFBD3zodiTAu9LqBHwuj1YCIRITlRd+cHeb8K55tVLwe5Lf7Hkq
//rTFPbSZ3CKjFzznYHHelpoMDvIul38rKMz0y3FEH8iO2Uyfb02sB4s+0D754BI
+ugGutjqqIaKASZyVyTmH0vsKM2pr+KiWJfJ7mrThJuYA4Qa8TPabAflooE0b71L
E3vf2fiTa7aKZzTqH4bQZn8jOopu5Nk59QNVJBaWg4G4BeL5KeIceMuIGlP14DnZ
BGiFYsiI9sRTwULr47JPkXbSAe96YzMUTtlfMU81N4AMiADbvKG65G06qlul6yqk
4XzBpthwr2dnNhdMpQBQ8egVDb+LPJ1ggBqOfF7y6i1HsxdRDJ6jA5mtNUA8kE9g
mTWqJXOJVOJAbOR2gRXYQeHcxXm1HCGaTXVHByOYNeywTY4eGYgcks1gGL8JJKOb
3L0KMw9Ucj56Wfp/nLUnRIo33jjy1Nt2Nji07A9/F1JCz0xT7haPrRFX19uNLuTp
93IgeJCyG9n0J7d6H769U0+UgQ64rhRK4NPBcVKwBubGOjMyx6UDEjJ76L20sZ/9
hYt/1vS1Hnq9fxGhCh40oMknFFQGkuu0h0S3tJiM9yBJSTcWsoGiTUpEZ5EkyKrY
lGq2YET4LBwyfhXKhJcX+QeOXIuOuBa+uuc5hf29UEI8wTN18y2K3lW3KjdDX0mz
7wbFCBVqZINZWeFL1Fg7AsUwfg1dHav4f9LYB8uTVb2BEQwkaddB0xddyKHZwa79
FSUWEjTtkHHJZvPyv/A3gRQU+GuuGHLBEF4mkQiOExPIrHFc0I5bU/RGJx5DhjC4
H5+7YDV4VyNzNdEwhBJrVQnKVyNQtOKwompY+ENJ7uVhBab9oZLTzDm31ceFuhlK
k1s5OmVVayi62SihmZfvaBxuKOhDC3sURc9jwPLszR0ZeU5d0EZpPmz68x69ORPh
RnDa8cbBItcU8av8UBO/DjZ69u6Wt6Z8ttm6SGZUuq0WprbUl+manK4WKIxHQk3m
ysHbV0zIlUwchlAv3YecYvnhgHK+ZiOVUWezGi+LqqTAhYFtpLP1NahGqHqeXngO
Zlz7mMJQ1X57lzlHulhkhARm0JVZoXxU1yOx9yjdpL6zsQAZcPjKeaanvNw2ROd3
JmvragsU3iLCM9aSOlWfP2nZ+cEWawDii+RLYQeuXwmnndpG03bx65Jep49tKZ7O
nCHjkg5h47rBusaTZqAwz3VI8/AFQjRF4+fwGg4PR2SP+/1evaSGe+TEK1+v/uJd
5cC+s6rMlx6jzn6jzs1sNB32wciIv7tk0Ry7RjDeLREkCzzQLixUpqtn05AMP4XS
B31p1lOQx7gCMxv9QAFyyPhMaPzVDQl1jXiOTQM43TyEXdMehwh950fs5iphPyJd
Glvl6tDnN/Kd47QcdGeAKmDqicsiEXqCewDnRWoAR6OTey+Nb7pxKvAnUxz+nGho
JI3sYuH+ThN18Wm6jNNX/2qTkMALqnDVk2CGn9I/C9fiDLQ9j0QK3PWN4a/2kWVN
daLaHUHuIpHbH7aipI4KmR+UA1/sQdB6DBd7lpnnaHMAtF85FxlNndajftdkYHhK
DQbhxDFrZVdeNqhktDDpC9ycM0c6Aqb4StEZKCFW1wsgXaUoSlgbzyEae7Ge9uEG
qnKTdyNDkeca8koFNJQHYcFvn/rc09dEngWWkhb0JCICCKFJ8SCX+VOqC5EL3R7P
zf81HSMOQkzd9SndkLvcdTXRcZwgHR9krpSzUmOnasc79gq0TU5EfuDbX4XBTRP6
VEENxeNGeBn1G+3geZso99iR1YyyWqoNew5gQXl25udrM/aWwMrwYpaGlP0FFzF1
PzIIaVDhbUsREIMiro2MdXtqY2MbcYFcU/R9utCmrNotMwd3bi1ws+IfwoXUk6Zy
01hosr9vH78zJTTEbt7N710DgWShuV1CF8WiFWGTGpakEasxOnkAyF0eU0NT6CWn
XHSnG8qRWJu5H9qazTzEZ+pqcHiIqSjULc5ZXn/QkEdJtbxljh3+o2gLQIYsZPzC
y7LxK6J74sR/N24ulnuHFS1rrY92818mA5qOxL5vY6xUdiWV3/LjdWf11hzdsjaT
aajGdFQc5Q3Y2QzOu3366wTAYxDpXRLVJobNFtaUEjtNDzWyfii+Va62K2CZyR+6
ClUHJ+dCxbOiqeXw4kT00hWzQfpetgsIAKFu3PAHlbXV3oHYsZuz+UtzSV/szsi5
LEucq5llsxeUnwSOLQWNjn1FYXW/blX/HhenFmlkHgZ51i4bA1lOkWX7yyoJ3QbA
PlP5M4NehNkWHQI2YNt+Yy9bt8LyLAPo2G+Sd0oJ2B2qYbiOmOF8cS2YW0Iw4UCX
xzJsBlIwUe2fcqJS0vRW7nosfBTjCEf4Rgd/YrGUFJGtPuZ8vIFyUKiemW3dUL6m
Zf2pHmLtufNDOhyxPxuTAgRE6h+yaCOgCpk9oL/3tgqaYlZ29WuR9+kBIN/f7JsU
7ODAI+wT6ShH6psmgOTNZBze45FJuPdORohWrBI3K9kxnVBHAEreWAHuuDOoKI74
EQgRl0vw/RM5086uBohNJ8yh87byxwyse/2mZ4rTx1+KbNAm+P6CJckxyHZ29PSP
VxK4jnhNIhiTgQ6jXXRg1+LpRGopXgA8ebHQNLQY4IBKsjN+HMxJ57mUtlhSNOV+
MOY+5QZYHAXlQYgVvK5G2Uir5QLXG+pHPOcczL6j6XHoAaA1BVNMjGlLNTaKM2y0
/xDfzl4Yg2EG0N7PB1DOohnuOFYBWe3GQKel4mMsCAshdlSxn2+ySa7Nz9lm6aR9
5jxTaJMhm/M+aXAXt+RNuANAdFrLTvK+e8zbcqXZtQHMfYCBZP9XhIpDID5Rni5e
Ucm9ORmDoM4wRUoIR5O03LNaV9tZV1r85j+yMM1FA/kkGeR+LfLXDDP/WfS0ENtf
ahQyi+db/UzHOz22c5zKE5nIe+oxqWyQwVvsdtG91uROVzmDMeTy4gidFzpDiN7/
oRm8opOcAYuXqTHoyP2KO+tOHnvx/Ohvo2NIUJVKxAMPjPcykLb38Rvzhv9wA/bx
Hp4fRcSzr15sF0z4Z1f7lB6BgRS3uEp07lkbJ+oJQYse9aOsF2MdnOLNA2YznH/b
8Tv1NtXkRQdfr6vj7u/FjdsmPnkeihidMUA1M9ljQfxmpfKEMk3P5AIV9hPKAAti
RR/ohWp1KyTtwiGRK1eNsVh0QA14a+F6P9ljfWa6rLxUtBdsrJ6+kEs5qSibPcqq
Ju29Kgt0ueLJpehh+sizT6V0htIal6sBIxLYGL20Pg88CkYaUlmORj8XkibJibg/
JqREZPAWvxFxlwO+3sWxVU7DFMS7VtIpwLdAelHCn9EBfpRmGB1irvYqairHt4Wu
5ma0uIPadkD9zzLmdX/hqih18rhEbqSDGeSeEOY5/HqpGehtkYw9WpS+3wzKVXIr
32HdmTgHX/BxSiwvJ+45LHLeuHgYtBqLlVSqR1eNiMJLmwHMDO/AQ6UCTBjXxjsB
UQs74Wb3fupkch38Y0bczO4s9rHW3gjT/Jj2HPD/wHsNych1tXQfeWaGvARWl9wT
HOBcUTlbbl72opwrZD0bhy+fAm6e+wUdjH4cnHdSubdkOGpjwUFHldZnXnChj/kF
C5dNyXp1BEqVGcVWJF7ik2yA2m2nYvzPbTfMrJly+On0detMkBKpYZlHF0R1HRl2
Gg1y8ENTIcxqVqXqufh/nlBn1NwzswEdST5YSBlA4t9ATo2ZFjgOnIgsexmHwodi
pBdK5M5ao54uFe7e3RJF87ubW2ULy9nP9rMYsU3BEBm9yD4j2Ebrcr2VPFoSyy8l
1v9xhgnvpQf8MkwSASr3NHMye1J3hdyzwpu6IBxXRxIne3wP7FFE6bg4D7Lt63h9
Hr9f3o6DCfUj5+1RcfdkKOjHe2Dut4LZ2WhpI8GwZbWlPQ9byENDIkQJQCRbbBAm
ZG2S4PDwXiTCFrmqgQ0I3DN2yXbJzMrSBtqPYndQnvkuromgxOrzwbYTKNkJZzNr
tt69GltcXtWlFl5WZFue0H4Ypdw/6k5zOJoCOpN0HBM+VLCaJ2Ue013LVyE6OEur
929PHPmdqvg5WEDzZBvLv4OuYNJ8HKWH+/GhFwLQQcUlLfjjmFbBnY0Gf53qJrMc
bH5LwR59HW4WPjryBvzbj/JjayHeCQhpHLqscW0pqpAO5eFjdfUiJPOB0ACeC37R
Wb/RGUriBE072PmcjPp+qSP2OSFXEY1rkwKs5w59kryHBv/WoYHtcE9IlQ7vKuZV
Mc6g2rXckUte+AW5Rq9eN5wS+69Uf7nE14tI7tIGIH1EckS/xzooIWrLHtJpQV/V
r2WnixrOv1hqtMotx88/w7FXYrZxi8nbuL1mSGfzumNc0U3ZSfr1SGBcqhSqks2N
wP2886ieJud4+zauT5SmrES13LU7T7KB+U3lae28MpkFwD9Nzt2CA722JwThB0hD
ifl/TpFWCBVyE+5kB1cSG6tX1kzxTYvmvy02ZDMn8nffAZCI6WDbkxomOfUeeS6j
19FL+EWrcNzmE87C1F7KQ4ewtrBZepsfWmC+hAdEXPLC8NH0AR3zl/B3sHS4NxRO
MExUyH/JuZ+beAx8cFcu6WdHnP7ikYwIhy/zzlUvXlue/lUmSiJRIwY9dCudtkPk
jVJDe8tWew8zatUKCEnoL6kG+YMPbHFmDSOz3L7DCZJBXJk7cRpm6Pl3L0l0i7cN
QboCv0ZLWGTFUoGjY0yO094yh3O/3j5ASWAlnrfMr+27F7SLeCIuyWn2jFq1lMU3
WHcqfM7tZf+13byOEszWdC+OurUM3/cBOBH87DDsjAp6wVs5bMhfaDeosp822EXH
DBnmmvvTkzJsf0+BnnlAPgbnuQzZer5AFSE1CG/vFOTcXlTt0Dn4JFhcV2vrY771
jR3f4N2hSnMQR7m5zLj9EmQqx3To2O2pxkup5DpiIyyq5MHctV4+rWAQPHjlZ+je
8qSCQCgnSmKIAVE8YsdPF27F2L1WmVT4m8fdOOQSqCa8DeK0wms/ArM13RbnU2vf
ZBWYzek6/nr9GWIAIXwkNnnwo1iE0dNJPSRz1vFiCutUmDX77tfpJPS5AiMuB5SW
vU9J6IDlmkWvnEHgBnX8av0c6WRwUhg1Ytz8SiOmuxsS1HT42LZ+CTYkUpFExvLF
H3J19aaESdrZ5ljgrHzXnvOGB6u0aBQUBt8WwmBrUIXWT1ltX8ZkWIaLFoSxT2Ye
6HHjjHHHRWimV+fcGNY5t0wGQa74a4wwgy+O4EQONPBuwhCbisAS2fKdSeIWv+8D
jxeUFsc7Hybo4O0lAunorWJ7fSvpfTggALiOVFIdDoRJ0ClCtJwWcbvLfQ7nrSoh
wYT6it6UMQfkW6pVi2eewwA2JU3NndkihZ32TqFqVKFnEgac0mdpSd6Lqtf7mEm2
vLKaYK6z7Bm1aKFCutQIm/xY+5Nfg0/955QZkxxuTolzCYFD76CoITjo0Xquryl7
haM5eQf6M8vSlIESV66HiQ2q1Fh0Ywvs4/5ukR/pF64j3BAeqI8tTaLHdZGYxuEb
3ejxNl2/tCGTh+SkTrOwMpgOchq18lSBuksCSHRhZoGGWytBv5YdJ5qPDcgPk7YB
CV4B1D3bYdeYIoVy5NQQkYwD6kxpTGvi3LO350ZdxBrauusB0kWI8nuiyfrakxgM
EPE3s1dNBJJBPHm1VYQ4txhM2w/c0PBfVsrmZLxCNL7jLei8KoYMvuA6OY1icLzd
xzhadKNuX7UvXmX1QUOJBXRqJ+QTlnuG5UslgQXYcLPzem+DTD3M4ToPjmK2HM7F
pi5IJR1jEGYaBEa9XxQStSUifUJeMlRP1mWpa/sk4mySLKJ40jn/n4NuwmqSKXVN
qnvtvTNoSXTOkiCf68qbb+7ROR+TZQKiYVboLg8O/7QD3ubtM4byhOXYkssDDZL0
x65KupQ0taCzbAcVk0xsFTmv0fH5ofGvOvPPzYeF/eqXkQxvlHnsQT3yvyD6664F
9jucycKII/GRLkdA9Ovz6+N4zpoOy/3zRPqdxJYwdBgn/MCuDpGkb4hXoh1bh3lo
RBw5QEP0kvXyGz/sNU++AzytuZVW4BIb1cIob3qVNfM1Aim0LooOQ6lK7Kt/l2eb
i1NYiQQ+i/n/HkxpOGh41iKLgqUkRECIpst6xQ8R/eBaYoyd77VoOUVzBjeToAwN
Wb7hfJRGgi0RQRThZgNIN3hgz06kUZYGZOEU9x293ItH66vZPRCCq3Trfhtw/GJP
PcEWaWSRFX2zX1uoD3MFRPcE8bIcN8fhWGl5/ovo1IQbVS3t/D+6pNv2Ueeh67CK
2D9Y7QjSD9FLvwY5fyhj6IqPoLCzk2/jVgVj8wM4bu8zm5Ws5PFCrquNOkppIy8/
g40te8iTvL+Du6JuOJrLizwHxq4bZ3h4WwNieJG7O2jGQkYB+QrFwOtdZ6Nq/SKv
iWrsgfT4XuBi+ybHOY9DlIX5BAa1qLb656KA4EMHvDk57SYiwS20M8OHrReQj9/u
d2oxbFyVFkhWp+T6OKTEw0ivSeMFEsKs1z5n+6RRPQt2TGtTgz82wU6rw2R71FRY
IbegW9t2Udejs/S6DzTotnRwE7u/bOdrodl9kcm7bWAG9FZ3yxwIv6T8hz0kdses
qxSk7bwOKFCimXTMw/bwVr07nkKA+CGkifEdIFlfGkGPqHrmyyGhbtaBk0FqQQLc
vNU1LDI71Frt5AKjNnP6EFoNZRTevn2qPdzHPiPt5T5Vogedq5QsUcE8Bddeknj3
zwZKOfRd6Ublfo+hXaSvMai12qpAb73ZOL3yPJ/XHxKJ3kcgJc1d1Zg6sdNsr8+L
Hi8z9a4cpc6ooX/34D90kz56y8K97FDUY+u/FelcrDcaNd4breIx689uMYVdyAgp
XY6q52IXX/CBlNzi7UFTivK79VBUu5LWUl0cjoAG+6zKR/ChyFAuE9ykzAn2Ry7y
JXr2o+t8ugrgXsXU+Quk2RkTTInfMnUZWDlMVEsmLOXkJY8OlW/L1PHJNKMaVC4J
c94cbeO/itsNgEUd5xegWpeDft4U2IvJkYR3wWPhClIH+vFhTMPAzBvFsAtUBY6C
HgDQI7XdvXrq7T/S8jPNoV2wZKn4xcUFM7b2iqOqUhJU8GfvrZroLemLLdsbvPaR
6tuM/w/cJBzZ/xvqKVapj94Qx24WnszLuxfw47bDzpSa/eDO4SGfq7Hv3a3vW1Gq
NeIclEjW1erhLYVx+UQd6WLuW36KMQ+lIqrRqiH/8AZkz/SkdmXHXJ1ntei0YmZ/
3gPEw5Pub+A4pWuKp2QhwyF/FX3fMmOPTBFOKC2Ylo6C20KhgFqUonAi/MYVYwZm
yk7m2nJNdCPecAkV+r5/DEBXUfIVskujZoP4m4Z4odLXmQWPmm7tMAfBqDcKG2WX
8Vq3m5Ao4DfRVsU6j7KVOQ+XcveUtMc/gxqiTyyZsCnUPjKRiQ3dxlaI7jwwzfqK
kO9q211JAQ4VGOrLGpGsXMG/DpM8mGDzT0MHE+qphm/edG3MLysMN6tivuHUCqNI
9pd1gQq6GGN3+o3H05wq6OVGLnh0XM/kP9IXCyrzwYcPbza8Z7JwX/MU0kvVxsS2
PBQOXP6x1zhg3vAavLvZiOLeOZMd5GL25dnK2doc8Y1MYw/v/DqxUUyxMwid6IWQ
ELiDkHxCEy3ynpyFFGKDdq+VWMgFbrHnh6pY0R7PAG1b/WL1gwl4E2R7U3g0QdTR
k+DB+GJ6ID9PakEp7EKAmSUTUOPqMNd0kkKT1vOl0/WC4T4aETXwmqAO5HiA88Oc
0W3dKKBeVlFtbyApxd+NodXyrwCG75LGbNQq3eQrjE5UuX3TAca1/7Wt3SjaBSYN
h8VGah5PIBhOIS13CQw1+nyZ0IO6dQLwLMuZ5vBLTPvqYiv51O058JHlHXYJ7vKp
ytcXLPYV95HUW6ot05xAeqLF5pJKBxqmP2NICIBfNAjtJ7LgusoVjvUFnDLTl4DZ
yZQxu+EqDNLGV6d9tr7U4N7rwzL0i9LQKWAmjhN6Yv3myY1J+lHyzPdAySzLpU0B
YNA9TbZtSFpGnYfVlI9PwCX10Nbp1KZ2tV5E+o7YZdaFYdQUFwtqU8c5BN0RIYmt
snC5HATOUTy1ljgl0Wi5m5jt7IUVvtFVjO9NmLGO769z1rPg5LIPhqzle67EHhYD
tAIhpZe30IRQW2jS4mFf5kXiRjEsrQ0yGyl8s5OCbp6O9d1ByskJPhx/8A4YGfWk
8gRJBHs+BofSJEUTpAoexTgDfSOqsf1abFr1qRoF3B67A4MEUfLCubZRLAZlgPDX
W+bUUS+t7tK3F3lEb5rCSUm4oiqvmOH0Fbncw100kcUqTxTD1NREPiWVuOWtXuIX
W2KxT548WxBmI/TaoMOKcZAtZO/Ff60AAApjkzn6XNshMH1x1h/jGOfXfmIC/b1E
W308dir575l7R4NWVL4pjFHiJkmr0c4WNX7DilBsj14x1MFOxAM99R73gJ8pajDP
27VkjGofoGWtaki6q59y8OFtZJ1RBhoT3n5eNCUr2VCozUCOXoM7zPlRmyvLsunz
4nGAnvBCarB6rJ4mVzsBxG9mU0I8p7PipLqj7I05O2s/yGNLcpz2j+Rsabx/5wNi
nSUS2nBA7leES6ic5a5kPZrsbhRnT1aAgsh1HxRxq5PdzTPm/RzuecFjN9hbnTVm
XrL6dQRbgdWppWh5x1WpS6KxhmhIMVQvGTLDEmkfeHETDci/35AZ8TJzzaeFOVfj
8m/VMUC96nvB59WxNwIkTsu9mdL+EQ3wR0/q0D2Kig3SXrPEunJXaibEnv/61BwF
XXLBmkV3n2G49QITgV0acPfAxVE6hdaADjxEsUX6wQSyF23OzWsYL69+BUX48nIZ
WRZlCp8ySG5HTvokN9Nqgib1aODpDLwNrpX487C3fMKhYRItdhOx4zb+HoFm/PHS
QQKL/XA024QtYs6YGERnXbZq+MezqJjM43jXK9KO1tYLvvfS0AQMTEpiwTedh7DP
0uPcfRya/XYcM4+V+QENQLayEhskAU/PybYayPjTa+oAJ/sCkCOdrGuwh6THLM7D
Y6WdAPfvLEx3GGdh+YYRmIDer4UETNriiY96LiRzFMPWKrSwfh7UC7uo6DY+EunZ
aWDynBozkT5RZYb7JdTLf5Fn+Kn6qX/9eKY/0v8PD1plk55saRlZFvTSsaYHiIFs
7q2z7ZbLXwUyfdxuZ4Y/TZOmngoCVSBddGA500tlb502Z/DUUnkXRNE5wBjXKv2d
tSj5B97MmDuJT+o5bWwUeDpoSb3Q177tNPbkbOi3ZoWsbj1Zo+hpP6dcWlTyLm7T
LeLEB6R5M2iI02qxE4YM6bZLuunYc4HJZZuM0vkhypS4rYAH48VVDahoZqdXWc1E
m8JxGjH2367KSw0aQIMMqRUO6lOVi2beM/HuvBgG7xX1LrS7hGNxXmPHdHqyFJ7i
3Vxj4nBGw+O9aQPQZHaoFfb5PuxMPDUo2JyDlYnHTHo5i0bQtBW+RZkoAAInGHJf
qfnPlwO8OKeIBpyC/w+29DGTpKthzz1sqlupiT4cdN9m7JCUFRYn+SjX90xMEGct
YsO0TA6beI75EeThET98pO9QxKRPX2sQAZQBUp7lbNld/PCVOYVBgMDcCrXhfPjQ
e/ZkZn8xZmUWBXJms6k3nJxV/Ts/GflCWSsr3OkIk0ersOPi/uvLMwA+1env40WB
v6LdQIelKxcvx9bqNz8Djjj1rkPWL3ov8gSkUs7sxQ9QAwJo8/Oibqo5NIou/APo
/e/fIi9zbiyQBPYUs288591ODF0+rRTWnPESFfobkbwSGr5+ZDcM4Do9uOH11Eq+
4m3r7pCT3Obg7x4CeZfF/74aU/9EwOaMsI5CWIk/aiPCz8VJ7wXcuKxNgvWcakVb
mICCGxJ45IWFGGz6zkN/o6STB2rk+bwweA5KxNBFXvFyBxBRRZQMEwG93SxaTpLk
TucozuNiQjhsKx9OkhuAG1GDn6pRze6MVNvMlSVvPxPUDJPLYsmT5yqKlm+2G4EK
GPh8w6+jHuYkSq5bAhKXeFFRo0WXf78Rg/wBlLziLQEK1GBjekwKBB7MgT3Of5F9
WLjA143op+6oYkUbTuDde9rRjb4O/WF+UnmtsUBFvaFD6rrzc3cQ7fmp1cUVcZo5
FZZ7LbF0oAfBKNsQRVmlZfVqa5c7wJCeiAys3GL3oGChPZsNEve30vddzDOnVl8q
+ngBbfj61IDjnIuW4j48/kKJiqF4lpCCRScD4ZAZb+qClKwGVA9phROOnsuadlCy
khyGiOfb38VFojkx+kSCx+6NlJO9jEvCPD26W/WUJ2TmSlxqWCr8Xrbc+WliG0VN
Z+VjyOICoiXOHXWUdviVn8DtmMXeNaeW1aMRLcY201mpkiGM7qv9BWEOQT9o9o/a
UyQx7OkqCPbuD2N+mYYi81yEfn30+LHC1y+r7eo+JBoZe4KF2eIcw5HJ8y6UZBPz
f4NmKz35TAAETuvO7lsslu47EgW4lEwsJ3L9v7Hfi8BXqf7LMAkhojhRSlL3VPBv
myXvYqSiSrYTF5AfRP6fDov6jQVUUxjj+RRb6YycqHwAplD/EcehQDr69IqJEo7h
Kc5u/nantRSGj9TcGjz0gfAPigP46hu1VFjkhg+rio3xTFeTnR2LUE/0dBsUiNum
vi6e6RlL7nxbgoUQYEUpvnjk0GDMKHvr3yEHSNqN9sCgvzeyGdhIMJAAy6gkLEbV
s1j7rISejdZl/wbGgzCm0u6e27vGn+uzD4pJZtFba23jRtOFwny0G0l6Gzr62eQe
fIxycU8iEnidezc9GPV77fGrHO4Ssa5u/PwFKALN4ksEXeAR7VmAB0mcQUIm5F0y
PhA9OXzEnJL8u8z+fGA5V9VprefF/sabYSWDgXJDfcyn7fyKtVtw5TA76jsj60KW
txAJcmwGCRHkx5Aggw85HTRa7tIX4xm3+wOWY2L/tj7ZO2cgOz+oqtxVYf6Xja/L
5UrTjTvPNzPQRJE7OW7OC/IIT7V/rf9e6vNLDoXQJ9txWBSTkqDGFtii7xx5uHc8
Wo1vzMM85MQdvn10dW4YlYw8KK2oVk0aBghpyOOVLGk7Iw8uXUG39lvtmZgEGivP
mI4IeiodE9i7G0JpAwP+uM3H1gQel/ZlZaUvRbCHKf5NWgS5R4DkqIVemGRKCFw0
7UqcsLiv9Y4s00Wn22Sy+IFeCiiZKE7H+Rr6pYefRLdUPttV2U+3EGVaIMvdM1kh
UkADl/oTInDTY3Ad3mK9Eb+mA9kqy+TDTIve4w4f2BWhAX5+Q4M2bou4pqYEAiUS
GQTqVomU+0Z0YF0hHeHv4G3eVbrHBRLR3kiU8mBVciWp9i+AHOedcfsMcuBYkEBY
6kSf9KS/+dONt13KQXe4NBC7LilrOuJgOIrlfTuy6PSNJ8VSWaIYzksY4Ts6WP/c
7HZbos3kEJGhV57z1RUTx94UZvC9Lg5JIcwz4/Xr2zI2daqIPXw+o4KGg1Qm10JC
9aF74xX3NnKZWoZN9UYBl383aWwA2Mg3penA7P5F3MBDf8EEysLlN3OVcB1sfqRZ
w8I3zXAbCa3YqCvKcJdXQWl6FVG096oUvZxHIoLsLwoLQJYG4ZqhYQunCSdtWWtY
MwDGMcj6jI8iFJ5LMVlLypX3ybun7zP8fpdl8vEdvOtVOXLsrTdQkAAY8VPo5VPa
e8bfV1q7xk+kHCOeo9TsRm7eIvhjxMW8PwiuEurXE3So6erK3Rkzm/dwcwoKg/E6
XLVbqiDbKDVPfOiZlfdkraOC00ov4ytMtzVYqlA+lKaSv/KjjKW6AjFiTDJZFRci
0RI4cJjsMdNVmchjqGul2bA1v1H4o0NnSN5DLpTgJG6FwK96djbbmDe5U00TKJBx
J2V1rtl+bUQigl2JAb73ij5SNFGA+dpr86O/Jn7J/HbHMySuLOE1Nu58vZvs5Ly/
+Wv4O9MAjkP8VwpgGJljMvhNN0tr2wuSAMpErKl5tGBfNS2czsOin3i7FaaVp5Y9
FTaqJKEDD6yBGr/Oo0EpKdiPVsNbZkMeswXoneOqHeKugQTswFT0vgR61yq5NfCN
hRhVffCCENZAsigDHpKaHbOrQcQs4eRKLYlFPYtORpVi7/Vqlfl1ZmQWJDW8k9Rm
F1icrTJUkamxWXhCZkmDCB8Cxlzgz1YANceGhlf/KwprIkUsRy8GbMFCBg8YHlge
9fjUZMsft2h+i4tY+2vCJNr9AVCRbJ4HLSZbApLQAiWQJcqbX7mW3VS/KmhEZT5W
DkNr6rQYiRtDGyamVapvtWaFGZI6CoygIBhyf7VzNU9dAQmI9ba2lDTYfRrVhNcf
cgU9Y/pPFMM3qG0GcNyyoZ7uW9M2QPvauKo+E5IiGrDYpnD9XvzDPR6R4SA/WAwk
GscJMI+7GTDuUzDjtcap7M7yaAaDucSgy1Pf4+OCAJLT72h85w5a6t8qUzFgRQAI
RLWpFmCgZ8hVuUaYSgz5ukA/OOMW3mu+7RzPc/gxbPycJ9JDSGh0CspT56V3ivIn
APupvoVwZng4aHlr5Xx2TOfe+fEWg/tWN6p0Aebwrp4kt/R9+wG0fGGmtcA8vS8f
HF2YIXjP1Jp9T7/tZ5VE6xC7ceuZUuCO/PIXt0hTrwp9HevfYP8CNP87dwvXbyOe
BxJW1DsIRBiB6k9K/7K/JUB2XRw4jzDLYAq6MPsq1EXE4W/HRUAI3w6Hn5ai/YCQ
qujajBlEqDGCVTzpsqIP5kBwybMceXWWr7TQKXjvT2Awe/kq+ydN+TP6IofCxDyt
sva0ce0AyEq/sPmlWc50O/Ou7iplWJc8R9iY+9iwrA3EejaNH7QsuthCqkQHvlUu
Sij+9QyG3SdMJ/B0Ct5uuDUVYxwpkarNANCBZoM8vupgEMrBGSMq//D94f/YAHRn
mqcPQ1jJKK4Q29FH3mygWP2JPYW3XwohnUUPfIS8I5wyghemPJoyZNLtr+7dNppD
5QuOz6estirhznr7N9W+n2NwgYySPsVnQRZDE4jjJEXLie/9/QsTtsWfVF3z7JCv
4IPbqaEZlosb5/ql4WV5yivUmk4miPax1DvUWkRCcezBymR1k+I/X0/6FnZEdSrS
6vvz8SE1Ju0DWiVjAvcdufEGw4fK9OCC9wd2iV6JrIA09OXSgxvJWYpe8E413JfO
soQDDUkNFHJdn+A4ap1fBUkA3bHa45j2L3ntXv3f6QfQT63bocfs5gDMybk5QXw/
DYycf05ZJ+OfFXoWrtupa2qHdHOSIWZLAIDNww8awQ/jqvWy67xn91NEwLUIh3rC
GtfiAEAMKNzyvYoiZsEN1rL46L1PTNV9Rg4x8qYBkWiynvZ+MNaU/2nYVynkB+FC
CpkeA5oKR11Cl8K4n97BY5BohtPnVlIP+mks0sMqc2SJZq6spbChvDbOImkM6Tic
EthrcEIRoRcXfJUTJBA6uFYzJL6w524GaPnDYfKuwxvxv7zjR368w3WfAIjGFVh4
mcBWgvyVO/yc7J/IZayBNQ+wAK2x3r/3EpU80hADoAUdpc6Ui5qYqYbRUU0hGZfo
aN46fPA+/XoQWyKfxYXoDvYcRyn73mAzOZDwHKKJuiDlrCzC5mGXqa1OGtBBa+bn
qBjZ2ioRe6zJWgLeUZjyw4TRvq8iqMR1l1eSMCqz5Kp6BRpPvCSjnMnhe9YDZZ+5
zw5Lnia4IWLCmB8i5dmSVH6heAygYTM1Kr4PUmYtoO6pgBob4tuxVq3JH/cncP2M
HL3gWhjWgTUNemMUzg2p+Cr2dWkcZDxmcNM8Fdnv3QWZ6buodROguhPFiiBssAqI
rX/zlEfWRl3/NEQzNT+RVwoRCTHa1h6FNwdbGQkC1iOttTFqJzF+SQsMuobNDLVG
+Oukc8ELHKAgLCniAhugxtDBwDl6+8+gtqs3H31IBwIQ+4GDsrZi1/gfIlJPhxjd
I8MYu0D+uY5uDq3MuID9uQh8cH2QJOycMWhGWd+s69emjhkcORWcitZg9boC7sWE
vqJYfFaGvnE2sG8NUIa8N59fwuycuJNSXmwdnZxW/dxxAq30/Xax9BEUVbsnBTt+
rNfNmHUw/syx1ydsJ5RBi6Sof7x2Zd7crbJi5JErtc67Lu2SP6EJKWrvPsHhV5lK
5kh1Ly2jLMyJUqYkaY6ITxPrCrJELXmURgHxEJBSK5biGOeqzjk2lsU2na4LIQFG
fuz4m9KLeF73brDjamGrykPuWzEgv/TOcT4a+VgRV4mMhlJ0eE8tyLi9mOb/fhgw
dg/qpV+386UORZj5m4YIaS+cyZJ2eMIX5+I+QIkkAZFRJaozNchvlSvph/9YStbm
UA813Rh0MyKReQE5/bcqFqksHmfLbLNpimLZ4O/Im3hj0igqzfsKLWWggVr3Xama
mPT9KpW+OXXly4XFkfcadq0VBNNAorYOjZJmuANeQ5UDkZl2gfFP1NUk6F9ub3Bc
B18kcBXLn6wzaYEVzjDNd2RKcU7zeF0fyS9rKQvOKnaDfAr8V7XmUFdJApSPkKgr
lpPqJ3jfQGPqml96oPtj51lQfv9xE4exCjTiN7frajhEiLX23rdaM1eUgHrYJ8ld
YzkKr+AxVQ4QRDksavj/ZRGBQBqNWc6OkqxUjvqeII8C+rkiRtZJof3T8uVol/sv
sh+UceDmcN7UBn9/lrErZchG6g1A9R0r6x7+xJSiLqDA00S9y7pVljp6Bffq7o4E
oNSAkdc1kyBqTt6eXlWmkPMfpjMWJbRz356oEmz5KsxJT+1T3kzKeA99KJ3TFMTu
oCKo3WAwgc1BuIvCxBFDe3cnPNdtk0Elc5ka5D7zvltyOwXfhsxn/vEI1VZrnU0S
PYCbz9JTGbvx6vxSjcx2GyrySDvGQHldw/wgm8rHil6MIpitYF4PTyMKE2aRNFIv
3S5KK32bKPD2CLyD2TyXZQ3N7uxFJEw3bzXcsccONymS8n7//tpKobl/0IG+8s6V
0mnoisgdh+zOfXuqoAQZSb2gOvUPnQX7oxysmXuTDEr0FBtreikLj7HyHf/4+dfq
LWjhVZXXEUY/grIIDoPiYACYrcRCh7s+rXLyaoyqOeJBG1YSjFlLBMwGkA3p+z/F
nZfC/gZlVVvWKbr1IM7FnU0X5XXYi7u0nZRBfrAScZVwtvNFkx+mL0E1E+JGvG3W
Sn3n/UJbA1Bo24BMxAQCV0rMs2SGKtJRfEZX0Ioso6Tpd+ZFzhfkFzUVgg5V8vTY
Xmzjg5sVsX8tVUBRqiZZ8A+SUetkbhhFDtCBgmkMPzZnXtwQ8K6rMjKOxqM/eX8n
jyUxST7e7pc31xoFVnsCH0yyk6F7vIQg7EBuQe2+Xq3Ty8YlEjDaOJzT9xDiTlWW
rgtSnyT61qwqG1f540uFsJOyn3sR5GZ8TrKtTR/uFyHXTTnZSTklLN1zekYeMN4r
8S2NUolVWH7fOlSJRMos8N6cSBWHKnmndswol34w+8koRAeB0jDFDH7yQPCufckI
aHaUSKoY1bnPW34IfOOKYw8Ra4NtCRU1U+s3RMROrMfzTriPddbnx9TvE8+qT/Eu
HpbDM9c50vn5lJli5yE3n8HOK3WWYIQuncwx/AaVDYGZ0kDPSIcxdCGB+wXnkf0a
5s8029tZqmSeGkcyHd7VHCg/SCZCZA/C3Alxg8khaotY0d34OfnTqsCvX4K8Nrw5
zbhaIV/iOQJKpV+a3iugxpiSgkqlHFaKhcuPR75OYNo7nBk/68nnNN678rlu3coz
OG52fA0EIOlqvGSPY3O3ArqgU+zjE2edqeCLwWuXbbAzFmE1uX86S2mrWc816/2c
9/m0NZdIJQwW57oNyenYxLA/AuvP+8Ip5aQyKkUYnRyLR5mJzwO5skx+bDX4Xn2x
/T3wcRfLTRUQi4omxBpNzoGN9FGVdKvhdk/GoIYvp2m87WFPW1fwrzFWzRIPa2oV
wdw5ZPCpBYX+UwlbK0v4LWTn2qw3/gxGsa+pgiZpLmbaGO6o3JkWeT0QKhRX0i/7
tAmZUVi3NCPSBfPdLS17le6nmH4pGlRO7nrVNWScj2zz4DVlvXWn2+qpYoJdJsFP
z6HY8eixcVGZVap8+4wTOwcErRU1HI7NfTpgGyNQtRjh1SGtXjDb18CbEYy/iP5m
66VtGLbF2jS3J1CBu+Cdav16wFtiAWpmLo5b1y7DdDf48BjJT/5eQtI6u4ll25fU
zsVmUaGaKpLZyDDBIIsJzrYUMWb5xYmQiv+N9/miEjbuefGA+bBFTtv7ECu/RL/K
3z1a0yHQE6eIyTyZ6eTysYpsKClGb8rm6rJx2CqqrfahTeakn+y5XwSaRDvnFoLE
pQfrX2dzwoWdJF/bw13ttv2R4YG75K+xPNsLox3+xvYp7bEIud1BF5MXhxd0EQfk
EZn1lg3T/hZzg57Yv80PyJbhcssw99f5RFaT5CADR/Nip0PCP0U5FdVRdQ9iCRRR
8afnWz2hCTlhGyigzXf1owGKrxbeTW4S3lCDdosDggMv9gA9miPXP9fQ6Y0Q3CKN
Y5ksI0VTgizTx+jiq+CIxYiT3fZYAKyNbkirpbWb5XLVAB7cBbSRSdbvF7/455Qp
3ohZK+STeARzigCFGCpg6HfJmgwRuYBMKRhQGM2b8bBynahBtRKxmL1GtjhG5hEX
cpaBcr4Y6TFVYuFLRtxW9A==
`protect END_PROTECTED
