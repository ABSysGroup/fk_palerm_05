`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l/FVEGETWgBDEhIAJ9Xj/E4TD++Y5Cfsdzw15FpbxvulW/e1+eaDKBw/kBpobPij
rpduj8Lkgwit+lGQMg8YuOWdu8/Tl2Oe/IKVBtS3Uh9vWC6xEA5NfayTgYZPqqwS
vStYRMk1Y6WWGvj8qpB+7lK3WgniXnPGjPfpJ3BA2G4SIkA0ZmQbckI0IETyiGt9
he7NdM9omcR0b3916/3/QEm4PZJLieLLHjs1hrWgVYboMzVEwCSzr+QIs5a6vscc
cxM8x86FyrR9jC+lc0NFIrzEbZCNwRebv+5W4yN5ut8naOiCDpKs9s1/l/iQyJF3
IZ2Ah5Krj2NQVabnbMqUWPO9xHIMtnmDRK9wT8UrSOP3kRl6RyldeSLbZuaZLCTB
HPvXcbevT/Cy3tdWKl3VGyRyoWzj982naA2rOS+LNcrn4Zeo1wgz4vub6ONJ0Si/
hzJrLBYuw0SNt62cNcPto0lvNE5IoL3qMCnW4WSENmHKsI+V9hF6naFWoxcXk+Xd
6Ky4zf3g/p/0pCPDsXtTgo/GrJeiw7aUfgdtbZ6feSkewSEPiCTmn03uYI95eIVD
PMJJXlniwDw9eqldpYKFlgNyZ1zz6NA5jUiGIHXhGuzA1w9oIYIm3KPRawGvodCe
mlZFO/ndYGojfx3XZqKKP894njBPQhfBUxp4Ln7Ieq1BZHelrkSlCmCYDECxwK9g
oEwS5XVgdY1usxLY+KvXzGVrci92CwqdUsXpP82FvVz40UN13e40aL72otUV6R1P
FVFGWFZWcoKly7W7vrK73vxZnHXVBXpMhfO89kYhxc7xO/l1tyUA9FwbpXDrPh6S
7n6DKcPgOc4NYUdlZdlV5hFCckQV3iMYEWYX8j0fjAmS/94kU/CAnnqM+rE7sN5Y
DshobN8Fh9KeOF50eFScwUOy/vPnTV1OFtcSeePpslqZ51zmC+FzrE8Mg5crrkfb
6v26YgaYKiIAiO+xsrl7G3f0eQc//CujgeP5ExD/W0NR/UDwvYZBZIgcWz+fcYuE
99KKSq9BHalqCLxDDb957MbkIoATE6zje24Jhs5SEUldDWCWQ9SnW9AoMMIh5rtO
tq56G7Y0y5kAzBZJOePdZ8yW+BW33Lyb9PWFkHODBzqXPJ6QtgzAv9V+bCu+zc+7
t5fg3p4PiXrRXJqVTsZoennyjoWaPRa1ikLtrYkHZYu3YIvLnoVxqD9QAc46JgiG
U1DzQ01h5qTYp/Uyxu3hYH5rSE7dgaCfSIvm1ZG7DLLBYqg9UhMOfpGC7gK57okN
ACylIyXVSkplxetUwQVhVoKFarx/drgMBVDyI9lXKzJGbKMTg791CnwomvViC91b
2bl572jzvw1QGDk+CKbXAEnibDmo7Jo8eEmygxw8Vq41vq7xGJv5OWlhSizc4HKj
TiB6z+TeS1cGxOLeGPuVxJQK7K8lOMfHRn9nH8lqq0X63QOGPimY+HT1wLmTbwdj
XDh0QiUA+9zr/wuKtNXowZyiGCjFnEycpnRIrHGgB4lDccabFo6+iZSO/HpCpyNz
pFQSM6KLfb9HsQdih4Eo4vlaq6Jqn3itgKl6n3NgEJCDNdfn/gGcvim6S7QU8DIa
/LJsI0QcFT36jLdpbJtNSG7Gr2GF1KbzKodf0+JCeUmGmdvzrfDHDlKktYkcoPW1
gZa0qCdZoVICcOXC8mvdtyta5/t9N4Z0hGi9qsZbSlyD9YYu3HC+cYg1nPoibtGa
2LnLJqSdwo9c+j1lsXTMf1MHBOVwQns1aJbe9aTiWC5JxjoUjO2wIxEfxJT8gIbe
pMbfuXsBa0VS4z4u26/tFsW2IwVb/pRU8dME4tlwJdDL+zZzjdrSwr2vw58Xp0wU
6KTecWwUQSXUtWbGo80jYeERxBramdMqPDop5WcoZT0JUfRmLDT3cko6xFL5VImw
jT9kT750q1E/O/f7Pdvx5aHKCDlEb0VlVKx+LnSoYNzQzluA/D93sZifz4wWMx+R
dNY2ik6f+fYOyJ16Nhl+0Ee4RNhfb34XEUNONj34WmFLlfUEKVq7wXwraUJgcn8f
YsozzV5bF9IMopZ8tYIXOs9MRXZ5zhvja9ozKoeDvMMvelyLdNDg7lGEEWYh+QBh
0b+jQXGWQ0XqcMFYraNqe8V+EZrHyqKwZfvoDE3vcnyEZVJqisFLIwO4/bG/lNCN
`protect END_PROTECTED
