`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nuh638ZxljTI/6iO0BtQYv8w1P4vCZ56PDS42UwVbA1W0qQX29+DLeDdRRFfazo0
XvcwZFiKz06f3LhJd3Ro0w3BsAnSU95LPom3L9oBvnxaF73fB6pa8OIUJoYOk+8F
Iqt944dJLyXnpMOGbNLhrsDq+dV4o0BzU9uYOn3mWI+o7il+rvJbvdbQok4GQnsf
UAj64d1ulBraA5pzcfKkypX0bd+dQ00GxKZ6bcq1ekPW/Vq3ZMuBdYNMQ6F75dG/
9c5sLdv7lM+IqZrmhFK/2FVBz2GNlHhDCoSsCKmSZ+DywLBRmOBnHNv8QqNuKEtX
HbUdZCLQ9PdQzWEWwsDXgq/bZVKB9NW+m+0wFIN9WuCd587cpMDEKSu+ILnJbiWV
2/wNk6iZxPZbTyUFKnX0aKzPwqLNgXRJBS2eFXRlSUUm8SUq4Bhir0YvaKH8a7Hx
z3b+YbpY48rEa+n0GoF95Qjjj7FXTNzv6fl2HsSt52sY6qzWwDmGAqPNnmy6+Ymh
3VrO1F6sR/UAU9W0GpHD8PDewoLUYx8p3SfR4kCTd9jia64YQMmZ1KseWKYY/bhM
gBFi0ElTJUQM0GaQ/v3g14ykP2sy4m5mo1X5j4Q+s9jeJ9xrcVt45trt9s1kCegf
W1WerBSS7w3kWXtmc7cgugDYRqkmaU5D431d6mXh8AUmo3VW1zFJclkyD8UmwmTK
Sn30VyzKV9/Dlen1CM76kc8+Wd2gIrSNUk/KdP1G0PdZL454SANNwn/CpETTtCsz
Mb4L1ihJYNKTIxrO3+8AH3iVQA9eAEuY34hNxU1kdjMbhgw/SSkZK9F8Q7oGtRjJ
HWEZCUm0OS9akKUm4rAeqDuhWxC18Mli/rIVtOwQsCsjS6q9X3A2yoBfxHXNzGln
D5XcE+aILSB9i97dApqrc7ElFWYMqRIOnY+Q7ET8eTWYsK4P1XJNuj0F/hMaKsW4
OGgojSZfkk8uFLZ79ILxGYety+4ec34SoDDC5soD1ZVIPWf8ukc5MsNHodNf1ydv
nkWCyqgVDvDV/eNFz69XANnMg5F3WSezs6kxYukPYqyd6OMIZ98heSHc7grvryx2
AlIeHH6LTRgtLSLd27hvrxzyAriuMJ/yvAfZDrCBW79e0wN2rjADCAbJyO4NtOpy
LvKsRQ++15gtnbfk+Ye7wna8lMORsZmj32V8CPFj8c+zDS2Ps7pas5HY/pW5i8JR
WezWcxchoz9uoZ8+IOobQesXYXbaWXKQ3A3MtGP92PPqYK1J4o4V7NSnGbaoKXZ6
Ur2aXBzI/LVgjxwSbZYA3RZIDvVOQp6L2jMthhCdkCMNtJSy9TwVzB194GcQrzA1
PkzZ075JuAgK0wgdtq0ibsa3cQ0it3J7Z/GkMCpclT+1iec9kpBwgjEmgjpGSFks
K3RJD4vTGMWOQnVGVcKXmFGzNaqMSPWiDAFtvm4aBDsbob6tHXy7aPC8NHV3svdu
gW70CBKb6FQjtuUATWnc7/JOnEf3/JToKX0YASaBQaY1cJqIVphH/7wtbSo/NnSC
`protect END_PROTECTED
