`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RhakF63kgBY/uy9MdV/N7TBJwXDzi4FXYUceOCdzDEmXAnyzDG7Do6Uw/HwrkHpM
D62/h9cocG2+jOh2LtZQgnQWEgX4H4M6nJW0o5sMYDO2GiYmxrkqteTuNc0RSJV1
86ZiWYikK0+uOrn8qbny/4BKNxamp2+Hi7V3a5t71xK6hry39E1boAGftn0aMmZ9
FzRksrSkgBJFALhWgEEv9hqgpjVgKGu3pk3SqsH4xloiWw5jgNWqcJIWb7mNcWpo
g2GkPFhV139mbXfyTRAiqAPAvNUQvM+kat3NxLkw2X1hMTW/FPNtdfD3YFG3/jxF
9sIleY6dMAuuv0PL2RczzUZVIvar3MQf0WCL+L0uWx6YWgp443nF/0zAyE+5R2JU
QE1cIvrYKSPNxAw4bEQ58b2A8/K4Ar72+oEbC9Jzr1Jav4NAl9yYvLW0SSWCDebr
K2Sh9pTkeccSxu4AWLoI1w==
`protect END_PROTECTED
