`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IGvap8sPd9VURiv/1oMD9SE2UG1CiJeJLq1ijB72aUI3uo1qoAM8Z08sTsmzI7Gz
RJZFT9ADpWnyhSknqWFOTHomFCtx+PeV/7VRfCbO8k2xrQWmoOjD9Oc91uf77QHO
zN1rPlmlXvJxg3G+w/PVuex95PmThbJ73kdEboKnM7xexBccDBB76QE2Ttc0tFcD
6zJ/mtlHXzaNGvRCEgTq57UUNf7wGlYNJ/VGKih7sG5uMLt+vQlwY3JsuYKpOzPd
c1o7qVOk9Bb+vGuOkaEcNIh5Wb73GqUz/JaJJe/VX/kFShhMxqD/0cjMzTUjVPOF
oW2M8TP8PwYTg2if+baPvUKhMNJDYALwVke1/Q68hxE/OXwQTvC721zIMAHU5/Ln
aA3rw9ZqnOSYvOJKRsnVv+VNxl3IZY1rRhoIACWuekPTEOjJbQKoXbj9hbLIsFOq
4O2RLX8kC4eFx+47g0VROM4q1s2gKCSs98wyalyeHcD7XayUh+91M+8KE6reKd+5
m3Fw3CONrvrwAa1miwhpTblDg6+85pBgLpFemxl+s2Ro2DnIkaTC3RQQQTBXzHok
g1NaMCpahFE2wJDXOiYY909iZ8M9j64+Du6KXYC/N0nVWHNntreIwNXIV+c8t2Nc
jWr+aRb7OzjFVauo17H0ueuNQesjYltvAreWCu28nAKI+yx+KzHAoWm6NHUchqXV
aoUkknefzsDC1Q4m2fii8QcPd95+HxUBzPJRFE79JTypFuy2U/MdbLIQsKRsgNo/
Sbwx5qcshSxqHtEmOioXhA==
`protect END_PROTECTED
