`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
djK3sd4HhDYUnNI3ZLPOZXJACtYN23Kx9VvmfJs62UvuWzilG0WwARLtYKnO2Y9Q
9mXjsTzQgLrbWHgOPAgMmUBcuOnuJgN/ZhsgBcvjs581GYLp7U4VF+rXEqUQjKOC
FQXMD0L5vEg8sYDROAElxwoFKA7cATJ28CxhFIJVBEqJ1vSiBwZFzVBHrUwzNqE+
yr6oN+UszUAzzaOGvrP8MfS8V56mapvq9AhQx/8K6MsL4GsOZrQnMrxngikvfQka
K/iSHe6SzqBhXOB4Zic/6OKFiHJgjiJrQndxqn0ViZIZqPS+Lw4FgJ0ejONJ6bTs
1TTVDyYOpZ0VSlQ1+mQI1gcA3Txyn0JLzzV6ckOczvCLjvKgjziJTCsYsTWN22AF
goVqg+UL/bDEC3z2TrFRYrXKV4Qg3ua27KcuEQM39AqHXmFVrB9Atvw6D5KI9s+H
av9hvZlUOVgK2f0P2CzlwRcQdhDFoBVzJP7rDagHN2ft8xzfcFShVRN+JPBxcmTa
oVrR4pXjI0sJzgo1KwXI2YaoStHcDNcQon01SdJ6w1L8OM6qfk1L0Wfs0p2k9Cli
zO6KZedA9apb9ZyPli5cARCrGVZtvWXFF5+G7ozcYAWGliHY0s/3kFVFU5rzsbaO
EnBwz+SBi4JgYzR13p+hng==
`protect END_PROTECTED
