`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rayl0UfVN3Ui3Old2LuXwXNzmlrKfNeVv4kIPDE3ARetg5NM8ve2rpHGKWtoSFsd
YZc2mmTVel4ebuRf/56GU2DUg+KSUlkBh2J+6VpJ3g9yDlbIiQi5Q81JlEDnvnrg
tiYZEZpxeb3dikjaZ/cFCFVL8KFSJYpmWKv0Id/yo8sOmHxbnVsNCYY+mGx0+Vif
Wj+0nzuTz18dFTE4EgXbDb6fTM6OsAdn/JkIqI6LP4VZ0HrhmOnmIDfH16KPFCjL
CWpv/5pxdANzeT6W7NLpozLDLey/KPvqOPD6Bxhjlec=
`protect END_PROTECTED
