`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U1TLOBA7rsuGD3vwGpVcWpsZlXHJKwarrbClQKtav6YAcQeem+FhVgZrMneuthO+
c06ryCYcaAw0a0Khx11KWlx0oSQtGa/ADREHgu7GdaaNSrvSLdVYNsSXiEArel+P
c2j4orpGwJd+8C1zlEe6Ht9IMK8K4k7b3RaPI06GmOGSJ+5lyhpU3MgiHg2zi+1P
HXIGvQ6nBEdOQw64lfGgDTX/PCruVkVGDPqpt7Id7VXnG+dT5T7mjUHuAbUYgof7
bJb+0JQ+Q8pR58pfMmQL/h8K+M7gZ3eBKtg1QLeeuXKBhHbBjPlkcecP1pzaF2Wo
dPsnBNrKQOBcE6VtYIBU6w==
`protect END_PROTECTED
