`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aa0JdmMHF8JNhBuJiTa3uHeCJ2++4IuhhPHZFKz/I0vl4i72uNRIxYddwXBmqX6H
OskAa8oWZQwJKSLF460NwjnV0qBq6U2QcPHPZ9di5VcDF0sTYwwRRyOxO6aMce4V
c/YDcMoaczaBYaTFNYjvUGOjwVDbSoGeKr2aYIndy0TEorS3g946TDZxjOZQMkYl
ubW0LmsXVEZl8+sKq4HLvTvhFfzWZQQb+/Ns43ao8l3j/KmeH7KKUq4ToUOKtB8K
+RcfckI5Eq+MSI5ELsv6MMpyyAWA4i6IXDSGnWi21Hl22fAE4+GGascqw2dQW9PQ
v0hA7oXa7tTBnqyTKh1xcOVcthZjjFGJTueV2welY3dpUhQQu2waxN8/QxW8IVJB
TZk3UMP1S42DiF8VH0GJgoybnq0KRK9Wa8AwHyv1PmJaaWSsgq3kR08glX/Gt5Hv
X62jAGTSBbVuEYAr4UiCe5KTaMFyp/BMZ3lVAfEHsx0Pm4Ip611mlC/vNYP9N61q
CuUr9Tp8ug4dgQaS8iJS67Eu3HfEvBiYZsFXc93xf5N7e0uOmn5wYT6DtlITHNf/
ZJ42SVofdnnZTCMmYaLXCqpaDLStMRhpb599SmQSeL/D/X8rI5HCgZyqS9MDHQ2l
hXlDKcFmJXMPBsg2z0efqGvA8w8b1hUeFtp28IqeGA40W/dAiqeUX2EsrTSymkZP
IMPHksiIhA7M27Zmda9giQ==
`protect END_PROTECTED
