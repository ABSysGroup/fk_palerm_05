`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/s60N/yh8h4o1b6z+rHmv4mBaSELsV1eyfesKw2JSFRo4/BPD1xiXQRe+gMimO9p
ya6cNAvcl2S+k6vCI89cRfZ0ewxuKjyqx9II0UKwSqwjW3/R7vohsniyJuffDzR2
XxMLgbu4OKRSuRpfinp+5ZsDe7A2TFHJGgJEimrbXGoGUrLZnCFvEvzbo9ys3gBg
gMpGKA3XE34szPd5Cx5UrklMzGRmqMfdk1HeSulWBUokaTDouEs2st+siSHmiqxs
OR4EXgUptBGPkGLRQLPU1YBTwEfFOfjJve0h23TmHvLgAsK0AIVR6mwoSeOU8v3c
p+wRBkY5GRJWYzPqQMZ05jRrZxFUIH7MpVMPbGLOPE3boN0Lke3+T6yeDH1OaBYE
`protect END_PROTECTED
