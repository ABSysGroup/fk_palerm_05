`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x7+8f67FLbsLAs/5r10n/g2e7TFMhvIgd/dhYW53cM4E02ojA2SKKSgs4LzIt4L3
74E+0KMlNnYENE2YarNGyIDM0Xokh9LxXObmA082rDBJY+YzBxbZvFieXBT8mCOy
p+ubPRZzfjQY1NUD0fbl7GOAp3AvqVGycD098tIcVJqHfhicBrG/BgaS/DQmAqww
dVPzu/wF2QzCDQ1+SX3sY3NO9hr/OGGwsa9kseCmp5U0xU5HW9QhNiubNxKNN6C4
LgZxbd1ccMdFEnZD4zcJGbFK6piCX9BbLoys2vKPV7WpAC59qWqZi/Vc/M3r0n0T
IH3ntF5Aohk9N8q4moOmKS+Kwn5K78a1WwjfAtx/sDMd6mAy2HP687uX7ezH9Add
dXTYXwG6X3mdzeJj55LYPf3SlBpcoIVUHWHqYgO+eNno76NCx+WyQS+euKLxOAeH
8k6YIm9Voq8z5uat3uXv+cXRls5KxwyFdpT7s1fFp7yP2A3FyzlpKE+CIU0FkcPO
wx7tMZas8IISyjYatCfZ24KVgxD4XO6M2Wvsgjtuz+hA3cZ8iFXfiuB/U5FVrwLO
kos2ymRy2smRkYf64bWY8IvDpJ/km3igY5F281F+h6x8VXxWzb3MvxmQ39Uynfzs
OG68yLLH0iwOVjXeEYsgQq+muNt4rLhFfkarqpLd+zAsFc0fKmFrE1r/TRDoWpa+
`protect END_PROTECTED
