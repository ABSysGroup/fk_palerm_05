`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Inng/AKhQCLocMxdMbtgwPA9O7Pr5POasJN4HmSSIXXL1t5hZcjGKlvfOYpOEATc
X1j791EXwTe4cncjQCaNVFDFzpHWQ3BZa5jJaB8bdCZ4L9FO37TG8tzW2BAQj60z
Gh+f4yPSwmFmwI0ne99eFO4rLEPy04sygddeWme8DmiWJd1+KQvh3rS4F8VoProI
MkIOIzd5AbkeVeeNODMktU7lBJq65vW6KWDfpgA628e01zLqR+thtrLdLE0PoHLK
Ovu1uQ6wikQzJWKxnN9eRBM8blTZwzS8eQf21InPPqXe40wrC+C2bd3IvMEzIPGX
cC0mmDySNCdmGmLc1SiDHQ==
`protect END_PROTECTED
