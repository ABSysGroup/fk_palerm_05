`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7+TIwlDi8j6mxde0BaTtLw3S7xKu0d7mD+qf8cTQtqqDPshwT1x+FWPoTWDU1rGH
0T3Pdm4aijSD9RZrAtDCog68A3DO0mX2d4v6oLgDSzEPf6x9M6n8uvlp7k/tP4Nf
dQscjefcWRx83XSPqqm1m551T6NAly/QvJJeuan/L2+m02VUVVGRNK7u2bWqQQ8W
cyLMEUsw9Sp3ZM1G6MZxfB9MgP2pkBgaL2ELjRHKqtumWE4f/4eUBmaOpyDeOCMP
g1YTERJ3j5hny383BYgkTbEWGi8bN+eef+CHL8w0dieJzOh7lab73GbqPHnL0hlE
mDj7AlL3dtJIbdl9rBO4p074Z0FHQ8uwgBQaUhE9uOT2ivD4w0FGWqe1omhXrU8e
zzG5NYULYt91cJPTUNlrwh12H83JmVlEfAsndJv0hwweOApaYnyoZNpZS29ikwuG
rtSG44CF9rTuLd34r6UZqrvqvBUyCfYGXRXi71GAdpu59TGJvEBqEh2eW3OEupXo
+pa0oCAAHELfoUxD1BGWZ8nhLLiy4JkYl1C8NI7S/kOx+epy8vvbiMtQEsDymFHi
Y5wThsEauqmv2pzHA3HZeFMndgt/uAuy0d40pGW7sfA=
`protect END_PROTECTED
