`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GL5V3uPrPZdj4NYXdA7HCh19FLK02mt4bWbUrDFBiXisbw8KEEhjp5FUH0Zm5uOg
NADDKo4hryO7CtPT8I4DD8jQ+4jbXY/nowSvsUFkuK8Qnq23Ki6mpXMgjPfWeoAp
Dj/y6t1OJILwRoW0L+S7NhDwe5qMta9QFbkoGkOjKFwHeUHPu9dkyGKLvb5fxKjY
m5KZpK5kxL788Kg61vJxVja325KhLOuBzQVsmf7+4g37j8m4g35iqC0M4aPnAsqu
MlK4LjanoLXNgcepTobyMes1+KZF3fY+YkWh84+LSN6xsDyfDeE0tExu36UQwzEO
PqsinzcpPDddIla4JcBLKbHLvVjFDKAFSa1yjVs+YGNFUf11CKUH6hMAGBfEK7gq
PACxucOB5ieakHrT4Dhju4z9n5B2BnjZKf8PEvx8KdPMUjG842P/8e8Q+VfIAiAa
pj3xbK5MFY0t9qOdwLdSFeFzNjvf05bkrYXOwsfiZ8gB/RlPwQ9t3SxwW3K9lZ3+
tEjigDymC+Cp75KvMEZDv7gKggh0qanno5bhX9ScU/Ojj0zR8esJDaabuTlIoAxU
QFRi9suF9ZMUkFsJNdwPAEfbkbKgqS6lijqaU7enfPOBmRYUJGvxAih5L4zGEBjB
Jv/+ISuFfVC8UBBF0lvU0J+qmx0KFn5JOc9Ty6aWi8AoBF4KerrC8K35nBrM0aQk
pRGFbygwqJnO7W0Roc3h09rEbeozsmuGSiCYNOB+g4IcB4/I/6T1XXQnoSjPsRer
Qf41t/KM9a53kH4ih2htKs3e7YyEKZ6MrwyQrtjAPW27fO2MqOP55GkowA1KGfLH
s9AjgZcv405GRnPWGYd7uOhmQgLHJcjUo1wZtAJviyoDJa/jUAE/wZ9FgIOBMpml
13QuHwUu4WLXATIKb/YKYyAvy0xHWv1Q76hPAVfQVQenxsN1+tPUZZ1vFk+hQTrl
Mr5AdfwdTZG1EBYdr058GR76L28lmjdgXYjF5VuBspSV/uGsVjdrlxXbLQsTO3K0
25dUlAXt907EQMcziCmu5FxjJKs3tOrJBQdG002pr186vPjD/2YdCmQmBPD320ad
hBJYDsxZqlf6+hWX5YGZGApA7JdUUbRoA6wI3GurzkHstawKqxquAZZIDPFSswXW
3IKmMIe1ANau9soyo7ESmyWDvxHtxY7mPtMnXxOb8pHg8my9Oj8GzLQSIONBnKxL
2+/6YHtb4o8hQm/+hIEyXEsr1pap5B84qqScEtpxy0xSH4oP62LHYHsfZGTpJzbh
UfWeOkXzI6aUESmHPWVsj5f+uyvsw4pM7jRa34O4zTQr9JfSx+s14fOLsWGmZ4R/
7EcesN8Khxo5Ccdr+E+AyCTxzJhE3lfv+Pb9SuvTKS9FisVH0QKmc8ReMpTc5ktF
kil7x62Ad4Wsb9KDSS20o0ICs1ptRJMi46BEFVUCNaIHzg7FyN4Oi8XUqnON2Daa
nFVfiNjrLvNj84xVPe8KQ/WW5GL/lbon9yU2vw1W0L2QroYE8YGvDkg5eWyv0qej
B6QXCtUqly/LvT1JLu2h8CT9LtIMUbZipdnIIJIQVosVY8a7a4uap8a1CkCuTe7+
t49dIC8QSBhCeL+ABHEafbOHWqmKZinRKoG9Utn8A5/zl4mnvoM2mv4zb/eIag6o
qQVJnHW8qkRHKqXRYxRkw6cYu5wZzfQY37E7S62WwzLxfVk2v9yatTqLrpW1UNR4
b88H070vSsRg9XGQLlpIfMb9EJ6sRuyU8gcWB5zGH3myof5xBDbMjzIUgGhH06n8
ficS31stqyPvQqzegKa37VOU88xA9ICzjFp2NDIH13+jHVNrVDzoKj/eDCw+P7XP
i5kQn60fnd/dya4gQ1GK45OwWsM7ONaDWYh8VWCXBXqqcsP2sNmwxYAReEt46Ovs
7NHVn9ngIDkYHJJCI7BzggO1J1QLZDSTnwpJRh6DS+0pMZ3hW+Dpnc3G47+YOsU1
ncDCkZCg6tizD/L1CoUyVgpbUUF8zUd1DtxgdKK/xW07SPmWqjpRFoC+zcHyZozb
Jcz6eb0VqDaYPWtP7mOOLGUVoCss58fXe2iONZ86xBHIKjZI5CHZnw7S/yBoeJaA
/Tn/6ODpucxJQG/4VZXhU2j79503Qn1No11Oq7HSrPDsy1r3hsRjK0LwoUcrHITF
3GjrxSaVierGsSxmVKrsAntR+hxxzYoMViut8L5mB9DTbxhROV8Qn1CKrtkDCwuK
Gb2jhnrjGspNGxoif8OstvRDVdTvZ08h+Qj2+bJEGkb/3/tFzq6/81bakvYBWVeJ
xdAHpvgSh4yhy7TMA6tnZejD7BXwrWvAB5dvziZsN1z1GXMgTJA88XjfnWhwypct
UW7zmG2JCxHw922iUFcO7JZgDyq0a/3hvxSSloAsL9o=
`protect END_PROTECTED
