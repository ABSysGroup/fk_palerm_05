`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FuvaurpWyIuKKMV+DQUzjzY/dGvp22KyV0lRWw+wII89IIFb2tjcpYC5apGD2d42
1lEjmfjzp7A29EjpksgL/S50zl4zCFGnn3jKrmhZzBWbV1m6oKMmqQDEnVp8Pr3t
8HIYdWpQJfXPO+bCIw5jbeR6Cir1a5LXhPoFEGpWBozrLUIrC399ufN2ubnnHcDq
3taJBXzEEC7oyvRI3Tg1G9UigsN2vKNJzeF6CZ6ZYLXA+Qi22uGYTmwhWSpnvImP
YV8wzmSvzwrVfESq0LCwig==
`protect END_PROTECTED
