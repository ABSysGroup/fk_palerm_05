`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tXR79JwMiJGKkXEMiLt1EWKAs5ANTePvH/MIJdOBToZbHyQgwCPgNY4SYpZFkn7u
zmW6e6lW5pF+HPycTyrfsbEcpbof/2aUktn0m+YjrWFP0BpFXafcP833dwAPbbow
CGMiycL5G4PuK78tjtK9RATx94seXPyyIUSlB3H15Pcc0nEBCjCWxXbVL1LsYmnx
LoqjCffJfMwg4xAmGjLHgXVrKPOPTw5OylLE6D2C+GmZ7eBu7KtGmGNfR7GOmGkb
uWulwH+eHP9puOQwiLuHUSyZUddn5OYSjO1SO68pnAPwisCINvKz+RF5swGOcvot
DjwPCwnsa/xbSfEvcxfCEkZbFzJ4L/iDF3yMW1GhRfZvSsm1zRYu2JqkiC82G6PN
dz9GMTsChF3txoTmJER2LkUVFui/BuFkllVK4vKWQx3NSidK6DWfOOvF5pKamrUh
KX5uI8UITEFxCjlJgti1NmdWCbhcarZ+vvMj1n8feOLxAUljlAGnp5gmQaQS8tNl
xfAKP4JsgzAaYrTKkyXciXCJ/STAbRQJG0CnMnN0XHdXQ1yIx7VA3bcRYFsSuUAB
YsJ449s7tYcBEITzDexOPLl+yms1woPvWlZ7OP6AGQ4vqN7Ev2wNHx/s3YztOzxP
Aqw+12hIhZ7Jm07RSJm5zHEoeG04SmpiwqYYxHmn0rKBSFWee3VoSEfPQBOsI3as
oiEdb2DphSq7KAtkmwws2CDLa6azsxECu/hbVa7eGXrSa43xtDJvPjoCpWnGKBZe
sK/YJkW34YKaua15FWQQcztUVPtwWG8KF6ZLqLWVfUmqdxhjhsFNuiDnRbhtRS1c
15xLgBfDN5Cki/BYSpFSJtq4WHW+ZBgWm3V3YMMghlwYTRjqPb3t4Qii2UBs4j8/
Z9a5bZpG6/vthoo1IhgbM7kF3Tt5P5Mbw3sjkkm1ajWLcI4tqkj1W3rWBSJD+Omc
ugySLzK9zs4h1eyEMfICH5vZRhJbK8cQ34/UNa8/FbmW4VSdDmg3NbDHle0zUe7X
PaxFkHh7OXblXQ4L/+/kEsDPosX8n565Wqh98zusYFhNyx02nrqz21f4bEU8cFC4
hT0FPuVxEKO75/mDTKBOw3GNHK/bCZcVJ3WcRNApmnNikHsmnl9oMM3HFmVYs+TL
gz+TVPuv6N6KcFy/3+CAqax/ob220LpuUbHnrPzNViOIszGgatmkgA7yyD58cjr7
3x5KBM0B+Vam9KwrJ+zsdTN1Ge3EqUQY/K1Vyf+A1qOn59zgOqNZxY1vKseBnK0o
MHczsnda1eGv5bzQtMzobK5W1mM1zsSUbP0UxUcgrjojXYIkPzbNgRAh+InR9Rrp
tipUargn7l4WVFI/7OSkdTBJbAiun9plKHwhbU0qSLy39jz6vL67oJhynl1spPo9
H0hpVnBtc/OuVWx2z00Tio/PhP1CNagWoodiZEmrCzyuZUKmnw0rC/9fMi+P8MP1
A9O3xXZAJdvQb4hEnlaS4AnjtXa3DwgyktGN32r79x4bmrbYxAh/vQg7hq9Kork3
B5q6hU1oW9U3I3UENsRsgUEo4Z3kka3Ero4A2Cb40vcaHm/5rR0kyZKE7xdpz/EG
bsxrv3O2fMFW3BdQyL7WBJfoOSeaNI3gzLTPaLRQqcac+asTHRnjAtBKE1grM1OC
Z//xH5dMdlJVFDzVgM6fI5dhejgaxa7Wa6zwaM0OXI+3Yh/SD+1y7H3Enqfqyskx
wyrvtG4R/Eyf4c5+xsjGSdAPKWOkFPDU/dVt/oF2k5pkZWV+9vrkmrM/+fiso+Mh
YP0RqYa7pSEWnt3Kx40dqxCLXuCz/x7zjOR/3HHXivGiNj0shwxyWZ4GpUliAIcf
AQREvmEhrZER/ZUxpgU5j62eeAJCh6jGHWcQsCE88HaP00vbcUzuds9CeS8T7TIh
xZ2NWwk93j95sBC+2qiTsCMnokjcGVw+EEX1v/SqKqzqFMKHL/knoTSLur3bwrgA
50AMuVazL3xhPPPkId6+1oQA0hzjd+g+9bZkUZWqhuYAxbj/gmmBv7zj18bMtW9N
uKJgJimXlztyqrdQuiKVUdnPvVGXM8CrHiQI1Fq7JPSB3qnFRqQPrFvr4xZ2FLfq
m4BVPk3eM0eCutVYI4nCaKgATdiENaGFQwVii3hxWoKUu84zCfTHZZqNfHzFhhof
sVPsyYZKD9pmVdX8kyKMIYx6IMgTeNNk3Y177de5ZEdPLb9TkLshCGNO0vmwUamN
2Gv15K7SDPBq7xXKeivIOi2EkmphdsNcWEXWm1BkqCRIL2wTADhYibPtQwKCVxlC
g9xzpw3reLKTVmkZSPCcU5YaBmtQSweZF2ZVqgV/aZzi7xwHwIAN80k7TafwrXNc
LVpFs6i8C+T+4pfyp7pqnU7Q8rlkLXtFNIDUpofzJpW+W8g2uedhSC4V6BAH6+YD
BmXqncGyvzrvZ6RKj0+d/AEJgh3I4K0YtnEJluJ6yE8qa/88qkwDccTdHCooDZ7+
MDB42scd99+QXSG+WemqKYRlJJcklGrPVQUPY9TIDHXZ9fW84QWKZKNJ9LEn0rC4
XYMUM0ELiQ9PUxd2fkfdWT2dakcFKZXCkSXgOJpns3AExPpd+sMhYJsOQXK4hZ+4
6PwgpFI7h1QRmY3eakFvF7LkZ2sJd5rdXrAJouV/Yzylv85tU+L9XyWePCGkRTT/
K0t4fspZ0T0ya6+5veGjLSAIAHLdvyaolIQ/VjvCV7MxaeIRHX4RUlecckqbezB3
yk4bn9M6cKqshAKJGKWTatDvyptU7ziUYRhIi1wazcGrat7dwWadYbL/drPcCwKJ
zYItoupJ1cP/riSGGmcwPmNStabOYFMrQAM/xYd3E49dtt94eBwV+IDVIyb498cZ
hj6FLYrzHur7WVtA3qMKrKGvtWWpi1IQzMhO/2XjGxJpS/Nl4WYy591dbGzRnxHC
z3GKBciDx8mvqLN8a4PdBXfdgiJMZKhe+y4lIOTEOObbHbeWbqVfQZtRoAUa8Sv5
qzRX56GI6tj5/eTVZuUSRabGWC7giN8U3tKcLgvtGf8rGAGfQwaNjlNKTu8K8fcv
bNP6oqqlHn0i+Fv2EwKbcPsuiNkpDBOme3bTALgUsxo=
`protect END_PROTECTED
