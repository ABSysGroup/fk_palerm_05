`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VZquuiymqmYmnWbKtAqbZnnQnn+D5P2v0n/+Z/jH5z+PNiYmJJggShHjxajUqNOH
1bxo02VlPp05jCATWfCcM8ywSQynCHQrbDECihQOzCMLbPAvWa/4/SwiBT3XUFKX
baOXeLdYSfcxf8i8DOPl7es+gJMXsPKJL5kVj6TeA4TGa9Y1eVuXOUIHY7Ub+f1x
qnCeA11LC5q/TpjSSztDu2xJ+WYgfLqSVlv1Yui1NeYrTIkQEUAzTCro52b208o3
0jTQibGcFU/LwReZkoezhIhYT2bBivNoUSXEp8PlFnubJAVQewMtrETD/d+rxMgg
76/isRiboTTgCVSGLxU9O5hof82y4zbIs6xfN33hIWiox2jKHHvHX2IfYrz0ZJvS
1++mL+95G/z8tgCcZ6N58SdYt69neB0jYmTCXnXsapYjEyGDo5nGQILFPQ3mSNlL
1TnGi3UKQcNLws4r0rpQ+tdNlF+l0HK44Y75QdeE6s9Jq7JTPd0yYsDoH5voqfGe
1Plx/Ms9MB93SGNPfIhykHih/xM4JlvdKHMnTwphNVnI4i57DT6o03zfTj61qqTy
Z9IqA5LrnzjqYJO8r2yzbWj8jWwINF0HpeZX8hsgxn0BQjWj0RpG4NLqb2vHSsFa
/OIOiwaX+i+yKkRIo4wvYeY7IomLnpZUNImI2mCpMXlOX8OvkDbJuVox+sSHqPnf
TPobxSauAzaFOJGj3uYeNb20kH1ID+emyIlVt4RDWIFjtF9RLpJT+PX/XsxCd6eE
SmcJltxf6MpOH1jtKQhqfHjY+Za0DF+VwANzfRzM0YHyKoKty4ZvNkGMiIpe0PMd
mBJTfrEDjsK/DpWDeILjk38ORYt8njd37BBzycSou8ep1Ny8C6Bz7zzw92l9umGX
vgc1OECanEa9lB5hJoDDj8R1K8BGNWzgEg/0ACJv4DhydSQwLPXIocXB/7SO4oAm
u7Yt9Y+fM+qQMIBnht1RY/5z+qCUkQ5GoRYYB+I8EYzELR8RqDikD7pQXAnLFfBD
8Bn7CneYPnh3gWZR6qwHgHtzELMGL3eSTqfHkJ9LMfnT1KrpeoZ+f6EMNlcw6BCy
lqZqtpcll2ar2xzt+NooG/Ox7PiLPmeBdJFDu8fwFbRa6dSfIX3GEtJPPSM5ucVL
J1lyLeRUsJsKnbRIJ0LwQSwpgXIaCyeZy3I4tRDh4PJUjuwNDY2WSWDXHkICc+Zx
iGZkyfS4UadDWpahTH//fjAI7bp9p1Izt5FJxYdAVVBf1OBRsgi1dNzeww9nvL9k
LKgPwf1OVEuw8+RocV80oNnRVQYp2Y77O/YsI0F4x/vVHnlXmR2mVi0Medo9b5sK
/eLz34gzNlCKAamgOsTJh5F5th+yyB2WjZReNg9fMZELMkUCcIHviMIRq/YKA95l
IPxolRUIYwxz7FeGTDrA5SHBLEY1i6HxKipxMmbtBTGmvkPYWeC0BBHAVq0b7ux3
F1/ilXzLGjfJKlWtExK91NR8Ppl4E4mOdWKkdchgSz/KsYrvCnvbT5svoPgPLhkt
vgqGrGnwzI0Fa3iwqCqU/5ozmJ+h544/XrnNCQdgsHqF1961U/ouzkOi60hS+6te
xo0JkJ5S3ptuTtxjVPw6yW4ieNzJZz7GbgSnYgvavswcYNTmohD6sr/+T/iA/f3/
j9EHrVXvS1RQABaBh1Yd/A1hR8s4A/6i1EpGdb0DNs+YKrPEg63u+wjBmGQEHZsm
HiGgkmNfFnJaNzDP3I8vhr+JfqHGstAWI97O8z66QAd0vn8DWa3XTZHzHlioU/7q
EhWAkG9riTs9VeBxfptBIdatUxFL9ma7QKguSkLDxrIXw0hA01VqY0Ae5NnH2JP/
eYgLF4o05PBWcwEWbLuNNzlZ11l6rhF08mGLejWnrsYz/MtvOg/G0CGu5+pUMQLq
1FaPHjwAuF3qPdYIDzySCPfi/ozrGhUvBtNBmtzVP5er+wQ8KpK/FdOSmfhZqBwC
5/MVGdj4kqV9NgSky4ctPWvC63GK2dKMIegFFpDhs4DC37wtjKEk9kvDm7FXCevn
h7gbtPhNRDbU7tkc8eLBwPmxzRvVuJwJLM6FVcbgf8GuzP4YzzidkfreWIOwliqb
aUSWyZXSqDX3nNRL4hxPQDBklPx8vfJ8/D3f/yUPzWt73TdNzmU8DlFK8l4nbN3k
MdkUMifuyl8g2w9jQtE3MYGBI2boNnFYdmrQJUgKjM0OaVFAiL3HTBnVLcdngPE9
Il4Xzey6qimBHeMgeCwZsRpBCsL9SLikMW4Y+cq8VsCbWPPL3BnaXO1wcMtAIDTk
605aIWacIhWFtI+hrpuBpgKWtOkW9VVeJwOZqYItr8g=
`protect END_PROTECTED
