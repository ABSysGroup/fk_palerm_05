`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NjVdLWrxdw4o1fdKhiO6VKdfwiZzKjyyVMS+t4UhFWV059XwS9uohXcJA+vNmKFd
xzSCAo+ptvzQWwVIQySe0TBPS/pbcF315dCG3kiA+aRXxKIHu7Hc4sl1K4g1FHtE
XLGdjprgerXzh6rfCpFC4RNRAokdjEaYnecwkXDhiPtcSxLtb/JLvlsOJ+duUYYm
6zqlBdZEmgBwZPrHyOi/HYPEYRroUIbVfbcPJIEED5ihYc3xsVUtSz3/tB4nlpBf
pNs1f2J0IGDanKu7Z3Un9HAI/YOqafvku6+yFZ+2QEnikpDULv+gyBenhAubgaS6
ZKUzCOW/NuIonFEM7p9Da3K4qLdIh6e64sdha50RzaJ4sQZPOgXZNj15bLQGaegK
uERf1qlQoSJHqQ+xweKXiHhRkcyyIpE9Fstr0Ybh6fZyFS85Z8e1I4vo9I7PK9VO
`protect END_PROTECTED
