`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bLsd0gcl8P5X8fB1QiWYmrnxNAL/z2hbhf58SGK3Ku/M44ys1bl1dR/ZzpkazYP6
zJv+yK4VSjhMAgDBe2tO9ASFdxvsnD4segFxqTQ5ZsExRXhvkB291zuHia+lC5RU
js90+8HoO90kgxbooqvc+lVRET+bvwCqZj5vTw9OPlmH0drxwKC+oN+Doz6pbR5B
WZo+fpQr8EDPritEvFdk0F7gvPa0Dwo72DpFYWjQ+j0T2gTBMXqhMNQFob9EtAmf
1P2EyNqmfa3L5ROJ1IMIOr3YVJEZ+8Xo3orISIlOmEDXjxjfGob+W4jMxsV7LQdn
s+X5D37PEuRVcI4IBuB8xkdKThGfGvSwNJEd3ExfrVTToHda+LtIM3OClukGw1Xc
l3THWwvxeAnsp8+laMgOZDxfM6V5ocHnXyjnlDrETgikhZ+vCuXa6M54+PmH7eTc
3O1r/ZfqTP+yP3qy80IC9JULKBmDC74yp82fhXCGhSUaFh71jQUIQpkh2JmQihHl
mAg65GGwlwK4DPBjPrWDaD9YIyyF/llsxAVNO6kvh/x3dqIFnInw06Lu6jr8pkMR
n3SFiIQT0073HuYJJHkU25qjF9xE65jFyHEgBQszjywI4XmmQiLgv0Iuvu8CVYaB
ro8kHCiewgWHhkF7hoeIJVJg8zTLPU4Dij5XBjVKqMfJajoVKwR7ou8vGRBMjYWb
y0mwRzGWn7YyTNXaMpyIeypb/ZBVDVO2c1kS8QFFPVuaHnf06AOfLghI2mmv3YXV
z6Woh1rCKTiEvNHiODSJ8i4nrfNcg5EkfeptJVUVGv9W2tqGa9baYY3quzcLgvM7
09Ldwo5Ocb1drYwgcTd5P1dfqv+L0o04RMYyErKOjc5aVqrB8MgpN146WB+wLjsh
wwRpES9A/rbq62nsDvRmKbjO8r7T+FaURBU1/HBnYI6pucelEf1FBypq3Sl2mySt
NklZZOttH6bndhTMMfco/ghmhU2OM7n98Nnu4bZD6+dwv0cL7NPSBdR9dMb5tf4n
wezvn1wVCCxPPxxlgSSESQA9cIUuCV6ahb2ucIYSjcMiGyieWWheDf0RU1ZBpYT8
R2tBKf8trxel5BNWqUZ+Bx2Q/cScM0r66hSV2wbnGP7ek6Idi6M3bshbdVr0xWYv
ADCtSneYa5HJ7rTsvDziprs9JkSqaqXR3aGBYLWYKmjv34aAGR4G/tHyuhhNExXy
BKS5MOU5cbvQDj74iwWUtuSZb+N5N7/7IQF2aW3mDyUnJVIQRcDHkrWfh7MzawM5
/QKEfhZkXFQdLXp6YxqAbzA3bBBQO0TxPusckNv4B/00JG9XoimyoFxPC4O7+84j
4N9E0lVGdMNdC2EWn0kja3C4K/oeyr4FAabCyE4P+XtZKjiPB/ukZHmHGlAsBRDR
KVODrUei+6c1N6blG92ng6uLoPGzj/2cwFMxoP2mrszV85PK9YhsKStqEWN/EpsL
MgWiz0q90Np7I7B8Xb2zYbHXDzYb+M+oNQBVIwYWSagdah1SOotlBWRdy1eJLhA/
gm5s1NI82ypk1pTvUkoBsId6+YlksDX42BtkUd3cjzYa9EoCPUWzjVuiLP/8ZZFD
uIgavQyHh5w9kJ6lxMGByCp2hIOENj0yMCP84JnUzshtrWVz2vMWmvMVK8Dlp+6W
hY4nPc1Ja+U22udgEnLF75jv1tT+H+8ry/Qg5EhGqdNjuA6nmWTAHudlZ/+DZy/V
GFh9EZKI8EEEuypJZH/hjkE0AsrFkDEvT9fEHtB6c++CrO4o6p2RO0F0XXV+XJfc
e2Z6F+vvxt3ppuLIgzNdj2310rCqC++naS75SWReSTxv+P19bXGYPvEAih2qQFta
iZgPXSz5J7sKWTaM1I2EZG23Hg3YceMhdWPKDdVUKis67o5Tdm7t3jNU8SHiZk+H
`protect END_PROTECTED
