`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FuK6TfHJAXY+CxpKaS2BQT6WTySdMMEhYVtmgcFefaToljsFR8EL2etg2h6sZE8E
v7gZB6sWrdeXoyGuatrBHYniAsJhoGHAljEignMM81wBezO+sgy0PLjArEZb3VQk
AtH+Dog69n/u3vbrMw9cqCz2a3zaaElLk0z8aiAQJ2pMvDjFycSXF0vIRfAgtnaL
Dfxvl/89hWDgoHUqtZJSzjqllPiM07wbqrW2VuYG1GEj1XsiUtuE4MFMMa3nDx9u
iRuQV1zn9NibFeJW7uEDXuu1brGl/1ZJGT68zr3I249JBhwCa8OWx8qHrOu+HSVj
djIbNeknPvULoshGrywgg5Zq3FjrHapXsmpjIeB871e5fNobAREm5Y+5PRbSHRsu
NtJeCbcmE9zg89WE+V0sLTJrt8tocv21MFQa8FxvNYsRTEW1CuhAwktk96LpwDQh
dEpA19/vliC0kW/AdsWs4Koedqx6sFilClNmzRgqBAkeh9kzwdUDMYAI0e4adZDG
e2j+j42EypFWJj8pzD3QslLnRvF/Uj8zAGjLYE5vFwh5N0bq7/oU5SYQ3sUIl+bv
l9bnaK8r7URy+c29KCGEe83O6nqxSO+eEqPBsYYbys4=
`protect END_PROTECTED
