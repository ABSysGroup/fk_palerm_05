`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c4sMmIb/WXZ0RJYXXQjaQO4MMwocJy6qc5B4Jmoi98vQyQ046HJqONNHh2altrea
5s8D0A3yY8+CTUz/foPdumy8tE/xOPpKUI7A2gntFpyr4JUS9NWE3dTt6mvUflqs
LcV1+pVoDtGS/rE9zD/5oyY7DsmAnQLjVX1C2WHncLzJf0lDiUik1NduwmHB+MBJ
4SA6mhy1jKLe6z30CcwtupvCGPg1FDr7p2fMWJqSPHZ25Oe/eynK84fWDlyBP5A3
`protect END_PROTECTED
