`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ut4F+VNN38V7L2hHuaNQ5sfT/ScrO/jqZTAS5DJ4C0IxnEfqK5KTQZB21W8LClFX
wbSjld90hlySgVI1YwAMeKbdweGv6vzqsjXcv4luIYO/MtWDI8lP5ynvKTFUa+TJ
KRDTuJjg7Qxa7M1TqUIMLyg4+Bwt5xx1mgMAR2pjCPHsQ4Rq2fCDwflCz62VZPyA
fH9jVFRlVf+F+uZMTkAFzg0yqNKHicqGiZYvcIfbMPNZ/jUzt3o+6Ts9obf6Fni0
nZteO+ffYG/36iIGplKqKJHRbHLyFxaXcJABRH4DOcnwXzNcwmrns4LSC9mJCNyr
/TFB01tvTjmYd+lPufL4lsvP5VjTi3dJAML727+W4wPhQWgX+zhhT8dwl12dIECC
OgrGxnK3PZIqzf+U7wOdAIy0t5Y36nGL1oMo14JvwNQhmGNp1oEr3CdCmUAH0Td3
4gOa5DkbBT4EZRv6ccHxv8uPBKW4x8LHJmOg0APTJhVTjSac2JajYmmbZC/pTVoe
8LQUbvID+PqR0qNN9+B7kSO0ZeGMOMRa46X1HDjN9HXaSe4VbmIk9XCODpTUG2t4
lhBxAsB3fZPY2QuggZUncwS9Jn/dbpTCCAp4t+YzfamsGEnWQXGJ035E9TEBYkQr
inact0Gw39Tf9x/w9yto0IGRYI3WE5vyFfyDeIr5cLigoOpw1tYRlO2BtBFdXU0U
KCUtAtNKTSRKGOYINvwAT65AB5sGPivLkYwxHax+tRZbeUFiUjbgFbek2M4g3iMK
uhQqqF17Cb1puCHLyYlgyhRod1yDaLuZWZ37Xtnd8J2rtGpC7FDCO7vX0B7cZ+m5
K3elqljuyOouUdWfqvmC48KmNKsiHzVbS45WB3L5WaIYYYpmiZ2wjva4/OFCQwSN
FpJUfAW9u6VcNgc5P9QWNEFtj3yYKV2wiRugRdyvN9zrNBNi5yFn2wSI9bdK/UXW
`protect END_PROTECTED
