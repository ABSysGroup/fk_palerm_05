`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZGgr2bTgKffzj4UyMNMLwd1Ab+vIdwLJ5+DmXmGN3SN8opIQ2rKL0MGumON+FtnI
UIfugKiCAo34HMk2uDeUmo9azLQ8S+jdBIDndHNDgN05J2kTktXOtRedUJGIa77w
18pTNF397FgxnKZkoMfOpo8oO098yZWrWJoI3s3Z/nBhMwVNjLw/INPJ3evWoVe6
ZrvWrU27pQgEd2rPI38P/RbkKHgCdAROgQL17CXxHYgxKjeSSP+j+J0y11vouZSx
nksIJjqsfPAeniWiTHPKylX53LXuA9IP3r4YYAaGsCUf1Ea4q1eZiMWe0ZG50mrN
owGf4AMe3Cq+yETEmngg0PKphSw2pykLztNccBGN4Os3rn3LZ8jlLY8qMqvN9caM
6v7J/K7/FPx0HVvMzpaBErh3QyMGD1c828jUBUyGksM2Ol+1sJ8aNxWC2HBiMj/B
zAFxLEp42i6eSDCyV28YSd/fpbc0E/fc2Grd63ep2Zm5zZqwCGosyCOJYPPsAtkw
8ML5eV6hrfl/hmZJboO+iye+8s2orSVGUCf911Bi1q4OwkC8fWMAOHpfqJxBfcaN
N3p5hNHcDoKXfNxsjiitTJmOIZeqIQ6VHUUbSKXmNlmz9rslQ8q2AVjofHg4nHqv
WiItMrXyNCHPLAp6OIoaBX0RsqcEENU0JJrz7VoFM+m8gkMM4RYiQ5OtjIZOO3hY
woISGh02cxZyYNUEciVz0zL1lc60Fx/wyaDUdPu4kH1OqiyKEDSbKwNYKp0J+pDJ
uXAuszpjS7Iw0utO3KLa2h6O8jSaQtIxK/XK9zrTWBFEkatGubUpdJcCkkVUS1ky
IPAXFCVltgZuxBBroPWEOmvBjvV4GN2itNXlxuSz9tBSO7Drq3JC7HFxyQUV/gyu
XYZvxYqHXeXplfBzlH8W8lJpiW8QYkNrqR2vZLZsApOvjw5Cldi6Wb3m4E4a7Kz6
`protect END_PROTECTED
