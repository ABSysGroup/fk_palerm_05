`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bcNdeMUtznQ2wZQ9910E04M96NA5UNFkMkUDp/VcGZ1KwiqPvhVzsr/QI8lrclEn
CyghVp2isPRfOp0VR7CcDgfVxV6m44sn6Dpy13KIjMBa92s1OoyxR1ufTyn3LCGG
RhurG/A3TCqczpB5XQJiboTye/XrOMNbkApnIp8ZiLH1iJLvfuosiq4lYurMF8Oo
WdFO0qHgPtOr1NWPTxbzybVD3hqX1msDLyyPgDWi+GNC+hVyQSBmzRcKwDapf9Ty
ZdBHYZ/G4Jod+h15x13Z2urA197wgUSFSalmHA48jh5yQr9NacdR6qig9+onrRn+
s0okyltazthicBoRlyXt0By79I74T3ZPHs+vVslMS1teBKRWzvCL/YdEQ8VfLFRB
oDPWxDLXrAPBsGjb9zcNpbpmvr3jB8SJB/6/OG1ac4g=
`protect END_PROTECTED
