`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bkkvbZhS9R07gXUjxl2WJvR7R6QURJldS2NzNjEXu/Dw4txjIubGzJLqdgmliz4I
1IrkFjaXNzWBsxKfgaK/5iBsvx3VhVsXvD/3D1KoZTO3V69VHeqtGw8V6+FeA8OW
LlKJGdQdunGdtfzp1Bxjnp5pqW07/Fczgchx78DTwoNmAuCASQCRsp+grilYvt4j
d2qWZLXNKfmjxTgTkbsxnJsUjqRIE5PwoYnJzqJkuqu/DlCgvyTy/fiZ20nrfU4/
vgzDi1ExUGHiz2pS98L76Jeg7VgaZbTjRv/eB7bjgN4i/O9JpEYhF9+wCAU1LtBs
9xlbYFcZIH90xgH8ciaGudzpPEwO7s94FTmBebJwUhBoE8S3Im5A9rtc/4DSEkgX
zerqyII0pbgiIkwl2bCF09RS0QT51vKqmjaTaEjt+1Lmk7fHw72EgX6lDVShLvX/
AVrFYiRSE6r/XqH/wHpuLj5YKtslMnWwTv2Q17fKuEvoodVL99gGX62uzqe99M5e
miIRV2C2xJppSxUouikj2u6Dd/cWs0cLQZ7HqZ4IhCk6X7N4AMIBvGSuh/yH0Wr9
3fyPd2uATYZKJndssoy9dDy7/ba3Uv4xVuKA9CfdpK6CXDr5VUmYbP5nzkYNf1A2
niWr+DCWYohm4EBhKzNVkC9fM0nUjvjcKgBfLqirk/uAE41xQhizxZf728VbtD0O
Dbl4GZsyzFkvzHXCtmKPeiUmqu/UIJvdu0B2upusGiG8vgBeFVkb2U5f//7f5ZYZ
pYKkTL6yWHMDX3CgrWjGXdpDwnWuoCK53L4ytafUlg+aGSBKQOFhmxR0XagYsxGF
Lai4SnNuMgBwWl6fAi3oFlk6R2ksiJXFsqocyj6puWxy/rHubJOa7kHVaCemkzZo
7v2Ojr0lc+RzKS1gLUgd9aUFXumqrEsmrsxyfzXMPmKM5Bqu/Ln3DSWWi4DKWAjj
Tnxot2Es4yrKImzrzTx9xjQID+O+AtBx1Wwvec/74WYTbsTB0cKg/96E4adju11o
3ahSoF3LtDn5tT9RY2n/5w==
`protect END_PROTECTED
