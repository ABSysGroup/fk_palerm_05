`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6x3M+guZ6Ic8DekR0MtRY4OgXl3h98AzGa48xM0y20IWO7M2a/BFXSBu4kfoSx3D
hXbCALRG1QFub998cO+Fa28jk4TVkyNn5VFMRmXQglVnJJvfNcwhbLEkfHHAnQw6
0dsxbqzJKYSJPnoM+Bpr1mBPyqZljo6WijMSdq6bURFVrvbuquA6hmzuWL+ZhQEs
/u4uIBuDdbtTzcIBJ5nQbevcUf98iJ/tpqhLZ7onm2Th3ZDnjHrVWvnaD33MRs0N
OBIoI0F2IkyF09hOy99EF72RGeBpiTetT9hKyTq0waSrLsdVn1ktcsBlIlBwwxf0
7dbq/5ooYJu1TxWUk22HCT3BBpvZ3MVIZMhy45mAazaqqX/TlCSEAJPusy42oJL1
oPQ7jiot6evDWuxH7YTqnj5yRRQq3oJLlXtnRFcqYvWCOccIMJeZPy+FNaxOgwuG
M8Y6iWqdUmlz2jE5efWJEozxzEj+sjFX+vqSqgf/vOwR8m3xWXfRKNpE+RQxXS0g
6cLUWfeL2TbsQm9x6zwF8qUgiWtpUgczQAeyTLKhoG8=
`protect END_PROTECTED
