`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R6NErDU4CtnToNLKHsS+LaUNBsdNSpC+SSLrCqUto7bC1uK2NJ2fm55FQRfChteO
je9IN9IKWm9mX/rtv4xGrAEAJxXFVER8GzqU8K2moFbHRgQSlJrjNVjj+7iYuPFW
bLPlKQ0K6hTdLBYjGkkE1aThqbl0Suf4a2VdyU774o4HZWogSaz+KQRpDNaOWKBs
QVH3jw8fNmropI8VWLhGNHmRBwLxVPU37Bw5ahpEYCl8zxrBKL41NHBfGX3QSDw5
Zebt6gcLfm6hX8tES9pBUzgyI0lHk48nE9p0/iz+qEzeHQg1f11c5eJtGBRKOWre
Rmea0cOEqDmkNC6LwdyFcIZrCrdFzrgGuGEKjeb+C2uPrnWRuHFyWj5RM3ST50ZD
JrO7xdkAr4kiMpotvxX00UtiCD8mMsQ/jo/BIz6xh/PAmcFG/4vAYd5io+h+SzzR
zVVpHIe8b8UbdjqjtZhtBfLIcxzQBZ9wXRn+taxAOfTD8kOJGOFaFDLcrenTVu5l
iK2+I2wRJlj66df81ElZ7bTQSBLJx6V5sCeSWTPu2kj8tluDGBa8zufBL00G/GUj
E/W+ZROi4/2KLJ71srshHrlXLSWnd2yBosx7mOQgg8ZuW9V8HoDMIuUtF+MG29h4
fC7JjG2pU2fHaZXLlBCIsQ==
`protect END_PROTECTED
