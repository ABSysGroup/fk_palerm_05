`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iy/ANmjUEQPvpRn+3VJR/iLX9aN6HWOH649hBuvTdZjMXvmuv0T55d4harkk0zKr
WBEpXnHG6vfXODe6TiiJlsAoG+GXRabYWng5ktTF0k+m4sKGLtvgbdXIZHex4uAm
YSdKfKNmX0QTHFiy/24VDIBJlK1/YL/6yp4OjvKWmHy1lmWe3m055hOAwyaH3TmQ
W8UunO0qiNa9Gy3IaSxKMXYBVYjsZ1uO7Vay7hUU2J2I229xV2CclQqjSJH/cvlw
De5MhvmwsnOBYuvDax0+Pg==
`protect END_PROTECTED
