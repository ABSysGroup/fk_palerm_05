`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
krF4xRsamQQdcsGmc1+o3Ih+1MlJZlW0VU4O9xuffAwiIW/DBnyChU4Ap420xepf
FXuEaLqNlnp3wHKKG1SBmyRmJhJorpht4KoWpWohBGBiRiG1XOHMDvGzX9ZKbASG
Ce65vS27dA32aLlRwSPzdC+zxF6MR88K3zvJ013SwePxpdFKTjpibkvkK0YqTZ5q
Ii/tj+JcUvXOolYWN878QRFUR2Cjeo9WTEADuskkgahhsMN2PcWmZogBDsi8Pcd+
0gW/iQ45AXm4EoqFkJe1OWhSM95sou6T9YeyqXPdoapy5U0y7ibl3i6cIMW5MSFq
13pSGgOXDiv71dSBHKRUsD9lKNHA6n7nfy5ARpwAakFuqwX505lqWxKrsBVjVdYE
G1sdVqOjkxcEkwXluJ4jl9YMU0X5axPeR1+Auu2Y6LkGCcKYoqLH9+ZbXD90cm6v
9eS62i5vDBS2N5K1h1uPONMmF8erapqFKXavSHaKYVGRLY8+ZISFaDL1BqEJbLvU
4BbspIZW1LnFLPEaTRHWDXhU4rBiWHrXNozRdWwdEEKMe8pg60zl01amcFx0k8wb
aWCKFubg5BwDZlzuNElvH8QbSLwgpopHnmuiLmsO0E9pzhdWm1Xw1QS+3D2mUi31
STNMoT/0PBRo1GYzOkM9SkYyuIBUHiuMxoSROwl3LlKLU0djs5Gi285ayk1+4Nb4
ShZH2QfOvt43JSC5zG9me7r85WRiPck6MkEwTVAkkIpUFrZi4X2AlaKt4ZQPceg6
vxH1AACJWcaz80MzIN8pgrbW+w90UGRDxl7ApD2I5B4Ql4ujGiDe7R5rHonsf9mR
0n0wSbOw5Sc6z0EtoLE9nPnzzwU3okTJJbjHBG8rLu1USxlu+5beX9CasqUpU1Pt
VkMIROuwalstfGAyxM5+geHSyJlTzu1blxrhEmOo6M/fug4EF6rPpruk+8sP1Yk6
3f9CVrvobgWeYuggXCn2f+gQm4Soj9pubUrohCuiHOGzQ+DcNLvAmxORXJAQ4hHE
AzRK6DourpNkSqnfEqNx7PeV/wY1K4+xgNIFcvnIVsH11w7xBurGMTujOaIhK/5x
kHzNopdZY161LtK+DiaoWLcuk/nodl8RR40NyqjSy+z8hmH6EsZDEHMeOdIvAKya
0dTnZUDU5LBKmXuPEDy/fyyRPAt9OATmD9DSyzZWU2asLXgy3BX/BjUjKJfl10Sq
/Lu5TdEXgpmm64PEnTx/huRsbEEIz58Q+na8a9U2Nn9qKEv7bYSjYdcvk+BkrVd/
V4IeUQUpbPjYdpH8C1d/3Pw8SDCIHZpw16W2GPIniS096ziHnV1f1rFlR/Z+4OTR
kh9XsscQgjf5wDw6O/gsXdzES6rMXQShLthJlt0CeCvR9cvi4DiA629CkScVBu4S
aJ9YjD+g5T2xuu334/OsOfQkpQNyJl56V+M6JKVUsBQn/0mwwnzPNfSfNVXz/Sln
kqiIoMv9sJ1Yz2xb7ccM/8Nc/Kz8gkbJ+2FitGqVq3lVF5RZC/baBLaJkbYKP0qy
hhvb0Lt35iH9DmfDQF+MUFGoPWQUdutASipVe/GS7RiJ85Vxwk1YD2hRFnp+ymSs
Ba8l8EhDxTsanNvxizqzfeRZJ2zLAE/nNFf5kFB+M2DFs2I0YN//d3TozZuPwAky
hTkUAeIbv7525CPoHYbR05TlcUI2pjXM4O6bwGIya1k=
`protect END_PROTECTED
