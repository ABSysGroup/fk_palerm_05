`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hUpEPe8ygrGwFiv8DxcJR7vLgZ84Hw4IeAXk0SxIjhPJ85S/6oc3H0c9v4IJdOSz
U8GB9LuZLr0feuGp/lKIvOfA53Nfv9uWA6BGUADlcjwHpXYFCt1vlKHqoOf+1ZGk
RzOn4GkaOyGteH9hyfLzCBO77ukuJHk6akwZdZ7iR64i/JpkEgkJ7QjjWkNhUPB5
aK/nN6odVNofMD+/cpp4Wmz2UhVKse9oExUleKjd6KeXnEsIL0nRnK8GewMFs4Ez
ISdKT38Gw3zIH9iXU3+S5gB8BA32AWMWsJxEy3+x+t1Ioad1sx3ukOFlYbfPGssG
ewy8tRyayqzOcbwtim7uF8m7lvZjf6RhW1YIPyutLjN8PRksG6DoIfSZjXU+xSd4
yKzfe/92y6GdW6swB+2yjTbCHMbCF1KA2qAKIvJ5OK8jh9YL5fIObv3fGBc2QcQG
XUtj0JRog9zyBI1AA5TiiTkEkOjYbxUhX15MS9SIUVTLIIp/OVxnt1mlq7JYBZ/C
7/9nt0fHt+449h9b4GEfw1uHzAmih1gsfHtpwuuDPgtss9QLsgk76q/kFYsC4+ZP
XT7fuNjNOC+Bk0YiwXUHs0w7It0hncCyouVZRVSwmz/oqP73iS2HofUwMGcMBKrB
FxgwWv9h6Vbh5zNIzqmMiXI6R+r7pcyvk+5PHdnMJ8ddyi4yZzzoosMjPfrvz3KU
z1vBF7d2zzdwV0llCW3+vgJly+aDLKaUMI8cCka+YgI0Z1J/Gwngb+TEJ9LxRTWo
0Dj1gdA+bdXSpVzDXQfeWFxrVx/kLPKmVWGzKCC/j6pQZkoF4ShDbq2aAn6baXlC
lmuMAQkMJGVYsIj0mMrQLz68P8E/3ctjLY+9oYdKZcO8drvSCxNr2MYkWP0ewFau
ko29UHlI4zAsENM1nOAp8R9Rv1gH+pvtEGAd/boNMf0JepquEDWRv3hAL6t1BO3V
LX5S5YwA3lPGl72lObTQWQWIWN6PhsKv4hQ/GkefWxG/QVDksVH7YN1VCBDthA4c
l/xfVQMiMdSePSErxQSpk+G6btuHZ8uhI6jcxkMLLDWQZV5vck494Bz8P4RScG30
YldV3W1T/CgiJxQhQFfgoLuLEgwdg3SCPG04gMDr2a61DKf5L+PzTp3bG1bVybiH
LFRVFHBwhYA2uqjeJhdGAVW9b0DnHuOcYv3LnhybuuxFrf5eKiRHd42mgwmVj8VJ
zqYN0JUUlj2YD28uxej+9Gh18wHLLul58BqbicN8yU56IH+kBR2qUyCdJz3LuaXv
zlpW1iGms4wMxq0UGXXaoqCJAbaLmFaY/C3hCu0Cev20iHQH7UC+kgI4con0a2Mq
ci+tyIKLwuLPAm53y+621eXcXRYU5yjEMnXBWwyOi8/gcnK/ecUTDsBZYIa+KpqD
hqbm8apNfd/3CF67trsQcwTcRjZqIKQH+W7qmCeKftq3xHxE3kuduV1fIPqigaJQ
drXrlObW1CXoFkobCTlIYolJ2ihx93aLcr3HrQ95C9emDC6PTgjZN7zhPUBnY5px
hOkuedypa1bOu6tD6ANUNKIuGdtSt31N4SJiUCYqFa/Zd5A4SjugDQiVjRaKbRjo
eQp5WetymkP37v8VjfE9dffoST8Q+t0u/JuqWNGp23QNyUwbfH0YxGgGPlwb/dQY
Hb9s8JJbqgEXs7tYEPDOgBx2nHs8oREOudLTCJQDfE58lJiiaYn+06D+W4aYyB/g
Kbaw1kSIGcOtbzLF+SyzzFFx0Xb+kJUElpoGxKVBiJB1pmrRarBE7/wBVIK98D/T
DTgcZbhiKCoikVpHnSCqq01zlNoHx5JxH0CCQrbtOyqdbJTn38qFtfpWy1PH9IQo
ocstRH0qw/mKIWKYct7ujif1aNifS/oIWUL0fJT30sIBch3KV2+RGkHcUwfWTEZw
VotJIFk/QVi9ZkisSdUIQkw7ZS8IEm0qj9DkC+jz+Z8JWVO1QQR40xtJeBIpnQQ0
4t9XQRRNT3p6ess3OxKscO5b5W2dCt8LWkmfk+u3c6kGn5X7LMq+2wJSMJlssqEh
DjKK2RvXADcXc7RW9dsUHKC91dGMCuJtzjcYSM+QiDQN9zWr/ZcimyTUf2SvCrjU
9Jn32tgbdmn3h2d4VYY90ph458SOGGIocxzSRmrKpfKSM+ppiQBvBqCkZ033eXuB
Lo3AXIahB5LhtdwHxAxIWyiBIsU5k/ry73pSpVlWHysQmSzOToUlqvArEQgzsqWf
6kWwTOunj9KMHz4BgJFJbsveAhu6lKlUpjZi8QKnycLVX1OCkbdRnl3JzXiWYLtJ
94swIGiobulfKxGn6GVQHQ7xwuI7xaUxSz/GqaPSFa+S/l+ek8cIlf1RbDtDn7IP
dAnYHEOm1jz0Wys3aWlMg1tSC4DgfSoUgjk3KoecnZae1KTgf1soIJJJhCqfl9zd
35Fm4fE/Or/Zf8HKp4eQABccjVqce/Y0qx8Tzw7KzezJnHoreW4ULGmkQnxxlbde
1EoI18fOSvI6yE+okSHCJAj0L9XVZoi+DX4IN1nuHYuJ/mcT3sED8/uWpPclpyJ6
0wP9B5yqlmZDhAC+OZjSB5Hj3HJq9E6Icfbw51H7dghIdP0/q9lye+rvM81wrajW
GPP6T5lMH4gQ/on+rnTDKc5XjdVJ+0hrIfIUdAerztwhMXu1rWdXXYZ4Jvh9Iuk+
GlYrl4HfzNyla3Z2OtnicA==
`protect END_PROTECTED
