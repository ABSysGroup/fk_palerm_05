`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ud3s5r3B56MeiVNLdXItpXkcz+3zJfaHukZl6HhakduJBSm+eo+6vnSIhzws3DK0
+QbGPxDDqyfGO3yACgWLv+iaaPjUBqpxmgMHzD1ZETSyUZ5qD+tPD8V7FfpkUsSz
SzYAf8TJSirpYwj6u1bTAaUBzI+qe/mIWbl0La+OPjBFPSkKgmXiDjG2drujIYKL
5G9UKQY87SQEplK2fA7sjy0A+bRnHZEW9ol+WnxdQTkch7IdAzRccDOkgIU2TfeB
M7/x88mQhC53u9GCGM0kq5XaTTACLdlzhKyEmj57dRxT7KXVfjDVZeUSHKqy+1P8
yQqKZI4Le4y98KTZSe6Sc6RvD3rejlhD+aNCjqGcSWzHVYYSO+1JysRhlT2EGtq0
IForY9jnd5QC3YtrpgDFxtb5oL01KH+niRyYB6/uYjZIE4RKPyRaTjr/uIi0VlB8
pkJym/mxVTpYN+/QP/5m2s5XzQQCGI1cp06hL0ZyWuyXoGhdOJfN4ScHBXwmXbme
rGpWxpnIg6LZ7UuApVq2Y9xLPy7sjB3J7/9E3MiQNL5PpWisHXwP9sBmlnNhgRPe
Q/KXJBYvVfeKJE0/TVohucRfbN8UOczhwnZbrvPm8h1nMLJ/Nu1jpZ7o4caZh/SC
TTrygtNWg14qjBmM4PVwSfzPJHSRPdpWPXfi+7TvQNFa8fmw5d3XLuN/mgaN3mHj
5ZBlYdZ+xEmxzjMcsv7ViUMTPKR9YM39kIXRZj3UOV8uZx63ma72V2+Vn/qDQxDj
5dotEKdMZGABlLsyJ1FS1mrlfVKROq++dT0IUJHhVRf6eHNGEu5AOzhoIxJcOCv0
AJj6i0Pig1y3WwKtG+rraR8BZHbUZFMAs478reVvnrIuXTjVQNfTshrzzFczjTbM
EdzXTbTGLmM9Jr1Q86HdxawJnoV/GIgha49fxyM069oG79cURZOVZilF4+m5GzZ2
65YngXASYViPaj45jQ/B5UbisjjcCLuJXEgVDLNEkBTl3YpXP3ki+hS7wWY6PsM7
sPpnHUzPW9zADxBUbn5xzWSlsiTny2uMI0pCOAUhSOuGtshv/dOKOYchQxuMHmwc
OjQpGaThUSh4jPEEcpocuf5L0dVI3vk3JMaSbefd1eH8HJANMziQBxDgaJNK4Xp9
WpKzv8PQu4xjXPNa9PrjhNhRziHeBBv3LvMcZc9mhVSdlRUJNT6jqUqr3+RnHLsf
d4iDhgOee+OE7mPJJ7TqNulXfbSPXVJa6dDp8JBNVc2M+K6YM0R4Y9uO25jtGU0j
8wDkdRVs3r+ogfvBKo77CYzg3lFNhGMhY5rYOl3OAD5BtJPcQPtYhWerePwB31rm
6e3rR+rWMfQ7/aI1Wb6YHAonLcs6wcStGOId4OXFEj1qWXv52NOoPJERiKitqZFQ
fZExSUzZ/mr9kIHFASeuUgm0PBGiMDS7qjBE5uspaua381nHTRzR1y8l0/Z75lff
ftD3ng6TB7KGp8977DSWY6adKXt69Xzd+/U5udnQQWFnU7q7Ei847fMWf7MZvwBu
drBIwZVoFcXUzkXozymqx5frSpxMU+ol0jtwp7lkcAU6WRVgvzPZaPlU7dXHNopa
NBYg7iAarm6rNl9CCb9N+SJBeGMQosMyj9ROiUxH6zonam+GE3LYvyynSTU8NRuz
bmi4J8aJpKiZjCfFEHiidJU8CQzN9NENpjBi8NrUp2UiJYWMEus7vvGrq89mjM4R
+ImRl5c/swWV6AqrNUBAZpmOR2yCrQu83O+PlDB4woB7KzTVWYsNIK3g/CFWmRkZ
lBuoLzTDIY9BS3T0lrPC1NglaqfiUuNb+16PTXZfPt2ozS/aS/PgTr0umRhdxqJI
F1lo3kaT5QGUfG9j84L8B0QcAaEV4GOKv7kO8TwKSbR6Yxwo46OR0AgkoYfE27gs
RiPPYTdVMIBugH9CLSeWcONQ21JmJnmVc+lRvdRtjSgw+12Q5bis91DOLWP9Z+3h
vWyfLYs58L4K1FDxcvVx0q2m0SDDn4hzMPgAbbEf+2kAqokVfsRqguTbqQ/JWAA7
v8Q5+tUcYiySguxrpMFWb8YPKXfsQEtRwEEMj9yRKTP29fEq04LaZgk4aaxTD1X/
TZurM4wjXR6dQVFpLep5fGtlQ0bFJx7/J6zY6ZFtg7sc8nMJafO/EW7NGimpLyed
X6JJRvDBPp8a2Kg0pYGqMsrfOC6gxQn0ZFI6nKFAuHH5XDPLQ5JWeQE28wXDmktR
eOS5b8tgrAD7J1HAoOx8/DJid6Q0gFItfmloSelFf8Hjie9FkFVBW1V7hyVASvZf
0+2r9DEz48Vb0+e8aQvba3TtZLWuEzviHQvcSMsAgOFc/+gkMA0RkAe/eBD0J7xI
Y3rC5AWtzrcZZ8mgORlnQ1+gG6iKSG78hR6Fj7dQqDA1vAdP4WZa6ngSk0pmZZwA
8u+TJ7bYqIYfVlhdJfNmKVnlnbqJmeR1RR9fSI+u0ar8hqZ29592RMF+q3M0vXVN
YV4I+1Vl8pJddb4Y8drUJgIb4xiOBUPLTtmZGMQ6P6xUyK8rJ9Vg/tnB8se5Gzz7
Cora3Nl+3vhqPAPUCqqlmEqqARAcpHFtdZnybgrBDm4YAij1TDk6A1Eli454H26/
Jp8RxU0HKqhD7sqOH7h0D9PaLJWHg9x1HDUGL53DK0hPrUsUZp3DCok5a8UxV3mW
dN0vDy5s+ubt99FgZm/PkP3f1GrBk3tP1uTH4EmRjmNrPjV2LTcb79uY5Ni2P6Qd
MwYZ4+4P+1Ii9Lc4rWjdpSZHUWy2WOfPSkFgqVmcEqmRJIKg0CFb566l47tLntk2
w6WS7GGWkKQmPcOvR/f3DcqkEJobHgQoGwXcLcQP9ODi3bf5GBCkg42kfh2BgEI5
NNspMAvEmOGtxXjaZeyr6cy7ZwqfI9y8uDM1+OkJvyVIWM2yD5zySpj5202lOnf1
O6nxRe1ySNpxiHSOyH9qcdRtkZEWFJVWe7eCfOUM8ChB81OFWDskKFwsh18lf+x2
y4IQh4dTvhJUgZaOOQZ46V6tnFOqaTThzKBWwXS2K2WU7UzcJFvXwqscOuZpuIKU
2r5Yz0h6/R7AQpHF7sE5f8TA6UjXNTK5g39saNN+et0Tw9ugSY2B7rO+xi1BUiVU
sExzoyk+rAP0U8/yMHVLDKYR/3NJxwi76YwUiGXVfhA6OpsNlMZS8DWyqiLQRE92
gyh8JLMxAqbQhaH/sZiTyiWaq0/4AD7DpPRZQmg1aRUzMJ9UhYJUjYBrugS5nuR7
0Y4Ys8wiz4J+xeGqmAYqwZjeHXoANxF/vrQ+I2mgI08rCJUKuKRkq+rxQ+Jx0GfZ
TJPyZ6RxVbw4Ae5XP654UpEd5wVwLe/PSUvUYiC2XXBAe5Z20H31DyIFrtfDsYDZ
XpS9afZnq3M19YJRPPzl4DBDAR4IiJtEHTudNkIdipNh5WzqWapT+UdtnlLAw4n3
hO9C23kulsPi3/VFKF9lqMDGlMnntPU2gvwB3Bvwqrqj+0C9/UquDilnXK9La330
iqT9Xw+DR3hKu4fA9G/lcz0zhLIzJfOJ3WW3Clx7JkPyiB1XPOB8SxM4P7k7Fcbo
FzRhjOAiYPBxZi6anjw4+w5Ef7jeAnfXbDUtqpHY+7nEBt7aOq8un44KykLuACI/
c05xV+C99tM4UU8frlTzAbr4kphDFpy5/1MRP92CTmyYDseVL4Wp/yJMrZb14H9S
Oa6IpybMj1//kalPDA54oogni+zdUyTzQhEH9GoPxHrvFkr4XvJoxqma0Kk15/l4
/XT3lVfIo/4wPneRgihJCssPjSLxBfk8T0AiPsJknDgpoFRQKrAXY0u0atSvcKNr
vGw2ZCjF79vVcKRoN07SAEVynKDuDFQvvk1P/PK0hDGPwzITh+ZENqTQ5DUdURVv
G6AJOjF4F5aLnj/oq/DgUiuuE1CLeU9TEZ70N/rOvrE2C58RvBMejnq+/Kekr/dF
Ifi7QioQMuzl+JQIAGb8SLFQEst8E9F/2tgGUyY3YRhuZO3xjGP2ouCSTvdcILbw
S5RhYffSpvRFTu8sLWJD7dTbMzlwPewXiUjP/J516mbtz1kZRbxrfXcP4q+BpM0V
jKic4ZnsUnQoMHoOiBiVbhombTCh0dKQBD/igXeBvxHyWvOLq1SPzuvzPRVfacC1
tHh1+EUXJk77tGF8tBqWYKRfbHGWYUgBE21EPLWQzz05T0qw2fZwl0GPTb6uZvA3
rd2T5ktvd3fFtjQz+lZ16XRz0RozkActDt4WwtSImztQ9e6Xh4h5UH9Z22hVYxIs
GlA/1dmkj72JwjYs+k59uOB72VezUSRNEql57szBeX9yHi5dG7+AWc3EF8TzknxW
TH3nTMX6zYM6mn9liSCytjtw1KxZ+paMrFzH4Ouns3WiCiaHQRa9slxeKta6a3Yd
LekVY68nfO6XYN3Yf4jGE1JZh5uivK0cMt8snUyeHQXj83ci6rOP0k21kWd4MWj0
urBmD9PADGaHx3pNZcf3YnP1DxhGU9RZqSq9sttud3XCTXK50L4j3xsTEMfPXhQ5
v+l1zvKQ7EtwWoUgrrIbugnPE3JO5kAADwE1sQsdVhfmVYVefXzEw7mIYuScA/FF
l9NdiM+2D3i/0LqcMNBVCEoXz2sZ3a2UDZjJ41IhCa0KQtbkQlYrW2yp8Zy9Kfb+
OHxsOawnMgr6uSwjwf3zSUk+X+mkx1xURkMcJsr1KwwTG5vyKX0ZaR182v0vXKJ6
/Lc/H3Zuyi6n3XS3UZygeSmHkoIP7d1EoQnrlNoFpcHHnfJp9iHUmom735ODDzOJ
0LXfPr1Rqjzvc+nsIwbfmg==
`protect END_PROTECTED
