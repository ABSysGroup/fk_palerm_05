`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pg/MXhl7kPI4zphhyJegcF1pDB9iwj8rOXeFyx84NZU/4JgHdPIi8NkpTUuMW812
EqXSL1Z5rbi/tSHDSLg0yECQQqqCYDq7QGgDVTa9rGT1kev7nruNgYXozVxdZ26D
wyvrmK+tQRP/h4F3gK1E9t7mAcWUgo3B/I6pbq4EPiNfSSd7BvYmco5ZKz6kpsuS
hycejtXTtyAVSglP+KmmVlyOXqsjLFC+EJsDzRHVsBRWbenN+dvXOTwnOyruRyGa
ka5tjSP8y4KkYUW3+66ZGA==
`protect END_PROTECTED
