`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z9svGQhiEq/Szrbcch3hK02puTC33IWB7WbpLo1k2hVAJWSYRoOrCyCcKnb/rXDd
385xFNsVMUbJ9fn6ly/B4AEOKPRT9CCybzX3u+M91ul6boigddLnu/AjTqDth2cT
F9CV2uQcQLgDSeIBV9wXfOhG2UlPla3IIjK9iTsxgLd8xyijz1ZT8zpouxw4qp4j
Rbryy5gph/7hubPT1NQwTDwz1LCSIoJPQSSZqrBv0/Cc9R8jRz7amF5D41/GD+oF
MEDYGR2Pa01HLK2t96cY57xvwKRlcziEIBDF7zIdGqsVlwVaO8Ihl0BjvxfRfOF5
FpUxdwTVn87A4UjN7MOGZakbYzCcneHRX4uU5GN4Zpb7jjTJn6JK4YXjomd38AQk
PQomhl1UyIoKzx9nrnwkM37cqCdh+/l8zz/QXz93+NkebEmC5wCG9hcy4UYsKNmz
3Gb4YnvOQgR0DsqbYjzFObKDHB7OxFlKIkGVEXIQ/ffbjKM+HL8bOrGqSEyy2rZx
5LAcT0TyVC/J/X9M8A5GoaXVQF9Zqefo1JOtHYYyooMDsHRkWX/ecCLI0QB3b+h4
iNxMZjhEft/r4i8Kgn9P99MvChTB3uqG89JIVhICnnr5J92/CW/2cd83DiYDSCno
H+9mdAkcVY/AUHncQrfIvRYgsnXOs+TEYYWtnvoeyTNjokf47XK4eD6r63AWORLe
Tmr26NAvilK1lpBrxYk7Q5SoulBHniATvQoYmaLRlYRz6qBQrtSAIf6qNIuJqWzy
cF7ZNLkPY22D2b2A/ni36GJdpDFwo7OIGEw6k5cTWz9jQyUNiwh6KwLuqbR/EtlI
O43jtNP81z098v6u8gbffC/0cjOow8RqIhU2lh8FULi8fegxDhGex7Mh8XhRS1lw
5pC2SoQWIw8UpYme1Y3Rze7kIajsVB4DLUWYuCiZ3K3a9/eVFpkHKE6ITNfIpPqH
dxVNpmp6vqXAIOX0y8UElVQJQf9xEqWhgoS1P2HErwOAvRRsftfefQK7TuozvNcx
S0RaM3qLMkvBdS3UfHwPxW20irktLVrbth3Mvncp9Qvu9Lnb5U/172L0zM0qiP1A
pBZxTZ9UbnEJ26rJVqC+Qu6wbIcb3nDb7+YguGRZTHwjkNoPw22d7tnS7ByzgibL
UDrnmxBqcJ4elqAdee2TG/TBtRi7T1J+crT6pIqYwyEidyoDqs4yevKI3q9kfZy5
SEhkmHeWAXZ1eC7Cm8+NOHFzvYhhlCBwLX+kbbHU8tcE1dBU6K7y3JZnW/s3be+3
8H4mXbji1/b2GFidQMjG5hIUE8dinL2YnmniqO+pwTuBCbQxeW+rAiVf0UOTjShA
N0yCE88t0D4EnLCa3UW8kjkFEXUOLIkYLoW4WIXvrkPGhdNZQeTPIKd0UIRAmYbH
T66ejCoIC+a9xWzaoSTslcvpT1YuBL9C2pbVGif1U20bVOvz0pIxkN9EzR6nlxLO
NwmkItW4hX22DlC5+6rfOA==
`protect END_PROTECTED
