`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EDedZ1uWQVVJc5OuJ2p3BwD+pHknf/MaWt7gsZYTAxkKfVVDBQWK9hy9hhwaXNdG
j0Q9VmJOK4Qk12XuZU4QlRUhFUyU5PaV1L5F+2yVAqELK4rzSE7O5kJYbI9VwYex
6y71L2Z13F2T8JU9Mnu6V/1gBaSN/vz1Z/yvxSf20qyEyI3eTwmeTjhZLr/zdTba
ZP/+3UlwWCwSW2RNkGzmyhh2eh2bOwuS4r6MaN7hf80bComsa1/Yj99haneQQBQf
BKrwVbQ/aUKpuK6jgcMv7rVDbT2TmwWHHBSYsnAQuOiZ7aPDEzaoTH7UWSUCNQ8B
BjdtB06l9IMuUVE/x8M2aA==
`protect END_PROTECTED
