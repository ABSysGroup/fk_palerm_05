`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PxIfabjcbcZJdxG+6yBEj6+NrdW1vp2RSRVt7Y9Ih4eN54X0W+PZv3ovw1qyFKD+
neOvq/5tlcDKG01rds2jD7u7BbKb21Q8HPoV5syA+qciZGQXuXHUDSdV/REzC6VN
fTGtd3JlHNfNV8iKm3f44zmk4Gv3IcgILcjIgthIjsp1woZbvFcMryD11cSrgKaE
3dp6xTh2nFqsA9PjSoOmIqgxzAiY6qYb9mOo8oyLU6jb70tANxdMY81MiClWLGLN
Uo5YUw4PSo2RQ0hSfRWiyMcyPqxYIjbyzFswwp18N11ipAmJMKzp0W+Cg5L41ij2
7S3jLqjQjZ48ej4wRC15scMtfty9XvWnQYS0H2G28D1czA8eW61XqPnzm9Kbh9xO
95D4rbsi9MdFmmDCbmd7r2+M02C8rh+3oPhAYYCUtlmNVVL3/WjOEYJjSET65/zL
A2f9b6zZ90SBCShuKBDBYuda3A2vrUS7qk10/O22sLH6+eAfVmu4SoUdHivVEXiy
3pzPqtA/8JSfvkr8x7/QL4c51TLI918b822LgN3/5fyTF97CJ188F4OfhyGMKTkc
iENhUiySF5SMJGL2kOB/G9XGaOI/nnOQ+LuxXNQ5JCA9zyRDLXLSCGvUkPFdTWVB
ol5jrT0VTqAibOP52wq3YRbt3C9tEg1BcyPZfQtbJGbORV7DUYuY4WEIOj1JLj+q
SmoDNZwhGh4WeFCdwpeYCyiH9VVKQLfq/p7iVBdcmGEYGPuPq4obs1nxstDRlcGF
0j3VsJmn8VayBQ51k7Jss+NerOWt3F9LxHIbVd7Jb2H6CoJh8DK8gscvmtBTOy6P
q+mr5CE5Rf+m1i/snt2Kz6oF4go6tV6vffiyW5IFopGhZzPS+VMmYJL+tgnjTXvp
3WIssIAYI0HI7B3f2JK73sEeSXJ3YXaEflG09B6bGOJgIVewLS8rr+icYBvwd/TI
`protect END_PROTECTED
