`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
poJ9RmPiLPkV0sv1+NsC/Rsao/XZoaQ7qI4QkSYVympph27ZqbCtzO0TXtyrugGS
GaVP57vagGf9+8XC5MrJrs8ox1+/TA7ZjhU/1nYn4XEo1J2DF6FCMYOH51yQEao2
yUZxySWIuYCA65fxE7/CTfhoIYvT/pTHBRw/cC0TyppQmePW2b69IGqRwxoX+YtW
FP/VdCbK8ub3+6B8rdXL6sjdb3YGnGPO/Rwo6cpwQWRYfilo8swQnZSJtTAsSKUJ
Dsds0WzCM/d6rrjHeY+6OrB5sQ9+++JnF67l2UtQ2uhRnKwVKIofc4KMWJhg7ZXI
H9Y5/etbOHn9GeWjf0tg0Mzb6ag51jTqvHBnGz4ZoeU1FAJV7zUiYkAynaoprmPd
vrJhL7PMER0jabV+E3Vu99EWFhjO/vjBVVIdsIOKqFXm+0UiTYaPGa/OQor1x5Cj
RuBTlczWkREjyIaj6T8xyD306lf8LcyEvesTWiup70z4tEDS1UHxFx5QyBWp6n4v
KL24zZ5Ft223LJQm/YniZX4xz0sSOCuwY+3c+bRq1vSySgJ++eYWG1UPaSzLzBec
eYU7CMYCHYzXkcHys6nG1KbNojbKzMn3PHocHlaWFD7xAIl0vDDMHE2X9VJhnX/4
cdZLOdZeKAztOjvuMYRq8814g8hjkH4+LRW8Wfy4nRae37G4ULSMtocq3oHh9Ae3
byt/JC6k+EcYiZLrxIzYNNy7V5ckRSKwwJ0Dk/raTiZLgI7iGwsddclWtwMlSUIY
pOvli24eeaSfk7AWhm9LH3ubm1aJJxR1QJ//o85rG6TCo7TmuY2IXhEjgvgh+q6b
ELMaUNRPv0+8JhJ93O5W4XU3+65xyyO/Axlnh2S39dWSmYlQ3DxA4FNRmwSzo2/B
XsoRAKR/RTFLEG4zKBYs14XUg5SkNrddy71ZrIcE1ySVD07NKrqwSLE5fbljg+0u
`protect END_PROTECTED
