`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MbzXoKdxGPl21kD07RuLHMbVlRGNBRh5H3xCYqIVFz4/x5MD19oAyyjrv82BcFi6
xTfl7J1LyxzWfwQK1SpxXyYitu7kja6eZX1tfnHWku807uup83JQ9mOdvTifZFPW
PqhuQqtF00KQD1m3QFV28/xu03mZ+px3M+fmiqTq0St/kwx1f8L+d6Zb8xydRkKv
qujgF002HD7IYVDDoEvBeW4vdr7uUVBStUEoLu5ju5r4Waw1KLD+MZ5wtLPGwsDp
znya4/c1iw0kEGRsywUZBfycSzqVmI4qz9CeIghwvUcs4DvD1w+pDC1sH1arTegT
XjVeo2J8/gTnXoM8tHRkIaQRFoAHdZzR72MM0hfQiJw=
`protect END_PROTECTED
