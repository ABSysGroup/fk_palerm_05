`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k36GmgZVAdRO/vJfnpZ0+CNbUhapR7k6Ky5kt+Y8DGcqXqp6OZ0RwDVZebnFG0mp
3wAeip6HvZbDw/nIzUz93uuosaZILkH2VyjZy5EqhhaY5OkOjjNWa4gK6tcBlCBh
5RKy24kNz5EHAQjSbLfr60FihulazC7dsnRrFVyNZCk5LRItv9fNX/sH23et9qKX
Nygx3Qu/7oiJV1bX60lA+omFDQ/k4ToLA3ZsefxCBIpE3FjHQu58LLs15aqcpDD8
oAE3y65erZLs12uMr8J3wUZV/F0M0ZF4qYFK5QZ55WGQGjF7QbZNlhs0G/omN4kH
gwGv4NffRcTqYB0PcOMvEmFyR7v59RlTE5UjNiZcDYY2flISUxVfK4j3aQ+mJa76
fvChQvhtksW+QhgArwFSzIHC1rz9VbSdhNJH45EDrHcoJoYdiav0JZpzPYZMX8ih
LoL7FdgzliZY4NeTyeq1FbwLC+R5BK0fHAexCo6nOFVnLF0mGcuBhvCFGjbt6lnB
`protect END_PROTECTED
