`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jGFjJzalqO5yEraHqW4IvV7Whku5c3TVEwH+jk+zMEl6IcNneJs0uBI77a4yc824
wjul/fAej2ZjLp3oCKS2y7daTpOVaTFb1iWBGDL3W0rMwae0zpeAi3EOxHePeP+H
Ymdj2+kSoFAC0Mz76jN5dJ8l3J9Ck75Dc6ylfSCUKL/GiMBal/mhFcHDPQTP4xf3
bppzpMzoFnq9aIjMmq4Ax4dyjc68zp4TuhYtMNWmB0UfPpDDJ0FATtE6ZGiOH/WA
Xy6+jV2zku8A61OVlWVAPSyynkoNVHukKvbKh2a5DNM=
`protect END_PROTECTED
