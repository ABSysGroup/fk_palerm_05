`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ybuYD2eVsLUpopsiZNHDhT7Vn0vEQpJZDbT0LhDloF1eUmdAmPlZlK/WE5hoLu0S
lLX+E2nuJ5w7Kku+6nNPhJOTKvszmPdyVdO7jKNebCuegO3IEaSlQXh0wbIM8Kba
tjvhleyKr+g94wefBOzI0l+NZ5TOcQW/8HCM9oeQFSDiJZ69UIrozJkBDjz10PHH
yB2A4fuxxlWhIhBi5yUdxKL1EY4XxXFuM/G4O8vU3cqjtBdSf3fHoqasC2zu7nis
YPxY9QE+l9QTfi08rnMdqzEjLeOLKCTYf4O3vDUyn7oKBhAfu6dsN31KBW4TpM0d
qaK7Cs2etIC71ckUXaDVu6pkdj96JzP+RRYmun6+64aS1YTPcGrac9PwtVBVALVM
+XHHkaAIF6VZJ6U+7BijjQ==
`protect END_PROTECTED
