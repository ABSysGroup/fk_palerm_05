`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NnF8CgqvaTTqH7KiG+nd8/ClVmBA1KZQkbPY+FNwF4nmd/KcUUFlZNZAL4IhZg8N
UHhdN+SDTrihU+aK600ceLEsTFsDddvTie34HtDwzftcnz2kE6f8DGkKBPdNThcT
QGlujfIquF5qc9QIgK9AWyKc7YKt39MCLu5eyk3PAeYsxtK0e1fBSHXCfLXaPc1S
0Nd8xfjjG6bVds86W7KPxDJ3wBt19FnfSZSIVqPP3KynOA2thJB51hNHHhyjfkqj
mP34u7I26IMei98S9prnYIxqyQ7NoBja/1XM1il95dixBGYvoqb5rnVLJQHjIa6p
LfwEgb1k8MnQSIdlzXfo7ozLOCnGIhTmFqzTRE2NnKkpzwg0aCeLwYQlxNb7P9n/
lI1wNUr+jAS3Cgt3IBMCmw==
`protect END_PROTECTED
