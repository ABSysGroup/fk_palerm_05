`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CpHHZZMTdtgzeywcRA5o+cwrBTEvHxrVEnIv4MeoT0aNMGwGEVn3lLJL0fMKnjU6
tAIfYrH6r6F2/MtXjjvAFzUSPyXzaucPW2iyxtNv1Li5gPt0/BGDCsoi32g0JMhK
e3tc0a0hrdOg0kiB+ErqfAG7APifuWbmku7pnxdKgML12ywjcSGs1hEVSIU4bksC
dTPqZYH7DG0k6ptrc4Zn1+UtMrHhs38AFdhqe1afmxFaV7P1ARDuUsgeST9s4/Pr
mLpwjl7auKT0UwOGdjZH8H6yHRTzBxiUjwf/OA20ezgFoGamsDxlka5wVHXGfGlM
9meUWv1SEWW0zCatU6Q03ajOuhLqQZbm1EH+e5wtSaU+emyMype2QzNTVW3urt2g
bE7/TrXRwTkzsW/Wz+0SnoAqMCk2JXWkyknlkWCzzihUx2qzRIdajb2jDgXNet2N
r/c33yzZ0Gj6omG3qxhDIMgAvB38+ePmYCLcMysLYLStL20iiyrCBGT8QStZpqnG
pMSdhAVd9YASPP3PMd6PXQ7q83OEXHkY16YDYSn5Hej09F0MpDHN6I0S/fhq3nUI
g+eYbYSp/bM7o4USUmHEZQhKcH2NI4iy+o4Z4zKCpj+cws9YnMrCZEwYiAPnml0G
cmCH/uPvBX6K5JJz4cFEnilzDJoYLPt3ZQDhBlqA7D0=
`protect END_PROTECTED
