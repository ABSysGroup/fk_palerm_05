`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P1meFxmUpZsfl8xbEZsS3IKadrPoHIF6qj/cEsdeYyXX6mkgSpgWUekjw1Ny0dPt
dqrfuUYcK8c1PvYQtEXlqm3wPBIm82NOHKX9PSN9lWqjCs7DuGSMuBD8Y5tSxH3x
bl30TAByMoMYvX9giK/44SZ/fetEn4wWsLI708p3wDPS4iwXR95eJBxQYaus83lB
ap9IpgL8qzN+/olgTgi8fxv0sqFeneXsaJkhTaEQn1sFFwBxPwsQw6/UJB//WyB9
tQpitRtndgN3COav4FFhsA==
`protect END_PROTECTED
