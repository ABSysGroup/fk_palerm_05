`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
43TWl+vbvbAf5nRiGRdRcIPEY++S6cVIKys4JGKYoHNyZ99fyvuNpT50PxjTLuKg
P8ZQrSF+2GOZC7AlbGKUVjldE8srBMzWyyU2KUr7wssHzJ1s5E0aiv+ZvpodvCro
L8R1o72WnqKXnXXfnnsDJ1XQ/jQY7+haxKJ+Cs1GdRTUdggsMpCZjbjcqN3Bsb+T
nvTb0ZB5r1gNxacYcWmm2nFyyBbWK/zoNxNsCG1JWVuquvyENm4kjA0CG7mdTg9w
SFdDNGYZGo0CpRgmwBfHQfEWLCr9fbd+NxdGCwEnxQrh5zx64wPSb6urix7SB38Q
wP8e5XVPgtrBQKh0SvkdeRYjiRwYCPSgJQBqGxhRj1z2bUrhK5BRNLkBo4k6LbA2
fe5SIM7YHygaoTdBI31hP/wPinf4lbpl1rZmhCGvWuRxFVLnmMY42XFQyKWpxa2y
PTW/dwlpzBBz7m6y2H3KJ+dvCC5BsND7YpZ9GY50IgJonV6NUfgrLr9FQ6GhIflG
PKrJgEsuNqENoVXA9gA5emPWRM5RuZOl3HJhNt7bMNZNzjkzpvs3zAnae99H0xHQ
HMyIMyIUovMN4KVKXoRgMtKHavtWkcnsEg0+HVI8jI9QsW3YnkhaXYFs/6GJww9I
S5hUwAJL8imN64pMd5R3GcgWL1N9vjaGlwPM19ghQTDFjyMSyaXTZ1lFXbrno43b
Ce9w3p69HEL4AQ0BEFSSaQ==
`protect END_PROTECTED
