`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KSwChpclOMX3YnooOW5new6x8s8aTexKCLj9MegVG7Eh7mDw3R27NiJUW/iRGkOP
dpXFfb1TWTu5tCIr5X0Wmai3S91tYmj3eLJvAdfS2LC0IN8A620Ihak9Vw3EtdIQ
IMfvP2YLwQe6HgeS6dNxCRxQLmKw4HwIFKiwtXDHHZVx5K55WIQnGMu9KY/H5v9c
2sx7BTMT6GYixQgmC9vGUfYZWTuiW6/+VBSXwWd8cYbyh0NnE6UHecXb2ldbanfC
p45r7+/PIwSPBCVEc9qpx9R5aVa9EoearkpmSFB7uOttMj3A4MTqFbtjSng9yM+a
cxyr4n0Tgs0AdXtlgGAL5YDn/Svp2N4BBEH/zEgDcyIYJ6CxitewsvA4pRJkK/HM
BBUEZCFlFQt6H+eou1kNqCp9qRifFuyfVm1oOAaZfy53nt9PJdgG38Yh5wkBANrX
Cvjc0ryXm4T02w+NaspZUCZaqa18lEegdE9u0pMLeq4C2EtdvQLJUOpjsIi0KGfb
7c4GyLcODP7yaGKYtOtfSLeTve8PwL3UYH6e/tZy6oXlzyd7sZLPOk1yuB4nieaV
daH5SxfhYAER3l3Tjt0HQ9fo67zlb3SviYKJSrd9PZrA6aubzRUOnPN9c59920uJ
E1n1Iqk/MXiyeIhX567OWdMMGLrtppVJflniuOyxOE9CaisWRlfF35ZqfdcGGYG2
MW3Oq4zHgPVNEhra/6BP0dIHX8kxgfp2iZ6TmbRL2fegs9S0F0FzQRukSU0ZWQDg
mpyn9AZvKSN1yDrMenmBIR5D6z9y31OIgxflA8Iz34nXqXITiCEBgsQ2Z41KaZfe
zX9PLMLfdJc0DrDIfpMiBnnyChdVdyYOlrVqJBh9JT+Uk+nwGD9bYySe0LdyEhma
dp6SSyB1RHiY8GDuZHGG1WGKUw7zRHasnDKcKTjY8KKhlbAsG1sYzVZRtOeqAC9v
DW9Qn+ljTDWACxTh72VqHyijcOSnjQYw/6UxMm+UHwG2C2KuhjlWs9wt8kxRyDGm
`protect END_PROTECTED
