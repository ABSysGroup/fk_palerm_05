`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DVH7Y7Hq0vgaYl4k2GKofgbp2MD6yd8b1stlQXZU/19O5njwDV42g6Hb5It2PYSa
4dsH7ByVBiPeyenxdtimEfpsxT5PTtpVKivysVBQzzz4NK0H/wIGqN++IaADsI2e
0B6xV8hEqVusAuVvlPPBsevFcXEsjYKwTq/uZEHnuF6VPIgU/8AhkhPeHZun2Pvu
/4W62MASZ1osgzZCR4BT57CsZSy5AfnTUuKkmPLW9JUeWiqFCQN6NjL527KcuUCA
sRVYoCy3uickptPApgQtSiw8n0GezkoZcPL8AF4GNcqej7kcshgKg+cPf9aakiI8
5B0hu9Km+npUod+EAxVhRt2XgJI3ba5XdYvE0iNSWzSARSrToAFB949UEExXqOHk
UjI4jQiWmI01QJEJQGPfnTYXePUcYDWt0i3sulSOUFkeAhCpNJ1VUpU9H6GuiP79
rPo4nf8rv4QJnAHXDQ1EHlEgG4UpVC9Bpl0KNxOPtsOUtobJF9Me52t4pSNtGTwb
dFw984X8YeZUS8GJeGpBgnAhCe7AxXjL/tzmoVmXFlpbWX9+IJIfN2F8nqqOhYm7
wLTPU+MUvEhxIB/no732Y8KgP6fkyMyk3CfncR5szKCJW5RO5botezFfaBFzzhkv
hbzx5dxOYB/7MoGJJ59qug6nht4WF9UJ+9VdyYq/ak1VmQ/Wn9AqSt9ih5ZjYGgP
OdFAQK6fSVeWZC84l89iUC+U1tSuGAyBx1vob6bMzA61tPGR4N/Hla/LSYuTkdds
HerQSBovW0z0BczVYZLMbYkmH/+g779JaSBp3WIk6Vcwr80xatNQOKYKsqn93j0h
nUlKLvPrma6muPRbksnSU7NdPkShhKr6nacFPEaiMPf5U0Cvh8yO3y5pVj40NwxM
/bLvVY3ubAT4Ht0MR3O6AR2Z8elHjog/ZP2deptl6ZiOHdHmRT98dt3w8gvK7B7Q
Rs0oNn5NmW+duo1Ujl4U96dEw2q3BvUmk6ytwKNL/B3zsmKxPTDXiT+rxb8aTS2h
Hfvu8Dlm4jzDnvN4rZqScNCOAJQBEuzjYzjPHx9n8huqCi4sYenU3VjXUK3Y6g6d
jYEAdpqjsdsCLIHK1nmt8A0NnbJxon1kI0RS9xS9R7+krHI59oZr/IOIJ+Cs15zs
rn+epDJx7kZGhjlvCbBVV00kds4PQtTBjWBlWwBPE0mq5r3yPwpIatL/1tHKNvaE
y0aat/ORoTnt/CfJO9/APpgCAH2g7xo8WiMjmow0XS0wolp/zYRtpMHHrdqGJiva
Xa7O6RWuFueQdbezC9+xZf/P7k7FQfekXNJ8QrYdCHyCq1Tx5yj+E4aMv8F5gEEk
LpjNbpXoU+uAVORTQxyT3+0ImvBy+SVOnwXNuBbSTK6fRps4iQdGGt7/fbp649If
6Ya5aqDcbiEQSZEozmRqD/p/NLVD+VOYD0ZF61NNso7OzGCrxcQn9ebh6TXvmToH
5tnFYofg/6Bb5fkMJpKQ5vBmN0roGC2FVKlzI4HEgLgEDqHxkV+yQnCpM13T1RVg
fqUlMJfE9aRtd7Gg2tiFKoy6Z5uE1UpP2I5gYf43ip/PvmRRoKXtcqO+f3sYeMrm
vOgM1qQpS5P9FgHvzQX8/UXdIyW5MK2giDFU/CXNHw1wV1XK2Rt65I8AELNQccQN
ikcJgqDP0HIZX2fB1Xauzz786flu0CpjgwS0WTP+o0Nu26x5nE5aVGLgO1RXinmh
3sdELFSUiPxkHOKUE2W5b2w5NcB1cIzH3HGKFdL75FDFHppgKXd8fEe/VyzN/pfX
VdHo9uvM0q9jT3cbqus40zoc6KCYpYhE8x/pnBeN2Fm+1x83C0jfpd8XYV58C6w1
UncB/CfvVz9aughf9/RxnflM/iyYfn8m2iaF81C8QxqHzA/5Z6krtnaDDUh6+PpX
XMvBfhOKlu4sTwdRS7Pa7pbOgezMs+NyYKJ5AP6Ob++UIc6EJq8uUyTEe27V8txe
jdTzhdIEDUEOuuj8fZsmzYZMZ9bpkR1kme64Tr2fJc7U+y8sHShdKVQ/Q7IQtCsK
NDb9DXb3uUD1Eqr8HCQa0hPEs7koONB5nPR5+YrH3plU1SCsi2CNRTPWW9GO80gT
U3qeGgq9lVOflH7/4CfMSGLYkGGhg3veJbeW9a4Da1XlAS12dNSJRDcqx+OSOgOr
iRBEccIJeO9bVMqkgYUvDukR6+xahPy1vQK6LMwBBQMyzMnd8KXrQXYhecgvzm3s
SGxWhBiD6TVjPJb0onMSBCDS1Rdblwic1KDvmcRcCxcCdqCJ9zBSj5IFkNmfj1cE
kjq2+qgXP6hWE3deQxW1VbF1W2m3RlmN44ChC07G2fL94cJJXvm6hn4wTvhfR0V3
BumK3iCDasqUZs8xvRgi0VftxLrmcjWry8XXnkpfwa44/QlE+BvwWniET8kW+/Md
AG8GSULuue5VHo5EnWi12bVm0hrLp+QgAVHxaGDCMrXX65t0+4hiiinETMEHgDDB
B4mxI57O4iCGQhs+apcBAVvQJXcqTWHfc/ZxBUn4OwGaLabWyzsxVyo9dBT/QYQv
HCvSwz+A8TzsFEqIOrAgSg+5xxDlt9PyO5rtZZXsNXAEE2Q7Y5EmZZjZHraRtqQi
R10Rzrh/jR/lknehNOc46mm2Eqp9SD5EZJY0AVgSqeAHiKzd9tMx7p8UuOoz/o75
bQ0zHWV4p1iXE91tBVy7lHZ8garMyR+iRiBm9oa2cC6qQtQ0RVFsnrqHXoNwtaHG
hYaTVI57B248Vl3aGAMIlOdwubhVnFvM5ftYPxIhPFY19hK6yoJLalJ98cPA/3Hk
7++s5Lkin8IGJk4TJ5ORawdKu3bD1E5hzBv3yIh6feP61oAU7/dm3T2lsW6ot5pS
CPpP6uECjfeNkjTS7xNelmXh2PqtW5VhH8IN/MqdSg6QrO3WOiHVHz/NMcGogTlE
`protect END_PROTECTED
