`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9kvbhcVwLA0h0hWZdetV9qMjJAOkRETwlaEW33u+ZK6Pn6QSzJ05BdMgH4B5YO7s
/vDEUApXOBkKcqos6jiOcQ7eWYzLzksadYC4zDeC+DQD95ORCNQX5VjpKG0RrNc/
T+voUBp/ezm7n4CzpMq4qbHnD2ysKcDgX4GVYSQ4GWR0te+k0xeSmtmkWIUY8aCV
2i/nCvDskrMfhz1SdPFURn4MC7ZGU5yVsFtMTYtpolNvSjgv/hQwyxa7CXsDQ6+7
kgo+mqRcM/XKE2/ofaS2TUTJ9r9Kq5RyrxOkz/CIDWuPn8idVvLGupnRfXzTKFBf
PXeJKtgbQ8yzMj0BrZ7/pRD8f6d5w1XZuwp+mBupXoieHiMQ+4zapqZ8rMs0WyIi
th1lOjfiFo9tBZ1ryb/15C74TkIGgSmotFVyphYQUSYfpXLpGJIPCsAX/V+hZz+u
EU6PYA4EwlBkPNEjpZQ5I6gej2Gc5i+PjCs3oZs3d7/iIqWaUl5myjm8NCQheD73
Kxnskwnx9lOxbmfFzysMo7Neu5S7rWoDz3FxD3IjRR1F+INW2NcVQkOAzL9lNXX8
5ptdXKxG/G5wzb4EKmqcLDTe5My/3sja8UvzBK65wwqMABw3Cb3sdQNLsD5thAhn
BG8WMQrhZjFh0huXVA22S6V0wVBn2AVvXa9c/0d4T0o4jSwfygrEj0S6wdbHS52e
EuNIs83MgAFQcqyLq5GU2Ci0RTs0OvVw5GYqrGQDikC2K/P+oGSiGQnZm4Kwgm/7
56XZ2i4HZRT6OYMr5sV3SLfKjkZTqRXCtslfvOf+0nx1Ccd3jDEKKNfdLLAQl2A4
FhuxswYviwn8gUd/koF5A3cMs5yXVuPSwlzpvMn+FA+4uPbQSZ5KMrmhbVXMLrLS
CjQKKRiA2wrdSoI2wHob/HrxudgKR0oB91Tkp6FbCKDGnOT3Dq7/OC+sy3Vira6F
IGmIafSfCdtsg+TV3udnicG+f5ECTq0S57HNECunRp8opyS2z+F7SP1VVAfXKZrf
6Y6tPudsJojR34hIFRokcWhoDjOVWwXk/iKm6akMZ129hFfqYnKC+CKkFfBFFlUE
stgh+lAnWawUhZxx7FelDLLsp/5wbKH+DeUiKeD8WcI=
`protect END_PROTECTED
