`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XjiP8NZ4qmz+68rzdorkp1dRR2RpO2SAS/1xTNdJ+dIc7N9Zn4W2dclbpXvuQ6py
mx1xA4de9/Apqx2YWrhuFQNLkDfTZ6344tiAmZNKXmMi0ab/LvOCvxIwx59pv0g3
KXvLamNEemS544FL1matR8Nl7pOE/U/cQ7jpPdZHljSFUE68ve1b+/Vk5vZxPua2
jwBm2NbsKeEV/wZyASwHUd4VfvI228MrE2gKULcnPWRVACtNGwl/yAw5AEXGZqJu
XDNbMzpZzj6ozdom4JzCZoS+CmOmwwDhgU+c3f84XHp03NwLa+7NOpMJ0nfXJJjH
lTkiRLbtJDJJD2I0i+rCjNR6kCi91IoRlm6+AvtcXVddUdcILynnCNc8deJWxDlX
BtHzfIMuOpniESFcaCk58Q==
`protect END_PROTECTED
