`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uBtvxmTI0+EZ9z3YfONebnfp5JZNLHRGVvfV7icGoWKvrfFswt+a0jbchX1x4IsF
kxcdzUi7EOJM1Yh6A7ppOfGlGjE3S3iO62p6CJ63YgprXsZH94vEZKdw/ypQmsJ0
Bwq1JSq+a6hCeWFOzNHRFHaoRFH2eggGn+tARTpuW3vgj4LTLdE14r2WACKOf2iH
//dWOcrRIcxLTL/jD+OC/cenzj9StPsd903lB4aFuQmsAdk8IdHIxLcXAqlpAkdS
t26dM9S9qgovt4gdYorFrxX4NYIHPTenEi71mcj06nc=
`protect END_PROTECTED
