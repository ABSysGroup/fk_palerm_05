`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6PHE2VFBt9uSOqZSsUnRfbecsG1iXXKDRdIUa2Hnz/iu+NZIVHKRxwAyDmtlJhe1
yX9CDplTrrnXnUgAkEcSNvet+0zzBvJpQbwo/q+Js2024zehqtr7NMT5C7IcKW/R
/GVHyyEkp1KvCWTk3AHF4deEp9afv50HhHY95OqA4qGscl9/vDyhD3NgQvuaEkUe
5L754UaThjFwxL2fYzCcWnAC7co3+iJQItkAjtE48gJgHOQ/7Vqa0c6pdLhe48F6
04Mf38Oy66NwFtAyCis4gjLXc1wFr8nllwNJGLQ6KFS6/+pLYIo6Khsw2f/1n2Ej
9b7Q6Quq5kc8LWRL3Ge3H00JC0RLM+sQli6AVL8fDDiTQfasI7HNhmVv6nys3fCR
zyIamDNYYE09OGpXyj/Ls3BbGNSLd0J1og7Rjf0tzO3vbHLW9q/2EMwOHEBvXX2u
zflTV1tIW4PM87dPdNMiYpZmh64YLXDP9A2GxtyzYLP6Gnz9PgzEEjDBGsM/WrfF
87IdhQjMDsOAnwsZCuSV2jyTFXtVr7uYtCbz5ssOVqvxf3fxYs4yaTZrEnZsW7tP
40mxu4csqAQ/uz+aXUf2iej3ZIax69JynAvpbQwkEhla1SyCaZMFkjxXHIhxBLC6
w94fYtjxAF2iVNGzSL8zFn/KUSmh6/6Vh5oHiRYjyAU=
`protect END_PROTECTED
