`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SuX9MbJUIQLH9lv7tuDkamTKQissMswM4xo4E4B3UpnMDd5DGuQ9k2A0ftEFbARO
XJWeEFsrkoxtOev8ftfbn4AUH4O3na2E2T2q1DENhjMX7TAlovO1pD4C7l70CAZC
Zmq205TtWkrl3U/No7EfRowRdWwSssRM7ztNrJviP8do5uETM4uQ0/KxEKcM7T4S
9Yz+1i9Ps+sMUhud1QUrQHSqaRT/ZtZBRl0BRUC29wTdL9fKjB2HmAaHZiMMOGKk
0UKrXHFvefo5RQSjhoLAK0zuKq3Rm/ITKpVlR8wyTHZ2NgQtXPM/77Ri+5OTUI6w
d0Dso53t0/c0E0VrCU4QrRmAvmifxX83QuK3U7Jsvx0I2CXI32UkvzKQ7AGQsgm2
FZmj0JDxMRUbjBd1UWXpKZUd+4W70pB6InbpivgInnSC0nM711fq9EXB3ofcZbmc
2gcmAKjb9l/6Sb3XFpTnwg==
`protect END_PROTECTED
