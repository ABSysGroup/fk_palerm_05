`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f9Cox4qaWeYhS3RyMT/kqvvajys+Tp0+sDhNs7Nf882X17vnHeaiDMUZaJpvghF/
C1PSiFtQcJXXeB30r2MrClDQmX/NE2CQte7qPOg3zIQoxfspjkkZFNXSF5NBmTfT
U69PjNfzd9v2a0DzzRK+LpBKDNfrSIif+O1U0+JU05+9UpKZ0Q5ZyjacfwJvZ/zh
mcPGNyzcrSU9rD7VjmpkSHUrnAygGgWRuDQfbgeiESo9jeLP3+raKgkb3uhiCPjv
NduP8KB2Fh2gX8/DIGt7fJiu9SrPkKEHW+zHb9WBLCDR+ak9TywU8INeTbIbRgpM
fy4KacW+cR+qe2iA9oxrp5GPA/nATek7STXfWfhV7A8qpIxu+ptj8hacpdhHx50f
gbw2I9ObQuPRv4r8OcbpeMGVJQdKjBbfsjaEDayq7C5yqhmYN4awhqTrO+X2dzMQ
wwLJnpbvugzOmFFCYHVhoMCM1kMUaQlz1HOAa31qfYnqbFbFJMejX/tuUEoGaYHQ
yekcU6bPQYpdu2KmhdWy+4GzCh9bSLsSDLZ0Z7wE4aK8yRDLq/6CaO71JH7Tjblk
Y/eANgsxejLfKav7WO234sr4wV2rTJrU3yUk7l85j6e1Gpb2ek37+FH3ZGj9DxnD
QduQV+zyWyfcUiIanle/o2BzQfGe+KH8LiWTOAmwWHo/Ts7g6hnqkqAzHt0w/57B
zFG9CaAR2IuTpqk7dw5qXhwFx0KqXhx0DoPUYXqynycHpa5Ty0NPyNtBi6QzdSdC
eTNfKkZAhkvwiCtw4t5yJ9RLQi+BhbTJql70iqW5maruPbhOTPgCdjZQrMNcRBZV
oGAzdPsgmPWQbIAZDvgIUHIL/8Ajl4B7N883e3eP1D/gpUktSrNVn+15CySkmG7e
bciQ+gjg9LTKmck2wh8NOUO7IBOsb+Jl8CKTjzEDa0gyL1/yYbFjKowfAHaOpqLs
5KFG+gPqyim4J+uvQ+qtvbvv9wR44+JmmOb2Veg63N2NvVd3bRGkk6orANoqrCMc
`protect END_PROTECTED
