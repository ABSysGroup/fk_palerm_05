`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1tqWuQxJkVli8Ov3E72+yGfsseAHob35lLNWdOha3d8bnxCA2stqKsQGyW7k8pkx
+hMk4/bY5R7nYY/33J+C3j4QGIZEbQXxaylSqtXVM44jTEZtxMozLNJZOCVS30Jx
fwTyXM6g4cMhrIbo1/BqwCsFspOEZAh70JkABURr3GzrXnhlOhcX2olxHlnmkQi8
52jcfAgxwlGb9yj5XioOxLcW11bVeV1g8wUPULOOHoe/7m3fZiYlzl8XIrO+F8Xd
hwItx/+rpxhHVbe7S3kZOPMY77izkPD87K6oboKrFAcAkx9+ZZzLpIQSxEn2Uu2k
t3Z8c8yvuc1XoMUnP1VHPcyBN+ND6j3rTErQrGzmfFOYpsAMjqxMtzPDy3dglWi9
rDwakZTvS7GexHBJQor2AC1/b88FVas6ylOsqgdfTUjU/KIJ+hNvgoxd0McHv2uP
4voCXzFzcmLn9Zqe4zoKPRL+HmDggKFd7HW+17OLXunBFgVCq4pT27IsbmD18hvq
2X/6otMSflSE5RyodJXSQoQIcFhJ+2zwryJVpG/eTEUWrTXM2AzPRiKnKlgzp4Rr
LSpvBmd4SIKturSPBXRMqgSIJZbxjWznrdtcKI81J0x26hldr5qUJALF8kiJqC/g
ZX5MjXgJ/xisQ6P1QLI+8IGjs4N9wVaZhB2qpnsB5U/d2CnKYGDkSAH2PgZK7waV
mN8mJ+aslOWa75GFbNMsjmzDcZfGuKo0pD/hYb/snmut/A7fHDl3k/GvhN2hCOQ0
TAbX+zCWelcCFvwkVSXoVQ==
`protect END_PROTECTED
