`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WjNc22XXoz3ZgxOZWnZ7PrPRhPk8aMKR7lRU8T0lpiigjbnxkpwdKvBtiBPUdC8v
YfYRQuQZXPli+Tc6UWblWwINHJgU8jPKKVYs1fKnytYNdAS16I54QgCk4SE17bd+
9atVnBA5jYRES3iefstaA1Pmmv36Og1i5LnZUMuozpHdhFCwH8I+pzkxsaBPtY4e
AfBRpoTaknTzdvx/hIcXWAtO2PWDGea4OTe+ct2IrFRInGXCnGPJ28f5xXxGHaTV
FEfLSaXx4gFoLHonq/waA4iM4QjTFQQi2SN6o9xrBE1xAymgdlcf5Lb6pym4++mt
ZekbPWc9v0rgX2zJqIPIHN2PTSMoZJW2/shcMv0aRZ+3+8JU3CfgG6b/XMP8iIYI
GWbFXz7KBSwca/AZnlLLjdAtWsPqWxA0FsLmxZB7DIX4f5XfeaKYYBXBwAnYnbwR
gRkaHdxWuptOkftpEcI/5LtTRkkZgwU7Bg3fiwAzGFHBpvgGc9CojA4B2EhXvGum
OsG041Ov1f05BxPslCkuaipMV2tMtrWkC2ApMt2tcz9/6/7lhk9aMnwb3AFYNQTz
BR1LndjmHpx9XhV/u7addv8bj+zGSr8s39lEE/6MiRsMEY4Tjz510qhqXYFrjocU
8Esip0GFF1Blc4kMF6jaxNxiCwVDuQMj2jm9up1IdBn51ojaY9DXRlFxv0CH873o
tlGDHZerJJQOT8uRD7Ho8pR7m4Uk1GThp8ZnF7iMVvou5pIyU/kjVjGzLBW6G6Pe
ecliuTMeiHLYbLobj7nHgPE5raqWPyg3eKmF8B60w7maAxfNNAzUGKjSGc3CS69C
0nCIROAwgOR7KKUDryyA57kMcYgintraXfM68ZNdGplGwEbpZ0Xb7rPb/yq6gby5
ZRnjSIQISr2ODS6ntwJ7PeyqAUV9L8+7JNUutiKqnjhJ/Yl11yW1Qs1bKs2hVRRo
h2/pR7EJ/5KGvF5mYKoPyRIE34Tv3vsjtIMXRsqm+rTcyaAhbhCXR4BFE8t2/+4j
Lg1ZcxPNMX4DG1sKiqjSyv8sINqS2VRylGv5s2gOO4CauS5oNT15lA7/JLCDhyFb
urc0kpw7a2iDokj7uLBujGT9JPfcZJY3AsZKDKxLPLoeN9HK3kSzYbbhh8wnVfLl
ajLfp8B8rRLNUcj145O+HkDuPJrVcmK80dmmXhNKowmcRQ/J/TUG/FHjZm4nMa8k
Dig5kVa2v+92z/HVuyRbpGNSWnrYqLOmLBiV66pvm7zKt+wtbavXBI/AyqZt19zL
1ZqtgODP+8AMP057c0O2Y62cfXBvl1VgdvT1jkDH0vQSEdGvD++gWhvUF+yV2a+c
gTGjWEcLaAhnvNVvGFc5mcv+e2BmpJCaqwJor4q1KqMXAPWEQAHzCQMt0k/SNZCh
7AndFJhA3qJZLZPZfZZhmeg2DolJGNUCn2WG4OfbSyDUEESYNc4Jv/WQPHXu+hqi
3anYsNAegzgpPS2zG0jkjoNonUaEET+EC4DHzkYm5oSLsofrb3zZBsCKubUFvUu7
M0mLxAtBjTn3Idguap5yVLpfz6/FJdBlPLgE3V81fb+VtKFy9IrKrusnowhtSlfv
beVevsF3ZowUhxXVKqq6sII1SCa9skmdosTP+PvgYlrzw3qYcI82C3jqbOHbSO1/
NAJwk0TsnsMqdgsFwcxT1YELJQticce/yJjK0vh5NSbyQ0/0JsXI9omd0jlxwg8b
+2hxrUWXRrbss3SKhKAE3SnD1G4dJZ+CjVKhworC72HkXPA+uT0r609ZTwwG0DdJ
cAG/wgRzcBgZcvqWQSZzCTCpOEFuiSyqk9TM/RkMs5kyjjBeFT+Q92GpMgYD9SLk
Nzk6BOsyGpqDZNhVwqlk89gbZX5lmk4Gh5jeMl1PSt95MX8IbdlhfKPKCTJN/3hE
ejBFd3CK1Be/XYqPbudsyyeRJo5XyA0BFQt8uMxcpUaS6RGun4KkfPTkoE9lH0cT
pQrLoKcOdApw4HtARwYIUwlmxi+W336LjHCHrHaQPdWl0CcakVZ0fQcWPvZEpv84
6g10H9mRwoYo+HcQ30sCQcTR5h51FZhqDRg8i9raPeE25kcomb9ZAJ3Eh9bSvZrV
i5ys2lWo3mic+IQZu4NJcghSM8KtFDpxMw+JgBQjEUlD5SEfKuaPjCUJ8F3kAynx
x8u+NB3JvGy1mUryolccTjgfxpDkigR7kyYDiCUDiBuYBUKl6MHV9j50HfojZ/7K
L+AfDpR72csyWtXLxfBb3uAT6WJtbW1UgLk53S4+I8pFoJb/7NhGG07c3oCykrdw
FRajvtMhRZoWC7ZVjx9zC41Pdymmw8Zhc0ZB5xKX5GqsLRHd4daD5dL+XdHSaVdn
2oOruD5NbO1a/TUdqQSS70SB3iz4CQRdDRZMCMEP/4lywL/sguVMAQcqqdR7k2Kp
KJwDeE5VKMDUmBsFJwFGcCxTMuLFjocvE+8OSNCp9kz8FQhHsbNMZOQVzwRzKg4U
cXhYMYU6mkWMZLXLgBseNTPLO6e8MQyAymdDMgITLbHnv1tlE3m1QcCRL9cGOIy2
wD3bNo1Hj5HzsUxN2xoSJkoZfQOlnoiWpc6BKySdj91yNdNe/+Qh1h/cb6kRAaAW
nbQo7QPsdgVJtXkw5rAHeySl9g3FNOIzsZauAXrV40Uw0YWHU6KDRj4qR2JxxZ34
468vn47L+hl0w19apTdyA1gqVigxxJAmmNKFDNNlJ4GJjM73ZA9y0oPAwbCbANLl
zGlxESMlYLJWWrNXCElWX+bRq/Q5k4Ejds2kQjjWEMEr6VRS+ulRUNPj3fte0fJD
jdtNXrYnjdmtM1LQZur8Q9dI3i2ajZ3jaOmdP+u6MYLorgCwmOYk7srTXFmxIziL
BkumDJSNhpB7hP0AIMrkSsusgJdTAk7mEUksPHRz67xo9wpZoCDaOejqBzxO+PKr
di6odZbSUuedlK3iEUb/+TeHfW05/kv03XO2dnvZ0Wxu46ek93vBLIiDYkfE6o9Z
euDeKmabmeDsFwZ0kOick4Vnd8DwOJB/mB0sOltVktbUlOT9dKqRW7gt/HCC/jhB
`protect END_PROTECTED
