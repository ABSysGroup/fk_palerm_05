`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n/5LHoRNCD8ZAxzIBX7+FoGnjEbmSS240yY2sfd2AvVh59asiTboY3RYZiXTv6vi
VuwIuhcFGhp0ViFfRWCCpg0turuGwjzS6w/SoNYguFH+B0MAHDH8UBBdNZtvFQJ0
bqB9k6uNS+sgm1ZlgH138lJM8zBOpozWY6pm0wsIyfKE2QYWYPfE3u/tT1/7ADGV
gOzWT+mPOiJgOr3vGi4zaQU/NjH87rrrZq+WkeKfzQwrY7MzSQPu+l2PudXdnqJm
aX6V/cYfIT4DOhDSSPDFzWRg46hj4qt13CNDzGbKYMx2cOZjKK7J18Q9hWlFvpmv
g7caRvNXByUmOlMCcpRlcsPXNB7HBhPiz8pdKAgDN3jF5se69Ge2Iq5sCKgM/4iX
IAxXdAndQPaCqpmASBAkT8qQrjw5BRb/YaXeebOhBmkUz9IsXv0mcYNZtLLrgBZz
HauYqlXAHP5Yn4kTt03DHrlF5/qH2JRHJnB2Itzgg7epCXlL9UAcY8mwPFaJ3F7Q
pvmONoVmb5kj2KCUgKypoV6TPnt2fa42zq8uyWENciMgRyYZsnYwiwypOpXdXm9d
HZMOQDDHtNjVF9AS86gsoUul/n9nTd/nETpX6nKtTWU0QVZPVHzzcIuqdV9JqEN9
ABLphHXTdiHGn/NLWc9s6sgG3j8zR+OHEkVXXhklkAVe0HVrwFbgUcImRhW2gp+P
LxniqiyK4kOg2zNy+SwixC9JrOYq8iWISBu4AA4OuFgi2/FynKpP1DjcEap/sCRg
pB3rDyFjVyhHRCSb61j56kQVFXm9LRQKPUoxkzXToiRxDYCjbCgl8lR/ZCv4WNz5
mZTfgw0e/PExcR9X0ipENjqubmPzvCQlpqgKRTX8mbPdZo3LV7diHZ+NFSX5jDGi
ewAltu/Y3Sn9uIlGHJEfq7buJWj8skj5TzcglA1coJQ7slQfcdZ7FaB7w0/ZIUGI
`protect END_PROTECTED
