`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nBMEQWI5PjRlL9muv6p21DGeqWcy7M/cIYoaPb0LMxFs2R8cOcan/m4+5w9w3t+9
D//2okXn9SjRf560BEiWSHR9/2BcKNxOl6zuWoTicrQ1gm27gkUrfarFhbk3DCt2
iXceQYH5/dEhkb9/dQj1gzd8EQGHr0F0ThQJ4WDFh9Ff5lPsu6VMWNIC11Z2NaYS
VnEUcx0AJjbfrHVsXzHNwPhm0l6OsJHv8K+vr/TwFaIPUof+6NXnDCDgC8KYnsoP
xMT8mDjACyWco47vj4USnkUgF+DSrECM3Twjda5u8mYZlt5iTH+KkhWB6iWd4HAf
2IQL5PzjZ8CE8a0YSHu7TkkYQh2u27wry42zVKbF6GtCYhn56fkc7vx/UZS1Y2r0
xfb+RU+ijkPX9jjBgsepqG4Ar44SAa66NtpiV0htqiITjnisr0cOfVMqcCvlmcKI
uqq5HVknLrFigiC32hYB7T3X7KzTppMzzMFu5DNXGgAyVWQn8AAqsGTBMghkvpZ6
1R5nHYW2uZFYUJuOCNeNIWPJTzC4MN7zxYFxoM4WtJLBzQZA1PoMqmwH8ywTyl9M
1rYbg7Lc3uoHKya+4Y+nu32h2uVzSiGuytVnevZIwdB7rcURLoi0lwyILczQRl+P
tfj3cbyed8aVgiA1c4CkBb1wKe4e1vW+4bm2v0KEadNPMwYVN8Us4OuuzBQOEwh8
C541PIdP/TFEDxKokquuNzDmRs+pwikKWBn8pxua2bAY4B/K81EWDJ07I0syciU4
1BYcjgj+xBAKD14H5LWfm0lxUXtJUyq83arbUKEJQIM=
`protect END_PROTECTED
