`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VETUh4+17ZCBWK4DljCsp93PFNe0d48Rc7T8qVuRG1rWp+HEI8xlKYcwPtXE21Bi
HqDZNlk0SdMLJtr44XiwmFZ38foQq5VnISNfqgABPP8IU0eVD3gVPTnr0etak3U7
G7pTZ0Q+heZ8KhA2fH75fGTW1DldgolBndYISTg4h1iVvkJKCGZFIfzZRCdlh6nZ
v0G32c5VRxGAqBuuGB7P21v2gAxC4bLrtMaXOyP7bxe/5FkuK2YxiGqbTJV4LU9b
EGKQbzzldEzXjc5FCgjTKkiWgzkhcr5bkXg/S3k5dmETZo84SZe/YGfTlksXXicA
ql0Xew5b22VPhJETUgVXaFK/VAtXA71XIkfSPMQgjih8uB6bGADhMIeVM3HJ/Ea1
5ez4UHbRn5za7JEt9XAw+C9v4wH9w+J8arpygQyXH3nCzYtl6m1HAybPoQj0gzrl
wY8bGLOIBiop/welcQxv7Wi70wuRFiKgLCe8md9iWPXULXrrWj0Vzdj3J0Kviung
lejTcnGjH4kmr5Umij303LpEzl0Y0PTo/ubodo1z40EI2JnGshORI2gytH4x9U69
1NjhIw4N5EobvRWiZEPYACQjctG3q+LpNmiJ4vh3iy9Z7hQUhuskj+bPJSIB41Hc
UQtXuR1DQuVVymq31rGSgUpXYVxbZUnlPgO75p3vxzFDZJKhIYSqnFJ/NhegLMy4
WQyxmCfEs7xRskm5sTv9efqlBmDSUoVyzZpZjv6SKoabF9M/zDDD42B1WnRchPkC
mUri1K+d3CqzSEllUqVsNfZT21Cwx53cEER7twYeBtxM3OVEJnRLprgcwLeEBTzV
6gBkzMDOql9wFdG//hgECz4AC+urZdwQwYazNuLAEaGEEUryRBM0ILJVRNKz/z+7
fO1dq9/+CO1q5YUlZjhjk6tMG8n0EqX8Y58ra/wCwgrB+QCP3BOLHwgPKf5w9T43
ruR13d0W7xl8aWZKX9hmLQ2iNUY3/gZ/rExFcjoIbh4QnG805HhmQ7NF0Z25SF9H
3WG2APgRvYvsBbPNur26d6t9jdKMipjUbpslANe0AUpvAahhJVpC8WzzVUnX4Ild
a+MQyWq7aqmUHwMrbt7wEw==
`protect END_PROTECTED
