`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OAHfTHjLB5ROcZbI5iNtSzIxPVf3rAL9dXEw5UmCAiBiJ2rINk6TGz2tvZuUvkzQ
1ue4pfzkodVn1OTPLDM//Y7q37eZCDhho1+C6kUXFgejwISSnhRZ3VIpAOXl6iO0
0ypAzropMlmAfWFxc7v42bnthhgsIglWi6DhqjOcg7KRZSby5dx5rz/ENivK+vVf
9AI0zTGJo0o9Raaokjn7vkffgMfVzceTcW8h6G11vn+YKfQhRIzVlKMGhBPID2uU
fw9Z15vwpcd0qkMQpIngvyZWNnq0UBCiFJO3sFwm/HP8Hqvvk7opppzSjyspfB9o
G0tX7mZhO07JlzSFOrHT7SwWVg+N0A9lbkMM4LR4BDli4p1bK/V7XfzHgL+QPmtS
w4EXR++3MWVeS9mGpC6qSIPNqCV0y1reteoU2dcEzOfiWklzjaRoAsgbCcpkR8ed
Rs4hR/htsSpjGse6sNfASvv7egaRtkC//02EXZvb8wwWBuU06HXPTSHjecFyX0JT
ZtZPB205io4KmTuRvU3G+W9zerCF59C8VorIlSxJGuGMvZMCT/358AqXZq6HqXtw
`protect END_PROTECTED
