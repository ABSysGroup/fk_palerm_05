`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8B1kHwQItRF9kAhaoGrv8xL5uLWKr+zoxR51G5+GEPx0vHaQuAPKsgQpnm0cn9F+
UXu6zF7/nshG2ZYN/2eKlTinbEsnEBlsuyOc7bxuOdcfgnoAlldFiRYk7wwCh/W9
o9DRs90XQCBdVwdqHQwdabc4npavTZ372K377jyCPdhjGU8+6xDvF9nDAUomBF+p
WB+8lI4HpqlF1jgOkMK/kmoSUFo5egy45NVwSs3L1b434JIvk4wM3roTx+6mcz64
sf2P0fefbPN9IEWErp2X/j9vqdl5fwm60gKRu1VUfhd7sMfncv7OquQy1Py2YlIE
Pw1qzH0SPXFjTk8j/A2MpMjr53kXWURktDEmt+q9amiPVDMUqZ9SFQC3S9SO86wf
kV0pZfrE9Gq/7gW7L5E+Ie8batEJtoIq9CAS1TeHZQGJhydtnkPJCSjtAyI6G+VA
6yNsOTvGpgmq7qWYjCk7yyhDufA8teHGn09pMWbQ4eLGmjlcbTKA1ZjTVWlXRWDs
dq0ZYLWXUva0UljIKUfccsfvle+u2vHfyo+X17xKQO7ho+LZYr32sXj9CgIvPIex
hT7NkMuPgge5+j4cb8RHE2oTBLkwftKe8G9v04kdqbE/rATvs2QEQ5wAk7vNATAL
gewQhC1v7e5wawrUP6a2RSeOocHsCyCaVjhqoKzXaSUEbHqqKuVxWCDtpkSjlmQU
1erIIniXEf9orLMDdwPZip3HvkIs39dDDxR+/HDNGOptNqjymYGLka6GbjEVG0/0
G+4B42qusFgAkuVmxkZVEGZl7CEkjO9kekmilNYMGOELKRuSflUYFY8C/Yr874ZV
10tWtp2onUpp8ZREnblPUZ/iwl8wnC2NasUQnWIBNkblvNdqAGhDq2sB9HXtjz01
qwaAKO0XM/79nRoxlNdTiC5QaRTXxpS8xukQV7mHjVhGwwiwtrXEvOl1yoivsuWU
`protect END_PROTECTED
