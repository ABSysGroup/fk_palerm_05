`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gxDpmfrkDJhrk+7Wf8IRGYh4OjBNwGCxI0bCvPssLmIzIvXbX0qEwRulYuHMyKJW
iFxcMgX2r7rQkdZsC/bAFGf60nuFeaDEdj94LR85+Cij6ziYax/OKBqZc1TN3AjJ
GijgWumL6lJAND8zC0F/y90szZ8I/8MuOgiq2DptehoQNLSIZFL/Y7QbaxPW4hng
SAopdwk2sypUetgS94W1ZJa3OG/p/UV+EBh6edCKPaJjr8euinr5x3KvdBiJsoIq
wuVY4RdmNRHCV4tJOulLuAwcMdqBmv+kz03CTV/3Cbxz+N3qwJk7bugCbiCT1lCu
QqCsoO5S9cgZ0PuMsjWX5HHjrDosheqrZQuUvA4UPtl9yPFSsU5PEMzbKpTtNOXg
e6ij0boLL41zSUiRRljYzOvplHSFGUE6XPO9KPhLotzJ5hh66zF0YOWTA38H5c4e
r7t202LxqhK//ALAi7t68kR2lbMba/wPhEcqYAs4Y7pf+NVJDacFA4nLahquaBSv
CI683M1jVsOZgVQbI+Pt2ziZltgGzVLwHDoMCgDD5HwpKlibimu+/u8+IDpyefFY
WZwH5zgKPC5GA+OFbcvVzBb36LSbZPbVcBdmgz/45hpLC436lIdLN1qXu6fQzk3A
Axsf4VdPinQZ7XBpit/exjxhd1t5jP/oKeuxt1vv/4Pcu8X6XpBsVlaaJtHrZI9U
A5p9OUYGMT98zQ3vOf6Ylc4zZLOzmoX1F4GWcLtmyzAbAMLVTXmrD/OSqpAkfazP
rxV+svSZJHZ83rGHU9EJ7L3yDkKMP1whxQchlucags8h8f8UpLkXz7eIysdqn0j8
5WQL6dE01H59FzsaHHDkivktIMp86QfI7d49Wz6sCeV2WPA+BXpZOz5t8PDw16op
zFkS25eBM3ge9/E3xYvdzEYXTVvaufx68tODDLQz6cI6+6NdlzBbUP/tT+f524hs
S9Dhwxe5kg6vWiZqvGt3ql2PHGGsxLA4NIHp74N7rtjxLzUeoi1zxiC14HbONv/B
9V2GI1PNQiU9kOV4XW5t6Po1LWFa6MoUxeyShTMWutUyrjtpDTZZZZTAg1hkxJ3x
w0yfl6PyzyazbPT8f5IMQRJCik13ayPlmARlUTHmL/1f+Ul4ruFn+he5Re1/z47B
4ycrOv0K4nzlu4h7s7Xl3nQ23kKNg9NPiaVmKyadQ3Cce5z+RgNS2Y3GNotudHba
LdzbpLBlnAjyIYRe2bBEp5kIiRenzEJjSJyw427XnPSNsv3N0D3DTIWVabSANYNY
W9B0l7sTBWBmVQGJvPz4n2OU8JQ96pm60WaGepstKMISGsxAAZUnkeyEj8956XFJ
C1UTS5nzaH7xuijuRI1LvYZU8wld0yYZURoLv5R+lQPMoleTYnDk25Yq8+DMFp95
KoGi+ypyhirBwa4/l+aSH/2J9dBpD6oYVXs0jH+x7QdPzCeBu2gqi9/wOL3NviqA
7ub2ldEQQoEPrUFtNstAJeHF44R/xw7II5euWCQLSK+q1Xv4AW2zIAdMv0DhSdiR
pPHe+iqsX4bUcAZAHZyh1rPTm9/qei5Szu6+l5/hK307BvMU0ANZteSMwAsE5rv5
lJ2sxS/iVC0K1akT5YhcySJKkp7GZqou6KKbhEhmT+1uyG60yolaWn0n/szkzZnv
Ct/fMC1Ue+us9Qx1o2zZ8pWs6hq7ge1H0RnRrqmjVXI=
`protect END_PROTECTED
