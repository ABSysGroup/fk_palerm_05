`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JWJXfsozrEyJOr0bRnpRiLh/Z3Nj5ubX38iBXDghV8O0G4OfV5Q7HRiSrRVKxspB
B/hipXMJ9tuFHmlk7eiDGK9qzealy1NDDI1FaAHYH4RZWEVn6E33XakqwGE7c5sM
KUe+YL+AdoTzHEEL9C8r8W44P61hdS+yhqvuQke1iyAG6xzRGsw92P0fPfcwA5u3
0Dtahu9+HBEnNhTiPkHf173EYSXhLQZFP9jj1sXYxI60T2KvkMc710JGwfgkRDL5
exercBjztsbigyBeNuhLsB9nJFSjQkopuTC1msmk3h6YSLJLo0gCOyoirSK3XZpz
0kwq4k4I7QTYWSpbZ1Bv3jhYSFZxWvwD3TORB/7aU6hXX5CBa/lcyyM9f344/WKc
qQS6YHd1w84DYoCl8IKD1UxFWOKOIkuIiMbx4P8k6PBZrZvOLmU0u9Jxzqynd4yu
0vFmGZSr5a1+jIhVpo5eyHuLhfqlFvDW+SGY2A/ekdY7mPmwJpuXMdAKt+PBbgbc
kyv82cmBw0WseQEVCMjU76xaLoFEH+KructgJx/bcq6crt/uM48PkMV/K0BaMHvE
Uyun6OehRmKd7a7rHRxJ9A==
`protect END_PROTECTED
