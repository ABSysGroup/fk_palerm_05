`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NVEjmfmqc+lWJtYwfpjRdrSO5CcvgARqOFrebN6cToIOBQbTBLjp+y7DXsKiV9MA
I3Fc8D0/GVyPWCHAlb5U6P/Q4yDvBbKcF8iv5BCH+MQF0MTAJ5ESGhcLmrRR+yDz
Kk6wOUyThQTmJeGfxBgGuMUNaGGeDfKJEyohxAFQZxnVZATqDEib0y/arGQRvvlP
j364AOhUs4ZYMRIIhUryiaaR742o5o+RRzJVMbRLblY7GcoPI334oNgGyFISDHtD
0liU2GczOAXc61gH3cuF0PORnKnITYu1BhKfNbpnnHYg5RwiQCqkYf0vOiEN/Pbu
1UiUVw34vCvJNDk4cr0I5ctsCnW083yGCYAsRtcSaCvNYFG85uwk5ycRvy+zPvS9
jgk0R9pM5xPNv9kcqJIuLuNKvD+LHn5rc52RN/wxvDYNFDmvmtzQ3NX1ep49pZHB
9UPXTb3KlC5h6mADr80reRIMI5M3fSR6yW/XZxwRsaKJBWyr7evpyhiG52NkKY1N
cnvgbg8QmWWr9xLt8BVS5wkTKI2Ah98pY2XyIKsSXWlIxFlyQjUZyKogc077KMGy
/fhDcH6N0YgxcLb00QfEiX2DyaiWfn1vBogMHluc9p9L5ALZr9HtrnJm+30Ewrts
/g6FKKgWWnfS48Bv6HE/UCSFpNFJXzXLyGUq6V65/bNQwU74jyH2uAQG7Ya0r8gu
JF3NAR3Q/IT/DLzMxuNA640u6my18y52FHiWAEFLS4TwwhGGMu0D5wWp7r9wwvZc
L+yY7WIIUHhdIc61QrtFTaEBK7eqI7WgF6n6sClcbqokdKGcQV4zat/XLPbErIr5
clN6wFMOk3OhN+5Vabpd45OM1c2WxiY4sBkmlUgb3ZSuc315duKlcLzRRKvLlpJx
zpn1XwibaDT0AZR6TVTg2Ye1hVBrWbBHkZB0PGLbzDjJW4+vlsGh7b1aXrnwa6PD
Vt1nzAY9Re2qz9gc/m7p92tLQR5uVLeJGWLS0G48M+Ulk6EDk1z5yYGgjkkreo5S
A4z44BFnm2q414B3/1Td+yBXYV2DrUFRImpdHxcYqYkN/eziDnBqobKkdjwg3skd
Nq8K+Ht/+nhvnQ4z6XST9rDDXlhxB3SQtg+PAB9Md4CHP6HtgKLVNU9ave1d6UsR
haljIC4QkcJGfarDP3aS9X1ow5S6npXR1tU7k1aAH+uk+9adb19j5m/w03vQxr7/
70gyMuzQDDsriKqRdIjWU25Ew+RDOtjQiI9B8uDvqQX1EMm/84BFyP7gHO4LoYFK
kAPo/7r7vwAKZWqZB1C85Sscftft2ZZr+YCl8bdd7TPLKG4jpZHRHPcvVC8r8WG4
ZgebFdqMLPnV+7YlJFTIDrq5FupB/n/z70q9ZzMB7+Ct4rxmu/POcU6ovMLpnYpc
bs8d9bILrMUlrBCpRMBmWscuNvCqfry6zAJJjWXY5+I/O3PIY5Gmw9Xrp4ljsHY4
0xRpNqI/aaNi7i1zjRe1MmlOVG5d7QX/ohAD5HC67PRPXAeiW14QIz4kpLov7w6g
jcQBO1Pi3BK/fgKQqBrkC/aTweKVYVBlA37EIPmb3jBIvOZ1ACV9pzpTXtoo2lmD
/FFoSzR7wwibe1Bpze+IStBI7Sx9prIzhYEoPTnzbCyFABxm3dxPpdMBuSytTgsh
7zNTrimqfvG1x0VKb3VxHkgq2g2X+rHgLkkgQxJ7EStCre8Z965HwLu8rQZoOpo4
ewxWKu8ddRYEUSANipjxffz7rggzZQmwdIplU7A+xp0=
`protect END_PROTECTED
