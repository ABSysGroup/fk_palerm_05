`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zt6eZ0d2SIFFYAc32h1so3iG3uf/VT+UXJua+cUjuHB6OP31R5KUgzCWNbjhpEhZ
XBDgjRr9By5Vy2TAlbDPi9abLH9Zgg0swAuqy5BMHsBgrkDBgqsm7KoNhOVk8ZgA
o55EMgSksy6aetUC6QvcfXdp7kDpuIoDYfr/prBKbcrn1tL2uu050NPEWm7BzdKJ
6Myw/UFOSHAAcbPi8CUZwY+x5/Lej+g9R+N5GIOLhUBRyOXK5b5uPKLEEWEi00OT
H0DJiZd2eqVTHuHDEEcuG+nHNcpXh/eRQlEKuIrpRh/pyunD3ptO9GTCasf1jiag
FV8W32Sib2Sd13JRG5/l/Z/oFDJKeajJ+R8JQZlsRWmw04EGzG6X7e/mvjzkdkuf
L21Yf2Ga4an3h7TKyckATTfDQ9l1dITrp4IbiPyJ83O9dOEODaw+tKi5mOhxVma1
774bfzUzZGXXd29PXDq0K14oVw0sMkvwMxhHsSUJGnZ0y7iLaCD+aZK5QTn+n81P
U+8wi7aUc8M7x7WCrZCY2jsYIs8QBMB4mQhwd87386oDoGZNtaonF0h5mmu5qaV/
W25PGP5Isf6raLp6gbwLx3npoTaQrhZKHE5qZsM2F/hVh7vfgwsA/8ka33O4uwNG
+4iUxouJjFwoSi2pVbonRYxsX3gT/wdZynMfZJs7ypw=
`protect END_PROTECTED
