`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tyQbmtEvGFFux0rwyh++t/Qoet2/fHP5zcfCKd7zL/1FdmQlkAK2CxhqpjHcpP+9
yeDwKSt8zDTugO2KpfqQL3D8bpDaA7qQku/lOGi33a6y5F2Enm4F2LVNuNIMQdJr
eAsWpaAhGkHcta3vw/oOGFWnblVWMpZX6Sj2dr6ysuZCOEEdjK7cLfBElkOlh6cT
RR7RYxcGpuNBBItSUxfCMD80IZsC4EDs7p8PEkJx4sdTSwLo6fRgs/jEx6tc2KCy
+zIzcw08UDe+vNS6KoE9sOSQ6JTEQHt94cWbyJSQ+nM=
`protect END_PROTECTED
