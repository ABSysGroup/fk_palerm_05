`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VmHxf7mIXemDT5nNFc29/gXJ+pzWkvzOK+MJL5EeqnA8lDXoA9x5OgOyB7NrF6QV
UO4a9N1jfJ69rMGT+Ng1BiS/IaTbEX/A+DlvMcYW2H8cLXt24GS1DRODnry1tbxK
U85F2449tTyHvh99Oq5gSwPkJs/G1VBQyX+zv7xuskhDHoOA+weFS0JFtzSoRlKr
PK+c6QUbX8qK6OV1eGTZHl95JCrQ3KxDf69N1gBs00ggw9j4FIxtWKaG+z7FgUCs
ZziMc5A18dTwvjIjCjTbZudxmsujowvPMvJUZmdev/Eg4DjEvujVNp+f9wayunOc
npL+DboLK7/wv6NQM83b7vE4Cl1Oipx2f4JFaiyODWRCWssSvoIGN7PKqmj73114
UptcP2UEGbnIG1CMuXhMKgIWY+tvcwVT/SwBl8KDDUliwwlj9G360GuNm5TREIL3
DrrgflkHu2LMxHZ8HMOlcUhO0oq/XxbhdOD9twEySTPImSZSP8pu8ufBFYRERafG
eIoQGvRadeWwYkDF2TFyjsaurbCO68SRsws4o8VyRqQIU1ZG81J02J4MNoP7hruf
jMhWXaNzA/iQJsAh378+N5NhD8k28d2UhfZj9Q4nJkYZrWVoAV1SeOBGx2CiCwRy
rFSXP5l/QLQETZfis2t2meqkYOsPwZoyK3ch5CkrPgqAKKg6YTETjgrnhHcNQmYK
qKAzVSXEp+r+hm7KWWyiaGRO94gmZMW1FOdhRRhJzfFXmc91J2cJttl42bwTFfxS
RZ/UCEiUQbtOcipXJHjIlniRE18pQaIdm063NolOfBVEnlhNENpmiiYZWtvIpDRX
aqVuNC4Xn2vb8ekZbJxDiuF3ww+6ZUekP1dl2GWnucOYwUPC2BvC1Kyu6pKnpCq8
FQQVNjWpg6cvR0QGpYC4k/sLKRv81GsNlmhyVOI+QFkQxgEep7kCIQuAx0ZqEPEr
SOpNLN6EEtN9FfHk8yKpBtXmbQ8ItCaYJzAAgSqjz1Ems9a8w1Cc0GxLinNpYxdj
qxPHcnhQY8ujj5+zsyFKUdD1sO7zYMFc+ptUylTpL/XvZ1fE0f26ADgzbc6MXNH1
QL/UCbJIgQlxnlTMyTu/SvHOEMtaADm14hWgzxBQz3lZSU032x89T2q9jTXTz0+/
RvRdr9W2xjCTzLYLu7JfFHqVv5bqetgxkHZ04IrE4seJoEVxKcN4VuKL5UHCm6zE
L5EWGOVnLG/IgSV5IyrPwyXA7X6F16yHPP90nHVwBlM=
`protect END_PROTECTED
