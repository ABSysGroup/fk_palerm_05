`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WTrFlE6cmuFg4sTybMLAUWghUxfASCWZXh4ry694PvbKXoM59MIdcxuIinaij2Wd
B0f3hrlFh5r8Np8K5xtjBlHtejLNsUA2xBIqV8uazcgl0IBBwiSa/2xoSK+rroPE
fvH4tvCdh8eLl+/m7Zd6jf07fINkwGaxxJ46gjQlELK48y1hSF10+Lf/Ywz+X9BR
8AlXv+cJhUwaPhbfpUa8RH2P88yd+TCDxSpXZl2yXRNDYDutWYpoa/k/j8UyDgvf
1aT0wSeTnuLvbx5rt5kFvzWtkFUKt0JbQVPlDU6G5ALm/MhL/8s8wNhWggkjgiR3
iQwhOj/7wBkzrGYYHP2Lzuo/BuSfm5j6TrLHQAC0TSl7T+qyqCzwUNDQhgoaMO/S
/Nk23SN6rb7hSX0x3eTVstgFn8KpRgUsNH4k+NAwGJyDQwBIqtKzkzK6gtd1X7Qa
6h+w3dAR6BRbv6Kk01X7c/vNThkWnomWYl2na2Spe6quS+n1eoe8Ywye4Icd/xtT
Ncrd29H6DD7agWwviv8Pa29WH9u8/PgyrKPe8RxyrD/2ilsqpQYz/Q+C7If7MmRM
fcdAMKoLfY31e0lfgoqrPNDP1FK7MQK5hOUN4Ff3HrjQYRldnJrhlrf0HtZzcRCf
saXTNxahXSmuFlZneiLMOmf1vuzGcHn5aoDloT7NCkc3GQrN/c/T++NrmtZK4x+d
AkuvaaK8ohLrvvZJgmisS3AY8voXbJZP5yY3bdTZHA5Or+kjpVwv6xZ3zxZzDwjs
VESWqVMyFpewUW5kpyTJ1dHrTQZux6tqbonP+QhVThtARl/tnlcU+Yz4unQJARLJ
gFXCWfPVOmy/pMhURiJV7qoBRcU5ApGiRFIvoQjQqW6JkyoxSe6Wutfzujmrga0x
CxPzMoAYz9++4uzNv1HTAPVGaXHoGO/dabNLAm4sRPUxPAR6bAVB6E1WI6nIR5Bo
/2O7QC1BypBs7PHr/6kjibwOMTz/IRBZKlfwlaoz1QbAviodiy8FZVLgERWv8Adf
Z7gRXW990mgTkTIPcDYsKfTMH5Wf4QJ60Gb7VcqC+JRbUVCT+qQzQGVqmYZxf7tO
SbsdYhWPkdXjZFyihX9c6NcTbH7XBMH8uHkghE3IMF0hmabzf14kliqMprKJnIjY
`protect END_PROTECTED
