`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
88shTw6W+Qa2V6KQl1zSCQNEExEWSpXK26HTlY5YPVg8O4Z3BLZw9E0I1k7sITRj
X/hCb0lM9kktp1Q/FfpiUgRNn7o6bsUuPqeoNsUvqIuke2eWcTRUsml2DJIjwCiF
1LEqui/6SABP+PcZVY5OutwZ6jgrjuVxqF+I4xLUoS4w/S1F29Os0UWRkhsQUGXZ
w8SWiYZl+nO3zQEWpEW5mbm5q39TkUhm0GkQaJ3aUGutx9j6OqcT52+7wRpPOjQf
hzTYj5OMcfIoaaWZYEkzqJiYuoAN3qGM1dm5K2mIOPCFjg+zQv+lHvM1CXk2B4XE
3aU9t+vCfGv3AFKRRR0zdABFUEFXeYDxc+EJ+Rah/rgHw9jnbYsxDlQduDQ8ZE4I
LxSBmD1QoHgPM4QAeERYZul6HDFbi7fxx+TLv1pTRE7P8HEuRPAjUUbMqh2ukBe9
B7QSxuc2gypT6Yt+4nBgSNWYaDdt/taKFyOFc6jLHDEMsxyo/7EGGVl3VT+VyDqd
sMSXz7jRM7Y9Wv94Lh4jf92pEKuIJRRcsdaiDweRJNkpoBXjXUXyAFhQV++RNzre
7/y3+6po4YQQ7/xU1sY7wKj7lxDCKYz1kYOl3FLmDHfKHlE4ugIz9P027caJ2QVv
4bZlWYKn8wj79LAF7EBAf646mo2f9NxCd01tvKNpwBNsN7bavJCsPgZ7O/cxAJJX
dhP8W2rtsAPWoZyjm35f8ZUIjJi+39WjdPEBUgAT7IsvbUWPyZRNEagNqsmM4Pli
sqM9izEBCr8Rj3erAB6q+xRm/Y7QaPytFzDmeW4bLtE=
`protect END_PROTECTED
