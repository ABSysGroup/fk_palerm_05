`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S796Gs5TLwrJcDzU6l1C9XCPn3kPE8I4Hg8jZstM4OKK/W3lqHRSm3otiQznVGMP
CWzH10jjCNrRkBPQe/8ZKrhAlX5nuIxMIwOGQk8DP2RVa8LnmHOnBTGE4urJwwcH
EJ323ZoACgyEdYNPGqXwaTCqVlNW5go4iKsszLfuYrkMqkyJsJN/FgWphQKOfrPx
ekHVmXU5fKpo3QI90zwmPHQ8J96OtrlRQphwkZFiwscAvcph5MaeuzRFTg7WSQeI
ugxaFdze610kY6kb2oiqFkBFy7JeUvsVLArJ8Pt/CYPjsARSAq8V3ulc6RzcQJdN
pAeNfc/uc7ePud++V1T61IGk4794A8xhZTDKd3thOJk=
`protect END_PROTECTED
