`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q5l3f70NfNpBeufnIIrV5DO6fSuufFdQ8rqa+li4wPtLwJr4Y1gS+wFngoyrCtd4
WXN/7gJaD2m/bSrMUs1l2hunpj6Fpn0/sQXbC6+ge2szB1Hv2f2/JiTBACFGoPQd
GBmFOitQTI2MNp1MnSmG5CBKc4/WZZT5LtBjN7P553hSue8Kl3dvZWw5hzg8ACOr
6rjPj2Vv2gJRxeDrzzhUye3qRkWAqccrybJ/xg+lSNGavNnMcEvVe3QqOYqf0r49
/hBqSn1b3t8TcKLKRjs3w1RrsKRHJcmqJXif5eSMH10c+VOtidQU0PDsZ20NCY0r
3dACF2Q5MrGTbBpYvCYx0xFhknXARjunLGTr4jdjWnLEBmyUaRuOswA4X5Op7dWU
OoKRCiiFvO8Nhyh5LUl/+m4G4+CeOgJyaHj5mSBXoSqKKQJHhGjBNuIADjx9JBAR
mVBl0jdIbcj0qSrp4lDKQAFP3fZLjK1tZvgWfD2NHt+GAvZizX5+kHPA0nfzZDnR
uGeTwUukXLXHsl1tabt48/E4GiNuPaJFhxozyl15VtkIRbciEVG7xH0uuUWqsQ6D
tRGwCJ94c1h7ICigwSEmAicssPRRZgNKwNtYP3Ig1url/NikorFd53Itx0xPdKJ3
lWm7r8U8WE5SsEnDduSEqb2bXb2HSrPhjOURjFPLrlJ09bP1sPfK6hhTtuXC6IUX
M+ADoVkw2huxcM9Td/NiNC5umajR3XE7y4W6QYT1D7eTR/e2Twy5arA0hRO2GaBW
8G+ga9i12GJZOn+3tSx5oQww0Z+EjuF4j6ivI0ILYCBdVqfkBnr8iFj4kmceabEV
u4lKWSXE2jWa1IOFL1FrwpXUn/oKoqHt150iWVVYoGEjbgHzGQSpwCfI7uxG/STm
KispsT644KaFmA8ujqJ4WJPEwJITT6CJ1P/Pme+D5M3SXAmr08d04/SARXZ+5y7Z
i5aieTYRqyVM+0wjPohaCq8MAGPDY72edjHklOQ5MI2EEXjc4IxFfRWAh13rdX+V
lD5Gj/xGmycpkazJLpG+bQiQSiKXGPb0uyde7oL5wVQB0V4S4hO0fFDd4+AD3cmw
DysLqzCO9jHhmgMeGTacaQqEVw7bTFbuIGtbiDCzcL92LL78dHJKHyQG09E1N7+i
obxIhFEes3ZTTJLvzzj21GE7YrN3nb3ALbDcPtdGzWU/vTpZQrCH89pnXksaUiXL
NNGOR6Zz/C+sDCcMiMn30rNI7m3c1p0Nh2VClLAZHoxwOtWai8cWATdkjrKis4Do
PyiKJQsm66x48qB+P/85BbQP+sZAXhUxMLy8pJtmVcgll4Oqh1rk7KV2y68ckHIP
t0qOdBVW+YBvJHnQeh6yrJOxNdTkw96Hlm5oc9QlYyGMfjmGbAquq9UwQsgoEBmK
`protect END_PROTECTED
