`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i2ktR+MIEth0IcUfBrXTzt09KN5J6f3Q6nokyZiWh/V6Ok2GapkSRT8s2vHkOMjw
y7cfDauf5teSY0DX8O5EEW4N/stK3TP/TLahfFUQJmRQTspu0v6m5zJVEDRTV61x
Y6mh9wxSJYD5wHV1+HwHJ2r8zYsiKEmuTpWuwZFhSm3mavB1BFIMfxrDtZqDzphq
MANSY6/eIT0Q81IZpDia9jRuu561lEUcbq4igUGxSlBnN8EMsgBezb3rDz7EcBbo
eZRPyXVN18I1ylJNe/QsDMrbyo3EJ+LAHv7vBtqU+zY8WrDCwAnWGCM04IEtCGo/
1F5S5lzWRwJbzMfZjNR8xTKmHRZgvM5xZu0aHfjXSgAZlr4DMiD+B+KvmeKdk0Tj
373z3+xdljs7gi7IMkMIY2UKBe7KEZyM5DZkd0r3Cx8=
`protect END_PROTECTED
