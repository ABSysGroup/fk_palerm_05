`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6knOLs0pQeEMa0gsD+S4xp3iF2v77bxHt3KA+pZrCg5qGsA+l7ZO0+wIA39bx27V
cXZH1nN/IQNqcePJjGd7831gclNqre/wIDnaTMcLthHXfpRzAoRZUeyDask6yQ6E
c5CA0ufoz+eqpgRm4/b5lplT0YNPDRF9S1/8Yw1InuKxrqw//mOHZf5ZAP1NZ5lN
4kDTwclV8p+n7s0aeBjcgf23rRgHrukk7O8RXqOXVV1Z0WGQDjYYH1rsi9AdJYKC
dP2lbC9ZF+stvKpHJI3dslXAUM55+XHuW219xUHR4vfXMhoWli8NtMktnLyDFN1Y
WbJC3VMoFoW/m7syOmD41LBpN5h9j1lLwaooyxtPCsLRryJiw15RS6BtVXs8CE+H
EQbOW5oCIgb33WCPdUSoZgvV3TguxkDi6pCxRABZLgcC5TSobzYVLsaGd0BH1urO
uwt3OzhUUpsoSo89sTGpcKVYaCIOSIwXVp8dSCmzcsOqrhOcgKQ12zmThmuxSyd2
vaqHhQETWGDhScFLaocDjr43PdYOyXHDwU9JzJrYXwWPuRweltJJLi2l99VolzCI
QIDphWxete331W5CtsqXUW1hlTemvye35midq68UBB3SQtyHKtptfQkZMCWpKEXm
YklN6IHsn6YjdBJ3SGQjh3qoOZ26gP6I9EIdW0XijoTamOYHBNWlRw7L4/0RYSTR
9Fjv14L+bZiG8tmp3yajhtJ4Pf4UQFRbwdsshnZa2wsZXANwMuqJcNEC4oLdRR5r
aYUbTl3ekGAwxndbbgL4aNAAnDm1p9y7gbsqtEavx33pmty79WnCWeyBmvnutq++
gE2MIIvi5+f0qXwoSxEHoKRRuqU9KIMTOJreKy2GBHY=
`protect END_PROTECTED
