`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ykMU0PC5Z3VTdqDwT2ryuUWT0pz6we9B9BsW1nBwQNvh1t2ujb5Af2lzo5bE9R/S
+uKLRbdrsIorlDLU2EKSLDe4nvYvpRsKkQxdFS9iooxCu9HZdqemdHSm83uuEe1P
MtoiZ6c65F1/bRIcA8OHH9esWC4YSsL/YXHLUHCsj39JA0/Dh+A9WNEioF8MsQhH
n0UA6ZOqOLQyCXHcfV3l9WgF2wpEItFmQ1KDrZTfAIf/t9YbWOoUJH4Y5CCorRfD
6Brr4kAGasgVXueLPWAlQEwU8eY8ZUaeoDS3EHctzeW1wAoxI6sZp26BEUi6pC2o
PAaZ7dJ7HkTKSg90jM1FMrjndO0tN1NP7qj+30KKQp2aplHCqlZsOP5aXQblVbxE
waZ+YD+7Ze6WCzMBOsuVZID98+rtNZxIf9iqXUPKwTwJo3TlRfeJHf/xXBFtQQH2
ppHw+mCNh+vGHYBs5nIV+PFhLdonic8eZi8Gbq53FZE=
`protect END_PROTECTED
