`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V27ZFVeUsZvbGA4LTi2EA/D45oNzy1uf/lp+vY2mrCtbUsbaRi3DldVWvv0VMKhP
F0oDCwL7pNd/LsTpemF5wEG/i6X2JywsUnTgAtRqoyOh+1FTQobczxavubXbT2gg
likwnkXZU4hMSiYlU5/GxW1rLaBF5n8GLfYv69DOpxxgFmK79YQowA5/b/4bE7UV
5l9Qajdv37xMe4fZTwiibrFD1h4BvPc009OA7UGfQ7UTPb16DDk4gw8QVpiqFp2R
sLOqNuB6lEaVF+SZ50YLsHU6QLG68yrO1DZb3DiUE6hzU2KATDGBtvq78ogNMVsB
UjpBRHG+8x3Od1Yhptyc7gDBp2AL4talhdlnaUs0M7NagdhhHUIk79hpjORlyZt+
v/us9cLhVYzw3FR2e5xkLhBsHNs0AQ2eQhLwzNRtFZ73UxKv6k6Wo90YHE3TU/ro
2x/N4fMedIyZZybICrGvOv0cm/3ILHxc74M6okjccd1WAEtNZTMyrXqPyf0s1Oe7
q77ha2Y+q8TfqZUXp1tucdqKPudkHUWErKZcNNVYqmfxNF0Lw3CaZ0CoJpWZJrap
2ET+QlaPDSWZOa17kqFUa0G3b0sNYc1yxJaMmim8dR7P0cuzVeJogjP4Fr9b6ldB
XRrtjbaiZZQxOSqFaNSMFw==
`protect END_PROTECTED
