`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NEwltpudPkB9PtCUg/dwRL3eBlNR4MvunPPyi32Rt6OZDRs8z/tr4O7s9H2UyPf1
8G983UqXpPpKO7Ol5qbzTWPT0I07JHnIQPhvSFVNWC5NJC/ry+WwLrCV2CVCJs+U
rDuD+iRzGGFWXmN58sDcKnfSBHJqO7C7g3UUJn/b4KUNR+cSznWksTCtcqLkQF19
fmmxr17cO4iek95id1O/JtfofzUFdoyHXmFhgTEAsdB6C3+NUQkZ3kQJVIYQkkiV
Xa2rLdqdTlYu2N+G9BRZDBRCZqfoqKpsIrsVYnrstbwtKWpG/Ub8vxTN17iPDKa3
Gf19VKoNpa4ntqRpi2WX3A==
`protect END_PROTECTED
