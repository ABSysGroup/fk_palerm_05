`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QYpIo29Y9iol2Yo1RXNmzQq5Z31wl6LvaucK1XN/ZJ1KKxMZ2nrokOS8eY08GNCA
URgs0e7kI8IcQOpvfecxesX0eFvd+OJfiHUkfrNDWoTkNn1o6+nzzvR+vmLHNOKP
DKYnNos/uIx4CkT35qjCebF6Jaysi2TggDwHGOT/ZIe6kOR8g2VM6bY3YzbTktA6
wc90JRQXD1mTwWDpjVn48zwY3g6XXzd2aR0sTK1yVCvIkwuIAbtY7nz1D+GYLkEA
qhImD7Rwm4X6jjyHaxAGJ2182tIzbG7rUN8DNG4U58g=
`protect END_PROTECTED
