`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BLecwDiacDNr1H1X7DsxJD/jyspbbNq4CGm4PTwA5pzbIu7SAjBxvye1CAT7HVUU
ulZ/9xHAWzfAPjPKeP/gLgDESQn0q5b4mXIBEYzVQe778jaowv2Pxd22E65Dbk6q
b9UFz9XfCNO0O1eYlBLvw90VfLBJR1ZBSlJDm0uV8R/PFNr35JFa2/+mMsWLBrk9
euM8prZVsCoqPE9sAR0S/wc0nzCMxHe15R7ETHSaa0POBXtG3H4/oj+NwuUw/zKJ
E4M4h0GRMv99T5l3mdJjjtly2i3bdu2VbIYlVVz7AZ856v/U1HLrF0k44G/Vbe1E
Tc70fmACwbcoLOo6xsJXsCd2tpoN/SS6sBItPtwNbVOG7cEGT7EYKpmHre+c8CDS
+qyj69s2x55ZKGMg4CDjut9DULr3LPJfj0j9mmagrah7QdFsgaaNMbH9rcJViTma
04I4gj2V6U1IXNPF9cncpcglALw8MPm55kqLtwYoffOdP60P/owXJTDLhM1xNh7P
uGslYhSfJJJWvkZwl0PRfhREqVv2V/yvhSxB0j6UYaUUys26oOT309utdoQaYqNq
8YxGwC/6u3ubynSVNyZrtNb7rbG3+YtKMelet5ugJ0NJ751E1XyOiJVRpEmJR29U
`protect END_PROTECTED
