`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QcD708cG/Ufm7danGwDB2EAz4elJW7cMoJqLq2d4yjEJQLr4JkqnhDqJHy/R+RH/
40+e0l5nuWitnknLC/EMKDYHLHjckqwSviDwVRG6RRT5AJwtijzrnycemdOFlqql
KhWYFysiqtxyZrhQSEmA9mon73FdA3bAM3wdpHPSxg5ySrwMmBAKA/Cnr28hoa/2
0Yl0GEyBqCV0FaVehNJc5cY9itTWrS5PVDGSkVtUGNdyee5nLoGOVxHSKuBX69H5
H9IRGnO3uzYDwpOr6GYl24z78JvSfp6HMD1tc7D75iB2OS8rbPzUYLHUmGDNY176
NushdhFlMQf7ywVkkApPE58s8Z3Vi7r8Z8B7BStoHJ+nJz/RkUYEBkR1a/DN1jSa
2w/CPfWjx+l4EKbi/+yiIKYyTT3Fuh3O5xfovmq1yKN2XK8VUMkliLWA+ciDsEZE
pzFm0d35HW2g6W8WdyD6w/8E/u2/bw1GXGAKnWRGcdUYZGVVi+Lz+GWZQq+N476q
s/07V/vnIV0/OW91I9dQN0wGV3Qlw5oQxLBxIbuu08ZQbzpslwHij3rRq723vOln
`protect END_PROTECTED
