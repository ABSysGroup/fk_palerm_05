`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8SO6wd6/arKyYhMPEvgaCd8FW2SYGHcwHrV+Lpm0FIn11P4PYiy5NvT/79dySxWN
OEgejvfj30e57hV3rx3r0j1EdxBTlZiJAdxk0SPO+taRiJyDw/DKJdwbtsa+8wcX
xQkZ/ublgt/VGeZ7QQC0VVNAYBf8hFGVaYOSDrD7jzYNd+HIRLGPifXhiSDzwigp
yX9I3aeQkM6+TQEUm52K4MTa1gRx6oXPmsmTsKFry93ZFvViM7ittFlZSVNgCb9Y
GktCR4OhbafE5hbcSRQiCH30H+h8H8jdInqI1KX97ogUILiWfEki5WlnogJI0uQR
cabt6I405Jt0WrsDp0Y9WetdaZ1jRN6lnjXrQ7yACGY/Jqd/ZRZSV8hKswmEfoNP
xYREgZV7uxMMJ0YjZLO6k2hxMfjiUT97rv6iSgMNvDWMbkflovCbRKu3T4GdJV5Q
boh3RbYc2JHftOxfdktb7dGqP7BPEejerL7UkzjNJ4SRlz5woKbetXdKHwtPtaTu
wijhQeBzPKbmYf0ukYJ1vkR1hFFOUc9HO/dFIBcm6RjEbC5SWkg+m/SJnbMRupnr
5hww6qC0zAHKmaW5qLWGosmaYRI6x7Ir7U1MleZ2HFb5c1cLtG90Z8ZNgRdQrqUe
hB73v6Ryp6B2IS7xhFwwmMhwoLT2yRZkxfs2pQbQQkvYq3yJLBttvt7wwa8C4Qrc
1lJKNaD4gfbzG4xA6ls/gmczWVCRJYkEEqOXl8nW1T87oUAytUqYBYhEq8iIYIxg
aW0V4pR6wap2z+bebboUaYRvc0HYWT7X+5bxb4GBwRq/iVdIOzxAr8VCgSVhmGmA
hpOIWYaYAiK/0r7wz0NlfCABlXUs+XG3+X1fXbXv0Kv8FnlWpfs/MtwRy/aGG/vF
4GtKHVVPWVjDuDeUYayp44/6WE2ZqKlTLxGjtB1nTzsxW5gF3rU9xUAb6LvuDVXC
a7KRnuc/bZT9uygjKQOiM4+GG8oOqP+LytbGzV7KGzVAZ1Vxx0xJ0J27RY9M5Wgj
3f4hmoRWNimuAHAfQM3q9Spp4bs8uZhZF5TxoleIsi9pqR46T2Z+1VntjQmtpurN
tr1lFNFqGGFSUWw9z8gbl8tQS5pJ/P8x8XHUJgbb1wGkfCqUF/z7E76ghMI0jfhS
7RzcI6IZ6SDGNOrSqKF1yyKWavf+qfTYbUj4rIRJTBy9IULzBQ2fYBnPVrKESSzs
H4DFtlszLOgghB4aY0bN7cg7vjng7DNm2RJuMNnFdou+Hj3gezW+A1CznbdNMbTg
M0NlVOrAX+hRHZbq9FRgTC4A9lL4afCCl1cS7R6yi0FAvPY+PZeGaJHYWPc5Q3hf
pKRZJzA7jyW6wZXaERu3DymTREh9++JzWEQa4mC0HOjGUECUDiYtzc81th14vBnC
2vUK+ZdZGdPYcohYaiKW5o7X8rF4skHVLiv0fBuHe0/ulCY56jgXCMLk12AFfhPK
Tb1C+HY+CDMPwBj8fxaF5//rIPK8QJP/CFxGILf74lpcMQFjwmcHGmONlsT6RkDN
nJdUi3FkFs+V/prJKLyN3RM+I4g5smsi7JX9kAWj2xRMmYEzTfSGiVw0ZtL1pXWI
ARgVlT7MMBRiJQHhsj/2cQHyFmC9rYWXDJ8NXjh+lyFBxZEMqL8zygmofv7YJcZz
ohuV5DvUrOS5QpYCKaU4VlAFtcXURiit+ThBBxJEfETpCJ933VparHvJhgl15J2/
lrbAxi23mkx9TkPL94loRflGB6GIv/w2AvAyDq0bqo/cbHLam45mIVMa2nUgSHnm
zIir4164wF+hVJZsQ+HJvj14LT7S4WkGkE7mP6yxVFItVpXA6P9GX87vR/0JXrd9
l/KlOETGCYjx94+2YC/xick+dr/kAxnsos8byzO7a/P/A2qsedE7fZL0PQMWry5i
13o6V88nzLg9Y+nxrKepJj18OEMhfMLIxE8LvAGXZyWOe3Gt7ivKwY1oy0j9YMh/
4ZS1H3VhQ8/+vCuxKQY7qYXv3y7/lwQPReQ7yINx1XEjyG0/mDYgyNdlAmFvKDO9
0koeP2k0FxWd/od31Za8jFsppTIUzrTZjuwEdHyASpoa0NuXyMgNFtBecqOizSQh
+H6f44WnXsojEJZSvzaL3D7AIII/Ovhk9DVCzrpHGC849isA1Y8ALvHcKv19ghAn
OrFaGsoXdZ3QdwdUSB29SG4PlUFXWsBCNcZxO+hDyI/mN8VTD/O192GAf8/1wI6G
FBD+cvvFLMFL7HXa8GIsPlysA40WuJGRpbBnQEmKBI49IFoUVKFieMdh1hM40F15
uFn+l1DuV4MjcbmyLd79ae6RD1I1o4AYh1zyQYk7qh8kIks6bYNOWfF6wmGIAYoK
H144OeeMBIiy4TUjLjOigwado+r5bNsltCe5Twv/2IPDmeuZ7NsnFJLl/nFAKrCG
7p4mi5BwvdvUkuXHG+wQEt4OQkjm2Ec+pYqnGUMZUzbDCK4H3ecqkZqTh0TpncJ6
x058sa5O/2wuuvxmJ2QL5RAOI6mk0/kmu5E9sGGJN8SL5VUCBisH3xl218B9rXzq
YcBRdPDuG+sWkUv1FLLl+Esvb3Zt68pWOWyYeB89dGS8nO98gBYth9F9Szx4LHXn
DVhj69h9/vhZe10c0tmOG2ZGo8aaaSUAmHt637DaTd7HdLOPTTAmFnyCP6tVX3ph
gBm/+Png741OjH+KCjpGU/qb2MCX+3aSCklkoXmkoXU1RcU42HMxZG2TBxuNQchP
fx0PBhpaDOCoxiH08rXccsrCCyOUuc7sez73Jf967bvNGsYTLYtHl9ghvWuqfUdN
cMBa+oX42WT0p4ZrB4Vsgbki7reV6OxtN85qbhFv2wG0ikLKEYXXJM11tT/bdDAM
4fXoW/oejBjKcRA0kOl2I7G0FcyoCfUGkhNoby47LTuo+SnsKtprR0XSZX/AV32J
KXm+bViYBnAkCFKfXd/ChT6NxoJx2OCz+ybBzLWadOeiCEEE34t2sN95MefxK/4H
4qmwTBZEBASABfM9p7vyqVoqG3AAmAgUHcBt0YbTN8WMejECm2TY1qZQY3TlHrN9
OfXjy9ruuXmLDeFEOuweB1m0BWamxXOgWcAiguP6rNvHHxD6og0F8l2jyvTVS2pM
FNowSVJOM2v1ye1fXgu77sD5mZHU3nkRnTtZa8X/iIEZVroeU6RpCDwc5CiOWjPJ
ha3GTB5Zt396Dz5hcFKQ2O+1M/0he4JLf6FFqbkq/mP8t5Uruwr3mevX3gASZenW
2rNsq9cZnhSk8D7DDPBpwGF4nKThN9Ty074V/fIYL+3AWKg6epmi6PW/gdb/KJ3T
tY85hvOxV8OpKXZwmQcwuibT04cQHjelhKBqEm6di+f+bcIysYqf559ffWmOH3oZ
TIU1wUye3wD9+UR7HAmC5ygN2oCjsXFPYW2wM5kkDXNlJcEXr2SpOY1NgDdbZQQO
TEnYWs1bzNQBhJWyEAhTPmqz54t6lQrnh3lfnIMW1KT8XW+341qust922POi3IgZ
TJqcdHdVuDCuxDUDfNgPWD4tHhRuLSgrKLK4ijh6f4XTzeoLbKH3CV0cH6jWndVe
2Qd2FypaYOl3pRubGFj8jMPSmLP/nB3LAetK5+okBR7dkcswVYtCh10W1E6Y871T
iMVHNDsE+1l9SZGfU65K6WXjPtoroe1grwvXG9rooGw7jTtWzU+fIVxDbvUllMz7
r7jYxTx9gTJKcbnlRNM4paM124Np/bq5AL0b7WmjUNjkR10DAkG/3NXIAw/xmRAq
ALrsnJuM6kabEdlwLTL6scX7QEZQO4Pr44m589UD9b0h0KvHqyy5ed7XxnaI9gQ0
bwKMUbW8gC0s23Z9NSt96oVZ+SO99Jom6qPhvmE5zztfWUBRGl/sbAgo6sspmcLj
A30TgfV2DYjUH4EMmadWrtY6QZjvKgB9HM/nWq9tC6lg4n1ExUG3gkOkqzA1k/Li
RExboROl7zhf7Sf1FJ+HLXScs3vZfTfJuZ+KtVk6hXm2Og6EVjcZsxS+vI0R+orh
WC4X8WHYfSZVTwWnFL9wzX30aHTIvhJZD1htzTAP24hKzNjJ2F4xIU6Vl450fD62
9i+LecSTNvPGrAzr4iPEfknPdtIsOKqTHh80V/75/4+dyDRIe64hQ6VUiaC/t8NN
47ggwAtZR3UeOGszs3h8pKCKMvVa4/h5ZjB4/xxUphi2SHni5YxpJmHVDOTamdr2
Y33e7J/jB0m9W3dpss+IuXM295pDVWOsXOQMUnfBDYmEqY0oKsVHxeLdX8GL1aiA
1Wz2Ynl2KrtDV/rGCoeBct6+6yUJvc34MOGi4KuIAEyvkZuerOtROVrpYwQGgvNa
UHNQ2y7+Ql72xvSDmuPizTQhjugwc/YGn8jVRCTBYIhBN7HNrnlI4bqv5zpu9Yzg
bOQMBvOtPiMaU+boXyxaNruztwGh3NpN1tViFPPj8J+P1xaoz5ofX0EMLG0QEWtk
WZ1Bk/3TwPUloPEQa7XZTfsgFItzQFjgWJ2+L45tVrFOzzXmDLCpVuxRCWKl7Jeq
pUnW3Xf21kCl5zs6Zg8hSU+GL1mDxtxrN6DN8GyA9Z6E5pR2dFZ/xxQKPJB/6PlX
z9cwch0yPe3s32eOwKwwZhB+ugQma7TBFRP7QadM50sUdnN9V8fsYS6nlMUDnuS3
5aJSAvqWb+0QgI5G0SSQePnd4bL+Dp7f1yMisggWFkkKrOhDs4Zp5L2gaa+JXngw
iPLkCzs54uOPl5iZN65xAeCiTSz1rEXSBcLtE17mEqfN55zKqyLUZprXJcNFXzBZ
r+YGMwN7Vv+x/fWpuMUWE2HDcBWks8HfeK76WdHlh2Ics4j6pjazrL++lmTMetca
SwM2AswUyTlzwj2lZsHLlaGgwXy5gP8/um/GONEIdLZrHhyj5dC/JG8NVsz0LoEC
5IPAHYcki835JL3dK05z4ynYfR6tFQvyi3y/ffLIen7gMzE5lKdRDVOXsJCCPpob
zFsk/DBufwMlQ1hJRnOJM+20Hd2kh9pFnsvHZyaA8+QkFfWr/o/kVi9LKppUICY1
xiP8gv++CZMkGZzdmI229KCRvUo3GmrVAXhExmUg4XGDIKBpP4PJQ/CV7xvuhQEq
4opSzlJIO6TYnzD7Vy1qk62923DZKBOgIlv6+GdF8IorkxspE/miKh124Sou4jpW
xadztfzgjfqSJZkK/9z3Wm17dLJ6orJNanfj7nqVAn65W2D9CxZyU7JlWD7BRVFR
mn1pRbqhonfgJcaa75uzJ0FGxATU2Sf1Ik2EUe4m7m8CkjRCiafI8r5Sgmgc00r0
tQ7A7ag0jq/jmeR0kXo+UDgdPArQCMCx+U2x7Hp3ALDJ5IGNwnX2SqPe6fxOV7QF
UZHLgxBZt1wMUA4GvUJlxg3AvVh/jmzt0GczuAQHruBhjp1ZoVmgNC2ng83WWUdL
QdZRAEVd1l1gfVvem2X4/OyXSre0+f7em8o7IX9rMn/5larokA3GfPfQAzdDAivj
L/+hh3XN0jT3CxYJUUgTZ6FlE3+jgcN/jhNGkX5T5OtEGjQy3/5uE1t+lE0A4tES
A2PG+4OJNRyVnmZPgR33V5K6eEz9f4INmHOh2icBoCu47TaUmUk/tiIKowLWuhJr
XpxvuSG7RleA4oPMDMRKzSLlL8NIk3Od9d4F/7LKEtfXAg+K8q9PJZ+bP9+rMYEd
6EySeNmUThyW/vEsrbu6HNfPHc9vpWygE32nPdGYZ5iBpvcQXCuyzYJdjg6S9w60
V2ZIOKpwyrX0DXQi/Cu4eh3QseqvPKjklieXEWSgUjzZHy4tLjDWQWHei0BGRKd8
+ONkqZ6NSAJBD1P10KqdpRbm4vqqFBWCfFuInPuyYspf21IPNtnVLkEply3ejpbc
SSQVpsl7+Gz6Gbsy46lC1atDLgBIcYOuA8uY5cfZ0hkmdtxrUW1uuZkislRSTjt/
MsHpLgu0HQbwHKvqrZJ/e6e4AE1AwicmJxfGdJ8RJ5y/GtDffxeCrQ0g//SfqeTs
OO8JXAl3XcWSLlgc491aUA==
`protect END_PROTECTED
