`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yC//fmLiWg2okhwlqPdrf2Fljv68FAkJlnrkieSxXymwzwFgelEp7d++JqCblPvn
jI5Dn56WzYaUV+UTUr9TrU6t7FP9k3Gap2r9PuBhSu+X8+T3pBnTMvxCMgkvYXmd
ErAWM0V8etxNnTbldLBcOfkscOAQOFsAjqx/Z9rRbVH8WsjLAczAqeF6tjbOQNFY
YXFw/CV2FMUzkcRMQXYUCXC9TRtwUZ3dcu34S8k8eM5OCO3JWRTq4w3h9ToZrXVi
CCxy/jjyCZ5tY0R0Y8DkuA6B18sCZxTFurcqANRdQtprVOXZw5bd5yNcWWJURYOV
mOc8IMBzJeA/uqvuS8SoenRHL7XNiN7FM1CdM9QBD0RAPNKGMmsNCWvMfwicZOoG
hbb8sg90/Oob+Ybf5R074PB+bS42O1Ucw7k9Iuf+P1l947673I5oXVUHJMC2b1eJ
Sp4sbw28g8S7cTp8SvUNI42m7r4kxGKHmAK5wQWYiM3FSqN2yiHCKfeepxAB/hFQ
u9K9KGMfyN2M7tR/JT3sr+0tFS+YKgTzi7fcJQOl8Eb5hh4OrJvzh6K6CQPDSpWv
QrpzCQXlLP25V72Im96v/BECDdO1tJxvWzg+8wDp2oEAyYhjJEHVNsasRcq/qm6w
K1qPPceskoUr6JfzJrUgCc+cAB1HIyjPU7wmPhWeFphp7gWHymvj1PU43yEaMzTf
1xp588JyJI1hCYPY/ZLk8n7Cv65lvmbW7ltNZpTUM8BnmsKMhgmEKmodXHIwwjWe
X9BurAiqflp+7T68E5TSz54vA+3fj2arCatGcjc9JiJ4Qx5qbCwhQJS0p69CgSjA
k78kypk4M5+kRxR3cwHYnaSPz4nHZhnRBZqL2C4tVBuR/eLBaedRQFqHC3wE4A5O
pZqywUvaGV+6gY+Q/7AttFIEAhCprknqteX6MjEQ3Dwd8NTIXUPiyYOsXuzBGAfD
379CFPecZLAHUh9Vp+16NNjm9SeIRflDEJJk2nwJlN4llHBveQNSrVjMqfJ1FWGv
Ed1lGK8nxspl2Nh+mHOt4eM0Slp4lwBq8Jjbgz7UFjEQBSLB7R9R4aUW+49vfp1/
6UhD0zfldcECwLFckuldfl7WpJ6Ssud46U6ZEEQ7n4xWX/6WJPCJSagEJnJ5lOL3
e+wVNsaV8tOmhf60KJaDPMCvR5nnOC7btn4sMxzff1NnIuzeVBH+IWttcWUHx5hO
Db+GuAn4qaF3DC/ZtbdCeXrRgtJ0CUOUTT5pZtzeZTCcCuXmvSkVWfSgVx/wZ5eO
`protect END_PROTECTED
