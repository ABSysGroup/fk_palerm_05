`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dSmE+1AWuLdiZZ5T0c0TvjYGnIInLmTAex5HnFlbvZCs7fhidp/EHWJJZ5qq/ASd
mkqnQ/Ht5ehPrGXtuHxWSDvu5eO0+2cvLKG6ePhAxPBG3rXzsC9ga06VnnxwzkZf
oDzDgdFazJDQiFAhBG3yHnNBVLlm4K+QLbqUYe/+o2qaZebYkYCllZfxO5Ryxqsa
vry6f0WU+sKxmXPJE/2yxrLH4z59Xo5cHxt2w1YLchyxqgUBbBVestoPNSoiLxRy
DiuXfjFPtFyf+mrEWDAT9g==
`protect END_PROTECTED
