`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hp3d+kjkJz1zHY3+RtDDhuuBc4YBGfjJzq46mNYpPIyhppBNHzf/bYFcn1zJP+k9
Zu56oG2cWZs4QXjG/fsZm5M2PDz2qG4nRxk3D7PZd5j0r/hvEUODH1j1NR4wvW1v
3ppupGGdZ6UxglTOMEib/A+gkw6Ctm+Q0C/Bp10nD6BkxxfjuAuVqevOCcyR9F+P
UrWW5xLDAlb7a4Lv8XRYZ34e8nk0Opx5dwyXxNA3lzs5floG3uFlzIyLH4bJ2rQ/
USDgss8EQIWxnDPnYEnFg5QoAtOFZY6Zp5Cg1k8wE8ckhvc+G8zjDfV55qJ7rNKQ
a3cSh5EW3xbNeC048gU1TtfJSUeepFmmIoX9OE5O7YTA8pQtNaJjpU7kD2Nv+WSP
jHNgEmKEKh4Zf+tvGNqXxFhdeW4fOP+4brKG0K/0Eckopy8kMLR75+hJje1kWysM
FON08EZQYBUD133okB5f1gQIhgg6fAiH1xPrvdZnNNfdVF0NCONCzbK+O6jZN34k
K8XN/ov842FsadihDBbCGOPaR/7RZaHnx5/DqGDDQJ2LCeojBWhCRpVu+wu7820p
o7fS57UwXkYoowJtpafKtfKdJtk1eF4fWwRRap/+0NyrB7/IHy/Z7pC8viSXoLSU
`protect END_PROTECTED
