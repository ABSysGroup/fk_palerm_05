`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OhZSXw6kYvekS1Aj0g9s7CsqrRBxliMlrQL04T1UZ0WwyBHznI+nuaG0PRj5LlA8
DrVjhsqZ/dJ1/FcAvsCtEwITsDQToC2opInAcnHypoSudacahmClF9ziLJ4dA2Lo
bIyNK80lyRJD+IHEMS4C+fySRi7+XKMe3OmdjafDrLMUXFiLWBy9VSsqlqY7QXdx
B5nGxP09GyUqXlIcDkKN9dANbVzAB/yaJsA5xg4vi2PbYjVspPrYnRV05mZppuiI
MPZXnRGmkCBgYrU5MOveNE5wYX0HuPvJjPhkToz/9LlRpg899e6ytPNFaN2kmhmE
i+XR7rm/FYuYzQrJgNOiefZ8Lj1FAlt8Ct7/0Go5v7LQb7Og4pduk1LYTBHTkrO2
cScV4Aw2gM4XxQWe7K5oUOKUzA+qm+SGpMBcMiHEyoGQoUWY3BtIsVox0gaPL37s
`protect END_PROTECTED
