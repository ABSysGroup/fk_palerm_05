`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
afBQzz9FEHgFXD92AP3ggHGTjwZe7sBJlay4BUfE7oSh6TEitlqpq8VHUVTqXvU2
eF33uxFHUYZzZm2xuvdP/v4ySZp45h6Vb9jfjIJ3FoDDsPt2bDIpKwBhWI/xzbO7
w9veb6Am7VRmt2XGhcGG/Pz3iWQuIWMwPyPHFtO7znb0OcsvSZ4MIpfF43ZC9jpc
J/E6mOO0Pza17QsD4q9i6qqSGJuyOU0EP1FvO+m8yAT088WHxqtNUY52l+AIinky
CXPpaquDJaMXOPwiDpER1gve7KifLiGmqaxoLvXaCHEKS95EW0VQWGM4+L8X5cT8
Z+3B0OEK2AAQnUO/WoW+HhTwRZjM802t4w/tjDKS7Jnp0GqD8HLHaCX42nBOd99b
+TpDgmlBRYAT79b27WaNiwHBP1qkFFb9U6B1bynnDTyCvu3ji/3lcY2xrNeVmeBO
xTQ2Hbe13+N4Qr3nRKTjoJRUcUz+arh1xuljPJPhp+0MIbI48Oqj396osQL14OZ4
A2YF9aRJg2jIByF7/+4ciJi0UICDP/gL/345u2Mo5DVFlqYMxjAg57ZOWuXPxCu+
ARxIqsTa9sE2KrEpsrNSuLP5jrbYphrK+vr/0qZO2ZWdm/6moOhKJSyN54RRW5uV
ltOkCETtF7BxGVcZzT91jw5FD9Fb3Wbf+7wisPJ3/OCxJT351PArRvd2LZhLdQbX
0RuHEGz2lJXYuvOMCB9lRGIgbB7dgs6xE8N9MwSyrMKP8rv4lWTub/olC9XGfbiC
LQM5chHMYPd2ce4yPQcm8etgnmHnb8ipMRSAeUttUD1z93oDiUhqU1ow+hLXeDRQ
x1819NuUoxQSaqNq7BdgL11C/P7RixIjbhQzLD/ZrSJkmq3xbrZ9xMKGQR0gEbuQ
4BX9tVu0Wz99Rprs5lKRnH3F2aGpwYknl2NfLrT0Ffjg+OkvHv2ma8bvocT2jl0q
IWz7ZEUL3r3KYyFuzL/2pzl4kRL6K0qogLUBLZmziDjqjVz4TD7XfOKKz4dGtCKn
wwP/lJ0c5rqlxJwVoVJb8w5CNHwvwpfvFi4Bm53qa5TwL1iVlTEXLFIq9f/Ibrkw
Qrwbj1x3zrvU4q37sjuzfILCTjIbuPZNE4In7iWTlbBd/PkVhqxgz1hKqYG8NiIL
ZvCfM4BtIv+dMbJg8hb7Is40lms20Cj38n9TOPcWPP/vxFrtEX9xkW7b2O/WxtsV
qnkCKqUOuotgvufvNCsWUUAZgpjpWSlpdvxkVEqv2D6P14uoyEfOZpBBJ/YPfvzo
9SkrPCMdmD5irWI06fNfiyOboJivX2GFthguLH+r/N96tPpjz6bhVAATRH7PUwTs
w5VDbvQSj7boHDyQ0iVfto/9e5hub4fOV36/7D/BqvynAvLdrLsNE6cct5jT2uH+
+MhD6X4JZqfbyLcFgG9oj1bKgm0gEbSc8ipB8JrDg3q+8mONlsr9OEgr8ES+Ani9
g2N8DNgMoOJ5xsUzp+MBk1dMnZawjbXW+GjosPgmYswDquaRS6NHceYuU/dyuYv+
LGy3wmrlIGFemCf0PsfYCq8RgFtxz1ETH1X2UwOb0aobGTSPRruk4/KegbmV9kid
Hosi6npu/XBT2+yreYoki88LUhYniY9O5Q/oyHgowx3SdZs4naDiS8vz5P3h3Y4P
tc1Q3bIxCrBMCZ0/Cekfglbt5VWLkkTPBsoVrBdK/Dx5I1AcCaXClhWKxdwUzIk9
kBbWQ/sSbgg+vV71AmCcUMdVyWji6Cqrvlsl5EZWAhxOXEWaEGjXG5FnCzjhiepv
9wMJfZufOdVeR3d7BWa7icW7arbSZZQ8IZI0ggRFPCdpKp2jJNnfmwBNxftFyi2G
5FWdA7v9MFUWu9doixP/44HHtNo93tTknSpZn/MuB36dC7LhhqF1OdPvaMPCmbag
2TjpiiC7TiMOQyUOhrFKTd5xE9LzaCfOFxUE7F+SYVmTmtzwZALAyvM49u9T4Qvz
S1yvUZszRDPEbrpfVnhO4Oxm1m41NxPLaYq/aHuwAf1zodzxhCAMwyqWc3YAhGIa
USDF05jcJH5wlQRfdLvbYeyRytojvHHUcZEGWsfdZR7a9h7tF8ZBavwDFLmtkM5j
nuNrAwUUuOtyf6Y9MKOkgI5CFnTnTjw5KYkR+90ijodbiIn0ipWQFvQz/xpwRhZ+
3ugCsPcmjCSqERQ5gCY4RAMF4Suc3EYEYNG1fta7yuk61yeoCLY4vXIm6o8+6xia
`protect END_PROTECTED
