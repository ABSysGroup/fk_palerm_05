`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0rwV3nuMAuiqt51o6bT6wDai/q74yz68JJriuckwzIVAMB4m2FH2edKXO36Mo5U4
lpVA/pPTBXqtRcrhLouZ4YSDWZ89QjHbzwE0xzBT5DzqRI+L/p+iZC+GWo/9V3O9
vaj2lW5oNC2tef+oDEv1z+LMGnS1rdVa3o5LeYqjjB4RwL+UfXU8xdbgoHsJM04K
BNJBFbK6hW7r/7c8DsqDFNPo+rCeS/IZgmXibeikO8I/L7/3c0DeNRhTtNDIQ2wC
yfhkhvqRSveruKhrjVg82u9QKs4c1rg4NfE9ofxRYqxkSeWw12SNjJ1fSM49mn3w
Ul54KxZzNXag9tWZ50amHF9x4weBfKJFrrIJHMHguDJEb2PD5APMWaQuPRAk+yrC
xn+502Erkbwxuc6DYNkVX4p+59p4IWsoGRDAfSKPWwubBhvp/eFvU+Z/tK12aigo
XTfpg78ggbkINEworn0lDgWE5nNOPfxoSXIQU4hD2G2M4WO1wy+o39hQOyf6SgLn
`protect END_PROTECTED
