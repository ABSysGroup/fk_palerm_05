`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N6s99g3QZWcBNkgdhIpQm0MYzyNUHECmQ8qCxdPeGdaazV/w7i9HPRp00+1d6KJe
5j9IudXcxmtkIzZxDegoIHIZWlBIDxWBMLyTCpAZFCENxpoz0r45W3LkV4wHdQrR
2d3ADLNh2ufV8Tc5bBm5CCoCW6zo1E6jmMNLN2KPig53iC++/sMpnlXVQzVkRLep
flVavzFW7B41SVDoKdo7r0H7zDsNnRq4igXxwRMl3Pin432+anH68VNmd8Ma7VIP
l2yra8vXC3ktixtaMMS/vwYoZ720EzPJv5lUvAs1DSslij4K3Wu8WUFdEtlMv/Er
599ZYgUqBzRKmKP3W9NFbecm6CfQop+lLkOCEexZ0vgIv+ZmhgD4ASVnbo8MW8MH
e2h+w3VXaIH4m0V2HVKRmDHRz0yo4xIT++MdSfLH0rbcIzDohedmyN/sZmDLCQDV
UB65vfWfA7JxA6wLGs+sfo8NuPCvjgMEeMCiBhzBgzmtWy2c8QYIeSVJcKdhqEq9
YVBXclYYpQUiqLQTBwCrpBPsXrsLM1nfzW3Mh35qQL4UE1NVu2FBn8op2MeCr70a
TNunPvZr7bz3HOc/PBS/IwGkW1zsbzpZiGO7aiwL/Y0U/xx3ohVEaWcxL8DrIv9/
5Ti1prJKxB1tSpLKk9vpjjqR0KvrCRLkbNF/2Alp7kpj65LV/LAdOLUyZY7OypRc
U3fy70eJ3SirsXc9Fxnb35oT6BIpywj/M+rjg+M7todhi3EImNBRTPCMDoUvTva1
B2tXiBskcHqyTLzho/AImE4UzK+mqw6+720QgwCrxzQgF9HgfZaHA8YXwjTHSCCx
Q9NWq0EBY9J+jjNU/B8jIIHq0UpDEVIIgmxUojkUou6Qd0c14RLKuHKlMb3ONby6
1/t+llEFWcJhD+zHXdIFRVlzdSMb/eOnxZiuWXcEXwUJbIqus9z3XoMy/e7N0YkJ
tgu0L9LhQMnepHlKnt4B4+QtdTWZ/NhVmWEduXa9GiXyfCFvJ3jJ22/sOfRq4KIc
forcf+niOFq5fJCOEqqFCw9Cv8EQUfZd5mU13Lz3eX87WKdcnzSICImvdfWNhY33
45pwV4zqr/Ka297TcSL5os25wWZAu0WWX5ECkAwIuyNzPPs24l0TKIoEHlaFL2JP
tfW+7dbgeIhxT6y+oxESWc8wtk6IEkbyCjUW7aFdqaGDawPwqlGfQwmjrJQNg2Q6
Znkl/mFZL/mYMutA4nFobk5Ho6pc9Kfoo4Y4Ikwx58SgqPEwGe2imk9EyM3FlJyO
AsCVnze0q/Go6bQzAfWmcGXNGS3M10vykSN5zjXYaUciaDeRUns0MFWn7BxKKGiZ
p5j/NrWLZZyKhiAjoA7HNVwkPEQKirbaBHxUzo4FNngEfdTnAT/QCH8eRiv/SSev
0JVRXmiiDl0Dv3yXdVj64ppsBfyis0lQHJpvACAsFl8IwbBRwrFT90IlbzlrlziY
pxMQta/u/v1XZUdcEf1n/ViA5Vjnv3Xy+sKOh4VT/sBKNMWB/Bp5u5tWXHNnVgIP
OZFaxrhu5S2X8I8763oUohbylT9d10SMbwYffebOkbMAb1gBI+HLuMWbxtgUi4d+
VKzP4g0lfj6ffsg+GdjSwtjtr0OaiaF6fN4BxGgdnmblJFDSmnq/BJ1Q6tGOUnJI
+Im2bXNSYsI2wPAlac+6GOhTWA23E41E6/Ji8LOE+1Al2umItMFDf5g3Xd1eBpSu
+sFhDWAfWvPNhSrDnuLfc1xy5woyMNw2Eo8IVv7NczpQ93lfpv4uGF+T1whMMiE5
77P90rhaq0eJxSka3DzBjIJmOe4Q/jVmFYwtgkcK5hH4ODLzebpo3po59SHjkoaU
sNn4b+OSrDtcTKyE4Mvm0LDvq8FXuER2mLaI2WPopMDvYEgm1N5uHB4uld4beF7y
3UTiarm0BPQMrnF9JzdPa2OIE/w8j7yHvW5Kd8hY20UI4zLcKvJzvB6RqMgRO/4b
jc+heCYvvv4FzMXlBDukSX6VPsKvsWCBRw9xarHkkM5KOfJ0BRFmHDCJ70XyTczP
DPvL1zpUxxvGHmy+iEJsSoyupGK8yT5xlH34HWEEx2OFyOCE7gkAWwXykEddDXmQ
qTthoeLE0e7YzEsNiyzp3sby0zKDG3qZyyTlsvi+xszKbJH2c9VFzTf2GGLmVIw4
mygYVkoiGLDfarexVVVtGznslOm4zouMLXuGSbJJD+JpJxI9YDThKHG1qkK6pUEc
MJQLWrejoCyZpbuGzq4g+40+r2q5rmPRPRRYQ0SMR2TP80sUHny0xGZ9Ju1Wwwbp
yMT6QYYz5OMXf8jQBpze4Xr9JJ+H4NgluSzpS2jhmupIOxIq4gWfQXT3EmzsFKwy
YRK/+5uqoO6t4g34z1BeO6D9ZXE6cat6Tk23OUOSq8dBjGKG07ci36ttK7zgFCFQ
9sqPT9Bc3NeXv+tmY1kU95YNUp3oGdgZewzVkHYV5k/VVJtcKPvWUxnbEp6IPlez
J6NTkaF65wvwCmTLn3WvBxpXlaSgSoD8rvtKupmUsWksb0FAFxMyqYD/d6OKI1H+
u/6NIuI03UzriYWVJyzDC36MR5sYZqCggFjNMrKIN10i+e8ZmJ7uQp03rLOXlKOg
CaPIxIOFbFvJ8do/Sbb2lhV0StHhfKxcT0+xu5vdzZ0nY7Y8FeU3rX/lbQwQbfI8
x+dvvRZNudum+8cnWJ2hjs+ZN0zOWnjRitujAfnLGdWasRtt7hlv8O10zEziqSLj
cQdzMeeSQloVof/F4tNx3W0EyOP7Kwh3JQh7cFxjRVNQ4+qWgTqkRdhmuzxqQU+1
VTL2g5M1gJ7T+lgm2lwJJD/VXYH5Qvli6tuDXGDe46l3f948Fj//hmiZIfMzP7EY
+Jx+arNU9YiLDDHaHCJSEn5010mtr6EvdP0zL5Itpwexj4XFBjt77e4Wli3v8aIf
JnnMqPYx4mlGRKpAAHDpsP/SVH0KUN6U5mF4o+4Yw4MPFuhq68di5BCM3GCjbWeB
SGNZPeyC+P7kP7XSMYYm2+c1wci/UK22+A7Tb2K5p7nR8Fz5wRCoE7iLGMdHEW01
uaNHwrpHbsBlZf/6IYUsO2DxNDoJviunc5MUydJJUC6Kg5792LcsFv52LLrTtwzd
tdOvndGc1iF0E1jZW9BURonnvya0vDq6UX+0WeI54r8oUH9D6XU7FoBlfp6RLlIf
H2UOqMIWy3daZLB6YjD13OoRZlhcK1XdgeZH0kVszyKo+borUt0EBHF2UK8B3mts
xMPp7PAWKPDriDbSGKoxXEsgKpC/Lw931aAIwRbpBem20flQC/ZQYOQG8GxJIX0G
HmLxOajPOIwuConGukhsJHcS8YL5nh4ysbI/T75Ct90pVyOIz+2u7RL6tKOfAfX0
Wz4zI02kjls+bm24MMKLLksQnzLv70j/KlXPU36PoaIdf+hFJS8kc/i+UCSY4UW8
TPRIDBm69tsMHjmj80hUs6R1pegMOvqjBGovOPhPoNz2kDyemACvbPdFK+/fg4XJ
Zlv6IZ2/kNIPv71ASEhV4IntmfX/Ie8uUgGIclZqPHjPwrZcLROIxCmh49400/5Y
KzzkqBvTE7+MHjpVmfz7aqzgKkGfdPBndFZda21YlymgFeOf4VIbf8CGQyxYsEIr
6CTFUShlMWEv5NzQDS8RkdAMc1QDzy7UR7w6ykBrfRR9ZOaZOiDPTqNuKCM+TgVH
vvO3T7MjN9WMMzvvBi/bAI+se3MFSX6jFuy1bxujA5+oIz3250w88832Vyj3LHVH
ScbS+v2ZgCcfqLnJsHzafxJtwkqrIiLgL7zk31Zq+LyZTCf7p0o6h8w0X1VBDjbu
YvHZip7P/Ml0IphbVpVh77bfVP67kXd/BICmBOpfT3DMQRdunBCbZ8qk5XI9WyIK
e8XXQ2OjkDbF4y0wIRZz0iMxst1YXrtvqq7GOKiiDBfhqTlK7qKf9RW6Pp2IjlmP
O6qGm7jS1svtE1KD7dH9SPT0ilOVTNqRU9AU/+0oeIzicAoCbi1BL2VHHTtNzjTD
IQNiDSJ30GZshyg4oBu2xg/tsUsBYEzpXm8EvO7K1O/t0vdCI6S6Kb7lznmDktLL
R7FYu8MtxzL/JRrif0RME0548oDyp37k75Mxrxy5o3ZxGPbE3YCMfQ/718Y4nySX
jGW98r/LxkHlXCovQCiqdYrZmcynOzPvGMphazrsIXe5nVvT0cBLLQm8tuTL9tNd
mQiLTRl5UYV4MOWlpRWd7/Ai/Vs96jPvxlO/StTR6U+Fkp7ZcgIqzT1x/CcuPVls
4LtV+k34mVOSFsp8x1tfXMSZrloNPK8zkOyZDThcIm4M6orOQBnhR1TGwdp81Yoc
X8zf+g0rUFeuEsAyysUJ+OlZC7y9yUHK1stBeKpQqNiL1BAdR34rApwuEFX9XYRQ
b5sF03NUkBLJ8R1wwWPZ+TJzwkC4d1lHdqVp31CDMVvkzp8YYE64EFkVsonSvawS
Wa67W42LTkTVxltpaISIn/bj3xvKu3C9hbqIercmTYkJ9neStQWpksoppt1x6L0g
t7z7mHC7iWcFVF01xjPn06P+ovYasN44u2tZo3APJuvm7lK+OXyIukOB9czMm7J1
e38AmHzl+SKYPEXicqIn8c50rarwRz0xPqUM4YLnRkMnYpUpPN3TNAP+zrMxGRx3
DUAsgn5A5sXMXfexcHJXnzPjUZxEvr4zA2II/pJmq9FHbw1v255PDUzDv1ZUxyql
es9FsnvRCOIAmrjoPpDaqJ0Jdi7wvNhYt88o4fOjdVQtcmuoRKMnjA2+8ANTOy/u
yJXTTCMuF7V+SOk2rgXgZwsn1JmW4sW8ptwQJoRfIUwg5H6GCwqPixm8qUYiB5i2
6UeLSYMxIEWUUo+tzrIrFZwt2Y9TiGyWIUnkVB2L9hvpg9z6AOZCF/AaeYpbDJiU
JaSUN6yY0zBT+9awULpE3NpWEcyTdBfFVa3Juq+y+bMMDNKjRz9Yf+dVBFmyj41G
zGxCD26yEtOcwuY7gK8j4PjEK6/wVhALfLSOYbs1fuy6UXfVN0G7AfjSBY/H+pYx
40FkPhgP9UJEt5fFQopnH14A9JNknpXfWaD0bCZTqrSmVLSddVjCKgLm6xieuFm4
DqsRnsGVtiUKSJvBzsPdIetem0pKphi3T8X4T0xxfZduAgxt1KU71UxuSTdwX05R
AGSUfg6ZVcHQvc2Vyq6THM/Fp4EAXy14aOJXJ4fkc/nw9ZxET9c9itgY41jRpoJD
GR2KYS4EYLJJ0PNmAtD9o39b+Iadc+2oC7tQYmPAsppPsSJWKvKgkC4lcjqFqDNG
3Djb6PT/ciajR6yUTxP7WBVe192lxjkW0IuUH6OdPw+I+FqgkdZ1dw322EwY2Fi4
sjY0uINK9TBC+JZ8y1wymPuzTYSTv7f5ImpKXin41fUmlL50ndXtNNA0UNTMilHx
zGYF0wJKIWKl+yB5Gvsk6V6Zven56Krsj8Y6EgXhTX70O0KWYxY0hhw7xFVhTyC2
x7C0IOXzsFAGVLUxeAfMf3WHd3jNyyj793M1Cwi4a+8Pjv705i9pkmb1fF4YYpfQ
b7iN17d290MqJUhzcqSN09Re4cP8hhEtIG/2fHlqrP6ipoIuSZrzwlZUud5uibUc
NUkMQSwSTALVeAlRGtAykDf1kXpG77cCKj3bPwk1DqkIL9vThEs2/B4jpysD1GpW
PGXgGTuNOpX7wKVusNiAfiC3ilk13etMNfK/ajqzf3zI6+NR1ONqejO/6VuC4j29
cMv1zx2M97r7/TXykZkywB0qrx+PuQBUv3+j9KvssPjEfMZrEVVcgZu+tKgTZ9k8
FWezTrCNTywaeQDsQkCryblvERE9JH7n0jUhKovEAbfMHeK9o5JPzzZYS2nryr+g
Zw16zcNNeIcr6tZcfss7sUPvU6C/W2A+ikpG0cEjmclAwGN2W5L4ikZqitIYGkWJ
ejxbSp+WqIuA+4Lkc3ezmLZHCO66rDPGgqbd3Dqxi0a6Q8WSCkWxkI8KBREcMpeS
VO0DkxlgZ024ZL33GuRb4cFPkC1ddinT41wClDRH8ZnCdOjlw7H7lwbb93YXE0GM
S62fGVji3bDQo0tcqevDupR/fiYaEN6y+Z1fA2wL3LRBVc4iaaY4rIEfJFF6LRWT
nHXy+i4S9JeUgIDPRT6lpwLTW/yKonO8VdLt1WC54bGiBuv2jDaL5s5YnA3kNrU3
wqCn1124oddigj7f4mNfu9fF1TLEObxPeXNQUNLAzYW7EJU9OQ8wJYF5OIG8tKa8
z1dMHyfbatdZcbDZIQXTD2YzLld+Vql2YZbKfujza3ytOvQXZ2hmjDzFBm3gDfig
k4/ectIVT7Tm2aSiM8VorOcjnqLdW7P/8YjhDBYyxABt+G7530LM7e0c2oO75Afu
fN/angPZqg53svj7rPxh/JKt1HJEWwxDeYwXS1VyrzmOdI9jhKxJfVJvmYBP92u/
nWPBXmQHKh6LUFtZAz0aEmpfUu30gHBbie/Z1OnPSGKZU+h8KpA48q88OX5pJMHu
L4oO0lSDnvBlautk/xRFe7+3bbkwpQ2tkSyhhhKtUBJiuVKgJbO8jrBR7hhbMHXr
RPb7MRXODQttgV/NliR28iWXUmmS4V1NaVwuGpOz17dXuhIirRDm4+caEpcbki4w
qXfzJr+Ud93qSeltxOJG+04lYV6ufO/xYoux29KHJc2th/b52JQCSzeHDYgvokSf
hCpNDe8rZwSC0RaqY/OKk2SPt6+0Q27QhZbRm2IVkja1BY28uSTAa3Xpqkc3DYoF
PPtM+lTHuwnNhQ4vshjruMy6JU5p4bPHKYaMurk+9FTcZJCrjV+4dHG1EDOiNxM+
2QQxIP8Gk5wYNZadcmoaqYfcvFAn7DWSDMIrSS2dX7QHaIe9im+ooIhB19TB7jja
ve1EGXPrIi8gi7MOzCKMNAnXmrHEGJ3xkqoN/mShJH1u5sZtmbBNweHFq4huEWqp
PXSBAkthxoGoaNKXTKBXl8Mse36MyUDww6tYdk6tXPPgLhxnFI5Ajeg66oxikMTl
yjKApYOdoG1lYs8y/YSjWJBGRIiG0oMaCBrfUXCCxXJ7dsplB7N37drJ+Irk+244
MLJxFMY2Ja646KqKchlWivwCxvvRRzbKj8lcTvp7h8lJOBXdZX1EREwckoA0rsuU
WnN9udH1wt/sypzDNkEPZS98TEx09JODDax6i6i2hU9b1fXfgUDj98WTc57VV3Tl
85pMaJ1rei8K9gspbY1j1hJkTLjAPBQLI60tQGenA9SLK0e4YZL8xZMI0bIaa11Q
rO0a/csWH3Xzq/3Bwq3myQG/z4Pk5IoZFMPJQFJE+xdgBLQ3aSQH+oMKUJXJ6pdi
R3DAGPH7D7rHXNglpyWyoEVISdypksaJMP1iz5oHs2Q6UsZvtExpXaXDFxbWExTw
0ZbpDoaCZhSSLjNh9qkP4RKuIzkLZAz8OVBm6JKDx+sGxQcAZwU2Zp3s/Ig0qQxy
PdxndcOOuFeIXssq/boX0KvgG1CHJsJbywPeviRjDlxTNYJ1Lm6ctwTHQHrZ7xon
9E1NMO37NJZur7FISP17QD9R/ub8IPOyTfXyhme4ImMlb3yk9F1ue/8zZ+XIswLc
JH1vBY94CnHvth6mMIrvw5xW2LHCKki06iqzNk6Yg9VYv1+/iqxvd3SWWc1Wh1Mc
2YXUod61l2lRsav2NAa9QMk5lnwoEPzoyGKSqcScCbi85bkCXujFUuipWTGE6ZzE
0OZH6OlDWz+w0/zBsGPso/4zOH4CKJ15nJKhn9SgcHCTxb2JU2J+o5KbNwi/AgJZ
4kLYRA1+h/6zag+9dxBTjtIcakjiCogElUGQw5niNP57Z2507KQkWKzieLnur24y
jptU+goq3CxBoPQdT45sslKQV3kdsRrroHKpkgL3GwZR2i9mmhkYhMcbII5XC1Zq
PUHIjNoHgPh708hKUJyhouffxZGrN9Qr2T6hBxPJzHOp5K2IE83E9jsXCevidsAv
9kfcAPpOFHkAoTztLOt6j9TAk4ucRIRBO0jwo9CCBn4yK1J+P/Q/YD1kVXSOwam5
IqJzhhpEm9DMhnA4aJoCABwTHcRiFyw4JsnrgJ+q45fNy4mHUzrD6+HTiIZTalU/
fewwAYdWidThb/UX0ond9JoUPD06N/FvXuCpWMl9l8AMF+vwIXFG8QcPz1MdPRhO
D5rtgKKlofxiVXWMxW+ReczWkIRylTISYx4qaThTNEdEZ3XCALZGOJx+6IF0mSoJ
/uULsMVzncKsxFUM6RMyMbCIoovnOZqyJ0IASEI8UxrsQCboiXt8KA47Mgm4T/3c
Q9nOsCySqWFl2+BsbLOM0UdrN5uWWL3tLXwcsjYRiRGQv1qAhDX1hkfQ96u9nWYI
8V5uddenrf5YqLpR4E9qiHnzG4z21LlrQK0OSpl35Qap7KZfqMavGzEdA296hHzs
zZHrp3aqumQUdBdXjMUcj9S8smSsKhaErgKJFotdtIZRJjg44dFFv+w/OYwYkJ7J
4H8IxdP28FRTkEVDFQy7QMutlwzjD8wJ4FRJ4WPcLAbknODWksjq4n66cGgwE7qO
4c75hv4t7hJqS03rY/imsYZxxIFcRT3eju8wUnJhvHn9b/mJ3FcXY+S1ryY2AK07
hkNNp+JYmEzY1wTdHTrDieoszWxyG49aSIs+G2MKGKFsBCvDZdWjmym7j0xuNLfF
AwEh3WrVSFaXhgCUhiaKZ85IDSMtFVn/TpnQGFhSdBZdmIL4qeMX5TOpmQbTvUHS
gRkfjc9aU5UN85pL71WaynpCfN5jyVWwU4ItupAkR5VCXSGrh29PTrQ7DCo7CjmG
0qv5ESmgbxxxfm6x0MIafy38+vEYD5zwTaWy4JqlMlQMgUZSUJeCPuvjq67ik4sn
FaRctHiSxj0gXbTVtX2jRvzRKXICXSXMOTY49/wQjqGxVMWMwwDjEUAPNcTCwj/V
IaK0/ioWzGPjxDcL7O68vp7Cmqhl1pxyU1H1BpAwekcnwGCGWq2B3vtNT3Iv16uG
Py0+l6GBb9sWKmhcL4Sjj8JmxEstEWU2e+0vI8EVo6paMUeLdikmK+rdnO8dvZog
C7nUJ6HeDTM6nt8lNhotswkKMHC+6rm5NgZ7hcYzSKLb21+2hT44CwAFO/EHVjZI
5IO4fOxWY77RHbQ9KjJPZ35hpJ4sdty2nsGJyW+6hBbABQz5E08KettHmv3Xx/oD
1Ki02EHRXoTlQeew+UvW1ul7dmZm+guwAGQWI6BmlzKZ1LFaxlj0zlQVc5F3NZwc
amy0U30JLd/dMud890/hu0xNkDesDcst45PRu+RiRk9FCOGlXDwOngwfO/k1IM08
ae3xNF35HjcrMMo6DwM8ZrXwmnO3TZw/ncPDctTwJtCwhrkKeFkzsiMJyAdyJGOU
+CDRTRDh5f1LvIV1Tm8kwrMhcG3uwmZHWZoWhTUhT2mcc0SmNQEtHC/8+xsti4Oy
QzyKynrMs7XntI3ZMykvt84q4xcRLPyTcvnrKFXKv8G5lmcHPPV9VVCp79b9b9z6
njPQOuav45w9aHk5gpXaxw0eIzd2/d0Tfn9rGaeYPJymUXHGatmLTD8NwgUy3Wlo
iiXzLKd69dJjUL2ApR9usBGPoEupNDvAFkjBt6FnlVbHIHGZoMvGOVJTIHH4AXQB
wogRBH4esGZTu7YxQxLOij6APaGzz1leZcgnaXKO7K5okdjkWzpr96ND6HcQvAqn
KBPed6U2NCHFZjcXiaSXJ5WE6u1yOgezXnxqA8HKre3Xpq/g4km9g38ph0pRbCWh
9vjSaN6ejIbLlMLM6KCZsWGhk+f+K9E1I6PWmcPPjhUb3q4RMs28LenvxJ56NRsm
UxA2AVwQ4GMJQnMbZtpl8dwLiEd0vM6bWt+xeiC1qJ9x0aYeI/PqaYK+K+EQTPpA
nXM0eLZFbO8uPUkzfmnGfjw9NE2f2uNhaWTSgLzKY+DJUwZ0i2Y8ZvYjr3bBFncP
mUMgUPahL5FOW6qL9chNU+q8lZtnkjkD2TCvDWPZhEQzGSbhiym+7vZJR9RIsiTv
c2LeWyYmADlgVfC+TzYP40sNocURB4q8Dwn9hNUkAkAkBkj0LsRutaJoYR7rX0ve
sXc1QYth0j8VIcY+DXwmKuKIPxS6FVIsDnnTBShUDzKAiz5tjGyDu2lm0Qa5ZNap
6hnEfJNDknwWiC1RI1Lvs/sJuiCDz+kVMGqlsJOLhspdr0Df9oorbb1tR6u8g5vy
rJAQZVOmggS11crhvVD6h1j1iL9oDC8hRzoMmRIsYQBq8Vw1/0vB03WqkiR87llA
Ltzk8L5fNP/dZ/vqtYL3srtBM+EaqkIZ02nf8KapNCXQLIz0UbKoPPqiB5doKmyO
wwafOd1aKMie5gXWJu+oqF3GmCwzQgre/A5FBXsdvw8b9Xfsf3mK4cbxwHr5hfEG
dD4kw1CKdUEKgVRro6E7nj3W0qrwPKANDhXvZLpum7SLQtuNCJ0yFskfCV5BJCvh
aJNKTI6HXW7IAXckPKxRawhq8fGb4fviL/TnFGOOLkjzEGxNmDEqy50oG4SQZBBM
LSJsnvU+OBYadZKfT+3lVIXZOz4bsYQgsRPAjmridQmMvmC6+GM478UzUcbW+QqC
SGIaszMSGzBU14Rzwb2Ml0v04PymvO4VCFDNVVeJDsQoaU1E/3VJjlCAeG4a3yCN
XjVMRdOb0HKSUZ0fMxmMhyIggzH1y3BsYsQrLGhIvzVI5E91SPNBm5qkOmk57biN
v2rClNTajG9MBitNHprWYD0aP4gvQ7zTXK25RG2j0OWZ3gF1ZN8YPab5lK8CY03d
sg5YaBXl3E580VuZYq0jLk7rhu7Eixpf3aNoDWoiZxde3bBzhxsvAzCG2W+tWh0r
jfPmq/OsKWRiTKxyGAdrtSnt7FxqfZ9EOnL+WsZZ10A3oZ9XnfnS7n/rAWwmDXls
Ys3/vyZVZ6CYGcSo1RaIPopry9HKPMW+LU5aMEstdoAjomrS5PFx9yjipQSvws3P
rohTZZFYfTRL8y9P9EzmKjmHoZt1209bGG+960BTHqQ=
`protect END_PROTECTED
