`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ynxp1IYOSwd579ZFlm2MZGjxt/rfhGu+7n97KTAV2i15Zc+kHeBNi0Hy2mJKraL
nUrqysglsoUzB/tIrDsXJTlKHnoED60X4jS69XF4lhH8h6plqhxOYKioYEC+f0/e
SNFzsHQchuq2IxAMGTAo2j+2nQtcaMynO7C/82FX6LszPQmSEyQq6iyn/S4pWzoL
bg5Q41knS7JeLAT7yQz8QxQGjr1zTTY3e6DfTaHy1Te/mbfmqdx9A89U9uJCP4A2
eGjjb4bebbUWpvRoyR52cHxXUVLznjShMibHiT7tajyZ6c7CSlZGm56bj0mEM5el
RGWUVH7ITiSqtlOCSf/vGy5qj+J+vIC6hDAaRpAzudhgR8xiieigIjeWS/UvmUxY
Br9te0WD8F6nVh1doNfV7o40Er4GhY8A4PwJGbUfqcbmcIJOzpsQXfaJUF1F21Uo
d+uktEUXOE6iOCZx8rRuo/x3uuKXU6PUTy2PhJ/ri5w=
`protect END_PROTECTED
