`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SMV9urOA4hM35DkVkEG/+9mn51yF8VBxq3/ALykrllmO3mgNa8D0uwSXn004caJG
z2UY0gaUJfP84PzRYnWQhrvXnx+P4puCQ+nkjjmpDKobdcWDKYmf2E2xOMMch8Xb
w/vfCxPKoDYTh1J49QYm2+XJy6DDxk9OKVzlDpfo7jxaj+4Bjal86hXPK87x2Z/h
cGVygStZvktD3C1rEnzWj+SAcMtAANyWO+E44kcsVDbT/3vtgLmdEJfVbLV9pqjS
Dbe6LKHi8TEQ+ORJwOKPsStryKdEQqJdxP7yHQEjHIxzWMKGy7eP/cdt/Jj13iJV
Hxx2gzVpcRd4GbRPSQXY4k0N3tSy5DdavTQUluYYfKMQMaO+Tx5WrgHdjHEpl80V
CUCG2YUFzq19XJiqxa4lQXhsb/zjFDeSma9chYDntyOlH44uukFbfs2Ut2CByTWS
8OYdQxqIsT7gnGFw66KcajPKpBQkHpZn/n/u6w3/ww0Ns/PstdWamcElXoCiXmMC
1FpcgDeb9Z1FtSz+sttP+Cj0TzEi8TMS73YamvHIMTzP7CaboYeVwvzykNpLrdON
QmCjYzR1LlvR1OXDLRr/5xJWtKJyf6m4sxwPhupfOePhu9tF1avfOFfhNN76stgF
Z26WU6qT6am19DBByXL4U6mDzrS66Q5s83IRwmTWs71ZwxBN5C0QWZd+AZXWm/vG
JXT7ZQymaaAtmGR+2fIi1QXgQrrRYnzGtC3HShuaJUTepiBYLmkBtFo5dWiZm5js
g0cyAuWYdxWt2EOBeCHonnVzIqY0xevQYkYo2ToJeKHL4cmUe7Oi3AUF48T0X5zF
fRUIYX7iFckzAlwghn2L51+Z0zrlQY87f6/qRdekTiNomY3WxAeB2xuURp/YW53h
Y4qeWcFxJfuSPo0E8ZAyWOH0x0I/SX5rQAao0L6l89icIN/Jg+RJZ29JamdZItFz
UDmCTQrabDOezyTPY8fCXUR7iFtVOHEogqkcxGx/BdZ3QwvnBHca5pWutPPJ0sK1
MIj4dqzU/5BFmY+gGg+RSclT2DrEZ05WTjtM7MkvFYnKwkCGseVf5B2s/itCe5/X
o+1a/ltlXZCYRBijCRU4eON5h6G9kSzvwN78JGVwmizATroFNGpM8P0hiRjXgR+o
Fo04BwfMWR6idLCkIHijUrWxwcFg+wqayf4nJnrrLbXKqr+niCWgAaAfwfdrcdnJ
kVKxlT7J4vCWGkAXiaUasMfHi4cAkx8IUxJfYfVquzYjQrlKyIDAV7jD/5WYUBJw
YbhiPS/D4qy7Jcq5iUARqikztLekYKgs/v2vUC5oVh2kG3E/m2bw2YFWCGoLPW22
zcTUx/OJhEfeXFQk/uhdruFy8zt0C3y5cel5yVG0qY6lf3Gb6PaMOzjd7yTGcLrP
es/x8hQaqcCFt+119VpUjrNhmZJTt/eerrq1j6bNEE18Ux2DwEMXqy4ms/5+v2pu
WBx7ba5i1AaTC3REYhTvzPqrMOvwo/9KF+GVcgI+gQ8ojZLddqpvoMSi5/3bbPkD
wPaNLki9urNfONqwS1UWy4IvpwvbddqINw7qq60dSGEzYk/abYzPE0uNMWv94oA9
2z1ZQ+KLUl38wiTxYbajJcpW2QIVgGWvrmA1cZgT4o+VW2L1sHXmCqv0r5tNF643
oNN6wUUklK+a2cKKP9RaBZeQMJwkOE1QsTgtFcCM7UoCTWGDDMB7aaZ/98b++BrU
V5Bg4xYYFS2ZXL/M2FWYMM9HScBrMYIqdDb2fBhfY6SM3F6FGdsemBpMMOlCP4Jz
IjTaytE6BbtnVy03SWNtJmoCRSfXRrrnziAMMlvi1/OY+PrSHAiD3T5rWudPCh8i
gkcE3Pm0sfcqLD8nte5Ojuezziy/yRoWFchjF5P+g3amqafXJWw3oBOUTbRPDi0z
EYWJSLGNCvLwtmLq/u2ODBGSTnQ849peOYa0bSIR5WPFoDAB23UvlqIKznDzKuM+
wUC1pwJMLRilGSAvfqE6RBfZ0/BC9aKI+VgohE8cpcVu+4Jyx0byzk0HDPP+q0GJ
6Au1oPfIC9IP0ut1emR2yi5nvhwqk9v1xrvjAVH7YlcHOifPL/a79jhUkNo+iTpu
emovQxhAr9T7zDg3qFnMVuBd7G7geWLHPut6GDGiTvwi6K5khzu2F/4uULbvV1mO
TwHBLavSNTSdDzd4PaBKfy3bGyZP4cfdq4t0XJTeAO5b1L1ciTTYuHS99V4tISDP
bbREvfL6FLppkPElW07qbp5HmXsHsE2TnzDpnZOJaPfWHpXSksmv733F1iNehdhw
YcUfyjirnTN1HSaJGBwmBg7zrtSquw4vHbjXD1T3XGXu8YtlYpk45C/A0XR10mdK
VZbRW9BcvaCFcan8YYK7+aH+EMqFDsEXL5fpXPmPW8YkFeD5YY7HXyqLHmU7Gf0H
bRIpkes8PAqvU92383tpXzt6XFVvzsQbE704jJVFN/iFeuQclCekS07HAiO66FKk
HUCzTa6P76jERwlaAOWLI38XzX29kgzwuPAyMzke64sxEVOSMTwd/hwZ2xUZukRk
4GydgfiNOXk3j1Vt69IFzHir5wKq3jiP5Aeo91NMPWEb3a/YIg6BbHb4lm7OUdIy
vgEQ3eD6FnZNsvh3Tv7hP7lVAjKfJ4xXtdkeH7MMxnnC3NOjBo2kue00Vki5S1DX
bICgLEL2B/0TU8ZwrYwZ0xcpEtWXvh+V4hYLkWaNe2DrJY6vGyFGlWMOtaFX+oS9
MhiUMEamh4JVYutbmAvc+hQ0sxmQPMuh6faZFrEu8Fl8qLkSBpS0E5UwiqKF6YLE
1PXBped7VzDpsKlKo3UQn86tkc7g9L5K1hx0utzz9Vd9K+I/tLZEFD0tHyXyFQyK
Z58JI81iYq36l7pmiEt4WtvMTqH1ShZfjGfLHyg6raTRU1BfCzvrGq3OFzXNSbq6
mrvjLV56mgRLjBPMG8+i/8q2dy7kt4Y6QHCzuVjYWKe7OyuIMJdsTiTgZglxffyc
YPu37LffgJISb4lCCmEToJ4wezPNF1/1PMBUCxfmlD1S8QTZ8vXWcQutAOwJy4su
u6ZuPbz5L0be9s6w7UJ8qhAlFTOoc8RDtHOYGcEblq0+3bL9YS4bGrhrppapDPzr
le4rKFtkOkEyN53M2mzkGzSRS9oeUoc2iYx1oyLaWFysgiHKMI3LwaTr3O6jXdU5
hq3/7bF2qwPyoJSB4ejAn52FzrYHTsTGQd0MFi3saQJ2djPIkbw5rNvjHo3SRhiF
DFULZKZTgMG4yqcJ+bbSOlpVxsqGvoFCoGcu2dHaR7Im4UUi/uQz4/e+clKGjacl
qeFlHwBaIKVZYBb9Fd4Yx5Sl0qjURauAT43gllYowecmV4Iw2/knHoyHrqZzDBC6
+wYy2Iq8iwiEzbhnnsHws8WFuggjs3UsTOrrOnH4NajR89Kh9ks0tLakpI/DoQNU
lp6JgNyiNz6RDixY98R2gHiv7YvfanuYPdJ1Kb6HqdSUURFfFsY20t9oIawd2cIK
biSaFrbTA43ODKDmZAEFnluUO1/wUFd8QEFIS8B2d2FRSYXLHcH1OLlZMs7nyidy
Hnc6kVwx2ic1+OnJdSr0ht0P/Qn/bLvX9y+WcPmvzK5j3cmX9hNUYZqNU1v+mo/3
CWStoHCo39JSPOWAVgU7QZ92CXR6UAbLyldGiTYVVzW+4c16tpuVBVJ9h66dvPe7
8Jj+1IGWzs9Jx120l/pEy+8aeIIfFtkJxG3RDRAKYrCIjS6oMonSXpvgPTIxVq3h
9Uwm7zJwdaZo8DcTLvIM6bRhAvfgbU4O7yiHC6rEHUjO5O+wOZhQxSgG9OhuQOyL
li+AenxA5huUYi7gqRLimItVPoWMmscShE3EMikKFkLyJdEzvGsMtBxh4vFSHT0g
/1Ohj+3szFROZnteF0XFQwL2tQsnC8TrOnDhbsHmC5IORxtOzwkRIUrVZnEfB6sT
yhZz3y/KvzIdqyKjg7ujUtmuBXP+1yBWSIZH/39BCYMQ9IF6Iohg9NY1C7nq/n+a
D1HnZn7vIeO0vnZIVH1yysXV7RDC6bFplX+ycmepYmwrowVZiPZCkYXZbJt0jY+N
FNEnO9iAjZ9euZ0gb+BNM7F+uJE/30iCjw+W1IWgkD9uYNm+xSrjMczQBL/Axxm2
rrgcIcR8XNuiEGTdTdvfgRWlxTNgJxHT6UoVT29DARgJ/5s9BMmCnvpMxudqOTY1
Y0vWhkaUXu+kQUSHxDHYvbdJuB/NqGYaFPCrUVZd8jhTwK/U+ueCy4Yd7SmCWEoh
OYYOvkins5yqIAKmX3MbhQhuBEFO3bvbJk3Mw2lXnowWpMi15qU0VGBibvdJXnxb
d6QASm7e2zhShVynIsbgitoacxrWL0H+lGYu/y8IhPcigEnIFxBzUZqlgbiIPTcD
66fUmxF/MKl1Ig7bv2Gj9IVX9pwXg6/ZTo+8tdT7r8s2mC1iRlYUSbgyGxVEGOc/
nD6gCGgWIEPGdn1UZ/gaXuDX0haTwlfNGsiYa1dZM0QHmjjVZen2CkwCKhmziIEi
RUifztgUBMZLwjLp2DrmAZquKD1UE51WDhEZCJYoXir/OKmXazap07adsyqb9ncD
a7nCfm9QrQRrtflC+OWjapJX7j1F/jRaXPL7khg8FyDLiYo4WDUV0PQeLh6SOX0g
2dYw34LRRO1oO57Et5fguGQWW7ZRvpiD6PYzvoMcFlxeNA6s2rRJLZm2V8lYGDAp
CGXlTsalkF/3xrsw2m6yz6+aR+biayQ7s8e0s4ouaJ9SYLb4tppAE+bIsBerXlxW
sKJvXqF5NYzi3j+fkCG0FvJcvm+a950RA87IZMl7MHgd5b1y3SDuxPfzLA4oYia1
h+1v3EbKkbvX4lfsUhjXA0xUByOCVOxmE4G0cSKnGXSDryWZl49lM9LROswdvcOD
/i9vRI2331tmKN9hWjvpZTtlit1P/mh1cTZMM5HjhTTgGaPxnk088XdOems6Is/C
SSDkcR54Tmgjo/waGYd8ZvcI+dq/KcMW4gXti5mQqik3xgKzlttIZ2A9x/5OgC7u
AaDZAlhmKGhaHTrdinEhsx6IsiEadV2+Owq+oNa2jO0avp9SMES0XvrB4Umg5BfR
vi4h2BRSMGcsNvD/euaxjj1m+QWsS6fMzT4Zl3tMAOZhFBfui59idGDA6wrQXYgn
i6RSzAJf6Wkl2xM3dd66mtcOt6rLCDub1S3SjqFsJw3P574IzTBIWyhqsxKqU0s2
PTI2qEcg1W3fjNSSP5b/5N7RTapDzJnbVL1VpyuC+4y9Epj7Urtikj8K09KJHiXt
OHyJe/+TMveJTrtaYpNqa0RpD4YFbLP6oVuqWQeEgB8QvwnhEzHTNMva7bLMlVq8
oUoPH+WUKjRqJJf4CqQgfeefcRc2A7Fymro1rs+ZZFNixJXnwjrnLpdrOCS0p3yf
JlkfonrpAxqCcvCYtNLVldBGP9RppCCmG1sdPwJu2O81ahe5GPYK5jpgp5xsBgxm
1H5qRx0cXsK10Mh7Cx67LCvfCt8NmDBZc/q4uRZLiodUZyGWgYMAQRHadJYRZugS
jFV9+yxOUBRlBjW2nw7r34racaLbbmsB1+3LPPNkXrkwnTQ6pqcgyTdnU7w4XSlo
zNY9FipyaFcyvozWUJpUDzaRSANdjTyhOmqCQrj00tNrireAKKYUVZgnKQH57hDA
tLOJAc4TUV0aVERbQu7ZjdaNK/tmLIQyzWesSU7qBIdXiEJIjUe4k3YywPV3cQdb
0aKuk02Zj+cJ45Ukp5Ogdrtsp/HDD/Ekgf3oIJZygr1c7YtGqR+FYuecEILnwlnR
iE859IjbRE34xzM6CfN9r3YJqKwvD5M/EkCFmMDjPT5maDHiyhL/ZyRk8/2byJXi
jRwCiyn7gSWvb/XLGYi/Qsv9IzSX1scASaEiFhYzTUZlMsPKseis2sGCkw1bLk3m
XMAHen0N+FloRSplrln8qL/uR8wauzg7e3d0EOzacBq20PAT5xgWwxHxExxMb8+3
OKS/gOMfoNRnCXm4k6jNb/u1+UxB8JfU50Ie4EKlQCaGgZH2QNuKJPREE/FRlgKX
rt3xRnt5zUO9jH4iQZkkjKtxzEA6VQWUb29XiqiucNMcCyuoyJLGd5qBhPsMpTsc
e/5oRHPXkZsJgipgTIN5ooucP83ijhlYu8JebW1O6ceNcH6keLPFdO+szxaPLiG3
guezsP/NZwUzzpmsjmBXykpJeVyUHJs3h+faiEdX6nuujQgfyqiyrjIUK8HNeNKk
HmNmzieV82mtjG0pmCMeSd8Ste72FdotCks8mdbQq6SG+4iQxlqK7I5qRE3OqL8o
3yQmY2Cgn+353+J5cLqqsEfJ0/NZxLQe+GLY2Twv+nytcIrbm2526ljEF7Pk7PLG
YN64UulO6rQ59qyAJ6vVNAACtpDo7TT9rhdLRXWwaJ2wCNvq+OZvOzLs7r3txF+3
E8Slz4s6zuRl29moyNbcO5d6kgbd230xcqVNE/KignhfRZgdGwEIFbsA5xqAY0pm
jqyrUvPTqGDz1AzkWXJUPMp5WYU4abwJOEdUd+uTb632v5AKHsvpJtQCixOqXFhP
grjIfI5P8rT5GM6XcQtitzH8NbXWdljPPYSP/FUWLJ+OgAkSG2AoJosE2zFUWZEb
cWxrqpXi5kq3804RwRNxrl6UYrq32lB7mmI176YD9D0hyC31FHtldCeFKCDqhsUI
JuCSCKG0AhjE+KVncKT8EIjM7/uxBpsSNSDWaJXiJtLGWIld/Vf9DHSLNUGhurmh
PjUoU7sXMzkx8saqiMOwQLykjjk88anS+PVhvf6119wlZkmerSL1xY5ibj/BaRnP
OHmO6H9/HB8SGoUz8BvJCbBk2S5Y0Y2a0sGkmJ8Ghpw+qpGr/Mc9LHfHGqikbGYm
qoN5J6mz1l1RH7IEyUqqPcdgQ3z7cdfEAPu1vh9QJ4UASfaVX3lt17+NdqCIKONZ
vPqRnKvM2EGssWz8rGWqXY9NFaeTXB6PpC0k8h+wvu++vgVszfo8pB7B8m+6hMJo
s2Drnxw36vVFF1X2bf4rGCTdy7jpz5lqPNnEpUlHrIfekW9lhDxTmzyCUgfh0/G6
CcOol+1cL7d8+p648ieqPbnfZc5Fm0l1JLIZl+FYuxTDJ3U4PwVsr/z4vLwV88J5
UbBdk8N0Wf4Z+NqRhl/UcTgaXgH6zIfJMUPJIfJmC+hq0yGbvpexgBSWuC3uSt0f
34r5BQM6JSBqQ5B8HEItv53h67/eE2gLdlr7rFaYoBRWX0YJcSFoQ7t31d0DXIGP
eqcBehEAUmUvV+Jj4TJh9W0lAyTb4BRX/R98/IAc2xTbxAdkzdxWsGUkmFseF7IV
6APfWuGUGhD45QDpNIHYdWTkPh8ETkdHa4H24nbWyhes6pD/gYHW/S/RULZ7bHmy
lDEbSbJhPoJblLHQTqqlr75Kflg7K+niy2166WMGTBqTj5WW/p+CpnZi1aT2IiVt
s1F6HvEP4E5J4kvuB2nPVI5h65rS3LHytsCZfyRsj/0kKI2E/HSFbNitHWHLZqDR
MKUKyakFBuT36VvumyzcbJqs35kl5IeIjdSz4EiTtCOhMIeA9o/ekql3WBrRKp2j
1VSWPoUbEjA23nnlqSsDZ02GVDZVe2UX+qdy7vMYowKNDAhWbbO8PT56UL5uMRjT
X5Pli5rg45n13sNX4KL0N0TtggzNPR9F3n4duN9fQMzyLnueALrgWJCar//+iVh4
6J5MsHoRIFTrrfD8rOwD5cH09n+U4yJAxkwkQ84vJ8thb81Oq+0pMP0NK32wPKrn
Qna8IxCSb9SeBV7/K+nZ6Ca6Cu63ev1t82mAmSN6L15ur67IQrOZY0fsWHLiwf7C
yKoD7rkqlQGQHVMBbi1bgXtGL2WlS1b+Z38Xh3zVGAg2urzGqkLFhStyntv++OmB
r9ObgC+CIFw2fjFEqZDX7JyQW9tOxJh7MAqhSrShrRWY5FtBMrgakHbD4JhWVVhg
CvjeJqAIU7D9iiE4QkoYK1HdmXUxStEK1zMckUfdyMSmOqynDiNBrI7HMXd50f7L
qnTmhriWeWaO68vUJa+EUsgpp4N9AWXhB8nkOVy4RdDtkmqD6wSay0Y+Zr9IfALd
W1UXDUjkRa0mNh7r64R4bRwym2aoK3UWc1GSSgztsE2iXJROY/zyWW+3bQ5ah+6G
8eafcqXGjyjP/ctZLwkpbX52wRdsjo03Q0fwUvhjXajtli2hVG6glH1qQgCrcZBa
jyJTn7Z46hgt5nsbTnPHAHXQFadU1NSOTJRdcSvIKjW2lJ6G5lc0M5cp8Gudef/T
Y8iJ7876p7lNCk/TkgMGQXoh20vej5bYKhDVBSK1BzR8r4Ht9jStmsMLZ4q15yyq
DxmLXENO5hHruUdxu0xCn5AGKvqwPP8aagO3EPav2f2sm/g75KG+thEtIXnTnFWp
37q+Ed15AcZ6Pp0OrmaMCLDNiQUjypEh7hLfPq0DzgmATSES1lZ3E8QkuuB62DVA
jmbkDPmUz2KrCLM/WECTX1hzFrwBpglgEHOiRORzsegdmxxObjOrwEslCwmIrOn7
IRmQ2hiuAWwZpHQX7RsdYgsh6g+qMgozh4L7CV1MD5yW7OhM+uyMXismfKFqrwVZ
Z9mGH2EhCSz7EO7A9TU35YzDLGA9/L1gw+sXWOdaCKob1CxzClTxxkxf/C8T3+uB
lULEwqyVL609BK+LZXiIKO5TCrTD84E1rpXiBwHbbD5BMXkXFUuRE/tAgbOZSXNR
8sUSR/LKEe6lGTVSBzHaxV1eyGYlM2OV20ZfRGtCmxgVIonro2GzV76/TRsDtF+D
2YPCP+uYgfBVajepAbsyRg2lpdhc5nqUWbTqYTm6DVLsgSttMQX8DCaCY1VhDq3W
zK8pqFCXYLMUpsdEJ7d0HxIGu6kopQJ4ew2Jsi9WYUQxD1N85QuNKd/9R/w5AFN3
lfDniGJyXUqa2V9WK9YNtX1+VHWsC2w2zBpKzw9+bCeKUVm7IFSaTDESmIQMVdua
I2LUYMyHuj1BUgh2qVqjj/lWOsOxLKyMIBvU14LAX7vRbWj2u8oSWjh9tj1wKo7c
N9ACqy9Xon0yIX/qWRrLfvQzh1YIaeYK5Wq/T2yXig7Ks/tLYr8IIShErcG9Qxfi
k6Kec/TeKjsdSpSgv1dVssgWlMGXlDLfo/Zt2TMQJg58Gy/akr/mrkjfceEbF+L8
O34afoC7VR2bBH6F2cDJxgoOYlyeLasrFgsx5uJv2PmyLsoMZXQ9ATgkNq1eLgwj
KHSRubZXPj6JqGP+EXV0ItIxMHqMli0jpB81ieveVE2+TA6HFGIv+wVtL0RQEiZE
+LEqYg9K6t+nya4inu24FU8ltriNAbQTHm/b2ke+mPrMpiyAKc/CnMy9zcI6FIxl
bmcXob6gTCNhk1iAwAxEzinZ/rjrQvdHVN+LaRjH8l2fv6Jc7NLiCST2jrqX3zgT
oLm/FyG2U0IVjA9YgHr62zzQtJ12e7KaPw6P0LxiALWNL+ZaLSfiukdNmC8ioRIp
57i8rQFE+WWyIB+7eAXNhojdncxfvXsO/rn3xCPbCkthhK/MedZsCzddyd2+OBut
0sqLvhId7aqvjUY+lhjUNlhLNGn85L7nvR9dok61gr1Uizi2GTUUhuQNghUGqeTb
yRw4/rOqeljrgYvsk0Xw/E7g7cNaQ8lYeWJeE3HeWD2cy+rzWUODB/yzDTmT0Ah7
3NGVrhIoImF12BnjDM10pBootKFlLo687hmsQHWZ45bOERPuS7UN8oEYFhDYMLEk
X8zSxFV5nYE0LKUV5YRCx5n++KCSF+Nwz+JrVOUU3w+KuI4YXoEoleCNHJl7EIap
5RqKHBoqn9/GBcUjPObNULNuM6iVGhtoK5sKoRua+SDupefWMm7kHZdK0Bgz48AQ
e4HYmBla/D97Xim4evFxBWmsl/S9LXzUbCnPTEZYtqYLYZL+rBhnQGl/ROa3u3Gx
UK03J/JrXurtlJELEG/Ndva91XgBQYL8TqqZctUehEK3m5Hqio9pNR3ZcvuzGtS4
bFLh/fV5j17B8VrbzhiBlsGwb3DZZps83bDSKTSr1Hb4rc5DP4AAwuIqyegUxora
y2dLSiHWB6MfU37BCOwFta2LryEc8nPOLrgEWmYBMIXkTFqWcpwf36/e5nZt4jlW
0NBh13sjlMqQy60f9hvM4dBTryYJEQsvpofl9c+ojetMXjgFDvia88z8bligHh9D
Qg1gvOv+Yp9HkXsMCl9KCydMbhaLLehPGPvzBl8+3fLEtCUCSJXtgCsyAzTVz7CN
VsSaqDK689juEJ3UnBDVZAE4EL4U3WAtZqLXVN2znzWDHtm1bxloRDZYEZT2puAl
5F0FXDjfkuihiKl0mVLjA8n6EGxLjmmlQu812HvUCvRYePJOwCUOqngFaYtDhC0V
d1mC5aw43wRwL9ttmXSgOwsqq3RSl92RqXwNepYwQZg4eGLch9uVCl/WtBHTfqy6
djSScdAhwu+oq7aQiMW8uw35CiYvppa3M+OhXmQza9rotcvaiESKxC4eE1SJC+1A
PBqGM1fL3RrDO3UqLadt+/q0qAcnLgmIp6t3ztNKS+tAZsAJjMrbDlDmmzcYKZRS
fgDBQkd7alRo89eFoF+Cag0Zap2EvbBqYvbFOayIg5yRaH8pYUFj6A3zd/o9wOeG
edT8Yh12GQhxfEDKhx/Q7JoGIK4NNyQ35Eodz0jim3nWL2PotMEYHULOu70xlMu/
jA+ZyJKFh9P/NP4xfrFRZ7THN6cceu0yu9bXbQNykalZ5TTxjjTRcw7XF8ur3vTZ
vAppBX1wplaOFvrH/MeHPuH7CNyRJyEhMEfT5ElfL9rF/G1zYZGkpF24rae5m6uN
2mwe5l0IKLoatqqaiGBADzfZ1H6sZjC6jMa956YSFm5C689ljc2uNVATMK6WKwru
azxZKM2+dMPfykCFGgFuE7UdxWKFQKUIhrjIRxEDkW8aBYTqwC4RluZkLIdTtoo5
5ngqtP/cAhFZJ3s3NfVaJbq2uvn5EUwdD+ReAutrllMnYKDoBrA6SGaxg3UeV3+E
3oci4xTa4KLAfnqIppD1iwJXWRMIypG9w0MuSOVo3UMcmSojDLlvjsipTuiIgzqA
V6BnV97N7jEVTbu2YefvzatfmsA9wQNOJKy8cEODhr2dePHrVMcuumB2lXx7xkAA
akrMHP4ipU+7yjf+NBe2F6W9muuvM41wL0mIDd8Czqq6qi7vW/V38Y1rrq05ySPp
KXnOVKufIPx4pR1r0yrtFpJbezgrQJQs+tHltJxaTd0Qa6E3hpx//WWfxlaQrty7
WJG15sjMbJICFVZDdrgvi1aBXSkX/fnHssP21QCsK/lg6fyGLJ6ut6ufzqh2/Mhm
A5JOs+SdRr2ZbEKwE0HQt0Yi9ZoVzfLbKQc263EIDYayWqMavtPlZvzO9RKFKgJM
y4+NtwGXrd9oIA8mRbA9NL7ODCRBd0Y0en2s6mDcV8u5SIuZymRO+bvK3jTKwC7E
RHe6wSphPqNRYSgrLChQqQYPqwkHcAXenaykEutZitX2qKJl8BpjnpELua1Y2Dvn
Shrx2AbIVFTvnEbFUK2YNjtIbaUHe5dcxhvrtk5KD4IHHaMHPpO4MM5shFkidlqd
6aLPK5H+5/DqT2tnY6E8DqlT++SyOM3oyoE8bEdB5cdQPUccGu3IqXyC/kFPe4dW
yConflGzPp/vBxAO2b27g/eXtZDpfoRTZmcvM2oqDyGS8FUcPwrV7pzxLZTH5bqP
XyAlU0bYlSHpn3siMicy39IlbHY6vyqs0SuyXHq5nA5k5FWlUrTrV/pVPA2jgfIH
Vs9+W7ls2DvcFiNn88CbQWZmGjltWdFEHfM2UqaVjn6IoyYUS+y+9EQjSj3dksbc
kCAYdF0ZzBWryHiB//hH2aCvQEZcfEH729/1UwzKqcqiqao3fL1Df1aqQKiLZ2TH
1+bQKVPndfZ54pF8id38LC/KlNVoSGtqBPr7ZJNzdXxNcHyqLBKmjqdU+m412tjw
Ut+pXkB4/9UWLcK5HVq0x+XViySMCg2R9RYDUI25MCFV/E1Xka0Dd6+oYPJnC46K
e430jstJLIfNPgZHH9Zztbc1VJsbBkufaRQ++UAnWMTk5CoyEZh6M3uQfLCrsUG2
fAiSmaQtpk8OplLvgdaxwbpWiUA3Aerggwz2PVeE8di6YHbGgQMfM4WkT0/x4+fI
6ZNVbJND4qlEDax42Xb+a37ncKbNdEWYKAAnlin4YO7RjVF5RU8czEX6ACNczmdM
AFPjLA+HVseMPWx5VT5tqEmFMhCqZ8qEZtMME/5H6y2ED3RSRIkxSF1vjhS3ETpu
IWST/DAF8k+u29Smgszj7j9XLqkc1fismdIvz2guQBynSJ8dYYROtNg9i4BokXNk
lPGlwZP+fwYJvjTlUxH346QOJvc4pTkyJiyznk7rjXJntjLtN7r5Wl0vbtciAK+4
u8f6rayE3FA9lI7XLTpygwg/tNTpQkVK68ezAUL4lzFcqjSybThwpF64oJ7bsWdT
mv33f+TfudKB9Ut1ElDeyZYVwpc/7NLyTkZ46/DHfz1dTjEqtae5QZCPlhW9d+Os
fHoxh1AWt/4+iz2kNIUqYOHKGVu3rFfaYp7bBLqr5DkCVRML4epZCHfR6YhWoMdX
y2rLEGK+c2zmk6LvGwKxnBYa3zRE+G4vtBeJbD12vuyXjyi0KPpAanb5vG6KYM0A
DetWRwDqOGxAzLJFIYt0TJ4kDKwntruHmAP8B4vSm7r/2NJhNXMdoekUKSp4w20H
JOE29CrM4VWY+868JQbBjaQuDFa6UEWF5YiZCAp7XUaxQCt05WKoo/uobPHyVQnf
62DiftJRwNjtoteDDI3YCou4EvXykXy7/9DxrpqcyW/HiX5NMJEJjZepiRo/rFxg
S/klSjfu5HcSVGaY+BKhgNau0nI6vR5FyEsmslcTfTN17DHqOhl7b6pprwhRYVEW
Z//jdtlqNx8UzeF8/8sb1805BhPKzjJcyl33lEncrnUJAuRnXUuxa9/GFxb2bkmi
ND3qZF54ZjSZv16hDNM7SrxEHHgeUf5TI6ZjpEqtOQy6KJ8yExU+8QgotwiCGXZ2
E6xJAEB7bPLkmHvP5lV34e7gGNymXF41aM5AE2iuB7r6tb8Ekfnj8wTyhYGKgWhk
PNju9AiP5zx1Xu8QW8YDNzH/7DffOgnzBRBIDUEgb6ZtDDNqtxohyDxZyTY5fhwZ
/9AcU49YVPecDZDM4r2NO5EwoqSi/EXO6+/9eK0rVFI7lechsLXeMVsRijM/H+CG
OdnoRVPD90VkFpH6NRXcGAH8qDQs6bh4lSsk7+vVaIwQ62ZH7vUu3BOT4mQZKlJr
8XhK2C9yoAblVC0JWaGi8iUSUsbtufehBeBUDcXUWkp1+nba3dmE0mtUywyn1Nym
EzJ/Y4j2xyxbSvH6PqPYOnyH+B+cBBGKV0NkdmB/PqkmkVbHXX3Dsw1o+kr7vQ2s
VqhV9dMiuHJtzdnnZTYm8hKtyIIrMvwYosm4UsN0+vatZ3U05inHUDvZZMexHM/e
P81W90zzCXUNAClgSdaS6232lNPayBEthMDQnQ0YYC2zky7QkqKsR0f7Qlt6O2JK
sL8ZgcArhJx/tDxlZLHbz1vlxBk1USKa4rI6ALRYFWv12URldvud85Ou1ej9r+9+
DR4Knaqho2oSUB612ltg5RQXSuGqIipJAz7MUliPQCgZ8x+StKErbU2zuNssDNBp
VWIU9jTRf6vbJ7Te27bEyFblALg42xK9OSittm5OwtKXeySrbr+OCYIF4mD2H7r+
89BhhIvfcbG1Ecr5RRzlVb7MdudGWrDixRjbPsbzOEBHlg0Z58S5WmLjd8v+vvxK
5hv8PifMAAFTaNN6g3X6oOWj/glAgynuB4pS+gZ9PA3MJWivecKlUt7gG838mlR0
/Pmi58GJo2FIVdMOb1B0cgX0umsAdXezba5jTaqtI4/mCIHV0cWwzo1GnztSeTzv
C5SAqfNJQU9iJOcH8vtTVyWfUENbBuOOdHPyXJ25NOuucfIsnLmy3Rvd3A34sGVx
bjI9gUGTE7K9Hg1vbU/tfHRyeD3VltWXRGVHx/SxqeSnqa6URG2KBcdNwTbXNyMB
jFG1AxK3vkbWxqWORwPocEFkfIEXbDTFQcZiWUd7xr3/k5XDmxsaH70ke8Vt6SOR
ShKXlCj4AJVLSMJbyWmW3hXYY3BNhW25ugKusLcBqPEBkh2uqogbxutdjC3Pjqnj
NANKVZ0JWXV39jsX8Oaw8p6RGGkGhWn4m39DKrDUOq+Qke1Wanf+/kWkbit7n2Bi
KtbRtUotHN34Kmoir329kvUgWRB3G+qLmUU9XgqZ5Mqz2bVK49qAldr9Ukey1Ak8
sMN9HT6k4r1WTSubPA+GO95xifY+8lVOhWQ0D1fUqm+BjmrznJWjKeT5KaM4eNJ2
b3ipPEZCQjDbFVuO3GQXV9GMRmV4z7+AgxA50fGpuESTdS1BD8hOVHGZ0NCjSTy8
4/gfIYtr2x20sDwgRB6S56Rvcv46oQAsS3qyzRywUqNTbIbOEQgmRpuzHNfOOvlv
loFnVr0mCdRJqNXhpnTh+asTj6sHYv8Z+h+Lze+GScE/yoMKvHYKBTyOCPmv1gQP
JNHV4lb4IhE92fFQcIGHpbIHRS3Wn7C9U210hh4ISRqpVfEIJSuTuKa5GR9EGfLr
5omyFZUsWSPlbvJAxQ7pDB4xZRHpB6upZ7VL+Wba3rKmoEo4EYVJPDTGPitZQSSD
AXroHLMj4pG/m2ytxczHKYsNLZwy7huUdTJ+Z7VWPsOMekJLEEBUNZB37c4QAqvd
8Y9pb1KVUotO4XID3OitWaK6HW3vSYMquMAL1RxPCRMh1uR4hthC8iYv7GOXFeeJ
br/WOjTRPWWws3CG/C5GnQKS4Z3NMr22ZLwCf4BLAD8HXZGgN709dcKVLFdxYREn
lE8V4CZqQdhMF1fq05MYScwqxjVhzzV86rqCi34GvR+EGHfSQc9evshj9i2HDYaJ
uWhuOzcmS9TG0nH+wJFINBsAGoB6B15LtaoFfbn143NHYtB/YxXWw2H3PCns1IBm
Kz5WYuVN7/6L3uLvYZqHo5YBQ16QCQDJkEafdsARDbmcOWj+A2ZzDW5a/nl37Yvd
O+n16X3aJVx7Z/NRPTmnlkdi6i8GHwbP6IXfB2spffMrdrZQzEYJ9Y2FkcoyVhN9
rDgv4IY4vRMB5YFT/XChD6mc6wrABOCHhPahXzVSDWdkYxcRbzVghBhnFf9hFRZn
rxwMRO3IEMyXSUXDffqjXtvKVZCSCzTn/XW/HT1kI6Ie5wPy6wVzZaSwC6/XvxHU
KjieXnojXPJhQ1AHMFLanj2ol7dcgiFpoMsxhlUYGQTvNEj9sW6VVXa3o2CblJkd
BmWAaNyaSASS1jXDTg1mz97BCO6+9aEFN28E0WbkmgfGoexY34ozxv8C/MkcsNBa
+xc+lKgt1UVvC40i2BjAbGn1jLdiCHeMIS86le1+XyOK6KE1dK6ggfLJYbj5MDOT
d5mRfRSvGCZTbmsSjSpMECLcVnWLLD8Q3GgbaAfh+H6NHpnGtcTfOBMzVgI7HEWX
LZtu6S4nDtibJu+DyFH+OJg0Ptu8AXtOmlcl3KzDJuWTiTjFwL/W+gJJYVE7f0wL
2jf9xiEUdykABJ4IgOy2b+IwYdp9FEW/ZFdpiSxlxBhfQa5tG5e47mxhYaont6kL
xPrcgRJmoHts3zi033HellBBt5+FMTcGc1UUucAlKu9M+l1dtvZqpvlAQxG5GMB+
vjGbsOdaQvFJUrcgwaNzTzbaE7pbQTJThz5+IR3jwMO/PO3UzC84x5wO4yKv6QdD
h6ZKuocO7/NSm8co+cfrQAvFrcweCpPaj+LbZML0La1oQAha0xxm3w/iH3acuPWj
WgzOZvGu1MB6IqBTACUV2ClFQS6G7XZ3sCICjTbzjvJO//tVcA0x8pDFcWQctxqA
727ZMXJqcdnU6sSu2kojPdI4Ll7+1uIkAvJbxjOsYSwf2EbqSQr2+lARzZM+27kI
PCC4O7OVqYbKgw5xrV0YOij8/lzp+bLkDpELoJAR8eILb0wDB5ouT5AoTiSMMsXb
ZyhYC9WZPslvy+9+d/Mif1piJf87Gdjn5qOpbwD4L6LVJvvdIpK2hsw9CXxNebaU
5sHDWt05nYyRCyPsDBvaH/WGstR68laVs1J5UBxxGgmsNjfy+AQNvPfHP9c5Q0RF
JkNWcNyDc9kuP9oP3Xh5yadXh43mQT974mxPxZMI6MyKgDhrqAdjmerO2FF8mStE
yp4KVUt0oMSBm8Ijz2K2XtN0Upoe7gr20+MCJH6Jd6m5+AcZIdbdH9ekExVZcPew
zjMtKLlmDJV3/pSD3+Pm59GrMjwCI14UI5Wsn38kuPrnaon8Pjc4hcP9COHgWGlM
+tRRqWHPnb8V07r7KpYsWMWOmjuj9YeaWFtIhEoWUXpu1tHE/yXDpIGhRFcINVAG
lOXOR5qyc5+OFTLq7Or8sntlGeIs0viqlQrkVRZCcIs0JVXLZnluEvS/uMZxoaiC
xv55E3MPnJgfl/R/+zQ9dw4+MYg4rCqc2CaFTCNhcpbCs9rc/H7l6xl6Ang/bQqz
s5ki42ZmHuwYLW1+pahSGsV3CNSZp2WgAo2fs1y5t4xNBBHtnS+Subw9wk9MxTKY
aqnTjl1ypMp0kAQoUG6aRMQ3tf4V9/e2/JUKBHtegr4sB7AvlndrszEOXczXTGge
kam3CQvmb/n0VCuhcUX02iLMWoYBVaAhYr/kIz5QSdMK9qiNJhsJAfquLImtdibe
UxaNYjLFam8/fXHzdif+o0DG6txB0Qj2VJqdIdQ5ZSDDrmWkvXdxiBgkeFDX0tlR
RA3rlwN6tWNYPRn9FCtxqFhfUIs+2/l6h+kBCWiQqRKAXd3w2NJcQmwLxABOJjn0
dWbVfPiBEENxpRK1tD7JPFtaeUBLk0O5BV4OzzuSMNmk7Ec5RSb01KHAAZUE7kZE
sJ61KTLnBWWuDL+bhrPJdaGhPanw4ZtnJ6NvgDITBr7i/Trm4p6rehCuvQ6FqxZf
aQS+jUf9Hm+O417l62pihDja/X0q/JNJPgKy+uP16X0RVZN4eT68YcgYrn8oDtTF
TB7EVX2GEJr4ksiIKt6pVE1KSNsrrnRZy2O2hCU8eG3MJlwLWlPmGo0sEWc340hY
FbJAe/gwajxI7rxUdGxnQAH5Be1FfpWrsN7Qo5K55WsFwEM8KXRDFBdgZ7HTfyVg
tixSPGISd6hf190NlLLrLoqJEL6d1El1ECC3VBE56/6U27cgaYDPP+fE/lQ9b/+r
sWnP2QvGAeLhq1lDyfIKsTQHXLrGCfQPogrIbtS4ABtaeyZAfz9zRmo/rCAbEi8a
afQyF9ggKFAbVhMpEoU6Hq1kRCyXbgJkkFIEjptCVZfm/kYa9xEXamweOJnpKfFY
6PYQviFq0XCKe+A+mPYEmmJ4uzF+k1CLlyLlhtmsVzja/FDeTbM6PIonB4IB9KPT
sSALbSmIk7n3dJpMQiZNjAlV+mjz37F4A29rRIkMC5SrEpLl8CwuI/CubccHUFNY
R2EAkSH6wLRaypm60ZIIayLQeApjdlaCCMEduag2uTUlfZyi9WXUI3iCL1g6kGqk
jdt1EgzqBAaJDpf6+SijeEGUpSoX28VWboFo00O0xD7vPqgc3ULkRW5eN0VZg10w
5N1YWkEySnMGil2nOKY0Qh7dGNFZjjTc+JRYY4ZXmNAdaAJczPgpr65UDi1O9aLz
rPcBjhmLc6YSIFt6cYFxA/Zu1J9zDNjcB9TVvd+5FOL838SlDNi0S0y+nyVkR693
PKzTkeQAKVvaCPP1tN51inFRmQ3fmyTb301yqYAy/1oyJdp3q0NMGWd2GjSUFrl3
1qmYDMHHV74lTeUQ60M0vshZ+wGsZR6w/sLS4CKrO9yXtbC8VNizsu41dFa4MH6i
RsPxk1X7RXCYK+5WpNBmggYmCo7CxzTFsD6HAHao6PessIN9EhmkNJEs3YcvXenx
Hfe2xPIPgsiH5uLqnY2L9jkGytPcHHuyUZgQzQ0GbCvhi2Dmd8glHr3FwakxU0LH
r7OUBj/k+NmCCg8RKY9LLn0vK2o7oJIgPjUQcQ6/SOhk8vy/nn/0fJiWop0n5EiJ
rXVPQ53sFX099U76TOMaax8UAuAhH2RgdB//3Oyvbxn5FywVJKjohSs+skj5JYzy
C76HiLrXqz7lv2Iixp+JTXYSabpHpNq+PSIPkH1/H0EUrWshWu/bS4bxcuzSNR7K
XWJUG4Z5sebEkQZ5fM13NqsRInZNiDwLs6bKiOoVyx5QW6Qox11ItHoOyrl41RwL
NB90YQ93DtnmFyIrXdjreZW2tKvSPavLOdONvS5mNIOFqp+hpCnAtJbeJ4LlH7Ug
/Fdehtwk+qOuxy4kwHKsNt75i4xMmN6OYxNmIAstfQ6+Rl9YMw+9B/jAsOAv1cJM
g2l7aATeA31hyFGA7BIqp/WtUEFhujCKQfRDJFsU+uEtm3X6irVe+MA2UwXJ2PXW
Uon1uk+mGsy+0opPI6lOIkog+HPn6EnW7cXTpxf+oxCO25o0Ar+MGDcUsDIPULQX
Z8UkF2w+q2XTfW7NZqD4gJvZVNt2Ir1YKoNuXL8EI2zEDipE22+WUGtJKlIVJUSN
2emMARFxklPYb5T0FIz+cd0Y4CFj9E/C7V9S0KH70C0GkNR8DeNMDGHq5veDSdUB
WgnN6ffZi+fIUXjVpZhv+s6g66YdCKTO/S9PM24o63YH7bpFzdhiyeU5N6cDn2OQ
aLG9y4kvRVAo17FG0w6Q07JasSgHdMgtzURziyrHIT8dhYZURkK494R+n2LaIwVu
mIFdhGO7wyJ6G7zyio+y1rS4P+xoB4M3Eyd4BgWGuLFzSAZvUQ6B5xTNoLFNFN9S
vSCve/MhevHpK9N1IO56ZbyClB/v6GXr5UZtWB/Mb6m0iLTdPTY3ueiNu8h8lvtj
TElKoGYV2zLTu8D8wBj/tDCc2I0DnZfqr1rOGkld/caG7EPoE3Al20bK5CmwxZXG
/1Lg8lxgS6/f757+/77u5FOS5X1uFUOVkDpFUuipQxSHEDWuQ5TQJof/OFVP2CLM
xk0FPko6y7jezUj/1oNWR2GpfLG3yVZGA88DApdMf8qC1SryLP7cxBE30B904WFc
x2c9lHpHtmIrbKEAFN3PG93SGutYzFUVQSZBu2LDbUo8YKd3K7BoVwL6o9hl8aOS
qJDs3R1NcnkXg2jfnRyYkvcWz8YnxCWD+kLRRHUumhm/dA0j18u+LD1XUu8c83+u
0QRBoEVoPbZs5ahTbagfsRRR/1wyBPEl9a4nOE3K9oSLar1go5yeprSvwopyn9T9
QstHQhDgW8Xgg5VpPs9s3MAwOhYbKK4UE0DH7HFfbGbjSjoeCHCW97x16QFkuZDb
RDOMXY12kWIxlgmCP5eaZjDKseS9rh2mnLG7josqhCTHjZkNc4vNTHLx1uCUH6gm
qV8JK1ZKbUp6M0kEPLcUBMYKGJvQ7xA+740DTFTABRp+B9cYCBKvKlN2vdbntoll
YJa0f/rSiESeCNFJpBH0Ma/cSv/tcU9TAAQ8sxHL6KGu4ZOBMp7bdAmxlLiYqP2j
b8NvOBvGJ2Q8hNTiXidRfT/CtbtRJVltliuIn312iKKJqhgA6AxzF9MG1m4LUKIY
AdzgqbUJSVxRqOgq9PehXoH8qR1bgLrOgFILDKA90xm+oWbGbm6yKYkjRs8+RZok
1HKVJimq2ymQ5is47SGJf0hWxtn/DPQZy8CZbtZIZo8GEIUjBJ7Fgz19KqeXbrAo
duMOHKmC5jIrrxN+qWFcovBbQOFlScDVcxSpdZHjyypLNiiMf7e7PMOnb1aF0vQC
l2OmXxYs5xvidTgIBgSeSiY4usHiRO3aUTvgTScYKZ0IBE/r32zHCle08G9CV8QM
3q2J+Fc0dgzhZT1jFFGc8nj8ue8RPmp3rRVxYV8jLbogkJ6hphinJxj0gnS7OP5m
x+fliedhHH1Tk5dCgIpyMl4eer2nGAAD+2SV9+5FpqoryrC4xcsPanvNN4pwnA9t
7Uy/Gc/KIj6BL/EfwCAdcN41h7ZnysxOJy4hll+4FKuoZM+ldIarpi58fDm/6xbj
vQo5VF6obe3MiiIeyMkMV+LPVC+F2Ox19qH7YoLiZ31iTHbCGfRt7M4EEhgGXP04
yoxEofJ5gmkNJ5u5W8auOJ/rMpzsnuKpNoLXFrOHTxFRhZdpwgt29+0ZNGBHYGsm
WlTV0BhXMnoIFMhby9dHY7siu/PHXslp3G1OVPA3y/aVpJfHpCv4UPvMfoNGAYJB
RXn+NaCnn0IjKjVQl+1tBzJjYWxVdGoL1Ajrtm2ljN5g43TiJOBIpXgzGYMK8ETr
zIkqqQm7ZCzjKzwIGpLwxF1alMFJtV4y4iejAB7U4mPs7GVIU3IZMkuy2FXVn1QC
5Wlj0a+pntqAKzBosZV9uVmsyfyxKhWTRps6mUvQzqaO5/Nwr0rnteMqenfKCl9W
YbkyRQpzdtKteTO/c+g9r5Uvv5x4gWISUI2+BArdArPv1YLLyu2/74cUyPuONCio
+PkXISkM/CqMrCqZmViRZULg1ttkdQSY0VoZwFXruUfyjDTR6pjh7hcIVa0DNlp8
wKcqTYLL8yPbtPrsGfC6lVNFuNETDl+pGFLbz+TZnxfr9xGEDFZzs2Keukf6SD9t
+IfJEjdRisZ8zArt29Se4n7wZG9xETRN3LkE8SyGyAEyFT/NF2TTEAvihCTmvswK
iDrMc+9zldWxOIDwSwuhtiq8J+zvqcr/TBCnl4+Gb51753NxwB67JkfJxGEWH8eu
zCB8XqPEzD3PeTSdYc72nPKeb85KNOCbbJGjR/l3xIMQR8BWckhNNc0f1rz2e3fm
3YmS9BUlPnwNqwfxDEqgDPIzcX0bzrRpp+Q2bmFkbpDHB0O5vlXTC2SDFTt7FZGe
fpV2W0VhJAMcNn+8aZQnwxh3BMx+3dcf/LzvliYsCjXFRHVYstIXr2tF2fvck+Pa
Js9sPwum24upBoljsCxgLfNb+gMKwBzn+5SD1JweYPd6IBabXxtAQ/Agw1d2/8Sg
bSXFH7S/9Ij7H5xtgEvn5Cs/8GFzYLZ3fDpkEOh/1E3xweTggoB19minmIZGati3
48TERFhOqXnpbV4K2A/6AYO9GrtFt6rxrJMhSTwXJSq/ijfykwZMfZc8IA6rBg6m
nn1yfnlEfh2ZeKC0ugksXUTTKqNIML3s5ksu5fDz2nqZXYjZV4pQJ104M2H0e8Lg
57XPEseN4oAyJ0ZBP/NyscUwXmsfjtYOXhlBKA7Arw1aJVUMHfsI5Fa7P2rue9MX
mJQIdSXMBFby3TpxtsiBgI/kmrJc1ZZdOEtsMz/bPaCTysg7mWBcaQYQoFd3FVL2
WVdK43/2WgeJkiW2V6bBpHlBcEOeN9B8V2TztVWAv+wyJGst4c9Zl0EDmuS95odV
xSpKsBqCCDhuZr52ljeysADB1kp/RJrVD37npIoDDRSPRve2wgK8WcT89kpJVJMo
JFYcUD/cHSeK99fkKGcQCN9w92xzRajAp16jsFvB+2qbB/HjAzW29LeZElJDJ6UE
gnqOZoSuZ7u/Tpfan3GGkblebu3PN6EQZp8oOHO3ddurei1I31jBJdyw1HV1Bsno
XP3wbahZomQvVyXQ5e6KqoO3++fn1s4f827SYUpRgL6GuCFJu6bhkmpHn4Q0sBV+
xFsCgVkLTAfN0gptuLlfOa/yaFBHdoG1XniSGa2qI6YTIAmrA665iceyR1IqzSs/
eleHBeBz0vaGPV9T9dn1pzVd9jicPTNwu2g58DwKrri+gH4NvGaGWSXd/H0kiN7G
Ud02JgVoBZXgZlVESc4n7tjExM96YcZTgrRRIzYbmn7AhRJ+YCQse2VifCqYrl+4
Om9jeV67kxGnzvBx3JIrIlkd2mh3x072cuP9hPC38UdN6zoRGu6MjfCcdPtQHUi2
fmVpnK94aKi6XF2DQu+EyjvC9tgN2WA7Cov8X6aLwz51VstuTrRa3vhxrsOApwuv
6acRD84bLktL1fHbPlwHIcb5CZw1aqwhP8ggQoFywq/FAW0sseUnAYl5X0RsKmkE
txYtY6IaDL3ng+M+wGIdAKoQvbpwqnhemnDhq4nzaT1It6GfDi+3PnpDsTx5YyQ7
TOPM6VzR1QUkNBoO6gHb9KUHZqntArzVizdO/R3sUEuus7jwLa+8OYhl4CAMQHik
`protect END_PROTECTED
