`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RXmj65Uk1mLVqgolegKvK9CMtu22DOsZKbncm24UeOoX5olgOmhv5ukwrDS9bsRv
aDPo//JvUndE7fw8qYxvqJRcnBRYSDmG+eTOdH00cv4ZsFVS0JO3lyMTA5bifksp
+PmtBx6i8XbSmdjqfinFh6cZRVWH+S+A9C0eR6b4l7t9DMTREdis05kYAzjOvwxA
NG29Fr+zZtC2UQ4PVOauDQv2S011CECSQkAGN7NgiCnQ1siDcNttTB/3prKVIskf
BrF917neMV5GVNUtDYbfy46RhCiUNXxlCV+6XHCzkP30ntxk7DgixMJKaVPu+lJL
j8acT/V1tjcmX5xHlgNAc4rzRdrv6Jd5GsYDhKAFCcMxnb2kaA0HbqTxv/Sz4jVb
q+d20mh+/nzhYoBi4FjnJmimy35L+bjj3FTSHf94viAwWebb/qScWhNbb+XWoQ4S
qhn9XnWlzZJVr9Ilk5L2j+UxhcfzIKGyZTPix7fClzr+pGT89waETfJTi3jmxQa1
vq7sN4caCKK+j0WmIInRDjrSK5Ftg8jJLRhNKRiaeEE1XX4yFcBJbtBtqEhA9LlG
SkUj0JG4OjlPfIqMYl6bH+gKLfnLZHLxtPtAC8uzgFCFksuVZFDPrpvniZ0lV+ps
Dd2R1Hqw5pOp4Iedl/MzkQ==
`protect END_PROTECTED
