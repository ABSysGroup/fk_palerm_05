`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xfYasZwkdzhXUR7qK7wIMRtu7xGIfQFHfJQ8Yxmc2LNX07QYFadyeNQgELY+vx0h
UtTygxXRhcO1NWHQiBzREQZuQk41nJtbvjuDt/kHill1Ju2rBMkPtAbYmTOn7xUQ
C2uDQwADCrFdyKyjUfQl9CYgGQv/GlvuarM33pCgHg/iBhh/SQubxRlyRwu16RXG
7dqZnMug9ZTDgXeiGIygU5UD2tkWKbf4tz+kQUUILLok/4ZLTc3nVIvIkLbcHGJ5
zV2sfwWVvZ50zV5aSnDqpp7Rvtnf/JAZnV4Q9naUU+gnM+UdfuR4TmTZ4tSv2DJ5
O76pw0uqM1jrz0QsqUcqvE1KDifcmzm5cNLq3SUWfA97m1cMoh7JE5UCD57UguGo
7KXdcwgRZDHpyiFWweeuhw==
`protect END_PROTECTED
