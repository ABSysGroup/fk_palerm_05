`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zT8RuOfJNwLtRdn2+iGNq8/NT2nry1V1EwBl3vByQL0I3EKdj7AE3TwRTKkA3myY
cvDBXmndJ286PZgJOgX6I1sUGIUNbUDNVZUwvk80fN356jGCQz+HtRmK0u6c0QUc
FBSJfjNbSh7rPx8kxdY81Dv2PzFlDqHr2wNkG/TO+4VcLI4LUsh0mueC6SJbzK1J
Ftx1jC5S2aYyjx0vQjwjbMiBMGVsIgOF6/qgChA4TpMx5cNKm+058tp+5Xbuhm/I
aAZQxQfzDCGCNzM5b5hAFy/2wfusCqpvOTuPrGM4P9Ib4KNY9V/TPJ9tLukL8hYo
rvxYQLAhJB5MvazHHEA1b6dRASVM1wJmDpT+0MeyurOmIXubybe++1yY1GDS5dfd
jF3BUpggD3q8AziGm9SbKv2UG/R9Ss/CCR2lewuHmmt/teptHD8iz/QfPMGHU3WX
y0lc/1pai4Beu4vwr4lbSLjjT6/Qe+iYYFJ2HVzHQa7ajliBStfJVdTARln0sdw4
`protect END_PROTECTED
