`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7UGVRStO2puBrrXQSiUEh/LiCm9GILHpjO/VDMcdeLW1ZG4ejUJgxTWsertk2y9i
NGETLnVhnH9SEF0x2cXLluARtJ2RlV0YsW2nbUIU6e8KqmpwUkJhWYHSClR26qnq
v8jTLTeC3vHdR6P+FEeXJxpFrS6odjzt2JCFncJUpco3F0DAvQAHE88kcpj0lToW
Od5V4Yj8IkMQBrFSRzbfcBRM4fuZ/5VNYtKOF2cZAQPaPdtx30Sm75gVMBLJ+uON
3d8uUi+6VwVO8bZyLx74WuckvV5vH4q1zSNrmKt/vAoZqxJZp+P4h7QcPNc3fyWf
FeJ8dXW3Tm5Tv5IeE5ljcT7omQXoh0CEZozPoHH8adfghk52YohH1QBHMSx3zHn4
crH7qkmD/xknIbvRQg2qQQTIwWd4zuxIpXgpgvXWIAM7zI7wf88hpnjXUtbCjFVU
k0rGswi4PejN4YFZ4HJCrg==
`protect END_PROTECTED
