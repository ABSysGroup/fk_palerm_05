`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g5XNFtJccW0SW0vbCzTVuup3o8UUBEG1rJ4G1tQHfu3EawXUOAZP+1Wiruty4sk0
esNOxwsvGRydX/ZwdIYrp8V1KpE1YjFz+MOnRDdr3OV0TrEQiZUQZ1I0dBPMCiO4
iRmw/RnZa22Nb5X7Ilc6d0G6OtwitbtDrTWUm81qkeTUZ+0onD+MC4h5fNEKBr7T
37Voc2GwBSva1qOg1725vSWmgw69kVKjFSRKDA9mzjn/Wnm+CsPGlC4diphy/0Je
`protect END_PROTECTED
