`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eal0MLGK/0HDHeW+vsM/1KrM8jwcqRU73A1fyp9AF+nBY0F2UrZZUVd4JxEVqjTj
O9hN1JKM+QPGDsLIdUOgoEet96CYOQI0zAv32NWnpkeIpOMYlXOoj+zlXNZkVrHM
qrPfyfrtfqfDwsgJPkDa5V8w02gKgwfa3L1Z8Kj+8Phv49cZtE0scy6BTFREHibs
pY3snWJXAHdk3wiHrNvtkn+obo7JQFkKFiqFRJhSLmWn7KOsyUFAdh5vIzNWmGbx
VKc32a0zO1zmLM3dT+OVjo6dGjjNMVxC8ZpNGU85fwnKYteAsqbAQr7ZqLRa53pA
`protect END_PROTECTED
