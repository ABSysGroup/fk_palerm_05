`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xbOPr8uXys+bP/PeLSE2e5y91b1t9plZD8pjgzHelBCiP2p/acBQMYNopOh+4rrP
0Nuq+0KaSAiX2p1QlF7H1YIIcMp7rsD7Z9PhwWPdsauf0Sjwii345JUrYpz6A6Fe
qvZrTx9A+hht6huNRfljWpKadUhj8X/5gQtdsoYfEC8i2Ip/ascEI9B42Lv589z7
TvB/7s3jcQTfzpFJgSjQS3WCvkj5KpIFje8hAHeR1rEJwRtrcIUKZ/8IJhPQ61Ae
wdHEbNIAHMItXZCIHACf/g==
`protect END_PROTECTED
