`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jhu1u/PhWWD0K+WVqmDfQ0oANR2sm2gsx3QtTVA+e382tFTOwp7O7NkBZMc9lrxH
HmsU1G/flXkquWXGesA/2SCJqZZMBC18n2H91XF4MEb+YSy79Rz5nkbVryG4fnUJ
eInQl162UN8tJDlcEigcXsM6jvVy9HbFnKIWFiojl6i0HkPEoccgD9tptIZBXZV+
R4cXBLAKO/YjdEl1dwQhjSSNE02wfCzA3WyYD8R0LoYIOQOYLbfSkn6NuQykFNIi
Exl5EFqhhBK/Q8C0wKdmh7CvIYgViZJqNhqtUPdca43YhBpgh8QgU0Aj08c1EfPR
4RVTCuCCOhkOlR7M28QkHwZpJ1YwQ2a5Tk3hq2UtXB5RKSFh9EL9mCSaAMJxMa0I
aK9X6QflHlXXwsqU1/Y3fKIadicQdEIHPwnEyn38lhQvrIDvd2z+EsUi4gWLO+1E
cPALrtuaRuGvnnH7HKfi8k1BkkZNtMBfzwOXh2k6HndTQCl3F1tFByGSEneU4DON
mnd2se7AsQ5rgP/KF1mh6ebeM9nGXRIN9hkSl61khDkOE65TzHL+JriLHlxJkTOp
uIddc899R8RdwDdqYJGmeLhBh0UOjFXkpW7Fws1atSw43o2xOORae0DbXSrh+tHj
kZnSAoLqlF6y5ymcwgductia4diuuU8tWEZy9vkz3wylI2JqHTTn+frtid0zvht4
EqwO2XT7MeuRk/NUVUthU2wvv9Ozl53EFn6H+AgrqerxGO2gxO/cD42R08ztYqFu
Uy7igq5lt4HP8McnBvrmlEVaZUllOZKW+xl9SvIwFwRpR9i0bx32ttgNWMCe7aRZ
9sp+r+RJ7i527hvlRufAzdbS4p7ufpkIb64nJ1ZXLnwdms1j0CAr+nnbGcAikEQ5
OLhJJ/i1EWvgzbTDGxPOgpcOBtdv4riltdy0NiQ+ZPA=
`protect END_PROTECTED
