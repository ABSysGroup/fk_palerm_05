`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U5Gn+9ohbgvZnWV9mrFzqdNhGOLk5ULA5gcO5swrxtZEoTe+daYc0JxgB77ZpmiK
aJKXzcGw44dZO5ogL39WxYtKqBNdxt/c2qPgrs+VwbdJbck8XaaWbV6DSCegPsGo
AIMRYFHiozc1n8eH2vSfUNjgA2OFOb7FJ7Iw3HMnS4pcADwddtmarUiTuZCeHnqb
ncWUnE50wilusAul+hYTeY4CSYFYyZ+9r7AlIcsKC963t3DWafXiTohQaMdQNUSi
QXidpmEi5bYWDFB9CEJGL1tinS1o8QPkPK8WsE3jTCKG+VkPt1atDGTF92JUz+t0
3S1T0rnS2EjWG4vGu0iFPFgqJ64SXI/dvC81/Nq5nRHHIY0BX4D0LxodFl6zo7Dj
X4LnJRoknWidQuvN8esjGUj1Nx+XhNvYAhSmLiTjewH+LsebaeY7pgtyjKt9iHs8
PobsKPtXEpguiEFPdEvxNbcjJQNbjybF7UathYDLbHsCq1iAcEsnhmOtJPgKeIl0
McXAq+ZxKefD0StlDsQMEib+Gy6NZ3mMQaokEgdjABiUd4Ov3NAWwBhBCCLYyNUT
2thSQB6lLDIYPItjOA9ivvLyf+ZX7Ne9XAlI2VLGL+DcqYgjJkWZEMU/PQnDi17G
oq/bYLHIlUnlA6nfDMZ5yElIgP76tin9VO8sd67kFqwdujf5RmjgyGQiyyn2yanh
sIR6cGq6rxiwXeH8GfojBSO2eV98pxWlyMZ5BIZdPtlzvu+qBqC3YRBbxzAfwwqx
q/XPsKMdnoVgyOXLLULXuKBIjjBHHlmg9V/3n3O8r7UZZPUBehgO4Ph66nR0A99i
hjTptnVU305bFpCa5ILR1WLv4ze5StNRj0FRJwFWNgSagG9FXrAQnG9A4jmr4wmL
60z+MBlh4oiq91T534Dr+zFDKJ1KbC3Xl4tSVPxL6+Dujj4TG1vMj0o2YxtDBjc6
YIQa1hCWuQEGSA364FnUxk1FAJfBu90cCzKUm67R7w3fmTaZOI8N+9yzOwNdroWF
OAkH7EIv0KLPz5juC52aQQ==
`protect END_PROTECTED
