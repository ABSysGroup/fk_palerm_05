`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l4N/pykHjB64UfiPWqx1aSsG0fcTfAPRWATweDZlfyl06sWGGWl1MbJkqj9oAmiF
aHcS8HIQWmurThbgBsD9M9NbAtMtFBvby+czLgw+CI7AnZJq3mUE7cu/G1w5ff1r
dXGjCNYeyrwsq2Q+IPuc8PzWEUvMvNVx2Ejpqu4POUxRRsaa+YSsk0EVH1W+FKCR
lNDDziCytfZ789rNBed5aIAyRMoeesIS82Y+d2WZFH/bJnsmzQWNxkG0CYtmlkdL
FqnUpaGmSpgSLzv4GUIh64XtQlQJX7D/tFBuA24dLST9RBalXNZy9v9vC0MAeMnO
xA1Luz2nv+mpsmmBVmrBH712Vl2hFtNc9vlsMWACn0ogdxeGyy67y6c2kn1YuCMu
`protect END_PROTECTED
