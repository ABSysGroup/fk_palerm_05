`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KqdawKH0ZV5GdD7O32bW6D18a09Qq6xT9p46lMBG7OsOJg4CIZ6lV7S/qa3VuUeb
gAyk0fLimnYv2CROJeXke/xUhY91qPS5HyH2ScryPiD8t8t9r7HSStrf2xrtu3x1
JjJbfZh5hyBrns/+7LUEvYNWPDzBsK1u8e3TxzXu2ayHgxrRCDXyXGKfiL9Gc20D
jySI71Ayz03mFqYlFy752toW0VI9xQ107XEXWpcZZa4w+LzI+rRvaxoDs+an0y1a
9/73DhVGCBNx5QPg2ewzsaz/N8cgN0FiqWoaFV6RKnw2mJO/LuAkRWmghVFA20fY
UM8oJ4FwXDLw1gb1f46Yfnk0D3e4ButqQogQgshVr8E49X92gmgSgkpyXK0EtSuC
2ALIIsM4rjONrCtY5GAdt8Z2ATriQat/jfyXPhiiD6+iQtyEj4fxK/4ygTeaGQiC
jWhVS11SelFz6NXukI8L4OCNK1fLMqqJVV5A3A3puGtbtun88UKIdDIE83Pi8iBE
xkFId7dtz26+tsDHnCGEIMBQmt7mlN/PLOOUI4LQDIyr9jGYqyz1RvDDF7PSZVA/
zo54PrM8bKi7BKZLYipw5+kBRhfZzjp+ihB/cS1VGxC8t4xcoVWw7WMm+NYEnaH8
SgzxjM0NqCpJjPtaLjZwdJKb4Iq8/gxb34nGd6v8LzqiIEjaEdaZO1fFC9b47E26
xk8P8V4XuEOH1sWOse/qjMeKj04XbSFZBfiDIF3IGmDSNLJkY4TTnP8dw55EeWfu
t3guhH7/p5lALJAQBoKa3Q==
`protect END_PROTECTED
