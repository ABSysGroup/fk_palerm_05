`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TqvNVoZ4XGTj2OTDYVo+hI8hNNcZvUU0W3xbXn3DMH5uYh6Dmjy9oOdsgQ/BDLw+
xgg5ti0b4DMKfkMJJjOUY3a+/cw6Z/jMzZYFQeXteibB/bs7fm4Lmoc0pJQp5lGq
BM0cwQBBUE3gKpWUTAF/onpeWbvtFycX06M1E8RyYlVjxCyzvpaYnIKGLNo8slj9
F/M9NWgm07PBy3/HOAVl8uL1zzuC1l3u2qfYbzUCQ22YztK/1gT2spokfJPzDRzU
FLV9L2JZaAMoq8dZtGVj4NWr1JC6t/yiW6WCP9yG5F7LNlCStS1VeVTf3qDdDVb+
E/jO7tSNJkqNI9emDsnoqhvjiVRz+tT4yuea9B8Bpl+WkcMEJFqQJSM80D/APTRA
eU8aPK1yDtCbfvAnNuE3zEkCWMRjgqE6GV3ao2FxKYQ=
`protect END_PROTECTED
