`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hRFxCReEertGrxNhWUYVZbFn7LT7kxzTki3oJqQKR2fpu45U2yg9TdOZsMW0C/CF
le0A//mu6HcDjYttP0FOqfzOh6Yn2i/070vkfWbHLqQo2kysV59pHHfwdNPDBYfP
ChG6bCfkyWT3g1Y0UZ+teBNd0qiHcmMP93xJvs+uATUHoTyjhUT3BAs5XhFganeD
WSsoDRa5iYP2C6g47b2m7aBxEp8/4pvONhoEUU0ob0fRT9c5rM/ZXfx6moUoO/nG
lGcYLQrkpAqdbx7nd4AlbXQGbEmvP32uVzvFXb1vcqKLbZvnHyhkm/ZcJ9XifZB+
6DYP9MPhMmU9Pir8Nb/AnTxwYzGAdkWU7viTokLo6sRDeiuqYFQEuEiSG0KstANm
EuWnUbnBL64i3+YIz5XAmbffOuvyZvGJb2097Auq3+tfkaDZS8AoKQvZN+nwsQei
QNi+vRK9Et1nkt9g6l/GYl4LQxL68eq9FHVClxI8Dgmj/FUkCVFX38w5agtzadP5
LvmmKcomznMa3gA45XiUJNj8zVC6OsyGwBwn71ShMku6gpQ/wn2eXCOTsprkGnlI
F25TDPmjrdHLtrsUW6Jvl3RWglevf5bqqS2sD37CbVed7dKDgEPhQIdq8dsBsi7H
9AHO/4snPprFi+9IHAHsc94r8CPdArrC/juPhZSaB1oM1N2wd2vTfcOPkks58TXd
/geHcR+RKlFTa1fu34H1zuFjfymIIGZCLl3q7M0nBEpEHb4JEYbTUvtHBBlEGfE6
AgVK1CiX9qE2FaQy1dcZlXVlYfExVFLM8DwUKRvBWRzirpbjRtja1h5QWVS8ddaq
WRu1dYYcHdH6hJJ2Rf3bQs1+kyeRQJQXzFUWBigHh8lgvoJZRsVdHVx49R/zy8+k
FJep5KtZPemH4oE/xMsF5g==
`protect END_PROTECTED
