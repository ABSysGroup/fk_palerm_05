`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MR5esDNhKwgCaYUjMe+9tj4iySFPNkzbEHs2v5lm8MOdzkDrBAOtas+tiyo27Cf2
/8avlfNi38B9/bPjCqDAgVFCaGpm1v7T0Yik118co/E2j5lZITVuhCwFmShciXLz
bY4FKTaycIxsxFWETc7+IGL83xaTgF1LAjpN78MSdNx2hxPNenbh4EI8nshK9n1f
aLg6yiiYSmCdnJgidpClkdIRMuYYqLQYk4oA+VbtPUgBvn8RY0IxQ1LMB2dBjz+7
ff/HHwZJ2v0rJREM9RXoFuNAvuuUzYwkkBByBGSezXSCtNeXy1xdATgD3viZn+hg
ujMKT8hNm3wW5zTfgq1poPtnqbXuTUrEWQzYLLvXCt8nJnp4shVK4kgNqmZlgyMZ
tLl/wpvJL5VPoYWXeFTtnx6c28/3K0L1TKUnSDNxQpA=
`protect END_PROTECTED
