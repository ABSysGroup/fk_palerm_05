`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B9FZveCrDIXEs7IgCdUhWlMq72+6L7hAcXgFlx5onw4trJOfsoOUmkA6fqA7V0RD
2GnEG7qkbkoTJ5sbaG9QPwsGVJKocnV6cWjUDeGuTdJQIpf8vYdrp6MRLzmqa7BF
afQXjGm+6XMp6fZSSin8WxYpGHJhDCyWacV9Z3EimaQnnxUOOCTqvKyK9qJbwVlB
XTGKO6gnk3fuPe/O1Pz9iiqRToEKoVEeWpDVMAlb8XP9N56W9CV+mJHPYqWkzv3n
QsuU25hjuYqxpHjH/f3BHHPNE+dU8acIz4XoDd1ELb5GMz2eygULE5PIk0bmCwr+
9r9ogxxnyb8fco1UsmVpH/hhetejl1h1y+DIxfWtWozivV9VcxVO9OO4wzMd7trb
SsUAvOgT78DtdqaXFLVnB0LmZJ4tm4pslllg76sHAIyr8lalrCnQD6dRqHdQboCH
`protect END_PROTECTED
