`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/10sBZ7SLqJSSacwoPhjU3vOxEu/IWzIbcNx1+QBkVk/Xuaksl4LZOohXFQ0EYVv
WCa98wQmx5okRKLswZ8FIL3mIFp+wuNS1B7ceyDuTqtcNl5TU9oGhaeNVnmIPBBM
XKuetTIpTyfFMf0fyXUx3VT2qIsotfJvSwCP4oskHSCQNNBenl32DmFK49HAPa3e
FZ1wXliERyoHtwNTsuOHmqfCYcH6YaGN0On/5jLcSR1iTWZ9BjOGfqluoEZs9eDG
sE6OnOi/3g4y6LXO1xxzFWXAUoKJkT/fcvtk7ZWIWFM=
`protect END_PROTECTED
