`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fKYxPNWCs6L2KTVXNRrt5XG1X9mOTCwUzBHZ44sAmBQ73HKWYMFGrvS2mKi53/67
FqC81PO7jz//bxh7HkqU/2ZbbDbCUKok8RRB2Wi+yLkLHMTqUgbHhYACv2LInyGW
xR3aE+Qjq437KgmRq+hPQFhhyPAIAVFqTR6ORiWS8iZPR44D7ux5aZajKrnlxNdV
vSCtrTnTclLsiH9ww0CF71YeWLHov5TmeX168fxlLqx3HUxzKLxHrFS4RvGt34fM
qkQp573+plvBrln3/EvYi/2OoIm84HDD1t8j8/NB981Smuiz+NZEyeddS7B3YMSL
pxuFWDvSjU06lt5SuK/tcQKv35TSVlCibk+OK+F09uAHO+/3ZxeBHI+sRhiQTFsL
3X9qvYSyIsTWfoN1TUL2F6O2InFrTd5kLaXE9UGnTE9sRmspFrZow9alf55Ja3Eb
df9vQwdG8n8MvFjLh8Tu6in818MPAHos5TE1k8JBPbhuWyL7kfRRzpXFeW3LUVgm
CDCgrR6Y3Qa7+znviofHogZdJ0CBH8JGJvosDJcTLnbimjyGtx6rfnQ7M/6EQRbv
OkxHa9FCrA9pElfzLaxToiaGsSBgBvc6zFjNwXtFAhey9PUi+MA/Sjbegt7uhizy
qnGwIWOaevb/v8XW5xp7oe3qKve3m4YXyQMQ/KPYxqSgUugghMilvoKqwU8d8JlT
+GJ0Ncg7hC4ay4kYYkVi/2b0/lt1IWrfSO0n73ITGzXpnvw72WKtNLe0EHVGyp5r
9ngcSuEkKzAGxEUSS7K3yEc/dhK/93UDVTbKC/BO6QWxpxmtIwqEqoPPJpUVsoub
FOOrSI+EWhvVRzHaLtpHucJU+G4UK+m75ycLN2uu0MAV5nT7rzWq9Amtyh0yn1mR
Yps4T68KsDqHmZPvRhzApWe5NkjuwM0ED1qTbibY3fGhh6fb1nqrMyErmu4pNW/T
iwYx4xrcoPxPRMmMta5JqdBii7KANhvuF4RmrJGRHEpLzIBuxqmhmuPK5KiBjoe6
B9DFshVvPXOVHjXvBjgy/2hMoZlYiuG/NoOzbADIbC5516+cUokBim4U8c8mXg5c
YOw/vW2JhnqyY4qCuD1NyEP264q0KP4twwxzL4T/F4t76SSrpTF09pZTi9VaHQ1H
GC+48D1U9otF1Nc1XXbPEKEp4DGoo8hQOLLQ3LDksRliwCvlZF0TMjshunoa4kyq
plhoxnkgFKjTH9CRYyG136bdtNA9PDwzsVwfHnPrx/0lbdNoIP02U+mt/USjPIa4
3tSIma9LQ/5aClYcKPgJe0JgoYR67944REzjKwb3EEnkBA7Ird24cuouxkdyMAlJ
/g8yZ1jNvwHX3lP0DgHp/fVbyypaLYBIDByXnrI3ej+lYWh0VRNuBgynU3lX/L2Q
rNIjcyYGJYJT0JiNGtrwUb02bo4NI1G3f0LSpo7fGeXOxFo+o/hSWG9uKx0yafqo
xNq9vmcnXcaXjUF2fEm7u/9Oq/Fnznos8GcqSwcMOggCLxWZqfHAq3g8KjIIzk1w
XMUZpQ82nz4NyAKi1Yk6dlWRX+DH05qvz3MJCEhxmora2YWQHunJLB0MUA9luneo
32KQdRvMHEQrw0ueerQUtINaHwbrm05jwZPpmqJwbqUsDuFJeuouTI0RMY5TjVb0
L1KF/CmRZwgBsd+oZZCWddHegRFTfDoeqqU4+9qLaT9xC48HV5ih1Huk5rWCAgKf
dS0qlSF9daalNZxIvKGScVKiRI5zqPsuVkt6Tt0fCvDwTrPBZWmobMAHYblRwnP0
C86MXtp3tCGo5lY8R9/XvkkgSxuU3fLZIX0hfC/44JPx/Y26epCmDc5DcdKzh09j
`protect END_PROTECTED
