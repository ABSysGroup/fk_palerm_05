`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aOSUolusVV7x/MIHDvTF+bPq2Xd4r0B/LkfLo0+q3LtGZt+UFmCwQ8JEXYo20R1q
alrjLAa5YjrKYL3kWtRZ1N5E5pxwL9pATJhjvRxdTYNmlxDd332EXBPgYU9/qW8Y
h+iV6HLBiuC3L6mKg/7AwMTy0caeE/mnY2C426z2XAs8JGAQAnFX4VDMUDYBDsCh
VLV1rbQNR803T/hLfPQAjpdg1FX7iZihLMMt1q2I7ydD12Jb5dykbCdv4LLKM42J
sh/67dsoz7mE37x/poCyeaP7G4zNuC1xiE4hwNFYCvArmzuhpohRRUEiJXgY/ny5
cDGGDJOqHhv2NJ/Dk5aYaRs4UGXbMTVvs1hODq/5MdMShjJr4leSGph+D50tRlgd
9m4qqjmNUnfxc8lw4Ee0/dYtkOQuhqLXyJzpMEkW8TaqscA3treXjnpFmKSJa0IP
Le9AKoejnLMHtBoPaqGzBrMd2VXiCAEZimeBp43wQ+YVNInU0/EfBNyrw2ekR5JE
zIyDurtyHolv9bebH46s6lZmyrieWGYE47YaLeUhBRtaS7hS93EZYd6sDWzVlRdJ
`protect END_PROTECTED
