`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BpFZ/UmBFWJEMHfPtQRdygUFvdMLOCRC3rukEAM4ysEuBw/G7aofaxZc5SKEsCPe
EV2cvF464kF0dlh3yALZ2JKW8W8pC4Lrcv6dYi1cEpsueKTVlWvfePfzNkpeOytZ
2a/4RBXxKXGzSBdnvu6iXWVolpQIigvntkF9kwakoQj+1amvgGzweoi5nZweI8Su
spiLvY6qwFv4iz41y388CJXULQPFhN9yQmUu42HlT4Xfg4KDbDoJp/BeRyr0zkcX
KTUPBuX6VAvq254XOOAItFc87zErtzdph1Linc2kCD18Xuqd2rJ/R3EPHZZjjoHO
gr8Si7IgqnsVWZMu5ijVcFHD6oAxVOobPs+6G3VoZuUFbreJogQtnUitF7aB5DOW
H2JISCdGEAzi13KHH4krburXkgvLaihwNcJlv+UwJ+SVsWydD+aDQLAdRmFTinwZ
UeuqKSF71a6KDwexOERmp+6yNJqusvD9xQJpSlV7NvXnuXRm8g5PP4NRRJIcs7Vk
mbESfIlieYh5FT4iFjwfdJT6+LC0ZDYYovdUFzClBRAdijpylwaU+IK4Has09cXx
PftbJI2XCR/Xyzk+bE25Fg==
`protect END_PROTECTED
