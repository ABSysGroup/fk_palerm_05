`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
srjuUdK9gxzYnOjzULPUks86dzOLDUXtBSSVeXcVo/Cv4jPyt13N3bomOqYxrrkd
u2esB5uGf7Tlr5TLrS/IQFjOurQdO7yMb6/6pEyn7NK205H2xnkdcT1REBYc8nuG
h3Z5P5sP61yT5woPlJ8G2RaNpawxPcv8hVi46pwu1JAGV1YKkOEuYyYCbH5ZaCQa
+Vo3WNVjpU6IxwsmZwlYlg==
`protect END_PROTECTED
