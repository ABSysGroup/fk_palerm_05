`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7cxZXFOpe8DJhss32JlekH/pbdZmjRTn50a6VcGvak+d6hXC2RC1PSiDULKLaRT/
p4a4YflQK/6YuMe9YW5QHvoq4gfnjX5VHpQJ6dNo/WvfqBI7GCqrkOeXNyv5ftnd
HsX9iYR+C58phHg/coTWKfKJfvs7mmlEeLrqVkzPK8LhzfwobzPUVkMaOW1p5hVn
/rZ+Xs/2OV0tmBuRlYNKG55QODYvgGFCl/fjfMG0tXdhrT/gTe+JPPFQFjxdqw7o
iKbezaQfLtmiT2CO5pplxBlP660ehjIdMifV8FMGKAijrwwQWGL/IwUS7ZizGbKV
sEIS228Ibm7Ty27jwqtidvRbk3LEIVruwCIshlVt7/SdflttgiIkT+he4VLoSrQd
OWdIeUJmOTmmg0hKh09WkiV6UdS3Es/BRTAW51SZLEc7uzm3SpMB3bYzUYrVzxr6
ZM7gzIUIr6YlLZNypztSFK/jtZ/VNXg1RXjMyEvKZHs47dDM5fHX29iz3pkhebn8
Y6Z7sNrCNqR7uPsQiX2ebLnW+gck1q3Xw0Fp/GpTMu/2saYGFC/3axuaGvSj6NZ7
gamHMGYHQAjcEzz7+oeI0t/66pz4kcLb+78bfq8bon1TS7xNVTKWsDvyinM9JVQt
msObH0O2Xn7tO44249lTL48Rbi27d6G0wsFGuu1YU1gw6l1yLg3jWCt3EhpaWNFt
eVNiotIG/MZAGFF5CC4pPaTzR0Q7TblG7HxtSU0WR15d25veOuixwaXz9XUgocEp
VWbsuLZYZvSJCMmDytHP693HmLzJnXZR9Bxgc0+fsaHEWAYs7awYmvM/uZWKxVOG
JFIzEI6+hvKzvoD+/MwIdP3PR8SN3+gmwDe6BxN0XFls0tJfOyWt0nOPrmqToxsc
Ssf20pLwfQ3CMmEdqCu4QEoRQIvST54UNTmHN02+6EAERs4rNOzQfGtbwrLUi+lh
`protect END_PROTECTED
