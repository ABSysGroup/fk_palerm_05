`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hcPHqI0gcUY+Tg3lvSILD3EQYH7PYherP1ljdBFmHwf60G0Rdy/xxfHjQZYHakLI
h17Z7PTC9n4mnIy4pwtQfOX3pacL62gXG3mhikddAgXa5WL1FU75skilw+8ehrcz
r7YxWTgaAgL1urBwoAzLCnHm+1t6OE2W2RgmU7DA8T3ukpbEZsgZ6efj2YCvF6Nq
Dt33UwXTSuQ6sIjUgsx0V3GZb453EbBJAvSSqlXA9KkuTRSW5q9K2TJH0VNlSFn0
O6IviC14VJ5mL3InJGe5mEuz+6avZNb5yTAZXu7IQpwAasaFNN+VkhTatF3vG3TG
9eI1zO5tKNlgxVZlFF7EGm5Ne5ZSUNpnVHBUhLLh68c9SrmqrKtEZnBnpcIs26Di
nT9ZoDV9ZhWyW23Nk6U26a4Rw9KDl4QaTbCK2wOtWheY4DccymK2DbPKUwPYKOxV
`protect END_PROTECTED
