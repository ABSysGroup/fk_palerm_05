`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cP24zzSpx0v8oVP+hcWzlzWAEcUWdeBKfJ/2+HT50mCRZsuEZFMdDpoaAbWfq8Bk
rOTCkvcjB+w9DNSCKbBoNY6Ax0iwllrwBdovFtaE7mry1IJ//P7kpg16T7xbbKSx
YQOPB/PWVsFZChdyFydvlsYOtlgkEkbuAimIH4Q5nISCAV5yxOqeH1jzSp1LJVaB
noKSBG2U2/zW4ETvGuMRbgQIJbOVtcGYuPmO89d5wre/PyX5q79sEEihJF4tpoNU
UfYqNULy8KUfl+Gp8Qi/8FcUiSGEPLx/mPk1kB4CDhS2BGmzj4kFyj2nr8edP6e+
fqEKXwto+px6hr1n09wESMj1+6LwNjNt8tF9WK5wBQn3yW6NllKIzCnQV065YiXx
3JIqdR+c0z6RgnocAsOBtiZcHUkyif2F9oBhVrrN525I1oKfgvS65xZFMPF9oVQZ
w0OAbnWeVjqQT9aCqH+VzrotRM5Y0yBYMou8l3m1KLIoaORZTsWoY7BDsw9EskIS
gik5q7Q4EQoCJD04/1QKGsCkC1mneRb38JVipTP0GUPjiMno0GjetB4ed4UtokIn
rwTbdA0B+6uD/4dRSm3e6mJfiqWp3KOSF4AKCBrZ+PpOCLXQUkgWIaSvM02DmBGu
thB/MqtOukwhb7+hTH7ETmEsqJYaCZ3fRgYUmXFZjVY=
`protect END_PROTECTED
