`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1waujnr00enEXN14u/5qU9wedjyyQ0WIb8+vAtWR1haWXSdb2iW5LfcGJTg2mAZR
eZbXMhLSMXU8ujXahprk0OYzLhSE+jk/tJrqfPyN7rLqUCvBY07cAR7unEEpBqDG
LhwAnRYgiNrd0yRtvustyIEbRbBxaypqBswcFnVSq82aBGwinYqIEOGEDLDYbZfs
XvYHboDwCuBS8bk/cxzb2ndQw18fHwU0YadQbtLDZt78+sOjBrSgQSRYEw2M/Hb7
v1t4W7l/DdKPA6gcOcPaIaGB+RebTS0naft74NquJ34=
`protect END_PROTECTED
