`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9VK4Ms8LAe1Vz3fGQD/sRgZ/SOhzyfkq6vI9qj0WQaFkVeq3vB3g5QJsG92mIDo
c2ZkZrNnqtWz84caJlktMCsECsLZJbxj7PRv0X0UOsvY/o1myaXrYtIsHOC8JBBM
N+a+ktlEwTfj272nBTVaXSbW9ncqPvG25nSGJS9yv/2kbzfwEcvPM0/Cs22KvHBO
FLUxwjTbbxH328ZUEAONlzAkrOY1GdPCdN2FWgEFtY/LJXDOtGVXN0dSM1VPj9Kn
ryJ9tAcprtE5N4Rnob3SPXYNq2HNF/bEzWu9nu777sknwto+Ec9pC1S3tcbjJwSf
vHa/PDBowMU+P/n54PtXon8+odMB0XPD1TRL4hGx7maKZH2IIp/3YMDIQS53gKoj
XrXAwxT6/mxTfaPFIhg4hYBVFUSqRqpDN0Pbsh7dXONlG4qjOBFRBdR5XHP/qvHb
hk5GyZcHe5o5DRSzcmSH6VClp90c2Kwklgde3f/bNqDb/Vqt937TqSw3MW0dmTsb
mCU5zYNvUUVaCz+YK17QrhvNVXtYDbx0UBBzso8h+/l8PQHz7W8tQBfDexCZxgQN
GkiVaBd7bRIDYNchhU2NLGfisiwIkmo8L5U0Y/ZRChXc/u9SLDqopy/WrXm57yQL
dfbFNvnvACo/CjiHtjX12AkSn6c2dIpnbsY1iYcFO+MVEp6GnGGQPjD65JNEJ4E6
HJBFNNdS4ltvg0Nof+IdvzB4ZG5vU1KYnExetapT1KV0GGnK2U3vfiDv9x+3t1qL
xIo2ZKOwQRVj5gxN59yCQRgL/wOFD3ImCB7E/h5babPwFvkep6lGmlZqfZ+SQzv1
W2GpvMJcyzHMMpzUbnITQl/aWPl26X7pJZWkMeOq5Ue9NdTY6EZDvj290VhkCYHr
jm8s8oKK2wibdylPdEIn8EUriVA1dzm/DWU69yBNvxc=
`protect END_PROTECTED
