`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xg1kRVSVlCxx59Xv+5gEb/vQm6JJkerTZtSOKWrWA5LvLzWRTuCotH43tqdcZisb
QXfrj15JbEweCtjZcSri2yA38NlUYlVVpVo/+zruSzznB2rBrJQTR1F3sTEkhnFK
0aCEc2zZxFqigzKlo20PeRDFsYkyjv22kBzdEm5xYy1+W/0mEIn08yUCnDTOliGk
ciwSb8VwlMXC4ojOuaHno/OKrxRGK6LAxclY4+JIoi7FGXMYh9XoCHhk419CBPUN
ZJ2YpJRsfZQh/xLEwTKYzFXib+ywpHvFKzSaE0zevCW4clSIF+2jF141pMhtQdMG
3Fa8+4lJNoBpw2rLgxaVXIsXlz/E24zKMVe0w8kz6wm2ok0tfCRHp9O7Mk1sDK0P
oFYpTQAW/zth/DG79hBJw9zQpSs3no0FXvGJslRWVCZJTyadZ/WOy2fxqfly9dPo
8M0pulJvkzMOia7pViDRqZkLkBopdtTfKYRP0YituEn1qgiST86vrNi9QVZJeBB7
0nBJpyo7zWO78yCnnv4wq7knv/el5AiJWHwson/4g+h0ECY1r+WcAs/dYh3Kw4BP
WrMMP1TZGRhWS3FaAHdpGvhhGTknU7CLtShTSnaO9DxL8zVDpIp0vShxbs53b4kO
xylYIe3zswHCNoSxEgJAdQ==
`protect END_PROTECTED
