`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M9QJxUxmNDd3lyeLHdRzydPrT56oob7VK7aJMdigATlMA+7bYqaDIrmhKPS+4RPT
4LXa5q8Iap5H+8o4O74uZqbOSkScHpojIHhOozxHufNoDZ+2pjRXif6SkdNlaz2n
7LbK6NqVntQNLEFT1vd9L53xK7w4sXyAPRv2+8IeLsMn5rGeMpo08kSDMOyifFc1
0hJg7fjSUVuzRUmIPACv6vUhyiIT/QS4ChcThdKIhNUhOueRVeOM2hzqoAZJHHN7
QV0KJtg/utwDDZKoElgRzI8sxtX9wtxIMCyhGLoiOpMfC9aRNlruf/S7D0RGxv98
eDsziIFoMrE6CKzB9kZ94LoKkO1uZQGdc/8gikfGpA350eRp5tv+AUrgzOfeCaml
PPobC0uxlmK489F55cRBpP3Q9c90Bzoo1uek2XV9T0k=
`protect END_PROTECTED
