`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1UCTe/aJ0FWS/dt9fDGQi1IlwTXzP7oOBqevopmncSevn9FFH+XOEQcs6iCjStrp
QyqVzlr5+0VKMilwZENcyFj8TVSWfxvw6k+vBD0rEWfxeoM9LdAVwzsi/4MYXKEr
5wEKdIxAcTS1SXJcSIBByqqyUOZAuK4iL8FAj77xvNlj+X1oiHEtVph9U6puFZON
c3aXnmuzdAqJ/0p6SRRf2F8hTmZQOSF2MuL8bne+ashuVyjgk4/Cypn19vxcbsRE
HRCUncihP38O/shkSpVI2vVPxQmXrW4t6EZPYIH762Ee2TleIofbDMMVpp3HqKEZ
CnKZMM8Do5cwML94cZpeKAiHZVZyBYyyieka6YEAUrMKZf2p7AdMsjMqBHTPidSp
ux/plHYj6Lix9sC4Jamc+jsZBscB37DdnY7YmfDofAwSeVaQqLzYOI3d01IKUvNw
J4RrwceBQUAT0Ni1SSzszZjF4VsxeO9BEOF60ufdhox4oBizVbAaqF4fGjTETpcN
`protect END_PROTECTED
