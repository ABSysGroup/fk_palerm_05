`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vOHHIUJ4yq0Xg2nzUfmMHNUxI8T0oVEUm0CZCgyV2wvzHVWb2fSpt6ef9ybmPf3R
Mv7VXDak9SwAefobeLADMVFqjNfaFrqrdctlAwMioeabthjxPTLnnxGpCT1lU7A2
SjmQGECuC6eeROBMqXKiRxe13YRaELx6d6tl0R+mgOE9fpzgOawfeIA0gKj3oXN2
1jiHqU/Kh4HCQOOool1gmZPrQNjAzZCG7Si/PSIKAvlSqhG/RepKv2+Wce1GquwN
6t3n0/frGJutKB3AsoWSJB218UFpm5BH3qSyRfmlzI9pc4CtKBVjJOK78aZlhrKw
V9sa7TOt3eNo6NaxxdRLO3DiwvRu0Zj+sCE67DrPC/sCccct/Bu6JD/m4u+PQKmD
HZvl0vIuSIS9q4KCI8mUqHMt8SHuZKNxzwEiT3/izhfEfWngqwGd0SBFlpqKgEOl
f4pA7r0hCGXC3Srb1jwZtPFGdyX8bmCzJQT7mhlOHazVy4+qwUFKrc+qKhzyR1If
F18EznOu8bCIQz2f5dH+x2xREHTWq9TW5PRAqDOv+SuwbKn5EVdpLA6jws1un56W
WT+2IHbDzrq0G94TJ+iACui9cL8ALjhtFZjQbYU6g1gCUyHrs1PsxEuzbWaopwCV
BzCrnj1rTb3XCJT9UC/kQuPu28qbxhjF2tBoWQoek12i0UHeq9W9C7pOwd1YA427
Xtz0sMmr2kV7Ct2O6PD78nruco+wKOG4bL+MsH5bv+A76sNVoQApkQ57qksxhy8o
D8szXhbxgVUPXVn31cOYVwwxW5ZnMSEuK/013Rz2/cjckE6VkU65Fz/CAOwLWHzS
T0CfXS3DgXOKw/tIDQ0lA5Zy0vpaBadN6nYEK/tcOXz5ifv3DmG7z84OI/9ATWLT
nUB3eaXh8Wd3UApMxshJRD1pYIMMsQpNAcF4zA50GHI=
`protect END_PROTECTED
