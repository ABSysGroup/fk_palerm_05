`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E+9n6mnpwhcVdiTgt7WNFkJXfwwy8xDQ9qzjxHYXYP09OeMSaDBoEXrKLA6gLf1V
wjC2ZU3zrrfAXBaB311jQjB+cCu5X3hvD0r6ZCZsOrQu7XZtSaZ9iHgYYwNDtcbT
DP6FJUiuD2GJ2us8Kf3l3FrTOeIE42Vqpd1XlwcRxJYZXVyfJZGdtvDcn00wYOij
5AfRCX5y2sKGyfuvjGnTukdJW14WCwPCiPI+X3QD8W7OWWjGOiOyWD8oeol6dnn4
9kAvDKwkEURmqSfWgtY1xBvRgfTzsH3vvxI07Hm5eyzwlhzsbaj/SdM8tnIokUl/
idCv/DJTvPGCUpVmxL+DcHJGZRyZOz+pxP4z/Pa3mNNZmqdTTFNhApHYgpoSMZKw
n0yDdSNvdWYbOH1SV+GohDDza7KdyMs7qzJU5ZZotmDkOCzPnJQMiJzeFAmGgEgk
GMtE6va1hBtXRiEdfC9Vzw==
`protect END_PROTECTED
