`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JqTsu7eTRFIQ0O3NnDFRsSzh0d4cwcvkq+lc3OJYvkLDD+435/9r/3KT+Ip8hLP2
Djp7DLvT4CDrd2oIelTSYAbDW5v0bdDJdLw4ZjGf63+yDgnxDIv/qUNhY/58Wrf2
zuGMmkNwCM281k/jhI7p3GnteSby534kqr5IgDcQn13/Zpr6zdh/se9bdEI8BYEq
juzZcdZikVSHsMyGECBMJXlcI9tvCGWV+TsyJcNvt6NNLIEIQR5csFeRIacNRnOX
N518mesR8dDc6vOTKeyLIO+ihAJwi5gLnmt8GIgsL2SF1QG1zCjL+ceJ8R2TYVVk
lmAHXhPVhQTTDXfKM0GK65XR3sDu2EW3GVbFHUSJkOLnwghaCFn+bIAoJx4gMjHy
Psbyae/m5WjdAL0hhVyMV+GC0cqEGh6m55hM4XakDn+0isf9UtImwl4WFk5EcDgs
gnlSCY6vkaAP3U/X3vjouQX4qw6I5brKXOB2j1ydO2zpHwRLPm0pa0JJiKlKLanZ
zxfA8602nxQgNvSiy79tAlxsCs8D+hMWH/SzAJt1nOWki9SyLJsoCoh3qynP1BB2
o/Nxy/7xYefAr10g2YSJI/EiFOZKxqXk/3Gc7j04v1wAks2xf2xDQsol+bqQ56yk
V8d2L42a4AxP+QeKRYimlZrxQa3153x7ZOFJIumbKMIO4WQm3mNTLn7KN6m2SEmX
yPX/Eza2f52r1O3Cs0S4kesBhGQCHylyY184N9s3YOSU3WZw+a12bdtViey4Ok+n
ZxjrLB1gkjpZJ/Bf72+cJnjO4kP0BK0Wi/XTsQFZD9PZL7R80dRFDcQBQfcutwiW
1TvDFGEugKexabt/8P+EI97HUn+lDD/tJbbcaaySwb44ScKlRJXxhLRdx1bUNoVE
h4/Juq7qgnRWjdZUfNDx3VvgUdanZ0c8rJWpY0o8gbrrZ2uV1UY5oweygfirvwZC
wrrAn/o7Sv2RKgOzSN4wW4I0WsopUbQOB4w+HkRJyElzmA00teUHMlqVqugsEi+o
FcThqHh/G9K1ctyyx5KLp0+TWu4F14huT5QYwdXcrbZQDG9b5NwjJDdTemhXsA9Z
1fdLHeqxdWvuO7T1UTXKS14VKkG8e4i/jUzyYfkvIo3CL9QXJNEDYNaB/Pxk1IiE
sMKXJXJ1OVzO7hyjsGRNhXCxW+d99KlHWnbEMC7WytZv0chJ58fCnbb/lTDoYCpC
jf4If513tQFqwh9xhXttQUB/wa3tD8szTJ4Nt+3fs8n74rqrdb2vpsz8IiOHzfva
bnTTsAXC0YM0sc3YTFAFbu+ycrOMl0lmACGBoP5lYiiMsG19UwQHUT/MllglAsA2
02r2CKmePGELrB0558IVdcLTp6uWFgqCiFWPW5xHxx5vvAadCPOasMRU78b0Lg7P
WKpsxaXKich976tDhtUtq4Yz/08jDDfAJtMUCOKBF3AJiqyZHj7KzmIomkC/gXv9
9cYAVGFdZ6Q/5IjeizjHi4oXKRUv1wqDUwfPdpCPB0pRdyC6bCpgC89ymOJyDzdK
2e6lKckDUMkKfK5P91+0z6zsprNaY9EhHR4I4EvvT7THsb0qPy1chm3E1PvdgMbJ
0yq38tUwBL2XFr5x/7Upx/yB2QBKWUN+vHfxz8zo3z1Zx0cmn+LW2dpHSn1sfdsH
XlpRkfKGbqfrcsWCCT9DFPSg+NSTlg8Fg3KLXS8ts47o2fKyGQIxqjIB8Tc4bMkW
zsMRdWb9+eyzgJgMNxbPZQv14+XLWX75ifMWxfq+6YP95edc2NJKHMASV6u7rIow
LGSbk3/rKyNQizzaKmvs02+xgj9lQnVKlvC9tdUcAZR8qKVxuxEGE4YYPOd+fA0j
UDChhyNlbKP97ZE/5sCsM6BXVqo7YAxoLHVo1SbEz3vH5GRLvedgNXPNciokKZI5
KeH5dRQtPu5uL/z8bJ+VYQEi5/u7kq2OqeAaPUvZuA7G4AUr3g/Z+PZd5d+TmD8r
kq/3vg46xAAq1z3cJEeSyv0xTg5ED6YaAJDx0NDYds9mo9rzl5WDLRCqOPawL4ZL
DhirSZP9IMhWaNeXYVqr1lv+LzX068xMIOyN+3v6Wbsyz5DflGCX4XBaALbjxv1N
UkXhbg4ENAyCsgh7Y1ig/kRr4lnvgRXjCTPHVTroDVXOVxddgqFh8/9T1vWSU0T7
iccgc+yfmEvi9GnGtFepDTx/CEpcs4pBy7EZJZ3KtBmn/UxiJnwxhXV43i8KnHLe
Q8J+KzCMwQ3P0FEtkZyxDSFBTZs7/kA8mDB4e8ht6iGSTn4+4qxUoh+bZPCVumFf
qUM2rnZjSKo359GyGsJcIujoNAe9EvLHOJj89ifk7AegT226mTLvPGrx39n7xysW
h1HWqWhzVUv1l2cUItIXc6LjNyU85Gq+1jOr4baurVRXYPEGzsG4iC4mMdsfCTdi
z0A+DMq5Fn4xIzxzemePMPgNs70bswGCbBZsoCpQ82YZaVndUaCgMI4Yh1YdmhZ1
BEKkvk5YFrugw3DdV5EwwyV1E5DymdIX+BQPTd1p0JcUwdSKOw7H7BX3mu7AjhSi
hAxyWXiUg+M44YrxO6mmbFCBUMb+dh2ht7xxck6VETMNWtqEeowiiZ6hibjNZXc3
/E4ZYQJcdEhdT72A0HJB7EF7YyHugcvvKetAHoSEuG89ybp3/uS8rbqwyS6KHP5h
Fg6ZhyJpzpKjq8Q7leLCgVexSh0B4Xr4Pu3tCUAJkQ1DkULO3MO2egBQpBYM3tLj
t0/zn2iSvL6+j+vzyFB9hJnS8NX8T50BvwfXHbMTJ/p/ifF7xwLSREymh96M3efA
+vNpOBlwG7Tv78wknrAAA6emWn1u9Km33I7T5WUSo95/8KfMGwPcOB3ZCnqtMSyS
qAwK3AFU4rtNS06pE8IqO4j1lhKnN/VRfwtf7/bMjWCkj/Y5vPm6gfuwaB/KOy8C
2XfUNaqeoov4bOLqf8AJqp6C/BqKFu+jyvPf49KGOBvMJKneYlbLdiCz59FjQpnF
FLkq0LaYx+BnHjmUSbEsuUtZ/Toi6z+Uy6Jhi1V2fZFF8bC2vOGr9X2R5hSeFFsd
rKfDHnAvjKRr7LQjD3+K89ug1/q/2ap5dzr+DLbgQ9fb3HES+KMuMshl40+w3KRH
u9SO3whsvEhDkRxj1otclj9oChXO5VrsMrt+wmn7sLvjAEur6yRDTsFyOfrYPqOq
MNHagMqEGxDK/mOM+xd515/+R53dP9ZleiGkbpl6ZpTL5BFdydtUntRelOHKtJAr
+X27Mbp2X7uvtjWQPzeQfef161TAN1s8K7cWTAPI5a/e6RMCnkxmqewX38cXrzyK
aA8kFlZj/HMOEsdDzeMJRxLyEI32TtXRpBW5Kztg9eyPmLs90MLUGWNrUaH07hc3
EK2d9HaLyeENeV7sYlZ3xz3Teo7dnl2+KMmcFIPAf9E+VAIYpiSz4sOhGswSBf22
u5mEiloL0Jf/tOa27RQ1LufAmVCacPLFT+jvD40IgQDCs0V74warPYJUDxpd0Ldj
xGwce7zrbp2QdLp6+5b27IIPGR0unzC4H9OoCHmWWuXBZqegNBlrO0FYMOzP186i
QczpBfrNFMGnrCaKtH8UcLvW5IbbDIMnntQT3hhcdtfulIONphKi/i7kIDB17MWh
tiJAVxktXcUOjwNeNaYeVyniERX2ku18fheeLHBJZLMKr+YKJnqim9LiSRczJWbd
ScWkTkIbfMUUgNCH7lDEMckQK7meIVQ5EinbunlSHnZdKtuPkwvZGikllQJcrYvq
WxaN07Y3d9djr9P5cEIlb43ZOfp+3hrAewf20uv7e51UdsVPzSbuPnw/ayQ1oWZi
2wBSX/+3sB8FBITpkRuK7arKalq4ogyDdFWYyxaJ9P3T00Um+YpY7gw4AuBbCoRi
ww485bds4XSUVTPmQcMlEfrZS1/iEkf6B1rsPNi/TCPjk0+Yh1Zosj6BTg09ZMrQ
pKwF1efN3HHlM371hXrtQMiyb8zsINvnxLW0CYTsP+O3nBkOgf2FTBHPOyhJGlU8
Y0clSWzVnX44mp0q0paiMVLI0SSSrGXduHhtcDC3dAi5H8GDbECDo/v0Cno5QUOy
HhcVbxKtSM5unW3RpKgBTQMSueW3p3YGsoFYqrrUertw4/lVq8jHzkxMPqmrScRF
iuQKTebGMiYkVGu9+4x6Ks/CmGozYXmDLBbukVy25gBszkOa9IhqROit/Sb1y03I
DU2KMjAbnCRqQ9qWFdM53fYN706RRSWezYMMMAtIIrmvoe4lhhG2gbaLzCzNDrMd
V2XvLy9DgwJQ65+TjCBEe/fn1QZL3ECh/nsBVUWTotccMcsjY40g64/A+8dWaYBg
+oUkBKCAy3YzBbPyNUGPHZV6e/FGDjDqo7g2K/sLJZZA3BKVLAx5Ao9HJZolzfL+
za5bMxj4dljQf1geZSDaxnjsGoCCwstr1IP3zOW0zQ2k/r5p/WODaiF9oFR7U9EA
nnmflOSueSdniJSR2aAdtGPLVAEvFzJsT5nbLKhX8YVYX+z0cOjqP0wNfmoyQIBK
OgJ285PkY8Vz2TY4yaJWe0l3LIM4DqzY9/lWjksaCR2AaVkhqMEJtugpMGkZUIHv
9golF/wxDpPJHXKkU/YMvhttCf0ziSua8JuJO1VWsAXykhYVhIL76ss4WHUfYWCk
dJgXIAN973gnjYZt8y1j1suWeDS0/+83ACfGCLqVNtRNDnR/KcqIIy3EQX8CeUMt
vxJ2NBFZIUWQjPenq3xNRSFzLqiPB2Iv77VlsdH0S9nu4QatViHYVjGKtMrIGhP4
zbuf/Hm/w8RK5gQXVK0xfBPeKG4p9rhpDNHqplqq0BGf2+3CJOE7W6YdqBBrSeM1
jy8Jrca6A0G6TMz53+TGdQil3jmdKUBeS80jrAVamDqaT2XVnGHAWqBe9ZKRJJtq
1oHlkRAiFkEjFs/Hf36eyafo7rsYDIf3VWFLnunljYX5hKg84L61cgFfr+An8wEL
Tck46Rl7kxJtzoqHzqsF/MphGe82yXaDxNzplc3hmZq9ESjj7c7XVWik+2NzzYoa
xS5WF5mKnS2ttb78B2eCl8H2AzhDwrsHOrxuyB6SPrdcu6hTzTNyOHjT1G6yjC1s
5qFMAaMlt3duREbOdESIxM3/RO0eXNHRifrAOHEclj+CCQ38vWqZ509OCUJAqebI
1FTeZmCtPMiKMDyAr1l53PudlCr2Y3KcZa3MDMRB1NRqayKZzAUO4miXzMcaxFB+
xafgvRZXmuKgv+TShHBptpmlgDp8+rfJN1o3wiSphmo69UnZ1Rc7Uu7EkuuMu/gC
Q7ZeLK548RuXfJNkxd1WyVilYuntM43TdtQQVIUkgQ4dI/ugOUEGZNPinfrlY802
lZZNcgc+ICX3tooves910Vgv0V4wgZ/HQzi0Txw7Bj+qNQEkzS8hPW/kJiIjbg7s
WjpZoHEelcGsjq2zmq7LajUP12ASKpSiqhTDLqIcCuL+DP24Z8O4Fs0/opbGYASu
dy8us1LUNSZdDTD+aWOjD0HKIktM9acS3ctMv0WNrt5Mw8bA8ckc9A+zCQ8lpxWj
HippcoikHu7qes1gtNHr6+15XrnjxNNax1dEBB2UTzsjADWMcyZxSr1pzXpqaBo+
vCYPKvgjtTfFBB7jh4/KozFcWUo2Ky4IwCcAq+QqiAmoX57MKeOgOOnLalQBCPHb
F7PIykK6GCrdyuo4Wlwl9Pq3V7m0isE1/1iwis4KGp0u6g5Ni4DOrJV48/lWvqeO
uVDtPtT+6kfYxLbWbyPZOWBKNyZAzqCz/C5mAShtHnWEgfeuCKxJkblqmyPT4nqh
2RH4uLeU6cYKT2euiLWd7ODrRbh90lCcXOZpqPq1GqBCsEE78BKizxevDX5FMY20
WrSwcckC1OBbXOOokLkFlILhwtumbwTUe6GkprUmEoTeYRmtggb0m8v5DeUuJeCr
nWi63HCRM6Bld+RyxxPg4Uk5V1r4kYh+nL3MHIn0AaLPGzc5wPxQGcPmS2DrYAfo
6u9+PKPaqMaOovsF1n7znwskamnxkiSBb0RAarScRWaoOUPhbIaGD4HLJ4SBwJf5
sFaZluoYLFjRLOF8nZ41mNWeTvvZTv+ieOLkedmlFR7nn8Xh9KJSPXgqZRxUsnhj
PcqO6mhsLYd0pJxDlo6xjXPG7Y919/BupHqBvUllZV9lYeJPnPVK3FNc1K6dLu/R
ZD8I4sgy45ZlYySHq1NN6BHfqtL0IOC2bTxDvubhlUzFC0A6AlZ/+3W3t1jG72QT
UEJ+gedy4w2wvq5wQwYgNz6qgUzPbLoXmP/Pz2Vx7MyB1k8ty9ArhGCsOpFBn784
Yi+y9z5/Rpkac1AOHQHUPwPRbqXpyga4/29mpTxIGaBh2SOHg5SrCng4DWiloC/r
hQpz7iP0Pl5Re5ZH+bb8ub5w1gHuLGr52IYENuxwYzDUqZ2gouYfqIHDY09nYV4C
btF+eqOHoDyWBxonoN4lX6mSm2F/9pnZ/bGvy4un6AlhSiSTCQj2DSPAWcUFTCc4
6CZGSTmLlJXN2sDAyaAZDgRk6Y1zQYoaf29uIVqsRmuBCQeyXTsJKAenLA4ajLv0
FLhqxVU1kKYnJ+j1khOScJbc6SvD1317EssELb5x1hjSboAxRGmnoXJW4brhBHhf
TL1YR4iKKWPIH4IqcbVh/eoDtx6GVSn0N+OdvZ33Zfs7cXxRL12c6Yo/iZ/g3JBG
Uje45f+POqGWgyt2V8SMiDQyn5RUimKXT6g99FVFOf409OxECCkx26wCybrepVrb
7YUkDYj1SPSDjwrLeEjd+VK2zDnQYP1avv47HWXJufSa2o3HiHeOV265ug0qMg3O
BpxGXmRfyI2IqY1ie3WFyZOah9ye3GHSy0KAuEnICAVf0ZCCHI/k8v7rkudlRNwh
qPe8D/PyRfZCLmCUxPZWmFExCAF/RJE5oSi97D9Ey2T5G9qxK9CgL6r6/5+humtN
OLmQlzh54LF2c39RIqTJ8k/WBYlE4xQuVfiXb2gsU12LvALC6neXBPTuujRDvley
2WkoehabwataTXAFPQW9aPOcy0ca6E5m45ZFoIhBEo3lkNxI79Ebd8LN6yQmXyx1
+KeqSjCbxlIxYcU+lOGTAa25HCxgatjAwNr1r9Kl+GMw3+RpalILe8JzRctW1MI6
eZ52Ch5PbRdvj0zON8MQQDBi+ZPY2j+vcn0oe6VlLPsJg7pHltW3PjRG1ltwzeVW
6VX+oqZAJgCXJNz3EmAwlFetI5NZ8IE8tpw5WveDFG42rSRQvOVtoalNeD9IbRKQ
Tt/EfQOa8YzgLJ8aoOzBNLUvyzIdZVCExoJC33QfjEpZUYjk7iWjFvKJIVyrsu+u
ibC2Mi/yPUAgzeal/qWfPI3aZKATpdZvORpkmVyioJQtFkaFGlfzd8F2GuB+OtbA
cGn/2ENIAtu7RdGj3o9CTmUhMtbcgvvN9+HlSh0lT5kviwRI0QsDZOYbwHP2Qajz
xLaE3Ge5B/ZW56rTs2dCxGOOlomlI4pdtKi0XlTgbqXwMWclvfJMIrKXvWNSB+cg
vUtZHge/gJLo38JDSeUrvFUhy/csecYFBOSY342Dti/7dKq6omDKzw7KlKIsvtpU
l9v2VUxTTkd6VjFctx6riNjgSwlriVXj9/R1QcKA0mR/e+szUQSKDtTrVq2Fd+Jr
le30ADx2ulta8HETwejsFVJ7BjBduqmBeqGlIur2d9FMXtTmN1afRYaCC5lmyDx5
MmZPtqARST1SXIXu1Q4WX8dFZKe4PTVwIVWMIK0Pd0XxQmT8znQHQbSvnmzYOakL
RzTfxtmrgTgFVI0jw2gnAvM3jnx7wP7gTIZ5anPvJYY1tYYRU0jUiGdOGlEt+bjr
pD0nJj0G2UmZep9TUM40h/M6aZ/XRtWJwGVWP/Gv6DfekjZJY3ORD6W/V4Fpx+cx
zbFXi7RHVhXf7xgUS0VgvWGDSzaFjfgBeq3BjvpCQBuZLIMP71d4ZRd7aWvzRFq1
N+pmtOx3VikI0R1kBMWDyYPnx46Vhu0BVVHM+OQtYW4bF+ujt83ruJa8gIIt8jUD
nIEbDEwr0UDlTyfZ7d6u77iVeDnbX+nUaRWTB1BwO1CQcbD8Gb8b2EXVF8ZdJZe4
DJaKHQ3Llbjiw5Qxddn2rU0i2ZLJcSYX9qDgMc4TA3TxVuSxPfJoUETeo+nQGldT
n+1D7WHQzdkvumDvfmMBlhYHJiZYdauTjiWiJmyEL0Clf23jrrVHIbenkXsGZ1SU
0KqujbkOqbRpWAYHtOz+lbuN66GeGaxf8z6UvbhOlz71ofvNxhUumPry5Q9Qp5FU
IxGX20oANTdEorDAcDtwLpPZ2yw/Ab20zBiL9VwcuzLfxMYlddTE1zGQeOY8KDWB
xGbpK64MJuQZ+CzbuS+d1ZvwhnIlVySYPD+l7iG0EVIAK3QHOmz2j8zaaUyzs2Qv
eL5w+Ll5PXxmtju2TOKr8M8yxOyUSnbr53bsrbG/2JHPqmHOnX45dg4ITG0ygyHo
TcgTNVMqE83broct9dHjvQrB4H3OgsFfRS4JQXafy5Yc8vRbNu8pX4aigQpsOV88
jv3fDauZdHVLeY9svcZgOwErGnYra44hGYY0GwVCzIp37EIMCZnR04WetYcHBM07
o6wLR85LUgY5eFCLcBxoUsHH27oHGaNjuidwOpZYGarMlgC3FVRDjXL7XGfRj45V
/psiQnxccp5vZwN0GQwAk8c+y9qRxzb3xxEtNSSC0v8Yk7gCaebimCJ2PV39EsrK
vNrleTthnALL3ETKPBLNrBo6YaKjw2puG3ZTKgAw8FyJHuIYwZtG5JmKxEINpDSj
sGHOBxngOBtfS8JcjoNRqaXTV0ORRRrzCAwI7URH7w02KdF+pKWT4utkMHNVwOEp
tLhFaqcwF0cRD8rQ6eJ2hf75v1oyfqbcRUwvMZI2aKu5JQ0FNVX7ZG9j7rHukAZ7
bnlEFXT+/TDAHsBGvG759LtcVgBqEkJEFa76dmPH3z/bBPku1eee0fPXx7uRin/5
cv8fQDDhSnPOpQFGw/SCQfIzZhbvGuH64OAGQu4g7K3zkaHy6wV2eTXe6EbSOXtR
oD/10/T1Wco2aMuK34Vw5jrc3BvCzPI8R1cNfcGF6679WkjXvrLlXW31g4AX07JM
Ez/dr6SyyWASfBu/0xV3kuYc+vRK5+EWtMW9rvIlSFlcJ1etla76aBG20lS6r4aL
RDH5VR7wUuqS5kl1QQWyVIQ2o4/3eOQVl1HFfLsnbmT8W85sG4uxVqBVNvVSEufT
mlwDyWOzCHUVTWzDghxVsbsPpZzlkT72xPYab8l/OtY/VZhJY0HCgRXWk+fflQTr
j7MgumrCYS/0QIJdEEJmG/rp/9hqSd3/5HwiI42qH2EdWACFjSMHWAsjvILSZ4V4
3Y8kME/Mnpknf3gsZHrldJqSWj82eZaHlB6AJp7i5vdoCjwQ0KyWgMUPnG0jsXO6
OhD9OXmwBl7MZnvsIque0mCl4h6ms9Lg4d3rPiGapLWaYGd+GWMIyHrH0H/UosFv
NcY8alVpXjK3rTiBIhxyIslADa8xi7J/PIrZ0AZZm7+mhdYY4KwGF2P/KTFZSjyz
B+2rmQAU0Oqu/F96iXmcIw2fX1NVzLmMFhj/8N7wu+Ug56kT6GgBzok2jdjomdrX
rNEKuXEfw0GRT/AtjhbMzQKdUVU9OOnzVWQADts4jArG/CQ7WTa2hq+iCYU0nE/2
5XlrTQ7Lfr4GQJjqKPPFN+aQCu465daPJ3MYm11Rp3bia2scsINbz/qD5pz8Qw2D
bcujhRq3yS1fFW/y/0DdIIlA61trZIf/iVXDZ0tdbL6A5+s5I0YyJBTSxCgQ12OK
i2FT7+GuXgmFqxDRYRmNNpTWZR3KZ/ewTWBAVKV4fAOGIdRPcDuJIUIYW83r8pz2
XzmhcCOVs2FHOHKRtaXBqHVTlArsO8FxivClE0tp5iHhWu4aNljO8282AlUmFm7d
kundyxuKsJ0Xymgin7AhusIZ4ShWmWq3XnGtF/zud0eg3xpcV4Kzs38tS7dTOfps
aKHPiwDwgiVgEQeY5btvnY95EF1BgPteXXbTTzOuhnfzUz6GpGCprargCxNetlQT
gOD6bQ3nSGkkAEQEuaSLL440MQxxdrQIGZ216YuuarQnwbXCt9A+Y2rlPtaayE3t
FC0VklackAC/1/8kfVOV4mjUzwXgPtbspXyWyZ0hAyvdYxGcattIFLB1y5SFQKfQ
EUqc/gtM88e8iLW18jpo9xG8O/hj/2gjBjcOE+Da1biIvQZqwidWAxDRhiAklAPy
3iZp0yJ3UCjR6w3LU2gKuG7lmALbQdwVoO3z6+qHZe/fZbTyMGXi9NF3l6WN5iO+
+p1JKTP9x98jkxLlKiKuRNqxjjjlBmpKWPLnfiWzB0sXa/aVA+I0u3+fSrgpL81a
9GrMzZqZOgECzz/39WYgFhznUK8OwTUWQJWNhj8OqDfRoOpXYE6ki20WXkduLTNm
MmzDDFGlQc4vPBjPNj35dkXlVEVoaE0JnxgJ5lhwKyqKvc3t4yktVBR9J/WJoLxQ
z1xCFwMcnNqcYqA0oPmVpItugiq/SAkOI/mL4xp+vDfN3HQNLf/zcxXWGL2J4x3V
Uhv6AVrY3BkarIpOAfsGjFVjPLzB5W8XWhpGFkg4XnrbJ3Zw7pjqSkSq6uak91ej
4R0ESXy2xLSoapjwUEemvK2WFKwlVFp/Zp0d8umrWYXzgytw9laNOUeVLrrHt9bp
Lv/95pNenZY586x4ghMksH92OHbry1+4Rc/iYTho6PHHUNDSh+EtuebHwBMqHuM6
r4u42tkv5gLxyNod4C8ezrZgEHrNsur5hSKBVEvc5dWxWwzYnry/A9ONCPVOwMDS
xoU/UXy2ETja+K/KkyN9/0TymytgXRE1gkh4WnON3iko5nzCoy7VI9WX4Bu6J14K
GZDL43bn/634DF2XAcevH/q9cQkuYI8y+/mmW770YL6utC+2cO7ZwbDZZSjXO57v
5fEdiA3d0akE+/4J1Eur79YJyu5tq3ONCSB7pRM7jpHaCkETu3cP6XgsepvMMtAN
21bIAIYIAVme+lhte9fBqf9CK0G2tEUZEnF9fnTT7kfOdkiEs8rndJk/GGGEO5Zu
7hLOUSkale42DIDS7efKBHH0A+T9m7pvzXJzK0IclVjULN+xn33IpoSInxhYH9NO
HfTcHRnVR3xdGRHfoxeR4j1XhbFSnl8RonKZ+dcL7U0DeSF29z83DspPbzKhAAso
o8iPdFQbf2eaoAzKMfDJ5PMYwrElmugUCo4LI4A3zEQk9TcQ6rzIDbhKoh9lEzYS
quzd5WSWVDcEQD7yfRnBlNpta1/V5cV7cv/0q7pShuGEeOVNAUIRGV6yzWyfFTud
2F+nQHR8P6gz8gTcfRQxcbM/RgyOodTmt4d3dAudNFT6vdrV1KvEovwdXnyLNOMG
zms8zesJ/TN1LXZE6GPJ7jpJ9yTQfQuHScnfay5tddWSGEBP8aBnalzbRV2CsUNE
KJ8baUZ5MoxJiFphgRgTJJS0EjWzKRTsIjCdpoeHMBmm8IEUtBJDhKh6GI3NZkmE
+J7Uf/NQus6PHv53vI2HCI110CI7QSyrjesJ6FhspV9a1QX2H/NLv6ZfW0FeT4z1
7qZbtSW1f1iSFZqeD8AGfELXksKVEQIBLegOIUya1V/LOXUFvo9h2nVwjFgZiIza
PRQqN1hyyko2CibICck+7qDgdD+Qzsj5D4KBGhBvOJsBFgEBKY3ubwXRMhG5r5Gr
3jAwDLXcA+e3quoD293iPK+CfmMn4g2RhnT/rL+k1//332iPhr1UwwgUUaOmnU3C
Kpa0uoHrW1A7aG8BU6e+gc8+db1K/OpfKO0nEKL1GiFW6xGdYkG+ZE4KAWFFjMrv
HNM2blLZcRxDD6daZsTrsNjg9NFuBFkojtG4pISQpcKfvPpMzkB35tKato1UFw/d
GmiFTQm8h7/LdBpZZPWkzqkKeRKFFHtuSFhRk7450B2a/u7GkCBMYgcrLz7gUbqX
6LbCphQe3JjHndja2u5RCrXTIiEXCu6ZnXWSllGACEYcQ/cknrYjhZSb3KdcX27D
BVaCUvej4y2/N0zH4uEozrOCGWStAoxZe1tjcKymxxo7MDnvjvWMu8udppP4ywMX
++6D+7uVTxmOJ5hQtiRMBuvubziEozXDxiYqEZimAOEx0ZgErnOeGVDpNWV/Qzfg
RDbSFWqtIvA5VNENA0GbT72hbhhWy06UDXgOPam6SKINyEUJkuRLwLPkkaxnicH2
OM9l8d84zsH4If5DvGL+xGgAgZn/bj3bmea4DEKvbzro5EhZWZH2NsO4IrPj0fcM
pg8C/PPw+ffloAI4bEukeZvpq2X9VNuG1lVb602Ir49sKPg6BFv2qVuMESpgNeiq
E5Cj3trr8dVj+NkP56GPXPkyDsI/9QVtZA9id+fref7kl93grwyylZuBRFG8fDaK
spC8Yp21ab9+VGPgsBEpcvh0nXupd1ebzx0ditrCUfzwn62FOl82jePxSSD69Tk4
6ZudcAzzHBRv2TlguoXVttMG8uqPsTEjuElD5trm+3DAkVoPVnjcpXqhosqkAefg
wHZ2LQmWkKNtBAF2HxGlYAzwparZivPg3uS7fTrsivysK3+XQkpSDX0pbST1UGB3
650p60UaIRQgqUe5vYAnPlmEONBXC57S0dwEZmDSvedUriEL12mbwhhlaaHQTwbg
DmqRMP6hlAzAL5dp2JJeOcfpb5g42qOwx+GDhWxc1HSMV86zzdh1sF7oLPeecxL4
SC9VixfIFiBUNm4e7SV3TMqMZPgPPwcrmcBDzpysIJx6ExWQqlgica4ZqDQsZVg7
vGtUNVO0LNsZQNRppY0PyCU1tmlrIg427lUd+G/q8kjtvy2c56xNrLB4gFgZMVGd
i49i7Wb7JirqHevFA2t/RswrKdu3p3/Rwx/4BF9C+wmsN3i+HSmWFmK+c9LVzkrG
DQz6aYBRlUqTt8oCBVsmhsAZ5/D+jg0LRPzlkzbNSu+bqZdiCdivBr7/IbZUeEd5
rGci5jZr90VCFsON+NwGLNc5eNBEkMd7B5Vu5mZao/ruvNyVlt0567i+yuEyLC2Y
CmHfewADNtnO8Z8vz+s1Q58KYnNAaZ7nT97H5Hu8F/W238Fp0gColr+lT52vudQ7
2IddXkz3X+50I0Wj0qUA9HaGOpjX0PuJ0tGe7u/fDI1hNowMqtq+9lKlKe5mHrTZ
jFDwizOR+LFCqOEEo/aSMHsHtRJxJCovRhNUcQDmCJTxoML2BiEfKlIfWcZr1ohv
hCwwAZHaoM7xDYSY5dOEq3tqfh4KlZQ1Hie6ffluq4MqEdzW4i3QWlWry7aCQKJ+
dB0OaNcLPcKpl/50qOJrpWDFwA7Jv14VTQYgmUP0HpVfV3Mjz1t0lHfWa+PtJCD1
MGnFy6hn+aeVOif9EYhV0wUOUgMj6UexYJdZFT5reeZLy6EajejZyulB8YoNa2gh
O52sZdND6hvy5K3jphpmDVReheJe1Y0JoCI7sJCJhwr0rHbNleVlZpOVDfCY+2CG
sExLgLgzfLabd+uL7pL2VlcOnoMsUC9s311MjhA2rPMMEB85O7VBX0M2DVylQcIN
9V9EdgW/ezH41LINopj22WV4lQRTxYLL8kvuUy8gP0F9MxlUgTC1f78wQO8P6puA
0KFbSNaUD6H40PDxhCruYpammkzZmA55jVPaJph7m93fGCXVRaGR2SA+yDBgHYVS
3FmF3UFx22ZPlIoe0PMlwmm4ZhwmihXPGOojXAi7DI48DklGE3czZ4U1Ne16mrU1
M8pFkUYOSoUYKPzDKkuofuCT32V5pxB4xoy3E0mH/OQgpnExfyX2+/ZJGvPqMyM+
UCL4URoLNCtJaBllTOzmwhK3+dyCPZKc2Sk7LK7IXnMD3n2EThuoYxTctoA6x34s
7ZuAZQQOWBcDe3e+SruKlNHIQo0C6sZYFVcQzpZ99ILtK+xNoiPq8+x5PfqqyGqv
u89sdr8zr4/rhP5JZvy1QOgnQHYxqLtSlf6VOfcWk4iREgoi4pdRxrE+XLkk6Pb/
2gIrshnuUhtBCzVc0IGIiRMCHUgbiJJD+jti9Edixes0Hc26STTH09pPnyZ9ulzF
aHmMQ1Nz7hm4anHAS2OV2i9HwX+/WDQEaJDEexcPHySc8wJeFdozndrO42aKpGfh
NQihAOOCzNfIjyqOVRhzwrxg9QMdIQHsLc51pxtOkd4SrxJ66QPesIG5tbH88lac
N5AoxJvK2R+RyCoNx/0BGWBsP3B4hckqK99tfuhnZKHhNf2e+kQmUpe978A14d5k
YPAiAv5InjTJzRLm1G9EgLoXceNYgJfdvb0yNejXF862gGI10smAIQTbvVxjvEnP
VjiL0fdwobk2Y+Ph+mQonTbdz6imgd4q1wqDwZNH5JMf+hPC+IvIfRlsW8LSzZp1
Wdh4APT1dgBKfAAyZ3OqEFlr9R4JVlYQDKUfXjfSxOti3SEOZbZeVGZ8h6Pu5Cno
rt+a+3a82iGDTRxM4aa3V0OIo3ppC714F68qucKUZpPoNJhefQhf5Lc1zL1jOcvo
0fX6QLdigL9Hkt4n5CRxqNNwzA+mbpIwr2DEz1UqW7AXh9eW4afq6RL9V8LnDkrH
irFidcHAZwEaxtCZgY4e3zogxplxrPBdP+MiYgO3Jz00Bl6uwxAfO9PyIZ9zO0Ry
V79q8TDTsrn5ndoPkI+s5YVioJX9dDqrxQVVvRnVp1mC1VtwczdH5jviiRVKzMX5
WmfiS9MwuLNMQt7txUBijW4Q6K8x++dGePbtkmI5xGlo8MbRUsCsVu3XgV6MhpI1
F0HQPMYewU5uwOd2MYpxhRSVOvuQlWE3WHjIhjbay7rfQ362STghUlKEBJih5Ow0
+F/jOeRYZeQ7MTacrEQrs6W2S8/Jvq6+N0tAK3g0IlO+ajfalz/d5Q5N1ElNHU95
OMDgFr3T9bT2orTP84b0pDSptL11OuJ7K7QVhUHC7qjKQ/CSggU5eY/Wo3aAELn+
d2gVnDQEeARV62tpbanhCQjoD0oyeZzAzrc+zN28s5LbmH8uTwOOwT50klfKI2wG
RmaOnRwivawtdlPtlBX0atUoFSe88ubZjknygsMHedMPaz47ITbF/LGbkxt3Jr7L
bTx+o1CQ62VlCl+Wakyzhp99wkP9hLEvhOLqSBI4el+qsTGspB0hylR6YNIJTWGk
aq2NryphP09zG/9374hJIKCMvQ4tcCrSYxe//sFWg2gFLIYrQ/Rd9lLqy89f6S9G
6+XGp4aRS3QceeqsZXeqP3u9R9ZyrX0EgQoXOKxh+2fPvLlDuDi+386BB9nVPfV3
z9FHdbCvgjdCg5m1L/rw0NVcEjELG9z7YZM7sheaONQcimJPczqch9wyX+Hupzpb
EZjJCsYBqNOQe4fUwj8wwaSjk+lOMIlULSV5K5yOkxeVcq8r9kb/eelDD+Qi3JuJ
j0rkXxtbcDw41WtLb9JeqaOxn86IUOb3rn80IoeGgl/7fUtB9PWXtqnjRKHT2ntc
f2Gxbgn9GK2dlcWOI9rM7h1mOVaAdbGw6+nXighZYECgH2XCfYCZGELZHptS/Pog
8/UC93Y50lPlm956GCgKF5GhH9Jpei0a/sizR4Lr3F4B16HyzNEpR0RulGxAiL0f
sU1i4xO3kexHeZGGH6OWaxHVdJmBTTM2EeZMAA6x/Wmaq8rFQ319ceyyezCwSG/2
m7OBwHS3YwQEnDPqFjvpV2SMREp0F6CMMmMLVHLd1iBO5Kk23MJuq80St3pUxhco
H8mtyCX8YDA/TqLvO1PHhpFXcVOg5+cqieA/9eXiibkBttEC1qWeEO/r/tpuui69
KTNZIIFZYHqwjmAXCkHBR8E+OjwCaiUBnZ56WlhumLsSP/R17e5Mwx+ElJEDASsk
MPFsb/65yZkj+Pf8xZHJoA7VcqsYsR+/4E3OwRrxwb64JoR042wBeDIHUP8471pV
6Xxg43VuWzCV3mohwiTBWlVx9Jn2ykOb/DL45BJVsYVz1KBNGC4KT9aHR4Weo9DR
aIhMAQ89jgQPB3dg9RaWA0T9ptMu6HMOpGj7O0QFqvXx15D+AT1VgkZytkIoFGBx
sPytm+fHdGguPXqorZ2e92T7oJkqA28be+li7R5PKMZFSYMBrFzEtc+qftU6kvwV
9MVOD6sfnJ529xBXK9LeaVdEMiwwidV9IktYYNRKIF2r6hu+RZS+6o9DyEUy2ENf
aWtNuC0nC6jA9cV4rZXbA7JdAemJry7GgmIZBiYsyKZjA1u5x32ueCvriEW73jgg
KWm04/T5kY8tMH35oxQ0o2D3futX6vUSJZxJFGCXRV+Pzu5RVh4hfah0mllvTiMQ
sBjsKBSIzrWKtnzphd2KA7pW049JkLdiZqigTm4Tp77yOCM8QwQia/eKvZpxCZ/g
vJqIcaY35nlB4U3mW+DWi0+XY5W1WQ4kqZ7cZ9x2qdzlHCqqQaEglfpS1dFVzKet
RGTBuIFMRBfKN0+uSffflpVIDUPxXIMWiehGkY2X+uPem5h81nqzhNovNARSOT6x
qQV7LokJopPT33wgkJuVonOXDd5SlIyzF+Pn4tRDwc+IHT9rVzEW8fviDng46VVi
+RxlANF+Gl7L6A58auft5QQG5DwILqEOenSeVNBCWPYTuw7EfZQk3urSImJf2CB5
4kbvmjaffQvt7Dzv5buql8zDLM2IifJLtm8U41QGqHSyi+5872++xlVQwTRwQtuC
1XtuLBsId/CUFvy75/i1nY0LiWb7Lx3MkolUhVSWKJ+F3YexG8ynmvkEXs850Yyd
6wActYJVL8FjIM3y58MgLHBZLvNqHL7IhPEpf0zTvbcGNg6c06dmEcapkU8vQVlK
cZgfJJ+gOEZhhEhaWg6axQq1m7HycYjGNN8wh7HSfzJ+hjZypS+cUushA4ttIsip
//GpInCcX05p4Urj6vOyHRlTspdgV0VtfWunx5eoyMgMC9Bl4C7Koo39UuE53FUl
Xc36/+E3ZgeVtgLaBavFMwtOQdGtfmgJLbgcr7gVz0aGpRiPq2Lu4/0g+48pYNB0
fSEp1KfCM/s+qLQnt8N84xTxsdlC8pbxDORB78rcWjEMC50fPzRDXl/ETRNirhpK
1M5Wteg5dRZViMwCfA+ykLmS+mbv0u6klw54dIKpHtwUxVVGWxgyvjsYcyVbN+cB
PzDUGIkdfF9EVrCkGfsLH+AFGqbJv+0poU+mUObmSOqYDr85OfNhKfWyROb1gW9Z
SFb8iJEi/dICqZ8weMtAYX4onvh4ykdnY7+AnuZ3QZReg+vm2CWkzL95aHWLQ+na
IqxwNYo6F41VTsYKJoPHC4fQ63i6dgAsT+J+gLRCi0YuTxbzv76/0ygUNQqAIut1
7cLvIt+RYt0YcWF/fdvq/ACsn1Eq+UJvTXmyJaZ2b+fvFIrD9R1u1lQ3xPQ8GgHT
t1BFoLc/VyeROsklwAEPvYMv+J+Qz6MmPias3Hf7/6SNMwbah2WfHjY+BGWDLww6
e+C7XA1Dmx/D4jezEyNJdR1YPXQtNL7xvZHUeO5GHV0mOqmjmW/1QUdVlDaHfAVE
vGWrC3/sZNhQHUKo/+qhNebX9ggpRWMZ+6XRKCsh7Ix9nKQAXhrmZdjf6jXPhVtW
USRj9p19UGyAqn+T7iQ9DaeVe28ybETvQyTmtWVuNhtf/KGnLce5cBj5YCtcoryL
tHsAKQbMyZAyoovcqfIA6p1ecqjCTV4aMuzmdJkIudhXIW0S5Ovy0Uf35f/xodMW
EMmev17qKOWgDoHsdZJuyjMJGVK5cWxBidd5kw25vxUF4NINI3Zj3DwQaJ0gTL68
sKfAIGvaAlYlAhMNNRZhDYUjscRKBDmXfwb1SPk2SUdK1X/X8/ekGJeUSwpepGF3
+BfznQFmJOcekKLO6VtNKEGva1qx0bAMK/QBrac18vGhWk9FtEaw+bJIYZ2688W3
cT2s9ixrhDDs5awow20wskxr00jAfiY8t5h8LIYpxH2v5acawXx4kz7sHNg/q7GW
YbesKMAlbqg8Uid+/JfHo0VV28yHf/xQuh8rP8Y2Oaoxwud7DIiig9OdrytL0SKF
7nwVfxTP0gZGUKb02NagbV7icxnHd5BVumCkVwa+BVZTYuNjlq7ur0n/YJP0Xh7I
Dsj9aFiuuhRtrVo8Bj7DLJN7kI1b0bgRKG/sR4fs/Nr4S/1fgdylHc7qcIRKZznD
xKiblSNGw1apgKKgyZUNBe+3LyAfK2NeLcGq19YzPWfI9QfgcftB53oWD2btde06
OCd75lTQ/9dg4jMtN65k+p6fb36KuutJf72nZSE5ht3HoleKSH4f4KNBRYiMn9rB
TQ3IEHIeCh/kXGIepZ+P7CvC4GoKWYCWlPujQ8BVfWlzwYzLmYgkD3eFBvB/FJrX
GJ98apuyDqF01Q0hjLGApsWtVpLYWD7UYjYpDPnzSUBczt3MyXfdsY0H3MK2blgE
4kXzc/lsfRpvDNDCK41oF0BgygPUcV/EWx8u5OBqUo6AkYvPtQmCGHVhOSdTj6RI
iq5iSTRvWILElVNWZCgyycZcu3mC4Yot5SKXUOIabpuT3Olxk6VzIVLUevs62o/h
bzIhIoxteIePX4fOobQRBc0jkubzx43MAU6SbN9frFG4wwFOvfyUnOLhZgk4WUGa
Yw3cbhgMIFlG4bLf0NatTIumPbTATZlthpUWzWbYSOiMXU2M2seGeGyj25E139pZ
l8Fc67udgqv0i5JThclpmSEm09GHl14dGlqw7lPsVFkLb9hOFjzID/5R58B7q6mY
nTzbwEU67KeXkIOU94ngA0wBGDfqrQQrH2C3z92R836rzHuTPT/spUNjwCuW1udF
126elgzoswvfLBMVe5wbsdsRQZSRH1BRa8H/umRWCQbca6sBO9fWmpTvdpVclsln
3N1rW51ZJxADGQdZxMoRRQ+E8mBOlgWytXWoecYxjWqIHtwFQu/CIWI5zFk25jzD
y/1M6HlogHGhgIy2hHmyh8A3a00nGT0Bl/UoOrT8zurt4oXLoq47MbXJgSYVsxzB
+nhGVuhKSNBzXgEWKUyfNFMl0bz42WDucQp0u/uW2ws8tIKYaMkAP68V+7mjBF0n
SPj41zgi5ccrCwSG8CMyhSgfkNhfQd0xaS68BdH2c9MwTo0w7tU7VS/AnW82cetb
e6IdIgUSCtz9ZNvEZNFlP96l+h1HBBTZo5K5333l5jN+SYOwgbe58Unzuh9Sn18p
y02T2ZPtIQATNJRRKQJqHYlOnago4ZjovxeXTT/lNHBj1kYxJ1ohltYP6OCqUS/K
rA1t0ivtnbwt94UQXwlE8DTH10Hxo69B9PGh36QEYyydtLfN/xR7ppn61FSiJjo2
tETqCvjSy1ACvc7nVAWT2Eq61hQsHcgVk3tX4Z5Sx3FCCAi1tiCoS7rLMnU//eUu
hNm462o/RSfC20+CjU4XIasumu3xRrJ00DDWFAXnYEaJ4qXYy0APxlN+xdvR9Pvz
Cew+oWYJLZ1qW0B/cmFdaWOuiXJDgr1puqa03cRBNtVXjHpYjUSk6jxzFsKU598s
Y5QVNUdffmZdBMpTPNR78oyPeG2uk4+SBEE6UPt3QH6L6RbZJ7O3S9hWISZSWlsa
bBzm+VkOuK1oJ7kliTGbCMKsb/+/IZFXera3TTs08rkHM+rKpTQhmP6xUw04C0hO
3/gpqzz+zHk3Io92BhwT6BEXqrbuTKFXjqbyZjLYlpkAMnRRGjgwTCOekbEIXnu5
EMegtvRATiSM8E9Mxh1HcQ5QYjNLVf04o/gftrSaAauVh7zQq7S4RPQdn5QYX576
eHJeSIpLIE37TionvDLc//HtHCJIJtLXUfRN75JTnU2oFLlHgY9R0FqLVhnAZ/7J
pewBeLdK+gnadkEhhgt+1CwpunWc6AD/WLW+2rKLLPGyNmY98gNTciaR3RYFGsOf
KppmBhUZohg7YCbBBhwLKiKkzt+rT3o9Y0PfkBXS5GT9Ml50edwao16vpDiBmikD
/f4n0g+YHCIz6RuVE4roe6JMDWeItR6Kr/yt0emVLrRhAAzbkugr/ViGeeGN0Nxk
MyC1fZGkr2YcXPkQnWER2ncw5Vs9uMxHXInsBGLEsoSktQ122AeYyYZKQcJl1CtO
Ftax0bAGx0qw6qd5cbLoS9uIaMK0LMqpF6vQpCbUlkijaRRYlBNzKyEIt3qhXCDb
McxK39LAd6U+CSE+ovO4WQqWy/P168iNULMU8zY379xeLkks4x+0kaLQcrUlKp/x
Oke+isg0Xo0RV+e5eifkP0gSNiYsjtdDKTC4U8SYcWqw+nlaH3dih19HFEwhPMyS
c0spXYfeOCsEg2mMqHc0LVFxg3y/ExLZpP3cIlCSud7QyZzNoYD2VWGGsoSNMLKK
q1GCaLfFMMIpMDeQdKmrAQM/s6mnmClL9lJ671n/a+y1BVqWdnhRE8cF1iJi4m9n
RT2AdOo1RoENmZCBb31RqbA7aQrecXhLae5tBKgTgG94LPSJ4LsL67EgX9WjEw7b
i1AfJgCwDZ1aBysQScsWx7A40BwYFETHp9rBKNQSAIRsPOP5eJEQUUkFF/zZZemm
p5wj7VSpZdjuwMnx0mr7B5DAwSUqA/3ZXS63vkoZSkvOx0DDdgYBElMczqo6zW9D
KHio8Zd27o8DpbGNpdh/jqJniypL7VZs8JtxUDQg2lkSwhxFq494hGkDxG31Z2kJ
tOBW1muj2HP888ggu+hi4lbK2PLZ5iq7ieAHesGmepdY/0cCpvXtJZYCDD5N62Gx
Fm0xbXnsRmuYuk7HIz7XTSRlhJLB6iwvgSmSQJa60IgzjUepWrLRurCcX1kif71c
9eJzyTX+pQ5xFFHsl8g5pygCKQsrVnfBPOegcZmV7Xgeg2PJvBmHLhcoUGkIs9YQ
EU+MXAyQmKyUGjccnrktmG6PAVo564/WAHItrpNMlA+WGbfwmt8wcBnPE5b2U9Pw
B6XjFCVFEgRPK/othjJIBkgkST/IZfIiDDres1PR1RME1hJkgWgG4mthgajwlJOB
vUFRHP7t4NJDESxNEstZltBM/YWZzQTrH2jmaweJxnCekVKzyLJJZJvmBQoB2vNd
whpsKZbxhSzc3k1YJ9TT9EbF4t6iRgLue4R1OQLkq21FsF+TnmOdCml6V5iXtsuA
ng1DRdc/uR+Eo9QLimsIpksNMjyGnnC0+FbZoEF/OO/oSsbf/NZH1P876HWq9VEY
YZHAfAXhMBcjOqwAOe3XiXqRW7M36wAYfQq0f9mALT9CnGgGF6o/5l0wgSI5Icsr
V1Er42o3cR9i8LPgTyNbT6e0WHD1d92dNZfp2V6VKSFUq5xO8z17PKDLIvRn+eJq
el458nskFlPOrKDmHkfTXbGZsSvO37NN7RNx6ZicJ1/ULrRxFrfQkW8XPy9EO3Mu
wE/VXwCyWhX9dXwRQAjzLmVxHX2/eVQfc+rB5gxn6qS/lQVS8xhN3w4h+Fk4or1d
42mk9MWXZKIYuthnVKp8Jt8GhLK52E1lBcWDIMlR3faagh984LIjLuEOaJWS9QZS
E1OES3XoswoWagg9tSnIRjbDB3EFAfA4pWMcYOYiSl4TuOoSXEwwsur5147SEHYm
pPyHWUu3j8S9cOIx8oQqDSTpWVJv5jzwFeaOzJwQQ7m4fHMmWdZhDsoVrJID6p8v
baKYGMbwHVAdvygXC1wOU/S7/JeY5O1t2y9eA9YH4Vh+0IR/WIDyYlrJQ51ApP1a
QDy2RAAJPw4/O2Yx21sLeD51KiypBSQmyOweG3QlfNhRsyq2zLTbIe31anpLemzu
Q2nPGyo+Dy4MqbfExYqI5JcGFkrDamP02XluMbQlG6gdsy4OsowdlOeTQ+WE3/A8
5WJQqcbcwuKXWOccF7uv+xxOQNMNFtepZYXgzKLyoItaAJR5FL+DEQ6HblxKwuqA
c+VISInjXvOzUsaUKRfmFk5nAfglWKJlyKRGegKJMzZYVKnCtbbLYSB6jOI/HFP/
sdVKj5DZi88ywDZO7WmqfNlUIp99d+t1XnE2oUrhgQvLF1Vg50qxzhM5HrPJw4R0
nKU0/VKiQba+9zxosPDU4+ni6VfG8/TouPUn4Fs+pnsdf2K/Y0hFalqxN1JXYEw1
MPjOrEuBITr5iJ7H09KmFH3vhgF9s/PCS462/P2lTVF4ia+2Ob4WFy7Gx7n70zwH
sHCboBTLXX0UkAfbucFncoZv2tQilIjfg5HxItcNH+49ZYCr1EQdaipb1sr1Za3w
i7D/USqvXqAQCcngveKFpwtgl8pGYsMoStuolL0lcDskXzogkZbnTRs12+Rd1sej
GHax3Zy+QMNcwTGA/BfKgrFqqb9h9HzO7ffU9igWBEeyGPr7f87m+qCTjdTgZ/4p
282EYlmFl7w0yHN8diNqnC6g76PbWUtso4BUr6yKjBTwUv8HhO8//u91OZn6WZV4
6k2mzkPM8V3ZK7Yndaa4fHtc13U+nSJpQ+AigatAk5QrHSewHaOWd7FSw3uMw5xf
rf3R8Hh/79HYS8GyBmgOZ8G5zKwEnv6WDg9JhegjwCCtY1eQAogOTWcHI6bVyXUq
HDobeZG/R4+0qTLRsKeUNwuhWbxyNxiCtSaPJQjM+8kJhKOW6pEcsrewxUuiZvWo
R7LycHb+iO6ZQKiUSqKLtXegvhxWImNqiY27v4mfcyFVXt2fcefZaLnZbhJxFGUf
1ugSz/FsOmLa7s2IAHhFjDaI5BLHGIrMeavNZLTxa9gU40wIaM6ZUuxNiWh9H+Ua
ndAX3s7U5izkRmumaBYd4atiujG3nkU0HYkUZ2vEO5fv3u+11OkONSryHzHCO3lh
mM5lEQ/QzTXZtQxYNB0OCe0ab7I4BCPWnsFe5aBrhxoH8Z32qlxcSxri4R/V3Qn6
Oodg+W6d0U0rRehMahX90yUm/FJZzllbPMFPC1Iur9/oXh0h/9A+Q7xdCL/I/uz7
w4PVFQUl6GXcbnopwpWkDO4BrDEz/EDi940S3ondJ65wnSBLVkgnSNe/oZSL0Ig5
8gXqk0g3yPTrDESd3yasd4eoZIQlfzW5co6cj2+LTEsbDD49LYC/ZXSJ9gN7lKzM
3ulPMDMPWZZ2R+0QgP3/NUX3j/q6QqlHspQ0mblbmvQDxZpFhFLp3t+k2zX88w+Z
m/eW01zgSEJ8AMxOj/TdZoy1aBn0ZCtX8oVPqm70+rfMUD2pkpEW9ZqYcg5m/KLB
71aeK3z2VZak8Gq7euAYj8v1i9yCI7Kyj78aDu9LAyqCbwq/CZr0SVKTobBZ7p5A
Xko2naXqPaJZooSo7JNxhQHYoMKN44hzWqQMf7gbxUmIP7e/ziWLYb2hSyCK6K/9
UuaRgXITGwsn01oTFPcgbQUNYdF1WqR58xi/AUgv9LLsxg16E25tl1DfcNUkXOtw
3lpOElyyx6oIyaGIFvcHvLd4BUvvKp9QvkWaZ/H/8gAyavgiAXB9UnNi/ZCNWt2y
G3bibgL7hRIcYGa1RNKBaCByvT765+5fra1oHFe2LmWVM3U7OK0ZjQz59Rvr3B30
Mkab0LsLVylPl1uiYiR9qX+cjL2ewksVXrrHEfIak72SLRzd3k9TP9tGJEpN2GfE
2RpnQUbfbkxSRQqAwWivZqxUftv7H7hzkXvz7MK/38mNaf0d49uACbl5I9bylpuS
xUNIufrwdjNKOFEpTwOx5IIL0YiRFsPiker5qBvauUPl2d5poaeUJG87WxsCLI3V
F6aYfOiB0f3eH8To5mmn9trZoSTtYOVQADbYjrYD2fefETtX1hdraLfQly+uV/EW
fiIh3m+ItMrj/J4sef+LYSeGqb9krWIyKKL9O/rQ31hfc7/YuOsCKVEkDd3g8ur0
mJFv2MunQyFUBHB0De73MC9Epxjfq1WEVc3gnBX3IwFk3YIGKgxw/GDlvlHvhUXu
5JIjSxSsz46TAENmU+u/64fM3J+/l+2bT22LXPqZ48I/geHU3wwN3bCojprZhnut
rtFP/Mt+m1SoMohuTMCjH6hFxQEmA/tU7fAXXH+BeIUg1xLPfTG0A3YJLFDyo3yI
ZkRCw6h66hgqrEtp8Mm17kv510r6y2A0dxnmv+EQPUVB/Qo4fKDN6ibrhqSsTak1
rJgK2SakYsRUlcbjIPGyONCmREFgsy9Yfk2rIYkfz8fdg0UELb3JMAJv283SfKmJ
86pxuUHOpBZPn8zVSeQlIA5/RGRYH3gwmBa9DIJTTHXWzxXrywYqii+zx+n6FK/h
9/V8lLhwDEqKhO9GshrHDoJ4lQI3w3FyyJP3w4IBpTYA9D66iFv09nhDruXGIYdZ
saXIanQga/Pyx0ih6sR+5G0dafkOjlOVqIlcKF9Z7ThoA/pB12XL1hy9TRr7LAXM
E5JJEWNkF+ptL8ZJtQRRjkgZiRQP6aIvv+YKAWATvrwsHywdstvDtgAVTFzuJcMS
l0fYCFYpgAhxuPhvWNd1ZKO4tdnounk1DRhJd2FG1gFJc6YYjpZdpzFOx4RNbptU
8v27Y5GoKiw/gWlUR3o37IN9611eTQEn3RGOzP0/sN0911HObfJ/y8Xl4cm9Jwbb
fVJt98Vp8tG32QCT46IZgFr/52wVHJCAib5rRsFo5zVf/1PwtwK5EXf6lCZjqIcb
Wi/ROjAoVJVsEO4gD+2zBo7yZboeZyCCMKTd4hT68z4YjgaiZkf1RfgCMrsywXyI
XxKzr2wMaXW/uVWwfU7w3PRSgZG/wRqoTWi6FDwJX32oWclDX8tMD2BUITrsyoeZ
9s0W4J3wk83tFBkO4I5CTlfcjfKGSKcLfZqByNVAGltphanS4YU6eRhU41+fhdMC
TyC84uOSV4T/+AVSmQcV+/gsLUURajIOLbF/y5dWYaQLgV1Dtv9MOIIZwXy7U+2v
dc+Z2jhNlo7m54MVx3e9bKO3uVB8Msr7G4id9TBhWwNlrsUW+JCD0rfeWvA/A8Z1
j8WQSngv27Z0OdwAp7Tq6Mh4qv0JWVQ+85/28BlG2l+jo+mkgcKEr0SZe+wzHWoF
OjA+PjjKcb1BUipyIBeQVjssdXNAeCgtkilpW0jSvumO0mHJTTZQuvvXDJutEdk+
gnbaKjKLG2bp0HwUtRnQIY+NlTyA/sfR2xMUsvy7h9LZXsCgFcGRJDk8tn1OxwTM
97GMMHg2K5jvkceBb+jy74rQ/fmtkEvbcH3hxbYbcVXuskNorruNsCBRRwy6KiCD
SWxY0YrZHV8q/jSoSjdRbXyEwqRGToG/hBMCskJtpm5/zB8684Mt+BZEFWIYjRuc
u9fWb0KVIGfpVtqFoD+DZPgJnBBYmTdwSaJLYF3fCRlv2eXoICU3rXrP4hJQ29+D
VM22rt+iyBj8n2CL2+mpnT2yJJxyom6Lq7EgW+LVMq0vBYHdkJypoSN7D+mSN/YT
8wq3CJqVOOuLuOnXP8f4Vkdl4oD4FTceAcdtkFaGoyFRbpEKcFzdP52cZdlLaTap
s8NGf/LhR1PW8shixMqxrVDi4QKimoi9wHWAWW3rWceas095VOicKfc+WDyVTxyz
7HilI5cJ5F/fFdiqYZjzNQwhtHGQESRLS8IHpYs2aTZCYywU7oBejYuPaI1HYEj5
RFbD6VnAVI90GYA0QDAOEkBvflQEljq2+WrN3UE24K0aT16apS1zdUHGx96rDfJK
2PGFDhEk1PTeaOQRuimtz8t/d4DQiN752MtwPsI8+B937HczMUX5ghxuz9Kzy4/Q
4122DInv2c+5NrvDTxm1UkR2HNS4lBRcfwVat3zoguhDXnWKBkAqJklG9BlZG+1W
edFsxlEI9fqzSmD9sX06c0R1gD+w64OZ3uUKKi5x1sxz4omFhksayZuGhI9yOf5u
ZbXxkg11tPzHghBHvWo7aEKGNvQGESZWyOuiIU6bgDLrCmqMLiA/8T0b+MUKnOsP
3vHrGjUD+k69rt1C4sln+Ws1zIitkPDqdGIKNRPGvYDZKkoO2d4LXlVh1qUJvqcb
KK7vrqqNn3L7y15s/0647izRTRTUvtppbc3sGkHNOeQ/3IENDMNgDXia5pMVYYaB
COBmzcjTM+5RM8kewiPUYjpJredTzr5Rljyf6gtkaFBmP2EZHWZlUgMEPMX9stiW
Nmv1Uxtj2AjiNEAG/ohbk70TgcWe3ZsPgEoUt1NQZzHE+VgFB6JUbmrJNiNwsZD1
firVw4Grr4Os5JAo3sPZLiWGKnWywFgXOcZaM2jL+q5md6y+Wp1dp14m7EMzK2c/
CWpPWzE42sPSomUsVisl32wUaiq7jhA7L9lSscQei/szJtnuCOzaOzfM7neMOBup
Qdpwd/G8ZSHXryUJKm8l1UCFdVluq9zPtU7uOeZH0AwwzIXLf7T83WTOHDjtsdYx
hh/DWdKst63/pdXvTN2qYyN4MdafoXqn5lA8081hnt/xHWDo0HVMVcKBA0dTrljh
k67V1BOhXmChVaLysAANSrrviPfuvdAWlipns42Sk021M+r1J+zZlCkZ7rBSHUm4
/wqpixh+s4NTLRQxRR6r6FLWFyGiUTY2MFJNX/irqg/xXN46RWOi7CUVGCmF/FDk
QXX9rqNqQh5tc1f1K41GIurKa+mDNG7LnPwxiD7FKaNUXHoteHFNK4g4fG+s9gGN
JAqf1IG1O9shbgWL4GDzDMRR2pujTklSs0qqzg4mMteM8YF3pywvDqEb/YjeVpCy
D25LZGbHAOGCQUiTe9+kN92s1lmEHoEECZiwMqrBa6nW3zKoW6t71qKWMfNM2N4t
QAiyFGMsPDizCXaQppUyiDjAufRYLegCdrjKMNFvIAmkso07uo5AJRU61SXIoRz+
6q6zCAcfD+oNnC4cBrkk0ojD4QrPyWo3d+n/CWYy9mw9/CiLOLwpF5Lgj3PqZdTP
Xi91+jgdZO073eQigJqw5aO7e71xuL5UXb5/o49HWr+5FObfeXBvxI5SlZ5y29ZN
eUNpu+UVTJtEzyMnPrFCsawD3kSml+zGwi60a9DTP6naa92926nMU5DlcqV7L734
BK+zeAZ+ZdxOAR+U8VtXZ/khtfuNFtJp80nMsksqc/DJtit7dearTpI7cN5kEYCJ
gs6r4xWFxda8rcdrA5YVwJAU2skz+Rp5dzWRTwZnTLMOG5e+fv1ULBcOzvNUagZW
ySKdmNzgWmX1S3nFYTdqeYrpBTf64ycQ5WnUHnWPj7PPjK3btHNEBMDnSUcX1HlR
CVXRpVhRiFVYOZFFb1n3Y2CC157yN97jjuT73Ujmb4xfV+nKocpBtxbqFsMeFtkt
tjP1K5tELXWNZSi3aMQD7Mb/uOSyB0hweJMOb5aQCvbaSo/GIifUX1dgAaW5s5tK
ADUFsP60DRW16pgfMqdq9/rXmL7LgW5e6a2zNPCGQYfuj0Qyv6rmNqHkAZ+GaWg/
MDhgu/b298rNHxYBh9MNkAPjFNpi2VCZX8m+HFcSxkJbubuuD02AuoB9jMBikoni
z8espPy3IzHKel248UwDtZ6mcCftCedZveXSNfdJG01dCxxwdy6xLOXQy2mTdPJA
ty9+P7oy6oC1Q3AnPIYz/4h5FWoxL8548mD1M3M1oXXLITLA9evG7KoW5fDN5YQT
Uklj0mbnJFQjuQFU11tOyTV51o16q5pzysodLI7/vHXtjza0z+yLNgr4N4npbaCP
bh1OeHsXwzkLX4xkFEKNvbTqU4e3pvgIvbaK9tKjV655KtxiyYrauHfX9dnW9meN
W7ZCvfTP7RM1qO4fz5p2hfauN+EXiOm44VjIkA6vNpRzVYkc+C9ybExYnRvZ3EH0
cgwgywbGnKfnRTLExpbTjEfAoa1yDWZOss1odVrWU9zVQ1p7AakdXFZfVH3osdd1
CmLiyZO62KbuUCA4g7itWyNu3SXntle/0IyCuNGFBP5Cpw/Nz9O8zQkaonzT13JX
eTgkVglPt5OBHFcCXHpZtJr8a/aPnIgamon668gUqiYPtk+sne6z6LXJTUFQoyJR
rxACtFBvOs9RbaaWmokfZxhX9QCi4BOxBxdUkr3gRTCWhX1CVKpfYMDBfqx6NxlX
/UtLKL9Mh0bX2EJofqkmC9pDWHwgrTAgBYf8vK35/LdsZ6ak8aS8/hT4IVTEEl90
dZzNf3QFGyf9Z2aG00mq2j5YR8mGrhSuiNv4HKPAP4RySCZIjf/6tgqWcUsCych+
HbAozBpaJj8Vnjb21ANN9fuDuFDsadbKiO7HuXg3zXAJMjNTYasP3FYy0w7bu7nQ
5yeLmadV3F0SG8WtAuIqfB0rPN4UYdMH7TIi8gYEjwB/QktZZssg21Q+AWELSGJV
PX0IX0SMaE3mb3C1m0ue1z+DkHCuQe2FWukQhE+itnHnRpzcQpG2wJgrIyQGat5z
jaseYHyzDm9jNvkOhS2u0U6JSKCw2oe1EY5KsPwJhBO7KwGHBtJ/97NhUxXcRVNz
L+B0VIAWCBt8BA06Ih9OPfi5ywTUyso1PBI2DVeOqdR8yUDnHRSPj/CgAGm8D+cX
sxqLmLEDmKFny40Voc7X8pU58Z4Jj6YjixmxNLkOMucUk1YhBE9woGg/+Xp0ihx7
MWHzJ1Ee9wsd183gDc2uPWYsLoB+RIYEcxfatIW0tVDYAy98BUvq/khPiOXwBcmB
3JEMqa6MVgbOuRHhutOvK1vqXPsDjPZdt9s4uBNgm7buPnMOvLcp7l6wdcao7bnz
9PsYDhfpd04Ex23TzJYUQRvPrZH50uCl2Uu5TRmMdz+5jgBw7PzAN2HtZHG08VoT
NyYx77/BLG6AhSYsScADvLwXSs7gCiQmFfrr0OIYPk0ye5A1Ag5wsqpNSadlCwam
/+H1Ggn6ZBjDYM4rL4FSLiY3TtAffXVvjgR+eSEL1u2Um+ur+QjVRoCJ/g9f6Rl8
p6Zp/fXDQa7/xIkZ24THckRKmLVDq67GaGBuKUjbTW6Yeupr09kxyNbAYg3XrnTY
L+q3ZvYf8/Qc78Y6pOxvBaUFM+OwaVIlm14yu2EShS/sjfE8UAwqLnY6SBqcSKui
5eMKLNKTY1MT63mL3YSId8v1Ef9x9R3XsTdM7eMyWa+UxzE5w3aYFcaLO7FroTPK
FFKSV2T2dLgXSGScFep9VqTr6YVQI/IRp3Adg5qZcXH4oJI5kQIqZJb/uAgMdn5w
JgADoMDSIHqFcRVTg3jYw9efRb/qhaa+PYQwpcfp5b/KmJCTBQlC476UK/YEgLZ4
TYMu9ITfjaO5/DiTf/n5xQaK4yAdEoilIuU6dflr+ePfmhKK57UvqcFNx69IWs9A
xuc/UNByfbs0jJs1VQbsWs7SD/JrKWe/kvFZtBPiZ3dOKwFef0KmX9AvLwZ4IKro
GomOb+5fC1D8HgmrZNlV9jZ7P9L9Ew8bC2/SHUeQXKDzlL+AVpROKVILL3AEOXs0
efi1rvqe6VMl0+hhcR6tZZerv6A/RRnW3v8FcJQKk5jDMmd6QmIzZdrXy93rfMLC
7Fyve8CwuFvgCO4oqI28hkAyYQXuT+o4EFPlBEmft4xZ5/BUxv2q5G0UWsSXNpy6
g6mBQpesLwJW514VkgTr7jAfN3xaOWT9SCiCWBBjC+lVJAiW6kMsog0LjMFBBZKI
HywaK3hkML4BQGTAKVVKB5Cco6b7LnK8Ee1wWBYkuZOB8lQXOmqtX6ecu8/PqFCe
LEs1i60uk0uH4OYY675B6ohkvnkHDFSX8ASl2RemjHir9c4L3SWt+nUpEHcLnw3/
oi6k1lNUlyBKUU8OJwNgB2xNd0JBxFoBZSJM/0AK+C+IkmJoSOHcqx3z9HmFuH6V
zfIuDbxAUZYHtLdyjMlBJgwFyarWtmSc3V4xcj8VYQBf89lg/1QTKPYIkbDn+GVw
noZeA1SLiYok2SG8HVTcSG1KqHcI3ksKspvV/bF8ofglIEpOnUwnJCdXgQ8JHPFA
o5xmtUKFFuwicS9tlzedgiAl04Gc8XwGDcN3TsJ2/wvXi0qYnI91chBse/pRGMnf
PDTgi0r1fUJPwUGqPOfAg8dlYp5VPlyh8UR7RpN8wLFrtKNZpyJUbQ/j3jKnwW3c
6ayDbu3ySG6gHxJHec9qD60QwNE89kjUFDlzipuD95UytHUIBq98lNrBl/pKbY/b
Yb1f483iXOdC4Gp0LjgfmEzHhGq6/afeoozDJtT8NffrE1vxJQaDAx8aDU3BDMNw
unLj+CsSOS4hQJRsTeK2HzGDBNmKkSZu/Gwf85sO3A94kCgOJJFOjyCKQK60V/om
UBWwBZdAoOPcJOjbOy7TYCFvR5UofOIz2Dg+LKFR7bxihfO3PEjbs30w1RK1+NV/
QJ0Ry1EVrsBzCqR6sQY8zsfnlBIaSNXKf2Cb/gpzRagKdA2Mbk1f+6dxDk3mdxei
Cc5OrP8X6JQ6I0IkiAwsms/4t3sZ7P06SR/hyEJX47jVd3FpS6H71Px+ffLztmgQ
H5dEaQ51fzHQcAQM3ujzAyQNRTOUnrXRHb1Dm4Jb8StpFhxBcOpSeWqFpmEKTdZh
sm6dbiAYahy/LJetBm4U6JZ3gSfNcoCPvR3brJcWVu083uNyGLYuYgDYNbYt47ZW
KjEiKkpR4DFaC6LZUhlIYZrNZ9LsJhxy6rO7LAV1p6//LNOCz0p0SrD6W+yjN8B4
6f+qMWqncTvwSp/thild6X3op+UETG3U9xtVP+G+Fqp/T4X10DMUMCcA46ySCdF+
hJtRz2MtryIy4pnJBdLukLb1Hn3zpe4P2x9FyNKtN9lGYolDyaEE34wNWMAB3LPe
ad+TGurTN35ryWmjoTvpEAp96wx4tgQVEdWOIvBtClZ7B2knL/ukNu+zjxAii7CE
SuBR1KLRiOQvKvlfjc5rYaX2GZgk4fbnZ1qO9GTHiLO2OjMoiTjIGa3pe/bEbes8
2XfqECr48Inr4sp9Vo3AE52IHvnHaHAYGk6Xxg47ONVLgmsUYyIUbwlvRIxIr6/0
lJKJaajGDGCIOcG5ZC+pWGBRWN9XrEK82syrMCok1og=
`protect END_PROTECTED
