`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JjNtPAXrtj8y7fcoDFzMGVc2T8hywNJoYSuHVo1miWCLG7c/QpvhrWD78kbwQw3X
L1r1LSXuwtX3rZyNo7VVSYQ5tiYuFi5W8XAaf1v4OU2SpX/nZFbroWPU3FXjcae7
pk+84GcrCDCqV4CSYS0ZZSuN15t5XBe7ZornONcPdP04bpDsWi9Pny1IDSupxnfG
MTbp4ru4FDgNQO0XNVgBjKzpo75exi5aSLmh34l1Qc5p6BgnB/VV1uJawKIVam2o
+7AkIVQBp4WtivjMhSrZVZVfdow8daVNk9wr3hiecBLHQ4tYWKwIs8ojsI0jqsyC
lfTMzvumAuRkwUnAxGGitKpGWRfAZ/oC2vGPuw8jyTCvqgZbNVSfAyWY65JogbYy
JK1N6qVkXuU9sEz62CyO3wlLKhF/Ku19iRVnxkTu8Qrb6gvD0IVJeiJfzEST85vx
so1b2ZSxGGCAxNRmKjC0XCfJ/g/PESQXaeY0bLf3k1LuZ0C1jMC5ukusOOAsMm/g
eUZudT4FHAILoTC7BzrRH871IgeNwg7U2cwPJA7vPK31E5e3QHrZjhVSdb+QXbsv
xbPW9y7GyRdAo0M5O/J+Hq3/zvcDnnb/3cS2Ddx8Jqd4f5a1NEql8P7+c4rrDhua
wCFXr4DmPQiMVJkUTvL3Ds9KUdFpO/QZ1WK37Ly5TkpLTQP8h6Hh1rmPwY2qY9bA
XuJeFfnuceHPStEYTC6eoEKRqjCivqkHF4xE0lhmPTyruu8BUtvb/xFEEuPT33u0
DpQqIrVixmsH2MFpduO8H0oKRXexuSx8xybpSxMgwmS2hMWB/Soum5WLkSZ/fyYC
ZposYT7eKX08OExfCzBzZAEFfnDCcLntUYRB+Q/3wEskVGBZI9xVDZI+ZlqaEyei
EaLOrXCRg8kvDlFV0NWjzGy8V89FMCzOOz7b1zBn2JDZevNCWdw0NWSzgknZAxCY
QHin9J4pByNzdiEzY2fL73nsq0hUJoDmiC18E7DuQDanTDlXqAYP1HzxYBODHiRC
GbGPv1BhaCoLHncpOGCccoVS1kytf8cMSaw8t0FKauc5vX+evtup0Uyqxq8N3U15
PLqo0Fy8b+NVVunEfYC7bnlsC95DOSfeO6i4IimGWyYUcSC2vjNwwZ4al3GC20gY
9uwXbapO04wF188uUK0izxElyKJCgSHHkK4JYSaN9F4loWYBtwLrB8wbXJZIp2+Q
yRO5UbQOCTBc0G8hQpxAWSLOvX38018Ok5Xzq20a2YHODAF4CKWvwvJDg3IIMpel
sHS4FF6dFwpFvjBYnM+3N218Sx0SN98AHIcXa6ZMwNcM6lpqBnGDgX/5U9PDxt/b
w4fjZJ1FHVTbgY92n5MYKbfs3M9YRYcdWMNvPiPb+wrhn5KS+Ues8V5I2JZLgy8d
tqsXJ1o2wAAdqdTgxRFFYjyq7vlgXwKWHF4+W4FWhfdXDygew6kmypCRYqF4Xbd+
SVJNSisaFQwl1LBOOI932dyOkvFFU+emq9A/aHiL/my6wNkKPFZqCYjyn7pNGQo5
0t1HEQ5Z0yXBfgE9rkrN3xySnldSVnXUuFjTt17VNAtxicg5BpHHCOHt3+HJ90yc
TVVVIbZ43V3SBaxX5O6vqS9Gi3PQLceNyh6b/tP73lHDDuIo0o9a8Afwx8svNYpQ
4GyQoHZlzYVqFMrkEQEpcFlEzaIlA9uF+1pR8fNbV2uf6q+prntD/BX9aKI3p0/C
iQzCrrzCT6SYZuyQAEm1DYhasSBpRQEKWvL8nh9n+nGkCKle+nsiEbRtnbDrnom3
+7/PdMR1Q+8m7jLwbfRs6vvfWtLaNUlyDSjkCvcw11mkDGBCJ6TYtg8G43xWkKRP
+dKGInWonGl1Phw93cPNoT8/h98y1QR8+veB8/wFAVLWXYD3ZOjegBcHYxMviMM2
dtuX1nsvpkBvhq23hWGZ/Az8uSY1D/z7Y8qYxgbFB7HlagY4/BaPqXfkUZ543CCw
F2Ym1cSH9Cn7VHkOLJviSEkv4b6nEcFnWTYdgTjLQBCVRdi64iyEwC2l/4p+cUWk
IqImwJV6tUhDEzuqSl1YWoQxvAI3VV16eKFpa08aKQkFXZ1jziCJXmhTaAYzvwTw
Y6MzNzEQ4MXiXypGdF/8Jo4IOtF8ATzXa4yEM7vdkImjeufN613dnlgjWA61ckfg
AKNi4qZEienRsZLffEYoPaouHjL/dP5+s7V54/l41yFI2/pcvQsQlzrK9nWaoUVO
OIj1CNf1k5S6eaKyBBII3i8aHAFE1VMprOB8mUKkuH3jkZA7V4DAZno6QqGfL43R
gsWAb5dSwnoELNvjP4EH+MmtUvJcMukYZBpeR8l+Kpji4hLnY8yb9ENmsLIU4hAO
6/0ZptEdp6+/WOiTUAXw9AeqlgqJqkxYMj980+68ea4ZDrxO51dEaFWOPms2ykgP
RCSLKjG1DmvDkP/4Wlc10+1lj3ZoA6f3hx8qnHlLUgwgoRyaIXUqkfldmG6oCb1j
ulUJgg6+lJa6FSxW9ZDXjtOSPtiv1UVyTit4qILtTNynjMw8WEixOlBoVNiXgFqz
1xgsPBYWPp2EVfZfFNq3IHWLnuPjXsWWPvLSr2hVxIdv/KQO1mmYqAlGm+2EgjwH
z4NiTDhRG/K6wFXL6Br2qfv3kY8oTN1ioiYEP0jJNcClVf+WtIHmLEBeiRr5fKmy
0kKcKfAni+T439j4M9sMFlBUh+Ijgbh09vC4Qq2k1sj34Dr2HXhIIJEyjhA6dYsZ
bze6hJP1gD0lnV/xrxQRAYm4kx9mrurcTG/zlHf0JU0IClZ/YKfeG7CxbIf6AHjr
0mMxadx8IrNHJALWy5uN9qwRqBHN9IKBGnjHkL+2zI2zfUhAbUVtSU3eDsPw/nFO
IzMJtHH/dkwYBCbBoP1xCiLghS6QPmMzE0T1pu1fY0T38JYv88MFPaHjJPgu7ECn
HWoDlU8PBewcaQklhMxtmGDa6mJ4FX+Xdeha2b5/n/WiVGZNOhqHC/N9GvvM52D9
NN/qK5AB/iSmlkv5yypRgwqD8vfzVmvuFfo7/Wjo6iDlV99ri7op+1vhtLIFxHuR
08AFm4CzzGcRKOD2MILfRdNLkkPZ287FOJr7xEM8/am2745d7ifU+YQJyyHlvzia
vwM1azt7iqf5r7YblsrNOZKJUc13sx8wI0g3vc2PyQyYgg//2uJkMOQkxTv2JAhh
qQIhQsrmKWxvVyDSSfOBCderaGsYHMkUA88tqwyR3mGiWj/mwFqIr2pYbeTXt8mG
YzR+w0StvtAyzCBzgZh/OQ8IOBJ772MIvoGqONrG1q4csL+Kf2Q9pnZJPR26V0lt
fOi62Oz1B9ytwUdUlmXk+xeLSkooI9WBQ8ZUwN6PR7H4bLXS4sxxARv1c6YfpWnx
0A5ioTrmemoZCO1mYYCa7w4NY8Xw7jHBL4T0Q/w1Iek3BjYzXWxvqXV6R0irYutC
w+QiQlJTnQPLP8c7O2Up55+MCY8AfPFn5/a7qbNK2zKtXyNvcSPFcWH34sUEEZHG
zbrPQsBky0zjASo+ZMMUja72DXf1j8Atcl8cNsSW4cwD8SEpSK4oJY361gMy7v4p
Rwv44zyKugFn4rjKu6Mqs7Oid4Z4gGk45HUn0DzKr+dnPQ2afaJN9l0bpGVddyoU
uLk4NtcGLsYgA7cWBF4gxe9x5fd/u5JkJTl94/e/dosDNF098Hm1+pUndRT4GDxN
91sUvrHTasZa7LAgZ+DgaKl4VTaaeOs+5horf+JNeXZ5eQCHuQxx6MHin8JXWjaj
v6GRX0ceAuGJuFuP3/Po1aCdG+giMyMmFlmci4Y+2MHBcrTgZ3J1+wJ6OzQR7wff
9cYFt5qt/fU4Te+TD/RKOF+pJuV2tq8LaNocRbdHZbfpj5foPoAOq7/CWGgwzwbQ
ChSDDr3sadkvf9CPxtuAqxjjpUP/TC36sF9xb9nfL0dupJtTSylsgrUr2oxYljE+
qFTrmfEnlv+N5JJYzsR7BRpMjuWWKyAvm4woXqC5PD7A6uuQeyVAycrNEIhjPaLk
LWXctS4z7hrVzXruBysQFdcX2u1Zlg5gNmbJVSIecINLU/jzajuMSOi3HGyL0zRu
J/7tFNQqLO/KAF+2/r73E77+VB61bBAdlQ6JGZfMqUrLzf4KRy0Eh3NtMzsf66YT
jaCvRGl/q0y2Kit5mxIFCQAbATjrDkxvGsw31XTvrfUJjhqguYKDr+cXJTbS76vz
2Ur/mfJt8WVy28WIWwVLlP1IS3k6V4Jfw4sjSgEJ3KAbLFlSyLudvzqGzzgaEFrv
z8VgT8TO0c13Ke9I8qP46tSqHi0h8jHWAdRKsKPYK+OxXBx8YeC1js6OFxJuYiW9
IFqk3W08Mulm1hZl4IMMGZvGfoy9xWWKQwsOxK30K92ZvexpJrMKslpn6lLIyqIP
4BVkiN9SMgk0DlTZFq3Km26nLe0XEtYX52S5QW2CjN7/lTiHF545/VstKYm2GumQ
fMzMEVf9wZLA8oeCO/ptMPEEZL8PFgA1fvDlLplX3Z2X0CB9S7Y27N3JGODmm2hZ
Ez28kqajW6lVynm/02SBbW64b+gbcHi0vmyoECpbQaclbNkr4w2B3BQtlVlc1++p
O720Z60FECV/MCs37SOv+mJ5eAzdv1+IoYKhu5dq9t4p+5s+0fp6TZKV9Bvlunnk
C90pGEqJbwmvEqhUrV9RTH7mggWbPWG+lTxIdRoWM8fPx0kyBFtvJsP/qSenhMIP
rb8cUJFAiAOFCl0rFgn1J0wLvllH2DMKk4CZmvJuAu6UJtFJyor83FPDDa4fPfXx
m3JbfmoL6mQObtFW/xUjwS1SYTJYreauJKVganbApHlyDao7jUz9ibbYnoZW3m6m
n2kLbqr+DrAVk6o6avvAborZwcKmeF9w2w6A1WPnUS2hWT+rknQdFpeolPmgNTUz
7OXfMsg4EQSf+vhI0Sc9MMOt5RQwgzgiJm7McRMkUx/kCSB22zK1rclNtYw6T4MB
Sjej0RIs957owMp/ct19/hg7wwEPQour3TT19hcI5KF6oW4hwtc8MuCuv+cVW3e9
Jq8FlKbyqjR71o3RdyIq0JswBYAZ0anP2dKT3CRzKgaMEMCFBJE9FGkepAKyq0xC
CH28RAq178pKu36W8DoJrBTJ2bPYLf81qWslk49QwtuxNh4Ipas7qmCZ6TFXIp/d
0TUl+jAp0+d0tFGUUkycPgBKa+q2Zoir3m6TUBUXiwF0S8gS8J1ep8LU6pXWtS5Q
8e/gKUHt5PPJ99rgxYubKfr/3/GKKAo2NyNuvudtHnw1zgXhy+cC5kmERymEd2ur
C8TmPdzpiH40B3OaGtnQS7tIaJNuJyAvv4tyqeWg7CX3v8hcp1+a2ICgXGl3diQU
tcGHG08Ehin6UTLZV1VeYaXpFRhl4c/iVROMzOWHHznydHu8nDxybJsJTCFaXoW/
YRAiFtx5DYJLEeskucG+lFRlPm57+M5jt53OR1FnRO3eKLSx0vXf8t0bii5wrzEb
oU7ZfcRE0+IJ3k/K3ylfqydGPEOrwZBiGMKXxpMwgyG3YYDjzqVcQrkT4ekeXGlv
RVwufb9zv1u0KzmuAd1Sqq5hHrtuRqsET8pkFK4eURM/i3tl5dyQ668xhZD7kFj5
8kIv197MgcDvN4n0te83+n7rxmfdd6ny24edtUsIvX4KqdR9qr5ON/AQ5I0BnM6k
ZWItwYFAKgjwws5WJMXBr4DQs4Wh479HOk+JK3K1Ui3yBA6POasrl8u+7DMbwt8+
dj95eUr6WVx1ryd977Jgz2hDWxvqNMVYe8p61KMr8GQb5LhWj8xAcuUNyrUB6/JY
p8qKsOakC1qwqVlmXsxEH0OifzVdmYVz0aF7zhP1k+KfCulRpROvhPeIL5UjgWj5
Fb2CdRRm4kW9f0qNPDmvr5YnUAiApijelONe1UFFW0706kYgwdHay6XGR+AN22iH
8F5Fi9jHorl/L9IVVFLkbEceFnfdDOcn4hkXx7AFTtyN6OoQ+cT51RvqWBD9An6B
AIwi0sOJ+5I2CHsqTC2SaLmBSpqDRXyhDvnZICjB9R9vTLT3ahcbcP1nHZ4kDGe3
61ATB1vFSyJlx5Lh0Fm+zLDam5ZKuaL/nlrpgXUyzNix7yjr98T3reRYM/ME1KDs
HUqdDVoHc9Kk0cFjTm7QgROIODz+cWVWVLkbxqOjVfCCaKsFMa23lg9ZTiE01hZa
ZRE7u7TzRWTvx7pkcrOF6mIyPygTfcqpduk5b/9G9SmDtMCEsB9l5qZlapR1OXDF
sWEgCZFE0P2nI6tb4cao4N7Nvl4fwdIOEtcwx/UU8XTNfB4ASY65EG6TABOjjvQY
P79+d5hQ8k9O8PyZH3jgsffMww7ZYpiPKR9Dr4hKR4u3qPidUjUqaMBD/aNcD+87
f9PWv81S+mUDcKC53BbGi4cG5y/YwKJ+hzKBY+TtUvO8hRDUE1X4trN9qWNX0W4F
mb8eHeCRFQWP2CrCSwj+6GSyTVBJZgSnYtaR6VjKQyvmO5XXMYR6L7kVf5YO4itX
/AmRlEOoRyCLc7eLWFNDkMcMzBdeNfSYav9DKR44keWB6hvRrZ0YckfsMb0+BtPP
Z2615zyOKHhZOY2ZupLwy4abUrAumI6n9R3ZnDns09VKFH8jqDjxbFz8c8WTEdTQ
NmvOSyIBggf24d3VCjOMiE2IpYmgfbzjOMDovI7Y2ra8Ttqfmh3AVVIgU7Sg+Knb
lplrsZ4s4F6I1i2V+TlchgskaOgmMFurUx1rVa8iltwIgzkZLgv6sfERV1xibeGF
TPpkiAT+T+5up6ibd1NDdPWUAYfaMNHFDEVUrMAN89JKqUDO0HQ1RsdaQjQlOK8z
VEcp1d8jBdWWDjgJIjAb4yHyW0GI4zFyh/knneZV4fTIyQ0eMDeTnd+E8/dnAxSs
AQtoSgw1t4Viv/WyIwAA2DosObKoQSwpelISzqxu/pnpNnZcnVmocUGYzoO3y/ZA
6LxatfQ4jTRNgEKKoGsc260SCixRZHDUCmyT1ivgObp5pu7vf2ApucfJYsGSuKI0
1nIq+3k8Ot6GagD+Dvw76Ku6cTlyyAAoontTq5rEEVdM52/U191Oy6AJbfLM2Rjz
ASG21ZZpJaC9cASM1nCnbYix2YDoyuIY1pSEthPfMyAo/3BYdXp7QZJF5jlVSOEY
Q6dmEYY5yuBsnh6NSxwG3qJZbzlczEGX5nJTBgeazm5Pt4L1Uh9+YFkWhojHZ0wP
FiNG/9+Skl1Ei2rj9oV8ORAV+IjBt/h5COw7Xo6wVrDgn+RwGYH8lH8VZa62xOAW
OJNuRaqypUpFOT6MflfjvopSWzr/7oGpbFeB5koCpRdAgT3+wlUODB3u37iqnr0b
AVhQ8riLHE55K+ke6B5Qqaz1EG1j/9oCSMBnGKE2eBiiO3Peyp+UeGMKTPaECbxG
TaXfWi6N3jOhcmy3jK1ncKZnen9+lv4Iyczo0aGYtVdfCxJPDqcrKCZcGqPN9eXc
XMq1glYwkpZZqrkMFXq5ZLf6ClIp8IlWhFyOnP71WT6Pu77Ef+M6ernkFKDdpEDk
VfHwFZ0Px1ZoQu5chqU6nh+xypX/DgD3JoBQ6iVW/l58/oD6p5o8wjyPsYCLD0B7
ZcfOoMtka6klqX8kID4c+9w4gXSMbxvMgekbr0bAc+s83W8ncJoj7Zafmnv51tes
tF1rgQ/uCY6RicbuQItYg2SY89+O6IVmDzlcgPfOFzHpzX/fe/yTnzwxY/r01xlT
7dsswO4TKMiS/Td5n7TlPTFGMlEHcV8vt7nZSEteatGwBOR/65HBVarKW22rTke/
2u5U+AbPpHDhEZwgQftA6YZ9bWBOVOLRK/1aqzV+f3Hp3G0NjzOLQUmPBKvwuKOi
DaC1N5wFRgiPf2rUVFOw4evq/+qySd+lfux4yh7pRqsrmnq1sPto3p7WlPK7gBju
L/Z/b4yewxLZJBPIIwfAzOfHD5UKxbNf5kWP4M0lah5Ep6AOdq3zbbnHD0najBVJ
js/sOgNZvsNsRizFgawNRKq8MjnffmUiM2Ed7ecsG7RcCONDW6PkyJxXRWtkFfSY
TtluHMplr09Fp3EXsAbPe2SA7D11RvLtlxHgpIw5XX7Lnz03oK56DUA0FISUXes1
CYQWolMOThvapbGUCvTs/suutlvZn3OvqEFX7rLqDW4Z6ktdo7SDc7WazW2EXvFX
DoDY2kiVsGt0DwBmm1iUlNQXeVZHIqX9qkdAMsSXD1/4thXUZ/XROSHek4mh/neB
J0kaRVWGjG8Ly6B2KtIBNY3dElG0s/vSRuCr2oAaVDCUL4ZjhWBIp/yed8TtpJeY
PmWIKh4KTXjXp8M+rEA9F8pl0unf8b/hA3Jyc/+vwaoWWqEDAr5XHzwf8yftM0wP
Lh6RUzu+fqhGDhIi0qaQ6KgGjV3d55rdhLihc/bSj0OFwLBixSMbM7ZvScIlDZUv
rX2rLs0mJuEnKVoAngu5Qz9DrjrmJkD85eRRJcVxnZBl9BWRsfHeYlQ79DmE97xi
LOYwu4W8ZZNAkmeiG0+NdSDLwqABQn8ixbaYCSNHZPSvvA1TxOXzVxe6EySuZdZ1
wNqGhYJe9/b5FzxovGwILBfB/S+W0MO4RnCV7bmAsq4MQZZpiy0LWq5r/O5Qkigg
bvAQhYU+92vx+Cxr384dddtL/334I/32s4ouOvK7ox5VHRgh8tHZvTs23oKbhJDz
dobHm0zx/ZDmzlg0a+JsQ4SV15DshLkOVl6Uu8x2MWTyEAVk03kUn9kR/2Hc3VOB
srCO1njA9Tkdd+ev2CZ+LVfMGTy6gXzZY6w4x3V7SfP/11mT2b1u1tszWgeX++gN
FKz1dTZaL0jq/Q93b+yIe40EB1bzsySXQ2/mfRoyQzOcvcVstnT/EFn8x7arGH6S
1sOjYXnsvnwArtuZzuINFjxQo7OSVfZXF+KJSD/5Vjkz3tRDiTwo/a3j4KUfls07
Ys98Zzh1qhEq8WMqtIK0+toMU9u2OT3RYCuveOJ2ID+6UZsUP7tnE3TicKJ+IIhh
Qgt+geixrekjRf2MO4RxWbMJL6TRpTk8Wm4zoQvk8lOo5Hhymj31oswAlRy/0SrF
He9M765+UW86LwGrvTODns0/pCsM2fDq8J7BQHR97ldvORupaLazLjZ7b66qfzn+
/467x6bi/iPG9ngUPuNR5/jgc95tJGzmncqnlDA+RRcHduiMp7yOAZDn6p0PDEYa
YILNzymDTYEoQBMd5c/ppnW1InzVu8p6W5ZWmsa2lazUDCGnCD5OX501njpOioLN
n/wMwudDwB8VxRLrFDBDEeRQ59takr1hOcHAD7t8wJjjU9NNJ2h6i8oPX85ah2D8
yclBmL9TuHQw8EsFi6/5vEHr5JfJck/Svabzs+nuZKPPHNhITAPGNdrqbpdr8xxr
bC7oc03maTXVO01powVEQC/eGzumLiZtVnoMiOncX+scCS6LCvkknVMrMlAMz/lM
7QElEGPrL5GL3EsxiDdQV7j0NxROn9Ug8X9F77Y0bszKeiCKSSRnfyXxgmTdsDZr
ufEMBVaFC7evp7CQ9KZ8bbxjR72G8YCXrvp8oZY7/tF0PGJpUPOFtPTb9F/kXmVZ
Ip5zFd6eNAgBXq4kMElYVmLzFyM3I89SR6BkPdCaQ0vAEjGjmoKpXil29i0iVefF
K0TYXRZSj4uP06LqibTsc3d9l06S08GNaDmAJawaWBCTPNR6FaAbYw321fauTTyc
R6H3vVicSViZVsvsBDBsBiSnwQb5T/vK8hdekRjc/Par8xHJ/dCe3C22OQA3k4Ip
0+BJZauj07e1jLPzzY8drXCc4/H/2W1FxgHrsCr8H1InT1XNPML0CjcgwoQsn5Xu
IEiP7R6CXQFWUDg5Zw+LafLbwMnQIOH+rbHriJeq017xsRFiYD+H1EMP0ZwDncBl
ai1oUd8kjxrzxKNCmu8kMwKYIk45y/5yuL7SipwsI+QMPTTyDV95WuSLm/KU3pat
jjipKMqgl+qXbECib0/0igO1z/oqaVYwmsr25XRDuHZLt8WpqExZnofy44ahJRCk
Gp0fMnpjT07qenb/flAupgCZz5ZAj8Vp0YaGWNLnJncV4hdWFzG4nH5T6pWrqfUJ
uTsd5l5Mr12JaC5ej4iDWoeIzk9iqoMdN8C9TyJEH31jMgU4eKbh+KI/uS+VLFhV
jAVC2rKBkz913Pb4yk6OJipp1OtIjdSeAQ6/YMwMPsw5xhda8gG4JgD1ONNIMwDH
U04F+q6uJuhTlSaFMhP2Szv+ijPPW2UENptPFfahy5bA9rmf38OuP7VfgXTqQCks
9iZQOaspZwaJnKdBgscNTVODWFjNdgm9konNbjQx6l6HoVSnf9jPknh9SLKJ3Jiz
Apogvx1uy2RKgHB29AokeOJ3epo+dsqpJ4hfltglQ1pGafO3tIG4vuBUWadnxOR1
sVLdg0+F+gWNE99Bhe7yQtumcHTvUdZ7HqaRX+9dKzuGrs8t6ArKHL2NuJeai0g5
bWn4X/gyYyE49uxrQVVOI8OKDR3pJ0lzyFcDHoS0Wb1IrW+Kw8dWQWMr3PFJNjdj
UByHZn5WDPUlEVpDqugJDbayU0l+YMsmt+cPxCHN3eEiZt5QKC3AbM4yYbLv88HS
XcoR1jAPMqiL0vdub+KmA0Hf9CDKcvJAq52vdkj/D9FSSJ5jA/kLUVWSjwvtSWtn
1AVzD0R9bS6uOnzW4U1oqvUFJH6B5NOmBtlCs8YbKhUqYPMXxqPNIZE+J7LHnIl3
GpCDx+VKBWSJ/UBwpOfs4UGmIozdR5v51O0/8pUivgu1yaT4I5kzYxnehapPl3us
GeC8hpC+0qMDwEjERFi56NrCjzXyJK8eBCgCosJObhvh6eCt0z0BpCkzu0ykds8p
0WvHUmyTBcnWSPO3SJX7O83T5dAPzQpZQvQQWUuO1PGACfK2wGNDHOvCUhOXdiKw
G3q0fX9AszXcFC820kjn/4cmJqsFBynwIj6fULk45ytnn0JtMZPeX7dgzVLV9j7W
oLKo8tbm9lDP+Un52sTVq1sMddhdCS8+gOyRkiX5OnsIQJHyiilfgB3YXMqIsJCr
34mp//V5JeNyR0h2y8Ce5KNdkL57CVOXLhGo9dySnMf4LZFSzF3+Tujx94IHb+t3
lgVK+fYJYdix72tPrvsVmMxzofd2q3667GaBRDnAWn500cUANvx3AJd/rjJ53NA8
AfYU6Bcy2HpLnRPGooDgl9sjXD/+lUAngACK6Z5fP7A1qPPjBwQNJe9LK4eVdEn3
H8D3Qv6ghHbJ8P5iHmgyCMHNsOvYuLK4zveigLpBd8+dh5lpB/WIlTMRektvEkJ1
pcfmkTAKuXSXQGmx6b/Yuaah+TQLomd4xJ367Wq7Sm7LlYRyjTtCXKuNE6bfJ4rF
Y8UlOKqDYQBoQmr/2m3NI2rS62pD/59T1+EU61mJiHBgbZJmMb6RZtQTUIJpCkbf
N2Pqh3PnsCZUCcvmcpR2XtiuhMSQCvuMYzQtdi4frKNjdbJxWq5fSOTe96szJRTC
V4pNM+gbpymrNgvMBccRVq6PZRU22HqCySTmxE68QFfqJRC2DlwKzhdVn7rNfsvV
2JIRdUPYm1yp2V5dsB1bOggKBo2o+3CpSb0AEvBGrV3E2rHrUJWfbVIKBNRmBVCl
lDvGiGAVIuJpzswKsnOp2Ph2BZCi0hq0NKwaoQH3dbwnZHU28cyN1pQiFPpBoE/H
/5ggeFbu8rf+oY92Vn7oYQCr1qQN4Hjd6qRgocUZ4rbxmAxUvCwP0CtIgmuYh+jx
DJ5V8PrzS5QzFH1DuP/t06pk6uf092SASlhNNNkBCij/2U1n4RXSkkekXUTyC1rP
aCPFVJFBAuSge5r9+SVNR148NRx081emIJzAQ69E+dS313j9TKMBeqsfjgg05bna
XoMmKmgBQrs+zuOjZ2KXJL41mXvJ5MZ4vbOWEtCsmXetrm5rxIgFtn9cXyicJZi/
IAraTyjixDkIYDxpir4rpktwdN0yiws75w3+ocA1AxHKPfyBDE/Q8/LS4b346OL7
QsXizKLLdY2j/+p20DNIVd5Mb9mcm/IT9OIHqvrA912x2yQ5sZ5+GBs4kCq8RXY6
JFRrilCuEYVp3pYcyPXLBnhjIdR4u3wsFJUr71xsEXIbV7edn7lmRTv1bpzx8D/q
7OMkRQ7KooAf82+F3yNfZTwCYxtmUA7HN1xbnBOti8QANNNXQkw6aB7OZLszFtli
R8RyssswstEGGnMmLgflpMLszzUc2CION1l+gr3FFNSgM8omGrD2h5S2EureWREo
Esu+chvqsS6J65NP4k5KpSzhRbGV9qVZ4gWpCbXrnW7z7E4if9uKZMPN2NC83mzU
m44yW7qa9D3qmaPgpf0rSc6C3q3vLImSQqMfhzK3W853Zcy2l5Y+mmHhNUpA8Eat
BMlrP3HsSGu+GLtwGu8g3YQ0GdIVjTYiURpk8DoDWe/eTwVeAIsSqHDYhl676yN1
z/rG1qtcGqg9AHTZF2esVuVLnREN40KfMBgRzAjNXbfA9ChWDCiYEgCAw4u022JU
OQ3SWDpiOvFT+PUeR5onz2n6YCvw0rvFpNA7cNk2KEHrm/HcS/4IjjviDrb1yXY1
W80R6okQeXYeAboo0M5FBS1DhvQ7Ypj9hpmsmS2PjECo7NGLVEpVzVsR0+ELoRRX
kRxJSaN75Z51KEJdCvBWu0r3iqLQ3H0lz0LmsviUxRZpUSwl0Sa4yMazzt7zSX93
TMS0oWwwE4UcvUMkMl9vSzEok4hsC72R7yj29RdFPbK8Onlcj265zxNuX9MPNpFn
XXjk+GMLX7mhPJ3kgJHWdWyvksGINf4spO4/ywHaAvwjaUsgMrbASYj7znMElsaT
nNmsQb2YrEEIjK0MssdOymykQq+ad46dngR1JQ+MV+X4fH7KCO5GMYdYLBtVuCwG
A6t1k49xBgv0reyiIMFpy+BsyxG8c4w1Jfqr2zZ3xjq7pbADiEZx8VnNQsrcs2eh
cykuxKyfoZYhc6cCns4pgi8QXIcALe2Q+s0D5ncraolwEDq+su0voOnjrbEueGh9
lzCW7PuTsYkq7e3I11TTqS8h4LBa0WW4e/1ZJAl1KwNxdeaPRU9XJ5TV4RYolS2y
2HR9tDk6UEn0n2Yl7r6ALrZWwBJ6PtkNrO4U0Q3sMGMDAm/2QsVDm4NJg8xXE09t
PrQJWEDXVuTs0AovXtgpI0Yy3H6p5r9tIgK5CvnaNGfSF7Xatam2bkV+HV1HkIx2
h731BFwjHSaHlUE1QShrrKFKcGPcfdLrsyFt9RVCdNfJr7d7RlrC+NWasAFOAcE+
hlpFawQTtqws/PAWpKgbH1mV3ztsYq1BkNIr54/3HS7H2uyTaC7CxqWLX5wtuliA
2DESCzQZ7bQht7FW7iqdEGb8lOIF3MiTz0IpGba/hU8JJ3kdDYgIxjo8OY938RyW
7N/IDWDoyGAvGfbp2Q1bCO8g1tb3REMpf/xSpn6xIcWOFcm7Bpw6KzYFlLY3/sdk
h0DzjRuESJ+Ux6jMfy4EBeEqiKjr1r9YsYq3tU5s91JEHPlPSMnBWRXT9CDLLpJ9
qcW3thcO2j8mBop6mXcj4bEvmljgNJo9IbA5VWUxBXMNth+LRqy50eR+aA9vzgWh
1Bcjkz87JSdgDt2KXpR9cBcyc72sqR2rLyT2vmMkiNEidbYVSETzO6deDwbNGqlI
JK/N5VMW5SCZZ1HP6ThXuAUDVTSn7Ab6oHdk+XjDL+3DlJRuTEaWgCigbgjBRYHT
3//AlPj6E8NP7HiYRuuz1H9UUcQDZHI7K2WxP1Fs2LbH2pVfeVgJ9rN4tM0zcwC2
9+IBYmry6JPSutMhw20CS9orKLVuQgJ5aAxqUpLFmDFWXQrDhmCpOgXKVw6I6C3u
q7/nt0OH6O8SWHiL2XCBYcP2nF+tZZh5jfas+k+JeN1b56vIfZT5Dyxb1WS3gW94
pHvLLn6QBPOdfLJhgIga8yj3ulOLKkJCRLO0CDf/wolvtamPysWkLpT0Xh0HeUjR
WZyvONxncctF7YTjwzUSpAanJuJiFoce0ngvfuYcSLYFMq1C0GtDU6BRPzCtysEp
AIz8T6K02XKCU8H7atWhSJxXEO9ZeB646ebESXh+tC8lUSrcjxP+Syrd44EfZJ2R
BIA0cBLMTBny5o9sEFup5pDl0VHSbSbH1SJyGNtmgTMpkNpd/EokotmDIKJnMCNG
zurdxzgNXeEvGBNA96/dXBys4n9TP2MvmkfAnCX/lGaVtPWJkLViNFOYrz2uL2d6
bRvNMBwLppobxsSnREq9wYTYxv+9nRE4/YVpe1COBXn76WK7nGZa/q90P4Nv1tgD
oZGOSXQdaLyd0Z7X4wpXziWU3Q1pC36gdlRFXCOzBWZrGcC7Xf+ccf9JMAMCRjWk
DAb9Xo2AIHbKJcscyky/GMJSYO00fcWcocMYLOIQVrNX8qj7xSZ5vysfZgOfGmBz
bURlKRGOAlYGMis7k3hosVccLweQY+kO4TeKNiaZNQ3OHCK14t/QVtf+ocYnynZc
46VZQOKCftlQpKVEX8PR63g+8tLGhbI3rLyL6rslYVmYoG+tSm3SQgDFI08UA7Fu
zeZFBLOLNbL9iH+UcVaDDj/ZmlrS9dd/ty48aOF6sqhx2IUh75SS6OPXiIVClwBQ
BP9nzTO86FJycgccKVBiLm0LWPofRxg/OHb0dcXXc+36850/M9tSzOmHjhId7BS4
b90dC3mzHKdGZe0f2a1h8fyKB/FsEXOcgtqNTAHzXzCARIEbOoNF4bqNN8cFsgFY
Sd8X8hT9bHCH6tXLcAq45hLeQ9MIbR2xLbLSRkN9nkndzY+wE4o8fsbEpjaNPd1j
jqm23r23Aag8vvcRuZ8c/doHY8hGe29syOKYPt17MmYwV6j+zqDmm7Cdo4SDYSC9
CtehdoMnRZwpa2xgWpXJ9HwU+jVg/zVRxZRKBYNVTqZFLcj3L7/HR3jgTVVX/Dxy
TzCxc119hI4sJ3IeLvLDYeXeseUiD1nPPu4n46Ijxv8HKcejW1BZbOyoYXtwbHWR
eD7AvmvlftUM5OpEvFcTldd75vRbhZ4hkisWa5GoG7UX/ocGYR7Or/scC0bRyJ2P
lewsvX6ITeIBShiVrCTN4DR1bMBHGmXhJDgE3182rS6pNl/nI9mPNSvTNTSGbCAG
T8OLowGCJAWpBN6Pakgbhf+IMl6GZpT4bM+NvX1NRQ0tnwhDqtUhpj8HaeeVRsME
BBXzGyYX0NPL6lYSNqX+i2G/KXbqwsZ3Lt1Ekhsd+Ry5YtrTqQ+KJmVNxqueJuq/
BOTNzKZe8lcfnGfvBfk/Yht88n9Q/CWHuVExIMKGqOrrmSdUl1O/m6KtZKO0++SP
f8fWPXl3h6WhJbp8eaN07jdbQ4aPpvAVOVB20HrscunDnClFC4T9+vZ/bxOC5QWA
2VIf7PuJwFJjH+j853nHwkxZtcY1c32sOuvzfPdwsEl4uKAtIEvX2lJRKiVTL7V3
LA/QqyPrBqbjMR6vpF35TgiFh06KK1YDhJP60YJygzaW0LuyluEwpDrWzBE8jV9g
fHnZXWf6pKNYmXj8BqJY+HkNsnIbIAGjiD0d/vifXGR4Tqfsm7tOcyyzlKKFC+On
ixDr9FTsgG9VEJluhvdnrvxIlWLOxW3OQUxtqBWjbGfkoTaSQO6WFj1nq812hqzD
iks3xFR3lr4Cptbi5eSF26B7YMKcDEFNUo6DCKBcxZzsF8+WjUPxp9b6IpV5waFF
29mIuNb6+lsUC1/rsh+cTlrxz0JJ/Q/EuDaMYUai5jDR1sFBD53MoryCmIT02ot9
atHqiNmdCz2LR5BFR90QbBTtkSDKq1TowWAh0d5YQ56EWFWpVQN/EKAtF5HRX1We
Pj5mnWMFegBBUqtO7xSiyc5hxDfnJA7/dChYXYoKu9KTq0FVe1E/Ljv9nqD8F3fA
w/t+SLOYIAgpJ094q5CrjIXHu6p9IzrDSCPJaf6ZgeRJDBBifgZjJf4uAOWT+Ohy
5jysHJSGvTCV+yyobsjT9EMYCxePFZXu/rRr+N1xKTPZxyuY4QGTjaK8+BJLP8er
p/zjhkzk7uRHGELt0trS31L2aQRoU0EBBiYsNQd1g4gyNfsu/cIEQ6vSvbG/8Mk0
OQYpIoVNmLQ242ffktP7196QRatNdrQ6VL1Nhhn9vrG2jPvvKlUJB2xSnD5yLb3L
GGeK2/LFnE9iFFCh1QKzMmSEErP2fi6Mdk/akTXlHPPVaiTzh+szdEQj/26uXaL6
B+H0ToCEG5LmrVmNtpYMbAeKWszq66GsOIhWzRKU8GbAgFSx0UdJtx3KzAkA0ZRj
/IFbVxHEQtSPGD4LWBbJ7xBOVCjH3FsQSaTbCVPS0O5CIw0wjN3f1hRXqfxEre9t
vxWJkUHJM4NtynXSKKPL/G61mo6ZvxGSHRpGcEQYARifaRLPC7440smrZmi8r1fS
XJcaDxCh76QpWQWewbydJHuL9mslqC644Mj0UfzDBKkgYLcc185z2DQA47DFs8CU
WbSnSaBse7Pm0trA29eHH/QafvYWrjVNGyyJjfGCAtJ3SVho7GEP6MXV0+/s406N
A8KGQEajDuDQnizik9xzOrPLbBAOJP4SjJGwUADUrsD/owfRbYd9w8v31GA7ZzNR
LPIB/DehL6j+WzJz038EEN+ijTllchLFR9THO2c1/nG8MIKRKZHN416ZwHv+LnKy
gn0X4kowaf8aKdhQlyoBVtbX/3TK4Zr+2GtqXl1BgKVDZOHOxV0HqqDtQI4JVDx0
zM0DV1ZxDBQ30t/RvndPWCb3VGvcOeQYhODcFjv/ILoosT/l32lCknzv0ShGNLMw
kp10jHskfuCrKixn5YOMlYUlcgWtYxAZDw4DZ9Yoqve1dEka7SXCKXcJszm4zdt3
m+OA9HznbkGrDBTJaybriykCLxas5oI0DfebHcF4T16E340Zf4JaNwz8WEf+kKPN
ZheYBQYKlzqmTj5b7+8iDSv36NHu+ni7/4BDxZOE9RXLo/hnuMMuLH03ag5ZRFWg
a2oFfP6pxGC3uEVuynOZ0Vq2KCNpRIVfYwvFm+qQSfKSsz6xRamt9niCtxaoQdEB
fJgzb/PQUkEKbts0om+x5sPNlxF5csEkITpvUbEn+rKhLp6ukwiiE4JOr9Nb9OI3
LapvM+gAJeXKm3MENqaxJuxdzq4jAY85uM1lTAonCNq2FkbT8AimJKeFA0o3VrVH
jgNvf4NXRX0HhXYFZ66qLL2+w/Z4wAsjAZ2r/vlRjHL7ywfvrMhvJOogOvsQ5JfR
XDSbfZYIVsJa/yCafDZpTbIHQ1lGTUCeZshjm6Pqd6cpDDne3kaiv9Jp9Sb01JW4
YXeroniyo9dIf7yBcFGIg9Zmft5F5POgb09D6VIqpfGLPZqJ15JC2jsKdctKq9JA
982jKHiK0yE6St20j9YoFSj3Wg91Fj9eeuU0+09lL+XxSRlMpbf8wOFv320kfu0W
1qaGx1DF8DP3QQHC2F6ClU//H3KG/3eyOxqBLzaG9dFBIjyf365uE/q85U/YlRUf
mvbGsxDdTnhYfWZvGDnyuhSSltyQZeVdxnxYSzc94W0WtaJQf0e7+6KhSO4N0zlN
pwh/7j9q68IiFO6PbeOV2SQMpT5ZqgfLwnUExtGbC8YisXmeE/xJRO9JLaAqJV6f
7jndTCL5VriHklmftgAOIcz/MVfaSVUPSXIukPkp/eIdz7X4Q8pNML10aZWfw6Nf
WCSZggsY+y1Ug76l+xOlr59D/snqg0g/aPsozrCecrwWfz1Af4Bbmpgd3RpjuvNs
EyidCT1SN4NYhZTMMU97IsqatA2G2WpPSqhzIgGL3OMoSdS6CyllO7kJ4RVBclNL
2ydQYtFUjteKmbGkKN98i89cNCA5ZgP2LLrfcqHyvUqzts/On2bWFKkyyLJPhm3m
ytJcsXjqU4gxZKZ8gkTXX6hF9UcrLpBUED49ovD9FCO+Qj1xu5Elf2qO5OOqgj0S
3UdteCHE4FFchgSDkk2ksPIm0BsPfsaTZkwGKyS5gPCV2CrPxoRsGQco0puxCoGF
n42bcPfLChSRe4X/RbTDr4qccGVbaabA8wcNGiazV8rXge5VchwCWOg7kAeMmdnf
NsrdK1QlXN6s/ahR+6r6SSk3aZfMmhLpsl8AJMuwxBRaoyV472kEqYcwsxgenUXa
c8vt6/HduyF2k3avvtzAA60XDx1RGJDVybRuydNvbMGXJ7RFyenY1CRGG5sotj4Z
82ZibxWO5LXM7Ik5Kcqzsm0N6YArC4Be86lOFnN1/dWF+uyKA+Q9mMddBssjz1xG
+9TvvwioNX8JjMP5LsLw8Z83GEqR8ZPct6HVw0QnQAkFzWdQoyBypHDFnWYZuVEf
oybto0TMZdIn176jO51O3euVydvbwc2IqmY+r2gqMFMNC3ujVMtsjWC6Ns1qFVze
dTefdn5/SrIRiZAPNx7diDDHdXu0bYodJKvIzfDhJXWZwRFPqX26cn8mAkNlTa7m
AjVnpPu+WhXbsZBAEr5oen7t+Z3CVlpRP63/Bn6/oslAbbzxuAbtixw68bH2C/hq
GaYg3zVRtJDX4IF6Ld0Uc00rOPKXDX8n4xy2N6xclHld1ZEiropjhY6wy/bLcN2J
kyOanmv9+X0/73HtIeSz0dFBa5L90uEp6o0Si/C54TO6w8uJVrXFTyzDrA/dpjlT
kRvWZcCuo2D31dwIlxmTfA==
`protect END_PROTECTED
