`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CoGYxOounXAEMeda3fh9ND3UitbxC57Pz+UvZebYDQ8he6ChK3329g78RwNVrzse
jnhjn7KjMcfb1RhfrD8KAQhDz8+L9UFeOUrL4diqO//POLOP5XjitpKS65Pvi9ms
5jDYKZXP20XpYCDLbY1qq/DqR67nepj4+Sy08QmM4aeVJABZ52eBttdTAwsSu2r2
sd9D4ewuae+KJopXPROS4a6xsO1tjGQsqJ1kTB6BxelMjX8sdhg+Soz40bGUNmNE
3Y6P51I5LN4WQeATgJmQDXu01pB0XhyPlXORn5j8bqkaa/0QcXWXqdWruSURjoKx
o49ikk8kJDyRtSA81YYpRYNjA3eDUCaafUX3Hv8qierSKC7uxyXb7SDR4Qb9P4cd
rGMvA/wLzK5Q+9C/WD6Wn1oBssWPeYp5mF1EC0VuH3DKNITMoVGckCcYcuzem0Rg
+hKxU/h2n/N4TKwfiyqsjx2j6fSS7PU4FULI0xh6xpuJGDyCHElaotpTpqqrxQNJ
QLs/NbpJ9O2g08UfdeDveFwE5kpu/iG0LDSlLLYVVmUssphtjrHgYIF9lWhRB/gP
WdaMPvfGwpVXMGnLAAHyuDtKCeI+o+5+nx1zv9O5Xu2byznSoux+angHz3hbf8Ff
AUwuTHTyXy1DzUIxjNn0k6f4uDliJcLqeipr5h3MNmfcT17uT7S9UlitwArrPDhI
`protect END_PROTECTED
