`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yzxrU493tklx2hrl4s9t+ZDh/Z6f/yBe0tj9qRVzo8DuCEYwTu+X0ksQPCGRR6WL
TqxoVINgCn+arvmx+C6WWrGeIAjhcmkwGUAbRjI+rcKdpG04Xf5NY0Fqb7Gw7Sm6
1UtZQ9/IzqP4PIMms/LHJnk3nn96BDbbWMoZ304PM3cfMZjJ3cjavRpM0C50Q6xz
wPv3VSAJLGxnxJtRvunW+gmzRyPYl4uy0hM1GFuKb41pljN/ZGzEXYhZ7pbhca18
8FYMGswCkrqxVF6zKWJkkq9MDItXisZEA/1fYPrE3m4VDyqDnG+fADR6ScgzHsPO
tmzxx/HSUPFIuN1gqAz5kHwgTcBdfYf9cIewu8tuG9nn2bnpYkGFwjkbS+2VmQvN
T4awZQfQQxmsxBTCVi/SIW/iaeBnbySasW88JHtGXin4F28/zGxPPUenPvabK6WB
9owY5r5DPtkirlD4nqdDP0/Uu8IsyU+ZKDfaAvQKbUTxuooKuWMiySEKqtIFQ84U
cQeXTOl2CggM1lYLrkoLtC1B1I8D8kcPlttTsTA0IG6c2rV5YLjBjnAY3r5C12GZ
s90UpNI+MHZTaPMobnhjiQ==
`protect END_PROTECTED
