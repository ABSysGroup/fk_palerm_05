`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PWeT4unYbDw8Y6211HaIa/py6f4jkDZ8AJaGBCKXgGfn3FY75IaKqIkjBQX94YHr
PJ7420AmX/sii33ksorIscAxeoeL/bcGEq+TXhzcHmMMcypsN161H87fVKWbXvAB
wxM94RGR+EDEXp+2mwR6nQveM6PiAlPdNbUBwJpwyx4K+V5/YsFUH0qL8jA7CaXt
uYnr3fQ5Yla1PE9d2lq9gHfQanrdGRVprBn+jAgYKdT0nyZgTNwfE0yPWYLhtpMf
`protect END_PROTECTED
