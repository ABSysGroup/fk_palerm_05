`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iRH2q5b/O5FqzINZOIITBi5ACUuz7oaYjOuG9d71FqfDS/sbmuHMQFpGel93gOJQ
ejp4WVy8f6g+zyOcx1wDKqc3Uru8soSYAc2LQ8qE/f3LFTjuFGrrKf85tHly88wO
H8Yj+LNhMyqORXqA/3/DtFIcz6yEDysbFbaEu+OoxuAw2p5t4DCGeddNVjEmma8p
ez67zzibr6VfIrZize/QUK6l7jmHk8dQf94xOxv0qp4hNu60JkZ1nrEN9eWsBtkg
fxV1rdrOmaCdbX0E/RX7/zP2Zv41glpPi7/ppBw73S2YGbK46ci89dRhPDF4+JMV
RVeYvHJSHTpg6vqfxC3OH5y6NdBwZSLkDw0UtLCx2M5gHsJLnMvl7oefiSEvr4Fq
`protect END_PROTECTED
