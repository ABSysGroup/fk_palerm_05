`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N4PMKsCB0B1KCJU75WoI4217oGKy/yBY/sz9wlSuRg35uNltKOtYh1zWP9lDtUYy
ePditsSzY8tndSUbBpvOZEyb9b+N3hVJ2tYSD9jaCf4qrQQGA2G/iBjqHsDZ4eGC
0iqgfKA++pizl1cgLSuXGL9/m6I3DAKo+scvMkeKvCv86pWkj+NXcHO3ja8H/kY9
AuYCOXgSLbrOJQ/G1WUmaWAUxWa7WyeIHCCBqY/KHLR+ngAtDUn+TKcYYm+Mfvr2
AUTFhtXRQCWmO7fH+aUdl8bKpH6qKT+ldyF1Vb5dYIg=
`protect END_PROTECTED
