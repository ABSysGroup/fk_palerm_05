`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n1b293Yj3bpWEqyFxlj33rprsPqZ2uDr8PGu8YcdIT2jE7PXM5dZR02pa2yCh6CI
reqakqaHvFQhu3IfvDGz0qLDOtri6sM0qZf2AAN0o/OXdv8lJJcYw/4RLZDtOIT2
hIbBrgmRpk4N4lfsf056zOJPk9ixVBhsKw4VfiUOVV+P69GrKy0v9PkJQLLBRZ30
I9aSRR3O7AGQzhi+TuGmfAmKSKG4wDlYAI2il3ZvH+UGMyTVDJNUVQXIX8huydLQ
ZqJjOwrw/pKWxuTykRvGqKFsKvVYaflD5vLVuaVqrVSzoJ67QesqyG01DWTGPTHS
2tnkFRebW2J0azU00A2Fp9WG9e5bsC0GYfMY0q3d52d9MS28zhnAgbQcAKMhxBBa
mb2ub996dgdbt/dq5h6XGHXQBA3J59UexmBaYOi8cXTEp+9M6CN9DTrFFGWuIoUr
RHD8qPKXbu6FgeARHnGC9kEpcUVheeJWNfmsKv4F7JJVLhZ9aP02OYIf3l4fFunH
vAIBE+tPTKtT1GW11xXLE6MOX2OirIAfDyuyV4RF42qYkmfp2Fji9q0dhphceMHt
GbFlqFobVLpW1VhXUv+bQBUdZTN8vbGCnfF6eW9iZcPQdZk82lG5YAA6w10CSNoO
O/d2qDqlbmXy4OGyUwKqNiWBnze0yxHMSu/95VVQApoYz/tjpa+/SBtkM4/eVQ5j
E7s2ACJzzvFKBfk8zxYY3/UZ/C8xr9TYjdzop6oQ7OC+KkBzKdTNoEZ1dtoH9Cpe
dp+uOoQD2/7pvlI4EhQVDEn6y3zDz6vuS0KdQs5WsFtut8UO46YnobLZHyFJPzYF
QyTX9Adh8g/zO0g4/8oeboZvpCFvMfkxHRnLSCZ1aLwuV6cHbs1cN3NudwNJJtJz
OzcWVj1HEzcqdCKXt3ADY9pgHc6f+/Foh8q8zQmTlE8181G97Y2er5bdDe+8s2MH
`protect END_PROTECTED
