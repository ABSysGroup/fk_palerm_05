`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GI1xkByct36WczO+gD5mzW1ImW8llVLMnHD0Fg1M6T+J14eCb3jTz0ibfGfS9iod
HE0MC1XH8Db5tXI/dzUmg6OWg6UuncssXI3xl2KQPh2DG3El3nHSteB0UVQxVrzt
uaFco0MV4eXAErKSGPbjJTfP8uF8y4z1Bmi8TKevnbPQSM98Dm9zwE+Ie2/VxmcZ
M322vIV2ZIA8SZcU2WO1VFlK+5W3Enq51dmK02di2Lc/NnBsSQz0u4Z3DOBqrrFh
2C/fcdsl43cjtSTibRuInyqf6M7bR0VxRuJ/JnJYhFhFBclCIrIImqQfsgC2m+Yb
bWdHtrNmlfG0sVUdbsJ2yvxi1ZXFlu1yavIs3m+Ab5gNHS8hA1GD9YcNvyRJnzW3
TW8fRYbpUz+kqkNc6z8lEaIKavv8noFsxykhgptoVE3qT87xw9SrmQxqFFV0We0q
/4kVpy05EwZpeboZPyx2sdwvQcylnjOdr41PcTfkWiS8ZT6aANacITkLkCv1Txhf
PLA+4EKiwOv4b/jeAPNy6YUH7RoVl8KlhiJni+7RJK+mO3FO05J/2T9JYH2o6wvR
Lj063p6F0J9Ks8NIN9lRIxsvOdG0Q8HcwMexRZpZAx6b7qBijF5eGU43j1V253dZ
R40WdMILfGxnfF/xJT9uWwdiRVy59HVdPFkG8kU2GbXzm2hdv6Gw+FkfGacXlhwK
xB7P6glJ6EHxgZ3jnyT4NEPLdbhcZ8Yme/HLquiMp8M0NU2Zj5FXYzTJy5At+lnf
bdfUQscaH69G7IUdioIAa4bY1wb7cfaYP3spVePgzsBWVk+iWkwN5LCRaIGJ1h4M
AS+uZdLOPZGASDEW81ROxmvrUwi49qZbfOX+3Wt2A70zJiLw1KYaKjz/Kqh2kr3w
+tg3hr1+/UQwYBZp+mxrwaTZZZRvrxwtaRDGgcVVtVi3iKY94oHyR4vH3+4+SbSn
`protect END_PROTECTED
