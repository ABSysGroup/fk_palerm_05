`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9bVxBqtkr+UdIGXejn2Ak/KJxMXtaFvzZXKyDbPFY1MIOa81KlJppt098Vka48ff
4of44HxuKZgxoOFpJXH0Z8Z7QVUvDweUoSbNOzFNZn8ssfPzNvv0r7fHpU7RSQJu
qkMmExqbAlPNRjzWkjbRFPF7LNoseuizQjbATdVZajfB//JzDcl3QfE/3bS+l3KA
9oT6KXqF6bTes1SUOuNRk6xQiI1SAoQ2M9E3sLSY005ClnNq21vi0j9GtHjVpP7b
PRWwKxVPH1p07+H9Uk91Ar3ZaBU0o7ITUEt61qcGAuTmGjvFklsFt66mYwmRfsuZ
SkHUg8PB50Yv6b0fHv0PpmeyAEICK/7r92BhXJT4QKQdeT/cuNoE0tF9SkcWERcu
QwCNvRuf6ZK5VBX769sFzP1qZRfTTU5hLaXZGeVDGM8ofl15J8NpTvjAYdVUACey
at0mmcNndD6wMGGIYM2hSo3lJjY45HMLmLOpxb6J8IRXC7pRJwVN52DVqf1CO/G5
W6mLfSKLpn1fyCdNVemNe6ny3EFzVO9FvBZnUxPHpgg5OPHcPTSun8WnPSEjm9ZX
k3P8B0ym8DwT0oS3uy7j0ZG7PLWnE+YrFdZB+gjkCu5haLfgnPQXg2eboNbVBz0z
q0fPKK1blr+6ThRPg8Xhg0ShAKV8bPKX5Q9cSXKQOpZ77XDxHZCFzLeQ7J5BRPob
23sbvNcxp4WsXiQO3pZkmRO3X5mswzANcEcQEMLADCEN6wrpR2XRTGMzSUN4kYTq
jd4PAfUwLwaghackf28r/QliLh7vsUOBCfCkBA0rcg7T7pMK6uwpC7OYIRSbLD/H
n0nTy7PDrdVPM6iwAHfbYYHr0QbqccsKreQaRIKbjTd+hb3x8n03R4WKwqQXpvm1
`protect END_PROTECTED
