`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hpXf0K19eTJ8Eu18f+slzFqjatltiZhTOqkBQYE5+1EwsSINbLHalrrO0d0atMR0
PoUOFa0Po2q1fo4erDb4CnrJC5XP3gU2QMEUbkegLSxSHMhfvDyqtmDN5aY4O5ru
TvmqD5XVNESgF+oc4AOjcCzn6szJJ8p7hIm+wxQ622yrCdxR64+z1s5tqH25EyxY
gSFo47gJB444eRRxn2Aq+rlUSY+/ECAa71kVe+eXl9LN9YLHQ7JCR0P2c/rFcQat
hOjt8L7Y7hGdt5LbJvqh9wU6rmHBl8yxTDi3CocJ5UDkAY5z65govbFPnpMKL2gJ
TyTWUWu60Zl3kFkO8pEOe5YOnp2SNil2a+3F3r6QgMDIM/Y2pyu5MdT04rSRUtmb
DnWqdTswS53Q5Hq9k66lIn3qKCaR/hbsB4QLCQDmBjkXN7dz2PKHiYKveh5G7EE/
k6U8JQbPeai2eYpSmAgApYWNwGWcNi/1D3P3A5+am1pY3MoMryzB4ZncR2rI3b4t
/1zHHH2mpNJHEDnM9sEGiqPsPKWypUtzWHhukGy4195J60svF6EWtudfVZB8V/iq
gutoNBDQjtEx7AMJex7anq/iSAdil7EAz9Fu5MP9aIRf0q+hdKcTtnGfZ1wNFe4H
B8hhED5MxSpD6pwv9uhDQdPHZ1L9rbu6msMk3xdRpeh5dAFESQaV6cR8i2+xyXtk
Gft2ekaM94PoNj/GsmmjSC3FpAXc6/5JXjLNSUzTNW8efKzX98fXkxHJae+uhrBT
Et/+nW39pfQelg63ZNLlUl/SDziq9olfhIGBtZY5YRXE4klNhCIBA5sDL85YBzT/
izDNBBogNOQBeG3yYlereV42WOsOqwUoBaGko8CHSaynyH5K88yq+gN1NDusDU4r
TF8mjwV4VvL4rVF5lZXJgTDVaoYDM7LYhp6YUMlbEHqHleMUmTJFKj0OclHdcrLF
/xqOrG4bgOaYKdmkUX3CFlhNyFzgE+9PtiJwCffi+Bn0znndz/BNZ4tXMa0qUCQl
O2Xs64yU6+0aCoNKJMc2A9W6cwF5dlNgRqLX3OVwg0+rFBNKTfFQa5PbSU4UTzLP
xvPvmru3DmD1A24qJ513btYOyr2t6YkTHAUPrQS7cKb96olR4djXoS41ZoI1qcgX
Ua6Fr5SelnuqIUbQ3rW5tIC87Z1AJOXlSPJHeurWHzXcgqxUYgbZR+PbJCJZvwul
7E3xL1Q+kVcVus5uHunfXgvtLFGRhd4s8BzTkN+4v4XxDMTj/77pbh0k/v2JpnQY
Pq1IpUQ2WtnrTbSEGmuwdQBzNh7rg5WNrla/yYocS4nPLAYpEL7ULYAf0i3eH9UG
K33NYovkh8Vv07lSqk9Q0d7f2eKSOlrGybUYAvgovVp0+1pm8bt4bsRC+KWCmgok
wCDgnYb910p7e3Bthep/7/PQBaUKNEv6GWBSCG+uDxAkCPV6vS7rH2W56lNdie6c
X9BrKEfU41wzaCubKRi82q/cR2ThnMurDnCECtjZfcstNH3rEmGDr/Kkwri1zV6N
b3UvbUAZxSDowzX78cOCgSvPO6oBtAgG6JeufUyQneA7PFXcLCrkyaxDDj0PQz/Z
7KeszoBIu1z7ezaK/AEVemhJZeJBKdhJGMzBDrXmRHY7h2pGfRjMbl62LeLoE44z
lTB1OrRXR2TZcxnKqkfKly05ThFyss69OYeGpUg3vX8kWDTm1qcXylfaJRso3WhI
p8aiQa+zCqkDHm4bsW4tqvTi+oE6bug6xAVHw7Ou5Vft2XpCVr0ihUDDDmEOZyG6
OPY/jL8rSDMH8Bc5W9BME1mO409rtsvorHX4hix2Ob4YflTSE6y69h2E2Yh488+Q
t2ba+wM3BR69yGnW3KMUyaUV82yr3MEjnsUGSmvnNq5VgpDDjDB181Lw8QihnZ0M
nzAFLsoVZzCc8lKpJWC60wU5jbxSR5o8PGM1zAohoIOZzJnfvhu33aIdf1NM//4m
KAHRTr/2/M5RapBEEvGiVMC2CnaXxdRKEe7hvEYFnDkJvx7MocINCa4glZKk7NdV
DH9jMON/6Lz1hP01BzH0c1c65vdcgkYkO0fQXv61BeW/vwhYMrxjxaKfjQLD3UKI
VoWWx48w618o2Lw+x+Kv2MQP1KoXSsY51bsNl454idncz4ftoiCQ62uEuS1g1jl4
92vn74tNgAL7LRRkjFrXWi2wUDEfKW2TZGSTSkO7Kt0pWZcJclmKTuCnf0javdqq
pUkMlzTMW47Shk2d1GenLTkLAexp9Ekbnq7L9BSCIutpdtsRRjufpLS8cWmEYMWr
tXPQ/gLgG2I8TwkzGkxCp4Pipn46BciHpddupamO9rLebe8ECSMNbUeow718ThsV
ozRjBPBWhRSkfV1yMxyHV34pTfG0G9XRoPGXMtyR4w7ntYzSxrDIAD29RE+VdNdm
UNRRy1OkBNXtWSJ3CWPwRiLRq822291oAxwcKp/nuRTo3M8gm/9rWMBsBThY3xD9
GpdXEQ34MyGm5L79H9CGjqkJH4G857F56gnnHR8AqDcDaTlseoi788+yEgYnib3v
mO/T3f1pbfuuNVBSC08EdmZjnFRx954KUHAgkJQBkgWkkyzJlmu9sqHuOYb4wLTw
fy44aRfoz9myww3ibKwtTUSNyyvWkrIm9PH8IdGw9HoNWvBTuZsJs8MMA0sZfSKu
XGuweBIj1HhM3YwtbJriBl81pUOmfYEh9Bb7QBYgf6TZZpYhNd/s0ai57YWw0KUp
XXN+al2Z3ut83m8lpZ+YkYxWY4W+ny1QD3t4kyP54Rvl8XWcSl+exHlpWERazSfi
ZwMSchWt4P+pcgjpYd/2HnstI3e20nAQ43aRtJ25tipyQ/ofNKXLORr0UyMoBRfO
hfxR99KC0w4VLQWta/tFZ640VmKcCeeCyE3ctZ3nfdXWPOSERPfbK6TjYVjNUnY1
YNN92UoXg5v2OPrpaGoz9aAy4zt6eyq+8S4telL/YhoSPQUEXFCx/SUyWpDcMEDO
NBXvQ6Vo5WGWCGKJJdVQSOFYl1QvVL5NNr+tCDFrHc0XrHZJPuGUy5sEn+hymtKe
k59WKUWJ0Y4NVitpkF0FsaQgkOfnGnxvnC4kaezFHD9IqU08nl39wJcpkJ1lfkS0
CCaDlAbmXU1nZNKY//9+IzuMhQa6dRXmx3k+hs+LdUEoitPSWRR5GxIlDRTnBUI/
r/m16ow11r0b9LaTlzT9YnUQt2wXilEPZ2YTSowRVRQow6DvdKRrTx3+gN4HUw2a
PbpHr5zJZwG7lsik+PtYy39c7zlhx+VK8F9HZb1pDwL6f3VtQ1mKwf1RVadptXVy
q8TIrw2AxgwPLP+1j9gorZXjZuT9V21dUsU5OPHIXr0WVaKNv94ghpn07E2KwIhu
DrgQAy2NIe+sRDdt6kdvx336Fhn1H7xu3nv248MR1Z8gHfDKAC3Igg1EoClvuGaR
ZDLWAVA6BhWAHb5b5LRrH3Ng6ODK/5LMBM+Nmc7CKVm6bgEI39WiZC/Yg6GnGMH+
72voYHvjkfbac4Aqy1AxFWB0X/hU4Ekjs4bw6FazE5oBoWT9GUJaIau8dcuaVs6a
zYEkMKV4ovLf/adZrl3Uj0um28mSVXXsyxipZoj7A5uyUdk9+O+j1Fpioji6raVo
sdNx/OZRrvxMskd1RlpgQTmu4RNXB0Ajbf8+gDWFhfRnxCd50y67mJCp8aSElJV5
r/O/5teFzjucWXq41T2dpoxuQjucop53WL7UvaYAKo/UP6CcWB5CIG+KJmeGkt8M
mDjWsMS8UQ4lOIxDyZfSTGgXYFewLOpdu6HcIiNbMrCu7cmHYozrcbZyfxccRASF
zI0qfzroR64RA8rWrzkcQvuADlOKP7N9SgTMv6L4p8KArbzczJNKJhwdEsuZBByu
/ZcGckXpP8AJzFCRi2HIKx0bPGSq9DL1bvXacPtmBhpGxCeLuYRzMznE+mGAQ7pg
Ki29k2zcKUYsopL3z7st+JEFGzB2OLRRtirMURJ6btRtv3LRdD5B9PzpxdfrZJG6
K3tGKouCCUFL4H1Jp83siLFtQNqVtIhm8K3BZficrzd7S7hi5CJ9UwQUqwYaBOUf
1tp4ApIATROROqCYpPIqAP40Bt0dMHy1Gi0Gh3Dji9Xuy2x0hTge5/hOzOP4IrFZ
e21oefxBzd5V7rNpvAhFWbeL+UNVtvKDIDpa9eqryS03/h6KQ73NCc+lI1lY0O09
P+zseA3jXyChMx2m4f0DR4uc+8de8JbkBrCusHF2P2l38+hFbnLIknC2bMNoXqmP
cf/fI8H2JuygzyOMCY51c3cKhPf9/+FSVRtmPawDTr+DWzgnYpc9pjoDagoyVR10
QXBsjqoHi7ssiykAhydP9idnQeR/ApGtgXEBQWLAyMOcJS2BD5NdLC9dxfhEYfnt
TwPjZdV8gjpc/KYqWn8v+rzw3gf8WlgxomapOMoCfcG3rmOIuL6pKpO9mGOT53OU
+Myu/CRMYJSTht3JTa8fwVejx67w5fdgq/fNDViRrwLxDbqf/6RnPqUql9Ps0+2U
1i4GniKY7U4/OdIIlhcYeABRlFmr7ZgjD4rAtxJj2sDpjms3AnCW9W3ZicuRrm6h
M169uAoCIUKrp5Z3qithnna6a6YYfKyEyX7z6qLFNE9VHFarMb9bY7IxD+xTauee
JffeDknvGGNwFJuufUuU9B/rJmAPGOaDeq6W8N9NG4JPcgs5edftovUhwcGIuhLe
L0HlLqCIJNbd39SmUdCr75Yy8JzTV5OLIqZZvS9ixjBMkRmCHRU7mnNyiWCKSq5T
eCXqbIxji4WMw+HISRG+9otekhcCu+TFFL9hn9C1VNZt1ejMUxLeZzIT75eSA4na
MQb2sBXaeAS+tFbGlPohN2X+AeTw+QbV0x5s6lD8KWtn4oAL9ESWBr575Af4M7z9
h+YoGA1nT3mg/264rbF4ykIlwxxl6lO5sMoLAAJiAYRpESto3DfNExa3xzWDjO4U
FaHlohPv9wNfzCjx1ZZnExfnRyyV2DHGJmAIiFdnjLalDmrWt6Rl1GIsOQ6wYLX8
HWY8H8I8Pw5dv/oSTgQzZd0jZK20niQsXU/LrWXrlIzbJKV0vEJoBkIIXTAN0FnM
7OCKafCtDbSXFYNOEDynZxnLcqkzgMctI9Q6zJakSzh8p7p+3+aahdEy3jcKX3s0
Ucqe+XXetgX6ovrAaK17LoyWHYUWDq2g8y/ugavXo3Hdn1i4LKy8WvzJDs5YDawS
dF0tu5FwWwU++r/IAe7o364o+02Ob0okUEQrWcUmN9YQ0zVk7hXorHSCHgxuFnqX
iW2mr0ZDEXLTnt1TQUyY2WKlg60QXm58qVABuZYcNfkKpNTIasl2riT/xmIDojQd
nilDoCOnBcyie5gmDOKm6Q6K86VIVvqIgo/fD3Ry55OB9yleM3nAIgasXCCMCDI5
Xv/UVeKNw0qk1v2YP6mf4jSvkYaiBqZ1wpkP98Jn24pUTkf2m/k93gHWJZUSfp7R
nI2386Q6y5UBSLiKn85PVP3kRq2Frfvl38leeevSWVuQEahgIz0g+ofGCDOC/9iw
5dPElPJgyguqvbIkVtCS2HvDkH6X131/ed4GDtM4advVFmyh6cbb4aSQkeNLA3sH
Pd998egs902swcc7K71cMpdfe+EnsZhPIqdlN60gv5Y60UPRDrSntaxArbvkxMmk
g9y0DswYZ0NMbzTDCjZcnR/Qfr+NpCFHdP3Sz8Bpaj78U1pZkk8wRoykcFm0RJr+
ijTlh6Itd/IAyp0gcfUPniCpxMioc8ZgxxEz7cgtblI=
`protect END_PROTECTED
