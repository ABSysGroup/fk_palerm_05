`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iQ9puPdDXuc58YibpCrvuYVh6W9JYq3IHMGmxcBXLLbAKDnkapF+oV+MygwKueMK
GZrjbVlFSRkFkBpfujww+JmyHlKbo2TaSXrGn/Zp+fias9bUK0rd/4wRV7vSvMMJ
xuAKIdlZl4oYLBdRdXj92aSCRpHeSSL2vyKFkpBoOMzK5Ho96qLN7+OcBudvotSl
0gUqkVFETsVMXohelQgz6Xf7NRcoGcKCYVEJPHclH2+d5GP70+5dnRC+JhDePWLV
N4PaWlyz9/cWH07vF6+z+cYJoLjA+Cuq2H5jXfDOB1IlS7A3gzWkioIxXLi79M/I
D7j2QFLal/teBQlkX6PG9A==
`protect END_PROTECTED
