`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oZp62IOMYxDQICvtfgSF17t5MeP4bGEPmnfL67k65+DaFFOmc9Tj/TxOQiIe+Mn9
FOCFqSvueZvKxV+OT1Lh2Nhznk8iz3/+rzCX/PXZSzb0eRLrVR2XA48yiyjqsrjM
gpVcK68X4wMsSfxJSVPTR+8iU+TIClURanFq6lPKh043nEcFwnS51m2F5/fFJXw4
KXleZD/84ePNNwof0Y41kC+ziXZRJ/O6HDQC4mCxJZJYy26ChGXn+J041VbkrCxs
`protect END_PROTECTED
