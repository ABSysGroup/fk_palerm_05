`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JAD98hdvA6jv0CYWxwkkJvPVIwNNMxWJ80gKFyoJiPwTRGU8LGTMPwHrKgE2rX1r
0xZ87lMCg05kZw7y4qQ/CvRo3JIIQJ/u/DzvAWuNd1dpIjutBzmOnlKY0lMFKwp8
SjI5A5bzmgVKAiReBx9f2XRx4i8VYDB7M/Eaxj9HHrnQVQRni5q6N33Ri93qoVxP
EKZuxZEf6uIR2JtroxZJHm6j4HNHSV5F9J/aL2K1+KinRkdY+oJTAwKzsmRKyJ/1
8j6NlVLu/vGTeTZxoM1+dr/l52xt1rGnKtb9aJcgBaL+wkKPkiWcuplApSKnEYq2
b2EDGxq8Hh6vi9bhadxPhoCkJ+8v6XqbTKFPfM2diodzAD5P3Y2TwABYV0OdNq+9
n+mWbyr48HUEQtdfX8FEjS6piZ6S1+MsMmFSpGEds84p1E8be3fnXX2WNnMVeVal
T6fWu8Y0r37BhQWRcXB8iuSBd1O2XlsfnI44UAvS2FlFqDh1virLGuD1iprWvx62
zRkhmqyk27MtrvMjOvVxYyJSrT5TIP83KJeKBUjbf1VDyk8+MKfkmxxXZsuu/qpD
HRNHfWG3i3XiQKy/zwELkhgS9qNpTBs1MHt9KJCacUJinfCCeyj8/4nv0IaXAjpx
`protect END_PROTECTED
