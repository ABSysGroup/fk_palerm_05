`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JQzzO9ghPqTf3qkWgQ1QYrNBOjY+UCcGMwn5QQ4lBjVZHlm9y+3G/eU8ncrcNrhc
AbR4j3EF401cIjyG1KQbg4eW7XEENHWZGuRf+/zqrh331smgJWqowUIGh3eK5vnc
YAohapO/uA5i274BTW3ZcuLkY5OUZC1JKIsRUh5XZKHMfVco5hcbWJQyT9Jv9Qw+
26dOGlIo7JEDizQmKcwXARENrK8r0zBa/AxJyQGNwfivMHymzkJ0Iykhm+p72PTU
uDbUaH2L3+h4kY2qheqORg/jyb0Cck9IURz8jqm/QPN8Bc2fshCPoRwxtzDXJHV0
`protect END_PROTECTED
