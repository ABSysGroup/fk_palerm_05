`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rtvoq65a453QRUhqmb8NVKjBqyywtmCQ5s/FLY5l0N9sB7+h5iK0RXf/Jc5aAWCe
4cLVxb6UvGaDyJKZnTlS/64pp8rxL+GUjA1V/V8xGumnWwfpQvj2dIfNbMpB5Nkk
fputEwBZDidCydOxr98x+fReiTvhcAowrRNvlYoIGTiY/h9bg9LvQMK/Ei36aSg5
q0da0QrWO25FlxPHMKmUAb7xCo5gjN7XadZvZv/JLfTxXHLq7WtSYqKzb8fl9gDy
JN2h0sb81m9MDKHWL3Lq6AgYCL8J2KEhouLcYwXIKzld3Fx5uzgN29f6cm1rLLQQ
iIBNgbz6CDKN3be1jLExUwAggSNfIMFKw012DT7rs4qp2X/PFDc5epuxYShq5IV1
bSe3NpeD6nqKKl7uu6HIHw==
`protect END_PROTECTED
