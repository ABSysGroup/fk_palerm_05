`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yKFLswky8/hlCiFps3Z+VEuK6jY03hWnnBiPHMDKSmSPF4z9WpFaYtfxghFEdrj8
ihgq+ahGJBt6BkvBdvZshG057me6zg3iGA1hG81W+xX9T803zEz3Dgnt3cjFqJJ3
TgOIFEM9JvV+s9pB7s9AvOg8hsL0QIJBMh7lEj3p/kqxR4mjzt4UcHNe0HYuPnyi
cqWKq6OLiurN8WzXIV5yV1Cq22Lt1JyqDhClUtYegkIcG8kNAbnheUXv9+yJl9Td
iIY8EJUUT5hR9/MNXoMX/q/tWoYIlAiFzcPW6P7Pn6tIoY2cPmtpYaAXUiu3M546
tyY8gf0TAiY5Q2cowjCQn1GVbAvJMffdfCbvgfh1DYn4I6yiHBIh1OfIx6z+NwGE
FQQPMMTifKR6UzuIwGF6KA==
`protect END_PROTECTED
