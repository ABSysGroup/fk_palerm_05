`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PHVErnXUxiAgw5dtGZ1QEY2tudvrovhlkVfQ52SE1inzbz5MdryfE1HHS7dVJWl3
SGkX5a8Vadewi0aPe3tfI+gfPZvvdeKvpAwpmKcQ2lLvZREYPXfZC6CYW7w/mGXv
yuoRvqvTW/gDxvlHrleNTR1vtH0sEVo7Vbf8ifJ8iKsj5pEL6TgwTcXAA64KTJ6G
612bpuT9Sds7Ka7FB+bAKX7tCtbdE0wZs0OHObEy+WLBpmwEdRxPHOhzYsIRCL5L
kK5PzvmAOdgNJ/koreMZedQksn5NLQMk1OEDQdAz19M712X3En0PvhJtGpWgO5bG
f6izim0OJwunStQPsxa7Jzl9xW8hc7CHpPUkkG+mcMc=
`protect END_PROTECTED
