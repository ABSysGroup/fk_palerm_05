`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4YNu+B01pF+G2rockkP+Lfte7NSS0abuSzbAbc5y/M+I0f5FQzuYzMrR4NuAb4qJ
B57nxCLrnx+djewHI3sHLdmjk2HMVN2huW7UdoV1hlUgBZRtSjcSYjMI5N9u/RXk
n6FZhlqTRthizdw3sB3MjsK5MbIk6qU50BspDhs9N4lERezZqf9wNWik89vFHr4j
+drwXJjNU74KGjgA5QsRcXkmxQ9raawblyznK6E7FGTAOLwuldeu61qTIfisalnA
CWQK64SmhusBJm0kqmtEIK4zMjnYl4b3ylT0wY7kSRl8aa20eqqOFZP0y3cjCk1w
yoWvsZMV3e0Fq0XwnglfujpefO0p5JBzOMd3yV5rbFshHwNojaSjT9v5To7BR50T
lUwRJ7wOnuFWgIqiTNlXHXvRytkknTWFvQNTpq1WXAHrZTNXdbuxP5EQK0dpr8wq
Dzd1kk9ME0lcCSHvJIu2YPRSAE3oraOfktzjCF0LO8dHUztHlU5mNQrO2DKpG/Jq
SQxCKOB3KHMtnTqDNmi7+BRAyqIhnS11HcCl/CW5jqy7J5CxiCwiGgX1GxW+KG++
ecr2M3ctaY7Cq9ZBnF+hlkS9Q6QTSdbv3YbMgF9gE4/fOHpqVxo3Xmnl2PiLBgzy
ddX42LIBbVdzQpCkwGT9C2vU0Ov/+lfwKP33JCVsH48=
`protect END_PROTECTED
