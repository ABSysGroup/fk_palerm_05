`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xKVeFwBlBrsct467HGBzQCXbCPSbHZn8mmU2dDztGtJIuc1WmQNx3K7fXeP1jG/j
WmifPiW6C9M3Sug2yqzAstw3DQA/QjYpJFtvuB07aMv5tiGAKCfdh0j2ue+gPo0P
7VHoy1yfi93nt9AkWeroeUVYekQidjxTJdKdV6mBpcr91Pm7EQ2uYLogXmEQE9Ld
DJZ42xB9eVtP0bkXvdaFUrDrVC0mHSdIIzFZ5BAvbfEIqOgWd1CVzbvicDpiNCUz
4I//IbsB4e0zpxdnybuCrkIIYl5/rGmowoyUC2dpBMhzaIimtkGiyC0CYtiHzSNh
sJf5dACzJAlehbMiWaZsEA==
`protect END_PROTECTED
