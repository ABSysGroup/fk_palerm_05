`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yOWndC8gdlBR9xGA+/P5T6/bCoXygTpOuDjk8+oEDGUXFls//Wr9ko5vocuszbwi
EAbk8gbHCtkhSgE59cy9Sb3WvgejtiHFn9mUNpsfrlsHhZ4EcKLVnJvS4OtGitJy
FqWGNbmVd8N1jP+DmrQHc0OnAgDuKnsfQNM2rijgsCHvIRR4Yo+sANtvYCWoe2KS
OEGhFv12COLVT+t90zTVuGO0M4lVkRgXN1tIOriJ/vlGqZ6Ecyxcnaamxxe2MpKq
OKWGH2CSdJXb0o7LzjpWA2nXBM5tyf+DGX2/M8mtimSA8rp99qbPpHs9aZQqqgvt
bSFo6BnvDwX1iPbam/PwaRKn3GcIZWzZX/qLaJpfwXaezKN87bhxJI+t4wcSVFTf
B22Pp8BHp2/9UOiUkRzC6hfyKkoZ7zATm5XXcMCEiwdj3HRGChuo26xjuROmyr9t
DNiu55PXlqW+JE4AT68erU+2iMJiFNtGb5kLZlDwjYXPHmKZFDd58StWpGrDOhmt
/u6yw/VyDYTmZ8w4x+a+LICOkcTFVMeo7RahmFkGCkq7qy8unDOSbSDPGWNbPpqb
5vNqqHNv76L926kVIV1yAx8GJHxMFePD7ISmFM06wmXku+dTPc+YY3u6lB1YzMFl
re6uL2e/GE5NqENT3TdwHf8bgzoyECf4bNfZOZlnpFcXYoj333l40lmOawbfaz7f
dSFofJKC7Di6A4LP44dVUvGswAsz7JBvJqQyiHOvtdwFa6rCbSXfM9fxN3ZyJ1Nb
Vuor0y0B5CssHzqJGiWiPA==
`protect END_PROTECTED
