`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3dNopAEi/hog+ikf8uYHUuDobD7p987VSNPwtAxIRagtXKGmOHruWWVGRZDEZRac
QD2YO7jwxsIwWTl4Ez5nQotEnJfWwuin27wHaNuw89r4vO3gSnDhNzY9OtoSb9vq
sORsYQfdX22DUALwtk00lCOUvpnkU+GdIAKPsem2f8ZGGlrQ0Ai0xdV1ktYbWpf/
8D/Q16DPsht9Q8Ov0p1qjPLJ/Q8oR8Q57eV6Vd8bhkkZnSA5z0YRT3NbBBlzRQTH
M4482Jjm8kdvZs1iPYVbZj/TsGHbZOJQXie943IsRLE+3noiOa4KzUNnjLC8e4P5
7cBwsBubk3J17E3NatoZR46vAXM8mtRrRm/9K+Y/I0k/p/hD8SelWy/S0fwuL3OF
bKAN6GZV8n2kCDzs9ATiog==
`protect END_PROTECTED
