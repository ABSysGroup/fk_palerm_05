`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SS3hPTtu+HW4pe0r85HbQ7HnFV2xUlEUNfNLDpNiXLSPf0RrdhdTXD/HD9SK6QTw
huR6ciwQcm5W598EWzYu8MiDl6lnOrTThTOEo7XcDr7NqVEYR8lube51af0H7KpS
gnBj1mfJ+U0hJmgC9SXXWiICoP48+uNI9ZgRRZD3RNxvBwMWNDSbsA9i7Gc9dlr2
59GMiBs6PU8WLIX5j58bXxP6HNl4/RkPMh6+60Kd0JV41vmVKWl90edV9YbLFEz2
/pP4eAkFQ9dgg5BndRUwP4LMQD3H+z77JWGbQhzemWNKjjjO88xV5nwbVPVJFO2D
D2w+Wt9ITEb8nzNgpZ5RVQ==
`protect END_PROTECTED
