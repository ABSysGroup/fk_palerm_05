`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fh1K6STIzPveApZPDW/EwFPq7I5hhTxi96NfYAKf+DuDLQFvpowwoPeTaoV/y5vZ
0O86VIb/Cc4Rpl1O0jvZP0RebPTM73a3knZEmG2rqDsmH4flD9ixgj+4m0KK18Jz
8r/Ye+tZBwQRmypn/Gn5H1Q8Rkuq07biIf9Ho2/oBHEmrzkNNxKtizl+NxoBLKpu
mpj55zMYiV5f6IIxXWb4KBhKRj6m/D05qSDlE2VBoBHLVjVbhveTGiE+reB2pFE5
yu/RwVAlU/OtuB6VSyPFuF/23MI8mn3P0OyvFWP0PWuQwNEp0LfmbESP3X2vnl8q
rcCqqShxSXfP2tByIK7q58Hx4ShkFl8PxUoYPurOQY/oTZUSaZocDiRglYfmpLj1
+aUQhmSLGEuTwstlFXWvvXyljzGekMamVkhdmSytMoyHyPdUGnPnAZTJOkIZHHoZ
5LzRDWuuQyML3uqY+5cAfZFv05A3xwG1e7RsVKpxZ2gSF5bpCXEyMrRItCPUsHZs
Fo0hx9ppkbqMQQDCVIgo0SVKoIq460TVldQV9/nt/Djv0uL5RJBvPkk6caibapj/
JBNOpGbIbqy6pqvLlZ5WxSwpHAdxn9S5Vqje9DD7Cu2uHD7Szf/bOePnDsKgaP0K
LYYpw27xLLWCMP903TYl4GDYLhgi+7ofSly/45TFxODHAeMb14eobsekN7p2U4Ei
`protect END_PROTECTED
