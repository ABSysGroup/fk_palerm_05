`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iFzxybXPC+7n58j3YDli8Vkx47OLXumvzzAmWf59rhPI1zUEwY4M4ouVX4g7d2AK
XO6VIU7EiEYmo0En+6t9oifyy/TGv/LONV4bmfG18430gGA40p274FpV9RKd6iVZ
2znjjBBDW8qTK2EoV076zTA8469VlAst4neCgmnwIzD4C+g+nQx9Ot4WxX7geIbE
ulsKDy4wb8qN0+qIHen03dePVv3OWqTh8QTEWYJvhBsHlle1l9E7m8GFj+xOZOP7
m9/977AgCQ28huo/lSR+KnSfJxRGS8FUou/6R0KETqV8+CiykPlLiRNkAUj/T8rJ
yMlvY7NH6z0Oy49mQ+IPxiYetOGrRjbwawxHCF6x/1BgRCoz18KrLxi5OdhqPAxf
sRxwBiwECOiZA4Spj5sytVnEtU7WNLhmaoCnfiN9UCl9ZcpIt1bE2l7ulOIJW2Ad
tkErT8GupwMYEXCrjLtvBv3eQIlDnfCtV0JPHegVLzw=
`protect END_PROTECTED
