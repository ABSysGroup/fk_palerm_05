`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tXppu1A+uDalvTJeoaxuU9qtioB6boeW/DnFT7ub8WamRkONdrlVO+Stdy3/C1Nj
B2Re68ARpDqxgfZw9/+taTOzJTb3tj7Yf3N1wykfACw2ebhKhXrPUo/q5UWae0Ei
Zd7Ba5W2qUpUjyKWQRx3moVgCwtl/nOPhY1A6FA+K4lpwZWgBhy0WLPxUaaBub3B
JVD5/X8FhrpbOcgynGYOg+t6OStWeTvE5OLc5MiQ+v8nCL1YEKax0JK9MLaAK/2R
VyZq6aodFqp5WFsqhVteowqu+bC0XSdQ+9DLNJwXENfihenHcYXFLeoFWd3YTERC
NiisZFsM6Ea1QUkc4UU4oprTI4M/ot8vcfH2igoXOiSUACKHkZmfMnTuLrNrfMmD
wkzvx//7aeP7CGYTA7114e9FBpvATaV2oWaFZqJDDuimcss7MfT8wXQ7gyY8cfhG
BHFTq2+SwEtSkHHzAxE2Yf6UzF2nBO1GzLi3q/9TSAkI5uMWwVUvk9w4uFIKvil8
pf293WmUWC6rzDSkfRejkYQNvFNbuHdHFTE4W85urwEheCDsd8+YCEwXEgww+yPu
XyG4tLbvsTZ8c06i12Y+kZ+5kLetT2PmXc7aH/WtDe2nkiJIjfbvsyHxvgcB7h4i
CZVs9dBrwepZQf59LQ6osGEtmN4NPTe9kZNWJBZnHuc5K3gYHt2SZLRoqxDvMWG4
LbgCbiqth8fvHTIkdPlKY5naS7rHb4QCFaFDDpiys+yKG7H92NQzu96RxXB9O7nc
dyxWl5etQ59s7E+mTVLhCv+sn6dnFCROmddh4BTs2nLjbockt9+DEasEAeSnhfOY
60tU3yyiythq6tePxBFlefJ6ScVjTuzEUobtSQb8CaJlILOnHyOA2qpRPPJIsX3p
f/0CFX2EEOsk7bV/lDxrmejxBaWvfl7rhGyfTlOYzHdf4sSis8MlOsTP2Mta0ltT
+UtPkS0Q56jzz8JAr5b/8Q3Q8xaifL/fojmbqYTt9Ff2ZxTml6Oke7fkCwTbezoB
uvXtrq3chG5tRGLAElNrvn0O34m2HdCHFXsPf6ZaviAzjJsppPWKpw70OrvGCuo4
Ebr9dWi0lw40vrvJ4G0+UPtpLgjrsweTLXAU5+NmLzqSFYSJMj35AumQdibl+sS6
Fu6CjlcSbE4A3X6l6vAb2qKEuNt2lfLXL9jkA8VkY9U7/nToIvz8tCn+c7KXr4Rw
/K+fEVg7p+b6Cahp7uE5s5m/Sv699ZHPAHSZr5TsFNtA5NWEYQksaSCvDpTAyM/8
oQQnjfsVLkQwAZ8rIPllC/5FMvlTHcz6On/SHPkmkrjovSUB3mJf4DmtWjnRCo4T
J10f3DLY3G3hu54Ni+81Uthz5NDNeSwOb5DVophxDUJ6X18vL7mXpRUaDv171Kr0
SdKUWcMskviM80O7A/g8bmdZWPV9qZZblsfYQqzVbjD5yoUENm+j3wMyjQkPqFzO
r8twAPvR1RXlInhU5TWqjFZbsWQrSaEayLn6ORXRSxR6+YFkD4zK/SfxCb5nVBjW
Wzpjem8YyaxAC5yCR3TW/JuFKL2QOoYXDh/CUOZ/ignToIBolmf0vTgpcoo+BGyR
A4fGt+s3LGZ7KS4kHXXhMXVIOzuE4iIJ9ppMeqH/Z7s+gR0fQl5vqppiWiNakQdN
zpC4pK4TlyIt/Ym62jSEpOfVzqzgwF0hg6LXMLQlYMf8QqK4/reyS6dwxVLzFw/n
BwZLIyKKzIq6LwEvaFbSRZ0+c4d7Piz0lWXOy7DT3sUf79bzvqCxMfK8YC/OMd/e
l7cFaMTdflp8z6SCq0Fm3tHTbQvDgkl6gmuLxH7CC1w/ZmHulgdvf24D4lCNxbuW
5sElAiryG6xqdur6eW9K6YmTBX8iZjTvSzoOxD6Pxx88TKs+firNkNdWTM8ez0bG
ZcepmBIpFLaF/dzybje++k4kLyWU0LNC968mBUqdl/Q/n5LYltzYnei7skY+kpah
tJwxrPbQ6bLaHZIp3BqqNQ7zcc52JOc22LvXu6kPdMMsv/vudC2ipXqJMTcvpIKF
Ip4ljoXUQsjxgS/m/xt1Jl6i0dcySV6UXU91Wu5802UIz5DuGTAKHr6TjPlCKeF4
BWu2FaxMw0gVj8cMc88seMuanhnTbjWhKNpaUKf9SY1kJtkDHcjipH6+2Yzt8D8x
QwMeNUaC3W2sKdvVLuSRP7ZeyshhKbZNiaY2/841RG2dT/5HNvc7ZqdIQvi+fw4J
JxJXJd9UWpzspX/dy2Y4zeKLmUSJTg244H2AT2k54rS3F09vZGWMslFGU/1KFsLT
6bvFzY+YCDX58qjx3IGfIt96dhVPOrsRTkO4BThJwMzsfOPaCARm7UEZ9oz1ToRu
6LHfinPCQcWOf7ZbF/OHNBFstxQpEwafX3BtEKLzBRqssO2o4KxPvzc5yF4dv/oG
Bl1Mg1e6oLwkKBl+SF9mxOR9J2V9jUL52MfMKPFjbr9VRnRi8BeRH8eXwliC7glU
aqR9BIzd4jAODjDulbW1QthAvhEuZrphdLAUMy/7OYNJZjM1078iF2tc715WCLVB
WqUr+ri0AJB0eBXmVROmcheScYc2rkk0Xv585/zWvojOwsAiMpLqMyvs5nUzNV4M
JVRRjD6rI1H9pV9umttAHezyObUvwLKVlEN6OJVvrFWR4P2yk7C7yk2Oimfu5qgk
N8o5hhOH5r/vbnzoGL1XbnXI49kdtJiMEhWB3NPiFQPBqDS0HmYwWav92pT5/Ost
TuJ/ZaVAhnvrj9TgHx71F3HRcfyXn8QPKPBd75iWGs05HXHP+gQDMGuguQ8/69DP
l+NHN/EzjvpDFkQThkGJD1FPTaJTgbnxLje5QQT+fBovfo6znwqbSDKa2GI4jsPl
rKttXZZn/fJmxRY4qy1ocIJvopiWZOyIjQFvCYzbhBhhQeAyZ2EwGzMRzWLN2bd/
pZA5fyaqd0kfQiPH0BKvaMHFXD9CUIYyiChtP39fAFPYgAeVfepRfd7Zhte9IXj0
jmY7WAB6+XMwGhX5njEFQ1lv7uyApUbQB7hix/jRMTznS4ZhKGBHFIkitOWtbBU7
p2r5GYBxEDNKpVkrXooBzmaalUnacprq8HpYvDZyyQgDeAlizAzB+vdmc4TNFxbi
V8apEw+pSLticuQ/9Wk5/b1smpUn9kPlEtOGJ5nCHAmz/Ti2yEX+AnwIHAGTaQN0
hJoY5VNtwJubkcNDnqfO2VBR6VALDtJauaLpePhccPOEqzc45T9fOV9xNMCMbRaW
RkE5M2dPrNJ4CUGbMkNAt1nBEVp1X2qTbgs5nfUTXBCXmdcMkAtsSG/mBdd5psYM
AGIrI8W/e6jIlX1mLGnzQUNHhiUQesll8HlKMxpgRmuESd7M0VeB2Iv8xPDSbWR1
+6EXMruZKqOyIPanZOU6Yn9iUdSU0chqQQsztMT2z28/vrkNNYYwQGjwA3sOggZD
f9/tqlJ5p5jbQn+XOexAwNSNEA10U2diSDPiZsOSnFcAQK6k0dBl8gN8ZfjXtZWZ
2PaFXmT61EoF61sX/pz9n56gCrOCV3QACb097InvkTQDdZVeGqPM74BZYZo0Pkgy
UnVqXm7EnlF6dwCHkVmcXpdbKWTcajYfHUtgac7m0P82Qz7KV2JY3RS/A2AmxzEX
Lzpv2CUUpRa1nXooeLC45ucj95TbLw9fMhns/OKUUwCTYGnCqB6WwR1IiMGzPd6b
gXi+8UrNGn58k0BXMlwJQULDtKGCQT9xqnIdLll+WnHgslNDSGneTV2Y11aTKqia
vvu5yG26NophMNPb09pxuLJ28D8QF/CQ8391LlwjfEDwzj6JzFSLc2uXQOTTt17P
hIJwE+ar0Wu3VhNkWlmBvDbPX0VX/HJA/V+gO6D0WxOfOC6Sxwq6Z55AoWn2JVYz
4ZyfA51/qSPLwMotiXrD3a8Z5ULQd3cEieVTnMyIhH5yUdRx4XILUH6OT9eemE5w
Om1xevdOpjQNFN0Bfxd9sTTPo1Y5dG73tW5a++LX8TjL6L1F5nSXQaxripYMp85l
M8w8Jq054MFwgkq/CrALsGLGSMDFtwzW8ZoSgh7u7KRXIQZ0m2Q1XDC1P0gXJ9Q+
pCYA60vgBbOuKwItVOT4FuycP7BUcdiC3i5jcpiEAPysCwhx44srIEWx7lUKmRJv
oDe512RrBVHVnn1RyMy3vAERLa7R4a3pELLt+x1XuE7TApo/RQ0uRiX/pSFIbC5W
+O9Ye5KbvBL5jmUVOArG40Dlsh4Z3kDjJeRw0F00WFPxa89gJvm5Ds2zhFkVKSw1
bfFfRGN4mtbNpYqHvKwog4ljZmpnsA8pZmRaSBclfH3efWTvyW3YxG38L0QwwHeH
JhbQ4NaAfHvkXqwRfFw3QqAvO3xwEZ+MwvVij4IlS31pu7ucF3kqh6qxIeTWalkb
wBbQgUfDla0/zgF9fssAbe1yzSmux4VXx1T0wox6XW8qChXhG3HSmBjwjlUScQlV
6DuNVWc4lmlJp946O+5qpNITcOn8K8TrRg7YqmlukqfKVjD2JDJTl8mxk9exPd63
hKIjBKhGbXQmeFtZUeSZF5mgcwRUnpnHK7b/okjjGVgIoHJvKnsAgvOquwo7CkGM
hyBKLrifnwqvFu3CoZz+XjFDJKX5VpDcwwDX9SbeeEHmoVdFR0iw6H1h440Yuzsk
MgoVQzKgbSNisUejgsBU1KQF4r1Hur2SIkxN+0m3E5NHYELzH8jRV4QIyz3fLPvW
6KkxDUGNg4ZubzBU9NyT2zLrAtRuAHnrhyfcoIECuLsonDy+Pa27YxUHQXjGhfVM
YyjHh1iS3k9+WrdQwsiYkA7BwMqv8+oHYMCsk6/dvopoYcggBrCDMtwkxXHjUK7V
olWpyO9+uvFLd+k2eFAxhK7ppd2GxouPWzDMgw/wG96+mY1dkMFdrazaaxeuX9cU
92GliHDIQXHr5BRbXs2hJgss959cDomnlj8VXzdQF+QerrLqlsrTOoM6/TgBZKvr
YFQFLaQzaMixAKEIDzmowXFtlmSd6qwysOVOaC0M730FZ631LBEk+14lAQm8w2ro
QsBymTnTVl4D73dLbBCqS304Qp5+kyG6V8SFo7O6DFdfneWWJduQhAQY4z3i+oe2
0UvQt5SKQtmUo/rRMlK1FzsCz6XihQVHNv4tvEPLiCveihK/LT4KuchT4LSjvN8p
TPCIlXcZ//bSpYQgJQTBTYVJ0n5MWZ9KIi30UDtfWGINp2DLUHREQtQ6HxsSwOVr
/qxJExzuvkpHU4IOT9u7ww7X0IunzkZQV7BqbjWu8xE9L3jcltGYRCN/l12Nsd6r
V+5BSbLxIQf2rzJfAsaHOL2pSmEJuWwLpm/xu06qTowDLaAiXVihZGN/5aAzQVvK
65CdSDtrSGAPSq9azb9VtU2ZSyfOCosAl8KR6VkRclKPyi3ezCEvBi78HjuS/hud
sey8fCbSjCqGj2r1fN9PGOObd8RPKpDd03T084wUVOGvkW7C5Ji2tOGcqTpofH67
wJcd5uUGPFmfuQd/If9W1NXEABkEPvbctNrbGxtzNe7MN1mphKTOrPl8e8HpXa8k
WTzYNLcZZzg8N0XAhQu3xPbvg90InNYYUG2yJZezxEfjGDtWU/P6bTHt+kjMxKei
MGeG0q9QIaSz049rtYZFmBIuLP1zgZXhUvI7qhPX6whFRG4AzLND8pB5Be2ei4u+
Z8TLqGwGv0whesDS98nabLpFLMvFp+pi4uJAtDnMwN1ZXF7ZhD6HTmnItA7Jl3H+
mXCuX4gh3zIGuvLFIWlXCGgizpyER3/LoA/0rnCThaw2IrpY0GlmuEqHURKeg2DL
1BBQL8DDWTOQN4lScRFpS26w3YCeApbLpINc+KZibrWcLpmuWYuJ8PtjHAP2rupB
d3BtLs6qZLQJw2G0CI1MrGcKudNRKytRWYmWxVIjewI4MKcv+GqtFwFFTeNmeX/C
86wDcOTkwcxwX+pXHDbKkiDmcAAzRpG2tMX0wfvcT0gfvTFjm5ntBO15SMddWnNL
cTh8WGPLTWI3Vm14eaNoApZOOCCHDyaLhhS97G5Gq9Wos6vug71ggv1DEi1qMOBx
ZHSwUHH164knGqFrp6uY7I93MAtKicWGhRdb2B5GtYeeCx4W5GIFKQTx8AT0blRO
gANjNbBbPWUz8I8pkK/hxrjWqklOC3BjyhxewXeqt91lxg+05JJOcwZXO8ndfgB/
IuSjFvEYUP4dgOFuBL+ywQlMp2iGfk7q9oouZoLvs6VMCgpKhS6456zTTqiklJU5
6hQW+CHRHxNkHlPt4Aodg3FugxEpzMIbtVSBr7N6W/Z4J34vp5YQKRm/OBJuVWg9
S0I3nHjElVyC5+HIsrLk0DXOJHyoKHjMJAW/1h56e9QDjYyEPhjS02N8br3mcW+7
sQ7H43FkqzanfLWI3XTw+2mihvkQLPbDRM93YmmcSJnWxpBkwaLthWcTRloqE/NR
66c3dIzsRYIIG40+5i/Hu95EKWleXc1uiFcMx6o0jT+xMqus+sfuSf3T96EmAZHa
OpWOQHIJVLEx/UsW+htrmVe5uMiQhniNdU/kCTtryQ/v5V5aYsSAtcMldCit7YPs
Nfpl0b4WZ5ueQkKu0boXqCYfO21Y0YACA/PhDnEcet3yrx68Gfog4CxeZHqlc1qo
MByj+QilInvy+xrMX+9wDQAzJ4F7s6++gHjdu18O5dvl+prgnZBI7DXKDUmS3Fma
BLFjLZiDKgiQC92g2AbBxEmdokss+UXYkNsYi2q+pqw/VZtACiVCz4EKDAZwsGJa
dpM2uiwRCApIbaUkXIwvtw56anUJSPGmtcaN1K64nEh+fSYvqST2vpMFNMbvpI6A
KOIy9CKedVZy1O5rbwj2xTYuRm8wZnNK7HHlGxju0rYvZl8jS731+rBU6AYHl3b8
EPTcRxPTTUDhNlmqVQuqVrL/145DrYwm4lFIeVIP0cmiXbpQq4XHhIvhbIIPkZoz
CxQi8fn3f90q3dTbcxnEJrKgGDD/ng+mgWAzVJbbXXgOcnJmM6RfVFO2H6rCEHRa
rxHS/WzxZoorOGe8V27p4tTYiF83P8be7jwI/QxK2xhu9qZRWf3HK0bzjIWFx/EN
HkiOqbppw+B/i0haI5jux4r5aXnX4D+qQ+lYxQOFo+dsyUW4qaDK2jmnVYfkOABa
Dp/FN4lfri4QzGEcheT/BDSOuL2L6MwJMqesdaoG2VdFeaNINSuZUZEaRntGeq/c
fV/B2h3dqaG6CqxD3YMMN0igUjX162tJY9//r8Mp5DR89eiV5v0qFDfvjlypWYFz
amyyfWoO17lrIW5c7eseWlDYkchRGSNNxycZ0BnSenC0rJUQJGz6RHvwNq9T0eDb
LO8u+enbR7/fMPMF77z+9hIOGmM8Zs83fsoFCbO/MaM7S86hAyleuWCyEn9Mc0eh
7u077lhOiBxvxatgCiP8jqnLS8Q96d3FS+SDJNFanLECxIPKQXFTRMjOj+pSH2m/
mFLuPdTv4cneTn2ILgpXR+RFJLfn7jQuIFX4zcirAsg9wX/+eOHdsUWQ41JsG99M
szFDvdRF1Sx9V+cowOyL7mcfgRqo12d0HiMdFYZybY3Rc5LYRbGA37w/O7xi8Vgi
7OEaynQxYhJKP/ymrMqohDvUduNNP4WV7CzehLT3W9ORQBGTx623Res3W6mtJ9Zb
aTW17s5F3551GT8bykc9xQc274XgkmWUdTw8EATPzGXILOMQsWVtrcgHTivlgjGP
29CJRNsuRbsqSxladq2yeOSw+eB2MZQbcxA8EcaQxB+sZWbUDLBhEDwAj0SFFIdS
BgghqiErX5GeJndMamjLqAODfkB3aPPxdT7oWcmOjAuIn5llbVC8WijQg8/9B3z8
1kwmfEciRxBfrtsUTzfetlBYuWze0P/Ajs/B/VCQiBi5oMuRfQbprLe0x8mYeKAn
mG4x0ZYzB11oxqXbiL5AsE7NW06ty92j/JAu2MAR/iAbgB8rWtxkFzZMxUu/B7sA
ya3SKP10NSwTpB1zydxEOzmzzJ3D/h4G1iyvZTiVBjKQ9yh+5+3mee4a9QF9JDVW
JTW7y3E7TxcFj+9FdWpyMHQ6AoGmMTmi2GJTA819XvUitMKVwtXsQLOgds+wePny
V58lUljC/dWAMmrZelwEZlLkBnKWROpdLQBEbojEG6HRSQG9cFauJBv47zcbZKlv
gc0n9gWMQQJ+LrnJeFCsHF24VD4M2WzSG/77FMa3KhmdFYIV8Yyee0/Oaslkc1US
MvOy6mimog2fOSZpIkF8ycdIwN6LXf4ZxoagVKk77vkCLaffo12or60EANolp3Rw
Oi6r3GQZ/Uu+JoNnF9DHsr4ohhhcC3NWA7lMGEIlmCcSyMi/xlJx8jgeg2W8rfZR
0dQrQgBsTwGkc50sC4jKHdVn3RXsWGRUvXcTgOV+w6UbI3jj8i7qnVPsRNnnUAJF
7fYH6NDnyZYQfI8ImMRK5FgHtWVvwtEGhyVUDk0fwKxPemM3JrWJ6Y13LqBe92SE
c4gvdoPY+Om9ccA2R5lG5Q4qePbHMB22vl8GjmycUvmdz8IlpGCBVkdpLF0SMr+j
20b+kiQYnnCcroOlQGBWPiD+Sr1CnZoDFblWn98Ni/9J05wCNJZ1kJ+59jRWYhEf
IliTu5NGns5CGhRukYWzXMfCXwL50g7szkTdByaMz+ZgjRby2ECTYoo67eLulkTm
dYGIgnnSZy9m+bAI+Yppnjz/+bGZ3CMPcbokFXa7NBPl21uBw72xqB6oMr7wvuuU
cMwUPfVxq2yuG/y2eEyly2mP2HVx99rKxcXxdZUd0OhcGojokdyvvrXOYGg2QuAE
0wHOR7Bk3NMB3bO7wYnCJ2gHRFk9ZWzAARHqZiRsxjrpfVAGpyMuwMAGkUbo883K
9EfMy0iru4PMmz0Qa9xjKgr1kqb0bhRAzG/4FnhyBZhirI+z91wEyrHpinFWBO5S
duSz/zyQdX4h2FhZRz95IOKMyywefls6NI4n5WpTzc0lyCtdWgzNSlDV0w5u85sM
12LOGFLerQDfUfNTK62jEKl5JyPeQyDgnlAR3qHb+PFWztBSfheKq4o0IudUCYoF
WYNRAL+E/usWH3a9mMkBeTSSqV+UN0zcYa+D2zh4mClHuVJy4Hk7bIPUJQzuIoL0
WP0Nb0xoD+hV6h3rfCQw4fHn3xm/905AGIuW0Q2illwyfKebqlFigvyeQFD8FgX9
nobwfZS95jc3xZYcVm1MqepDHJZrUaa0ocLpN6bt5AToc8oPUFCSzZN1QyIUx8RS
z7UcgYlfD1K9hlaKpvAuAVTsCDw5Khc+YiZaBdeoNv2yNZyltwskg+Qh4vZs0E3a
HVvihfN0xMM9Sflc8pNF4oL3Cv7HtnFfUVxpgUnWYSv8vMbyDkCT7IlyAd3NbPsR
+vAWx+FiAVnIYebLryxgk7bLVBaIR9aSHx5Kl+zSA+8ex0hnNjvD5/7bOmGieeB8
Ab7XuwmoWdIjpdHOMPY+oq+KbfYg2xz6KMAEEREhbeJGi6BShEkno8omj8N6l4PE
FAfx65tH9SRBFcnGfKSdkNks9XQeohhNkVdIuEtlqi/uaiYHb04Va5wyjDsPte3X
TYUyFwo6hKizjWFQ4wUWWyWZofBEVdWcECS8p/LS5+atdU/pTeVK03k1GAaAEfUC
WtyUhTD9/gqkYtM7h2QW53TV1Sowo0y1p0iooqaLkIOVFvMok2y8NS4oxsb3eGhi
QN+Kf+GJNv2QkBPmTZ3muwrtVrU1TfXptR2wXvYrlKEeFxuJRmpd+q7m0TArb7T+
RwygPWzh12cCE5cQDNqIkIEJgnmtYYK/uBmul/mxYuarV260i5nHgSMkWZrmrA0i
vRWcQ4kSLPbGdE3JITsCOoMa/MnNuogn3jYBu3P2J7oQLyWZiETiNzSU5g5Wj2ca
YT3LlmAEZ6cCDwf0u59jEsEPlVDQESDl3dR7ijG2M9svlTZXRETe9FNnGEA1q2Sw
oAou2JDKTRV8wUcmZvq/XxKb8eBYi/WIpg5IOqDb6G8rOMb/rz9YpOUtebaagmtF
JD3mmmyZMp+X/uclhBBgz39fHv/lGoeaLmH8EC/E776EEXfelVnb+tePl8Ao/6R3
gZUfCJwugJ4LFexkEVbGPS9VFzuBQSkVtW8ursJ0F785VdpINdnLxXXrnGI9E0S4
2t2EbVy2ngQ2OUZG3NUmWxBDPYQQMrmDdr0oP3RToFtUieDDRbBP8NVBNEV41pCe
NalbD/gSx1uYz9fMoUPwX2rJtLbnmlVEy3pdziS+IZi2MsxmMPVSRB6Ta0P26C+2
PdOW4twoQJCh2Io2q+CjOhCmoGHDs68q67z9kuop7Se7v1x5owWBpQghsV9tynfH
jAO9kIrfeHIFV6syPpe655mpaJTbon0TYPUa7grSZPaAH9fPXom7RNt5EW5LAyDi
Vd+8+nnnhrk97Aj4s3r9DzYfOsGqd2mdRES+PG6AY5wxqeyV4cl8IX8Y1uWU/zLY
KnZBCcLgANNUbST9zVaUku24ZLik8TyW0fGGk55at2jbFvNMjKrF4qDMrhZ8qcPl
CUHViBB/BGoACxFBoXriz2Bh9yKBoUEiMMqZOGh8uxdnZQNHfL2CsSpLB4cewJ9V
4JtEonAVhUFlW1DGRDVx/xNxlSyxfXyTsNVUTdu+cEQA9TwtJoPsXbnB6ixBcDUu
dDlXG7dKpANH5xeMy+Ctz9Xl94kQ3Uu8Egbav7Z4YOkHx8v1fnK0aeIwWv+Ra3Iw
IKWwSikT9TzW7687Lt+r0lSF01Eb9xAI54uVmxKTjfl0sya6uaIqqg0zzW8GXQ3N
ANPZAsOQsbbZ+I2Mt8x2thfXn0aLUTqQcFnshAKdll4zn8k7QWtN7l/nsoWFA1JI
oc2FHpgRzEJh15jVbjjRNGAPiDQUaIG2CYTFIFRdTNTpg3/5IwT6rfK5LYZ9xzVf
K9dJuENztk0chcNJN5nZnE5urRS/S9T1RUbdmAjNYouneqQ3QleFA3Vhb/NNGL0Q
QbUvIeDcjotbqFG0P6eH426Ox9pCL/4MDqUM1GjbnApt+wK4CAxpi8MpnW/aU/wu
tCQf2jXjbRQtinT34ntSK+0cTuNOvlhGEGkSQLtpHZiFI4q0uQpAv20qNqp6B0Ic
O1xZX4OW0Q9xwwcJJqemATY5n5NRbpNu4r7rCvQ3TSYqPTSdYRROSmGh8iQgRUio
Li+zVBI73vQddj0siWdL428QIVv/uQ5ots4RLgP9DHqWarwiaZvzkgzvyE7vT1o+
2IIlHWcX6KXaX77TKA5fYeH0VLDyNEesT+IDzpysCISaEa41yw6FGfJtOZxN1FWj
LLSv+qOhDPt3fYC1cOGDPwqzyLh5+w8sdr8KRZQuX53nTP5vSgeiJOqLlBWNZ4El
IaF2AnE2rgrEZ3q09y08AQ5oxKsv3JH26aabYM09UNRRk1Y0kJ7s2WVBnnerliHK
pOEEI7x2MXgV5YoItgo2D7NiNJYdFS347ADT6KismXMFBhjW3mp8xKaWQSWUmYEc
omch1iJpBNYy56Vx/7I2LZJmOXTpZ4uSdToM06TsGW5Wq1UT8z+9z9wPcrfm0r63
qeRCW7S8iZq1qOZYYfwBHE4LzPRW7ekuHy9L+sXWifJN8e1pR8gMO4r1C9XVCXTc
pvy0XY45PHjF3+ZXrvEAr/xU+pKDrfXaj/yGcoYbJrdRET19wNtdUGXEsWbhZOR2
g34cahzAxpN0kBS/Ywc6pC4yikohpwxfRQEtf/z0sjSjUkVrDDytc4/kIAMSpolP
zMjzAcGxY5US7fgiBN2hJYECH63pUcCyD/xGx4NndzobA40HL4QaspSIQoTybg2R
AZ/dKUEWn5hyTGLodoW50OOrewgydtm1YsqgxekqOOSAfBeIcKjFFlUIZek5Z+Ew
HO8gGsIKEuSPFgRys3m4qlGqrd5WBaQk1+GCj8y/i5kQWDfMk5OM3vP7dmmkNYy4
tQVsv2tBGK6SBWs8Dd7ADDNqpcf3hrS0bY0UGD1bCySlVBJeWnedoWUNcMlQyjE9
Xzv/IzemFqPOafZUUqyt0zKEqRVhKn+CDUVIGHUmvPX0ZtXDZR2LHuUjxNuLO+9E
ooFJ7Pvzwg98hXX+NJs3wlKgi0c2mY8M4byldIQGyO2Y8r9J0qwg7cjQFY+qI6lJ
y/xccaL7+aWRcgLuVa5IaweMZxP5s7dutSU+HUyqh5SL7XnWyyQhGYMozcTSvLm5
o/vOboHHOVgvpb3cRIJt2333VauSAsegOV2J8wYJXgYZE3AQJgYQbf6qBAk7QcPS
N083+aV2sZX4JYZZO9Epe0jBfi6J0SIqyq6mXh0UPmyFuW1ixre8isB8oYKcOV9e
o9WebROr+8tWHqth6pHPhH0YoRwsEVCEl39IyE9E132f6J7sLvFazq70uDydCvm0
Mh9cRaPM2wfuhjW9OsneAdVrz5CipePXRpN8FR6rAJGHKzO/LAfD+UqoLJX5wxdK
C3XsZefwHP8jADg8LXTiZdsoswkegVRcNpmQpHdnOIcFxmj+5iXYQffry5b5YtmQ
ZUgTv8wYOTQ7/fp4XTkx0kylpl2V2mJnpam5E7LpBHrp3xngsQjOmt13bJs8xklq
oZiw1rkt6UK7p83qzXqhkILfhiufcu7zX829uu1aZEBP8lh0k2SfPwLw5BD/o91G
ItrYXuGam2DcIzBaRCYA4IlCaQBuZS48mn9vL9JTPpOCMvj7NxsG3G0ecRF5ZL4D
3fLqX8LrCmO9rl+h2vkObTWN8d+xLb+jytF7J+f3XpImgRiZjU86b9jXQVXhbwTk
OGZv8ET9soEOfIlQb2vX9oSQ2wqDoGx+RpEMrEguKeXqAxM0B+XZ0SKgF+sOi+z0
8/4BPRhIPcEvt4knpxFvh8B1yY/G3qdU7dzxtAstCJz+S+RnPFQ2TNzOUSka6Hd/
Jba7zInPRD31f6/Qige7FhzAulUml+mtbOhLAp6xLECe+bITp2NN+LDBI3TmkIXo
yDYJeiK9y5GhK2Z2TZ+vUE5FgPmtKAB8Hvj0BQQ8kqa+xa9tyr2XJt91SOgoOupi
HZ+pHydqh3TXrt1G5b3MJSvvaBqsJWvt+tmP8OjbcLCvC/101N801aq9MEKbbdH4
w+68aN5MD4J6xxZ2BUqru40+5oKjnLy7lNoKGwIAAyOTTEcy7YhPR3uBAYaIUg7F
XijHnV00gzfUmHO8GOY06qgflT2S+g/n/8dhkaz7Dzg3P4iZV5IkZAG9aJyz5WJ1
kNptR4KJXAyfZnzBNzHHENTScyxx+tVNEjllbI5dOzvqrG2aaW9QTgrYB/2nyWPO
nePwiX2CNrjde9k80qNx0ebsfCQUj9BY7eWfGqqb1Kc/YJk++a6Q/cc4fh8Blw9Q
TNe051vxD8WRgV/CQyOu8wL0sznoGJ5RAEP8OMtlHFKbHXfNEdPdy2oGiM1yD9UD
Qg6RnmflCCkfL5KJyFz/Bd308C40nuYzGECLIbDAklXRyerylSPfccUTjdJ0y7v0
q5xKoS9Zy79CJOj5Iwa54AXvUjQNnlg8oKe0gNx4EIr1A9BkcTfn7U8qZytEqQSw
tJ277TPtSuIqhCaQvyeSGGSahCbzGY3A2Uxtu8Ok5eCndhckgWlnczoYbau6JDyO
z2GogmmBFv0MmCfTcMmForNocISPEWwjs2S/mKy3BImUw9XjhUnovsHfE+MioxlX
mzDdkyl9111KiWe9Id3HKVYExmJeDUyEooGiI7FpT+OMqIx5ZEZV7su5WrcZNBZr
CGKUckpy51ahiuJxIuZZ4dVOXrHI0dYeaz+ZZqtA4EqlVJ7N27N+XlU6LRPsElNH
w+CA4x1FQnhTml/gwDHwY1SidXjENSw1h24sJa1CwdUntk3wXThcjtKRj/JBeHTq
VGSTmSj7gdF13vxqyecIVDBpwhgkJL7vXRDElX7bSNjOlSuyI0Mncc6k2LguXiSF
6CN08GVCcQmaaoZ5VhE5gylox0EK2Q2mpGVHuHBUnd2sZxZIyUYbmqhP8USazHEy
RSq4WStjT1jllb3tU3onMzH6Lcesk+Mk9GoGZrVBlXP3J5xUgEHk8SnqhzeNIdo9
vcWIK7SqEqQ/c3c5l63aKVZk6z0FCgHmGzRgOUB3Z+ZnkZ6IQDjYOAu0V8bNTwOP
eNopjQUaeFzsjpSJNUGBLqP5hmszUU5bmjLMhAOUA05Bay3q1svmFrDDSMbvB1MP
OEoD5iYWLTz2/1Yz+nprUsaVUyBQyA5gJ8ba7yVQbK9FAMQ9p5gHBxeSnU0fzJYY
QZn/D/leRFJluXunCCNaJBHyo6FAyMBn2UHHjNJxLxsulgZnfsCd3qDoIs9rnlx9
+GBzXlXIOcYdzkGYOna+8dOxR91H8LSauXwwmhRKtghiJBTDFuhCwnBhIvDDBNWF
1Z/SaarMaAeBnqyz2JfDvR34SfIdSS2W61JSIOUJtOHoesG7SB6mvir0/+TuIyl/
0dj8s0+9UftpimcYh3uy4A2w9Xr8Acj9sDbyJxA0m5LWfnDMqR2XsKPcqMD7jEX/
UXYJFv01tn6jWrzTLbL5M0ilzD+ZAkDqJLVWP8jd/KVVaorbDQpIwgk1MfM+xqoy
6Rtrcgk2RjOkY+vM+e8pOWaHLj2Q7iMhHh2r/r8RO9naUTaYxam27LsO5x2grk2P
Vae0VzyvGVM1f45E+vOS25XY5foRfLStIs8Cwp+INb5vX2QkJL+rs0DPrscSRnPD
/iuBV+rIM3DSaPHM0LNFbCN+nAtXzZRQ0zuJY7ugifsBxLDc5sk8BjEqOrw/D8Ha
AOtS+lzkJZBTes6eVAuZHMPRuVTF+LiuShUaxCAbaUZAmNuTUpbuU9nSTsUimIM5
ooQwjVBqrZXNh7+IZ/fBnOGpdlSSZgTBGi+zlF0uuaF8wUpLOYf8zexkA/OgkvCs
J6E0a8GZSYOnX73T12PWEfVrwhm7WD0SvajgOsfvgBMTlwMVu5ge38STryL/anTR
CCB4uqc8RYiEHq9oi20GsyK2B14awWQeDokZju5hwVo4l8ToNjGj58RRXh1mxhJS
ccXQjtGeVNLFUyXs6DD+UsP3DFlZpGKJWIdOUPRMTYFKJsrGq7vQqBF1+39v8fyf
xodZbSOrUmtfIloc4L8idw1gKwT0p4Y7akKkcgNaa4I0PfenkmBnP+4sHHyyCQte
lDzyQHYjeRogXxQmxuH4Tynb5bpdPkFFSo2f5E9B/TqlPXb847dzmFR0T7mZXByY
R4qjk7Ayohcvo9P97RkTwoofSMLZyhaHUyJYUp+ta/8LH1ODNtTiuo5No15TYz14
83G5jO+eBgyFGOyFk5tYd/2NJaNZvA42D/irpKSq8W9EiW5lXWaFmFszuRi+UqSc
cXMaHPf8iqXxcEVNUisviOPJDuqUQ11FYeM2MXzvOtUWu/JAlLGCPE1EiDAB2BiY
mwJ18FLecUvH8VR4wYK5ce6CxImEvY5VWB20OsySZ6kfkWzJLd1PCgqgrsfP6mul
5/bZRNs8sx1LgDgoPYpF+rW52kRdQcmnMFLP7b9SYi2+1P/VPqStbJuIbjaQ7IZx
0/iKWDdv99oXpbwITcfNYQ1rLVpsknN7tZ3Y5rKGmAvO15tG69OIv6YR+IadUGLL
ERNjQQ4Hx87sproq/JvqTEaC2xpNl/bbjfHa15CPHHh6N+R7DCkKeCyh/5HBkdlb
6gPMHLID0a4QxDCeOoy2Ljfie7UoJzQq6y73ew9auX9FTHwPLvJOSRumYwYVQUNg
imSaq1w10yDksGggcCgvK5+fcewh2/2keFnNf6aXGtUuar7ljZDApVQ71mO8oyZl
qSkqEPmBGgRL+qP1I4Q6OyCo+XJ0w5toIeCWxEKHk8tC64bjvSeK1CDr260RxyHy
Y7UKDBM1ARtQ/ugYbwAoBCIoHo2sYFg6dbkv0iofOHTGR1Lac0MCODkfJzVq19Rt
g6RmgxbgDrnTn5I/tfJn3aWakCHlEokXHGlaaF7hM8syqNtY5E+Zw8lSW02cu3Tz
4MiWRaZQCtARii8Bwk5e2vLKUSBz+ONuKkA9uwTkg/x9MzqX4z7Eamx9hrfzQycN
8SkyuAIQVhXd+9xLM5Mgg5GxyPit4YZRGfaaTY0VdQn9LyBgioFTOv0w1GPnC3b7
l3bv71HDAMLXNb6O9bXC3jG3PjY/Zw/oRqlq+SbS3kGLbKkFPX985vmreXpbzRUR
5Q0FD1K7BQPiJ3J5bQtyqmQ1muQnSCxN6CZhMkzMr01T+XJ4BvjsDwj0JgOgPTm8
M1BDMQFDdELFyWhI8mQjmffkSk6lkMJbeaqVFn+gucZCZRdsQcglKUrKTyIpawut
QYoWeQAhR+IGsilDVKCYqwPZB8FzBP0JjpElIi/b3rX2dJ7F5wz+Y+LnkQDhko3Z
Qgxjnxqb9sdpdOQkf8s1qkPEQwHslB+YyOPuJDLJsbju0zIyUC9BJC+l6TrzvrQN
4Ns/5dfTewJnsCIT+LdYGBUgn431kPOYJPbrTglth/JjXiiN7MHRgrvL6BE6EZt8
reDdsipyA+OyooIGTWW9UtGE3tImAkNvj4UhdblKkU4GOzSWkX7/Nxkuy0bS2Eek
ZE6JRwuFW0+KFVW8NfQEDBNrSHd32t3bUjs9LMCRO48R4YVnbGRiiQL3DQ2VWDU2
y1q0Fa+/wf2dtMVv0WmYklqoIYS3BGMGLix1CnpwP1Uv3qNZtMOeWEj0uxu0k8ba
hr2EB/QHBkm9jyl55RZgoAmS2tDVPIykzBhX+le1V2bGMrxrHylhViauxXJxjknp
qbB1QQnUm9r4T6LK/zhtf3SJeYCOKznm15LytDbbRoaprYx6t/X+lQF+dsuLMi4M
YRz0r4KhgD/J5gOA6EqQu+2HOz45+nSq/bOZOXiPqQBOjsyf6d5qq5PMDBwhEDnd
Wf+91FsC3fZo8+xS838z4bp5Cq8pBPTSthYPkFEgcmQp1KO7E4lOs6bUkCckbyJ/
Y70OIcFTgXTGieg/Fsiavrq/iuihelfEGP5LHTX9Mts=
`protect END_PROTECTED
