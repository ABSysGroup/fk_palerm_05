`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rEvcDD3Aqp0kaIQqUxuUKcaZplnQu3wugu00JQPl7yRTTxHb5qAug2d49EQV216z
Rz5RuHaOV/wMOBmFKT2kjb5JYvNxMyTodwL9IQo53m7oRDOptRgYekjZxEM4WKrk
OKI1Zj55CDzcLSSyZBNDxUwsp5t42gBGNYNrjtHfx9m31NwGE7zDwmkB+JpzKBDG
+kgRTGSDDCJrvQSBapRTpdzp3kgzNXnYuASS7Kve2TdQeUXx55aFE44pFM3pSeCS
QWcpQ0bkdNyUi3Xx0C3M7vDrP6erYRqFfGWGkgWdAL6Sv6IG7A1hiereNNOG9ucB
uAbj3C2eWGdcceqyCXviFCIMXnWkBF9HoChVX2jgX2JwatT991yhPdwOLyhgk7dM
tLyMNkg/vX7FfDpUXeTk3S5FMgY4v7s6jnxHLCspWavP9mLTzuC7k5t2U9IcBsxo
tz4EN6HzJJSO62ryRfp4QEqbC/INy7bvZoY5xv6heSUHhYyBnNiL10AxItqIoiD4
LMxk7W5a2YjvrQJCtSnn21z0X/rJbOVgf0KY9TkN7YvIwOHehOxeRlApNFinHD3S
eXM3vFsvbRHxB5zoLzmzuRQBYvhcnxPXUoVCPYdwWv3iQs8Wuwm4uD0HNkNXWUUj
jMWg4tvDMZwkO5aEjiOL4yqaiq9YQeOT3R1e62zqfeVIiuMsGyYe0YT0QxkYDZLS
jVXdxaO0YvHDL6L+/0R/V7rkPqgmfEnFs7M/hrvqtOujUfetKbdN2PRR94dL9ZZL
nFV8Gr33zFJEHrGaDkQjBRbxUrXbkEb1mPZhcCo7nmv+CEuY7T6OGhkkWpN5Psn9
HV3ExYPqz6SmxO6TXJcqCv8Z/Bs+F/Yy+xPn1cf2D336z3cQ9S2vyADycN3W4Nz9
jdtvtMHpk7JhNCw6OLL9xKP4y7/F+ZEgpb3tkYlLMxkjy/9nrkRxXng0JcmoGMmC
6mkfSVus2+mu/QIcVYjTxd43gFGECvCC6g3qt3aGOqbQDyS0hSSCj5+u+Wxpx2lE
nIW1Bs7lAfCUpC48Ws50K9Y4tbOo+fl/w9dHrPgZopkfAsLPDVJmRW2dyYhNVEn4
fbp8aV0ObWV0CWz8Ppi0FZp9Lb9eJ35ltIDG7qMfe2+KTEI2i6a0V/bPHhF0poes
k6jTq3LKsxF2qfY8E7s/g5pg0S0gip/u7e9FCaVBEZ9MW/z9M9cr4imtNIB6JePJ
UuipVp39PlzaD5BMUk7xV46gaQhjJvewBC9MsQ7IPm+GEIGuvIBR2gVq7l3kBZt/
W681xqIdLVznhSPCzYP2NXMZyUNwBNkR6pfgGrhlhNuZwWlBmiO+fWaLb9gE1WJM
OTrsN3Co/YtH+50EHZkEsQeJkCbJfa8QAiNlcpAeXaAKJ5g+ftBxiK+y4s5nfwSg
vZ+scQ68o/7Q8Wrm0fc2FXFguSe3JxPDVdqUf+onRyiOJh/AR77bowTdMJCxR8bP
kcb7IeqgI4b/gpxGdqBFGBEwT/wPjXW06zPWhYda8ZQX3mLIOg8ftGqKKAuFNVxw
gS4LDIxIeR7BFG6uq8/SnNfIKzLl3c0NIK9nvrIBLncjn/1n2oqN6d9Bjhocyeq0
X350o1hmN7srNDiByMJwvzAWCrQWBCXHge5r7sui4u6sXTSyI0kqTm9ZgiRy/Rvz
6POFbOV+uzCesq7xH3INeebjby3CFew5sQbxmqFTwbCgziWIeX0BBMVDDJJlZLj9
u91gk3W8qYY1+OFThtUMuUtxeO501nnmZmILTdpyJPGRIYminhuashlPnaNo8DSD
U4O9VogoGdqbubkd+4Ip7u+NHvNVx7SeaNgD2V/+zNDXie9Y9+BPFICLFvShtg7+
8j1nO0c9nuYJHkfd9LTDtR5lTmHiy9qBhRRL7qXUvwB4KNW/f2F4FskzcuZMa7rh
Ufewx2Nn7j8cwcMA0C6R2xArQnR8nXPKXPmEQQ7h/l/JkK//R1VrPZ/icVsmrsB7
4O92DNzYTQ/bvVFHCeZEIQmNG+YWukNekHB6QH1OTwkIAhB/LLBxihSYYfTlOI1o
mR93pBF8phNgODQ6Xf/wgd2IWIlXp06Gl1ptIfzVT85waMAbG9iKNo7m+I2726d9
XlaJaoFH40TTAoMVJA79yFkQ0sHuO4XAdEGI0GonFrAdcEEpdMRQ2CCzyddUNTrt
4DuPAMt/cVHIK1EoziftSp5jbbkACcY6VEyvLrkUSVqcc9prLgVAiwxbm05ZlDLX
DhnY98q4hmlOD8V4B4oHPu9lGkzHosUwsdqES5W2ZSvoI3OryJ1I49zX/Yd0zVJL
hOXFR1YYtlfyRdw3b4hPxeSGimky01RvhZ3Xy7ZwMD6bgX/LHW3D5fajuPgAS/BH
NR8Ldy6Ck0yK6j9nKvO2mbqrza1MwQkkaUdosy+Gh6Md3QQuE5C5/2BcHUvLusi3
s95FUnvRwKI3KROvt+LrY1dtNSsp/kw/3WygahUmGlAOfAkl0joqYS3AdGYYop5N
Ieog/Ry/Ub/MrqAPa5rbbneA6nhJSBcWPmQR+cY1BnnE99IuLElt9cMDh6hOJQWU
aX9lqUEIhb8Im07WWrE34fLTZSw0FqUtWwj9RmDg+DB4tbvzb5qBPIF+dy819orq
YCoT/zSXjav84/0onlEg9eBPXptlpLQL7Keyc8vrHKz149aZHt3bffh90/53FDaX
8NEbAqOxR9gyVVOXV6rtwb9GUk0DVqXCQQg/ni/qXzXfJUBnWNgLjmdquiMI1xGx
FsRi7qztNO3QT59vYY07ygnqDHoD1+dkZ+Hin4nql2xXShkuHJQ8vtShVPnFTJBV
/oHwynf3PasPgsjMnvd1QIUF3mqugIoE90kQjulQ1q8n3iQRjdFps4pujnQTZHA4
K1RDsUQdx9s7ZeFpWczB/63+DxDMYCGCEZ84nBePTkrxZn2Y4XmCoXdZA/T14p/l
+yQmSTyWccc8HaigkaG/Gk2AyTLcLhEt4KDL3Pj80CCqfK6XHA0YwE+0+ZLzrWCT
BzhMWklw/qw4IVI+7R4XHzyAyLzOAS5FroKB/rd3ebkaCtxrxK19SY/RiR74v8O3
kmTIYQiVDEEnXNuuA5ieB0nRbjEVKCq8t3r6YkUoTFA3gZQiLjvkCTUFligfzlOD
ToBTRYuELo4/x+a+GeVZi3Urx91f6sMSRTdBA550xpA1XAXkBzPHTfGfa8EOb26H
K/nSrY3FMUlPF9AcvjWl7U5mNv45GdQ/GXvG1YV0jSOsorC2bl5rITDT9zOvN+bH
gZXm7WdMFv4bCgseYi1nHDHiNjRlkmc3yI9q6EyDJ79INUakdlhOayfXxUrRiCj4
6jqBmQDaZAVvTT1wZGlOi9v3NLh8Iv1/qDHybo6+1vtgkTH4i5dkLxKcES6LWyME
VuJkGLR3oR5ahl8IEdaFQDdiDQV+D2uP9VhmCmMhiIcsNawFnwcv7IiyhxnkdwBH
dE6U+s18WJ69w3Yq+4YubuCgAfIfK0/zjfbk7QRX4tFUHWdeiQoftd0IxldMKf7W
4ysPlMh25b5YxPWyMAId9cryrgQWgMcaMjM4UarQK2m7ZJZfqlT4RAEqS/9NylNH
WWgo3dOCiFFvZZ5WyNmF8cvW2ozwp/90p6YWyV4o+2a3Xx3jXj4Ld71sh9LGe34/
XI17CnDUZoxGEyTB69EIIUYcIL5a5Wi26PbdsBAjKohmoykWFjyJH4ht0Mn6lqPb
HSCc58+21ERRJ/oJCIKNrAljcap+OhGw60g+JOFiMFLO2lJx45B+JCqStztH2ztq
Q+HGi46GoB+9OVZxgHav1pcUtPfbEe5phxFIS9tA7vXT8PxRkvzs/gD0xSN6E48O
wm9q5svsxKDMkeKpJmUYUFnMa+vrux2vGRsHhlG2qDYdYXBnYqfzZnYIrdQMvCqq
bd0kwnoVtE1Xd8ci582FSYxDB/yZd+rtXJ7L908atUrUo76vo+gSO4bptYPqbOnJ
9xtcZ5zeEXYB/PfZLr6T6o/bvZo8dADLVQi2biFte/LZIbwApR7HD8kePnED4T+w
UTu15u9sddButLi995LwMF2o4DbljJXcvviPaXykVZ43WT4VqNxrY9bRTOZRCma2
5LcArSHpWMr6wcoiESUk7/MpBu1iwdl+kyzdSEEX9PzJaToMB43v1+xhsSnXbghH
Xkf9SXBYOX/kEfbfXMjZRTcyw7fpSjH73yilP4Uw6dymNeeG90XUMzUCzrudP0Gp
IWmVRItkdncjtStot95+pOlHRvJrGd2OVssJk/kMMkZo5QjFlDpQPQFBHcyJublO
SpA4USC6qtE/f2XxD+vq9QUVnYtqpNAb4H7kwc1BNHqzdNPVlIifcntGypzh1xmB
PBLRWFuCFmGE8zAq2gpccCEpUdoMDM+CqnsdmV/0NzgSWGbtbCK/VOwOx3iJFvEM
gU9zqmdQ+U/RlruSxzZLZGZwE+n10lSvsKRF2dm5wPUm9jzoi/frHM5ZzW6somJ5
C5F64wWVs5GDUYIGnjF0t8PlKurs/5tj0H7d0EtkN4pTnUuPytL0IZoxD+1qvbUS
sYW1w6eH/5ZrxJ7v7HCLJSAhymD03M+ebDn+/cHDITkTi5ffTs+O5WjH3/QVcXwv
UpYTNcmQ5oB0BMWZtr8fEmEfDwh9xbu1eFSm8sD9Y7NnoDwXiyTJ+m2uSRIjArba
NNYV/pTF5LgELakVXX/BSDf+34hAHRFNgmUvgUHmW1OMILouid0RNeJ9xSANB9rf
GBx47lgY3hFYuueVMInB05UsYMW5nIoa5OV+r6gV8VNNMO8Emr0lc3a/7erskGZS
403fdgParFNJgZS6tX3DZ3F4+2qEnQZKiUggnX7aCNASQyuu7HjJ887m5mqFhxvx
RiF9wlWyDJcVrKjAhmtq4d/7C9AkGaesFjJfbJL9y0RTiEBijutR9h2W72PGbNyI
oFomvE5aAjErgRlIVcexMyOlREeIfOhmv+ez7XeJbbQbqVABR/6hPDDMQ+hXBHak
CYNI3ezFEAv3tB+K9PhBXm9HW0sINeCRxJE405V3Gnkdg93aj3uRw+tBG7NeIHJD
0Pr1CCAbPou+/kEWgMY07srq2OCLwws1I5l0+BT1HGYzh3ukPzMZvWxVw5S8qgiK
8UaKKoMsWYNCrs3u3gqiCdmB1SmP3yHDPnImRQSoemL9q11jp7a+Y7fyfiQzCj0x
gwqAmjAGXkq1nOTMihejh/7cKk+0rxVhRBFNIeobZQGCAGoOLm64keaKMSteiVna
mW0fTGwpIfyyeS7BzGmjax6bhh2x9Wrux4jA+hnBkdLEI5KshBSqKZWLIr0K+H5l
0KwZih4Kyc2i6MCDJrb98++5cosYKX2vaYF/aZ5khKXwL9NFufwZjAATW1RUHiGi
oeB3+968shhaAUpq7lN7QK/coFaAbkYfyCmaPbB5R6Yn/vsgNRPl209HpNj8aqtM
fFoQXkp225J/1k/oNo8Q9/PyNjxh7Y6zHwtHSZHbpGlffl5H2Rwg6bO812Thk2QQ
rDS1cFUOHgqkcLO9No8dt+g+QDMbUhSPu7Gs7rPO/Bau24cBFXQSps16qs58+xco
v4K0o8UtWAS0M4DQ8//jNTXpcTbuoxCnRdMSSGOeCNcM8ZbiaATLIVd8t+1iZz/L
bJdrQop+DIMV2wfss/Pk+GtDy/p1AK2nO5ch+3foJHKspreW+mSoIPFhJslNVYq2
UTdj0XEdhZ9FIhgFDVxcNYWEafell3QwHfpa39w1Bdejs70u4nKF3nS8d5v8oXEW
DrJ5YTl/1C4/MoNzAIswId+eJ+Cj1ys0KQFU8gFYCvj+PyH2wm8zTtgKpr4rWP6t
7erYokl8EE3qoQSxKMY00qubk/blylelbt6LGpvHMi47Zqu+l26aKaq3VJgOlO73
F3ZiciaEdlyfQYfWKauVe+DJmXsMyrcH6mrHWjib9vFm3vJeexaqR+/9rumQ+NMy
mQ1frE01ZU2YOWUY4P7jhNfNsLBaK1yqV1qYdGzawOcvRq6vDfajMaqnY1924bhN
Ie9wevTlR8x50cnB0f3AELf3TQgHY8dsxG0R5t8Qpfa0TLfn0uv79eZSZDIFJWjE
pGNx7Oo6+Ao/SmbrcBKqnI2jMCYCL5lvg/KKZeSqAXycIfA6gW+9Yo8jnnG4dk0r
9kUJKDUbGBZMu1QiSxs5AG+jQssx90HkqoYggRMxzsLn4n0iB9o/jQ1GZQ/ozezW
/OfZAHQIirOpRU4P1WRC/OwJyYbcMruiLxB+VRW6QSR17Hwif10Y/x7tfxmxX9/G
tHUdcDfVE36fndpB8UvLzL6aiJxSzYootYqkXqjYo8m70lYhQX0TZ/N+gTXbqICh
dWPXChHfAxII62avU4/rSHui10RHjDch57nQnBYBgUDn83Uk5ou6DhPTLJ6UmjXP
zNcyxJ4vaTczFdCmXbpgFWZSu0MvmiKeeUBLx5worAU1NuT692wS/+XfWFXJEy+A
Tbgct4bqyrqzX2acSk5LUfCAAdilfSYMPR2/DyTi/kE0ygldry4p+yPzdoJaZT5x
886AHUxU0xfIXL8mVpND0t8m1hFHqzs06JBkjaVvBlq5yUq5ypL/b8DZHxtedJhm
6yDGjoDVDYxE+LtdukqpLnDfRJVcYUVESxxNvaKO6BbPqmFE/Vx/76BZEEWSKWMZ
h9PKv4UXG3UGJIwTRx5UwlhU9Gor0do/ehC6PaPNawTikNO905DEa/dSL60Ti2NE
+TP9jYvn8329Xr79AqX+yMG3xy69yymfnXQe3+CmKiDTXYnluiVkaXITHDiq7Lx5
1fK/iDYygBqE3CdeIxXy2Ejzx0/Q+J+nEtr8eXXy8aO4ke9QcXpTHZkWyc5P3DKz
zyQ8gw0w+VX29Cpxzo22Tsl5eDDu26uGKpgqBbGdVxTnnSvnI3xiD/OZoaQE1IbU
AvudlX6cNkBQH+Dp0IjeLiiXqB11vU8bZxviXrHwa3IMmQL+4Fzylbdw7TUD0AWX
aT3AB+2KiU/QB2kxzAlA+E1VMannfvbsqc3LdP3caLzTEug38iN/zME2l9TNjG6Z
AaU13zsZtl6OTJLK4ZQ2EB1NEihITU9pU5Euz3vcz44BHLRYtOCX/om4SuTrAyE9
Iie8IoRkhbUkQG0NDRTN7eeTU3UtL/VX0DeYvowV8xR2WeglnrM+l3Tcna8NO9sR
qvqV557oHqy8/H/9TlC57qvhwniuwMTxAFSh01c5aO5YXEAxUJjRv2uYoJycIkWQ
MiTnt9XvtHhxRYpEEgzZNRi4+oBQOvMIKPt/F2Njwu056eS6bMvsvvIisn1qKxTA
k6V2xW+f1+EycEBVFLwYBhGXoOXfALhNgd/cqZ329WY32dQf/Q363iWdLa+0AcU0
VIIOJG4JtGk0QtYpc1wZDJVEAgE4+mcN97gzWReMhLUerqOUwLEmk7Fxha3lWKMp
Yx+WKZ6SHjCtk1sNLQnWDrudbByrTw+IeUikrUUEMBc9dFm76C71KR4iASvFC+ic
pxLxubxoLRODCV0ZJCGUFkQyMCVqwxGyfxyKUWD6z7I/XHVnBJ5rHDHMmrXNjVTB
ITRMy/uTEFP/ras25aU4HZojzioINgCMZyuL1KXixF7OO4ohW9piqV6hXWuFyx+T
oEG4r9LfpRbazeUQVxb+1W+2s9/7IrU1tE8VfldgZVwzinEnrPmmRD5Obv50NsTv
HN6s1/qeli2tLa4iUqdvit68CR6NkFdG1vM4FtavtLAEaExbIDrcmVp/V7wFwmSG
bpNmXUOUMGInXjcvkM3Pv1R2+fFiU4aSrWsUiI5R0bGUDXORBum03360PtZS4UP9
mfNFwFIQGZNa1kdisWpKPqiTT7KUV5W3kk4uXOnuJDFyy1xgDja3JH3qYr+FAqeU
jlESA1Er7dBB3ahDax1WZbnVShsr48656niuRyeLciG+E7epbYzLRFmsHIwpSXfJ
HPrdLzvhRbGxcE/6P4kk6fnn7BwofQImS0W49KEepWo8K3OBpNlQZWEqfNmugAxl
KTL40m3ssOKR7T7w377FfXKd0L4mCC8ipjqcU7INGZQuYMU/l+YEVaoXMnEGFrA/
Dwq8XXeIhZBf5h0OcZRtkpBZWDieUsTjRaaCGCPHngMMzYywDK8LuuE/0tcDL2iH
fHhtCFslp9A5alsmWvd/KX89IFM4q9+3zQSP9F79zKkJ/Slyylq8ePJhhs3ozHXq
l0UgHqp/jIkwuhur0JO4rs8C3gujTpRa0qa3pe8hX7d9F3W/TUaE8H3js/+Tzfks
Ahg6HQ1BLXvkPog8jiI4PDSJhMIEeNR2+HjWP5yuxXAV0OJmtVWKCkY2bgmA7BnY
dSdnvYpygIXKumETmZZiiZG7Q6KmZADli1AFmFlHa6ICvr5KtdXO+TlOTlswVJw7
PNf+ZVkfvgzKF4hSQGl7d43TSQ3NbsChQmkQxxB+OT28e1+pYuronU58pM/tCGoI
B2udOh525xV9lsCyT+Hw7wgrPrDYtT8D4S6XqZ6A3esSfrwXccmiXfsJJaDlOD1/
LOqJiuZuO5YEsH9V26xhj7Vqg9k2qcNdMra2prXsr9FfNrd+5b322IFgHzpo3t4F
uZUZeUTMQDaAOnPpBa+uoLOPETF7NQptIPkU9ClY/qdOnvrYHqVwyXtEUrGYcyiq
RjP3uj6KnfLxFYRaSEcMgwqvGSZQ86cEOzD7ddTjPuxmCTa1KvApBVI+HfHDF3Oh
2OE4q+WIoeoD//ghjH7I2Uhtt9Yk6xLGcMl0+FI701oTMuj4kL/SKHmsHgmTbQQT
1Q/roiPTllPlbIVZoyhK0OF6/YCPi8TmdwJDtS3ZqmuWfHt5S6uy99mjCP7vXdyB
SRznvOOtsWGTYRG20oYyAN8HBA61tOtwt0QihszI3pNrgjlfRYjBlbIloKwb+yXB
Hyi+a4DajCET3zkUTcrTZdeL3C5mJc+MTM8T3zeBDvO+iYvWIEYh1CeOi9gTlTFm
+IzniTPkXqvu2lyuQtxZg9YJvWLG/VY4jApiDZBEl+y1Gfe55AM6VRT2lDpOB15X
hje4VKjQeIFYFZEVQLNWk8OzH33YrmwQDjzkHtgo2sq0wsPBEGkm6vEbaPSGId4c
G8MbKnZU05LYypKSn5JBNfR/iIVd1/G7hed/YTn1Oo9H76ybhohbanN3nIiowI8A
PSLGOhROnwxusSDt/2GYbeCE8ph7UVKdMpCmF0xIRCXSTGb/qWTq2AGvNT35WlLC
Q8tsXAqKl9VQU9YoYOKJT6/H4RL5/DrXHOkFaFe7QUapCRdWObbgsnbmcxI3IstY
fd2zmpXXJHiPJhxEQ5NQ99vt/Zk57wUCAZV63PaiYI/pNW+1z68iwZ3Z6zeorXGU
U9wXePrWmyvoLi88ZE5BCxYqXMLE8YLrHvkgB1NZbbdSccqeHjrSmJZI/29GKXnv
4OIwnHZrZoHCTsbIYOyQbb10tzIx02oZqXKarQhTclTek++6DGxi+bWavqF1eJkE
Qv0rZ7nAdVEpUaUIDq8BQ5zFv0v9PU5sRjjqOHge9E+1PcOW0lbFObIf6xD9GN89
/88g1LgMNNLxmpGCciCZJI3mUDIDxUNaFmQo2CrK8lftD+o7C4efLPvdHG5t3wNl
bNGW3GubWxu/7AqLRkbIaAjHDUj0urNfuwmf8HZ63XfOq5fEIka88NHojO3vZUSO
C0Qtfs+YOHAiJI5L7jQAvQoOx1VcqY1EdifG3wtt5RahaLntXtj7sS1X42kSPxg1
c7IxT5NFFc1tjVq78br2imvWzhgzlF7AK4Y3D/FmD8YfPqd3OuYictCG1QNBjWzO
upai3J1mGMoCyDR1geVWGNvnNkfTb704pdw8cbHti6h5nkJ/FWwyic11zJHVGEkJ
ts0mZqBZeXhG79v6BlcZ8SjBRXcQM847fk0J6CbjHri/sbXLp/je8Ye4WMkILFGJ
dYMQ7ybt1P/kIeC4Qqd1t0gRzZ/Qh/avHyCHyHdBNfv1AxUqtYRP2eKxISL/jNR2
kHFhKWFMGuqR+BtijVgMBw==
`protect END_PROTECTED
