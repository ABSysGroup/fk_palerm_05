`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NStQf+TVjSnzLTKPT48Bp7hdswzY7e6DBFYvIIhwOsLzWejSdDhquiJ3DTbHZIYo
B/GfOlFKx8Kz9k1OfR2Gsk2gwWu+LZDIcmsg0cOiDn+G6hAE6VUnC0WIBj++UHtb
It0VB+LiBVSsCfEjgek74PcOwGkCJ8FDfagVvCwy65wdr7sDYyZ0WC7pDWeKahfy
TkxPWkLWL7fqrMDuOvifHRbbUldceOGzcvgShu2jYd/eMDZ80HTmgJhCSwZSRfVc
5G4lYJqjSvymxUKthZ7Kv+OUjTJ5J5JCNXahdcR4KvSJeoPJKKB3YHpZiV31aRO3
ov4Ycddto49FUbRvoO/D3U+lDv2e9m2W3zbYnmVxQWe0OcO9zDMxF0e7DWq8h/0e
aVqLFRHukdHwQlg6BGKxWFTO7VsPZ5V1ic/6Z2ScCOt06GE5LR1r4bfVYNWKcuLk
kcVBfmy91znYu9tCgaqrwhCIG9/+oNqHtgLHWgWeuHU81ym9/ERuTxnUon2vrrV7
PZvVoaYM9/VrJUxup/eUywY9fSeQRJ5hp1FJWampYfMh8+IKigtFUPF3maqz0Ir+
NJTqoM5q8CgJ1MmbRPWvkEqnb5xAapzyzs8BvoqsxsCH3ulEzfQe8oHcu6roWzJE
39l4Uqo7IIay2xTBdt/QU0MfaE4ALrXJL22MQyWIdetajUx1hlsWQZRWJIOaFXqO
z98O9qOY6o50Q2q6bB9CaF4nUpFDN204T1jCA1JAEt6Nchag1Y/PguIR+lACFv7p
nROi+I6FXjB4ZsGDwKTM1V+SHBhnwAG82I7/ewJ7A42hCZO0PW0m2ekaiglVXzNT
DNpRo9L5/F7a62VogbS31PHPhi6O9pVbVCu0pifXK6OqTo4eFDY7MCF8HgBdFhHg
XQkP7jDnukIX0kg2i1ItdroVijzK36JFy7/OmQrUCTxJjNmIpAZ+2diMW4hHceLl
bcy4gnVQawo6EhrCIcVBWl/gxdHG98BqLeaN6DF16ncPa2rH85Cvs02a7hYThiLe
32SdG+3pXMwzhCy14MTW9cU2mJ9e6u6rdN5aDaZz3tRzok70KzaR0fEZXW7/jt/k
I1iof9cxsoZhq8rjuAiwdQ==
`protect END_PROTECTED
