`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hPkv0qzAkg+I6SjvdzuibDoG6914GTY+/svJAsFEtSijGACOD7FpoO6EM6ssq4zF
NawUr4FshRJdklsSPkw9TiKFEiNAXwC36ABOpfR9uO4doJIQ3lpLhYAvKZkJznIY
/P1FfL+eks5ElQ5UEp9Ldsl2oYS694/UScH9dNkFKv8y6p7UbmLSVZTw9gmvBzf5
24ZWwXLMzcczEukyWAWXWY7zDxQ/fvQCjLOAEfuTZvC2Db0xcyTOTrraURMeiovr
0Aol7TuPWXjIwyg8H03UVQ==
`protect END_PROTECTED
