`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TmS5DUeQud126IxYgfWHn6d4aYE7zZ05bONF3YWhvNfN3Rq8lhbFejays3largba
bKI4+u3xVLsRuKjq4XmYMiDPBBcVrp9/DztLi5i8UlykYAsg/M12NlBGJxFkE6s6
OTp2JPGGASqsoVj/scVvgPs974bP1h3gCNWOUUFKXJJaZOwNjQ13JAxdmjfVHHAj
wBVMotNlgyx7yAy/vuVIUr6/+sLa59S2Y6pRebqmQg0Ouh8rqrKNzD9+TdytvfkO
mXgisGnizs8cvNPUgGmZtKPcvj8jN+izz3zAcZDwGIpK0y9s56YBCM4VbjTNr3ls
8/UaUQDWr0tizHX8k0a+AVpbw5zmw4iGRpodOIFlPXueO4Aj+JG5ibj0yprqGXti
kI0yzCgyORiBPWE0Pe5fJCzwmRxX/Ju60Vvl+SSPs6vaJ6gC3DTFAwRVuPOVQeLj
U1VWU2ICdXA3fJHU1R8zWMnPh+qEvtHGmzDboggH9oEguQ1gha8fUA1sBwJ0e4qZ
mAvH6rj2mRwrqKULiq3nfuQ3htZ0O/B+DFB3X4A31d1lcTOtu1FBWJi86nl8Gl0C
SYj8DCRMWzsmaCcoRrj32E48aENeONUew5Y8w6q8R3VKYT7iAztRt0btMEPLvCcw
WKnC08unKi0ExZtj58JD4hiC+LJNbK0RE1Bt7uPs3zeXQ0qpCFecysW999PHE4bU
jCe+wpb7YPlGx+QV4B0jmPZejR1QHIpPB+FnKqnVFAaZf0jqT4xHQejGDegtULZ1
RGS5sUHHe9MFqOyV4zogF9rfUyDPwbqC2HmADn0QTaY=
`protect END_PROTECTED
