`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1cmHQQV51jujTF6hsWP9JL/imsw4YSHj/gxM72NWK7DjQDgAmsKugKXoXjVM/Zv3
2515lAZPj2jaAeTb/FrMFac6bSumVqix8bA7d3PqK/lWHARbUpT4cxpttun7CWU3
NpA0ZXnpgikdLz8zpgZKGGKqkq6M40HwoCOasndD5C/0PjtfvsvkTsAnzgJHkgLi
8yktqSE7fgKJxEK798oK4f/LD7DDswmFmGkksQmStOnjI/yqs7aM25fW+F3ufVRz
2TIraeXKPY6VJ8DRzzRYe+w7yr5fCHhaxc8stBCPus4XUHVzAK8a68EF9xyEAWKw
gxbmwY82Lntyw0JHrYz8wVybpjFuDUcthH45GnQ8pmdOaATrBlS7ZTAbK8nxITQa
StkFAkq7COF0hTLhKW6FonEks+Ykc1GH8Y8Oas+bk69/aGorf0ILXE9HFMFwzprh
qiTCg3idcGLRrT2BuipyQzI9UnVo6ySeIw+3Pz7q8OFoC7MG+oyGIX7BMFG/SBg6
7fL/LWsDkDdcrKY5BrEMwsxh5hg1QHcmEGQHkfmUdr77u2sq8iwdFrF+P3i1TPm+
ElcErpT84y8OKBcCIS/jFYlZQ8+7K7G4OR8e430SbFx7dQnztn0+tDxXZnzFSM8n
oNrQxNq69F8Hg0Qr5D43jA==
`protect END_PROTECTED
