`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
chhEpkN6dikOmZvE537704AohFXB7qnYkgV5/vj07EEgjftiRb/w3GOD0yK/fWG2
GVBh2kScehKcDfrlJW1Hkp4q2kV89b3cpM8uMJjpwK8LlzWFtx8jch43HbEBlvlQ
dFMCGgRoa8LO6x/MSj0HhIiETtib8gL6/VxeLNoihMa1/fS4tse9abkCv1BbmLFk
KTcrMLahRgKlpPz/mIxJrE7Ahr4ucr4+HV2/FQzfCs8M7zFPW1P7FvIW9dJrNIif
JLzGAFN8orIESJ4hawXFARr7rNuU2q+EVia2O7cmOSrGbm5/Ep7VXU+AOneTXQXU
D+HRnyk6jm0NCA7vQtSuRiVX4mXLoU75plY+3i3qD4uMtsxEXZZNJPvhezZI6Q8G
mRV9spz8hHNndgo9jSc0y10lkaG33DJZ7AMwAHJ7MUFWpH6z3HjbTftajlbtPCh8
E6XO7n1QRDdJbVj6ZUnixkWP4fDqmVSFAjGSAAdoSicSPr3G6sA5VvCohGdfzh1Y
KIqAmd8Lp3mV1hDVM4Awmk6ZtQyY4zefqdgXhoDgg45Q5zpQl15OLKfxd4v9AL5e
UCp01SiQXewxQz547tpy6nSGLKOPA9RknS6vf4rRQiuD+nbDZLn22+7C5IXrrwbR
uwEDF6DZ1a+SDt6pAs4qVfy65YvkqYpU/4xxMdmppZ9gy0AZG/6JoFsy0xYxqxlN
`protect END_PROTECTED
