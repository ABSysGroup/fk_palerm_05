`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nAPmcUp83LPM079IUMJ5kCGKN8IbTL3Mc/qrKQLqnEOvHq8nre+6Y+BJxc9dyLSU
me6TRsX6HBxyJ7HQYrf8sjVHFdMTjWCZZrFoX5CiECxvtxYT35Bhzt006+UkCKOd
FudSUbQstwe6Wj1TkDWb013oATlWRB1eGoAK5ZwhkwuFQBHJAcQWyZ3eNgqW9eaD
y/7L5DB5T3gtq0/wNeSNZO8qVe86h6XdG+3DWummiT7YrqVN9wg4PeX4pLjX3GnM
5U9mpVA/HcP5W4QjgppRyg==
`protect END_PROTECTED
