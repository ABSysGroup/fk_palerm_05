`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x1q2x60WgMaM39S4dljI337/our+0R20gMZFHcnO5WVJlbbny0SSwK0skkBRvYFz
n8C+3vY5ycFShVAWNgxMqHnSZN4xVmu5BKChKWSCaGC02mPNR3aB55IMjH/XTsRN
/Hg/SMzD3+UVT8Wa1HYpZXwklfK5LMNaSGKGVe3jsXzvEGNAj34iw7KKTYc/ygI3
w637xFA8k7Rw+Y/Llcq1tKExPyXTZXYY8o7iew86E3Cfju6kcL5ZKEhWY4yi9Kz2
SCViwKeeX2gWDK95A7z6dgGfxQtCrQFU86beIlfZDBnUsAhohcOqDiVWuttejhSj
8kPYwZw3dOOCTD8XYSEeng==
`protect END_PROTECTED
