`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L7BU+IUikUPhQnfDjT4U4PrMmsRKYIF+k/nJnvmZQ9mU8SwBszAufcMzhNXotuPb
ve3xMlejJdz1ZR6XoW+o3M9EpN7AAfwZlDsdSCfcRkhG5ppWyttswdcc7gUukStz
+JLM+d2+fnJ1ZNaydYA15gddExTIGuA3IUqYy3JVYGgnXe/+WNce3SGuOWMVvWE+
fsCCxlYun9xN0mfFY/i14xotzI9isFkX7sV5bInawE/PKciRT1XGadia2KlFn6op
`protect END_PROTECTED
