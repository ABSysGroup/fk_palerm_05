`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kIC3l9eC3Dgo4o9eshVXuvVCef1OkqYzRbHxA2MfQ5Ys4HFhX2rgrX10ItyVvjT1
UfBY56QrPZ96xCZlWvP5n7Ds7/XyzC/cokeuR4D9tdhhMe1P1LSuV7mYxow+3V6z
KPb4NDi3GxeCXZ6m4NdoUboPjqT79zmpCBf4obn+1jQv+S9NwQBusUjamGfkjvpd
ZFGeo1WFfEoEe8xbGAHocrX7Y/r3VVADXm05ubhU4akPwGv3mluQE2UaHl6WIWiY
BK7AuQkHanst5la8KzyApWX+JWKCkXS9G+cXENGbkrUDMs2nmGaLlyb1FGb2aGTg
elwR4ZN29HaODk08LUSofeOBv7IwleSZkl/gKMIVlVK6xzl3dMuQ2RNW35dAV22b
lflqvzdR6ET+k4AjAKdJFW7O4vHrKjsxtF3sANDXVgqcLYmiZ/z/unjGH6bcD+gP
yGqPFCpZspuAAsdZhO3DWCigskIFl0CVJ61G/aV2XgdHyFl40ZPesm3HkwQxFIWW
z2GilakQx9amfUmoqyDK+oRtJtl6GoktfJqoKZrY5Ew8AqTk78alZJtYngdceR2N
MJqsqjLDmTD9wKcWVUdbguAKidSLFHaxG/bWnkDc3jfYooBjEaxn1T+QYqB8RUh7
cHuO+QDKd/9u/Loc4oVIwHN6nimZaX4IXU0875tWTTw6aRh4uT8NPE6Oy9qzW6OA
GXUxya6aOZ9ptnMJ16DrPXn6gGKZMXU8lctBAe/w1pIFcHAgMuzfBInMYNiEwcEl
ZuYwEh2M0Lti6oAX2lWerg==
`protect END_PROTECTED
