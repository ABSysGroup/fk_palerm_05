`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bBegNYQ+h2tCmQpKiliY3E8Mc4Hf9jW9cPqiGwx9vjug4hjsQwNcrbN5vuAa5A8n
VNnfIVwx8ipsFQhqtHzDbZKYNXd7cGoQWhbZcVjy4CE9dwRZgD2RNIocQ+HkGdV/
TbMl3YrrbZe0L/QTEvI3TyJTNnUz3diaZjQj2K0w/7HOJHvS+yIzX8/hJpzt1NMN
khnrONdn//XOOfB02PpIzRKeu9zUxbMPioa9xjq2oSf/1PMVPNg35lgxry6FOvT+
JIsqokPudIQHdnPT/fPP3FszwYl3pEp3bt5WRpKbqJT60c526TceyKuuOaqraEYg
MZGb+7JdjW0zWj4n1/P7LdmgGxf7fTTI5Ly+6oJS+fmUcScHeTOhFXh+lEAs5yFf
lES9BYbpwwW87dXBZe0Gu5QTrgTK1o8MPLSNEn1kORujic91qggBDBm/l2K2eZSi
yHB7zEsybvonf+wjDlrHuFdbL9ThR6kERTJsbwXC7+Xa4qpKq4sexRfer5A0SI9Z
23pDwwItfjTfoorjIn5nvhCQl/0IP7ZAsb9FAueTafL/UYuCMTbqSYLvEueLhbf9
VMy6eoOEcyRhRoEoBQ9bsO9Mam/NxIr5fcReSyUwAnI95QDvMbYlJCFwcKu0c9j/
EgW0CTKwSBbG1FwP/cFPiVclKiwJ/jDHtKBtrbt5yY170yn5pQ7ghf6vN2qH9U7F
tfuaMtcYU0+nLJTtj6SGlRcL9cR9ExHbC+UbTNMqq8/NyCBocV9sOITXA6hwjuE9
QIu1CLMUL+wz7O5true84bNWngAGqadm4G1MxcUrXhQ1ZQ3+CuIbGMbyDfgO6Yjz
aGf9CDKBsfRIYOaTy7H46LeGOd9YgRhbBDqHPQAcF1HnX2eK0c8AJyqqD/W4J/Kd
CZ8XQJkBS2RFAcuKBThv1EUAqghU1jJ/G8ZK++sGkmiF0ewoJl+7N+6dFS5jmhgm
RMkc5FKpO3W6LPVnXEXaN4mePqO1n1udFwnpdFzlRxkIy8DkA6Gl1j+/DHxXQ1Us
OP9v4r8cE8QBzUX+r56ykuhD0fOX3tGOYYNOrZyjtqg9fLJT9X4ZFUbz0Zz7h2sc
vnp3T1CDR87IKfCCzhLxqMqJBZ+/HMdfyukSv5Lc9DkVG6bwLlx/NJRrdMZAopBC
1dYXIZiIxDzuB6vQM4brrdF0DNBZgWhnoZVCjIxVlRbWTH49C124D0lYE9Jk7/Li
k5quZFHU2qFqunGyEnfyqpKOiXqI1sEQ5LcqQpVyz0tOJHDlgFm/ijcS2J8banvH
UsXlq4OhN5q/pUIDmtkf2nD5G8tFBpr2ZCJJDkJDy/dPT8wDdcNf8DaUX0onAt/B
1+2aRO6LB/9+dhE2349f0P0yKk7A7+wHVrqCAzr3RcJBlaGIfZhZD0bi8J11XzrM
FVv6TDf6kP5RRt8DZJY8w1eLpCM/tK52grEipLA+ZgkSv574BTUETvF/gsdY+wa9
UWo/PIo9wr55/8rCewQbTgIN+RdUDPf14/O3KzWZG688mXopzZAiGyiTaSLWxhUb
DkE4aQJGTCQqCYdSnjAaV2XvQFUiZcwxETI0y/birP1jRweN7bxmF9jLx8Aguhpc
EE0MsWtHlNQ6ALMpCeZtHVY2EvHpXLVSl+aX8bfCJPzd56/BmckdNLnNe4g2sHwH
z26f4rvcIcH5JHpsi3igM/Mwtr37UB8ZK0Rj/+pvyvZ0XT7HRtwTmXl+U33h/rKl
PKx2FMouKYVRl5o7uw+CgYxqOLACLw3CfLNLxj1V4Hx7WxC1rWqJ7V0Hlxf/hqkS
e5d+FQWUpcJ0b049yDNx+To5Y59XK1SuH8ifzuVyrjQftnws2l9Fepdn3HObS3ne
3qnFUgWVgofB6oBgbRSEfO+rh1wTzILWswqjKoA0BVD7w5umEvfF5Sp8N8dAxDSz
vCNIZtsmdZWhhPtyWeDBziLuoVGw5eai5uq4klB8UYUzsyjkfyucfOfsGTQLyV1a
mklmJ5/lNhhxlR5IHNJrfr1eJ6yRorvcC66c4kTSYz2wmGB65Y/IRcMpwxN6s/EP
65hhcSYuupwtGt5YutHUxcisHwEtyJIPK/yJvHf3kLh6yu4jsL7e+McilPYXgd5U
jyOYdVukIo32jx/AKXf8Ff250sjIxRYUJ8sxidUbwwUw1HOIpXBNUSeMYA/Vt0Ze
EBAdEHZszXEtKuS74l59UflE0yf+LeIkE38EQ37uLa5t9BTNTqZxsC5audj3oJ0K
Zu51Aoa3nBhCv4y0htMj8kKDrOgbfqZQjA4mqT+JOUeOLkRVTgl9Lrc47E1h3KE6
OXUpCd7Kj7Ym7oH3BFFxUeM83e6TefCtSkkrt3e6E+nt0aY2+vcIIHrjusvaWoSG
M1pV1pqPKv1cjDTvlKezc5WlMygmwgdBuQII/9aT1tEoljb5d6o9qms55jVFvOxF
IQ5LMlcUX6BvBIE5LzVrr+m692h4AhbId9w6fCf82albuYPSpGddO6ROJjTDlyMe
IqT79FHhuG3qsRKXagobj20COiyMm9cJz3+2zK84aIAxGFWV/2hA5+ctu4GMZZap
hckidFnkK0sB8YP1H+EOUyvJyF/jB81cbS+0a/nBpXmuqFaciIBI+Rusm1lGIBO8
zySRfV/K9DHjN6IXdwo3yRiz/heR/w4g5JAfKG36tpE18+Cwp9V2LIf9IelFGekT
TmL9EDDCKasAJUbiebU3rJWeLufrQdOahnFVKp7/t8KkH/sHpovC6cqfZe3psFIX
2B+N0p3vCyD4wZW9wFITCrB4PmKsikyNyrKBjoireAywhY8N+qBIAF+Bfy7ff5E4
3UDv5mGL8NwGunFeUhgsnxlY75pvBwd7g36jH96pxEiisYmHRtyWJY5Z2QUNnJpN
km+6bPyMGacug4krF/dNPSHFMgqHpvAs1a837ihqh3Y2do6fRozBMUhraCu+jeQb
tNmKYeqQDd9IGq08gK90yvTl4oq8lPm7N0iSKa7KI++8WYnpgyPLMyfgmiarBLXG
yuau6cfG0b3WHqsiB1D50pDPOdUyl9LgwiflSuIsSrXSSPlB2c6xQw19rhSfy7iH
nguLHlgcNt/DcQLTgqBk+Czq0DlnIOzJKmXaWhEuYxTF5XGADeRUMp45+HzLP52x
ak2+KkMplr2PKgYt3j7VkAvoT/X7bdq/fSLakUrRfoJlUMG5IGc0AK9R5jSEOlTj
5bJNdY/Z5N0TDh6fycvV2vLMuJOzQH2ez3PniwtqwO1S0MIvoa3AEcBIWB6QD57k
9g/ZAc1gErt+2M/4Jfeyre7/iWQgJQi2wYcdcuOSZB3KkXVqsaCqtswol3un5VjB
qtggZNE217X28vDNcgZHj4Qve9wSJSVBxXoDuiRVYscsKkrQGTDrG1PJGiIZ79MU
b1nzCkOlYLoytOLWQLf8NQ==
`protect END_PROTECTED
