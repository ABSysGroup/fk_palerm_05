`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nlji+c9M6c8QRjNxJUhLJj2dSYpkKSCLtga5o9sF3kMJNYfMoRHCY0S+zEgMPaRe
UwzjvPce6whhnVszGbAwgoGuPnPiN4o3Si9GSm/gQ+Gv2YP7FaSPn5UJwpFaj9jA
952vnNUgMy0la9V23n/fmHZYLcEQA99KF6p9FnU4ZT/HZF7TVkH5BZlK/dfn0JZQ
xz2PcHxr/tGgNOmf7Co+DlRjm9cqbNN9vfg5a8LL4AQMI4fhXO4xx07r7+fnGZwG
Jw55bSSl/HlALDW9YSk1MPF/fbI+zt3+KhY4YNoUe3cXI+dzxHEiDN/+dCp6QiBx
7cQMLY2QB+uoa3D89gFbSvZ6UmnUamXOSnykRM5yyCrUwVVs6OvevNIP+mObOZ1i
V9rxLBQ8G4hOF1jWzaQAogKs3oZyP5Zj9l5vREBeNswBO2Yz42428wtF5ysSIzdq
M2YwKO4PKZ9lUGi+J8oC4wWFjhVvmvfxi0MsPzOWOBN+tsUuVD6fZDXIHzeGI4vZ
4TtkmYdbtY99c5BAtlEeH6NMrZKICpKBs0/4V4t+I3LEeaoIrfxLb80/H8Kn7ZlE
TiP1cmuG8aYDZCECPMFDv2Vd8f6JfPlLV4R9dDrMEUXS//ngAOxIqeSXaANmXiNW
pQRY1OL0pJpwM9wOliQsePaezWYiE3KbATUA8jWEYgb5GkjYb4HWQ5+BR2+1Ren7
azxZAFunbJh9c/MBsEa6jAoJNCIetbG9fkWieAN0LI3KtSYnA0OubDTwI/XD1VBu
88Rk4TESAHj+7fe/ASBbHwJ7A5qZrtgX1X/A5Ir7d3Pf1AuBi8rjhuqPwxjXUDiF
LBBDT+gvyY6tLGDQm799P2tIYyGTZOdXGaU45hNXshbZKbA2HqdEU9eZNs/fDz+f
cuyPiwQ2XABN2vGN4t1JMyGf0QJN+yiW0xmzZG/kc1qz+1DDYhGgW0PyZy+K372G
eQ9zshIlI8JYhlO1kKBQ2KDu0jaQXnHGAPoY33e8+r0E5zlLHxkH1Ax/nW8YYela
7FODlfXBy0xhXZfMLom4A9wwz65WSJIynEItYLqBS/PEdlKJWmkrNMtu4vB9HSsg
DABxCABOtpEFWTiqpz98EO7OvMXrWvk4cROBTJZPql4HvonNq56WsjubQYp2fKdQ
d/0GXtgmm8RLO9c0FyVjZzsv0zvpiwZCKyzopqZJ9XTOJPZZhrrvfcy7+zPqhhbp
kYCnQJxAkhI+Xbvfwki2MFqmzr2ROeNrU9RAQAd5BPcHm7ekROc+jb/8hROGB5Ed
8Y2PBWSE01+Bkvm3qwZ1CkCVibhwF2CKdhp5z7pBeoueE466Ek4IYM9Q23mu+f5M
KcPyyzdCZ9B2dT2PYFa8iN0/zPn9rM5PFdNYWrFnABIsSxcalRi73e7f7kpHWlqr
gbwFtPGNJsBvoEhVcoIB6LAWcCVYv6WrdZqsBW+hPSFYzBduX3eyrLRcv//JCARO
oG3CH/gWAXp5OJ7iW74Fb66IHr3N0H0hKyptCXLmVQYrK3T+gpSlYPCCLLd7o2A+
zripsLYQgjxGrYrgFWXWTGsSyauIXKrnQpzi+I7YI2yrBZ1/hClBuJnn9gnaIMDv
xzKGZj31gT611xPwZ+VwYuZ4xWv7yOgI2ogjCHDcS+Jl2sZezzGJeY0SDpk6quDG
ZFB+RJBD5pH+ExL1nHqj0MsZFS04dcbhKmZuzWhlJwduHOWiR8JvEW24k/Fntu3O
Icgy8jMtidI0b1a6J4Vjk+nU4B25gtc3J7n2WeC5BCPfpP99w/H4mqVnJy0xiphk
vk2wMbngDUtHPqa8QQgWFO0iN2s1DyaKUjZleD56h0Vhf/vrEfqnlbDOdJV0/yzS
NTxf2bI7YlsGxlS91hEZw+C7/Lgcz1ELKiM55wCC1qGiel8ngKNXM+sfrY2QX7iU
09anz92LdyiSk2tNBAHfqXMG/QtTsKStoznHRkbqZiFD6qGNRUcX/bZb1gofE7H3
+rXG3LCYcPIZWswexD4igeNLR6mpjvwfZXJkioNgcA7VmUAF2phnC0Lsu8bB3tyS
JvR3tzlUP2FP7eDU012ozvtGbf28EoGYpsUtOfG4Pc4e+ZLpujg2CDhpR1Mtztj6
k1WbJE3Hp9lOWL0SdwrXitBdLu5bkNvidga5AqQjtaX95za3XkquUFoeOrvJTCH8
uTMR3nYjjBq0xlNgtUbAibI9XSCI9Wy3gF5reMl92K+CCR6sv5oITTQ/T6ZC5Zwj
KD2DEQLC7TRSho6J8Ui9m/SmwjnsxD0cfErPEWxcgxU=
`protect END_PROTECTED
