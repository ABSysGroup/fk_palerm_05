`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PObJfidgwfDKsFaHBydC17oaD7nAbZekUWwgEV798BAet7WDw5Ik+K977ns0A8W8
7tM7AvmSshGTjSAoW4r/30DNc4lsibdvIFnLpxusE3K1CSKafY03AgcIXdlUOEXF
0/hM21iPVo8HJzmCKvMvSytmh/fFYSYTb7SsrGCNsEXYSrW9a6CVki4CDsiTX733
kyJz706LlMdA7yI6BjUeHuR+UqjHCNIxq9U0UNvYDVqnZSTwwD4QtPc/Z3Sm1soV
a8N/z6hNLCWCyjIbWVbB1JKBDFxthzRgfHUJJHKfQBY2v5a4tKh011f25B1ocivX
gf6Kj1BDtb+cnSbWCMMack5CaYr9f5LQE0D3bcK8e3O49A9MH34tOZRw1P/m83Kq
xIoajVmJeC63KVXNkaen9WmoXvAP2ct2i3OYCkBospuvxhTHTV2mrvlDkehd8XU+
`protect END_PROTECTED
