`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Idv2IjLHOXXyWfhrH92Jdtt1G1E6nUY5oI8fpuVLORUqj6pVERZ1pPUScwLO+j0w
FeAsDNTJW77uAjSPuVyyWkGjATQibAkTkNp2Qy1rGcroNHFrngaAdXXb/YnUJdlS
2I0vkmYUaRBlqL0KksawCcHb+hNwT2WiGdabT04dH44JR4db9BNdTR+C4nbhfXPE
LG6PpSkv+wchwIPQclvg3AT8o26TSbgX7oanIJ7oQ3l3MJkRcN8XPKbVyjadN0jR
0eFh8yWyKVAcZm04AoaQg0fheyAFvFSO0nTf6zaafl2awCzJAB53amKjJfOVVVwN
VFu5LhVb6KLNo7beqozVO11uCy9dXe2aW5K6v6AcnBz+HvXRu6NE5CgYktpJkIpl
etZj7z0PNNI56gOyJa2T0oc4fhOLXCgbEGwi3ZXrMYtouND6scwh0hHFq7rV7yZ/
3ekrVkp5TLlUw24jNziFQYm4N6aqogwdsexylXQhxsl9lV/Ay9SWQ7lRAVu8eb5m
arRoSjG469+xgrFZrsAvYXLQl4ZNOubf1uBRvh1dYNE=
`protect END_PROTECTED
