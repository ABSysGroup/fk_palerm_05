`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9e/iXVVFqnPiWJkVFp1HS16p/rDnDV2k38a4ZBMy2FnnsPM0GZWwrfVrIliGuezh
IOo+4DM4++Dp2jtQ50N8UbVxk3EHWUMlCsXb/YgOQvxLiAGWgWSVAHgleZu5fzue
a4uBCu0J7SdjVojkA/wT/5SvkNA3mbXUXu4yurTrhRxddTwjOUAEC5V7F3YApC7q
+Mj2SxwTkUAKFRJwPNLqRFwxvL2RdIRmYsibBwsZxi9CLYWtDHbi46d8crwB56Xo
NYOl60KDQn11GTtAPbHhTx/kxl6na6b6LCw5vA1W/croddgMoN4HY3UFbF74bqeC
0YNh0x7ZNsvq/6dpTCSFBu88p1GY/oqObDOT5+JTI1SeRe7BrCb3FKzpa0pTqoU4
vwrLtA4ZQGdRtyXbLZRhbA==
`protect END_PROTECTED
