`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/16ZZnk2CeyEJ6vouqRqHZH4n4+gOzrY1+gJE9btBTHfo/XakmrhNf9Ft8nCIzyr
GmecFs2Dhb8JC2Hq6lhBhgfHbGZhaxvGrWjVBD3Ys/t9rJ0lp8CRZsluSodp5Nbr
P4tyUSMmDAu0j+VoSHm1NKm7UvGAFiIyrPHHlnTDyoiJs+jll1BaiNNrkVJanq29
ottW47OHfN3UquUesigRki02isXnRzGMBfHiOOzqvDzuT2vgLVwm90wilKtOcmmm
OvnLLLNdrWFWw1uCgl66G6fB5bO0xEp+3iL5//9Qv9PsRk+meAgv5uTU71a1svbw
uJR16ZDShLuPO5nv+VmODz7SGrqXpAGK2aH3u6JcYn/CJHLyDBe5pWZv20l2euoz
GX1j6SF6wETy6n6PDc+I/ebu/zdggsIS2oBB86iYPxM8j3iHuBS32JGJ94CZBiCc
Saecw70CP19YvPjrJj7EsK+1jQhr+x1uCnRmKYOO1O/QPOIoae7lz6qqOeQiJVVV
SzsS8s4IlfLCSA91qCuAE3Vq3w8stmLmVU6pajz39Q9scf+Qzke38cyE/c7eABUD
D/WHvHUfaMaf8cIO2qB3e6bXJNMVDbw6JdVqygvfwKBDvxoZwk3jniYa/8ncb0TC
`protect END_PROTECTED
