`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K9rFWtCN1ZXKMqz2DhkFxn4FY7Vf35bCev+P/Aa3YkiQzAj3QIMo2wLlMzrPYSdq
KFHQDB8qwGhNLYhXcJerqDe0isaBF7mJUGaTKf3+tGEhCXuQRuz/Cey1xYV8LDrI
9M5Gd+IpTsYIttEYE1f8v87HTEITQjE6uXy/zKuI2qWkGjXVHTnhMctjgTZjnEha
Y9cQ0+Pc+uXoENR9NSYNzGlhBAfHR9mTzhlObn+nRyKG0k6D9YeJKNV8gLQ67qi/
yxgePZ5tlewpGbM3qmGSOKA4CCaDyOWKLciQn34MvnQQAek831BZ0+h2qn5VUMpe
CFB+xvYQ/nvvRr3rvTW67g==
`protect END_PROTECTED
