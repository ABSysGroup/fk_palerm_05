`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sbelEGhlyWAGSgKbuBNU7qX4Db7UjKfnJxoIXA6SmuvXvMQ6Soob629jhseB3rmF
P+Bs/QMNYZ+71sdF4P7r9ngRDACYtgwerhJvPBvYO74dMRKuvgVcXY3k7KWTUAEw
t2kOVDanA9a4IEBz4MBIqSnNbbvmfigvtddz5Ru1FOmKZwpCvtc+g5DbatzkeQBg
bLmSJsdY0GMdLDMThuWWukyVc2RxDrNHLEDIRS/rSOCThfXG5wgI5iKP9DpDxBW3
k9R19ddoMRpXfIGwCHXn/uRI8ymFlNYFbAs3cvCFndFxxFGSQeXZrURZaS0vdSiF
YadacEtzLL3WcO98q/uTvIfWY5XCvOdqPj89nxDNALTQX/wTTmUaS/QYmsJsqK73
R1M2ZODgQAtW/sC/QRVar7Kv0Dy2X64ANHjekOubHFCoUggZEfzkPAUM1VZBQoTu
UKMH3NiVRlgiMAM+mlJmtGy8wd13ImB/U45LIAv5iETg6AwVJdKbOStMC0h1AGoD
B/j5aCtFh84vyjQ3Q7TzkSiOlN7DX/edFq8ea3qKoyT2XU/jcY7Xo/0Zrlxuzko3
hJX7oJfqicilDR/cOc0eOe87U/UWrsVXDrcndgNctkZLe/JUX8X3eysuq0s4dGcF
0sodnWrWtDu82D5GrIHcvN1R21VSndQr2dKR4+HhZcc=
`protect END_PROTECTED
