`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pkEi37unc/R5NYeaxki1NmYmu5oXwfYPRVvh4iZ+Q+o0IoOaFTHX3lV0P7jZeGJj
RWEdSYM/Y9LTBc7GjmcoXRdn58VkxAKTIycoCodGzh7lQrsJ3Y/QVEtKeeyfUrlg
sub2B/DdnvJpIrBKF63Oq+bNJjtiK/TQtadT+fUsx6GSE85isyBs9C9KT5B4CRZh
/eswQ4z+fewkEUmeiIje5n7zXDLvcnAGcjz8+RxonK830vVPHUK0lSMoskvVdkCv
78crka+LG7OjjHpypDyXPKvxZjMc1WWPVOIUkNFU5xQAUqbUzse4cHuvSWKedsv3
pxPyu/QuzQuZSr10mzheG8IPmZE4RMKeD9pS6gIb2ziWGoCNAJNjpWHyliFL1VZi
JvufL0VlsQ/Zzm3xk332Wdvg5BWppI42M1Nuz5FID14+VAn1m38IiD0pflWnrRqJ
yVlfLJ5KEqfKxgwwqUIBWT3ANfSSQCAcyiMHvBkfTCchmPpEsq/Wtf5osB9B0MIa
N6gCTcuHZryA2S3YY8qETcQ2kfO+fuhByndLLGlZDa1K31Jq6ysqDcVSQwBCK30K
5Fjv3UbA0oFzgDA6cTcDXF38nFFY1+6zXD8EEJ9esTIbGm1kF4aUV+7Rq5+vorlM
KooHuvZUny3RZupV0dmCMn9PIOuhGjXqVXTYQ+E9csFRQG8e+WpN/BlB9UW1pKUw
`protect END_PROTECTED
