`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vqTcJbj7yqPcVibs80RvTgKKm9ztkCCIkcq4JPS73TGHrqtHwDuI5CwwEL+Y1TNY
xS48zteERLP+QfdqAGv6BtO7vVXqCMk+Y6DJlQCQgIeryMG4cygdLxJuTQ8Gu6KO
ag338upErMyMRj8BRBFf73di4OyOQ85jiKen3X8J1l13Qzy98mAo7VS3c3QBxxDE
VJ0xy/XkRool+pCi3jmL7t9rd5xAw1fqxnkGyn5BTb9st+zWXVplh1AM4+jS9qDT
3xXiAuBuWF+otMr9g1nYXJt4xRhcucAMynMQNkpCvBCc2Ad2WZyuZZ5wrFPFGGgi
URAM5E4CCp3Q5l6jB2fMZQ==
`protect END_PROTECTED
