`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dxpHx003SZ07k1xOLIINTJb907nwfHCq24rrJUwJa8ZY//Jr89G0Rh/h3GBGEoHr
VwRAOCEBgtURzuGrl+/qqU0FJtR+joH+vKwfMtTJxXa3ROALKdO3RbJFy/HlIRE0
X8FeyYQB7HPxWcTGzxZrEIE8A9jmo+FabYqfGR68oBBvX+w7zdnAJJ4uZEJUGVAd
m3vfpa7spUUZEbrEZbMAxfyxAPffJPiTom7KRddtbbEb8yOebi0FoElqWxaZ+jtj
77vrfmwff6VSMAk8XDJ/UcKo22m3AJlDL4RH6/9bxVD6sqEQ7+YMZ/D9Xohyh3VW
xhEXbgZ+EhFQJQh3guAYStGcvAUAGYIkjiSsWaEc5KjASDEJ4apEmxhEIozWjlSR
kbG/5AKdipIMW7UxcShkHF/QUJJgzvf2rPEPldWt1qo5AHl5RHYS2PPbkauTBnWl
LcfdQgfKNeidzHAcqGok+dbPv8TxOhaAyz4SrQ+P/BU1jQDDMpS/o351xBxybZaS
8TKYw9/aP7zxjvY65BiHCsB/wvThaSEM6EshvKvcEZ9awCaf3RCsY+QnhqxR/Ifz
EOItgqnPj3F9MVsOkNBl15HIgkci1MWFDcq5Tt3A3M7LK3BXJWhG12vg48mPln6M
57UvJbNgdT8j+IWNcZEQKVd58a7DfVq9qjcjcTwFbHnYbOgSn3cU/BaK3vTNbrjP
BnKavA9FUJd2u7fFX3vTb7HONVsa5SZhnzUF8CYtECszwYR9cfCz7YUw40aQpXv+
hvdS+m10GZjkCO/HpLkr1ZtVqZ34/6Yp2EnXyvRuLLvJy1H9se8hahHHIkkCVPvp
07fS6NTqqJLsF98rr1fCMUA+JuPZKS/XgcaH0jVnujcVPQjinWRg0M1U1zGjTx4Y
WN6JpEagkNokHtDdVZ5auDoMxnEOaRVZ4P4K/xd3LNjwd7obZK7O//rDo7pigONT
bRrl6w9HG03+Fq80g3k8IMweiYMkLrXgpFx0p2S1jti8voCCmKjJVvUKfpLVpQsi
f3kL5aGOO5261TT8d3pjo3sNbKWkc4jR+BS9j4hBgRM7cXnZWwQbtyfit8bEEHT1
zADmlsi7slr2PcWud+aJ3DBWo/NzS1dRVMTcIHVjhds09zLLa4hN0Qf782N6U8yZ
ARSw2SwAGlIYiWCnVtEm0SfqmlD0v6xClMRdzdRWCYt4t0TnVWDQekV5OgpEuJHE
FsyKIff4PisL1U3YhIbXeG39j7p1hiTKxb7gXveQdou8ruT8JeBRkjBMfutPTXL7
BqyBmWy0zs1/RhuKo5lTXkJraFYETAxLFQN5dfYmiBiCYI88HmKgV2UXMqVJDKDg
DY4gK/Q+y7s2JoOBA/Adqy5qkjxtLLakgRusxkDi27XMiCgePFu+zk5lnNqRzY4G
D7efXKabUnrjeqz4fivpdjOzRqIRg3S7pPr9WrCUY55BkiDHY2pgWT81DoveuT7Q
KdzxrSzY4ePoZkRJaTHg5Ga8IETVtkuv0Tios+hQ8NGUj0u6k0U1/8G37HD8hgYa
ZVeQtNM/PeE75FTuibFFmkOWbbvdjHgjv8OB3DCVytUn7mFvxIw+dMmu9pMKwkwh
to8IXPsxs7JI93XHqy7QSCwcg/0pob0ghCoEaA7H+SMI/Es5ecSADXapt7fXTcQv
JDmKdDANm4Qg3babmnxT3RsjbUnMv7hIpOXhkxJiypVSAqze80jsXxxWR9FzqmFL
Q5Moaf735iX+xSBE+bZeWmeCYLaJAGkO839b4VR6TFOoEEhFl76eyhxpbopkBsNQ
r1aaxdyGD7X6IQWegkF6jlrugEQGITeTkDA4Vmrkvd2aZGxgUrDPX0VIS6OKNJDU
4jSn7+R3jzvppyYTuTo99KcRUPGSwxtPImunCA/I4Zk8ymLx1OjjGdU4Igrrselz
RKxPOUEldRuQx7+VtFUFyQ==
`protect END_PROTECTED
