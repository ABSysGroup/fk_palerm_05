`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DTQJTR0EU8KccvQVqYWzE6B0EH38yGsEDo6XjYCLIbKdILAtI1ZD0wtl+cnfZOo8
E/r/U/zHGRp+iatSEBairwJktpfEUycF4o2SQyQ6uY8y4QlNabARxtFsVMhTtM9P
iR9A8VHXXekSnIzGtLJaM5WmmZmt6fKHMBDp7rmTNBdWyPoLWr9TETs2QtrmgiOy
4ORHeqGZcmZ56IJB4KuD9TPZe4djJOwmjYM7qiIs0Y3v3USMXW0DbrbxkJK1AyQO
hwH2eqtB1e20JBHOC92BOdkiM6cL3oFHouuNU4PUMnH8dS5re0l8DFUCifUO8NAb
qIofcE7pfstsBCnLoE++IR/A2frmn+c4MBZljTgTPLdk6SByNCDMggxDauEqwT2Z
jJjZGB3VxcLJ4r5zLl4a6hCHL60daXuZogaVpZR+Ii/iq/LDNOlVzb07FbFWzc0V
aqqucm+2Jaa/zmzUlCgU+4CjCLTtj/LlNKTUSDTYW5Fi24g+EZM1LaYz6hrd5n95
8JI26mATruVSDTMVy98abOXtVcjI4Xoirsw+QOFn1nVY09umiR5STreq7gZaY3hf
7TxrPRRN/ilnO0tLrgTj3IQLX+1MjJyHXgQoPzvIxD4Ive+x5QqKnPzI12fokENR
/ktUI5/9FtoNraDbTlSl5OaLnajLy0aRU6kOcH6cYSrgjlPvVjW9qdermv+y9lNy
xlwrP88r3oKkcOPommuyJuZ3MP7gklFej+YkBHbGT1QjCa4mHqYlgLN+ZCi8oSEH
DCszzffnueuFiD40sQjyfXDcDBeJN6F6I0iu3fNLEz675RD9ZFoCotWdmgxQsLX9
d/d9qrYbshpS8kBp+cVzYJYwViQmqx7x1uE/qyxVp5bBL+vJYR1do4FK3PfstQAf
MHSCI2Np6GfVlWljzXZgV+bFryktVLn+hW0KHaa5D0g9YVCtyruefi80R/KbxVHi
niyTirfGbhVtHBPlxC9KPV/zqU84eJymRDzZ5yho26e1ZSVRN8SUsVdJc7i8O4o6
nYEAlwuYmtseakfGuIbqGWOawqfBGzrbpiCQy2Ox7BPbC4N+xKcUEjSo9pudCLAL
vrv4AkD9EGMsfZpyt/OeH/o+Ad+mnLZDMUEiboIVCUZssIjZwe6HteRphxL+/xBw
jvn7yZJF0J3CXTN52SkV76rNr51Uc8FP3Iv0tJYjstSCXX58lOVuJzTrFZkHDpnT
SGwIYjnnEAZeSkWR6hTreA4NBCuG92EJSI198tLMqiCqWFSLL+w8kBUAgnT0VS/B
8yUgwzxGsqu1cfjyNqECrhBAU/TPrds0x1E3DINt7xFYVdsVwqPrvT4TEJRJ3DoS
xEB8QYw/sRH1rBbCHGZVhQJiSfomsVpwRmr2DYMTVWxBR/3B1ICOt3zM02VFJnpe
8NP+XCP2Qg9jOh4fB4IJj3dbkedJP88qkrXFzhHHivVS4CkgyjPpvPucXtSdGBB2
ljpeZvhvKbsBaFzJrYBVV3jvSc7vOcj1Xg+3oX7Yf7RVB/f/13xySBCgL4KyK6C9
KCH0JIH/ty0UrVZ2/P22jlt7G/BnyaJ6suEtLXqVVqKlskF6LtTVmU1qnD188Ios
JzSXF0NTwJVyvG6z008wpwOAKbr0OhrNhfn1hbDfEp4b4rZJUxIGEU/0f7T4gUoo
wm19OSynR9n1YLeDtb0+I50KJZTdQqyucf1fmR2ovbAirw0+uJJUaKxbjc/5/0dU
qapaunpC4FeJaT7fVqn7sQsCDQEVDU/RAwI7gCNWWFtAMSlyq/4zLwWMBjq+weUZ
0VLmD0XQ2Z1E+l0kfzgqI2L4OlGQOjPsu/XlsGn+rg71b5dtfwq4gPZD0gzy9TU+
smntKbNGy/lAwwMh0S/wkw2uPvk2Kg4e6QQn7upQlBL2/pS97mvOqbdm9py5AcO9
VjTR6jbAfkuhgd8RdXJAkbUClEPcdAjcDpGo5wO6FolrZeYiRWed5FmkLpVt2AEW
jTsKt73rqCSmvGwYPvpPfLaK/ljG0T5ZtBoWKdkm9dPu1SycWDqnPgAPEXN8vVXn
S2MUpd5pIFYXTZgRySpqZY8y+tJ+YISu0RGWXJ0BofLeayjrLXor8pYqbmiR5zZM
6EKVOjlJCC1korvD9ni+7MkG8o//P/Bx3TlKRnDzR7ZCyCMwHqdzA6ADSKiOMX5O
VsfSHJwbXXj0nvC60k2lptH1qrtuV24+frP/m42vvkU2aAyRoNDoFBlhV/6U0ikb
AlXieci2t4qGtMjis9E0NnD0aoCuWy5tP1o/Vc9GzcGFIaTGpwCVv0k2xig8t+pt
FgxEK+jYYSnJ5zrbB676feS7ESEFydsgxx2fgFqiewCMk5gtnJ7dttNWUvsroofn
4Kv9gOE1GEwA3Sufe4LLIyydiehvH6Tv9VSMavCs3sUZYNPTcZT6F4FaJ861eOHC
s4n3fJ+hzd389ZiOBzo9jekgxJ7zW2N3gs//f18IUa05JocRWFgwbeg6SdffCrUY
IFy9Ty6gEviBeHPj6+1ptRZM6Jn1XDjXLAMqtxckZA5DO7Dc9kll0zzSToBk7rGP
kr3hWeFnFpCdQFimdbSQ+OuMc9WAIgdaiFoTPFCkiLXuzcq6uRQTUwA7NAmAQ7wy
br2Xo1Io0dgaOgqlFiNGVj1U0dxtxicDfM9j0Z+v1rWFf+z4V98qPWrDs5QIOf5e
W2jfnO48F8OREZsZwpEXfHAkPgA+FXV1CF3kz9DrBFj+uHGwDgjBQUBPT6Ff5FhM
jVbIdhIsf08tG5BMxtmc6qW3O6VxZm1ifmJirpTTQx4iQr5iIPK1nZ3rKfESYbv9
8cPcTJhWKlp25O5XgDZaNasO4NHGVSbk3W8P13o6wcXH2Kf+iiWiFdZR6+0rdeOa
7AeE0AeOs06exVVvn36eWyX6/tgg/EnCYq5gMhTpQP3LkXSTqYzy+F0KpsBe7+ig
FPtoA8wfH4rZpe5CsLea+VLq0Dj8OzRSMH8YhKdFaFJDgqVFhIqoz5fIMBo2ufTw
l9wFHvGmNGQdokXsQM7iWfvWJtshp4fa4jHcAz6ODmPI/zo34Vn2ecr8XyHozYEN
Y1lDrw0qVQbucbg4h4V3q3l2SMcUpPnlRafHDNzagKHhP4F6b6QyVrfYq45fZgpM
q7QlLjAqW5aC8wuYr82UZGrtjqiW/LVxdQI+320CPoEIoX1xd+vkKRssAr3UwaJ7
5cRq/EBIaVKcJjf87brylYQin4bd1vY+1CD68DJNR7NpYCjnPLlmy3M0gz64COS9
ZwLFWxw2ZEJE47MtxgfjqcEm2ktIXKNym0c6hM4hI/XueFsfsAWZH38GOaEig0E/
Tp1fPmH3AR/21IY2xuc2yQToAKwySvFvmoyhWvfarLQmrIh/L65pi0zbj3jONRzr
cbzyZ/BIA2nSbr8m0piTWEDQjC4uCwVaEBIdKUjm+gOpmyvsMMaTCMrikaNFRHtE
bP6Cr+qMdV5SbhKZRDdBEsbsrxP3jR0l+IFN3cLEG36acsaeIl9pf3NCD+xM62mT
Zs0T8WMFQe5mx+slXrkCkGawa2FDY+6+1UXPW0FO9N6u2U6oosd5scmYWSV2mZr+
hqLcHySgSOXdoldVVVVoVgY/Aq9ItqrrCITteklOehKg+q65ALUnWukTL1vlgDBS
8KC8SvPEDyGvNlcAw7ZeabIVCt5rNg2ejcirE0HxV6dQ+xhGYkL24y4prZYH1MQz
nkO3Tq+0Mj5KYXSYRP1Rl9nbTHnYPhI6uxfvI1wxjZZ4D9R8c0U1t03h445MPlZo
tpMjRcbthLL2xL4xUVItpxKdSULFMrAHyRXob9m1HgGi8u1effekQVDMAiWukXGs
a/5NgNTx0oqDkk2/aBBcwc6q5lIzpUK8E0ZZw7B1G7H60qwwxJbiPA2IhegLXc70
xIsKSlJminnaZE1890IobZc2WuNvbKM9nvErAUx790AlsfetykihC5+A5/hnbAhI
tPtm6IRbz1ixTZqOjQmRmVDMEOZKh2/mAg4dPxeqvByC0gyLpWb9nA97SAGmAS6R
18pLwjg3QBIaqCbtm3UXqoA275RKKOX8tEZeIXjcVBRcZ9BSu/X/UjBB5HabqMcw
xlb53mv0x9D4zOlM0qRc/Qj6xlIZ+nG090OQBdSKk9M4UnlfKLedgo0Wuu0ZXXew
c63Scei2jXc6m6YQi8z9g0oKvAkb3FR24a0Yx5LTfKMXcNA/ZykBlL6jaT3UfNMX
KnAd8cziEhjNIQiRh/dUvT6H9zT4HbAYn7A9vGylkVRXFr9/mB60zzIqCiK76CGK
D9BFZzFvAwc9ps1Bq3QvHOs0fEErCnUeXYNMb8b/bSZrEFafT6fxdoYOCHDE9WjC
h9PEewJIh6W/dRagk0JlsS6kkleLUTicZzt/ehSrlOQ4YW0tAJe4trniCIHzPGCo
LMLECjOI4BwcA2xyWEnX20ZSHukPxSaykrv2DSdpPLzIDjDJCoHcQaF/GHatoNNU
Rv4SP78XxcYNr35pnk/1hmA1uCjooxB2wh4x1N/9u6qHYr36qYyMcrh2pQEaYJzn
WU8SIhgAXYJEdvh6KzIKZdi84V5bkYXq68uM0u9meRNQb3JvC9P18MFV5w5XgJYb
4HFkV8bFeP4aYBIwLJlAU2XrtyhbpeVBvOBelu20N1JfLjpWRc2Re4UuTFO7H5aY
nFt0ndxpmepanSaEvRfhpNL8txGgp/pHfNLk1QkR05DwLz0GOJKnYxIbP9tPdsWu
7iG+JNeipKGkPIzbNeenntJ5atUc0x8D5mmfXIEI0MQY1jTvPR4GxeOfGvJrkDPJ
3wFqfLTGI9OzSErTkPd7Wcin4Rbo9a5wWBusI9ZfKSL8Ga9ZOqi2mNshS3xRZawZ
93TwCiE8bAJHVD1zqFuHCpZhNXqpb0/cymW4catMo5U23yHElNc3Sp+xvBnWLMYO
V6YRPxHcLEQ/pGJl2MdTOtiWXnTiM3jOENOh+IKb3j6vsXKIwT820QSesDpIwiIW
RMMMozl2dLr0zO4MuDG1CmqhI+GygnJNwD6kXDfxKRKoLJXNKSQzF+FDEVTVR+rs
BbrYvTwQqOyVskkhkew5276zUVaLciSccchYP9hVwUwUUm07wdfgqIhQ8H3dUfyg
FRaD0oKzOt3M0Dwm12LoIGX0XmCrUuasj+opfeaAgJP4QLLJbgIZzdbPsZoIjNwF
eoT8VAPIUHTRHF2CnSehr/VYH3omzKOlPymMvD2WrFgt1mxUvFqaYYVNwzLRdfZ+
vML4qEaE7Cc1qvlIDtllIydiblLIdVnIJwwekzrJlfF6iuMR+g1mECBssS32vfRr
Zd8oGUj+ZaLhOL3v5jTrez2nj07SOGAqVtOtu6MjmyIH01Rl/GwW6HknCXAmbeqP
L7nowhwUtMj8pUEa9800+7hZfJnpPniWV74LCwefkqSQ2XLy0LGIfST7pfbjOiaT
cqmfA8PERMRLaLmJdc7tqzgkzEJLZJVE4movEL2e2oLDiG4gu7+4bQP2OdNBzyr6
Z2wp+6J1sxaCQyWrWirKL2km8OhHrohTtock16BBaZvlUKPSeXrzw/CNcJ5VficT
f6xRVH5LFje8WmQ6iP69lDN0D0PKLZcGvt16UOpGH9nAkZY3KKvxDbbX5GDDLgCR
JmGuoZxlxTbckZB+oto4oM021DiK2DI70rhuuX5JJnD8t/VTsccyTo0AYcDx8hcm
2lehESqKjaxwG/D7a9/MkQSCQR7UexIZTiT5NTuFm/PpNYb9Yrblvd+r0obg2uX8
3dAzdlENiWXYoyQUDhOCk7x8j+Cr9OSEDCk/2GGGa1M46GXcdlqpMG12govbq/OA
kln9SRt0W2oA51zZAKoinqV/xqXY91XpjWuI3uLtG+UDzMjPX3NOVOc0SW0jlDNC
bjFb0DtMfgJDQf8O16jxnC8DU7G0ZkIcRq1hpzstlEiKWUgWJr4df04R6/Tp1glL
HFkeOkucO7sq+zuInAbadyNMwFfhkPQKubMmfceI65PM/Mva6J2XZH5a0Mr580OW
sEq7sz2aIczGAHjoqqiiRQkC8Ey2iydCFNLWuQtvSv+/F8Amdn/+ELpvcWnPPL08
qEUjZt6fF8N51VUOvxVXEYLSjK68dwXbSC+IGwqbvGfmg19hEehvS7vZHc/bisQc
Erk2e7wsArjumI2TI0ltRs0oDyvbvD9WWZGTTK2OuuuTt/XhROwpks6jRdWnBqCw
ZhcZXXu4GSYQRFSDUiG1QwUIDB3YApQSe9Ss4D/wPkjiGlmol3JFhTUXY6IVG67s
JdvY8TWpVPuIKZgkc0YES29Kw7oGGxglaFMzqSwXO+pw28MPRtOSo844mO9YwmFm
gtLoEw1vG3YUTnuo5LSJ2ELHjR3fBYr/ZA8sRAnfTjNj5d82648f/r2mr/rSpAsZ
x5ZFvVnBTnFSxaihK+biwW/AwgRJjC1J/1f2RfS6+RW8QdjiAzmmVnBtFj2oQznM
PNr5bqQndKc+d+a3QKsReUzxkh7Yh/z1xl3Xtbd7Jwjf5Qy63t4P8iugIb/GQZ8D
DLZcYbjhQJ10YWu9KOsvNOucbksHn8Lgzly+mrPomM35EVYmnWpmc/DQ0NEEpkqN
vfmaTfhoOmSagJBLi9K0dYw/DFwhuTI47r+79j50z593pGhftF0r6ZqLZhqzN35n
hLni1kFcP7yu+PhfaHGdZtpDP2lkbyYTj4ksrVK41pha25YwagRbxL0PpW/XO6bT
u4838bC9DvqWaqUkJJopXKp9oEKJ7zQYloBPDtzuI2zD7N87TqO9PQTyke7iUs1P
js+HvbJ/mHkE9pTWsmRTch0wThYJsU/gyZApDmi3CbIbLjO2NCn+En+VLQ359H7i
nAYiSTljqH60gD4NSntPonm4iIpwLs40xftKhKAhm90Jt1ZoBalrd88eAOwDpz89
HE9l2+iRY6LPc04FZQBwPh1Tk/lTXDQpyOuhFcQpU6vNYbQiNGxM3W0om6Y/wXnZ
CevDsvGLVfYVmxdxSm8ocEYrW6mw9C3H0ewmYS0Po3XeMn3Fikodu0bE/VX0d1qs
D+7ngW944WRBs+hYiBVK59/QczSDn/f+o0JbkrwUQ/iR8mDc8U7tvZ22mea9AxAM
4i9xXeBZtXbMT/5q7wDmsGxc94w39aeqMGG2QCntU++neO7AeTuP3qyiUhMboRDG
p8HRucPHYA8oBrl35hlB4WKY7Trfa+caDxwWTb+jjLQ6LSb2exp8oEzCm8bMAgI+
OsNpY1w/UWKU+0j5EReF5CcFjjUuGbbHMp6iRULaGnWoPMcmn0LlYn0ZvgHn+HYr
ZPWuZNViCmSEqr1pvENCtTIRuQCjeIWH4zR4dpMU6X6K4ukYSMnbo9D6oruOuC/i
79VxDjTQT1RW/oufHmZ9hGCh1wECpBGh0DMDaGNe9HUaAUVLc/KbrAzBLAHAp0l6
cscqu51/8A6HCZ1bjJqsaSYeVYz8DWzJ2tqEu+aRn6VAqO5I6iJlteNW3zaUiHxp
nm867BgfMQ0xHyC0sMdqzApHFH79hnv+COvgpY3K6QNYOFHylKd+zUc6krLUqWIt
YHdodQmihzIaWtoSCIKZPkaTEGNpXeXBwiV60DBGAHX3CK5GObfvDoSpe23B4UQd
53RCzE/hMPsVya9A34ggTWV9mhqseYpociJ/cBdoFE3br3losEhVxw3TOfj+NHfE
8ZoW6zV1Xi/VYdq+DEx96XFCPWSkRPQiOWK3BX0ypzs1fXgVDK1CkgXZiHMWNNOh
5NK1ZfXs7rFJ5hBcUj3H2AJfITQlLAA3EsSbm7ZgiB5zIktFk4nuVbd0rchhXmGj
9BgbbvZW08EV6WRgHTirXkUa+7mKQRKv8soICF3pAF2HMpa0cpoamY3c238Z06zv
fQU8+BOIBKVLHj8tNSuS3wHbxSiuFWClrDDZ7xFXuSP9DkgL8RVDk/kIQzdVd1TY
StzyuWFJeN3yg9J20rpXcQOUwDJoH8dyjv3jr9eAhHnOxhqR0+XmUD6O5XlbTON/
PwGc9EfIJTxfjPSXWfmJaOE+MQBnc04FWBDixl9pWTXfCdzFSznQXOkeTWtvwYio
WOJWlZjkC5dwpVYeF/RE3CGNy/E7M+/iECUJWF4f/R2hljvv1dhP64IFtSSaQZcE
JmotKS0ltIJurMuIE1d+8xUVwnIVw0/+FF42Psw0LSFDfEBe6uUXAAj2ntVWO3V6
mNIB0bOoG7GhCAOaZuPis41VwyesCGUv9TloBVTLEbXECfz5LcdBHnLe1r9bk6YQ
jinQIXz8oYwTNk6d3Igb7EwL3NBxmjM0OyUKHT3xB7XE+kinZe9NF+y0iCpCSost
1JYPDCBpFTAIJ6JrzhEtIJL2QBDk944y91TrMhLWGkpwmS11RfPGNUXwURY4YNgZ
KcwbJWLDiNo4nbvLCFIc7KzdjXuLdpb5EY2E0qSPFkwCmW7amRRYZUTi0Gzntgq+
CUlSg7wT+mgvzK7fak4Kr3LUTx+ipbpuBvllLC4ICnBB9KMZZu6XVoOQf3aRmf0S
ErPtYkcuEhoPn/+ZF0WWFRlr+1MMBLmLMTl6l652ehSsh9X9BrWbnVrSWWd2TDNR
QjgziwJMsc3f9veQhGqFmLzK3EhX8V7yH9kMBPhAUE+RousyFAf4Xv7baQbWESDJ
YkyKbs+u1T4JqWK0aUq4nArdq6UZcCy3GWZcIA11btvb68Wmwq2GmZ+x5orao+4k
fgSUe7D8TVu8Xb25+Cj6wljD8/7+srmoIdO9z1T6A1E7P77hpM5OfaovALKkZUed
ugzeTmz2Wt7dG5xC3qCZYFav7AMkGeFYFGefZfy7URuZk26HAFZLs0+xO9Sc/CLH
Ql/xxKIwhXAC4RG3dYSP4YewYRSvqYtEB/9TzttiEeoC6X5gIySFEN8+93WoiQ19
2rlhJsLwijKImVu/aLMIDmuAehunWhLglYphHlA+bEoslQDPlGO0QBuY40EERAd7
soeOnahSR1jAbnJVKXxuWszdj4d7T2SzLG+IxrcXJFgPXpyH7QO9Wo29IiVBtqBb
sZw15jqe7qSppueXu+ypopKq6RXhzMWnaiy3LkoGCEOeH0SZArXpoa1HU4k5OLyj
pkUbZVD4NFbj4boBaZYPpz2yny/9KWFvbV4CQxqGHShLPbr3/67Z+Pw0wfOTW5cO
SUKQauWjc2s0n5INj+e3KH7p6VVODNMIw/KHCxEuC/q168hFIuiRyViPQzgQvq1R
DXT8cSv91CCGxl01DAgaFtC3xtfbyfkkWiATpMQJEzXh/o4BS7gXrFLfHiDFWQ2o
V28KvaX0qDnmpGE94ttV/YIDHdDyi10qKesaJS2hxW+qzIOaMkj+drp1MN/3VJaM
Hm7Dmy1MmdYQ/TKB3+1VqRnp1GiSCvKnaU/bvxTJN1DOAJyiQpTNsoO3KGHmO1s1
Hv2m7Qso0EV56TZpUHCQgiCeaHBl0gLmgMVfMw+tKaUJZ1J+0cQke6Bgedn7xCz+
odTD2AyX04KDQx/G5j86vm4DtseGY3gIDdFzy6X3aXgLrEDMbSvgxRSwwdVVggNK
VF0hqfqw3JeolMYp7fgDUDQsSGNWZ/klSp2grf2W7RvqqXf0rgvr85wgqXsHqmeT
YXiGY9hn+4VepBAVH8Iq14E6oODqWdFNjSpVgWkGCdoLsFF4JgVPdpxrWJ1WITPp
/holH1IdeorSx38/FoZsRKKA5SbH/G1Pqn/vSngyCIuKSGo4YNhpgAPBSjVIYQFl
JWMWgeMse6xnY2M4ieEVKHmOduwob/iFvk3MG0hSdqbzXs2qWXA/fPhhlNZdNUpM
lWqIfM22PAHkj7YFb7//9DIn7rB9j3YzthL9U7JvxiJARvPtc9om7n4qk1Pl4XrR
q9V92HZh8M7QegNCR3YPoAKZurKI92hFmeafaA2GgYh8geEIFRsCbb7dCLdzUQtE
G6FzYhtB6nWV4Xie3sJCnNeM81Xci+owmS/EefWKpp9cKVRsbFQ1p0MJvKU7JyeS
LAs+2wR4sI1B+R+2xPnNFaUD2PnHfYPN2yYohtgCm48FYd8iVoSj0K5looYyTwyM
H5q53mykOFinOJ25xyJLm6IdB9oKT2RTlrx0kPWFI2cKEZcBc7xS+TeawmWXdUnC
27rQ2IdN8nvgB5CX3iiHhB+e3ju1OAWI9zQJcbtIyJ5Ddot4+L38BRCnb+WpPNRD
4R21deU4E9o3lfgCzWk8Y8Ph2XAMxsSilkUhffDOpgkEFjBYjAdFH8vBA6Pz0/j4
DzHUwlv6yXWlk9Z/CJD/s3S2pCAdPN6Vo4yN/XE3UdHxrTD2K+4jwHneOjQb6bJ6
AQTvM1inQlmh/jaZsYGm1fSzCy3b0njaWZfccaRLQQHItfBa4mbTzWtu70MCGpsx
d1e2eubZn7j+UwTEgGGhWMO3xLbm1cM5TbNhRYY/tpNYB6ZaIBrst2AzoBip2cA9
ShQ04grB7/+VGfTS4usSTqlaI5Zq1NTMISD5LTAt5r3tIxOY4p/GoaDr/uXLXp4I
/9kbA5KCiuCYeesNqoifcTbcfakiRaCX2GQRlO2ho1SyIb1HMDK+5Blfliom2x07
yJBhKmBuN8yhqlWIJfEOhro8TdKUTP9czTmwoHGJWabe8P4Plii7uZ4WHngxMHp6
WokPdd5O/U59X27g3OPn/hHJSgFfclCn0ll8HtbeK54A+lUIXFWTjSjNfTsktkYa
sKa0+pMVhgCp8M1Fmp1yGMkdXx908aqPAAa86cxEqBu3RuvRiXUMwELreSCsFqU1
hXaACesxv7QVs7sbNPNdqE3M2SOL66qxbeoUHZrMs46CgRjKDP5pBxfOYUOc9MEL
e94HpB+YL/SSqrKl+1gevoVujxuRkzk6SCLd0HLoeEkVfj0KIJoND/UZ8yTnRSlc
89b1qv8AHRH/5JtKdugJAUMYKsPB04EDDuHlZJsM6ge6+st++DEsYrIIaiPDbzsH
6udFvO0HTd1392F8VGuAR0/jAPntJA6AusYkStjzrHOmUf1GVIpRVRwmC35ET6y3
Ddl4r2y+0p7XZBfcJjTfWjHCTwLjjrTX+I1yLnebSTdRorh0r2oQfWF9RmW4FkXm
aB8jQpvb7FB0o1y3gmDxGQJC/5RKkTh79i3nmxVoVLpbcvQG96Bhn7Hq/FVGdrhq
Q0B+9QDa3IqqFtfVRPZC2jS90lOTP/F25gmKFNYf7FavQTddZEvQKcymGUkyXI9Q
f3ZHfEi+dvXD0DRgMZolNXw9jwxXXliiY5GbUGN1BnGVEm6CZilx/yOD2tMdTQVH
T0vDvYlZ1mi4XoEM+z/A8LnfthmMTYgrSde5wMCCzabgR2/h8yUn+7npRGrlxFx7
lCNJdKxggm80eM4Rt8fiEieGVmbdrOgep2k2gBwDXRIjjxfjYspPpkybn5I5+6Gz
ltxydO5gVJiNhwzNjJfn/oXZ0MOw5WGrtuOpCPF2AckZ1G/5wgwzXKljlH5Z27Ge
66JdRs1FpJ4FNWZmkP4Q9CUkIziLtgWcbeVudQwNAs7qujYPtkf+dsedGLQxSrBQ
5sOdXrcYPdYEypuByNKgR3RvjEZS20NG4zJle0PpeO+Nf+AR+v6P2y988+WRzst4
Edd23ZOymnkcRydfy7+ugDM/9UTZkxWsTJIpsLJ4nAg98Rkh2FQ+XFdjake5ZqUt
Pix+Ov+axwVPxikA91f+ONTvi9EzRsgYzCC2rJMkhT3+0/a3SivdHWZ9nAqprQjC
I90ZinAkPiTk7mbiFuEMJCRv8V5VfW2mzut16mPzIerpx+RFI7igS5/pxaYcBozm
cpRf2b9JLdIPRujkvuJMhlwcmg14hP6jeNiR+pM74nlorYxP8aP3MiQaW+oFEPc+
nv7p/XIjSRf3ABLPKptPHyaSjKBoRxJcKUDoCE1/vFPYiqqO6gkTIW2bri97M2po
I11Yss1PDhpHjshIccNlEhzc1DAHl/FtVFCCbog08oYjVi4aljiH083SEdN+GEqY
5RiW4KkHZBJqjPE2lj81MEoOQ/ap+HcebkCBYaRN5a+b3bC0/flzpE6dpUoXA9MT
az6BQn4MKmcYTc97PJlwD7rGEWft5PGW6TX32F1T9MMG0qNBMY1Tjn+BwaWYDGXy
yekBhB3dnF/wWm1Y40/WidHqIcu6oZBXIJiGBf0/6vHyYS8fIgX1xGHwinJVaK8n
SNuqOyDw0sNkcpILbQ4LIOOrH6OLfveb1RRv7v6UZt+VRtmFJ30hfYfVu/MK4WLz
s3CaYBMkaheDo5CCzzS8lwmf5womWVZKVD5oMMQt51pp2K9RlwKoITSYXt1F5r1l
MQYvuN+BQLhz3fVIzPUBmNaH+eVajSb7yY7EyMSCnaK8CFbmMscvUqtmZUqP6Zqn
tBZmOwZVCHNgfi+oLTaadJ09uB4o23BVDcPmo/MgqoXTPz+1YqjOdtr1alH4QKIp
79rnZBTw3v7pLYD0gmh9wiziQiFyOaMfcSvpa+SFta8X2Elops1Dkgux64eveeos
jDOhya9sJoh0m8de7daG7S506dbRfRwhTP0dREErRsLicKOkM+W9S2w61cN7wghy
9R08EvBw0FpIj6a1Frr7mmjbgrRDzUDZaF0SMVXUjEBqpwJEQyBPMrLZeiIYMmR/
G6cmTEZRMUB3jGbjkYp8rIKGxiiv0J4DGZb9wYhPmY93WzEiKobRNHtIQgy0+c6h
5+1KM35nLXwPhMXxAVqdBJsG4+smZU0JjoAYiZmZ1kDRtxkdtA+Mo6/r+Ol5YCfj
H4jqJg/IMQx/K1LUKUlQkw1NQFw7vHEWdnJ1wurTzah/NNPPvmXQ20BEGr+X8wh3
yV5WBUkZ4n4d2AA37hCjqf0YTYK3UwPptXBmKUiGp7mtlWnsVfzH02rmbVvgHyeb
8fRa3SSlhbsnqCZMl/g0ZY+EQJI3b4ZtJHM4P06B+11Do9/i1XZOZAe4PEQzEwOs
58rluAPFIAWpeOju9OmlHVzUruF58PHOooCgeqZliCaZmQaPyo1tB+wbtVt36zsB
I+KqfEy3WHEeVdyfvIm4nrxW19/TI2SrNNbk7/duySGAaM6cHcpubf2iqsovyWmO
uyNQaoouOwJynQ6ifRCxW1gyZgGloG/DYiFyAHk3snZypSsskE36Hlx4A582jwRP
8Wi8J0MTyEoIK03zmZ31Nbh3QqJXI/BT8KIeJBKTgKTIekyRLqdysjcZB8k/eaO3
ABdtbK+Jk08XEiwvmQV8+8JL8XIBwHkXun7htRbuMPmODzCkStGqTF5uPwqvsEO2
/2yO97sNVQF5ynzkL6RhttmljUfPuqGzE+Ysj8BnVx1yOJjqUxoweWCpmlVTDCcX
20LigNLdijuUkqwoEDvREfxEedyAibVVlnEe/jnbIzv0AA5FRSnLxl9wqSeXwxtT
XKJmgMRS5thwHwUaqphDS6JlmzO5GkBv+EZ1C5VK/FW+dIjE6Csy6pHk6aPJAxTl
nA8pFCM56+KGIOlP8moYAWA6J+dociAY3wa7+2xwxv+Hd0gy0QHY93tPopDPFKXU
gN/fGrW0Dmhox2l2QWK7GwgLzqnfh7VgQ47BvhW/HnNaPkTsm25VposhjE/RO/iY
XIwUTLkL60HEGjp7q+pfW82bfhaZdWMcsbbY/lBrfXV8/p2LV6ZAntT6vjs4P6cg
s2A8Y5ofJ7QYzbI4K0k0NgLTOIGknffdYF78AoVC6LLpsts4kQ2euZJ6mp3hm/8t
r7u0t4/CTu2v66L2xSVFCc1O5T8XD9MUJqrGcBVzJR5jSCT8EjZW4odGSzafq47v
LwSaeSPFu6aBHf9wWmXZ5wbqZyyrNlLyz0MBB+juz7q8AKi6aHBMMkrSaf88BYjn
+U7zMniJyQcLyTczCnOmJejbpAWQyPGOlaih2mv0a2Z0s4HOtpb5461WPwuRP6E2
kqVtIkG1Lptua+xXZ1S9ygBAhoAcpm5cnVl7XYiPEgtnyibIC9r3EraegoXDptbF
WysOGJWnTPIVk36s1EMvCQuTNWrtcohslGRRf0Wkp0Hh3Db7rC+gCn2jgUhwiqE9
3LTgcTN6/CS4Z7JyzeqKA2k2HEUR9Tdjfai41tmNCcRLAglLgOtCSozLYS0kE3Kl
Nvx4CD+dZnpBcRmvLiZFvgg1G8VCMpoMPd96PoPMDuMhgSTpiYFrpyE3shBMsk2J
GGnmqleIEnxrtMandtOfQlXEZB5x8YbF3N0jcn1WX0hXUhQV9LQpEiHTJLd3Moxt
NQiI36rnfl0wf5MuMaRsHu+rjgSE8MrEFh72EOVVWsTtHdkW1YojclPnx98NQ7FU
KaXi8lR3Ldu1uBfcNM+jKPZBAaF3obb+It6RizFy/3GL2GJxpIAgN2nCMCTVpXAX
LPOxW2PqAGMqNZz85FKW5QRrdZ2UlzBp7BgO8CA4VL16iwtsej3FWhDBdCHxH3TE
le90LMVMyWptZ9Ka/OlCclcRP3LsEGHllS+P0AAAQfw83cCCyOvT9S7lHcAjwAOw
8AyCev3HKnQ8EoiTSJh6rNN4I78SO8Q7c/iSAsTzhSNtMHER8C7i33eJOMNEqNu1
oRDt4bnzY6UgzIyN8NVrXFDEdhVOCl9s4+oLfkOr2CWAYOCkJukHqTuu+2CvAayJ
FFXgfgk/nwSpw0IAQoCC/KD/MVznI+8A6IhgG3xh1F4YvhkqdEt0KCYpKUTQSS5j
REY6q5QDwbUgPMBCuTRJ922r/9+NjJP+xYEVgw46g5OCp6sF+IhNZQF1X0hUaxMI
y6Klk/MVhvq4Bd/UP37HlZiF4r/Xj6CpGgxwACh/mtQzbedLpZkKuazvgomJddTP
irEBViFVAx+IQdlgeIfbo/ZznWNuS4FvTdmeUMl1rL6uKFGyUj64zOirTLZE91q0
uW4K8QeZDRe9/xesJqcFRC4gJFneCem/rYzHFyp0CWZOypTKB00DKIH5W1AVF5vY
4mcGpUAE7fm4yzOkCndmD/W7snfCE07L/SfuC3qcRGqsk0pDOzCi5mguvOaECvmH
+9XexHEOvLrhor4BjSHRp+If03kIZCepIefPTjPW+4FAd0U19vEh1lJVy3HSlRiA
3aPD9y9+nxVLbkAPq/gBMojOjniRdWQhMrIUVw3PQGAXEbR/goDHkbdIiH7wt8KH
z1t9cIL1Y08kmdy/XBBueLbJlLVSjpxWXEYYgIM0FM+3TVN6+MEQbHNgfp4Ao8/M
nGiq7Et6uEGheuGer3uBWxMaSOA1wxl2A2LgSXPsNf8/JjZw2EbNsRL5l07/8R8C
sHYmD569VN9T6zEbR7iWM4okKZaIp4tpLhOdNVVp+3aT49DUOoV/s2EjeKF/pqxK
qKHZQ2ZgtJxLx7tdVoFZFFfv7rs6FSKlTXsKWUoeRDhReucJRY9gKg38aQmMUj+o
b5QGhD2V45apreUx0+8pCCZK39710DNTmp1SPE/PKD9b/VGYJslWPznG6bpHYaPz
13tmbcsEwv7EEYQr3Bj8YXy+a2kQvp5M1FlPLdUU4QZSDNyPFEI5W6KE6fvIJbjB
CXD/7+ZwjtrpeFe1uZMZLYoVsRvvD23S4yvztIC6LDZR7iyVHjY2r70dsZ2wiLsR
xFfaRYbrzaV4WxR49jEKwfMA9XEkPZNsTA21yefqpcFQuCQoDCexPlYq72o7SQQe
jBsugFQ5M2JzwV5OpO2r43gQbxxBPeczseO6/pfRdcUUbCAaSaui1uRbYdhK7Uj9
mmJNWB73HwKpMEWjjhz+1ygtXBZ+Jxt7BKCff2sellmxcEEvKP2OUjC3DtdIhWbT
QgfI/Ahe4CHWfCA3XKyRQ0TEQubc4myPqX0uHE8dnMFZfPEJDUutxRgFuuEkcVd7
L51NMdSWFE/3sFDXd0KnZZP+PJX5iTKpRpxuHESh0UW+GirZ9xH1UVEPhArIFjse
+PmbsjWtoQwpJncKzyEl2ID6kitmmlh7b8aYZlBx3bwge1824/O1qUM7/vC4NNwB
roDgT8PBl/cd5F6O2Hj4MxhrlZCcKlkyrQMwTyypXVHKquRdwTGTvy/ZxojUGvsr
rMOhxIbeccSVxoyV6gru3owLLhNadYSLLjDeA+8O2wzhhV/3MU5g3i9ya3KXTgQU
gX1Rgar6dVP6ChNFk6ypg1k8wRxf8dhEZUiPb6toMxfscUyOG//P7FVShkO39gGN
14VlhvBdxBeZRze5+nqMCJGMdiVFrftYpUbsFicKybbIu/D7ncRHBXWiLKfmUTFy
+hrw3YIonHAG85AUcA9paVhXUCNziX+f6fhnpnDVPvXc8d6mgvzj9mpIv/IWAp+6
AtusA7DeOVgdNfi3UIw7/qhAUSOLjLRPrBk0r7MZpKgvcVPx8xZG6zk7Pr2tnlYf
vSWZF9Rj3GDHIikmYBWq29N3BxIboBeF3L8aMQiqkkn4tW6l58ZjO85UxR0Mu+SK
rTD9PNyJEXeS0u8w5M3hvqcJ3gcVapeautC/15gCve0uh9sBfLxjEzL0YUIY5asf
nQunKjabo6W4ntXC4trSMGbmOHkU7xy+dHWJHFq3KyR0UxBfHxAYY/coNLPMSfLD
mRThs8w8fSRecs1KjZcReKqfyGos9yl3H+bcvw9d0ecOfs1OGTQp71i1tOdV5YNc
hW9yVd5612KCSujyX1DfBlRtwgXP+lAHIvIYMrnVz2aDpIPwsogRmAZtIizFyuYw
xcTD3j5w+G/h2DktFbhVaBP14IPPXyqXYtlM3+6KoPWenZcQO5x7tLcuYb8j7MWX
s90pt5J8hqaI12/MBakCwnF+pjVgDhJL0ufJubCVlr9sWlbSpfX1T64380sIPVCw
aYMVQt3PqG7hiVRpy2ueOmlPjqEBV4t6R53CzGT8pgy43/1yElYuDkNQKWZlAS+7
nms8qX7K/hpHmwQDZjY6clg/pAzEokDjjVynKGcuPOmVgkT0+3lKeviRBkkaT89R
VlckL36kFBWY+F9Eq3LpXJwTxdIB12tjjUa0iBUzvOyINACapthXLw2SHAldltIW
evpAlJVRd68aUb1d6Spdhf24siRsuV4ZhrGg+8VJb3kyq7PVoKaYn0jd/UMGseds
fxTRg/yJ6qmKynfSnYVeytpO8IliYY0yYQComZUq4tIGiovNODxsJY2sk3bsF49N
iCOOi3YNaHq5PftX1rfKwClggixeDDgtHKZi1dT8ay3K4TDoqaKpV+sXe8tgHrTQ
qR6b9RC6QlHATWnh3cw0r6y+/DlSUFfKLANP0faSPIcRpEt4gU+rHubeIkP2Ab7u
X/ODDDxx0IADiuxxAOpH+O7ssii83MUAdUw4nZSWv+YaxTv+pnfZ2KYlc7jnWVsM
PLU7nvXsadIo/HJQsU1edTg/VXkzDZFvtzILWkUOCNislao0J3VHNBHmvIJ30gZ2
efN7rojXG+V83PA0vz7z6OIBQJNcWFTwexVtFLk761iRlWuNJlO8neTCJY9+oz5Z
ELkmGXssahROiOoSolYcl8Sqma6v7ltKKuHavSTMdE97WogzCcx8mERCXF/1q0Xl
XJNAO5f4aYj0oc5S+4kK7YrydgmS3/LW+HzFcxWQvXtb+/PYCiQulOCYO1pZx+iM
4+Ps/6OyZyiR3tD0ihOcxhg5vYHB1FmTBSb2vJjLW67g5Qr9uXOLTSQIMcRoYMnO
jcIaTNxiu3gwa40P1YMH0PWLH/hbdN/G+wbHzNQMzQXaVRM86eiN29HSyc2dvFan
VTfg16wk4hxUHmHr6WGK/rVAiWNBfJzEyTxRZy/oShus21Q30xoWN2cbNLWS5n/4
hzRd6en06ZMGqm2Vu99oXlWGjG54JRgQLvd/bK8ubflnzKNbSCsRxK52uWTCcxnm
nCn4i9Sddiek8GrUMGWyUrfyI8lNyqYQoSX28mEkvvT8ncKInraO8CXfVvCnBnMf
SktrhAcifCkYpTX/qowRV/yqw2EBd37AfA0lUYvd/L7MAE7U51UmodiPdyyV9zsO
6CUzHhhTOIiOMAQXVqqut3xEJoZw5mUEBUx/fRO6VNygMMBA9ID9rzmMNE82kq3d
XREWVvXOP58zZWpnuivGx0S+DRzktUR9IwhL1rmUwmPFxnj06mcAwMTzIqF1zSMJ
fCemfTD/uljQokhV2pvonk7IKityUznK6nTsuVcEn/WQzNDiuoMdGyMdk9OptRs8
e0lAp0a+BG+pUrN97sro4QqogOs7X0iHiACmid3zA3m6rKlfI3KgXdNJ77XwnvMJ
6rS9qAM+xta/hkvTE25hIZNj+58PQhS6nACUMN+cgaBI2wVJ4kdflR6IFL5AHy7C
asSn2J6jPqitA+QWODImzdzGw53uxyNtb19AcxTXkbGJlw/M02zJb/OLjIuT70Ox
W0p76ojzjCAHqf0uZ5O20w9Xnyx6qW27/B7bU7XCRqikkWFtNBQTlyhBKAHR3R29
c7jCrA0G301jAwk8yxZoOKR1T02WykX0CbzqYc8EDrToPlYBUVZcCtjgwLStsyLt
6/j64DOSHFTM/4ya6xrSyPHT8nYtP5S/iXiFyJON5n02bS1BNAUIKimG4cetETAZ
gcTW1EK1Him0WMBGlfHmt6hOk2eJYUcwrG4JdVrPI1bQ9EX95G/H8Sx0NJN0I1Jk
LNTSpMXz86jsBbhMWRb0z+fW0PxJryYCc/FOPq+/0phScr5awG1CE1dxZPx1SJc7
GcVgxAg2vo6TSE/pCAItP5qZ0fQVV4yFmefZTDPEQCRm4lcxF6nlcA5/yIxf6/lX
UZZXxHd7aYrab3xBFz4wMjDH/SSOmb5WkcCeTxtOXKSAxcAVVbvgO8Knsq1/fGZI
j3PYhVZCuyTldHs7+yPfQA/xwM2e2VeYPdLIt50mbDNd2JJbm1IKrve5k9Dcfr3F
t47hlOrKlZ5xf04LymFVEiUXZQnM9jxQH29qh8zyfTL7QTWl8wSLdCpErCZqneAt
ZTeVAcvEn9bGloB1jRCc57kFqjT2oo01Vu6dLsIBOoJ1KXIcXuz709mLTbn/P2vp
aICCwfpJujtXsh5v42ls2CVv7lmfo9i9lhlluVHFXUTLwCFarqkhsO/x6PvPAzcp
B+VSdjnCBmFT3Hxsn8sOGMhaBp5maQqq74yF06BY5vl7GrEPv0assPYkYSu4UjpO
QXiax2NFr249wAh0cnYEZf//yDrtWlMlHMTXchM/SBo/k8XRAzsddgODwKGFredU
9C4BWRdJ8dw4EhCk8qrly75KoSbobs2lQmK8p0g6Wmxnj2germvG9M2pFlt7lMKP
Mr8YX4O2md86QLBNOllIaBrFTm0iXopLgCbfUKS1NSLMcZFpIx3/K/+OvgLDAxla
Vl0zQKpzaNCHP2za6nJNjdsT5JzayLrnBgjZ2SeY3QV5UZAzPXMb0Nn7MMtJHwTG
BU+Xan20OgmY3gMihuYuc7xkHpoJCxp7FxI3l4pJ3WhN72OqklQAK2iFhgLmSOU/
16rPOaT0rlDLwpc6Lzws5jR6Vt0SOgVK1f/lyaNiY01CJN4z3R/zh3L1IgCDcY27
RaDOGw1VNrljuvC2zLOWvYTtKL8Z6NVqg4AnRCcp8h7ieXXk06nC6DS7BxaprFDB
4GF3EvEmFkhZTLOkSA3GwXV7TlD4WsI6wNNZgZgM/E9f7kbNAnuHckk+ypIRRW8M
Fm1sc0/14vIZ70YDHVE0vg8OTKUQevbcLatMWcbjkbCFId5nnpJqp+geWi3qoZLl
7fBmxFWvZsLoDiqQ5+nYLvB4fTfBDbLxBFBqgmCEX721B3jfKMMo1qU/EUQ83juC
uvhfDqJ1M7q5mS9jeHXE7sODG7gLoxzYT5G60cQQ62QmR0gVydFPLRdrymZzu2QB
iRPMdIg3Kij7fwwidOpxPlDcumKnU8EiKGO/MK5LOO71Rt4JE/EKZ6RQA4NCiDXm
4xaN1c1WNG/P7dJJlYmbVGErMeFodKpnFR7gkT2xFZnBBkpzBRIx1e7NdBZTzyow
SZ6Oj/oaY/NE3Vr5dwOe6u340FrHE6MZaP76tt5n1eBkD3d2RcBPMemr2qqUfMaq
+78eBarPmDktNZg7YqA/6u21WVJCyUNUt7xfGGjhu+/Q+/akt5yf3RkRm+RXG1ey
V6TbbQBZLPTY2oLpHkxrvxfb/GOULQ5Ku2DmZT4z6u2PVB5nObPzJfkSpNi9FsYF
T5bZDqCz3+1BWRQ5XQtepaP7W4U9TK56/KBdCCD/NoIrWJTwwcGSFSKtyfcQF7Lg
awtmgiPKLfnhJAVb88GWdbPb1rAt91w7kov1pcZfG9qIC1cGeAVYnnL7fviS1zWm
NxkaCe3KrArWVcByOCypbVeYcsSeb0VzYXTTEcvNh1FRI4pOOsG0LycjkykYCq/L
bIh8HZ6a0IfOgjXyMcZr1gDWtGd6SeU2UcwFmM1x3e7FVOcyhrbXXU6gNhnu4qEu
akimRwwFFSReFbL07dqFHEfEqra+I2DD4Vbop4II+jftv/XBBR5S13OWWSYfbeT2
pFjt7RbFSlyVNZrKyE2XnYDQCrxuMBQ+DeW+Ko1JMB8SW/U0MQ5nCnxx3oVzKeZK
5Eyk2kHim8fMWlrPxFSN9bdnSNyNUVbqI7yTxFWEigfvdRKRZhBgRaxDjPQQg/R8
+pcw/dswC/qENlygLWt52MpeIVk1ncc9eH+kBNG6eFxGu0K4/SExJ4uNti3St1VQ
6budoMevmaRWL54kRx/yId+hCWS4kbP010URReyf1rvR3RID3K0hJrXzXOCZt3LW
3ehXBfjkN981CbBPDAn3kaSCyRz1KYNHDzoIFE7DOWTrNnH2CJPQTMuClwr5BaVu
832aNpmxZ6TSMKCjFVlDli19ENfDRewadhvATRQ14WkCAD3tuezdtCb+/bz0joeL
PN/8UFUciO3jUVVg/Z6IBk/JwvpcOvUqBmzhhL+xrkCtalnu7ybfuYt9J1XS7vAK
aoudbG1wSs7pdamFibMA2vOJN+m8i12A+Wb9AWtIuqwXNTm7uBVSureiTntWfgFr
xG3l0H2tgQJ/w+XeUuLAGUWgya8LWR052C37wZxsCLyWdvv4HVH90Yt1v0/xp0SH
bOVaxhEgUgCKejOLpFFCIrY4g4vkkC/6Flqf5UrWxiwI7RMtORZjv+GjZif9ZkV8
7irwkG0tTBSmw9kbQO65Ar/WllSAVDkIQQv1qp6AiG9tho1NZyrTQDa4XZzF4w9a
6iiF6U3Zo9Ao+wStjWToczYJOQ3UmdwYa9CorqQPrDeZQgu13CokSDqsw+8dRQFA
0isgSWVEaslVHW4lrh/aTxhCl37gcoWIz6O8MexgRA6aLdXJGJ16xAXe5Fh04+yZ
FCKoj0CsSRfAAZN3eEw00ZjK9C0y9a7AhMOJW1YUXUFaqC44TAtRDuz2DcKAUadt
tIHqQyQoqP1nKlIPYwI1nZ6n8NSiF+3FEob1mGKNDHbNKKKIWAzxS82RNrXT9Zv6
huFwid2xlCohoQquQ723hFFeIOb+WUzc8DG+cNv/yHLE16tDSZP7rL2M0j+VFMlI
CH/62h3QzUt7lgEvKDt4BhbL3l5iO3fG36ts7xPd/Ks7roZRfDq7HIC1mq2QtFb5
kdJ312pv8HVG+lrYRSNW6Aw2pDCvmAs4znMIqfShz8+A9KCL4gPzv5gd4o0kL73J
vOuXle+0JdMs3usHBSAgjTLjwXK0cWlmagb+U2GJSABcyNpcMkK4KMLspYW3Sgt9
tFooU8F74+t8gSJUhprpYEfmo2bGQflUT0EtZ9yTVW8xwiB6odWpua9BcMM1WJgo
GnA2icgABA7dG4W5480f9V9PfE3hG//pmmSvPre+HwS+kWifK1yZtYw5QwzeKKeI
m8TXVrZIzweOdpQou+Y9/W3AdIPzORzMLdXYcA334lLRpiRM27/yrCyy4I6CYUGa
IYcF3Dzz4CvKJpYtJA3141d42h9BDL6IIo/4KMZtIff6o5tbM3vEAaVfZ+jYQcjv
14Szj4gL7EnApYNdjmDZP2m/wwv9ESwpolDyGyeppUBTIxdPtidvsSdP/grgPHyH
L+WawQnkbBWEcN1sHK7XdW5/poHWmk27R3FGIb4S/ynoAmSUeit0kQ1mLnXk3iZt
6AXi+KlInFnYvRkgEE0ny/I/Ru/QdvKMmAAoZ7uAXUQseLIVvmQVQBY45SQpNO9r
kmPEJB5veQaOD7Mo6l8XFLELuytIlQ4VYyzdY1ML6UAoMyUICKwndd67R22GHw3q
TYj5phXTliZPGAA9YQoxlaZrlMprk+TkPO8aFJNx6li3pxOjpI2+t4F9gpPQHOra
QTEHxtbhACGQPZfycMcgIz0Z76pue4UobRkgZt5rB5u79FQuX7Pq6fitng3CH4lp
d4MI466wXvLqkuzECJqfhmRlB7ePKmWIvGmAR2sLgykTcRdhO7V+PHYQOYwlg/r5
I/9tqtz+oNYs6AjSH4yAU86aUyAM8eqvLMztXIAUnBncaCgfT3jdjBB+n8/f1nAd
92o4hbRgHUmN7sWJWX03E5aLCu7g9Bw1idJ7Sn8WUpZQxOEQ+UDz3eyLiZYalLN3
LjUYzBa5o+mLDdHSX54praeqK43xTNlsW0XcMupbCjVeUQq6dEuPgzFqr7waCuan
dCLZu/ISXR8uUJ8RQwZMSfstqXNhKAix99CLQWJTBNDYH4hUP48/vwiXGFU/LDyi
9S1YDAYWcU2jnLJuYVcbOSyMwJ7JAEf3IpyrSwubPyQ+PNmLgCEQSq1yobttNPyW
VJsS+SuxAbrv5IsYtJen+RInHt+hSBXC/E56dHxZW2JtlwC5GI/Ht0iipuUWEhZT
QMQJgzfhnpMq4dmL1SxwtGZpNvUDhwFnc/cfHNMO/82UGsi+uEz/9m7yOTRIqa9G
wVtANkdqhxH41sxVswn01+aXjVjj5P4vzTP5EG/T0J+kyQrBNP68U4tIve8yybAt
skG33y75MvlzCtStdQFrUL/j3C/pkoP8AVDRHnVFTANfqWh2EuYBVD7mT3TVgZL0
P2z6GkhyxpRR97xP4JAehYojY8wvEUUb6tpMmJS0OCLpYC1MBr3C2Cgh00DLG1cQ
iJ+6RnqMm1bBnK/OROvx+8Cs1IR5LTfWKDbGAe7RvPcUNzd1rXBialtYpwrWiVkh
BSJhkVt/hgkPP9Se2FBrtVLRqTUlhwON3U53qCXUcvTlRBrS3rdydhEKkiWYAgVC
+imoSjNu4oid8WhKNBWe4YJWBgs/FChnrohbgfpEu3q9AGgYcQzqtEljrQtkSCTV
tDzMpgZfS8TTX376kQHeRyO15U1OJHY8UQMGKOVYQRvczBwj1QcDE4MoTI92rbUI
+clVXFRXceREFbynoOtumnz6aNlFgFmJfoThCVSG4tAdtQLjHtkgtE0j5O3hzYXW
CaOgvPH4ueAz39dFMVwpoNxj+CO4bWhq/q2TYmsBPrM75kllxt8revHee+XVQ5H1
EtqKVo2i2NfJ0rFfxhCikW4WSQojRy3+9qEcEWcoeUC6XGavJVVaLgJ4vObaCP97
ZoAMQ4kqacwLQTMnj+SAk2lxksIr6yHBPtbV7Gky7Xljv+fGp6Q8rd+pYcok0so8
JDh4fX/HN1T6TQXKcXZahGOiZXdMN1pf4hBpXWZhOtEG/9QRdj0PfuTgWRgm6JN1
u0qnM3BWj2D4T7t89JcJu8CjhsF2Fdr9ZJfGNa+0OjnaAnzi/vRo1Vksoi+CfI9i
xX2H4hM8OwUcJVBezARzqqLu4Lyu+fwaJrfwkncdMWhJ3vJgTS6cNM7SytT+GkxC
8qiKeClGbRX47fys1xuqQLQ6IF32oyxJYGnzixBfhBUqRjXFXjLpC09O1SlhngFo
3xUuBR95SrSJ3DAFIHLUtXfn+I710BFaaNuqND6zJeSRmDvW/klTUJ2rik5XpNPH
z0HP8AYK6ocP29L7WX0UYE7O+BRQ+hiET8fxyKfospLYQqX2P3pCx2epXAlMkeg3
6jqki7hNQE3CQwz3fqrr2bnWr0AdN0mYf+uNKypPmS/eNjf+QGJZGZyIg8Fn+fYM
LLBGdfvaVJYp/Vj4Y2686e4l6O3xUZHVBKeFu02uSij45TpKUqcTzCuzhIyPXGe4
u7XXNu82nh9chdrX8LmHazAPIDx4hi/cT/6uY1bYPzUBw8YU/VclGi75PJEf59qD
wTcGih5LcsHHYTctItRCwu40mJ1g1qkovJLtGLsgiBuD9y/YU7UeAo7wR2rkJOIE
1W+7gLsW5yXt1eqNDzTtgopDih0m1d4MXSX/9YYt3j3HD/OWoFkUJ3k1J0lgmhMO
GcL3ODFPcp/N9yoaeg8uZxtjp4r1FSA1/9jlB/vZvqiWLRRYvxmHISGf/pt5cNCV
tP+KWbqm5zXFdpLG1OMvE7SUZkf7NkSW7lJFX507Eufyu2bOAZt/zJ/Nbbv9M8s4
T+36vEaCDNflDBS1mg43G058uZ6hYPmpAvSb430l57BvPSc62RKk60F4ZJ5Io4Tp
db34B0GP5wBPfmOg+71shn1W9qiRjC0UoPc+k0bTwlov9ofsC/1776K8TVFTrmAF
r0BtBeRbeKNQj70ioPSgCxznM44j8rWUqqkSlo15zPudErhN7u+xUG1MIZ0XrAYH
t0jxbeSmlwYHrm00TE7zIX1tDrW7oLynD006xbKxE8iM+RXiI0ljBkLMWNl2aTv0
ZSGlkttvs5FLf8DqyQFAHl4BVbRkoNbXEelCdSuRS16BVYv3aA/WLmUgjp1rNsA2
jO+VM27MMMa6SSh0kyH5a5yOcS9PaHpHQfhMZDpEtCHBomROGvoLokN+DaAFwoUC
jmq0GVyVCWdUuW++yqbV2kzUW57ehJM/Ww5u9/Ud+i0rcHN+7cVDqFy4f4ghUZ47
6aX6mBVUcShRW3KwMqhKlx6abOdjBl19uBOj9bEaLNHGMJb0rE4BLbt0n0pxL/0f
9KPx2Un02XZ8uwDDSpPfj4zlIPRu1Eldj94qEGATfJ9TIx26Y3c61xiZC+paNM9s
9KzLAMEEVPRBDfnHqNCqP+IPVHpb0vtZU6MxrSwYqy68PPDOL96IHDrOVPXoDdiw
i6olfiEh4JPmB3qmv0dsxvrLLfWMnfhUH9ZiABPFg6xi3eeFIyEtQsH28TP/JSeE
dgNlB5XNGDnz01414mgWE50hbVCztMsxylsgE0okcIZqZfI7CqI4SVoNSetnf01Q
8Br3CkekHJ1+18a1bPeO7msZoEw/0mGx0IuX/A6BbaE6rh36d5gSZBJX3LsmGoHR
Qggm51+nO/EMykvxmSNrV9ZZabtjKvZm4PuSNC1JbPdfQv2mzW+Kmbl6vENlkQX7
lbC0JjpfWvOpTVJO8bJrto6iET7rtslNr8jjNhfyTyA+lhuN7U4SKCWrGQQADFT7
aN1ts6DXw4wp8+LKv9kiA/FraXVCORVYRNqJkJfw/1YQ8ps1vCCmCWcs8KOfm0YM
LZexJSBiycH98ahoV3Xcb4LnNZcpadC2PoNjqI3G2bv5M9eaGjFe1HMq8nqbI91b
xALGAqfrSuHqMWgvsRAONNacfUrJ9wjUadBgaCJ4nh/tuiJMVbVzITIIkhAxPWoK
WBleCqCEpq4To4OW1zdq7fXIkNsNcBv1Kh1gY53qLBOXTNsZOwzzQfda1AL0shcP
H4oFRvOVfnEawWMLu7byHTMKNg+Forze7mK+s3s4xJ/mx2LthwjRXIlelx1FAKKg
uCVzvW2jJS2Lw3NeyD+jNcp0AxT+BS3sM1qlWLYdf7W2YOPhHOpacfZ9Sexwbl3V
nb6oATTWI891Xnv4/y2lZEkIMusikoJP6m2YiOyv3BBUZhL43iAL9fw+Z7OMPeFL
Tk5IjRzhvlF3iPUFBLrDDoqZZABXxnOwFa8qeb4M+6ci0OzIHmqdLjJWOLzXXAiA
OxFBvopivLxSPe9CTWalxZY3uiMwtEv9G91yPtMk3mT29eAaEKAPJbJ8DGQqoyQa
evxex3ENJVr+0zYW3cdYTNIwRWrAxvvlaunYtrtAtLItm1Ovysmc0x6u+aSEAm+a
1D+n10ANe6Gub0eYpBduO3dJ4shXvHxkxDcahobK0luSJSYtaTsF6GEOzcmvQH5U
6xdoPP/t4uqA+e017uydreSDuSPR5NcpdB4R9K+RaFe/Y201FNdr5hruzESu7jeM
yu26rkcyJKCVqPImkbjE2P5ZXD6pwMhIau7f6qtGMY/PJJdio5CAo8A1+r8wTE8k
Wny6Fv0348hOsBSsfaa/iYX3NChw3IIQcTEbvycnPzgwy2UUEzkG3UM0mchGvSrN
mGfpa/ATIYa2oxQO7BaCSxEjtyb7xZ/wBcZWA0d9BYV9kkCnH2wNDHbBf21XdZwx
eCAlBOW85iLVf+mmKvj/tlVGgq3xY60SEn15ObWE3Dp2vwvWNFVHLk7x+lKHfCAj
AD/bwhY0skhRTiNYe0OcuUHvseFeaxVqFepSo4Bb4hrHvqw3Rf/SkSD6QNeBtF23
d76XdH9TDauBwVtLFsp2qzymZAUiOsfYCvrgAxDT7d+2mzVhoz4yRPjMk3/7+iSz
AFtlXd5zoUhZLe+5ZTPwdQPi/oJX14cM1cgS+IdWzssUOa8M/FlfgdYslNRnF0HR
ah5dnJ9BsmC9hL/RfjP/RTeYzNxvh7h781v1R8zPvCbEFcwnaZ7glLX6AxbrDSA2
H/C0TTbCeBA3Tf2hjqnzgv/gx5dsyPRuk/uTFof+xaYDwaMv6WYeOKxBT9F5QznN
JIjlmRRA5G59pxdTnKTg01XZNaz9t8mNK/S0k9Xu7pSWJsjuohj7nO6lWeTPMGbN
xmKLg+FnfyMWeVgJNSV633kxgse8Bq1HzMTMqMxRLzNTyjtDvyx63NLwXv8jM3eP
3CYI0gZYR8cS1iI8Wh4SzvOKttB6bfY8cp/zWxpAfXabVpWcHWN/YG+Wwk5ifynk
xgcyYjv3KQMd9oWXP/F+ft4YvJ27aRPUO+KSzgSfPXqR547WgXRxwE8qD4xd2Jnr
9j3SNS2Yh+a1ryH78xJyYXa85rO1W2kWbt0VFz+6iVOs9km9tnEclIE+GzSqByA/
XYE4W8dfqEHlGO+e6o2dNu4zk+4sk+SxbLN6sePPiOZQFGxbgMZgRM4VqsQKSpGu
+U8/+Z/bib5qPBPRnyZDR9yT54nJnrr4tUCiKsWz3CnGXgSMDqy6pILFjb9R9O8o
tvfTJeaxaQsg1Vy7wZQ1zAjaIC9vnaEWNxWrWY50MZ6n4Z7baxlP6Drr1ik4BAaJ
E04qLf/m4c9s5Ns/KCR/TuZgtRpEkGgErR4gws6zaKnGZ4v21OGFY6flpjstwRPj
pcxRYXMMW3cDwQiBNp0hD1QHsoB26qoVoxbtxDjljXHb0RvEhCz4/QqjlS8C1FRl
ZsUUOPa7uHc9eaAjI9yKry/havBsBo39TevS73FQ+0C/vk3wWvrA15n+b0J7KdvM
LISuhwVtmLr+BkrOea6PNu8jD+awVIOn5qCegsyKBdm0YHi+aLauEPCX3SDuLRxU
TCyF4eJZtUz38kj6CFpNRK3hhbMGtKfJM20gkF9kK6flkd2ty24pry9R/w/D1sGI
n4pjxc9zwx3Tm0gBwdrnePdyZqnoRVCaaIPTFbOvHoerXsPKfIM0Yv5ygGvpwB16
ReWTwN4NqLelYj3E+riacv3LCzaVgu4mXMkfHEazCIIaGZlMwWWoRzTudiwu8CIh
rCY+oLu1C+x9MO46vSIOGOn4OmN8tAwrgd0IHn5a17wUADSzXuDD+vrAEa3wtzO+
G93V6hPKlM3K/apPL0G2MUhZ6iOsGkdM60xjkpSBXfoesDiG79iSEPv2DBL8kaps
ex4xWsnQwXbx/D7InFzyYTZLWBcWxnwQhE4lp8LeyRGXRmSrLiZvUcCNXGkFJvjq
gP4xolZOLTe5SiBMzQtjvUn7fbOFrd1rWOB/u8hDXOmLJMvr9tl1JEFsS//c1XtO
Mo8i8AcRlL86GsDwglK3JAcFQlQeLMVTwC6pWed2ZAMcZyFr9htDrZhB4QMU+LAY
+aKuiZpvT1gaWRTBgKYcfv5OTOzQMrTlikoUkWO4Mc43HIJU7vJpdRGL3xvZ1Z4I
twjd6Y2hskvC+ETfq5SGl4xZqHqlktG1SBjRZwIgshecT4WMIu3DEzv7vYauHeam
qmwIYqYoDC3uqdNc4EkCyoXJEgyXMVhuGkRluNvgWmDZcDCRyo+eXuiB9XqGd7wy
cCAowI67MbPDBtrOtCmxp2SHa1GBwGP1HDjkzvhIQ73nto8ZB1pb/RY4lsdnPL0i
RS2WZtXg8jPwijLJrYhbVtkhAfxaw+m4VJ7zKsXnoYpY/7DGzBemOhnm1G1HNp1O
CtFouidgN3do2nHAzcB6pGKuM/p5AWfzgZ01xTSvbA2JAsq5C7CXXqIKswvLHe4G
jrSnY0JTyxe6zWuatXH9TXwK+m25qOLYRgRAngoyldxDPZbtwv3K/i4dl1ypy4HB
gCyTXtBXC5q1GZTuLKHXbQfrfn6CI5yavIrJJX7D4EISQfLtydr1vCxIzNxg0PLz
2yHXZYE9kY7nZIIryorpYLaFTqpmNP+f3eCenOPs6Ols4vL0c8HRoKkLF+Dv2BuJ
E4YZ/LPfLUn9fb295+vqt7g8mWzG0MeIMcdlL66ECbaUI/daYPeqzO0/akUvO0yS
YsurUjjSIdgQKllUPg9IXOneuNKG8BK6ZzYyo70F1MKYmx2f5NNnN2jYhoSHwmiT
vhlRPul/e5I1p3W9rMuszE9FyMTQNk4LngoTjmvcTIPMOp6abbICeoHLTaBPv0hs
K4VcAeQrxZ/3feyEsQdbuj4zgVzjRz0qqfu+Xw+iugIYDT37UtdPRCqX4f5Z/bWF
hI0CkbsBsBnx/mX6gq18jZqCvfVExzTlmQtq9Oa8aKs6KFsQcRPJhfRpT1LCgAnS
CnwHEbSJRkR3//bl89AE/0FRAHr8JoA0SI4bD2KtEwFOotvgU8uFnLY3rWOCmGuf
lZ7gyxP3JeIIhQ9Vs2KHL8kRawQY5qzzfVdPYA7qsngD+M1cSK8IdSoda0IOwRdO
Fb+Br9JC7gcUe8onXZSFXAhxtL+Gs7iAqna3dcWNgg/yThQhUv0fR5wy/j01BB8e
gem7yJ5qVmHq2NzFNozEWpkWtXn4i+H9NAxLpEyGrSGsi/QONmcBE+czLVl0eL0C
cc7uaSdMsJWTh/Ituu0Cu//CZfIGOct8j4yvcfNxxGXuVX42FS/oAmAESLSsPCKa
JukQoNR1V9+Y3c/dX31Sr+nk+zWebArcl5nOnLkAcvDaANmI4R9DTu+8X017ojaS
Klf34WR5DPYaZXMrczfKSxS7wLBBlvBhYPJlGL8a3TdyU+PetyfFZiwkW2+wNiq1
We3Pl4Z64TKX/fibD40uLgRocElQvkF8XCyRu5kmQ4lGqGQGTHoJ2R/eu6Fti5Jo
2VYrtKj4BveA8i7OB8H1epXCNcPQCa1O4SzHwE0HABYLA42XY9q3f4TaYzTC4cwZ
PK7mVn34LYWdwwW5MnNDFfNO+clKE3XrPfcyE3rpK/3dU4rRR9hWLsY6tJCunsel
IReYTDvpR4QO3Z8qblqVg35Puvk/ZlJ4g6aRlCoLAfascLO7miHt+Ihy4YWb4EKI
ZwKgbpqxBiZ7LY4rd9YW1RaLN63DbxnXg20azBnUFKEcPemn/Q/YBsbMRKrOrq1p
uLVumwi4G+rXUw7ZoTMIhp5oF0YeKYRaw9ix3kTD2WTrhTnowLQGuVdAUxrBm8Wm
WrLBEUCeHNCeVHaFGXpU7GLKZc7qJ7fdNRSEady9E2Ut7EoM/dfwLujxkaTVNBOf
2jQ5amYjEgZkCpIQYwAe+7Y0RFhQS9CjnVerOwhu4DMhnai8SMSU4yKZC5Dd9yik
Vgb8mILlq0aMyiIVHoaKRsXtrbS8x16KKpPLmLvQTiGVt38qCbScSNJR1Vm/XISs
OGFDwyRL0iu10EZWtKbYmcqa/NQv2lksYw+4hrsYw0peKKUj3W4/Rt8hFuaLX6L/
VRLJbvmRfdLKd8D54MNd2ayWk6zHnu2s4oSvPHcktkvWtq/2Ov8O0FexD8Tl88py
TjavgdOuccMrdFMZChtofq1z1NFga1wGhKuq8cyF6XLm6u8owXHOmwEGJm24OnyJ
pd4pKDEH5Wn66iUFsY6Hgpl1tolbOYK7YoGdU+jDrr2LBcjrNBlSephYQOdzWNWR
K/dhuo/BeohcutKKCgmkt4QqKwcbRdm3wv8RRPMvPrF/Gqa9C1xFigmsZ8MfDAPy
I3lMX6+ypCdTwCLuuQ4KnYhBX6b/1fPQcsN1gPi23tmA1kUtopRgGu8nAXiU5wz/
QdpyzMR+9z9pbj98IwQVCL/qh1fgwa2/aXoVK7hlxqWjXDF4ryOW4zzxs7XvUpQM
foRjBGp8FcdRuS+AootXssl3jAD4bYarkHk7Lx1w7I8r4lOFZm3QwjiaIJJlpdwK
m1OHv6ZbbuyZSi8rzuhzaArEMa+PoS6tDIf4hB7wjaRZgMx2MtrrQMYDvVnxmUWe
bOslHq2mn5+ngJUTPtKzD5ZbmpbbZoN4E0Ls/yN3NmdHUTc0/EUO2ksOCSeFqZGS
Ig60SckzSoIL8AZjs4UHbL9VWTJtkKy0pqmFuX6kGzNgSivBK5vFpkjSZhY1cTBz
gARLfy1ih6sVD+7BdjTx4FgcMjPLvgyLn4HH2g7QCGJcLXxgy8aAfumZruo2Tff+
8LmkrykWIFJ0XLkNPhv9I/4yopdWVwtBGBq6v6CK9AaeizIui1om2KEiiu67i2T9
B5CIntdHvX9R1COh/5bFadnatWRfVMrAKvNi5ZNItVfAyqzJuhc97c7Csx8FU/v+
dCn/yJ17wJF2gFmXYmWHYtbL2k9RPOi1cWQ0B/vPdGLQOCGQ4G7Vey26KeDdHyx2
3xE7fn9182/QowEywTJ6HRi2j/YrehhZmMP3PQD5SS/RJlR+DlhLT8OSvO0wnL4H
bOKSlHgIa4KQg9gAFpMTts8KQv3DBlERPrGtHYgNxDIFNE05BLZp0J2pyDHfrTnL
pma7mC1Fp/Yk0iFzr3P/1Mb1ELr/qRs8lrRdiUnTuleG2SNKZXP3JwF+C4YCT3pN
8UrZcgrZ/u73/0tdOH34xGPw/5m1Gn71ldPspqqurvBxJMsAIO8TlTPGvjw5rRfG
utiBd3psNHOrozJGBACiOm/g0rnFzH39SCBECzvplVedspECiTsXSJtDNQu1NHiN
mlzxHrciLRefWF1iytjse6dVVadC1F1rmsUzbL0toEl/WDj+EeMlsk4J1oqncx/S
WprLiZiGuejIXoHXHm/y8W0/h504ZBtTAgV+avLFLPw+wtd/gKIzPvtI6e6potIy
UFPo7yvQdcUiTkuFdMq+So6ok42qjaY1A2fFeFxv3blYgUaMGv1VNxOCIyWaDdgc
IeruAYM8TAA9kn6WXJ5j0yhaO5r316tlKINBmLPwVVjUPfU0CdXdjYhBEXNRJbmG
uG50NIzEjF7j1Gvl8+P9pU+zlU9dXbq2avYF6I0CEHrzJw3lNQdTLrVg39AGoiIj
/8QXoIrkQeJ9bzgJOyrLgk6Nc71mjZIhqZFodkmtIqz0hqO9YJXPpmugNNm1b2kR
vr58hPLfdYvJP/iCe+PaIGO3WfsIJuR3HFV9DZEjwUPuRI4PvbYEDFV39eVPYx5V
PainAljsr/JjySh6uOvNMVlPJJT3V6uh86rOIr7yJWM1lOijYJ5LyEZcalqqXve0
/6DQ0HScCVkxKCupTZIFATtPX1JVNgsewOzkSIsA7yu3XoFbja2zdJqItF9atCej
9xZqEFoPGx2h9HYvyoyOL4FHmmj0r3LFJLTfFgs5A/mbJW6bcV/rrW6Jndi1niRK
iJQSmJzORbkK+OdmMj9fi/t3QQjvKNZMjDAEeqNKZYWSD2vP5RaQ5+E56WuAkZsU
0fxOkYnpOAfWukcAvFJFS9JHRiC/5utPg3TzEHXEuHWXq0AzUqUZjKv/P0HpaVKZ
ghQgXzpRAkss8QEJU36OOYrs/ttX5n6MEd6WUfqFmyM5yQDvjqtFNsqREkYEa/R5
UgK4a4VXPY1IfClxMHKgi5d9/UgVwB9QKoZ7Mfk8pj/BSQ3iRp9LAl1xJYVQu6Lp
l5uzYZaBKaS14QTgfcaE74ksINgEejFFDAlB+HSDluDnUoo8/HwLpimijSwEaLtJ
EcGcAiZyXfcDYkYBV08vfFjkJ4kK+inoVUoClQsCTbBuvj+1u6OUsKEXHA0kHpsP
9FZluqi23M0IDa+Cwd9Me3IDOf7jVl6W30c9Mx2c8wITW9sRqo47BiVz7EwrXtzl
lVg0htR4ADC9tnK9uH8fQL3dHpmRVspKzizowuVwc+IEwQSm0Y4zjfBGuSXYdu3j
Wdmykg+/INiYEP4BI8XfwY+KZBlZulnjIzkt43AzRyyiMTz/e+VNlYpuyn39FsNA
Z+H7osHlKeEgXhBUEq5iQ9tw8wWntIzQAaK0H02YpA0fbGvN6Hxk1ZNBBFKwfRMA
kiXCCbLQfLzWzmE8Vjro3x8YqsEQ8tAWA61ezRdHvIxE55iQ8XRRz6hQtLjjMZiO
qec/8tgD3u91QFB5esDutHRfVI/I4dXTmRmFhaoJuwYKtJU1ALKd1tLOvlN8YZLK
LIqdJ4jf9xBj+uT7iC618zgXsFa/L3naLACvZ/GncGfEJtV3JBYBVKYa7uXpXqx4
On8UYruDKcslS6nMun1d1rl5XOVHcw+447268MdKdQdHUsphqvLtetv+O2xw1DkN
9/JooIvEKg8Z0GTSPSxT0DFg0AbUmvG3I/TDZKCZIZy79dUrlc9xIBsA1XXc1Up6
fXI1Nltab430bpaNzVsQoWNKdsXAo9gBhTn5roeuZJzgTW3i5m0PzxIRd0B7Vv3S
WjKZOPrW6LDrZT/mESl+nJ23P3gseTAn/9T8H6ygbWVmaITVNRiG9/dj248Q7+xJ
giv34NenAs60IynlafQ+lAEQlUk3qfIykbtGR6ewFPl6RaOPbzxKwrqry0Vn5oWI
FTL4XVR6WS05YEP1i4ru9OoFJlYNrZ+fnRmfaGKoPGvk4Pzh0f06VQtXZAvTHhMC
HT2h1PHsLksBHeFu2s5t3lWxKXAX1lyTcMhmEuJxt62ykDUdLkBZ2b1mp6X0WJdh
dOQSHjwaKYtDcqTTUYAwGRBJJiLOTIDfEaK97nv3V4MXdDGVoYJzDY+AmOuECJZu
7SitSdiFsj2KjPKrFX5SZtGMfYNKKC2v8jhLvSzq5xCVc/iy2h3hFfp8PMgOSwo5
luTQwE93JJnHM7DzTQ4dc1cLRkgIg78nbuwsq67Mg7ZvQAUMdrdgIbU7GdIUP0Ja
chxRw2dO1nF2zIo8Ix0pz5X7wBN8VfrhS/DGKjRiZtHyDDFRSaJGakF0Lgg7OTbl
F1kArrgidw5DAkvDPfL27qaJwgx0c8nTnrtXl7FQa0s0SKlPL9RBGe/1ObIAJMwj
R92SN+gWnp4x4VygUBosbRQUIH7/+utjyf0CDiXI0XdVIj8l3Pxr5l306zPXpGiD
90k69Az42a/mNr/Lt+SHBdkIS8ODk9n1IFTiqEz0pnDOO4I+4pOKgDJMJWTDLgT8
zTZvgbatRS4wLyVmmeneR2Ju9DUxdCYmOpd+hc8PyDPiYyWq6TlR/MIelGLCcr2W
4RGYBcKlXgbXOKW6QBANaiUuQxzELQbBA5goSHVvLvhvI/14/K+17nZWUeyqMogd
+hJu5vyPrTzKrYuazUB9C56ol4UuCqxJACqRK9NJFSzHNCAnmyojHXiV6iqMXQel
sSnuxseogZke3Tgc4i0GR1pHXteVh/u/5T0Gy6FTRyLcirovYW2R4YU8ysbz3oAc
8LF9lAXrDsiw11m6YwLXC61nP9aIf/iJfpLQ3OtVbH137MkPnpZ7BSlpRuVQE9Wy
G5MZcI8jV3Hf9nj2+LMd/XgME78jKEFoEPfnJq26O+eSctlPVd0NfANNDB2asIA3
vc3X/j2StXD8ZVbh9Rp/f/gqHFVAsVdxGRK2yOKbLMjVR+29eH/XEOUvIop6P1MS
9wJrtfC9tdyudA448P6AA71EVclTSjlDHPn255k+43KsAdPhMXO0jVgF2nc3FB3c
47hHN9RPcXFLVDIOelYHecaCDIJfopsf3/xFioA0c6zfFqYhDxKC3RaOSUq3/4/B
SvSmtYFBFuRALqOiheUg/1qi6405IqOI8/tZL1i5ecv2f4YHMYhB9+VGk9+K0PIy
G+0EvLK7s4ch9/sJ+ZNd0egyJcNOhuXcA0YMqqLVC35f729C1iAkmlfmBQeiCtLD
suz+4R5TeyIHFvjWU5GY8aU+drVHKG8LdLI2MVVeJopYnMOqOl+EMTW3EUj5RPdV
2Zl2N4hbERaj0bRFkxt534mOtRHZyzyJZnrFe3J+kkDiz5dyOBxRnbZvAhB6Z+nC
4yuxjSsSD4tzOrLkfQvz2ABzdEyKXtPg7dU/MMisMm8sCWado2w8UTTJYOkZMPEj
4SGph0uRxw1Y2bEbf0XLqX//jNn6barf2qW7QwH1SnHKfHrzjWFUbQnU6vS9nPlg
4uKh8bMSAhiMWO5LnHn8iSuKjfNwguj7zbp04drPtkCjdvlsSnO/xE5+T/gvWpG3
LpZnDl0+gMYN2khsACg2+54uCxe87lwJYz0VWiKxt/b2NFEFYdnM0THlXqUkJyr4
zRyVc8URMGZXavf6VA2nL6xuFUZpXlY9TXYTgG2qs+2exrMN5+vpdsdJeyPkXlH6
Qsu9h7rKxQXzv15j1P5eMgaSa9/FINj1xkYKIJDV0YB8ZI7mFAs8bsLbG3A5iHJ6
pLmgQNunC1mXozoCTS8NHE01oSrCoohTtuJoaRnVQe8GbZiaTG056Y/ZGa7lIXQD
HqKVdn+OHCv/l5HmBOdN+SNbzNUAmjKzP/YUnorvqDjABe/CCuBZg1KRNlRUBKGj
INoU2A7s2KGGkpg003ukN4rq2lToAgS3Yl31Rx1n90N6SGQFjbRwVxVkgCWKpovz
OUdPZUBxUKwmKDUEqgpfUis2ZEsA35QP6vtCjiIJmCxYh3zGI6NmOYD554TGAtij
Mb7lPrZmcq4armrZHyNwpSsLa7ozYATdnELv57fuWEFIxDq+PBMDgx/UTg+4Ul2m
JBbTlWZifqRA48GDy4Jn2RL4QawrFvEHgyFEQ2XMMD8VZ2CeIJmmTWjYV6DR/uGe
tnme0/JSFl/otOVLA3gXBdcY1NSV+dDbUkqoudIBINyOtm327U+7gH046hyjEsI7
1Ay/5YgCepSkw92cZxeBFfYCJsfNB9yPuJf/wUr2lnKR16/tTpAWZJt9Kr+5AYo9
3VKuVgRp8IA176xT97GkxAXI0B6bEpBuoHNcwpMUo475HvDFTr3dFeo+/kZKOMF6
MP+SkRocAyUKfS0ASOnBxgMLyxF2/GGnJKid3xIctS/qR9DuqNTtG9UWE5N8HsnD
JY4MQIwf8va02F0AGouY5oMY83szRzMDZG9hrUZxDD0691oDLrZ5OJlIUzuAxsaN
KonyDqNfRvYjPX4UXedBR2Rx3nwVcXoAB4dtOwN/v8kxa/SWkJntACrobWPpxK76
Zkx0TlZZajXiD2DIJbOxNJriwNSKNEZtIPxsc3KP2okyEG9U7fV7Qb++zvOmi9TH
toxaKcfzVrnFm7aBwn2x+7uzpg36AN+x/FfUfhtSnS2nHNjvMgxIShwj/ToyCtj1
9UwGZVwt5OI/vfhjB8cVQILhVFd5jy8MesgEoixG/n39rB7uM2+3V6FPuKpy9lQ2
Sl3IwbcDkUfljPICXdXr6ILY6hndyYw13k0U7iTagVt0G5GxML2dOmHH4gwXsA/H
CLh3KlIZzneQudGA2nPOQratdvdcNE8sCZDwSxkOshieKBE//RSeJsavslorpD4E
YxKiQbIgQ9+NX400dHvxT6kYAUmwr363sD7CYqj/IrOBLdZgR/96ySDYv5uiTb17
usvJ5UkW6pnzXndUxYaGUo3bW085bKiU791uRXEY/syXalFZkSnxDAJrFaFXKhfP
prrkBXBzDGucIafT6GqhQhjEOkUNbsxdR1hhnex8zJAuXHoqbfQbnVaRrAWc9uaR
/0beqJ6p3Xrd3PUfkPz9yYUjdyCWpXQSCEQL9voc6+LcFJmPPJieMd3u7ucSWilv
InBFmZ+KJgUpna6yRyc8Pq/uaGsKUs4eMrDzZWPJtZ2+EDiIsda6emjJMVuQ7TLN
0O+zVDUfrxbULaY28CxMSqzQU/pa48JSoH1K6WFTLEJ/NuqRR5QI3K+I2+YAz9ot
Htn/xyuSzyRLhq8JzpF1B8cgygE7ipwfaJsNy0WQ1ddL6jBCCM1c4AkqSFIcaYO0
WN3WDvEosBwz6y2ZEIX+YdLaKIj4sPINpPYu16doxrR7WnTH+NfSHUPwCoOBKBas
g87nS+PuPRqQdJjCMgJHQI07HDNElAZy6tAj7utmsn/3rl+7wS9vBodRhtkjYnoH
la/hPLgyKtvQTPmgkLusOymqsYB6iT0piOvM1M0z558Qjpx1yPVhJhCHRoxuzpqL
apBH/bh87nzUMuTz3eP12ZkYaoa3I6bE8BOIfHAY3o3Bs1hLq2eZlI3W+zAAISrn
9Q5Pm+rSNQzfO8h5TvWcEpVi2kkNuJ1ATi+qKoRkXN1m7p9+NwZuGPwcWIkId6ty
l7TzihtfsijICSy+heEz6SH02uRZJvevadWtJLVZkuglip6w07kBRI3QYtIcZF1o
N/ZFpMsHr9ndlQ8Pn/ngv4RgVCla+Ml5pKe2jshUdJFlB7l2ccBR8NiAI3NdIL46
f98mif2DhRTPyweLlxNDRDXq9E89VAFSCNmO6unxrroeSSrr+21a6/esXwx3lRjg
l3p381rZN2oGul8fY1SXSa7T8qOm1qHbOWdJeDx7UyxH+gQndjHLJOWhNbdh1e4+
nMDfllIc7waWl7o6oqyKE3akikC2n/nf4SrGzt9tyX7Qk75EHGc+JQZmx8m4J7O0
9xCTU9tdqsqdx531F/CcMm0mj7iov9e/2aCdJB42EbDBYbIYmeQfbkeMhuZXMBn9
4k+Q3dVtwEq0uqXjThVEdEfTpjG7QsRkGVI/rt6F9UlaRHh0+jcyd3J0w2XulECV
gam7gMfyul+NdloFQedipXRIU6QKSopJ4KhyD8YzuBly/cBta67+Ig+tR5ndERxX
RX4QZDIKBKxgkYhbFQD0F1BTFBpIds0mEvUmxnh/FWUITqzzahCN27xfZjc+L7Dc
3WqXImOgCj202REZvh1EjdoiHlSc04jwZllEnchcLFanrG4vbGyiKwLZa3JE2L7v
5CPXiOkka6uustdiLBvuoaUKT6yVMjQw7eyhh437iPC1hGjbp1L74970XkU0XV+B
rVtJXKCoZgnO+Zy3CwhnTs4nzpKWXQhJjj9mJCy5RyqxSDIXxaxdC4KyKPQG6bpi
5501zPkZ/vERVFUJpp2+vfpRIlcKopcbB1AlbtkOVCoESze2xU3PDPX23aUqSMWl
XLSX6W9OmvzG1KLDgw14RYiRujxfUHT5mcvdnvFq4l2zRPkxZMzdRMQy2KHdKZTq
rIldiKm6aX+HzPrqRHuVGuE9XMFLHXdos4a6qbtOf4uruXpT/hGE66V2SptKEllt
/o2p6MW1y7wbYGrbZWZiHpOWmF+T35E3vW/l515LdxWVvvPyELBhIXxOhzeTH5tC
L9shpu/HVuuDuLN/6wk6Bz8UOVT0WQPvt+ZhkOo+TaBU/0E4MGWorgixwrLLt6Z+
F6H0xYcI0FgKDwxEy6s8pFkWbK8/vLdvPw1fS77mhDn72o2NV+G8jnBVKzzuampN
oVI5Qc8y5X/Dh0hLGj9edO+4vK656aUWsxT6u8bEuUUx9xlgp4qvjX/Fe+uEWHGD
S5XZuknVht3aQCaiVLflGkv3wJI49oQaYYWg6zaTFfNgjjw0uQ3YMvlTcL7YE5Hg
mRw5tex8TMWk6RQgz2vN/8eQXMZq9lEhYjToW8YPfWbKn4t79ky1aEAbAUivwA+Y
lNlnSdXq3aSoZqhonVI0PHKtldJ77VMKYLzhgDkg6q2oigwYB0ofRM7wPsrljYPl
OYIyroWDihaIPx1RZ14L4TPvnemSF8mO5fDl7913UmZL9fyLnox+48D94+dVWwSj
Pb0enjMk6i4ZapJ3CtcZ/WeqHBAMkMocMYTjzgUsukZXmXaqUgTaqKsobH+z7QOG
Ce40kMFn9blZCR+NlnxPG1pyVYnzonGzaStEavOzCVYbM5ysX8XJtyvXMh8LSJtK
hlXKb2QFUsGnaFCE+AbaHhBJTBKL2Kwcro/Go6a1KKjlkfrC2unfMX34kEFykTsf
UMsBZFWqvv1u5o1Xmv2ko3FT0Wjp/3bMdujNw/LHKd+KaUuKnwwyTANIfiBMai0a
Gs6FPmwcHnebxm/59ecuGrN0d0y/wznQIe5++mXpmEkJZKc2KrQ8afuY2PkOWjBq
HGOahnFqES2XblhxhTpLiYFdPzDeB+671FcIp2Ndd9AkdKTASDVoJWHcOX6dG0BC
Vu9YVZsjVew+1mjuRZEG/iZc01KIw5brVTVNZ0yyVHZBrwp0dXz6y20TtNAYTrwr
7ySbNArCFk4S8FBesJ1rgB0rdFCt5t9W6ZPwr7UalUnP+8U2qgb+iFd6b+SjyCh3
9/s7nOLVTtKDiYnx5SJqFIm84I1Bj461BPsZEUrLPeYbALRVf4Tzqhe/o0wytKZA
mDae7zgT8TYONrKmW9N9V66xXsZlwn6QRWlXJkX75eD7X7anxbOcc6+JL7mb9lhi
qnFi2HVa1VnI2Hnabhud8JPXQYHSWCb0CZyXD6eUTzVCVvprx1NiV04QK2qJzMnB
4zINuCZyPenPfPMnOlgbTexIJCloBPdagPNloe1QGQ7Tf8UkfnIQMz9AM+rN7CRN
+F48dao5oAyVnttPUO7yWu60ZtfmHopZRaOqwPrQ08stY2NaEIwMo/+HPhicghRS
DNu8TrYA69e/d2VBiafUci7/67omzo/eizsFFDr3x0EQsBaLZ6j0t33gpcX93ySj
SQ9WKlBN7BZbgasLUd/KDYhU8Y0nhQ9BJ57b+H7Q9CdCtJFmvdPKLquoP+BqA2kd
MDCoS1eHG9fpro7D/TS8tmhyHLVBsCOw1y29ZMkvQUdodSC6heaKGNsU4KSmQqLs
w4Su+XWyRV00WGkfX/dtz5sO4r9bclwI1iKIPAk1ymPp/gZujQb3GfAhCi+gzFT6
TWd9iwuH05oHnfzgof59SFTttR7T3K5yiES3UaChnImOmGpJLBELwGOVi3YpzDv5
ESKFjjt1+WZk/CIoPqLUDGvRAWueKASADIyuCQQhxfp/KyLQZMIp2k5QuLPiflJd
CsSlWlgNQJCZvXTeSxDe2ZhLsff4PbauuGT+bgUapXfeSlOOKzx3+Wp+qxKG+qiL
bs3BGSyOz4zw2XBw7mPea1osfN6CdmQ4bnqIZWudhS/jnZT12brgQFOYN+HIdlrO
1AAM+52nxmF24MH3qpXhuU3CczcMza9QwwPH5Uy/2znP19HE9QJLL3rz93LqHC74
j3LLCrnJJ4ya2Eh9LUuSrSJB+6LyismwhlyyR2FNkXrwDOr/76eEq7ETJWnNfZ0U
IeM7cQEB5PBjL9UnOTjoKGOk99RkkLecIjyFIwohIuKeZU+YjblBCf2OUbwnNClb
a9ebWR8gTd6u5Inc+KEw2FU+MV6ymSYdJDRvC5d6D+VisSn47B0lAn0LyV/L9Gry
VALEQx+yZu6VFlMBci9hWnNmCW3PitYkfzviNrSmFtlCknVzV1vACbBg/O18dITP
ThfFS27jTaK/2+v1It77fIAkQDRHEWpDczd91k0wftclTMi0cxrGVtYhw6wC7AvY
iKCCu1/sF6xAlMkF4Ow0TbaaXnpRKTE+0MY/iwZwzSEanKigpMw/SzjdnZ38kkNT
unxnaLVvtDzdQyDRjVx+T+zvh/Nq2/DgiK7Y+fnkDfcHEiD7lKizGRiH5Lu1ugEA
hQyuyxlp2IVY8QwuwjIat/6fMhauinIqvoO1J61YYzTUedsBhRDscKTZyigAsZbn
dfk/hvqbhZW27pc0EXs/iXCx17DV5giWE6AImNgGcMv+b4G3ouuTGb+aOjvf9idw
M+xThELZSfd89mM2UUZfONvyJprBtSvwZy8w7d7pfBbuxa3goMBQnFb78cv1M5QA
YW9EOCnBE4unZYzI+ZyCGZKjfHAYc6qzq+HwuQDUiONHl1Ij0tBWVucGySOAzRaz
jaawk5AdTc1iVywDxpz7AhwIVRe+LM7/JsRSVSVpA2xlOY7xFprQUakIh7UAZvPI
Ymm/BvsgQlpernvysRIwKLlOjb3t/2PM98wOEe5bgetS9JyILG0gCfmlB87hM3l8
SoHqzWSBxU4WS8amM0s4yoFhrcu+TwmHTGrJApPjRbulOeL4vdGtmVbQKbwgqiM0
6n0DdUPd6s5yb1x1G6/Z4xuXjlVm5Z0F3G3QZXqshSdKiiFNZ+KONmJp4CqQ58xb
exxClTUyVz3HTz84pHYgEJNBtofvLR4uJxg51ThDQNumj9pytJDNiGL8aenlpls1
rsdHSBzUymsx5EKcg4zDS6p+2ljfMWnF0QAtMS97mCyRiM7iaDvnW39TQYqHGPZK
vsUa72RZbvpVn3VvZaqRXjJ4Opk2VG4a0XTca0XpHcDgO3AOZJ67U4zpai6f1z/f
PNZoTiOCTvdi6ym5/fueCjf/5IAatgcRX9Xrfzu8QhA2LIpHwvLn1gJGkSFJ/ELd
LS7rdkXbj/RefCqC3ZCM45XHLThSAn9ZedQik366IOuKGj0+9ClPK79FXqQRx++Y
7t0g7P29p5PHSY6wmDiIwn+Bm48Tt1kl2RqscBO4uZxUF+kegJhM0/rHoJrrdGbS
GrkyB6dgux/rD37KO4jKPap43H2Q9+awYda8NKL/so69+fVx0U7EpA8wq/Umx+cn
qapHgHP419PSb+yTvZySg/oT0flz42Q8EjKcPTm8LEhLD0lAY46l7Aw8n6Su5bbL
GHjRBzhv1/XFMqg3C49uEEeeRRKs7olNlvyD19jcPIQIidpUqoSCOl+KWhaupRFY
PIEsZTDTa566qggfhObeUklJiOw9g8+sxFlCOD++HWf6XJBbsW7QyDEZBcA0D4eX
I32FsANL8cx7RMbgmiyx4ZVyBB2YPivMvZBATjq+DIpVp0YJTM947Q9nxhdAmvoO
96CAgjbr0o9rPmlHEavB1mYp394yjW7gKCkkW/b2+9N5HYYDgEM8tIf5nPMhwpSX
aOfXFnJlFzdV5K2U59vSI9aS3X9H/zS0lFxdha4wY01+w285z5ygA2fk3ORj5Yki
HIRLt3R8x1BRqx4gnprD2dg9oqUI+afvGih3QZfoopZQRTDGqF1o+Bw4fV8X97vf
3dJWgcrpA35hK6hWpgRSjgb04O9PnmeMB8Pa+O/QjZP1mRdfHrmGKfGF/3piQpCn
3QXED5VHHk3Denl7rMleWZ+FiBIfOkqsekzwoc8ycabLy2RIpeO3UOuRTtroSWHj
xAW7PbL5lRIwpj6tnYcKodEDAc5R5TxvHhCsR4WbYaoE2Of9zvOVfTPyNxain6rV
0vVNotuUd4tHuCfxFCjPJ0RznT8NmNBN2M6gPtSNNCzNczqHYqidwF6BofamcZyW
4ySWdusJtgsuQcY+5RbiiH0vX57BhgmFvn1hqwHuktUC38Ap6DF2eBp4xPLDZK8y
1FBzBoWYYPIOU+8g2uy8r3DWv2IpMal2ywR/sEnjez2ggsvtyYU+lQWEh8lVCsSm
7CtcGpXOrDyWnGQ1Y4yanymhO7FcS6K8hoAgFAlsEUvYpMneyK0JACJq9Q85ducI
78ctEU7hr/ZFJp3fbImuuVSqf2jS9t8D4dF1VGb1FUMfhP42ujrJvki/R+9TS3IU
8gHty53vSgHd1csh+emrCGlxISeRjaK8cgVx6PBRBUpFz2qj/TN48IW1jT6bKINu
NyeAMETsSnIVoRaWFqFhXexN+cX5bfQt9HLqyqWksEgR67Z14ABQk3f40MxjNBEm
vrdVyLTZ+IyPDCqDs3xhgh70YXKJ6muht6nyQaErcyXfZHyHhdI4SXh7+KDB3Qnk
JwLHehjphyqIiXezqj61z6ivY4REKhKxmYpPpH7ZeF6mLHZh8IVOt0FDF2Un/HG4
X7N+qj5+tdqfDj4rhEPLhbWVk0ExfhsiggkX1mcO9K+Qg1N1sT4ZkOpJ1VVWXBze
dOG9PZbIIj6cvBI0EzvzfaInSS1v0sjimXISGekgcyYxBjLYao/Z1X4fOQbH7uJ0
yewJ2Put6uBPmhvl+axs33Osf2Nr8neGtSrrR1yxPK12QVvqdVIWa+sL9YKIsc7g
C2YBVL1I4LDg/LQH+G4nTZ4t7lf2fkjDMAhRS54UsP+cpfdfTz3HTgoMzmGpFuxS
c4OJ1dK7oJzaK4uUJ5tlhbn0g2ZPQJzSw1oaiGdqAw613DOJ8AV/bUgSx/9zvY45
NnjHif4DDMs1c6OdPPfzvpVeHiuExzBRyA3jSH08yVObcuYcFmRG4mI8WxWXz5G8
xYsrWyT27HkaXxBU08drLQLyAPEz4UWRwzQFWPN1OL8OgATsWTYrI7FlQqvqe0Vs
fXU/tdI1pp06WvEfPZK/AE+VoCBGY2R2fPH0cWvVk4ZBqFGJT/wtFhX3xPHVUqLR
4RXAfdmjVodw0Ikkqk61wYDjT2M+McT1B2+AtT/bmO+WspeQa2X7JSCyYeZijJur
sfFPPcHADIqRgFDL1szvGEmGNJiSs8Sj0Hgc17UjflHG0akUYT14QMV9vg8NqK9+
n76XTAAaZDRdZXFoX3sjDNgRqQUGc3xZ6UEEbm0WQbfonyt4XGtwzz14pYIpU1dR
Qcf7j3cpqrL7zEdH5GT5a3UKattGYCX+DOB6vu53kctPyETewtqUfUx8Z2S/N1vI
KvZFhzG+ISsfJPfHnNX2boAxbBH//wjyeAHwBBJ0fAitYTMQGnDCp5GMd4NpGJh+
uJZElknvpcU4cBmUhc0dQwIIP/3mGE1s6APnY+CCbTPT4z6A7i2rGvMwmdEONXsL
ihW9YDV/gt+dYYFbePBUf0wUGZF1cBM7x54hYjZU+El8qExrMS7U2fPLpIQtSmRQ
bKMQ+1HRYn4Is8XCe2C2L6CyduZWbkZ9gzP+1iG1Nehre0LvrJ6duVXg7usszw+4
3O7XuCNuIWkXHqIfKkXMSqX6iF95P7w3nlKP0VnD3/Lqj24KhCth08A9m6yMtg4Y
u3t/DD2CNBCzCF0ovWUFbCF6ODyzcCfYQULnIStOvJgsyXTBh24yVcvCBvwPk640
dd2NIGQ7t4N84IPJm9SCAxJs/uGbQb1bAUl/q/JAcOp/2vu/TxWcRV92ZySgBzSW
+tRPh+oAWZmNRuyR4Xz45XKbGd1t+pxFj0wSo8aK5Wol28XcUn2/WSOqBCnT+Nhi
aUmN0Yql7Rr5tbXmfIxKRwlQtpfW8ucR9hzM8Cdoo1VccA/BgaM0HMHPIk9Y2k9P
RmKJLIEyxTdGRHg0hk8SbwfNmSVN0sVYMUCDv9OFqCLhVnvAROdlalYlZ7Mt6ktD
xB9VFG+n2R4TfvVaCeHPdRY3kWRmLgHgUWmbnRHd3RveC3hAPGmvq3Ho6S2+e2Vj
HLuHXUJkoJpY+xeniTl2u3HERx5GGVZBQ4+5vY4vsayrFegcHPgDeDxyu0fpcKLj
Zt7VXptNzd6AZ2GNIDju21eiCa/uDrTA+x4EwJACYoTZIsIa0R/RSFF+TgNUHDBb
3Yd6wYCNydx7ncZ6Rr3tdIqxJr2HkyZlnHCyB8p5YQefcqmLW2rwOmHDAAlj0HEO
4h8kydECxqHGPAQ5KwulXYUpN2+vizbsecb9BxlUn+2hr2MtopsOQiJ0Nzov0Im7
lDHr3EYSJDtD1EIAvcuL5ymmMUaTt6Kc6JfZQSaHNuZdfUEhu/t/GQTtiE9SIGdx
7bjQ3T/RIzbzrIoakBRezOuy9SsxDD0SB6zz+Aln2R8FSb02xU4WGFTswtkcsE6O
rxk/Sga8LS9gVl68/jJwSaq1X/TNXFTU8g3MkcAxtzjesE2Zwi5iGyLKw7WBwpT4
+Azc56ltf0IKDdjZJb5Xd30iVXhkLTqijM43GFzAxd3Qci+zV4S1hfIZd1kI7NtB
twCWYsdARigJ93yLGw7JRTThz313LwkteJGcybR0504ZDcCF6R0au4E+JLmG1H2x
9h4SELlBSRZwEMcoOYFTbVYoEX+Vd1zJ1CovwY67mGUuwEpl/f0G3kK4QG+66GS5
A0kTNhPt5UmQtmBK68TCMLUE6tA+tuIQWeGgZxhWwYkINzFFdlErztR+4j5o2tWa
xK0BSKEn3oOC11D/J4mOFXFL9ru5bW61iCa/HS8qjxP5CgW9F5/2H8K8xuiZEcUf
Ub22l3Ojpg8Y+B7FKhFWELbyfP6cBb8V8dgZjkEsNHxeLx1VPElbrzR2sP741yIb
z97r3tzWJFOgnQuu8cr9tZk30gatI8tX82MVaFK8kawWgE/oylvrXNOKnQjtGa/G
cEunSEqRbilV7D8zAaunwNOeiK1cWsnnah0ADpjlKpDLeZ2cnIO4VHKA/KiJEnRJ
rfawUABBxh+zFiKpBSYJ8IKxFnhyNBg0fmz7snyPSrJxGxiFTKxc6uSGoKj5lXPw
+Hfe5OibL1g4rDeaCwV4X2hhHXmADDeUxvvfxS2PgrXhtaOZJoQcmWK3U7Tm+vIm
rmYNrhFqOly8Wgm+piei+nA/fT/u1wyEp6XXWW2IzJVpIOC/acdpeRsXtAlTAe7C
7FejgCbfyTFVimXKs9dWihduBYoFLO5ECwvDqr/wuzwl5bv0afdPYMxejH6ujBXf
ktpC6OMaUkC415BXeUSAvBGA1nkFkp0VLHA2NapwmgXnVB+kzP6gzQeIDLgm5lVs
lKbo0S127SdfFogb1+3OqlClXmVu0h87bFKL/KeXyJEUR3IL48zBb5PLCHpZ10k/
27/ZSnAsJc+3DDAkxV1ynSzp1yJZFmf4mmuLf7uGjIV++uRgKuYBqQXSqBPH5QNN
Bj8KfMZnJCuvbcRLjiIlmjy3RBUVF5BaDK+FohnytAlNTdvqhkUnTqbvspje4gpj
SfoYS/MfCNOFvsuwkiZybzRTq5qev+r7/oR4JNpUPUCsHZBy4OY5Bz8uKCAqMU7o
njIpifqyD6NthisXa2FzgulaPu4WGxyuktoWS2jxvjRuUmsZqa7WvSyDuHDIEvyf
ErScYWChZqda5H07oLnEGeWUMWICuMfkPdIvsFiELmOABNqFGRMMcTSE2MROvn82
FUfAPcqXE8TAJp6ag9qfVN4zWm+0GY2REGag8Y4Zs1YQkeT0lK3T7zdIskV59k5g
/eR1s3eqpPu013fqtw1JxVQqYCEKotXjnkC2wMQKVsjQ/pqBzEJJQwcUHLKuTfFY
FD2hLDCoTkIoTkjDON++67M7pkUUGv9KKbUcuh4o/XBjNMuDZiVCZN7C565ILpZT
XIuFNSTpdNYb/IgTTk0bNefIWwcW854p2yaKHJugF91kCNhOJX0DY9Uyoghj5/G0
pSZ5/ti3t2CSxdjQmiBKDddVIFbMZJzNv51itEstXM3B6cBmhyJbdzAjUY/khM7p
/1jb1lZU8NMt9K3pYUG9Xti1K8UfqlZHztacYTdeoWTIuvqjs4DW/ZxLh9bZCVqv
1NDYY2Z7Rru+NPGsORKgH0d+Eao/zbiSRYHl2rPpdwgus1ssWSZ6GviLvaA2fnox
DOH2zqRPL34bzQA6KUF3y1eN1UM7ZXvqOQT9GBllq+u2soquPNADIZOjhbXZTx4Y
xQvpzXat9hFF0l3rUAaTyZ6oDjy9Nj7M7+1DAxvfsFpZkfj7Rl2kWRKz2O/k8q+Y
Nr1GnOy6rkRdfAX7uky/yuECVOm39V7HsgfBI+OuBXSfrZrZaamBH46d+MbIIAY2
9t+GEeMyM7O/7DmXbgo2CBpnR0saEK/SAZar8WmXdmiYOU6EtAALGXEKea3rvbyL
xUB13WrcxlFbuQFfJI2phTzmmE64r20dMI+N6e9zaGy6iCM7DD34dfxx85T2Gjt8
Xvr6aXCucCHS0ayoN0SQONOXw3SQk3mVCdZeD3fKNYjyxz3pyFqvQCngaru6UvYm
ZebiOrTuLC+Wu1xydIYcjJriXvGW9lqJ+i+SNy5o0ynkx1xoVYy/Eak1kbvrC8dd
VZioqJ4wdISWZZs7PjbpgnwpQmDardiCTWKnaO7LHe9LWqm9ex46pIS1uphCiL9G
3T5y0ZIvULw0bMzPfAQJSRWNiy6naitHTzOoUUZdVOC/R7dONF2FsUnX1dE0UFq8
G2GISrS1X7ZqTutcO6QITh4Ak14RXHH5lWZ/+fFeBp4O2B+wjynkezDiJrugB+aB
p3YchVSegecmYisuspVKfLQaedx/ICclmaMZRofXOG9Rsd84lEZcgxN2LggPKptw
7obyJXow1gupI4MlPnkCiJInx1cUWeaK9hki6wRmrJAQTpaYxPkWrql3DheBb6KM
+QzwQ1WwrZRyVgcp9VfmZBLxUC6RCSDWQ18cjE/U/hWcvkAQ78VraJFTqB0aougt
SZLn7Ee1Vv03iTfVNP/adsmGUghIW9gXuLzHdGk6qsKP42WQWwRAcDHx2LQC6Gf8
UU/GckxmIo1DZxeVKq4VAOGlSb9CBhfv+JkDlYzMyIH7OugHpHCkQaWbnW6IsmiL
D2AwLnkLDbNdHZ0LVkQ2AdtzHdBTmpyc2+XBPTob7/oY1981Rdfm/Osc0wVN/A7D
ZVMHInhyicPup5iPuYL9VBf9e8bQWrCZoiDRdckliGrMcd4BS33HR7tb30zDRDCS
ikySV1iR3bMVw/3XuxFZtmB1B51BAPdForc3X+XFQOTBtNj70owirf3OebBrASj8
G9ky05WtAaPQq27yc51iwjD23mcRbZkS96A6+A85ggGoU3L4WzT7qQDY5q32p4jZ
mffqz7yaFbAkri8ZA9jMaAsdDhSslEvmUD3mBVUG+jTeNf2En9iNRp+h1p5oHttR
oplWgW5tqlM/DM2Ge/E/xFrINpS2nrSIeOlO8B9npl5SyR3VcAivcMMROYjbBb5R
F84d1KtHrsJquMAvB9OejvMspf0B/7v91wQdWZM2X6NH4He3AzLtd0xByYvGaZWy
SriJc7wZvibOAI7O7XkniaPKIkYImXnlYha2XUyg2z3ntzWcNKSETsMO5KWjUpiB
+06GIlxNSzxFQNSmgNUsjCDfLJWSScPl0B+HnMPMNAKf7piFiTio+c7UOpJrd4zQ
g6rT4XZJBQCCZzi3WhNl6zsGMTLpd3zx9clbdeef2sxxrXMzhLRJTv26uIvvV6yc
9UecesIoTAo/lTR4e5UjGUVV+qswsjO/maVxTcvLwamrQ95SlXbj2kru1iVJXFxg
OKPwaloJ6HClq4njW7TEnwciB75hAGZckpVXEytdJIIptk0vJILILz3qfC15TVtT
2RweKdL90bptmgpFFXfE6xba1/9DZtVe8UcZlPh3pS7pNvRau1MoNJ58/3PMHKdV
X1zjtZj2ekz+IuMpZ78CCmNWBc4Wm/ivuRQLOz6pwxLZNL4R3Yw1/s7dfvTLqX1K
t2szaPGI25orm1VPXA9Rwqxh5Pcgqm2MCw+1WcN63715rKQQMJfo4fm8bz1VMJWZ
SdTFj5JzSLceUVCkYmhUWCwELt4jlDm4yGKI1LwAN3BfjuG/a7A9P+E8UjZQXoyg
OILwN77szFdj9ggzJ/ycl0rAzRRHgjlq1FGNuLhkEFyiHOpk2FXvw60x4A6xlMPe
rw5NZ+OYrnqV2bG7J60ZFXDP8iqzOx5q+ngsMZ/dH9sfBOYTLbQi6Qz9f7npsS+n
dBiRyjK2jHKxGoDuM8rhJ2ZlBB94gIYFZdkRpN0/YRl0MhMi1W4nhrrUqgfrHX2E
Jb2fzw4CJhP+mIUE2aR5fTwg+fX4shm82LxBuHJUkuGRm2x5A82W44/Lfzp7qLzh
4yzv+6YPHXf6wXVXx23FrTK31nXbMjZJhlTZNsAUxt0QD+qTBilAfiPPyEq3NOmn
YTxyxDnluim3X8IAC97Vn+bGBtv+u+Y0iVyXWcmzAZdz2sFE+pBmlF0Qv2Th/hhB
8D7bO1SBP8VkvZTkIFlHmvF3bwX4X7IusIVXFlaZoUJObWEEe7VC7zqVLkE9sHUC
AcfArZ3XB77YxRBig7aqGptRgVIMTw5koDKe24+zlmHY+RKDYlk+QQXf00oHSV3D
slakhDDhthzFe+Gopb1ITji+0MpjPZraDZ7djdUHh7hvc1jJ6M2HBSwEUYcL1/Rs
iiJ95kHbt2UVgpkwhyYFcFd9tlt1VJPTyUJn6AsW2Ha4mPZIbIzdF23W8kKMwxLF
JavAtIx/z1oleuiZNSQbcksB/8XaafdZI7ig+/6XBtPrNsmvbCChtXP2IUaXTZNG
VZwnxdP3trCNApS3o2U3IrAU0Tn1ACje1FH3zOn+YmFoY7/1Agy+NkqUwgUMMinP
spLzSWZ9N4yVl5rrczHvOijOWn+Pu2rVd6KDFC72c4G/b4Iw7LSq54xn8R22pMHS
B5jkASZrhoqX6X/pTGnLIZcR8rdKysSxUvd7cWz+SXiBDSlphJgz/uiPJlheDmlG
swJ+HBtco1aBecDEg7kJ/Ww98x07qrJckPDG0cMdd5vgGWf0xQgRfFeO7t8y0oWt
MmyatiGzWdXdK6jNRihGQXepPhJF/QpHWnWLVMPnPWkq/QlczaGH+A92vApsFmlg
FnlXsJjyUKsmiUGyXdjdyZD7O7TJxVvFp2tOggAKB6DLIsZ9uCKejHXd4u5JR+6y
xEXfiUnurnDFfyol4Gux70edOyXmJqYAMAdJXJ8UYgveUNdlHFg1A8nosK+DpEQK
J5Zi60pnojGSz5ZGzPWKrlYaurieSgR66HIDgUaAhor0pkhBcsJ/TJT3fVqy+Zbr
63Nemdt7B1LHYxRjt8WBf4RgD+2cOT7vuTT7bCfbVm6JcSmAjrucbAhWsa0lg8fr
BzmTeI1VaDSIqwTgXgvsX6HoQqjSvRZZh8YsqmrN1gvenY5uX601akRgB9Zn6Zv+
7wxrgQT13pEXBANGJoAKAyFA+LmWk3ALw1zVHWigOM6A06fkEz0IfhtV/gYtvPkr
E5LywPwH9Gz5o2MXxGIQfVni8ym7xKWuxx9spQV3k0nVK+3cAQNH1iaHnVihBOLj
ozbwYd2lqmdm2fZPF++UUfYFESTi/DbiRVbd/PqtpIlDVo4Now7p0GRkE1PAYYx0
FHOmDLr7EbcHNzmnq3Uq05SUj0Twf1pnMgVUouX9kSmXK0KyMbm/LkC8WaHu5oay
Yay+I3JxNEx/89apNeK7gY8NTLKcdSLlJhh4uolvkKWl49ZvpMZ+coQfNtFI62Qs
yuEIZgQkqTxwIAdFso2pGSPAwOfgbOPXhrLqOrtvYLfQ0B+K3o3svZXrcexrp0OE
oMSzOpnGewGQ8G4A8n07xgeJoB5zXzZfpfhk3j8Bce1HjbnO2fFzeyqoINTblchQ
CNtfu2Vpndlu0OTLreD+5gQeyLSrj5PHNs6Jheb1vKrXOL5F/AvXNSrjdEW7uyii
Mp6tSYRecaWhmUUtFn8724SUzuVHduFtJEodCMyc3HIg0L2AxEnl/jXBRr2ylZ2+
gk0TyDUdakh5R5OLoLQTbI4e89tKyUZMvANXAxxYMSJwYBwNqrSz3WhOiipmp2Ry
FdGqc4y61fu198YW1R4E2qdAuDFdl8N4awJbsPVsocgJJ1MIzetMC9bGcnMU40pX
OAzQlBmZaeNXlbfzZfpn+FdEJiqFpBPuwT3GvvPYLx1URnW4lZ6IvuGF7nvvO6Ss
7jJdnnGRKFxINyhKQngcbte0Och70K7NCLRlpqPrYDmFxY2KAZaNps+gjVKvUcut
TbHs7+8aWCzGZKv9yxmA5FQ8Q9SGkKvXnHKe2m0sI6jf74R9chs+FtrVeAvPxj7B
InDZsO8mmWj37GvRuBmqtGR0rGHcRcUP/+A6l25S7Z2Mvo47T29mpMmtBsfYb9wA
Mm/K1U6o8bcpF9VcoF9OoyZ9+r+V3RuAOSu6ncoXIJYjqS+YjjcRxHqD8mVX7f41
NIlcrn9Sx+7/xVpSPHmTDF1EUSTrlLA6YBLTMikhj+5SenUcCfnbTgyHaz7Odiu2
aLlgJ5cTf1Lc3hmuzBZIx2x7oEgqsUVsmShtejNH4KiD3VJvQ2wTjHCH4Oa6uc7+
lNBywheOmjW4mpvhlxhcQ85d4LXt2DICvZcWc4JnCDiGuafFANmY5kMdzKJqLYMj
XHu6jTVu06L8kf8MiYe1m6GOcKDmLr/9+trVxDjRbczHhs0pR9A+2FcAboOtEqo2
voIqRgzEe6jJV59EC1iCTtZ9djPldWuFJnoQOvscgXceW//x2NEHBzrHuv9HvPjT
BpAmZkYethgtArDkRy+Tflm8S+As8HEqgLWddW0jjnwsxNU+N1LsiS5PewgDLcwN
j9/L2pQ/Ry3YO0oAB5n0wdTdqYUAJY1iaiFw/CGqNIWuIFPrYKscpj93OxTNFEYC
kAXVC7xUUcRIjFEZ3P2pHtvw9+NXgdaK3h9FoaTfGHJMPwuR15J9N8WfCfhEq1n+
kSk12fy0sTv5JoznE1NefqOnPC6mSrQuv+KfdtUotUJfAlkV38lyI624qs7wS9d5
tIo6LHOME5AeBNVIiEXESRgLQe2ktlJwIi5FxdedfpoijPCHmdAfgPxiFz4V4nl5
e0Ijq8eYQjl7M9A8XkXSB489Bz/NTxiFzNLGOdYCMkKV7YcxrPkGxtjH9DugpghZ
H2AIEgZ14iH6JkTCKDA9dMGfbNpH3FN4DKTiwfrrVbi8SWCwRIevg1qK4+nuzkaU
VKV83hoVCKRqIDktdil7L0sA1VMvFyofnxh0z4Dr6PUgQ7x4GYrIGJ6izhSIMcCb
bmaudwS85QPWBics1VIcs2iq3XhNK4y6qI/0rJ304PIvF7b09s5uaqvUrWRguPUY
ouqX0kgkJQDbqypAw96GTUrhODqQ+F3UVQENlimmo5zz93omrP9YOQMJVpZHxwlX
WWG6r47qgeYrE3sHOE9ta+azGeBPI79qI2MidEwx5x1Uud7OZPxkRTODSdID5Hd4
EDgMN5bdYtQf8DnGpSIRnIl4Jk+OPNJwMvwkZzo5dZKyX6CeEmNsL3p65j7Z1f9B
AgXzegQRJPHDYYP8LTOV4480rWxqX7duFmshj/zIXXa/ah0yScZNjG30DbiywIbn
RCrHpclSwzEhvLNLFmKNlP8COWhV15ql3SpYWOX4aETWYIjw2e2oSYZj8Wx01Dm3
H9LZK99ctTlZC5huBharZuPMalrgJjAhHZENNW9OE+2Dfnkf9LAMWs6O6SECFEKc
B0V5DyPCFTzrhg9Nl4Br+UYaLUzhcZ4s5Wgg+cEZ3ZJ+uYyVCXEuB1dC15MP7hp5
xrt/6CQ0ks7+EnT1knxfg7+63+dDCLJGxVY5xeR22M8BqVs2Ijh1VLBTTxB7q8wp
nBtE6qeYlqPprh1sim+VJY8CA+d3P2flFbyQc1oYppolEbu2RohOC5Y0RtrbkFe4
NPM79QpAWWG0PFZ3kvMfIjXlK+DX2r6mxigXQY+XoT2BSi6lVdhPcNJ42vPDl3WU
wRFl2R5gLlfqwk1uY0E6vdelSkX+5WuGXKiu73qDl0tDsdN7PsfaTUNuvjvaYakL
5HiUCBjiTVAF+VUc/DUZWMSi/nLPuBYLbkoQ477iKK0hXON1FEPCTLKnxf2ndpvn
ZGgz9LSyvMFLVH7n6ITwzx7UuLc1uIR82WgXDbmnWEocEr83Olyd2uNf7pyNlQ46
5gdiPi3uZ4LK7Ndv3g/WGeGXfPeu3968V/CzYLTmpv2K2Ju57+8841Cv79F2TGXI
uG0OSMRy3q7LwwDbiP68MTJKdDdk7L1Jw95CEAyaX+IcRMUltHfGDyqisHqcV5FY
Xv/Ir80EKdxKlPb8m0ymg++wh1XlY6v20DVF2St/0BGNTCx86jNF6ixDhoedftjX
mYIDkQfiuHkycDY/y/gU43X6/eYXa+wg66hjrFZ2cQ3FZgPRVC1D3Th8Gyl0yaOP
r5UQn3ud9+XQqlZzWCQpJzeqj/rNY5hXBm+eJJ+CzMM7ucS5jtO/dyA2pEUzYc7i
UUuLS75eLtZE4v7uC4TAKTn1ykOpAiPzk1949R3uWekhW7zZYWTbxRFdXypJBs7O
EHSwOsV4YQUVmweuKlpVt064q3MbUnUTzHgbKp/BfoN/ULS13RuwsQyy+9gTBf9s
grL4Z1ghdztkPrXB/k1W0wi+dA9W09vmIi8BonBMaIR8HoOv4E2JlPpoVwHeSEQJ
QqbszfQ4qAM+sarvW8fXPWLvaoEM81kqGDto96sAD7EFySvX8xjwYVkFZpVbfMKE
sgn4fK02FP9TMBC7gSpZdqbfFjPPTUs7eFwTpCFS49xqL7hdXkFwH+CV9mk2My59
SI9uVA41kK0xijmv8F4E5B6IgOi8NXTwqDdhIDQ5Q/EiAjFgqVIVIMrbBcPUtVUC
XUrjs7caSagjw0BAkCiGy9UifiGBV/yoqiqNNAnTPAB7+6aoa4AnOUSR9CPfc6aL
JYGaw7Up8M0Gt9nAfURn7ASHF7a8dZurtOW2BMiI+oO7jDXTxFCh6gSw8+iOt9UO
PUhtRz+jATv/yLQfvYon7j2H8oFxwbA2rQKaNt1SBZ7+lmJsOejO1ENY1iSpe4I8
chUMP0pC4YTKOZsuhQdGTc7kM6wXExUjnv12K8PCWWX5g75lA61JIXE0Zo4hCHsn
9Gij8QUzoNALz+aDP50IBWQtxTbyyw+hpgTf+GRqc3IZ4dU01SZAv9ClOcgMR3p4
b1kgMYEnowhCakSNasbRpmMgiHDZYQHPnlbk2BYHj5oI9bAzKAYix45RBQ+3Bm2K
qDoUWljyhYuJjhbikTBYpWqaePkG8Sk7Mznd3/DaXe0MUenJcdmAV2F5Uu9mKgTA
liT9Wv2G5/0l2g6YTgl+2aPwSQjuL1EXWnVpu3RI9wVYMHbkvhFZXxzWwUwbwNbk
BOhe33sYcU+2OW2sSXzc4ppUHtk5v2R2dYe8g3ExwimgKIPoaMeCp78uglaxCB5X
ZV3hWfK5e7yKXmVpy/0Jt2oGZRZSRASS/Ujpgvt/194tXH2ASWnB2NdgTOaD+Wn4
5OgfvtbUUHHZG3XpZao9QGbUSzmzii+kiF+sNlmW++PmVBORxfAsNotvI9GohThV
NT3FcBoo+OQmuJ6SCeKNK4sBCyddbp+O0dWsOCr3Ut9bInwRK5n2IdFz+RzncAh6
1QUBTgq3ObP37T+z/hnmIZKzUp12iw9NVf72GoT0ttTZDNq+3pku2RQssoRLTe5Q
vDA9GZ1c9/CVKf/g6Ik2HQMdtG4rSHXLEsOnwYHbTYd7Mc3KKlNFl0Gw/GiCCZx7
MAMrEGsv3+DE8PIw39RKJliMZJugFw88DZcfOmOMO9Qm+AAPvD5Nof52GQQ7YKfA
NqwusrWla+v8YGsrYMqJ9ZyVCdSUsg/4RKvwqey1eXOaHvYhotH0BNmuHpvqL0EK
5GzDlCiLkzo0p06ZM+dH0goBDDCgiPbjZB8fw8GPS4pvGUGa9jBAhyYbPRk95JIk
W2boE4Lcp0WhnIzcDGv/wwBA7UoITzPeX74yPh3uVX4ksnPOW8zqFLneop8iNSmv
xcRUabppk6Nh3CAMmJZr+up9MCWVK1lEBbebUBO4DEQdX1KfKHRdVW8uJh1nUcww
iQOu4pKlZ1DPRIJtLMdLawV4Ap28B5VJ93zr8v4M95kKFpdNCAjpPBLgOLamF8AP
N4qqLw5nROYwikw8k1mO++Xdgzrkn+SWqwfj8S4D4SmEAB81z/ZHD0VskJV7LqLw
f9b76d0YvFOAW/w8CVHn6ox2h6zbQVQnG7gL12z1Tn7WiV7VJ5yeeHQJYfaw/590
aAnwAsCWOUf9fuBa4q4U2w0HHaGiLY1dcp5XXUR32duuhBGJLGL6Zj2AxT7xtnmy
3+vR9oM+mm8hz+CfAjntRsos9DsP0N6XRIkQInYBk73u0aCMNziFeXpr2MB9EE0g
ErjSt95SGJmTDRJaT/v2gD52Mwlu1Bn8Kt9jDnSlnrHzWoqeJZFb+njM5wTZyQ2P
tzAgfOzZDsB064+R8SG+vV/hfYkJzO+Nf6jFr6YQxn5tWJdi5X/hpfoeOjWl3bCs
vHgYHgNBqnOmXWd7VEtsnJVC490WnB37AvZ7r7pZbJ8bc7DVoNaDGkzCkDUhbu8W
gGApc1P9Tzyf0b6owKTzxzvAQhlDaPiemwrFlm3Ol4CxgGgjYE1oAgoMQYNnYpJK
C6mf+p0VP3+7R4drhGxrAli1PpgA+OAKuAEJzosb+vDtu+zIlTwCTeWTZGke/K5D
ZIOxdtt7SUP1mzO3RRAQ1dEMRAWfkioEqMOna7dDNXjbRVgRGlHvP88ahlNt/854
ldNb7h7Cvjm7JU/efEOpkXmMI5iNjgyUx5G7YilB50v7SmC41+iSj0Li+hLH4X2N
3hAcxW+5csqQFavah0Wpq28lEJrRLBsqY9YEzbfMiNJpw19yJDJfoVHH0LP8t240
WIQ01DDOJzsUxVvlXew8eZNw04DwAUxS0vHN+OS9GEHCjrqhV6hUBdsZ0edbKa95
vpJJNOlT1RSHJJwmhXMwg7rWtNw6qBXset2uEQo7pOYupLAx0SxbtN6uoT8gCZ1v
aT6iFjwY4j5FGzb+OGE1iL/1Vplf3N5+IxSTSswyYRYaOgD6vZrM/WOfXRa8Csn2
XB2ZpA2oDlUE5e0Nul2Gql3Jpr4w70PNFzaV+dxrK1WTvKeAbkDzg8xuzzSYzedD
HwxcRvmdo1/ZWzAfybdDw1X7pC8+iF0DZqjp539dqP0TXzSv+hmneAp9/7/BSpGb
JRQqvfw5mRVjaCDr6q4PaA7v1So8eBUdt17C1ty3LmRh+Lw9xGnpKD3D149SzuXD
FSE6lr/OlQEac1W2HnGFsM3jstiYeM8pNkPTTGXVvm99FIW7Nxg1014+r3vJ9Bs1
6YYWmrDoKEkZRFlDP+XBcwiGezV8dfvKr7mU2JV2K4q20zZIVoh33LzxFz7fnTqG
MSRLcff7UpktuG7iEZ/22olsciHWzrBQ2c2g11sWp5ONHJ4u/WFczp0DHgN8WaQi
xA+Yd0MB5yfHzI5a6e8UeXNMogfKrqBOHb1pXeoDcRVsQriUUtT+kCagpmnsbRaO
Uvc3r5PN/20V1QrfIhU8e+g3wdkJZKnmcy74Yq8IFAEgP8a/c+V+YiQDHzlIotAV
6zYFC4okpSU8Gr692Ax31B8mW5mab/sXAQI7ZFdEmepNugxuy/FAJCpJa3JDjjGE
gqrkMaYXDLfYLXxyzcNsr5VTwxSwYosfmwuZ09vaBGWdr7P0zAfFC1K9c4ZfootQ
YSIhRJ0jT8+3/VmnmMEZtbmDldzdKdBMZSs9qzOBbkTE88WQz4FVMcLCg4mVVTm9
qiqDIM6U7wbOPzjvL3hNpBBAxwONX7w8FIZ35q78hIZ+zgLYOsEzap6A3SsjoCUe
Cef7ToxpCdkLCCdhuaHng3E4j8VwIdi3n3aLE4mMMNehbz3INrhmCeItxxbOgB4X
5PwMtWawO/QURqtcNDjyixGtdGeh5AAHE6N6+b7nVGtL6EjGKOVKQa2OAuJoDzak
XXwIdBW0VEaJcTP7+ag3FrhfDUVafZuSUJ470Gc+R2Zv5/tGU6vuGf1806B2/9or
t7JijOETNZDR9vo4oJ7aYbr7xslVhorfEUFtPjZqYHvpE3e0+3Ko2QQxv4ErFK6m
uggFA6CoC6CJWqdHk+sazPBr576U4Namy64QfpxjAybSpZKfm4Q4ek38mYAQLbVk
v6oiUNbxVx/rjmbYjisVWxj+nGMWRZ8MYzBHgmEYRnqt9FyZgZdlAODyJkwe7yzy
OKHuaOBS+dpqZa668PIPL3VFGFm6H6ENtfzxyoiLKFKDZ202xzhUm8fK/3sPbwZa
DsG3CheQaB3EygAr3mV/6+O9EgRsNo0xaKqPkCZ2lIokSAnzJAuNIFs8E5ySSbp4
VZiyJlRTVJaBOqI5iddzg4My4icVg3kocEJFc91r4zO3wvk4Qob3+UD5G+8tJSAH
+HZ8MDX5q0ay3424z07+DC866MGTWjL7BTowWCeR+LQ/cWuPcASVyLlAnteQipPu
4lbqQax480E/B/suXuUvU4PuR6T6Np9EIMs5vdtN1OLxoBzUwsvl0Sy5fwuygX66
2Y9Gl+jOxLk5d78kSNI7CW34QJACEH+oL3yQGbPw1Yu5dI01kPQU57TkiWWX8iP/
ai2qm1/tFUztYAaXzyy3YMQ7oZ6qNW1aYt4lsYV7bT8CBENle7nBETY+WRcmaEJc
bM5rV+Tffe7Htm4pLUUV5T/y6xOpnrLS/an7M+bKYeQ9fq1FpNPVfV0UkFfhzqVb
nuDqq3BN55RO2mDV4hWZyn77+7OJ/MEkvD8WWkDMLsqlvv120Wnm4FIJOb4272Of
7P3ebUFvVjwp3mBEKmaPPsI0wXfnBioG8A7GHset9nIPNyTm0jGpcGc0I5aqjpfp
DuSEh+PwwEuof/3FGZCpowKHW3hINUH3rz9cftmDsj3+egiRGMJGgnEUUs3kv2QL
afMl6lxJsZ4BWOhG8Ut8PLnReFKLX9VyyE5y2T96iwkOLFIFD7pAXrJRINWCFD/s
mXpoUcqVYKp1Mr/sYL7/t1cAoXpm39dCfgRmgEJkpirvVQucZn8KiPtn4LPdHF8L
kcNe2vUPzB2o7jQwvKfLx/Srau9oW+SJqbUItyd1kkX0V1z2ZOdTjkRSBUdhiYnH
jQKSglVZEtbfNYpOQAbXvmX9hGDq7nU1L9tnFWhrZsgLi7KB+Zesq4+iJld07Cne
4EcR9Q0S0HncnzafFMWV8eP1ZuG9eAotpm6dGyCTiAIbC7m19oIT6ZZF8u1iJ87K
BbLPO3X6K4aEdZCxoME1ZB5L7JQpbolBWBAbev6A8+Qm/VOwmrjAi2Yiw0ra58Jd
ixfVQMxlOSXH1jXTc+OaiYmEvVPaHTrNM+GdIoVDmSxcYiuE6wfqAOSCKgF0z2MM
/dKusR/N/nnPMSYU6BzNn8ZBI64YcMcKqMZoyi5vHr2ORhD7IoOlbpsTFleHyx3W
8bGNbXt4gORUcy07no7shVLQzLYSx+DqRGJhMWG/EPSRnpQivlFxQv+bLNK8wtd6
MYNTEcWufz1z9fwXFHaUcXwkLx6HDCnAp5T6TLYqebjg6VE7k+5X3pRqq4+/mVeQ
7iWoHXQZK+C6Dc0Tekm7KgXgFCxuL8gowvmymAO3+vR+aw3zPLUw3L2ob/BKs4J/
dQKnsYmgbfgskSK993sd24GdfUm/js6Jvb5w6Xq6p2CV6ZBVC7p3m4yvEOkoVlWu
gFReRkYhpfiQvmKqbyfHmMv44fZqXYheEAZutXBHUoF54w++ho1VjjBcj6SkZDwA
uHQCEWluW9QlNduVevy3iCFRpH7AS/6v3xzoYwlZHUBYtbOOvKwqJ7axmFjOGT52
onn38BjX11qjleB8nRcqUH2iRhD//Up4jX5r95BUDYBa4rj4hkiYEtsE9vsP11iS
4Qj0cVY3nFIPwz/5++JSe7C5Mx3M5onGUki9KvxD8khswhsydkugG9fjHhokZKMZ
NTYW+RbXhrEQfmS+sk6AT/+bRMvDV8VDShpa46Rb/guBXosMasmzJzk4rsEHVI+6
Pb2ZZZN8EcfLVLcWHCzL+RLkx6vmPUeImyPpBrE3zAiB64Jf8HfpeJ4rLu5NXHpV
iV709zSSn++b00lzo5mPA5dARHYnV5N1BYmS0gTExSxZbAjMjvvJO3a+AGQyFMIL
J3DRcSiuN99lp8M7GGbLC8y1hRo/cCtNoD6Udi0BIlF2f/ewhlGr0+dDP2uXCv0q
3p+HjiHwN1zxFC0bhIzGZeuhKWQAJTsa7s5vUnsKdKCgSNgXVlTy7FkcgYDw6rro
LLDCs+8yIGKRUVaKzVmL1kebAsgfxdMEjP+h6LsHhSlFf0deeXLsG1c9qb13Sk6k
nlMnmh1ROD/YQRRK/48XQOdMyDGSESOCT+E1mMPYv8iTihaH0l95KnB9/s0w26o2
vCUEJcrOtVFGJyifYX7ymLJMn8eX3WhrUqvmyI2t3pojJNQ3rKPYUMBF/hygiQwC
8pbHj9CbAapkDPbya1ZAUGiKci+86OO8ZGxtWL5WFMrfuAFH/b5xQb6by5nYkphP
BNHlagXVC4vfxaqE1nIXxGFJZ7pRQBf8SmqzOZy5z64+raQ+dk7cmc31Fr5U9/w3
hplsk9eaPMsiENcvFPJ2vYWWtr9CibdtSrw9EQ6AN8GOpiwtvLbp/CcvccHTPwbE
vVn853zyql2aPuVZ2ZiqMR94kTKYUNPxFcGoZUiiwOpNbev3+XXsSLl+n18sZ0La
IIzISfeHmOZARKpMfHOtzj/VHFrEPva+yYUHRiYSzaqXCQ/+kaRedQeLcKg++4pU
AbmCTPc+Wj3ieryxfXGwJ9s+K7pdUfhRkzK5Vynr7MWNDV8F3+StY5V815/HFxE8
rRqInlrpCEIBv/kpf8pNC1jbLxqTI8x44isUoeBaqUHLFWBTGxRQYivCrqSV9L/R
Z3gACfRdf7Gvu5hvtFh1pl/+qZlG5hvKaqxmEa2ESwD5w/sFo4AjB+2IFTqcOHMn
BSsG35FUEt00HWfCC0dEzsLREb3QgjdDm4xNyVqHopPHw96c4vZrnVRCShVoTXnS
0VJhPAM1rgw9KetJvfE51J2wg8q37lPFSHIOnx5H1I0eNCIGLHpL24du2/TXLoaG
qB3RfXsYty7oGmaCo5ICoIu9G5Rd87pfeTjig2i/phhHIpsnX5welfW6ZgMwOluG
gFfnJldENmXEDJ+0BxuNLykgWFF9zPcs09a5FMIDaQrsKuM6aUpvkOkeklrJRk6j
7l/+yIHtthlxl9xLo/TmtVN77Rsye8IZbpZo0iUBQ5HX5oEdS0KpZ5H1JePaXyWR
p8as3c0Ws88kQ7S7PhAxwIfJpxiIBoCrDY2CE5LbcHy2USnMDwIs4JLjwLS6tL+s
edvLbeTdG+ulT+ba1xXiCT+sD0920e5hYE3GDWipCKkz5dfQJ0tb2ULEVnOQx5df
8NAJHWxbg5g6Pldq/C7PlVKaocRhXOOyxf9Movngo9A=
`protect END_PROTECTED
