`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N9hovZ5AxqeVtY+mVOR94bTcHye1LGXo85oOVx6ieL1lGIQwuJoRYmox2Rnsl5Ux
9sqU0k6PHFpDCnCOsvuuL9Wz2379FB4qR1ACAlMoNXaMCWytMjVhMOdfcqUT1qgK
KdeqMqJ2gUFD43t/lK/EATchojugQo43+BVgfrejr1jW9HfVGI9lfIfWcEMfvkDX
uk7FYDY4RHMq+ymxjMat5hPakAh/23W3gqpeQWHaxmMTtV7BL6OeVMb+OmR2ueJl
CVmf4K35nm5ylgIh9+GaL1zxZLhITG/gS6kO/IOTZeiyCq+Pfn5puOfqthXg5o6J
WpgcVYQZqlJ0Hq7ggm9V13CZR34h37WWoTMc1BTbE7uSCHfQtvoIXvDhaogitMm9
5wVCcAPoOj0tSq9EA/p90y9Pr25hA1lKUnn2G10o4Wiywo5ewmA34Oo10voOwfqT
xgz8SmYKiEA5bSBuAUpW0MVaWK/lIMQJvoGEQxNNSRz3Xe+ONmq8dlEshVZfw5LG
Wc3GG4NmJKIug94vynlcEFV3pNa17qaapm3pPWxmmLm/6abioCqZSnROLqO3h3wn
ybMlqizc+6f4Qv92Mq14Wo7CTftYITYuuhKPOPhcczhwglYdDZgLXg9D95OlTCpi
Als2QsV1kkZ4v2sxPeaBJSbXw+7xVxbO1itMyLP26mITbRomGluF3XSjG+PdfOkN
SuryfpQpMbblonAgcGKHSK1jv3M8FD26/o5NWft4N7HRWIaAl4I/e95S6OMxHyRS
Fhzvu1mKjoTGroi1/0xs59feArYtOwoD9Bf9EuhKVFBHKB0AUP6kzcdUNabvzESm
IWPkL8uNDw5GC1aEEe4VV6ZS1/8CsZVMvu1o5yrIEbtghz0mLyP+NPLhxxlNUhJi
REGho3fwPWKatL4YJlmmMzLF4Z7XIWqqDlSvPrX+jskYdNTlT+vurEJczeeKZoDZ
veWepKTQyDSOGBdxUZPwLB7vhkjyFmLqh76p9eZ+WdqxCW0m41Ukmj43nfW87h9H
a8q/jCSTMCx+TBLi0nmFOlI24Rr9h02XEh+bxOZBb9qyMa+zoM8D4o74cMkN0+di
VbydJmD2Nlr93rE7uWmL4ZHEUDJ7ysLWEN0OpqMrxtdAbjsH0PDsucGpFijk6h6Z
X69dkrCCN7wMA/4nP3mV7Cl1aPj2KuoIGZka7s8Xq/ZzBUzdHIPWfZ3N++QiREST
qSFE5sGUjPI4+KSJoYLHxjJnbgaA4HFZojFA7CEcMAEccHp7AycmeXtZCX2Ey9+i
U8s4Fphh/d3WPeOFkUQfP/BtFx6MHd1FNu/ZJ6ZVGuiysVx+8CIgBOZf6MfPUU0v
gS/R0IkHrGLrWAhZmJmQa5JK1W000k2wWub30rpWXQUXvZ0MJQR8me4S6h4rGBmV
WrzT/NMlWOufBrzJEFHNypEcr2AsMsTEqzSFmy3LIgCI/MCiTm+isYNEjjQ36Zd6
KiR4G162Mg2hPLNeWn5ogd+cZbv3Mthh+coXLgPUZaDiycYmRJsHwSV2bqkO+CY6
SOiWVof8GZUG3uFm19Z66jaL26rQ2MHv3gttzuF+GaViFIBjsPphezw18gsFhmH1
Pc0VtLKaZpPmenM2DhxBXdHBy50I1OjvE+SKeJ0i//a3IuuEEmy7GDrObMYG5VWg
k0nXKpt9KGyladoABU9sy2xjTKf8ENqlk7fASOsHD6WQXqCD9CtjsUq0moGuWiWG
Moh1t41PR05EHybowpojuxrwv0LkehIeoFWuKMZzorMCHcj/ss8S1b4+vr2/Svgc
LDVRAFWvj60TOyscBlPVMsQ5ce3hafmGH9IDG6Cpz0ORPW1fAu5e4tm/XVJLrHbJ
qiUhxnRThJ1kBcQPZswG3/jxrJx6ggq5iLc+RB+a7Q6BJA5Nmcs2ofGidD4KEqz3
XlWIZIUku28a/YjU4EjRAtAGwbcivthQ/b2loavmIMzAEudysWsNl7TtTy7O73e6
RHsAVXV7R7r/ORFATrbYd/DSHBSAgXpk4iytwZcqQDOcaoZx9Y7m6E/0qOKBSIs1
`protect END_PROTECTED
