`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NAF+KftEdXxIyrE7Haa0aBKy5MxOArEoBF5PjbIpGiP28YPQK3koMwNak7d6N+D9
OcvhQb5bjKB27+CzT/EpWvRI0zzRZB+vGUlaW3SrezSh1qQQ/3KlUEetVYGRuFJ1
S/890N/TXWkkiPBhKOpeTCH+Jvcn5YYT+99Xzl6wQbN9fl0UitNfDas9YLxVqyRe
k3H5IrLaTEa5/fP+frZY42Y11unL/4ZHm3B/zJl5sBeXT1tODXfcVw7Ggrjuuo0X
CA1LDz6zMx6GB10XOyP3qYcmFLVR4D452UQ8dVPoplqcKrhuPi+ImRY5M0O37HEh
QAUL84vq6wSXzTxl7HB3PlyzKLIMoUz7XuKPp8hp+dK4aOjL4DJA978dGd1YUotK
OzpMDt0mESMI3HF2yFyGROA3hPjUA2s0zjq2YkseNxjGMk+V1h0i/yw+ytVea7Z9
UDH+8daq3OmFNnzX3ZIgB4ArVBFASA7r7vupwAdE5t8NIj1AXbn430ZoNacHRJH7
kfR0V6QAXNKa0DpZJygjkA==
`protect END_PROTECTED
