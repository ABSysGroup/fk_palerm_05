`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c6IKfSvE7b/0aXHq2zh26Mk+tC4E3XUbeAv0lSRzFiZ5PHbNSnEiQCH3XV69JmAj
c+j2UkYnEwz13r6S8zTBF8lP7Vgu7MbfvQgbuoetXbeRmEFCsgNgujDiaz/IBDor
tyhKf0Lgwf2p/X10/9CTNTQI8GmvqSSbNwNj5V87HPrE9aXKAAn0f/V582bwoYRc
KNoEOTCRiz5uxsa0EL2GcvOhJIpdS1SH33t6MON4nrLcZmIk8cGDzdOwXFEILpKQ
hz84tmApg6pj2OjzNoaCafr7QqX8yzpzkreBMd+beAER4lyo/u+BL5zXbVzFv2+w
E3E91RnLTeod/aDQYXcz7snnM6UYBAEoIx6gthI1kaBduN9huy7iz5nlbdnHcomd
dzIdI8PeohjU0wKkRQSdGNWXomja+q1YQm3Zri0mHzZpUWthXDYZ8XeqyetnE3rk
0GrGU34QHT5ucd4EIN8pXUk6kNEuXLdnIIC1GPu0k8Q=
`protect END_PROTECTED
