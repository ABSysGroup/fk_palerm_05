`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f92gaOHc1MUO8qYpJAgyV+xxIleee9wc+yzEDsSCUUToZD2nnnHSJZA/QM3JJRTI
plzNQPYIF+dDKrVIVopHKfvxJ4y54HUfdN6CYBuUT3ZJuHThnzjKDygSWc3UuZI/
PdEUZH9Ht3mEsCTAcj4LQh4oOE18IVZvFQFcQGc7FHKiCkZ0LxWb9WSue7PFnzTu
L07gpVvFnJ/tVRW0uvWkSZYgWw+gXzgcDgZuN1RhjS9idkyZZkud/t5ssi1+nqPa
EOhkJ6AAeVTsNr6K5MnhSywHEqAcxxJhA79YiEnxQz5SEAhwUwGnNMUtQ9qptIu8
IykwDhvNYdviIc9a1+/U9AlFbbn/q4S0CHwBFnWvsMTFbHB9hDG4hkPWPj4ocjCf
SOWsLKm41znXK6ue/hf1k98jw3oSHb1+KzEZem1AJHvJn3Anbox3TIu6pgEMr7M/
tjj27BV6MUjMvyFH7747lyt5pCygY0DUO0SdOLPUETM=
`protect END_PROTECTED
