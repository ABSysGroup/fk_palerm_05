`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SKQqDzkVJJiS0Wst8OWapP1mdqIPACC5+xmsW8g+zB2ouvOa6+bLX5BDywmJ9JS2
WVhABoZ0AQiWcesO1ZHaTJtPJqaoni57lLbeblkgUe7/AgrOQHsfZUf99auVWYMc
LRigD7vkOL8kgOfaDJ6twBRJvkkZOsXa3Ve6umIz/2hzM+yW/ipms5edtR0gKER0
gcjLFraqxId8ucjT9wVLR9T7/MuszToIiEpJxmWgMRrpidZvGf1rfKzgHXG1wuuv
NVfwn/XMeyBHtAjxXtUbEglpW2pBThZJo72EszeDUSw=
`protect END_PROTECTED
