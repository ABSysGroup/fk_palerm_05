`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qW2spVg1olCHEcq4ACNO/VK1B+rRZ+B0sBZFAY+/XwpDHJWBoZuyDLGZBtpBgxkK
WTRTqdr3ntaq1d/vl0ejjzKzKTut2VB70b7R2cWNEn+Co2GkX1SWX8wcixYJMxkn
MUaHyN9m6rYHyDPm9BTUlCoq1w9u0nK2Od7/eJQyzSNr7jHtF8daGmoO9otCRPTo
jRXDdfht5fKNB/kHO6AuaQSfx5SNtkz90R92gaJYYqkF/SE91+0tzFSErDMJSmoO
hCQhcE2C8bhckOXPY4gsT/ET6ITRYrnHqABbqcq5ivNfpqXGceOE4ySfsjTrz0Mj
PmUL9ZEeClVDBlmBiT4VoPkDahDee7BCcPPbM8assAxlC36N57Rl1hv7MdFkvD+f
NJQHNu0fgtUUKdEVaSRllCH6W4X6MpEM7zQlSVZFr0MHnRXd7CbkYGvIJOF6mV5N
pXjDcn8YWnb0v3yzosC0baXNS310uT4sISrMhXMGaYDGsLzjqU2SIHo0PCprWPRf
fBvdIorfUnvxVbMPjOZ9Mp9f+TfC6Ooho6xz0oEhY7mVK0GmTJ3+l1+TYfAS4yAR
YzE/HMZMKy7kBUqbrqr47D6TzslgzBPQOU9KixMv6Sbwzj5RHfa/kMWuXMiQuahF
7H8AMsQvDXhSN0OA/Ts5tyAtj+ZJi3UJI4Acj4FLGiCljD2aETIqF0rGJ4WWlZnt
jDLk4Z02dkLXBq5K+RNtvLhgbgEaDmTdHww+5QGemeLk8jthG2GnAbNkS/igXGW1
LWwE68P6n3Rqk6MJFvoNTurIZhST/SZQnBzYD8Qx1mKzOEF8x2gkQPSJSE2qKiuH
k0v/fTyArZIxPT1fKhm8smntjw9P6xrpOOpM4jd14POQ0CpkQfYaPT0mM+ux/FYx
h1rJ2PdGstPXQJH3biAJqQQZluwlzR31WZS2EPz4rZTcIlgqg+cTZRvN2F/BbdMs
fJtKKjJYl+zYyCcCTYKp0AM7IOB1VqdeU4mqNxhj5kCMY8lhF/3TGejoXNTcQ3DP
tAKct1RnS+B9IItAP36IrQ9x63YXdooWyIjdqCX54MgZen0AY2JQBqKMA7wznD4a
TADLATV8zRTBPHryz8/V6biq1dalH1Eh90sDZLsV9HmhysHfSUhocZf21hTzH7Ws
zhsUqOlfbwdffy5XCOTKPMb9DBeGftbvzkFEqQZCeI/0o7iDyLkelpDJIm9OPesQ
1IUscOivnow74S/WRNG/gsb4FtfhHKHNaIdjod5ZqCe3EfkdHzqWYnoRCJUbuoIs
nj1jP+Ofz/efbCNAHPNv5C+psgisjVeiTCHMN9niT9OkRxGw4+we+IDxFXxvJddw
SBspkhORpx4LjmLFGaf37lVB0rTSI3ED1HjH6spWA46UUxXB2HkMvBlbGtCMahdN
9s0TfDm79u0chJDKXPH+Dhgh3spnwd57oeRudXYf6J5OIk05ssu4omfF98QvIeBp
P7C8dsY/ZYUp7Jsv+d/q0iFtb2FImHxMZi4FSS58Udwo2CvQ3dgE3qjyYyNUqjId
6iciTQrtwL3vD7g3pZt2V2Fi+K5f3U4uoZ/9mXwSpG22XHEoerNpBNbDJ7YQMygh
`protect END_PROTECTED
