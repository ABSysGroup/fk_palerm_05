`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rtnr8Eh9bP2r3QP+tiYqzHqyLpvxMZBiQtJT593v+HaYs9A8iBz5tsGIdL8wqzoj
M4eMmT3tbBVSUOPWJeoX7VahRR6gjt/khypiPAoXFEZW78OsFnGgyY7ZTjkP1Cno
IREPuXcxZLTAXbEfDaHBqtDalLyNclXc96NjqyPs2YMMKPFVuyhn3MSNL75Bz0pp
9qHZJfP6J1EqeSx2BIeXN855rNXO8FWqkMdy5gK/hZo8Wlu79bUyjI7yOllOqJjg
yITH7WDZ0WGKuysAnOJQ/H0K7oDlnnGQzKZs+K5qVLFFjw8ITAg48bK8N6RpO8sa
BMvV8kusC5WvNVUNoM3OzmDB9t0Mn15nIsU9OarUvBXG5cdSLikN4ztRQfblB33b
x6nxyi3Lu5aP4HR+OzUeUg==
`protect END_PROTECTED
