`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nyMr2dfZL0/4l9Xl9G6Q8pPLZz9pz58e8LlR7Cx4KtHjmjPUZnzsZdC73dHbDkq5
nGKE2dOcIiIK+XD64j1kdbFaTNJp62bv+WD30TDeCzKw5NlBNimp45leVhAzowUK
63ShNNzHVWOQ+tqWt2AEeEAUCOGrZongUgaHav2xKfOkT5e4/bgkLTA54F/B5n0V
8/9rG71L+WdkyE6r2rguMZbCUzA1jbCcNDq3hPIoVhGrxnyzXCoWhgnmm2E7UjlE
p66IQQY9iRoVVNNW93oC4oHMx+7KMgdbtTyz2dUCsLvaeXThao7pGKS9TnGk2/t1
RQwhvsxMkvXUKmGhRKdDtIYcD8gcdqVqgt7Poqu6H9R5FbWnp52MPgNeJimVi/QH
frmTYevMK+IW8ftuP/HlwmXqEfifeHJNZIU9XpFPdcFIIc9egOw54wESvhLD9Pqt
64vGdLYyLbWEABEp3cSy4g==
`protect END_PROTECTED
