`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j96Si+Ui5vf03IPyJHmkKAQ4r0aokArFePIBZOLRIj0VDBaO9ADf5DVQMhemX0FL
iD61Kby5DCARW4avs9qcv9JQt6PCjqeCJYKhhH2+CElhMrNEx1gPRaFB4oka8u+i
2EowkszCPwgumLdRHRcIzGMynso55PijQoU/R6kdx9dn5Uj05ik1IwtWCm8tdugG
30Jh6ZvBsa/VpESv+IqeHBQAoxyrFkqbkSo85Sqrt9+uJSWBl80HbmMUgiELOL2P
24INtAwomdH8CNkTEGNwUoVOaWamOHYwJz/shbimxsn9oS5JLB5+sMasKxpWMUby
RU82CSKLpu/lCJ44UfryvfZcI4hhuRmu1U0ym2YEr8fx52ObG3MJ6J4y/JRvYNAH
RuCHyJjT8MogDQlYndSCc8X1dMJ5EiVbHEkp9W/QU3B8bs1h8i0n7qWDwa6MYF7M
W3E72pZeS1IV1xL9jyEqtvObNN7jHYrhXURoc4DUvx8PfM7hHu0bnsLUeQko6h+r
PJdPG3xkfL6v/ItT0clAY5S0JX9GMI2/u1izJRsEQnFDkGTiIgOzpt9fJ1sUFHXT
OpkUTWfE19GBIA8nnF1kZUkKJvB+38oNh/kOteFU11JJwJnp+ABvRedRMimjW8m3
2SwsoEjlXVWJ2LZwoqDO7iOtFTqEPow3+hc2djcH85NHcdKKFONneyWCbvnLKfyB
2a5zw7huXoD9Bj+ad617MULkwQkFv9Jvx9Fg3iRfJQ4XzwucqjnQv/X50LzN337W
WSGv45VDSb/ljAO06cPURUkTdganaOAMBlfuH/ZoIOU38k0Yscdvnw0RAx5VSFu5
KjP+YQl4r9d4PIAZ41HqiW1ATxQbyzEZLtd5E7Vpp+CRdjX85b9BudbmXuklEf/W
Wh3vcilNjEFRJVZGwnO1dHio2hrP53Dqgm/48/LLJjOp9v3TBEofhw16m8m1AWZa
8NA7srUcMqAqyEudItLuw47sOLolzbC0soRmVJWBg/TPU4feGb2ZVi4fGUunfGZc
BhY4pmYjUmrIKNxs4xxcnE2wy44dt/Py0XCfSgkeUAnsQXhqddzCsCoHX4FiYU3k
7/w6KJTg59Mcllmnf9T+eGUZYoZ5pStU/4GC4q4gnP7H3B+9iUVyxybxrdtTCdDH
4O9e2QpTc+nxLDynGhH4vrZkz4Hk3qmsZZBVbQ7WHutNoeQP+0VCKcnmg+VQH7tO
W9HjaUdEa62o/RKhcDZvs0GJHFgA2dKEspOwra4Nr9IBgKThssW3c24nBNlk41iE
Ce84y7PFIQVQQzhyEB82tU/iCVyggdyVW8pJnD8mqfrIDCB+x3h/yS7PJPCOAZlf
rCkDN22dTSmPG7j1LSt0wsAc8Uclv482n1cM8hAuF75DBIptyi8V6Vnd71K9ZejI
T66WHvI26TtobE0g+sOBDolH3ZmN9xRt1DI6WlGsTeaS10RRmoH+40WKN21A0RRv
/ZQ3PCWJqYyUk7q2v6XrhuQBhtTeHzKRzae7N2vB6VWlHd+w96/EP+wyjcU4Wb2i
N/NJAsdL9U/22jQVSfF4gKnRsC7FWJEqiKmzEnfmAoegL53zsQQTjq8STHn3T/6f
dPkjaYBr2SPIDmQrEVDohxh4VYYkd4V10HtEHNl62AbemwdrduZ6NvJZ0nm7iYI0
52P7GyXYJcjnDkkRjzo3n7BUcUyvWrGbiB75udn0dUZAeF8+bHdfb+u3gey0toL3
JjT2L46mkZRP6wqoAr/VM7wDTmtQ0BmxQGN3Jl8Sl+iEUOPjJKaGtsqJ5lxlzosz
vY8o2wIUpHuPsw1HsGrDn8+5bhvXxn/+qEWWnAxYKKh7M6RAHVl/SCllMxvzmH4L
S1IbRoQPs9/nx1Bvg/y0cp3IYOXUyulPoU6Vjxm6futkuUER39O48acN2xunOowM
2nFophftrrJVE4XCTjzaBsxhSW9oyjB1huwI0USP+0zJkAyt16qR2+m7yu37726S
sA1uZEqLRekQnFj6sAKMB74ltooXdh/Dv0251Oj0OYxV7AAL8TguHt2FH7k+cFQF
DkdgaVAzCUn7+S5+Q7skVbbsEjTiAwRQ9FJRCYIqdc4khpXTj1Z4PDGSlUXrEExK
5PE6z6fzk/9LuDnpsS0q3GkN+ugyzpVHm26bwpfP/hiQ8I7eW2zbGmZzAUHut7MH
yZwr3bPHaBzemJB+czXUwTLHtZKE/rmo0D+qh7I75aL6eG6cvHf6QGzF2iJ/J9Fe
z78zyoJnhzH+JGDEP4gXOTEoZagOH+NaUN+mo8Oil6K5Mhg1G1rpFf7qmG+j2+0b
kN4q42E7kHAbylyf3wVqsMUkLaWHt5fDeoY6H2oA4DHKcQjfLnlgPKh6GUT/uQ5J
34Gfz3l30cM6/6U+w6DmWz7T1AoUuOpnDN4ejYXgsuwAPzUvjKxOL7h+xdAe9YbB
YIKeQTtK8u6Epeapf7L48TbdLNnVfNvcGjob17yuw3q5cJs4S/xywmNTS3omE8wa
OtefsBpJpNqinm1fB0JfdLSULv9hFKEdau/0dGroHUUw3EYDBgJdlws5MichS+Lw
X2U2TdLeD5b8Lt7KBtZcC6rWcKovZmL672hNggMT9fuXGDz+2QlwZoazds+SH+Ob
kGpXdQ2tZwSGkrSdbfwdNaoBfasE19RoPDRZq9kIErlMff4DDfY3s1iQnVS560Ap
V6yAm71z/fUqDYh6NfvuWky0gkPpWxJ1F3R/HBKweAykVGdgKV+RMYDdQXDt4gze
Nz4LXDtV8YCvncmroy4Gt+lcMB3+DIvV1j6p/LTvJD9vF/YVEoddz4Osf8WerMo2
iTqfsr612WGhyd/efBJz1r8rV281eUwgByq2OfFVFxmc8KDnLUcuwOMhnxaa+SCx
GWpSb/uy6AQVrKPC30NFeNPTQycRn5SVaRZrUorBgLMHLwqlnh3WCDyIMh2Oy+LZ
uM2inYq7u6BwRR2HZl1wzz5rNLTFdZMHNTDeXmk0Cf25/rED7kiPNHp0WxTfDPv1
sEiZuO/8KnfK49VMtx8z1Rocx5bsRS7KmxYPYtR2ZXBbtiLLhLfFMnDfrvM0GBUq
AC8aNJgqCkYtGnfsdZMtOV2wdKrN+m3IbwOgowHHKIDTic1Skx1p71Cv4MRmldSj
JZpZ2l1fV+0KZ2/dLpaprpqlxGak0GI+dohjQExlAu5jaKflVZTJZa50bitCZPjX
RjYh3TJhLo9fG+44FauxQusjs/Hx6lwGAtFcdD4aEpTzIJusCmflnXxVxMXG1K65
aM0nt/xhG8gRqyjLJUd/gzgcIDsmInlb3dXxYfkRlKq0zRtqkwmo6mErFwEy3Zz1
PHsuZcb8FEGrZwZkPsG1jPqc9ITKnEzfjQmtoticogNAn4Dit4YFAjwrIvKH3KxN
2Lzf1a8yf4Brp/EHzPQOgptAlmjgG0bp6WuJNH5PEDab8CixdnEp0b6EKTnVJdIH
FwgR9YvNumtlKnupXBwUam4GAr7AZdi4FeExdMoj5dgJTcUtJVUUiabxfezvQJPg
HrNdtcCPNCpPuYPp6vNwvIzM09Si3LNZPpY8PG4ddgtymkOQpaoMHcw5b5emADuK
4+t1n40wH3Vfq459rqTYV0nhgSCHos3UD8Ez7VfKm/mYk3XKq8VzesgDdwltvZJc
TTwbajisOVPzNUsiGM+GP17MOms3rhcRaJHgGzSKGyIDl18BAr2UbzV6xA+Cz8fn
6JkFDVOKI3tJxjg3kLOdhysJQfk6svs2aOod9cbl866y0Dq5fRIB1Z2M3Ze2CBSR
SbQBH/Wlsr29DppFKLjRoP4zO4VfdzFIEmL6CnGoMcz+u8rZdXkaNIM9yn6DRsER
tMxzDMnWd8K3SwEbGXVO5H3OeFTUdka4dfSqrkR1xf7+4ROTXphmnj/pryOVSyqx
laEuq6+O/qbdcpcginlQ0EE7gZVZUMhg0nQgNo0/M//0cODlz7keZ8cEcp6oT0n8
mfKHKf8Osc0oIVywKR8y9NITXY4ZWIPrFXLbymcYt894J1vh/UcD66CpIlVowPwg
0/ef/I9eZPSJmWrOvJL5jvh+ZTZ27zbTTPrvbIA0Ognz05ZeV1eZKU9kRKPIe9Mg
OKqs39o2AMDG+zgO3t6E98I1FQ4MLWYmzrgpaJqt2+sd+3+u8KLBcxt9naGoK54D
4my9AumY6JP5i/9b5vRAzTjuQSyWz5N64ngjfSpEpJ/Stqw6ImcctCRGfBmUC1TY
TeWJ6+ccOVfzf40QvXWZjCMUslyecJT17iIr0Jns3rJveY8MPRHPZcPbSV5Dmll8
rWo9wd74D/SAZRZrN+w6xm11G2Ajbaw6+PLAD45SSoBaZYktOf29Bp5z5qcVGozc
cPIpq4JSwQVvjsCnWg/1yVCqglBtsNNPdF3MAUbTWNHLh/lD18equYSsb7R5+KZq
FT/WOh8GeVD57XEju0M4LMsmNBC9p0dz5tLD9rpXC+vW34tAlpvzrB9AQAr2nLz/
86j5UwT2bXHQtw9fkNXyzgdW8N8qO+22YFN78QfDaHtARoHcMYcH5WAK1V2LQjiH
HHDkDUwi4HP4TfcGeeA0o1RqPBd47JVG7yCR9E5lel1NsdchXM+fVy01h+d7Nqed
n3UTv+kQRBZfCEJexmWIT773VmfBbUpxVil90XUd8cCiWUt7Q6i5b+SGDPSRctaM
vL6hdRtlWpuXT9c3fr3j0BrOfYKshrIwbIIPRqT6PF8nSaYXnzQsi1x41XpvSFxm
XbRtd864d+Jy7TB/giI/lvtd72VV4E5w/1CGrjOLhRXO8eg/z0N3h+yvdCTgHEda
dEABfqrmQnOE1zgZEba7o0g2GiJlOhOPOyp/EiXmSpiLHbCYJ24sptqHMqv+8xrX
A/0oWsPGnhb2irFy397oK9pAvpUFI7Kjrh8uKT+XOIad2srLEmN5uDfZwHA7XlPA
r18/5rhXBEjrKtYoUWz8AkrzHcqkDIlOFkAn6+0A8YQpPdOnO4vlLz86l4Be8a4N
jmz6AEnnj9UewqQ7vj0n5LLVrbDi6qLqCZ7zVxNavjUYhQKaBcVor/URE8zvmXMS
IYkcpM+z3DSCsFCjhBNFnBp9BYvsoyY7q3VbUbWFaO0TDgg813125KmXTXr+KK9d
2gnb1+NFEY15vgP0OVxmjNrdBHN5NkgJo+p8A5pVB8WrO1jjGNlllYdU2C0JBF8v
T7x6XoT4At3qNydQVthMzmeu/7HsKubVIIZ8abZsXF0Ff5lUH2HlwZoSVg7fTO73
9VjXA+i2hLkfKbFLlTFTdQgDLEH/Fd6MzMZMrttn3iCXX5eFyAaLa3+JJKs3Gbto
QmizdPCAs/C4JRgKe4pF4v25oeCqivWtdVDkUfhuiEw7VBTRD3fyHGvQ7rhxIR7G
+wPODZQWRNKXgU24wRqphJJMntWAsX6wUxbGO6ZN2tQWmBXeKLVmmZrLSme8QP+n
0YlHtxOfTcobhOjXQ1cpZhWjJ1pjAqYJL7kfPKw//XvbPIp+SGpk4sPasGMBUbOg
aAVFbCOaGdlzArdy8SpyjVMYnylWGcsOXphF5MN76CtS8dqoY3owiBzAKysuLLp+
cUUiVwlM4YUtpQPUGZpv4nAEYoiUID816k4aqDq5hA0=
`protect END_PROTECTED
