`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9xwYdaBaHAg8fG1MM/DSsfBOyyQ46goo2Z0+UGFTO2gN+uKSc4p0pBqnl12QApH
7hVk2ZZPEDm3Kd6IsVcfeh1EpqqrBiPuIB+TVdUW8b9a/gJBWu8Lv3bSOVY1+bCA
pTBulTqydEQmvVu4wFSMWfks95Bg2HnswzFNYmLAk9wUydB+6+zIpktBKSw6pBQe
Sv/bnyAJvwmd4K/BcxxGehnTtvn7ZwkVxVjiLGX+WU/GOWv5ld2xLOJKaHu0VtMr
gQL72sF4oJy9XK3mIhdK6RNkF+80qJZ5isyxscvsCuEvzGcRrQnHG93bSIleFKyM
S9Uld0iv3d8994Kp2ey4uAdYTQu4ws973ICisY+5LcOL5EwLCs6C2AB4RZ1DmSVP
mayUOa4qLmHdrRpXiHdzexfcv+CsmIL+MFbgLxbabDbODj9MGg8up65oqgWODM89
f9FxzIR2AtcqblrWdb0NmHM6nq++wDCfdQcIKaZLpeic4VoFBxJ/d2kBHwG2e1Mj
xMje494+50LaGh+ui2MVNaittjKe5FMWb0LG6CdVa7kemWwhwOHF2+vMQ9WzHkYA
3kK+DgXka08qOiBgZ9TOW6ufIKCk9EMlER+CyEDjVScgd6gbBqV4/+7lsD3v2/Ou
0/M6nYbmteiYFn/XMpCleu5jWSSp/xE4laKbtOemMCwi3DZL3dz55JtDdks6bDUZ
3kQ3FhXdhrXEFptd+xkD0uZx+5Px4sseIEBHGfbV5HmD5cw2xA5Xr58nOMZIX9yF
KDgJHROdiJbLHnwWy9BcLP/vo0VWsyntBH2/lOx08WD8/yJkmfa7X1etK8nQhYty
OImBOpcdG+gbMGcEG7r6+f0B5BvZkRVPwgfQNCd1Se0BA4gnDWT2wMIf0K+mrDOt
WglH5jtZ+MumsIeHZ9F0Vvlqc972jw+aBBDTcJ8MNLuEJtIHC2X3Vknj5opxPsD+
jY3IQ8OyE0vs3jG/v9nKdnwmyqbtWp8CMOqzfj38QrYodnDV4tGSxG64uuZAs3vA
ficTzZdqwct43rIN1W+7Tg==
`protect END_PROTECTED
