`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4xHrzgTWmAZAeUkOOWmxdZ6Rc/l4RLbyIRmCAJ6ciRKj8n0uii0tYPLHFzRIdpBi
/8vYBJpHfxy6rtAFwk61UEvl4itgeKnok4mF7SQQ3x2uM76p20uiri1AiNnnMgX+
r4tgi7vrBW8f3csDipykDWBuo2p39/+kOWNtF0eTNOMPByLmmH9Ha8ArN6WnMAX+
654oeYzZ0/pH9Fq17CpDgcxxeo1NmSq4AqdWxfMbjBfxMNEXfLBY2FwsbZaVBkwu
HNzVRVzQoHMoaHRpV0X+ySGcAwUrFxtEcjMX25Xd90bPVI6KJz7+2eQpRe6BBIwO
RGmgLZYKmUXc5cIBldEraR2GJVYfaUlFXWFvAj876uXiqy6V5IgQfZyDBo2XjY0/
Wdgj+9fKivP8CYpssDMcEOoXrz/BkRYG53K4MMcNqfk=
`protect END_PROTECTED
