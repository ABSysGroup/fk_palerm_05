`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jfH2cqsxefpXkWfZ3b64Gc9AR69jqmPmDzGu3dtx/QmNjqev0/5IYiqCou6k2+0s
BrX+DAu6uh157MGafjaI8S708fdxNe8Mxv3gbqsDPFMSIcOK0hQjB3XZ2BlYEhQL
TH/XsnC3GIkwlCapfESh6bv7t6B1M6WHlyGUlTPMEN8qOjOHXmzi6/kt061XvEEo
yVoAEJx4mMAjTByuNdIHyvrKtG44kcK3YLN8uOOyjO9DcrpbzWXM6rhsbr1OiYQQ
TlxfxfEdiSqqrYR0FsmyIESWAMSeP2XonlQiVFq+wafFQj3SnBnblZdmKLbyxsSc
bLdRbg2G+VgJJVuy+5s5x4XxoQ7aQoz0p2sJ7hzSwRAr489258Ao3mwfCZvk4uBI
3xNgWk1l+M2yCz8ofysLYTKB4d1hocLpcEBc+rdoiVc=
`protect END_PROTECTED
