`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
17B+9WnjI96/+oIazb3rJ3u35de8bgN2/5Kvnm+Pp99x+VUkp/BIr1btT4LK+kN0
ihn//aymofj8dqE2eAf4gwwLKeHBRdD9CeZW9LiP/lOAg8D6DUOiLLJDkOtHdNsY
09YMY10UvgBFN426adtMMmP8s3guXaBPbWcOsR8ihXx+MVoWgEkB/aOM9VlFveMq
0ZKF5agyb49J1WZqCHNEC9L8kwhQorMDyAd09kOcdbw7uZByLRBvJP5tXdeqVdmd
NLnkS8NtJIA5WChoILbpYW9ypINIxzRess7dauTEqxWSB2mVbGSPce59ASnszvUA
osKl0UohE+DCfPGH73bMsg==
`protect END_PROTECTED
