`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/JYdVmfMYU0n1XCdaPyfvJc3SYp1aTIR2zwbXsEIqlxU3Cmo5lSVlaXoKV8X9P7p
WU/wuNorLRD9SG/iUjVZzHfaHxloEqEpoo2C2eG9YQv77uJzfOKvJBUayfrj/vum
I6+bTMDatI9EYtSSo68MscvNep4+wAYSd1pzGBV/ElDGtmBKO3GohgZFCv4q9Wkq
xt+Mx47iy/IL6ARc0m6DwbZqJwWNmnLGURjhTTt2E+dNpJUPMLPQa04Lwl4AD6IO
KdmhsWUAfxfXBbl/yNhV/8zBaXRTlTStembhflgbzLJKyKNnKu5ypio5yMNrsE2L
bq0Tb7WTn+U/cIZ4PL/kObz1t+51VBQWa2xNwuUNdwO3+T4Kw8AwD4gBylRUNSDW
26Jq2kzHJrcsowoYOyzcwA==
`protect END_PROTECTED
