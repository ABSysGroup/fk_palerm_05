`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GBGngaAonoVvK/E6vPZCjJHj5dtlRtIj4Dv7fQRvEezlISk5ZPffQkZSVfzFqZsT
Dkb/E/8DPFIjURdvpGY08K5ljIJm8gWlqkTsukRxzS3yn55gAaftzV7e+q4nxfJs
QO02aRWuKCUWU2e1fZLQBmYMQuRgDcveGw5AhRGud0Y1/PhsQ2IhjdxknmQ0hJ7T
6yeqkl+QiH8SJicH3il+D7SnOeI/kMp9j9YgqtIc6kp76/YdMLXHaKQA1NzEtDTm
Zjm/Ocu6MTxesAI8wcDw8MFZra7s69nZ86c1b0p9LQjUxziWJbZ4fcNF9cvUJfpb
9FM+cCvZdtVEhDnLnoITHIxvFdu4NyisRbzHlDpNk95j53PDMYjjiRmmoEneXj71
w7P5Ai19mvNeLn0CK2cqn3nq5BOyo2Z6zqpZTqK83qt0Opk/r9boKOZKzJfCkG6x
s/s6zbCXwwvKSOXPHgkFHXF9si0CB6JqCtXNescfUZZ+y+3XibWRfMzNWNjOVBae
`protect END_PROTECTED
