`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
olMBP3zaa5d3yr/SSDrbz5mXDzv1UxWsDM/M110jFONRzMdWQjmp7lDlag1WXKsN
l/ZAX1OHRyuXtYJ/SQnEluZn+kfd9ECx7jd3W2Tkcfv82UcKGU3/B3Eiyq+GTfU6
rc+euyLAjxX94rmQ5EjCTRFbddmXyhNt6yNK2h9Zy30vY8Tsi5qf5+K3W7xGOuHG
rFLL9A/41Z7BPEsqWfjfgbii6T7LR40nVxjD5SydhYNXdenUQ44mqUpgmiXfRnJ5
HHKtG2x1Qp3L9LXjsgvPNd/UcfQCAqsYory1AL9k2ia0iIMHVDVnTTLW+BkhBapU
douMh2s+6uDT+QipoYPfYLI2fAx+fMhFHlPa0f3T8OSN5XI/zqpesTRz4tStnN3i
Se1lXUtswQCkPX5GoVqkvTKzp5BXHBev85SvfH+OqlCUvdKQIWod7dgDfcGPUzdf
kQTCUS/GCFMzE/On8gqGo60JbjHvq7apDz7VKu3IA6+evYjfz45TjpOxOsrw7XYE
mlZeu0EUL1uV7RQp6NzyBOLuRomNm/ZQupd4Hmcyo34ymyvPpd/367TGNNDEZb2L
8c6IkibujmYA7ogdiKRD2ClYzHHhjG0pme72IK15GMJ0vMGkHAnFa3NK1fHRPs/r
9ZIBYuBgtdeqlxIIxzALQskGQzIb7uIdi0RmdN8RmkSJ25WSPGujXiwRIOMgUVd8
JQCSDc7vk5DDaN8OPa7HSt2CO5gmiNgsF9shbkzumQ3RzOEiiJqGni+okvphMMRz
5KnhaMHd9PyGnFYN3RWbRTZpg0s4ffKCIti4aF0JH4TUTb1DZxKmam5HmH2GGmcv
FeunPuc/u0IYIUIPpd/ctaN4JJ9K2J8UkjxTGLhEe8ImKPAWxjG2rzMo7ORW5gA2
sh5EmdBJh5Y1HcVxMWzP3l9T/NXF5AnFXnylNe/1FARf7vBTDTUFVQyj89CuETIN
UktBCKrqpdfZ4T3X+FmsAUc1LdPlc5hzKAjUb88bWkPNzuGcQ9O+CWPxcMoe2AvS
kILQKJhf7sz3HISc7M8hl2bU6h0kDJH6ohDDsYHYhTHBNYz7D/Q03P+YJZAhio1+
XJLYSuUxSMVfwLAyPKclMcsufleDQdQ0j73yUGY/f2xRCPUXf4yOUVMrY8KkibYJ
ded8N/QwwxF4fRWTEbTaWLb11ncwV/0p+v3oRuaXnSh/uZ3/K0yhu9a25cuCDbVd
yk6dAzeJTx3Bew8nKi71RNm6U7COmFraBTcOnYzrMLJwVDED0vbUUUJUjROeyJ62
9Y5qgJ9c3jz64w9gBjFR/xNp6VGhaLEtTBK21MW9fdUb0lzok+hbvPo+XVNB1tex
u2ieLBBXmfAr8h9t5MeCuUpkidqCk/fjup08KIQrnHj+5WDhMZVla626DFrXAk2w
kf6zzLPVN+iYEbkYU7Kh+98v1pxs3q5qbFCVWxOB7XEWNitYJFMm96Dr7l8IMZrW
iKkp9l1xlgZ/d0lbs50l6FFvbchEUrf2HKxt39zc95aycislX+2zICfeknKSzooO
KY9aFCfBFr/LDpg9VJv30gDpieleoRMr2Wn/G8pJd485KhMpiCcqeF5XhM20jObz
cXo+2xxKta1FjfxPaUvT+OCea1VUuqOyaEjT5epxX8uvBRUJlWLlSGPg91cj0VHz
WQhZw6CzChOfUP46ZAIVLLidhgxnEU/YPMH+wD8ZebD8DIkAyX8tVcaAwqR1QJbW
mN82d1e7x5YYapIDYma9Wh9KcKHKnPsNCLRAA9QPTqiq7I2RHqFz2GYYl+YWNaEi
hnLR0xbywMh00MlKPvKtK8e7T1thKIeXAoaH7LLgL3HV2jzQ07/NEUju8B9jXxGB
ScTq6BPLybUlW1m04RGWW10e2UQsVbSbwUYOBG0crCFrb5Td72cJ6PSVs+QwIcXl
GYD5kyjPU/MwG3xoCtlZ9UE7Y2xA0lkMrQ39mkpz07crUixCzhpA4owPgfcX00+v
n/OmAlOeHrJxsA5TaQl1np4kLG7165HKQPYE2oSEoZhsN5H6vtWg0UMqm24RHzxm
NMUAOazfiwhPbDlitYC4Iv+5ec0iTdLH0t2T4WL54ficDllxkUFtHhMVWY0LWo7b
8zpfqBTvTTp73hKZbXBcGh/gmts3tnBf2XZq1gfdou2mgfhiXbb6/y62Dn2zKfJF
tt+EISo0YP39nUezAOKGMS259y9UaDlpZkqQnYL72DOAfA8fiebyKZGFSx1I1Hfx
7c7AWOEpqjuvfgSKdDRPJRYn4A7z0eU/hhlFN2FAaWvWi87seU7tDYfiWBsdCqeu
eSgVbdrPasdJYApTAVp9iI5fl3EKne7SK+SWO8BAZ3bagP6gdLX+h+oERJCfLsAN
Fr8iQOiRos7GSirfZbOnYgSFI9QZXvCLoWTFa9Vc08O7umFAT8GY5wEcTDDrf4X3
prmfUpUn7C0HkoFjkF9kt4VzhBJaF3t9ituG95z+7H8A+wSOPhNwZbI0t/2xZmNh
MDFTvIJJaBm2NIHihhDWvlmryPW/BZ40lON9o+HaKJ/VO6l4ixbwGlw4fSgRsHqb
LsqW1r2hMf9lb4hGyEmzxqBoQK3ufvPw4k1Ts07bqHfp+i/FTfyeTS5asrAuwwbN
lmXL//saQJgQDO4gDDCLrORQsCf7slcs6iO8ObmWVQrvNAhknsf6bSoxDkMdskXO
7ggFxsrHyiZYn06BxAQfWkGoZFul5rRyU0cnqAZGPb7F//aqBMpAym2auDa77pzu
QmgOQtzhapW1wziez+31eGjFjn2yQ/5L1/x1LamIfuWUJZcFxPGWGkV9dLh0gmhF
/izr4pjFrJRVcgeK83GASDIqgsWi5kGsSXFOE+PDGEsoTK0EWa0Zit2gLY79YNjt
rFLWAIVhqkqneusOPeTue30yY7RlA7Fb00mgucOTwcddZ/LNXVUJholWWrAMzWjW
+vmP5AwdGaoL/wRQOldvLEkGi7UGst/Yk4XQ63e2AuO2kVsj6NzoK74xTgj8VRfJ
MHwjd1GakViOXSg1EJDpNYHJjSU6MGDAVozHauj9dcUPWCnQkNKrn26mNCIq9mrd
0RYDk2xr8qa5oUE0MQlZSkLxuYHRvsLUQmaGQgtt6WpSOpY3gS/4EEKkqBCxjLwF
GZ7rC+JdmvAxMbNf0PVCWacBr2jMw/td+VT/4CnojDcHQyft0JLVoV27Ul3Le4gS
gq0Ode7dqL9W4MysvlcUNcYuGj5bbnaAKjswC/Nfn9K8Qm6/LPv1r/NVrB4b78L2
tYeY2DhZfgJL5jR/85TCvH5NxBjGrl80KxkUmotv8JEE6kb55UbsMO5KcUffe/L0
bOgibD0ka4/vHVqHxD/ROl3zyU5cb2iX/vuHogO2I143j9ma0SAE5+mcE1/RUm7Y
igDAJm33j33xzoTtT7e6YcR7NXPwwLhebTj8WdL/An7m3tzHZiaRLsj2cK6tzXGE
QPgBCF9Z3+dFMs3pT6viPTOIrk331nIl/CTbHIQctQJqgn9bA+SdvTxj/5+0Uv9e
BBHBmB7FtAtvkadU8OtKKK/uP/ziZczGxGSYT/RSsiiCHx7dvWdZXO8nRUDBDXF6
czWuHGC89sx7pJw8cR574zeG1tR3tMw+l9sXfEx4vLshtphRg/tu0fWlNkJ/rb+D
Tbeb6bkzbhJ/qXmg3m5US7ZL81QLHygxGH2apATznBb54Kmmk/wss6wwyuIAU+/S
h6ALAK4OfmOPaoFcElPh9JNSGqscfRtCV7Df3k8ibSUCYFwIKnl3gMZsojG672A/
0hyp4OBWBMaYyLnC8nK9MXe1gvRCoqLTYM4FvYOarEeZVNYmMxD7xjftugbu49s7
ntjQJnmiACkxRXv5eFkPCF1CFdknNCeDDP822J6BbGZOP9P5rZAxXBbX399ix9Ty
rANPHggAlHPUioymiTU4tRHyWJinKP8i925R6C7tBEEWBzOko8aglcBn4LVEgHHb
qh4II+ahKyAEglHAZHfe6l2A12yfSD6KBDLl6oi1aOjjedl6veL7wl7NGbuJmB3M
Oo3zNzrRQc30b2kBotSPkD1qxzProa0Ic1RWOR+iW2tkNFlVjlnMoWDbga2CU+oI
BVenyH8TdN7cHTRoNoCSlu71cBnW8MtPLeXGe64SgUjb7y4KOoxZDU6RMw/Th2vH
xDNDOogyqEfe8ATMhKhRc87zhbfU3XZHFWxCQbc5kI+8ouAuBX0O4Ibbn4EdiOy1
LDz9bPlOgOPbhE1/CKMKhHGOl8edcUuqb2mzm4R9ECMeirL0+C+Cd4DO7illyOWE
AysMSwrcfzacrih4zqkDzgUujhH9k0yQjKjuVnCTnaoBV3/GvlqWmKus0Dw4uSIo
EjSLvn3i0GrnuOsU+6yNGR54Ahrtkqi6imhq9MEKZfBDi2WFJdUnhzIRK2QtFPKm
mnqVhM4Ep/TwoOwdUEY45vZSbw1CUx9AsNGgFA4X2L6xpdOMkL0Ycyy69Z8ZwyN6
xARqW9FDqjiU8U5+0glE8JEQeDgwMtBunmNZNqi3ahDBbDWmay+TRSPcd+EjpMpi
G8uhtY2FkgEGQ+xwxKF9B9HWzr8z0HGcGiOfai3RKscQAkedKU1bDNZUEJZyyDCk
vibjLOUAb7avR6MIEU4IlRkoVDmiSggDHFaMebzB6Ud1jtPOLBsEwTaBUEKXOJP7
chvGIAnQQg8aWrn5ZAlQYVhASiB0WxwZhKg7iTYC6DPAR5PU6LIcQHOQ2lRlCYcW
Q8nofd54KyR4jI8M1DjOfR8ZlUmwxXzKkUqRQh0dgnfHN6zW93fMCyO2qkwMgZOq
OVc9ildYM8vAw1yeVmhSe981xswl83zsGkQstmJm4qNKI1Rk/2+vPz1BTRA3b8Dr
+MNhChzD89x6iQ6LLjiebaGUejF3MkqGOXsvJ0S0MMXatpLNe0pdbtr5GHro6lY1
/TxjhWY1pzOgDDMh66LnzeeeDHoBH9CS0QuZs4VbrqY46hmV0fjBW4h54p/GOkb5
HJKJjlg6A2jfYksPrHf1z6KEfP5tqQBNsel63FhaC/LvfTo+vilYMSga0ZyUfDQM
lbEC7IYu2p0L7Rc6yBzte4HvIwheHEYKP68lmcE9Avn3HEMlZEysRPUgbiuOqMau
OJLwlE8YGuc3FT4uGQ3BTqBNpKslajAOSVZgGRWPp1NzNJEOArC5+eOxerpz5aaS
u2XjWbcqP8hJ8XpxA8NSuj1p5kTuXzJB4fADhkSZSDI213Pa0nYpNYAo5RTM64y/
w5MjQ4AKQ6CJye8E/UgEpLJLaVyQwHsNnQfXeOLRJbAGaPkSx3eisQqYLuhNClqT
CtorO/rtTRFdMF/Bp1KEbTCfiNyVkG9T+F4sT288MkFJzxA6/7FfbKkSd7fzz6pJ
IwIV4MRJw6QH9qK2fSYS4p77BX1fGc9MhW/bL2Va/72lU/d+voxO2E0k4aMfbsDq
bb8p4zwBle27QM8OKsf2TbNipS9ocG7CL798hRM5ZRqMNlXdnExx5j1Q8zMOKUx2
N34CRHo2YgMZ6VUyYbo6WTRKiWb4qqQ66v4CZLOVz8JO60Rb61E6p0WnNa8qkCO/
I8vJH2L8sPhKNQchmXyDkSk55gON3+kCGqUVAToJwt5bbbs+vfxGNbwjoa8cdjmY
iPP6WMKc3QCDlxC9xWaUFWR2pLGSFzB9kEthbg2O7PCenQyvo7FdOan38igaOYMA
wz6V102ZQQaeaQ56fdWY0VNx+cAOjmr1Bl4n7LzoGqhky7tBfWDNpUDl6jWdHxDA
6+3IZOKKRw57YvEZraO0PgOMPpqd2fJLxouPNAYscJxY4heR1uZ2pvz86MnHkLFw
Sdoh0NR2AibCSZ24eaRgwg+s31/VeOsSlXGvHsfg2FaMMEFhQsAm4+LDqVMZe9dr
Yv77qAOr875dVSIFdLamd6tX4W9aoTW7TAd5tRTdVojpICpyhWxKT+rJCwKue5kR
+3DO1V2BKyLilgltR3+x5yLpUQjUS5fLTdSTtZVXPcvbcN2tCdDGxiiYB1Gb85x3
6NhoBV2WlUlEYP57exlEiYAJYn1DZAH/RJ/Ic5zIMpR+3Ej681NvHFlxWpicB8Bc
slflpqKrByUC3w/CiKbvVVXuLkERwMPLj+B1fNkfwn/VzV0qpROhmp7cBDKbNjXx
uGRQCZPoF9fm8FYUTko1o4QxvVfnZwRtXb0EomC0PVcCM38sT9ybusXqcBuilNfs
kfvl3A4MLOlf+j6pG4i9QLGdEMTySAK2e5+tpjXd9F0E7McmNNiO1WVTDYAiihIr
U0Zxte8WTa0XXbbQukh9JcxViz3rkOuiqlXOi4QWuxZ5/i8rb3b/81SfebA3mCdp
pGCESaoJX7NQ1HltcJTzaNpV5Tz0Ai8qIN0uTxfC7g0ds1YYgS6h6qO8uNU0HfXn
qpvbYmS+ZcXOTrvCiJmyusSCVoci3q/FKijTmI+X2vcO8oVdNLRhdbg7eEPPKs7g
uxnLEeJ+GlfVsbOEzNn//tY6t3iDDuJj9YE0HvDj06V3zeNDN/TBvAxdlxrSeHZQ
P2Majnle2OLdxBB0aVMGmKIFDQwlQmnAaEBtDgi3M3AMvUWiMLCB3wbpNMOxrOIL
6QiP9vpjNWiA+OygoH3zsvrNkwHJ3bntf5qnCyJaDeqmw//DsYNJ+owOS4ljD94I
UhjHXWKuBuGRH0W7HYkJdzN/w5bCpDNPIH1OZTh1yQNIeCaFtqylPwgrtjt0hdT4
ZA6duu/1NpT1nyBTOLa6Hn6E3LAVvw4SRvlah6tCDMbHiNmERfhhhiRoTbiDXptu
9jFut93mRaD6JOQ1Q0ZBe/twIdSyuK+/fWsvuBgi3FKoO0lLMSdg0E/QrssrMyWE
1hg2z8ytBjbzjJroDVgxNTlVxZ4bRQm12at2v8h+8DIzWiSDlW4j1+vTjMmWtbuS
R2RiplZzBIV4MC20ZOm8VJBn94ppbYyRDIi9r0TmEt8fafKi17oQfbkr6mwAbvsn
dKSvJPJpsFEb0yJoxHNfoayjVCdNXgkwx4r0CpUzoHNxvUC+g7XidHuQB6BstQh9
z6posdMezcN9YRh2geh8ii0FOlWbs+GviP7scvneVc1vGUJeEs6pnqJyihgXjvQO
2dbjp4LzjCR5f54PQu7Oa9GhwDpJJpOpUs52Zy4G7Yo+KFbXsrro9FJTu1CMHyQX
MvV8/3VLdzSGc59AuamC5+4lpCuazuRxDuWtnDvB/Krz0h6FkingpJWK7uj5tgEx
QXDk/K/zXGh+L1+ku1+P4ZVTyWJbF2i5+M1YcpL+5NbrdDHAosKRw/V4KsLWZM+Y
3uZLy2IY5G2EEXi+3Kq3RPznv9CEWkXnKyE+niTgpV4wb4IYi9Pkyf/iHxQEcUCQ
OFc7AoAjD1720t+Ff11FeWAuxcgbuE16DwFGE3kGZumiGAyQw3aRqOsM42/0WJXx
yt9J4ZwjGI104Xr/EPhJSTsyivfXLH8F6TwAi7pn87DH8GfsR34iQ35gQ4v4UzMe
BmDoV6DapCWNNoyNRC0Zx/xpgbi3a6ikp7sGydvjzPVRpi9CuhbGdGZuA92Cemfp
41UZ7rBVtYfjX9oB1Y7VtPUM/Q1ccJtbnxLPcUbYAsT2wx8w5bmWPbn/5D5G08cV
6b/ErTzczLv0X3Hfa1uVSkY6uMarNLIX1avFqaB4yPc7QE9y4FhZwz4uWTRhT2nn
Kqnd+VQQpQNU8FIrQgj17/4XACkPet6otsDmVqaAkUepiWGCuNVfvOeGc7R94T2m
jBNW/7Ejcjgmmz7pm3Yb2Wr9F5C3EQPek8blqQ2l2/Kn4ea4ugBZiPzKexQJ9TUA
rHw5Jdfg+zBfThu9ZvGPenmRQyCcy85rmvxd6Bgy3lL6eVIyZyj+qKi98xgvxYng
W3vxv2G/8y+tNLbD8GH0Oxdg53wS9m1nVvmJ0yZmFdnyMgEyVuB90F/xsRjj50OH
f+gN8pmY2Iu3SGy/OmvWRiAu3O8grvOFe6tUv+nVR3fzTK1XE2sTYvNMjWLDTxKs
GkrIte+Pxu+ORTrVP3wUkfxGA5/u0Dk9AFOEh3Tejkk2b6XMrGE3Ox5nuB4o+poD
+CYj1UT2DuqkzKNyGCH/hGtJNtUtBq7WWo+bt60QYw3UKfib8t38Vcfkx4YUtmaG
kI5sKRDTSFyKuPcYksss8+4ASebw9jD7aHKX3LfYazHxEtiweuJhZaKwAceYXSnj
l+hzvHUm5FDMuyhEXVnTDJIsWPqQ+vB6gHU2pv1B9SOxgw3v2QNzyDx+cTsBKDC9
7nR7F1oXt7XMDyeox/SZoZUA++LcomVpKRZr5/67EiTrvxzdVa7RDuBgGpgGeUCh
uuilST2EfY++KhJds4FS44HKnKNqB34zuNCi/ovl42TiWK1wDMFT6yQjS8yS1aRt
1tqyWOEFq3WLytAZdu/7pqUGFowAyNYZXpsTOAOlNwz1cCducp6wJjz1GqPHQwdk
+5KG9KWPaCP6e75hpk8BGvPQZcNROCWzXfNqXGQFncH7hgMaew3Zy+NZk+khiuVI
NxIjgT2PUFTu3wejZwWvXUFnFWUQ7UDgQOLzQo71XHv6Ua7GR2zecTeXSdENtYq2
bt6WFYhmo5kUFk3ank4AQJyFTnfP+wJxD5rMHBj4Cn/gD7HILsX+oxFtOPiap07/
IjmvcHMh4etoqrueRp+WNuvNTdBJjgsnrQnBf3AmFHSZ0Drn4EIPHqrJQLiFCQRs
EFYZ4+5F3Q2RCZS45oLytMHqdEr+KGciELR6YmkpA2WN+PTYZQKR5mea4RKNs4RV
QlYx4ej/a+8ptYP6ztp+L77xa1JkS+9iLk4q96SoQuy66NsXkxKCbngGY7MehGjn
06QiyBipa6jziDQ8Jrnc1RaSc7ha5KNwbSuBWCJP6kK97x3K9MTADhTnj+tx20CR
3+0sfkR2LQ660V3LRRGdrPYatRxrIJairA1oAJhB1pZt/Texu+v6rEwbf5tHTKJ2
Rt6pzF7YUNwz6kP2a15ADM7aiC5xwBYatJnJHwBwAF+05rIn5LIhSdXPDw2ULShB
EZe1aCbs9nItBmrdppRCKULlhMU8jUuHCBnzJMWas4BfoQX5cSaaSnlwH1MAcbmR
OytX3BYcKj97nu6fcpMEdZaSQPH40JJ+8We8LiV7HBCmo+goTBSKXGlCWnRNgiWi
ME6E+BSRhuIlEWqeneM0Fnuf0c2FbVWcOnm2bIOtw/GrsB4hkWpBoWxeTqSQ7Sw2
KmRfOGmmNFS6oleGJCiU2AqdYiWosyK8gd4kE3QG5VQ8GUU5LEgST7bWAqbUjbhb
yzRdpXMtWpQ9qbSvY+SLp8xv/dbIrF1wU90vYHFq5QM3AFG04q/uGhkvs4w+adao
v/0x0F0sll4LjGZfzAoQk1xzN5f7VPyhDgS113l4PtYh5wbGu/UK00+VBPW4fGfy
LAjwejUlhe7Eam/NZ9Foh2981XFbDA1Vt8i86YdjbmMfUqNLizsA50WeFMCTwLEv
pew/5hRGjQ6HXRaAkOPWfa5b2ugvWis0tvQmCdWeg/hA4Z8lKWYiROUDoyQMI8qr
9A0O5BktTKm14ZUbsPct0wHikX4/Qum7q2977l//D6QJzszzMYS0EcEels6JQHBK
+txXOLojbJbEFGgCRRtzjA0nn/+Eg0EQiDRVaHrDONplSsJlyM374PjBI6McaBrL
U93TB5HsJTVaGxcDUE6kmgL7cKYGcQwWVg+gTBTo4na4lvURmnw3yGcbmBnaO7oi
aa28XnOmKQiyPRTd0YmAklMe1O/QF9i1stEVUcwDhYEXho8jcu2maxdWrHr609l7
0PaSs9vhC1qPvfIT+VwItobzhxaP7/o3299CuUCLnfeMVGP7zJXdNEyDLPgZu9CH
APApOYWM06QKA00VyQAUF3fFUNMcvg8q4M6nvkyx/hKgrg8Bcvt6/Z3O1vSbMAvx
Z2EFBLWxs009wofBmibVSpIH6XG+AbnuB/nFIz6Wdx4im2n4HjoxNA0KicY+Zp8f
uYKS/I09YL4+xeU6p3GR66kz3EC5yTZ+qLyvUMmbt8v/cutKpBo7OUdF+JJWiGV/
bgkbnshaaaWVLq+dF/pS6LTfs69+6dbvaLiKornBV9FLVPkYLNn6SEc3/j39MvvD
Xesu/BkcZTXSlCeLaqTTxxrRRr4pU/Z+k6iol1Lz6SY/DqKGWGHHFD1tVhyTviGY
mvZwbBQv4LFwugdT2/zNqUdRQpbno7O7/sva/3/RH/XZ0EiX6jFf7stM7UtAMgQX
Lq4dvUfZuWhK5F8TtlxWtpbdh1LZ58bdmJRQ3X49vyB7vjWUj7/PzaSDT6Nd9iwD
mwZz0KXFac6Esrl8V2kxCXDOWvOYDLDehR1Ypt4bUD4V9ObKXINtQS6buLHcTrf5
UsM384RjXDeRMWLNArK9zuCUxiHiY90gcbt7QBdY6Z8IAwAKoxV3OS8fWjdP7sZB
rC6IhKf0fwLmFpzk17CxFtHi7fI3L6lLpWNYtCz+jFEMybH+Boe37fPh0miuLsvz
y5z2lv1ZExozozBkc9lfiE1mcbP41jKlPS7sISh8iIL10XpZJ33UkjiX95c+VcQz
CYSRy3gSzkWXUPVh4MvXJLC7EYxAybdmpSBemUjn5LYGdUlS8IhFHHGKdgI86V70
c9SgLjDXuLQfNg/uKbD2xrumjE0myhM3byYUhULUjYlxakK+ZU1L+u34HFuJDGHQ
0gVEFbtpOaOvDEXIp0jH01MjvBxeZgGnFclXoQvk4j70wQwQxJUo5ep6KyTq0FDX
N33XiEq1VTnd7xbigVj+SyRt46X49BYNAu3DuW43DfcfaIgc06Jx+tB9jGaqYHEU
i2RC+IKhT1jibpJs3m/hJKWibEyDtAWKqaIoj3BIl7gaJqkD78d5nZzjaafgMKbs
DkSEfOtDTkyucMYbp+Bt8udJ1E2EOmeLQqJMOyyoxZnFelQZoyRXSe0ewH4cQyZn
8wkrITyRANGa3mg6caEuof48+tbqgDwoPXVD64I5jLG6f3UoLjlWn/PlC8riGFUv
zbBLV1by1qyLsS7Ek/K8u7Btot9q8QnhV8eCpDE+CrGtJdM29voEN4P03btJa5q1
MEWTRMSGJ6v88DByxmLB5ykIrinjOEeO4bBobYRm5rTsVh77i+bCQAijU8R5ONlh
uyTAD9oUOChLVgr5BlHxwm9q3BrlY66tVvleVxDw9JTgar6TRk6oJE5GQMBBoXyF
c8tnw3uhMdEY/yJHNhHzbjBRDPzPodq1lMXd8qf9LBgwI5/sTxbEroYmiljOjBxO
Bnwpf9j/5UKjV9pY5lW+UW7SxEIjdMkVZWc0NaENvEcxfTv0HQr+DIxtqyj+XRpD
4n64WPPhhVrXe7MtFSYVDJ3/SKDRNLWgdkVM/jsx3wAtXmVFQzRW44R48CSdKAo+
Ze+3rNDHCQhqLViDurzhmn6bUsKJQ/yKcxzrF6zzc44lVgAsMD5Qe36ggqn11wA2
QZbUI6pkusc734ilDMoXfbuHCUWA3ik/BkASsdAJRujy8LeTZz1E3fSJBoJ/dST8
U+UagskwbmMgCwR2xE3zt1wU1Nbu+a9n5aNdrUFNeMxXsbJrdK6/XUkJvoA9b2I+
tB1pU6WOFllpyx9XB2gQz5AfVegljsdr0ePz+U3eE/j3WBHYWcSEc6uU1szWTXlU
ZqTJzdEjc6K5S/Yc2y4PFYeaDp9xxRjwAYkkENbq+11LrXawMmacMaJ9Bf3EFl/Q
m26SAK6lXrNo7+PyL8EkDd9G1sP/naja52mFV+CSBqk80u7g240uk2RiFeGbMfs2
yDsimCOSlR4M6Yr9w91US/SHTr8T9jnTZsCg2VKIZkqw6Ux9fRsaJG3PlqpwLhWn
CHJ+d3wJC5vqjklbx1StH2rGuFoZqKOab1PaFRqZPkCPCzJ889XcIzH2XaYz9Tc6
+bG/lAY2V4sHQtYvCVsSeoqxSFVOEaEp/5LPb3VN3UVyTYfTGQreJshgJK/vbxoQ
AEp86cMz42OG5aSri3ceVZxjM9c13qU3KjNmSlWIXudLRTxHh3w1g/p1dmDzoTVv
PEaexvZsNtAp++Yc/AKR2Cm/WVE1xCMD3PeNlNIGno+R/M12V7UOqd5ybxobgFP5
mNsE5KQDo97SK+q6hAfSHU/N2cpfHqlYh3PX9lvDlBFUIPBDQQ7L5A1Mms8MK80Z
7UtNxcoaSUirVSW+1rtrXN1Sh+tyVwNVDilk3KtT1Q6FmJr5KYajes23jThX3kdv
YABFehCTdicqhMSGeSa1NCklVdYVk+nEm4CIHZfF3nipAu0OWPuHg0xYfcMSiR/g
BWLnZvRD0kGf8wXc24AC5whaKCPBY7Bij/oYlqRLm5mCZxRvERvmFZIqQMslwp4O
n+NSYxPpHMYIBJcJrYb25JnFKx4f3LY0ugZCStIHYqVfFGIn51pMt9MP+nbiE16J
2wMq6Mt+3F6Q5dO5pAGZYuZA2cpc13q3TV3sBCliGpgtudBnE9usRRfdcaatJ7l3
9hryUPt78kkTYlhfnEgRp9xLMZ+Jm1L8jUWpndKPj0yt3DNmVrFIN8RaSmED3g7+
Y0id4Tscn+I/NLB1gdJA5teCPdfSiOd24Mb2+2qNGMsuTIaSeWmOMqUt2qCHkLGO
iqGkFv+3Zf6pr6pR4JhdqsB/UUDOd5fQQmU/BgWeUUuhmbKseW49QRBDRdieyswq
hV5Y9JIxafU++4VNnbwyQj8dRslw4Tu90Pbk3hlNANi6KsfKub4crzlDbjmgxs68
EWfrBqX+1VevSkcvudohvVkac0Hun7QpLVkcuDx6GmXNFVBx/lFqqYEr8P/VMu3H
tI4in2GM7ppKQwWGbSqYziYRRTt+gbhLg0lcn34XN/vpzruB9h8G9S2KM4no4p6j
cudkRJKWiKMxA9ci+mRZS3/kjXOuWKWXjy3cgCYiNkKFdRCwmMErpEWMuRDoe2zK
d4M6hm+9K18cZb+R9koXeyGV96RaDYeBfeh4gMBAv4X2EUObJWvLz3Qp9cZXdFmY
n3ojCsTAUJYPhPaEg7dnvRdNA43P/megde0PnkAwUPjGhZ9t65l5g+9/qH104j8r
ZRtD1umMDT100H5/sga89CsjNghHbRWPdZxjg5Dt+c2PIcfy8nqwicIDbDL0Xycv
5UyDz1zSUR++POn27cx1dn4aJLIMXlcAaDD4E9calg/eCMBNcvJlRyXjz5f4xpRj
OIX7ZXzgt4z6KzjEuJCjPGYS5ugKfMF8N4+do0QiRappSQsQe1sB/mszQHz+wRhV
OGCJ9Wn1bdWzjY9ssUGCyXTIJkB/uD5rXbWTY6VJSxJNuN/Koq5akCvPefqEEn/q
CPEGT4+2VoxvCcrEXL0W7rxdtWPf7llL1pfleC2vPKuykQq0EWs78phLCVAniHWq
KEfZ1zw82RHTd9PGsjUKgLCRyPnoNq2EuafabIbNpBr8QCuyadl7ZLiceuHf0slQ
TIYxkwYYXPAsNbClPJn9ZxSKjlDhYcCpHiz4tnYlMvW2TE0sJ8FE4loSxGqZ4K/x
W9Mz8Wce2+rVzh7imx91DbxnGGLx06zngdHl2n1l0oQ+GBfveN+aVLXNhGkzOyct
hIb4KP6jxRT2qMFl+Y9QdyEUAXyjIyvoAsOx6C/6D2j4sqxd6RZgPhwA/u08N1wV
y4t/gzKbeVS3JJG5ksF3p7CZn7vR/xtpWjKT8+gDHEKnOZRhjToheuPQy1Acx5RW
t/qDYa9XmqNOZ76CFXxhQCmNE3RoyZpzj4vJL7DVGGSTvP4UX5vdsysOoHXarVOK
sW0zj7L4nVa9ETOXTry2mkdFZ+xl6HEaWAIJlCTd758F35l6Dri+LVLKbli0zGM3
DkbDGqUOihGKXnlSqQObnJlHfzfPddiaETkf6qgq+lCo+/VICRz3cSGjkFZ+pJCV
EW7KaQGnK8kH221YWpIlgD7fzgp2ytfqZ3Vj3Or0emNt7SSesJj9dnLBaa59kekO
Px60zLUGQEIcBInRvtC7RbMnZ2IJRP1cCHvEaMK1Pe7qwsUmQcJIoVZkppBylbnt
c55sDZY0kwhScFGDsAbrwJQ10bjywql/Qx2SZ7UHqW/WoN6LtcDRwmCbAMAhobZW
emAtsbDpIDbi2/BZyZJaO19SbGrElvYsYQsY12wcTfojNER1OTdNg5fgXuVdh6Ns
lmbLi80HT4OsY/jTbLIggT69W8pGGTdRx0+2UQhdgisupuECe7ySyxredVOpTeep
Fk0PGqkoL4rV1cPrOmbr+Mk9uFRHuLONlLwDkpEbi3TLRKPDYOf8nJ9/MJb8XxUY
mI2adjC+gsU9txx8tyAt4iqu1cl9R6X2rwI2MRk/H21RJ3xYfIdEGDWreumftKGy
bKp57s3nFImUETkYjH7KjU+909ifMh5OJP/YosE61IZSzHrXH2zSNg/q33X9V0bT
h2FZhBNbdwMnIcQKon0CW5stvJS0lwrJWJH0NUaCTLiQt0+T9JWeO1YQmp+bFh0f
zPXQnucqxQ9G1diiySW6k8GgeCcZbWIwyeH6jVEfpKzuzzGOFo4EaUg2BXQP9t7U
N8MRRf+BlckiQQpda1KrNFVcL6meXvSX/FMgd1l2e9E4cv7or8dXZoJncoPXUpvp
UPQH7eDtRGkfDve0VDd36QoKXRE3gtnkbA8m9akN0rRvlS21WdBwjNE0FHMmqF0r
KE5WE2zLf3QLWSu+I4uWjfxyfV04JROj+8TxfPHseH6mepNJFyNzi5lr2vTaGn8o
Sj7/EFLTBv7X7w70FIQEVIlRW0NfiSbxq8Xsn0H5y8Pj3GvZx9rafjO/VpyJTgo4
db9MbosmE6tCY5tDl4Bf03pm6amS64QR4RCLI1TAQN47RkZFEMwFqcrjIij7Tgx9
zN57lKLkeHUJJg+I+kX3O3kgTKnDL77SbQ4EEaI9L8hEicnHBj+r75jVyDSXJJN0
+61EhHW2x5Nnn+U+mvsXriDEEzGanzkeU91FpdIJjUusxaA5ek0W01hKsbmfSR2M
yfj9AyuDLaezB29kZcY75CL4C1au7gGeM+fwozYmKaWuVYT7x7g8KOj0CQrJ/pcN
954ETowgs1wokHLHpGDg+u/E8old4CCw8IdkEamTNoTlWZjZTzXT4gRTYB4euHe9
fUtN07U5bGEWygybO67P3HUbodiLTJ6W6LBEiugysIfeNiwy5mrjifbqkwTMHs5f
EExxhi0Y9eCpmZk3fPDiRyguzrGDcQ8E6SS0vpBlBZA7ErZoAbC+JqmDpyLLvWWL
8d030Ywm51gtd3uN9EJeLtXovf8itoUFilOx3Esv6Xa0APPtBZKj/VAioqqJHr5l
451TNXvZ0hgR7/ovT7AUGcZDloPo4zvQCDfUWF06dsbq6tRCnujPOTxJAPOu7UvM
RnKe9I5vnI+mA5757ZSHYlmt+zW3SQ4tPLvCxULXllyuaHfD79IKaLd2EovELBWr
VjZNMdb2zlIvgWyP1EJkS1LPOh5CXnNatoUIh2cuDxjEdn3WK/xT3vKtNNmK7g/V
xWsndChwGmEE1zBPVshfgOXzfCl0hx9ZQPxTHjSJ30HPSY9b2awOW5UujY7us80Y
XWG92Q5v/dVb72tNxhJuyq/LRMpR8TgjDiliOTt708kFg/CtwN7MZwk3SCvnIBbn
9qW1S1oJaquT/cL7fZNhxnf77AgSV9sF6WDfDOfaCiGmjcQSFcmSDR05zV8Hdyg2
GhUrVT7ptLGkWOO5DJXmQK7dRm1z8D3HzsqVbQYC4HAn2mIhSXVQ7bEHKvVe88hW
bOQBXrzRnsJcukkopPe9L/zXEeUNC6uJUgAHjX7LOUnRjIaBLnQS8R9D07Wgov5P
Qm7i0yaA8s5Xvz8PjhA+iNy5Yb+80pBWoIz2+w+ghyi+EBQUAW3LHw9zzEXCZk2k
DFYXiLmxiWCUZFhk5UQLzRyiD0YBzUyVh/1te4HHRzr+md0AygD0Wzb2RgKQeGGR
rG7fu+yt/k34KSHUgaNWZjYBiH+FtnyqMYdjYL1goEiL+sfiRnMnOqVTjj0Qs2tn
T4hTfBUn1kdz/LIHkylEfympL4nTNfc/Jn9HoZ8IwWX+hnFxZ7WPqOgprnXMVCEB
M6MyQ0B3CORsGL+u/25Xl/k46K1GVXLnXPD+PI4cEk+x8isjUFVhFTc3Vdx4QDPp
n5F2ZV7Bt7pnF5+t8h3LyvM2iIO9dEXPPnqFPeYP550yCSZDYReMEkFw/4ExBJyv
SSOT23qHu4BngOPXqGagS5q2gheVw0L2NEhrmJqIG+Th+NP0SSITx9nOaahyO3mW
9eliADgwPBrUT4VUaS6Kcw78LAxPx8WbSpnXyAwJWJ4IkwopAYVmeq/FLKJ2OsKv
ZGt706bhHWqQkWMvV8p+22QmyM6jyor09YDLuoJzH/QEdER2Hzqpv/ssYyI483Hs
++h8uMkr/qI6ydr0HyJxPA+2TfNgcrSEzO71FjaLLr2DxXTXXRBa62rgF+jGuVyI
G1dvLa/YinB9XDbdMr45UvhMO+KNnQSeysV9oFMCgL6dYE0V8X60oSQSmbYPnpP1
1XHxlMc330VGyM2x+MTdGC2jv6jYt2UVFkHePmIiC8DHtG54jFftc3d7QxaK5vzt
SJklopMgp7gUzvBOxrilPfpqs7/WljUq0xNg1nNignYnb9MvNniBeGMd7Ur9jBpS
CbWozpi+eXc54xj/dG7liC0GUgkRvwDnx9p7KBG/V1hzqBVS0rf5ZEVZyMJh4J9u
M0qbmasapgxBPlFWw9sn0vitexC11Qb69jVYBkjwbrkN0A+xEaawjjH1c43cTno8
AfwKR0e9atZEFL6QDyRvwJObMQfhkGsRWak75iPpldO1w3deYgz4u3mDjDJ5WltN
8zgbIuqNLuaUQeGupiIbiIrAOhFqP4Q3rmwsvKSEb47FrMm3wdtBJCeW4dqNkYuQ
/e1DxmzY9vyrFAJvcSfOqH0Ec8WHI1JA3TWSQNDCPRkP6nonmRxjhd2UrVAB0pLC
pampxxdI89TN2c4NC3dN4D2Bpp3bfAXrOjI3hjNJJXAL4llAfM7cujS1CHjFOGTu
FSI10h0NPmBgFrcDiCQboUo2lIV6nuGHFLgYir3WuPtJAKgP/TTdBMmrtBsonpG3
EasUkr1J55qSFHQsdrhF7C2ZoCdo5Puq7of3DtdD2rQOg1YBAzAcMhkh3c+VOHsl
B7Si/qNikQIbhdl6aUQrzttrl1Twi9vL5P12OD5ihC8Rq01niGpJgPhP1dotxy3t
5lq/fhZn2LVDbthGL2hvNhLpD/U5Tv6B6xRbdi18QF435sqrFEjYAueSgZ2wpxxn
tjZkQVmVOgyXJL9yHfUCrABCdC/+qhaI/H5vFoVv5GMOUCZOVNE09tTYqPgXq6Py
sqt6yyiaOYe7PTIr5Zo2nyIH4iUyCLCII1O5lVWskkfszQ5ZYN8ZPVv1NK/FfdB3
adzm/d5FevxqAELel5REnOuht11aSjn7yh7uqcH8PCnj9adXbSlNIZj/zRLi0p9N
xMWq3b+jx9+6trNFTbIHOWwn1Nv2Eo6IQvKYdVJj7J8bYPVvKl12z+TXMbHfYbdh
Dxmwaixa+CUSpiviODfTEee+YpopQcRH//SQtHKC0H4Q84WwF9205o/2mpMN2txc
BtudXDp8fGibSSwXWbnIvF/bAdnYRtpYcJjZwsDl5kOln4tLT0gjScYSGutxi0lQ
mRzvgj+UDFp+dQ+NZn7dxBsoRxEZ20uRFZrA4udc3NimCsH78wAvUhr5GOc0clw0
j0CT35Ft6XxGWKAM+EIEeknn2XvT01GF/qD+I13/LUgAraBB51wc5RtBseForFqZ
uiW67xvSHa8UMxHVBJB1BPsUkCJlSUpwmP6u3p7EkKE0M9NHAOR4t3rrns5B3QJM
fHL60j+WLdFsZ+wyUkgMZQ1G+j9JUqZuZEon2K6e6k4vsxnuNL3JJsqKcaYd3SnT
yBb7pUasZ7pn1jVn5eMe6pwGKVhPp+xGfc9bGRQGVEI8J5XCxhyoBKcwZfrxjFDP
HTDpuvYWBNM5rgGkOFuFhI3dzRp4gnZ+iA6LmKV47+yVqL406nKxqmEGcc1Y1Lek
xf4h2+7ZQhokI9ltRnQAB+m5xbT4yNSAoa0Ik8mCgGgRYIq/v3Xk0TCWdOk0eupG
ZSKaLw4oeKArRs0sbBOV7wxRRUUPiOuFNjFthIjmBUl9Q7NlT/QbvO7BUjQ9z2kK
l4b6JXUBM1T4z23tyaOD3FgWwUExQ6JxSMrM6epRk1Ru1bOyZlD2voGjXyFFk/hu
Ia3NGBuzKWaat0yf5UE70s+RSeb4rWRY5yNPR+o7fGEiO26KDzTPzSC6FIPE9EM/
O8oZY+6cmjyXuqGcRalbfbiI8VF1UfzcXhogAbOt7La0Yb/nHx8zYXpOGQNZuvZ0
XiFzILBzD+Ikwjv/3iAlJxkEWbtE7KquBiXZ2LjpNIBr9/HgaPgzxM9fSpQ1JZ28
FA2sF2IHIbbgL8xvnpRqJt4bC9ouDf8d6frH9mf0Zpe7W66wBYaXL8imurrsHkc+
Bfd0BpsKVRPcOjwj2damdYewpDQzy1mdWQCxDMzRlQ+XQc+ziC/xQG5aY0GWXSPk
gUAhwpbPawYbd2X0feCnEqM4tYAgcw06byireskaE0F92wZR+FURTvd1gxhZOocg
iDDpLUCzK650rT8zXF0H6DF5CxzBkBeNmkpC5gFWVblhJepLt62NxpAZLV07L13L
A+sXkZlD8XXiT+BnR1knz0nSsCGhEuM4hHLJ4lQ/6p2NogbeYAZypseKaf+Umw+3
pl4qFcx5ippoEVhr4IDBD5VUW0L6H5d1TND75ODr0Nl4Dw79Q0zzrCwLSACdIMG7
bFnDRomWCc4Oz2FYU7WW8c+aCBkQlExxReMf1rDizGL4DUtsi2HOhFCXVuerdgrf
2jZ7k7F3JxMBJUa4WKd0ixeMf8d6tvDoYghk/5WElaGF6IFn4kQRSrUR5vvxh0X9
QRWYLCHE5c5PmwwPFgh7uAzm/bbHiA1R5kwijxcSMtWj3QZN/etTgc2MVs9l+YAY
xFwyKz1uxfUU8EKQmD2/reoK3T4n3uYhb+1mvFGB+bXkRP9wsaEoko8f0OlDEVLE
XOA7OYiM9WsEhjrjOFPnTRiqaDBAffyNeQQmP0llUnFMsATaGS+omuVBtrdhdabT
w+HhRU4vo91GihNrLNCXwk27CDt0qBilSxoJr/YkZhAjUPlbQitOoD2Ofwgvld7c
8xsmqsvGMYCx++cKo5SDqZ4KCHtVhySzllREXz7rUzOcSFmJCLUpdjKUS9RrYnW/
60OpZcJan3Cvx/MKi42ccZSKyOQLmOOO3vWOGV4gfKtA0PDlC1Xw5keNrXToakva
lROHTXCFTeFyNt4KUCrbb22hYoVaFKduMY4PazZpVz7suFQLN2/aTIZoX6cGUAkr
E8tthlRtjZBPG0kjIMSj8/kGZ05DIQgObLyWmiTUX6b/9sCteRbASGCweHmhctVq
4pbPRlvVJs61PstdN/aKKGk0rSaimRSlyqNrd4GUiPmEGgv3KaVDHyrTp6YPaXS3
QXanwTz6beRbllv5jV7y9vMjRWqkyE2CCu2qCOGT60ymQQcKgUX/oC/M9NUhO/kC
XDEN4V+eTwqzIC35boCwveVqYGPryCsr3jOmgl3HPwKYEXKFMsO9ZvG/8JvvgNd4
9ow4f5jmaP4Y2xrZJJ5EId+NnsqpHq6r6iRwuiMkLMHac6Ci8ztpWYEWde91n6+e
p5F6Sfb0we+e+rT0Xcd/0uBA+olxinrTAA4hR6i5eGaZrXXTzQx3TA18fqEngB1s
O5A7trVrMK2QxjCvU8cVWH/TGMt8PTDROgQ7g/pvMaQXcf1Mv8NDvfUAnyrSvTWI
ENbzcAn9u9oN3EdSfkyh6f5R0riT8z1U7x6lX3nLNFsRRd2HCKqL6tz0SE6Oj2ZX
NLc9moZRQZQePEQYgsfVnValVzRJil2sgOYTEV9fWd/AjBsYxC+wSZdT8WpPk336
gRMijyX8V08PABCCUcUVwXVBSJ+KMttsrTlnxlQFJEuUEkOmaUE8SwuL+4Bf31za
qA+ohNrfl/pf6cMKaic9FFfQpkboOpmiKKhzF2rVCvOkKtKxaz01hu1f1CGfG87N
uXo/I0HQ9Y1brIOV+dev4iDXEuX11Xb2VhSr3tLGsVnTaGb5D0NVm0qjSX7bVtLz
v30m9jatH9CEDqoYUy35SiGxfMo5aV8xoa15C/WVntyTW2EZREGASXFwsfDbCcVq
9q6txHNUVrMTAUWUPoHInaEzkrBMyXAUJ9XgRSVOKbX7F/mYDgJ1LZ6yLFfxzWJi
amppPrni+CK3BC3r+fLAHCaVSyz3SXtBzTZbROoSY/zN/+s+mhbH2UVwB+YWrS7U
d86BLeLlBZ1o8tqva6kBSbgaj/oDyDoG/WooJLJgCjh2IXIInXkDGS/16sApfRX7
jsGC5vVHGlTo1c4hZQ3sQVcf4aiQ4Gtw/Ibt01ToGyymCH5jKjiK3ghvhDGu8Xv5
Evc20kzB93BrmyqJrkcqISnrHWuDig69nkXkRviNryBvxvrQ0V45nNCIHfhAAmZI
XOEpqE1jF4OrP9J1JTsYwW85Ep2TfMwFrA2jq6AZXWYWxTJdCK5Na9XG7cyVNxQQ
LSHe8U92BFCMvPTyNmTsR3SnAGgO4NHuv9OYa5SparoZjFPgMwjNojM7XFoIVxyd
RYV7FnkhackQ0FR64Tb8XeW27xVgHHvi3sjOVUZtUcN40UBv3tOHFMe3pvNg9qRk
3JVxoDSRp9t9agF9OvjEbd5c60aADGo8bVc7tbPfQ1TqWiSWrq/zw40ty0T6C9vE
m0mcqBHkYvbh4pXR7BMqffs5cHxT7gGtsPCZ0b3xqaJxHVj3HoL7BovVraBIbur/
P38jd6lRbwu1zwUI7ZLgt7eV8Rhks92RjK88w+tXmIJi8qCmZvJpDPvjHK+xqliJ
LWzenEIIt+qUe7kUMziNC7JOn4Ve7Sk9TG2AkH5tXDOCsPxB53b1W4zH3Un5CwYv
ZcfG3L0WLuIJnrrdHHr+Jou3rEuGNIaq9RnH4eYmgkMSt9wdUmcE0S5QIFo2fZLU
kB4tHxoBAZaR+Spj6phENPGK9ljJN+aXePT/0Wp3zR7X+ny86BGsUHMSGp/r5q17
xNx6BrnJ7HBEtrJRGM4gmkgh3h/g2jvheSSLJ6IclrophlmfxUCbc75zPf3aQ1P3
HMn5bQZsgbSDWQmW8MM1RdsXA58v8URPyaVTaYXfL3aTAz7OlbQ+/C0AXEMKzAHl
K7OPYSV8xVjkhyaCpQQv31BCBitwKswBbLujreyX6bVz5nU1rJC1k3bvdc884wpS
3W8F0b33hElQJeJUwoy7xUrO1aE3fZGfznxQNRUbItPqmLm1NKr/ZrO8AvMBsBua
Q1ZuOjIX9yUriVDeitsXKLHhuBAfEKHGBk/PIybHPBf3vJfO3txxNnBcyk8ThWzE
AErOVo+EwS8yGiOmcSh1MqkzuEeddL04J+W6PDvi5xzjXq5hjzB58fs36u/qFIg4
dah2Qecm65OEVkauAaVeOjuLjNzLwIfHfSlSnIUOPkbHGetv6/CqF3nuAi7NmC+R
FwoZOwLrhd/rfT5LCqdTxRzpaWBNO8YPS2mPTcVz/UIscewqrTGx9lqOlCvBik4A
yM8ZDNmThyuEb0u+nrJyOEe+hMUmszSYtxh4fsPWz9Os9pax0x7Cb92gA1WzWs3J
46vt6xFpoZqS5ywMVHAq6Rtxmg7QZdIqJGGyKEkETOtEumJaRjAAAEQanI7/qLX8
A625s8Xd5r13QEuJMbbpx0JiGK3t8NdO94VruHzeSOkkpgmDZNsov0J4rXmfNn2F
3a9npULYn7zV4Ale2m16+tT4NfptFk0iNbksRcD+NxJ265pS3KTlWvQ7gxhRFZGj
DHjO7JwBG6iIcn47S4o2n0GxRH22CDX/wydmgTk+d8BJfpb0pEZB922q/QoKnVw+
KYY3MNURImQWDazhVZPUIqTZyWracuM8UpIqJMgY4Q//v57b8IzDUuxl3tJMbl3v
JAFCEpIqDFmGh9kkoXnC8ko2MxbmjTXMZf98FJbz4HA+CrvGNbs5Oee3tSgPgIBB
rHGWhGidVtOpxxcLNA+YSRjpruMmHrLChaxVadZ/JGKZrTOK/mUa1UZW1EemWkCW
t9GD/8U94BT90dOIf3V+iiSXcdW1GP/1M4eIReuVOKM0BbMxVKLQqKgpfcPk21ml
M+gmJRnTWpWeLYzhVuHK+wZGP3lbfyyr/XvsDU8MTlO4fIkNymXNiMGFG/k0MPyS
FaOqWie/DWBvnnrmRz/e74mMbJ05XlmYzVLJfPKfMDbnAAZrczN21lzW2p4xkkMQ
rLuoeKiPfIq+KuAVDqJZadZfGkjiX01fsjToffexCt4DnEgdy56cdmK7MatmSuT7
QndcQGd42ZyM5P5VJkaFACd6zclkmovBeIFjhYtwX115+v1P6DNq7tcsnpQ2AuMc
/KcjCfdCee7AriP2GPu/EtZkNjYcFQIIaV7q6kJA2ICkgwE49a4FMwufG1AIq6nZ
uTByYE7bbtWJp+gepT0l8AgNp80OEKWgz+sUwDFFz2a4uth1YGHgCO7fPrfJtBVe
rSQP9wPr7HrZGX4ZLdgkdJmo2EQoS/Fj5UI7AP/aQAT4+PHxwMOxNI5TSNrWzkIO
l2fg4i1+2uEPofywujFy0Tlh/AIZwUR8nqCTcw68ruWlL0HxasHzYCCA5Q/1z9fE
IU0X/KZVVLOdHEuivHPpAON+i4HeUEmCrKXM30b8zjrYiSaBb9elQMhb8Jjsuvk6
uWnETy1e5HFmxg8dqqhfU6P5waQpsBmQEFRUxgifF1yuf7B0yJLm9lSCTMVslXjg
iTbn5TA41Vgrawm3Ww6kWi6dyi5lc0ZDsvVtVnlT8H5hO/XvyZUruwvWh0iCrWSy
bmWIru8DfXY/1yEH2CqxuuTqOaiGYtzGQ60NNeDGU/Y0PTjzICoR/RdKD8F0p6xM
K73+aZRw0mfmJJmddF2IchUtwk4KNoAGNsILJx8psQ68lJoXHq1F59+R6K838O3S
maVTqCI53NZ/OugnUXagWV4y5moosP5sB3iRBKeLQXjrAFDS3ZUytQ3OFU8bD/cK
DawCY1mm7Wd2qXhbm6WH6y97TxJD561FT9AfXLm65b8dLb3SrbPuwJACJEjlAAX8
4bkQNiW83aYpVBDCAwFnw1PLOyiP5hwNqabEuVnNduUQfHmcdSwHgEabQwaTGLWW
t8Xlr0dGH0Mqd8NUQw6uWDbypCqgPimil47dH3ttWcvtpQ+fvgduzj3y2zoVDCja
npshRImgTG9Eq9fo4PW+BRXTgkhJIx8z8zGtakh2p2U3pFvXu90qOkxwlJYix6Eb
x5SLE+lQ0mmxep/Th1nqaBXuWgOpmcGBMURDEcZWIp+u5W7GoNOkkpNflKa03Sy0
0C1+HuXOJ38pZnXIvU5yWmGs2Uvl3jehmkvEMBT7VWllXm48i9roDNTLUDZlhIXD
hEeHlKtccYpa/pptMo+N+C0RDu+60FZGt6iQ80p/a3nfD4MIls1n6PryxPG7jE1z
q/K8vqX40mO9MfPBeieuiRHTcfeucURtBDcRFrhYWTj3JikHioNwKW0nD3kyc+o3
MSA+Gb4krxyKVtIteVgpzVApxBqPKS4L2jG5WlRhVA6LBaI2TZ9EF4QT2CkrYsDz
RRGiUb6Drj5OzCeG8pkhpqWN6zotb9t3G2YYF5ys/R9pM8eeVCTJpzYclqT90hZf
bPXIEZ4icLBAa5oTmiOj3Lyhp9OkhbAHhBhAa2kDWjcq1ukNVgk5g4u3vzM/y0cy
tQJgrrzbziJpcUAx7m3XZNyAHbXeotwWsTFPExHbEmeUGDUta6JRsk3gCtkKArfW
klXeLd+jfkqAiJ/iqPmJm0XXeW3AIUXryJH+p7ZDtKS3Nxr/D3lJcTehXxjvAB5q
tk3yfm/NZFi7zdej0rClsrT6846rxDMZeFiXbj3Xrpwrkh4OSYNqQ1YyVn2RyQeN
q6DqqbRs5QQtoobmBgJJp+o7m76jXB2hKC3k8EA8zWPpz9qFTTwp06lO7rNNCUu4
5hyc0SWXaQnhD6EmLOfngHWKNjknrvx3uSIxUo76wpFOisxvGKc1iRZVFFrTCjiN
GBcVpFJ2NnLpj4OpXdoqVwvbFtdx+pIMCp9SP8DOIxR8SXAnkfEllt0PrRBZgSN2
p+k1HOtH5Scbx6nsVlNbM/Fonhg3rNLnf6fTt3cq6yDeUlOwSVVyqzzh2jVqWhVo
zzvwkjpmdQlgHAa3X45a+qHnkojkPT3Rt6t14IYp6l53H0FkuKmCEn1XxiRb72xs
YR8KmGGJ/CTlDJ99T4QcC+VV7qvXGdPue+xK8QPc2cxpzA+jS4O7KIOGqDzHOYC+
gcDuUlWeHDoMKhkopDXqAZNByG3icEklW4U/2WJjR8elULRDfX8G+0HYL1mmnLAh
ii+nEcwQYOPG3gqu1KAaranYQdASH8VsVffeae52/F60mvblOIdnccmdv0e0YfBk
3lqRtLMmn55ZSBGwemWayHKYphbsPIuMmZUw5ud3cjAQ1tS/yiHrUwbsKFT2Jh4M
bj9Dh7LaiFz5eGdbU4PuXn4FoQrnNJ/XIxfbW9ulRrgazCLARllzX85WWMSYUJq9
rdMj5Op7sZ9uXu/0hj+rm4d8yjrPwSC+g2YSLgjpvWvuTZONJSgIazdhmIdGODda
YvyO6Q7qRYuChLaYl/9a8Uvx9vL8YmVGlYXvfq8DPxN1wMzFQlzs2waC/syE4qzw
j5wPl1RqoNXZIVsra7Nrjgh6V2zPOGt/LQN+S/iFnYltwvOtGcwYgEfkyXlIhqL4
QpXNauJvYOi5SpKl/XWZImnHVmZQikqMXSp4T0bVe4Q+DeV/tT0rzeNc1Tj5uS19
pAeKJ0jyAmFSYMOdukHilAS4LSYh2S9/rrMyHZEy+eD1pnqfhk5FKUJrRM8NvI1d
dgHVVC+NnIEqEN8dtmM66/qlz+vh1KHFWHJifmUveGNvPVdNQ8tNsO06ojinCV5V
gle7y08W1J1Glv3bnCaBrr2rv6nYvg53wy92IOO91bNC7+2x90mGm3vDEYKR6kUl
W/O2l9tuo9hqrohxDTbPmlFjYLBYYoM0XmBLb4/HoM3GlvYuLZFWw1ZPxl4Qz+J/
PEV/SfmrtOdhjuaMEU9OoqiLgdVrGIGxelY1meg3px++vqfxUTNc7fxOEmKoSko4
8TdwTdtl7i5SFqYoyOOKvuOR6VcnNvXlmqqCU1hhro4fumauH0oYJEPIBlW9LwBz
tTpDVFp3YKbRNkZJq4+q+Dj6c3HUgK1FxyAVfFjR8R6bWY673eJk4+X9fXX9aaYN
UHSrwyhJG4umm3/OMabZtyr1YzLzgUN2B2CzXqhDpMRxoroIzxqTKHWwJIYvB4kq
SDT2eT0RVSpW6x1YrSAgs6QnffiRbvYKh7l/RWt+xifC6iYzBC/DL1vZeMTf5ZkN
yQ3yvogdBPFl7WuDLa7v5t6fTFb4dQnAzE6WtpR31tcg+0rNNS3am7ynFAatOyZv
S+n9mS2gaAONRtGBvI/kI4MhsIxh1aqv62izKro14oVbuJ2F3K9Fp+37wb6+gB84
zGTV7isruerK6JIbCfEKDtCDV6iAqmTKWnnjfTzyCIosZFGPW2EGbzp+f+tZ4Nxh
tMhVa6nRbR/+hMBU20LuIYyaC4HxG4TqcIRkyPc3PPP51VblYu0BfM2o3r1xJuoq
ECIjw1P6XMbpFh0L/BSn8H20PlEnOdYE0e49LtfX7MTxfYeOlLq2iMtL/ohsECF6
9vY0VpgjbEYNymwGWu933DUKPdIqkBSauo0JyxmcxRq01fvg2kMnvOYKvkqbE7s4
yGXdpIv7K6UDKdpOEdSUbLQtAzse86+17BtgVsrgFCWTktfj+/hr39tdc0xn0QA3
/zwFGzuDeKmZySTHV9PEEAn4NsPrLtZAYt77LtcNhq5dqfM8tjIDyH52yycylsrB
iYmHVRl9sOMNE9+f2VsFl4BnoEj7WnbwpPBF13TdJN2OUolQZMAgY9a7AL0zjssZ
EZgcmw+BosGgBn9VQ7lONjy8cBL2sipsV2/lyIvMaxWD/nO4w/BuxuMkpYebWPwB
uYBQig78FanSAxTj1NYrqBg/LvnZXTDhpnVeMER9k9V6HJdHtX+t1U9wU7YQcnoi
XuMZ3K01GEjr4bUXHDfhy5JZjW0qWBpGPYY+9jbYzofDInHQnbvb8b4tNpqYtKNz
TdxPcaZdgpmEQkbBhPWNz7OTuoazftKd6UE2592iru7dKFaL0f7T+/ek1U8xBnUs
xOuLnncmnGocZ0zNNbP2goYsd50w1m13InHZjkpOo/S8hSHUH6nTyK7SuhcZWHr5
aljNcg6eOnS+W7327w+6078NOgEnan21qvA3CYllq8ZrJ/Vd4OBlNyHcctC0lPim
anfxR+vgPCYZ2zdpKUycBLc+OnYZ4PkSg78wZk5U5O2PyMLPxReDN7l8OhsTfGjv
9iVeDctFUWyz6dGU/t5MHZe2t1GihZhaBSgFwlBz7yhqdAI5zq8pH4IOPQUZkVmS
vDhJOb0xliHuuK/WElJ6XGp6WNm++nWeTxsxD0IBFWY0Eh3rgr3q2gmcVSPJRC4m
b7StUzDJOcpUxG7F9MVk94o2+TevdsmjTz6klBQydXNS8bH1lUX38b1iHOUqLKwH
PwlP5g7r+WpMT0/9oIVgUsQOH7UsdOfP9VOxHpDA7BKndYf+QuhP3G3KfEpdbrLq
z+gE0ybw3NLpuNlZu51ljj5OIccajy7/3GcQjzeBaPCCCnb0WGTV/TBwBH0y4Z+Q
2HobXVltIB3NQtFuxK3lAr+2kTVZhdtd6FCTkVJ4i5XKK49DaEddUUQu6HA7bf0r
3RaQ1Z+fbDb8gfgu5vZ5aErCCrHD1bQw4eSiNtdbdwDex0AlYA87yNSDsZmoWoYA
4jFfN0T/jlUzEKmogMgYmgtOyvwbfciB/rqj1MigioVrmiRofbyz6yUz4uLUEVwo
4o+2XaVle1PrULoPuDcuWJZ6iwKRAukpWW68dnOhf1te3RVIW4pP5ujiV6NzhLel
dkW5BbaUOC+l9vDVh+q3v8Z322wKJmDPCI7IaNcEkMuW47szEzPqOSgthbO9i9cs
ofQTtV6baAJnnPK22EvR0KIYAsKFJ8epVOTyN26866Abxih/rYEy+AifvullzzHk
iuLiXC2o8awopWFaOso+KE56L7pWwC+MGN20ssOdNjmyClrRSCplMCXTI6xuGVlb
kYcjQFL59fQxTWw5vqQpGkXfvhG5o60e6reyx02nomgjxbXudfAyTRIqp0Bp+pYb
BgUYGg14lR4hFFW/yTc743J8ra529SD9J8prqp8mSZF2HaPYH4Nteh12UFjyZs6p
8+Pe7zIPaAd+P68HduKkyun4rkLGNac690d4ENAuEgo2d82+VXwEZP7sRJoMx4x/
jJqk4RFKkOzzkzIrcrJxuopPlsnYq0YG6asd/bIsejA61DTlOBw64lA6aL4MGByp
Oo5uN+qNHvB0X8qy+sVj9/pwh8ggVODB3RluQsBDmKmQJi/Em53/TTftBGahvnY3
rRvtHRz2shm8Y5C2OrUC3OI1v17NeZgwDh6m8/bF2jAQYrPEp5E0wnMHFnKCyLRX
bqS6CMNQ5hjrI+twwV4QD8DodkOufsdZCtdPRZoKoXE1dhZCXwAfJWzFh1NzZvEl
WvGRqtaN0ooqZKxyEZD9yTHI5hNL9wsaLbBtAnkcAQSXSpP+8ORtG35U0I4tGC0a
a4XwFfHUL1FQfEi0ZPFY6LwEqzO++aoUwVtKzE3rZU7IEDb91PSGoMQcfpR4kJ0X
gnYOllSROEnnwzM8LPi6AJ8t/n2+2Yb4dVH+UcQ129XII2w1BzI3eyETRiJRI3ws
cEzunjHURJGX22kyWD9Nyxx7TYEBnApK7gvRfV+rasg6sBDVQVV7AgBYOBImtpX2
gufsZAGFjf93I2AiJzeVV7VbX0vgNzWRFxUqLw5Db0KrtlwhyEE5CObGoktXfZQs
oPLc3wRehdqNmtr6sgNQ/k3CFhEy4cO76eXGCieblcdk7GG/HZlhzlH96oyA0Tls
jFdtM6fUO0mdemBeuv4ui0HEmlv7vK6LyEjfNne19JxobLNS16gQVTiGB3cJbzn3
4lB7aeFh9wpdAGaJJ7Ca4djnSwWfYulkNfHmZaiaqiNJBolPqVEurZUDLM08uwyH
/o0Up3KacOZuT5+solnQ8HL+/IwhJkqNXa0nYFoO8qkfsL16opxWTGuDzi2qzPBQ
nQmqiFyzIzwYFfgB+XWXT27WgvuNFY0J6MB2s6FYDtXklPlsu6RYMAQGN03uat6s
MEHHOSM5IWbYFPobjrMBtMx/EOyRFVU/PPTS99rtuWuDxZ+CvVXMebWtxI7rjUL9
/f2XEQejB2aSdgUjyZliiiNCGDJPmifvUz3/eTaZUPo7gopy1jaf7bv1WV7VnlJh
j9WLMjjbHxjraFwsfi177ObLbUbxpoY1fq0YSsdvmqn/wYg+1rNTYwERk9M8hDBc
UwCptXyR/t1ss2vGGF3TfAEQ6UWi/sF/JXb3uAGpUlquoZcl80+244sK2etBh6Hu
2md+D1bcZuWbNV17gGrNGtxiNPbJyh4SBbQNP0qjtguEL3He1Aw/f2Co2gQI9rpC
EGlP5bySchi3C6AnYQo9dML+/jHjTCNEIFIVSORT+D43c6gLYn0LSYwLv1Z7xHG+
JNR0tkw0kIZdplR6uzFPsuMyFiXtX8egN1WER/Cw3UcXNOHV6Fksb6E/nfMiVQOT
USmAkdgxLrJYh9wYoFhyQhBDX4BMKhP7sS5qy9yQ6Z6MVvD11auw3xZ6VUJnuzbu
Zb2sHJ2hihHoSUREWrJVm79wxpDYjE4ImFjRRXCanvrN6+iDrw9PGfwr0kgysBdG
17HgYFzRwCQ5HbPp73nW2Dh6j5dvqcnWd0OyZWdmIxTsT8u/skNCrFYUxNkhVeNB
/JLFwISPXlAbM0ayu0aai1OewnMJ79xgJjlreLVDdArJTPeQqSt5esGAuLW3ivQn
GCuCEI/S/+vcyLXdPY4OYeJj2w0Tyx3LW3V5kQvaKC3RYQ/fHrNTjQ6EwGlvaDK2
aZaI09ovoWetvTKnBY3lp756IfFwuQYFRPOWMYoflzzC4RwvnWTW8czjaZQY6DG1
5ZSTFPa3SdkWkvGR7fHWzXsVgQv7c4li4cxcgH5C/3bexE6UKsjXyUtBNvZXK1wv
ahnVthpMZ0KBW+MUwCmELGFaEdx+q+Uzj+T4+WCQCauDszy2wPX7W4ZRzQOd0vuZ
MqAZ6DojG7PrRu6M0r/bWBwd0WezGGpWO58GjCPOeaItG6vjN5pGZdYYmAUmeCxK
mW4QRB+FdvnygTY/IrV2ucwMb/5BzN4VcxyNcDCh3AUiQd9hZXVrgv5km0/gdPtn
RzFDMYvRgq6PFhc9popXNVg/iKWHCpSak85xu4v2+G1rG7CYfv7H3UfO5l2UZIGB
1NMyw0ijUmLfxN5sC7y5V7ik09lsuZFQCR6Sjl9XcakE1FLxk8c+ILNyGv9EIo8o
aQl58QgH383LITaCm3dlMo3Bz213i2PBOApJ4/QY9axe2uc5B9DEBvY5N2hmogKU
dJDs3BRY5PG5dChaivRfM7O98cYLX3roLsZQnSnXKDHxLKZMq6xsDzD7WrpjVMj6
X74okLnIzQ/BDePMmz0fMJH5C5SGtUXYGZg6kxxol2pVEfsmT+VDquld6rBgUazL
TbsKaPz4II130phqxfXX1wBkxACnhEulPvMWCjW0BjemwFLrESXYLNlOeTm8/gQs
RYZAcv8kkpP1ihX+nJGFIq4lgdPF3AeiY8gXhLS3F++PZzCbuRao7MfBcwYrAI2x
RrkNXyJ3ilLu2e65Sk2vEIPJXICW4/mF4gdYjI6h2yaZu/L85kgjGGSKTHzkeb2i
qD5jClP8S/LLt+u0mHWg4QULiVX+90StWwGq0q2oSUR9IXZ1X7//K4MKyNF1bRPA
woAuTT9BB81RTU51iejviEXUHo7qrAgxPUFSr5YBA/+UlomUqHvYjmgKcngo0hfz
eFg5vd9X+R/4Gxnk7PWsIAOy4q56tRyEg4E6JYRi4lHxrtp/iPKwgwcHQ8YjdyZS
yfiPQQRHl9jhD6gBvJs+dbxDk90Q4ty2sJEGJ4UkxNzNkp636fOQI8jUgrezKw+0
90KuuLtQR9kfIkjzFJQdIoQ6qeobgcXlvf6c2A2YzzUZm24woVh7PIl/SncnR5rc
RJ1I0P16HrxzlFiYvQO3XWJpEPVh025JEtX5636BK3jue9ok/zursOGSQEqfDfid
LsxGQDALU9wI8OHZVMsreeydD05WQWjEc7eSuD9VXj8zwWTWWxRl7/N5cZf8c7Fe
iFIZSz9+VbOiEQiGwGT7AcF1A+IVh1Nz11ejPuIc656V2+aOSQi+KZzhRsjPD8mt
12lwyLb4Ly5JO9K7XUpvXMTAyweRzOfS/Tq7hKGWpqaxfkVNlP15YBbZdQgmp7yp
vDAqOOwkF/+nA3poaOkfJDAUi/5vqiZkMfLwLB+hY8hpcwFShs4Vo9pscsJ8H9J6
aVUwqyL1/GmQRVZP43xiW6+N9pjYzQTZzOmskaDzN7+x6UwkAg7Cx3L96Yb7MJyW
GNOTr2RHYb304P+kxJMqEUK3AwHEiqHHH6A1N/7xTclQeMU4XIrIo9DSnBmEEjTx
jnzLDncMyAPJWwGq9cU0J6Ex4We/5mgaBE6YuY5bCeGRFdo2AdcUzXmKS1co31AI
E/pW5eDAFb4ZAmKQq8cM5vZz3IAoZtY6pzsvIexX75s0eQ9+wjqZRvIbccRs/EYf
4V3c5U1WyHIcjrofPyiyRUYrpAbAnku8vaEhvHqZXQsbOdGuKD16iPrYV8fH5Tjl
IMT71wWydqcAxquXCDX8qlBIujWxo2Sv5rb8yaqA2x/Ig1NmzSCEgS4nu85/Rojs
Fs/ozIjG0ILdCUHHO9x6LmtHryL88dDyLKFUyod1FMcQVFBKe1Ol4+7pUWE5jEx5
YBnxvvX2QJW2lo3/WsE/PGppIjyuQ8xUrf0dPeFW4t82llqRPzkcCkTTJdiY+2q8
uBrIqll8JlfM1ysgjeFhbkYrJ2S0Ry4olk4c+ZVJ12evokiLnHZLwbhXXKeySXG7
RgCeRPrdx0/UlWw6yJ//rgRTHzqEFbPzYpP8qIWt/DS7mYnSVqGNLLTje/ED6unP
Up/EXK2ewyG+xSpzLaKREplw533tj/vKkx2G1fORDNRpBLYgqykvrDwl3ASv4ig7
13ptPskJvj8t2eyqpHu1OyLr0iI3wQAqUGV6P6E55vHY40VPLjXKb4N6RfpyMqnv
PNfkmZPzTVDBLEEG0xFjUqJO18TI+2AZ90cGjlYDSZl9y5V3ThP9/iXy/q8Vzb7w
XSsCA3iOE3yAUDG4rX7EZjdzTdUodNnsnRNQndNs6dkV+3+Azmudt5CefHMlsBIR
Uq/ffJi3JkZQbJyiNE2kmPgL6BJyFDq7IvAhHdh5Caq76Tp9QyLOlUZdOcon8aWv
iIRhlrRywClAiUKBM4XJFj5Jn2yM8pP9elpdGIfNM9kkMDLyVDF5mVuSSu91S9dv
Ll2Q/AmYZWhGqgt1vX3wVblxgYty4FTN0D7XZbrkihmy8JnuX5+jRtJNl9FZE70O
Hx0Ayjb4teDqa9KuofoNs/YtK7WsuUZwFp+aZ/BL9au/pEHZNC3YxsfhZEhgwU2n
g50kte/NmKgkantOPObpJ2kDtNpViJKN/S9xUkxpPqiR3ljkZZfGowHHJy2ccj6H
eVDmOpQrAKh1LDD9OR6uVWvMOg0ZgLUv3ji+VuGv2SjiWcagi3t068UhEHAJr9xW
teJ1ei8NlMJyhk0MjYh9ViRTsmmD0GDkU0hsKhXobuA6w7wOtHSaACOzwoJi/pmu
76RQxhyhax2h3dFpi089vVXmOcQuuMCi5R0FLyXJ0cO2qOeFQM3ssUVJu1weOwKj
IDejKNWk/ZfnZc0ljtdKf1vlbSkBNQxVQZezxKp5P3Hxldzeo/VYYbE7YcT0xlez
nTEL8kM60K2UxE57TEKc4GXfa63Xmq4/g2wOl2md++cHYp8Wu9GVONqrB0Kc1J+h
LGValfzc+foUKmy6clL4Z1FnWuPu9nuoX2HaLs1EzIyTypETc8PzUatqBBqUqFsV
orLB5ZtS7qxCRir9EHMqyW9U3WkeZFGm0n/rdacsBlwkBgNTAVhZBxJwOmphacpn
cXMfoYmjXDSu8MOjxqxWS3W5sk3Hr14yRkWv0Q7F6RgBa4AhPAdHjAbEWz5uhIg+
nM2L1VPdOR1RHIg7rDCn5F2rPSQcbAjlGp+OdjTlR3P7ogssFX84DVRuqdRzhlXB
fT5OkEjwd7VGEQMcP/pvN8dF8gp6QaEMmzWpmNoxvF0ys25lkkAAX/ekqZ4A7A1t
ZE036xNXwOjw6wBeYB6HI/uaPin3tk4tK/iL5AIJ0qUgiQOdbpj6h4VC/gKUUnsV
wcb9Ln3CIsstPfiX0ZTGSY1hZkrWnLlf5174dWSYxPlZXaaL68nj9pyiee40IivV
VJndHUTfiVQduYHBYxLPgvQUtTVqOuDtiLdl+l1VzE1KE5lppdtnoLDJxxxwKFom
BarIXCXr2T1ZZqc/tCbqEPRnMFY0WzlItTfS3VjxncM4qRq5XPCNjPFT30ydI4jj
NVNYZscwW9BMYSgtLwq4bsrF0Iwsd4xDZsHZbxz9mMXoxSIxVXwAO19DdjuKnyc9
gccABy+wNCkJj1IZb+RpJUuVE2IJpwGCf8cy4EtM7rV5H6xn0it6RZy35zchBKsM
zQe4faQ6sNMCc5ZNx8Itsr+kolkGX7X09UfFNYY7CeMsfjrPJ+EKqfGqEH/m5opz
0eSvSONmrj3RBGoosaqGkmkc0h0a5ZzFnWuzi3LYd2XxAxLh8unaWUVTvYca4YGO
7kGF/qwcv62RxBNr02CnGsplYGd973MLiBHwU9MIwwvFEF7YJGdufgxWU9Kl+YbL
oZJnaX8K/wVWUHpgg0jyiCFUTBA62WsbORFuqAVD+dJ4tKzM0oP/zO9V6H1Zl2KC
IkIp6tT76VO+vuH62sOs+PsTBraMYbfaSsQkY/KSEmxVuv6xkXzYdq279smUPlsD
GDto1iAECKjtUbsGVqSyUyfKjVRC+fAQBtx5x7Q2ROlXSjD7XCKXiPBv69tyATYh
mINalbJHAiQ1Y1oUNkeGJFwX8qYQxKeyMdlKfEf4vX4vEaly1BZxsYYtY3RORqkG
BjlGoikRF38wk4vdQa7C5lQHiR/aFWzgHfZfi15DpeCATMEAn+d0/MOGu0V9935l
Ckqbn3wiHC/LH3pxx2PVL+dBO1Ubg22OC9K/3GUL0Jt1F1f/pQk07RJ7ow+Epqrg
AkcrlQL9Zye/HyJw5WK8uPPk3/8fW4WC5KsTLOys0lx2DZXBqG8aY0yr5fuLGeRF
VJMbyDUtU5yFHAy0/F4Yb6NWr8hikXMRJ6uLsdqYnrYQvEamhf5JdorXprYHgZlq
ZF/cx0DnODGCN6YwzLzW6pPaRKg+9JD13/tGGimS5LB8qlCrm6vLGWk2LFwMQeUt
osLR6TYONQMmLNNHiXk8PlaOv4A4tfMz5zDG7Jk8X2+aa9Nru+VTKP44UZHD2t1t
JlnF3Ctg5E/uhQFCZLaDyndhvia7VZwRFN35zjonKtaxwQllM1vHiwbWZIqvZ4qQ
RK26kF0ELzPWkO2/vXOPTaG3o9R0Z/EQM3K7v4ZKoLb9LlZrfKrfe8tW7tZx1XnA
G+m1UwxyshGqF3grNoDX9cinU+AK7AuAfCDtnK5jN1SyG9RocwoNfyUMrmUvfR7q
HwCGdni8O60nOw39XMkWOhONa+4bs0OFX7eN79mY1uV9vmax10+l895oa3PjFQeh
AJPco0hos782bjg7ee8aJzlOZnD7duepKWIDZ9LR0oq1D6lRgHuD8w5X3lJOhhvq
Rcwyk0D5ObMe470OSr4jzufAJMCekoHKNTKm29A7I1UgSqnliolCYxUP6L0PXMXz
sHVmlFhPn2c2Vf/WhX8UGjFlhi8jSAJrOhP+N/HaxjAVxBocT2bN0VkchDJjrzDJ
yRjPzprpkZJAKPKW6mBX0c+pO3mHYN/kOYuN9WQ8Z41HzezzRXPMP348N2QHfO3o
qtEq6ItpQinP8H1fg0TRBR6GI/4GlhPruwBAmzs2akg3RRzvozV37apJXNBs/7M2
KGUc5x64t9R9con+FcBjSQaBTNgAS/VA+UHwGXqNlNNgu100tUq2gESoMvw+Q3yk
WfHs+IqOC39VPfFCT14dNc2cIcb8CfSkMDzlSWjUtmPPNZ+79kR4eqq9+IVQ/MOO
DuFsQpd5elzBrdCRna+ePDWcuNrLs+p18F7rL7AoettILmH+gEuW+iCje+X06AVt
qAl6F3TJDTGYxIaPbbIexvnDsLLgin/JCiPOkQOtiZTkgZl9VVXUNfe34bWqXWTV
VvFc9jnGKjFQTaoNlkpu1Qcgbj6DqvNdOObZJ/jYI8FpNOBWUtFmmDIEu502LlgN
8CaZ+zRifDyn74KsclGQzKoSuR2dH3VMbg8xyKiG3YCjUtLiGjA0YvE1NT2EygQ3
NLoxpFlLS3iStjZ6xAO8S1Y9QuASPkhO8SRBK0NyWZXHSmh2p16qfP67ArbfOU5H
MdIN8iy2pCI4ijj32tioJlqFOTXv4s2YVkaeoSr+ygp1mvbwtw6Jf8BHz4IBcY3e
L3ZTA8k26j3TrduflspJ4HPMrMcGqrxf252JbXgfCAgZxvQGtagpWV2V99oUU0SD
awqyRK4d2MO9MCCthUBmksVTh/Lo3KPukAc2Zkpv/Fn1ALNgknSIKyoyOrf4WaSn
T4ulJ5H/Bfg7ionq2lVSwpEFRTCKTPqx96EqKHlJh4GMcsxY7GkAZn++TLPxKys6
Ms5qbzzDcW2tGftXV65FdrWWLHGb06k+tm2iJRDPqXlkXzYvgGaS3I9knJEW5bPw
NU0VflQjpjNeFBCtKsJscmW6Da/FMn81ciiGRR1SUnq9O98/h1LvVn59FiH23tD7
CdBihXIWFObe6BbdwnwHxDlT8yYPYm3hBb1uKzCr0dMfnCCqgaOxG/uHKQbHzKH5
NwMYbMA48lmSivhwby8eUPiGm0t6VvhS0NSqtXqiRiXFLxx4532ydtkzJl4GzqKt
s2zZ3deIwdbKL23W1LU2dTYDdiompLU5B3McoZjHfnsgyz6/aftfTDUKAiYar5CJ
ggeSx0KdZ1RiJBREy5D4K9kZwsTXj/9Fsg5IGsIK94kpTpj6mrYXew48xD/j/j/D
/IrCq4m337ItKtgCPjz9lR1aSTvs/1lkWFzMnHJRiNvvO+NjCoJ5CxeszjKDyLc2
W3J0wSECsig2oBBQmaIN58B6GGEkJuXkVNTXw8sRBEkLBchn3+n5ZoxjeFy4cvTe
NWCms06RrhNRxSds0CP+JuiwWasIGQFLRbFxd83zExfxfOIJX1e6fuoUXC+Gvjtp
d+HycldKqv9GUzxDi+JUbIuX0RcMdHaxWl+W5xxpn7IkXdKquVpzvnEIOqD3OvoT
2urZW2/Lc1HtHvuc9Wx3j3xa5dX/0vsMH7TssES+O+PU+37F7jJTk4COEPqKkj/H
5apy+PhBsAlltvJ9ULdSIm9rBKGsBL/WvzdybGV9auzy88UNJ1wtmQOQk13LVy74
ufyK5O3wSkkQacmysnJE31QkWdHuWcQUJqnKymRFqM8DEGZoqLhkVWfPXzKKKGK9
RHgo/GlSpW0O8xE+9L2QOCjh9OoGIYAiEhlov1K7FDjsAjrvS0b4JWimIFf4LeKM
K7YxOCvIdn2pTVt4YKOzqa7odL7M9Jf8r/K2hIXki7y+bnmcFlpdbU7h68qnaqzE
vTVz1pWGlTY+2x+V4hE6Jkio4jrX+RYet/9KmVlCDQgxhZqf9opzbOSlVXvxF0bZ
o6yAEYeIHCxYcyiHzUE9kje+9UoUZ5ss2WuDBMRQKpyU66A6OIAioBpLBU/NIHKw
hggKZNDkUwdbz6CFMTsD/cTQyDwfCNGlKCjToZ915Ix8YjBUbPfq0ILXcVnm1YRT
HexefZYOLpVgFtX20Pz+mc/fufQC82op0ALFoyg0unamujUFxkvgOCrw2OmT3of1
43qwFVHtr91fSIZe8pusmftgbDFCCvp021taGg4bEDcqRf1vIdNhf7ZPTf7buW1W
iIsIQkSVs27gxFP98bDIevDGXzVSpwktZrfUtaUjmMwdchtJwTwxDukWOqoRvMFS
IQQ+eP756+ZAlTtmmOnJaFTQI3V5lLzPN6vRCndJYi8smnjUDPE1j5O2tVEC0RBG
blIg5es+ZRJqdnQWll5dlOnnr1k7B8q6bjj8vWaqOFnTcMJcFZ0dbY+ARQT/v/N9
5KgdIaZ9Wuua5nLTQ6vP0g5aoJEyVSs6SnPS2yIDkU6z5iMyTnHJA6/36NVkynwE
SqipANwipWuItXRcHZVhOtshmIUEGEW2nTvI9rkeAuCUNNV2bztcqS2UiCiOyrao
PDulEXCSMHpmW3vIEH22XqgyxTPRVcbyakbPN25e8EPikP96KtJbfincsfMWV3xO
B2vNEXbddXWrNL4zNHMS1TI9HCnaQ5xHOendP+VVL1UDV4Xe0TQviEQ6zs60pPaJ
addU6xcLqvxtDOlVVEr9bePxq232+xEk27iY31/7Dr66Y/i2Wu82CHt4h2jm+heu
0d5eWoX0Y3F0J7pq8Slu/YA37o8IK0OhXz3EhPocHTxAGw9XrTF/5PiP1/z4xw82
dGmkXExdOVhNqwQDGxFwPeBDgM92X4MnuWeg4vbV4G/FThh1MULONZuQMxsQK0tc
IZx4OIe7+ulfIyoJPi03Nc8SruY83x86z896jRlntfB7JSRoWg6Nag07M7V4QpZN
VCAEN4PE2Y1N8n8AKMnu7Gljs8qmCV+mOorBv/4Lg/6KmStGUX0xdISYS5HaPc8l
i5KP9/HffKPrRZmPjNc8LdkDnC5YhpWOphZgZJv2gomVl5Vzf/gePvFZvuj9SQeg
A+i04FsNhzw+ZKWRPKFOgBxPUvQn1TT27t7zyauJzCRm+171UK41RbK6cEuub3Kl
ALboym9Xi3c/O0A2WSlxUrJSMWB5pKlMpZ5LHnCSSFdXSUDqVm7EGe3b5APnnbiy
nYtp4FyRe9Q7otIHAvVQIqiOo4b8MhiQyMCN5UmOMg5Sgyebz8ql2AEytyuNtOuf
gOMMqLQG3u8Hmb1mEsflcbk0RPZK/qNlXermoSfnbaJc7ompqJlMS/Y6JvYLYm1s
IUk6BSx4N5AmwoaR1R2bmHr1x2x6AlTonc72csdveIUC7gf7v9x0+RZ5aIjmzw77
FRRwWWDH5D1lvlayIBjDbOCnWie8tM8qfPWRfWfG7AsPF5KJ1jOjvqrRd0vwT1d6
Q+OtOdzszXjdQ2bx3o55sBO9OJMBd8EGlkicplph2jlG/tFAU0QJTJHzlwVEWp0D
0rQQqLx01fW4Gm30Db+wbHFVChvphgWSga6nNALT7oPxlfBMJn3RgT1Wjll5AFGz
f7iJFrol1keFgMv+stw3kmijE/6KJebosFy7Cr3xCR5QwXNemOXiF3znVlCs3ey4
ZDZwILUcHfS9RyAhRZidI9rU8Iyz65VinocTLiJbjrz3sJFV97cj9xapxhu8bsNp
S3z+VN8IymQdjIcewfAqKiPIqMBMGSuIBazfsR0C8xI4wip7XoRvmzPxDtrrSMNG
aV5nr93pKoEsoaARhLERVaDO4sULB3rtjYEvWyL2FSyVv7CXebvSNKTSeCVa9DYH
B8hKMujz0WatPBEES5RAsQ+QiE0bnNfrPOD6+3AW8qez/FsLQL1GVPWWMzw3QZQp
CCRFCgrG+15OnhZh0C3D9TuacJ5v76SNHWR1UFxe9VWWxpvstuf4PPpHiD2uUU6b
3hD6E4vqrE39q1hjsNmfSjPuhCwUgpNMtooZJCVkuiG8HMizKm/tVcDFH9EvkcSR
j26QptDlbAC4CX0EPQKX6zvhouFEWkGwrTOtjSn1UJDaCa6UN8YEi/aFTurnJ11/
okDa7Bp1BlvG+C9FVyfQb/GkZfsdhD0tYmRkbfrrYxzcTamhlHg/QFf82oseSjcP
ynYclDMXRkxj2FhJwjIIs3m5c7iI80RymS0BzPw2Uf806htb7njYmPMxZSZwJuCw
3p31l8WTybMZnBNLzLW1QIjYBnMaEneD+ZG5gsaPR1m3QKXr+jwmv5lJBAVFCMOi
jczEpQB0q8uO52QFSQ1XDShRTuAgzjedCgqSKi/4Nk8ohuNtZv4UuwIzLgqHoNJy
i0xn/QmwPxjhURcQ1JiS5GTjEK8AXNp4mKC9fXmPx0ABq0w0YPRRAaOSWdUkNhlX
L1Mlbe4EZXwSzygJn+nbc2dDqgPdJHq9IcCBagGjlgNqMJ7/CWLjSe61M5adGOH/
fRaUH7vsF4PGeGcWDTZFz7NvkbJz3Eim3cag97AzZ1/5YmaxQLgEnuR2mJIDkH1a
R57o8e9VMkzTftk3MewuvZs7jQl5+VoVHFWQUJQ4JyNiiLsf/Wwn2GiFtZanBJRN
/glfsLM0i1v3lmvuoy5y6B3DVOtZUbq9CMn9wBaYD2eQOD3xq26hfLH6mgZDyCDL
mDc6mBNnhkdqy+UqKszc76X6+813+eIcI/URakFtjOc4Cnu6W1lix7kNzMfM6f15
m/QJelZA9phYqvLHh9Qc8clmx1EiVxmHuYIHcxmYhAahH3fI8SPrveihoHyHRxeA
XPRNBwAUUhdgTqzrxkuNtz6S08aWgAY0j80lBZs7HFYJ0m9qxbW3OnYKIUW9qflz
GCogZjFZxs8xY8e2814QRCj4FIRcu0oisR9sG3oGegtFllRjxyC60g3BBozBpNz0
uHTa4PJVxdl5U0bypOB91rshM1MjvUZN2XUpqc8ktCJ5ekw6aZvptgLwFQrd26zF
ZFKDAGeSNgvgYCyLa2F7pgfCW94Y2G4jLVGJhP9/Y0yOvLTvkMETUl9P4e5ybJYf
7dvAZKTPq0WcuN70+UDhIUiaob2SlrKpiHlzpgyLRpgvcVovHK4697ura25WLjgK
3+x9u2r1Cth7VUP/4t5OWv/xF22jEUe33oBoYimXFD+GObsTs0piVRVRcG8niKeU
ZcDMEAKiAGewsv2SB2brrRdw4UfRjs7sPUULKvtp6DDZfBB33J4PjAQNnohSobrj
UDlGfAKdHRPj7HbvoR3KCom/hx8M8NJxqXIas4G1iFRmYd95HVbeDDRO8GLVKkho
QB6fx19n2zdEkNhjx/c/KpKrKe/Ej2rj4QDlYxTfDxP8/aVXFG956yb9bSa47EXI
Ba7j2iFisxHgv0FeITfiaQSpW1W9+UiwGACJo0WR4jpI+PtKC3jl4KYlR47E9/Bt
S2svsCmyPCV2eHlX2Rx20t+vCsbHOoE21McJXExLtvl71IfOBEJbav9UkdNnDfgk
qCsmovD5zbeKQngOp532nq1ms9QrS5LnHO2IIc277gLwmkIZkK3gp4YKCCK6cnbx
Qe+u9J3tRRsp6z8SG0jRE0P8EHXX8v//uBY4crbk0AYf5gfoUnAMt7SpfPLuu2Jf
cg6kIS7gMCdO0vP0FLE5ngKwPVBAy9NXmgBjHb+/nx9WSx0Ng3RqLz7bXJ4G0qLC
55U8+n0ra+k9VXh6apQ1cVPrHsBQ+jxWQH4Dgy7iFzPz00Apx8Hyqr2CC3Jwd4yp
K2O4FTIIGagHqKzWGTSkFfu/1FNbirONPx5M9l5QNJjFyiWKMvNWMdQKpx+Z2fsa
/Ec081VdqbENXESqkA7L7L94lh3FWZMA/iVVM/muBxEt5fexpdn+k/nkqbBzPfAM
NYgO1mzUwdPkpgYbjZPusCok3LfKNrLBFiLccZukhHwpPnNaJhlDovWr+9UmTdan
f1CTwKNm8ZN1AuenKAzFy00cGqWe1QnTQ8R0jGvQMmH16aEr4f+mMV1OaWKWIiaB
p53Plg1QIMrYkg42Apkh/4KljQM9s7G6/dNCs+Y2mA+ihnG7JcrMiimynevUjyLo
MHW5KgUzCH5nL5JPiDPtv+W1Pn+f1nIx3S7OCFSjH3zqogfcdOQupV0qsOWRZQ2M
wuBLjEE4+K2dvWjvSJtQ4mu7epRT5/uI2w4rCWFh3/DmVrhkm+cn/Tj4xwVeAWEU
BE0trYrf/n/QDAhG4pp2NQyRBD2+UTCr0jnkhzKQhxgbKkgpSFWFEmBEFZu1u9vD
iOYxKUaa6Bt9sSILI6aTU0fuIPLUXmCP4lSqHiL3k1JyRpdHduvW6lkLCe4n0OQa
Csj1BCKmeebyzFk69c9UqiZzeBywp/vTkpTTxDqWg0K2GxbHymSz79IhCLP7KpSF
cQ3bbApk3ninNOumZlztfTeeMgof+qLRTn9Fom9tZriYBokk0r5IEh3yy2PeP1Y5
9S+V/X6p27lq3AqEQH0kyFuSxXBuCTjO5Y6IBgaoD2htkDHvFMVGtYVXshmnezJO
rqmqg9NmiN5h6/G/txcSSs8Z0vtbyBziPDHBnkFfogYXI3Okk5eaJH6jivUj4UbH
UWTLWRnQFEb8v47vbksFgQ5yOyEhxSPpJk1Qoh7AS6c2ED6z8idebaQFWmy/PIfM
aQgF7f6S57vnh+z/kGHWEq2l4YcTQFvX+OrId1aUyoOTQBukaNGSbLI0yzf/Ym5y
XI9oxjtva/WRCmbTWxvApqitQb1LIMu4fd3jhfYvrYzftTiCWoiQ3+ushjjzC5U0
ItU8uVxM6xCD3hTRAUpHVSDsZHJqxQ7fIu2lZO/oEr+J4fTyv08iQ23GPWmbTLmP
4rfsrnP++0nLnTtyU3cCoyO3HouW5ME3YLsZoIrcHdT4rMjWZSkgXz5l/Yz5hYVd
6yHFnAl+tp5OpHo8LNq4T67zmmdB+iydpjonbA7vM0oHRlym+iJLNnPDkkXVE5dR
ihta+CmRMY+QSAIW8B/NFR1cQRmLny8TGyGuT1fLHbIbUMdlE+69j8lARGyxSNIz
nfYqewfGfeYPH/STmNamrrSpfdJax/HL0aEyY04vSc6BGmb0aGcjcp91XwXmy8/q
n7xClfIimNKDNybmFZ/vR44SEIuwnoGxNCOvqtotmyLlU77M6giJAnWWkS7TpEwV
KiyzevMA0DfQbbgJAKOLCx5P2ONSo3oyBOdYRJbJukhsqL4F52oC/hEByxdg44qG
vfTZ5ymQFd/quqARkAb3KLocFgsION555kq4S0y3BINi4QN44pvAWwXfgjxr9Nr4
jjNUodD8yf8TuCXdJlfJVmjZ1Gm5KzoO8NDk99zLbUKGfiJCm2YBzEl/daAFqO3/
zWR9KljpzbmihZEwk9QXeXiB3PI1labcbRwQBIcq3KQHTqWlXSOsE7K+sSmoVaAF
WB0uMqEMupnbgu1YZMUBSWue3TjE8QyqxCz7gIHk1mfoeXR1gPjJCwzBcif7Eihi
/nBuZy5hQYGihAaKp3IDMr2iNgLD7fdQKXO6YOZ4ORrNC0F2H0BM8S5Ht1+NLx4P
3Z3dS45neHQN1+jAoZ3bWyzvu/kuQ1bRDawhxzxQSdbkj4wylxMXCLwrYnyLsurs
t2wyIvJgGN2SJkrTJzbSofEr8GePBmGv+rENil6oPkTYgHzzsegxNtwKU/BE+j1E
IYg5KcroKj1MFp1NVhhTPg3N/I2uePMLHEbz1XZYy5U92rMMeKxM1oVlbcD3AiSS
BZfKXnvwJioyV7ICYe6kzW0lGGicU4M+RjWW/5iZ97G1VeN6aOjXxmXtzZ63Pupe
YCIA17MOP8a6Gyp8HCjk2FK38q5tb604sGhWkBl5w8Pt8cEDZ0yeR+7APXFnMpGb
edn/OfUPP76BFrDIrjQiWctCO3FJUanMH/odEBtKogyI2k2YtJ4wJXKMrFNQwCxA
EKRfwu5lL+7iaqHSb8mW3XtwE8SXiFclzenS5rBfctSSUa/JeeFwymeNXxGhgNn8
M3wGkGJkNx19m+/T4+ETZYqlt9y+XuDGh7UknxEwAchQ9uVgz4wchN7cYyrcgxpH
rh0Fl+s3ucA1wsUa+FAH5dJhSn9yqQ4V9k03xdTOW59DIWs9o/RM2sB9xn9Fhs1V
YuUn4jDrBVzKXCnl3xzt/dSyOnaARiqUC9ewMRjA6eKUdAlFZJC2pcKpymueLUwc
ZN6g3hPag6hIPtf/Hd6C6jeu4AwQyXxpKZb6zpLozFL+dmkJVPjw8fEmEfRXcVzC
K7T5SvLucmDYk6ryXS2dMPMGdEW9zlCm+K17j5eQANblA/s92CrJ2yCLATqQuv34
v9UoLBqh5HjMFb9cMWcOltTMafacEjWdarHlF/GhFOfXdZ0x3y98JfA/mEdhy7aV
TuLfsxEb1NVgihVEK5ZHkAocgWtsPiZx8zTR4fDT4NWUuduWEPWqk2DGj4G+mTd/
IN1jSz5Ydf9TG9k/GfDODxb72Dk9KqPAyLuKkvysejgzRTfotulNY4FR9Y4z6uej
OaqrqamXtxQ0Ydcp5AhE8INRSkrSla8ntlhSARG2pz4JveCPJXONoSP/biiuEj//
vGPrtvUNiC6pDriiALxn9P5MJd8rQ8/VEL9uQfD5xebad7GsvvE0HXAeqqOmhX71
izIUuOX/WPo2//GwXwjoxbbyz8uuZA+lRL1Pkj6ZwDbCVbDo91dvhiw6kEcAPTgA
BPMroWlDVTnPYnobaw02ZaXwvIoAba8ILTg2cj1Jk/dVPkjYkw3n1YbFGSgXdjH8
N2CgXq+mkOJO9eY6gv+JL6lPHOiO9hEZvBLeA+3BcR/vB1ukbteaV2nu0H2Z6U9b
J+7g5r2xLrEHMYcD5QdX+gybUloDldzP12I+Mc3Xwy229PLqIfYRS/hJjUui6+yx
l5JpgSXLspRz7y6oMoA8o/IrfSlFZDyGwF4eAlEl2EjGwTA97Zyp09dTAOzY7kh9
uUyWW574t8ghBwL4NqX6y5hweXd0as12ZE08/o8W0AyrofdGWfwN3CVpZb9cXplL
ucV8J+R9xnm1465btCrzQFeqOM/vIDVImW1gC/NPEdcju6cMbJTjAGIQoMqsSJt0
lsejTc0g5SX5wbW/M0ufgr/vxrDQqAz2DsJqLFEGgr3XZUW2NZca3Ph8PdJibNbh
M0jgR3lv4tr7l7j3+f5MZw==
`protect END_PROTECTED
