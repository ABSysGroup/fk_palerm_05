`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H1DkORSVVpEW61Rvv2neMu9jQOUHi7ue46lnXZR6AkaXYRZ9qSEx9Co8TcckmKjB
5gRl6pfcd/fFv8VkRRdIQAdOKPbsYTrH8LP4BOytSRYMGTqG6/ACBtrWYfCBZIlA
JtrE6/ZzdOTJ2EUveNT70I9cDXtzkRbuf9gBIjYNue1l6RcURfNE14+p0bfixVCj
WaBfqYcz2VEdWFkjj1cgseD9m8avOSzeFKQolnhyPWBm8DAL2M5Po+kklZ8hNDhH
4Apx+zC2FkOviNogD+YqtEybq1QCx+VZxXyNawSYyw2azeRKpzRAv1PmnLRjiA/K
oW3G2ej7xvUaCP/30hcW+PmVuxOtR2c8I+uiqOEEb2+VAcGaxG/fvn0KM29raKfB
zzwd1kCIBFYVTwAjYC8enoIdECTw0oQ6o915SXh41UDlbq15dUIDc6LlO+H1RYAF
C9tuyUwQq8pFLBpOQN/VsEz2RTD/R7Y5ZKyv5mug3rKbCLY6YyRmOtQUH0j86gh5
ohsZV8596L1M3dzmk3nRLmmzrSrTwScLUseok9BzXRP6rTKPh4t98CX5JbqOB9Ay
Rj8YAKEqeDYePL5KRjf9N9zNJGooIn21bioZ0QXUtazjI4ZgA/XLarOwaiyBFXDY
68soVP78vOf2edn4gyCpkkIgGs9mWntQIyPqVILxPPBvh5R890FDTlS6guoWaDfn
77fVlwdIJgjs72HW6vzEQPpNtbq9buOTmQGju/DWMKTnVBIFY68U8Mxq52V4SaIj
/C/XbhU9XkM0AlJTdHugh1EEJurYJxNp0FRr39R2DOj8ixnqKB4QumuV8HaUdYEC
UIBNziKWpskSjI+LgM6IuO9q/+WLu4LzC54nK6OHE1e9ZLsvR4U9qpzTXD9vEfgZ
6sBOT4n901LdHOrP/Oiyp85M9TYY1bPJ5qCW70C5jaicE5UCWRHvBMRrYf8DO4h4
HgsRRlthE1bqSvn46YovWrqE24HkFMKALtItGLEH4PwvwT63pMNwmPjq2B1Ri60G
4GXAToNjzEV/nklUTHB5ujEm4uzxk+pSOhGUjiFYODeSG8QkF69e6SC2DiUUrOVG
1N2pYlbfcaImZlXrBVHCZ8PTYWgHsNbmG2z/Z+lTM5tcVXc+X47uOFds4MTMsKMt
5xbLpyraQOhbNOXNX+eGdJfeSnhKcwdYx9bM0SKeTMTwwZ1XboJPyi5cIKKXdpGX
2IPZpn9FZOhW2VH7yQJJiUZU/PBcn/u3ecGbhWi+yYgA3+iDrA7DLg/pc3Mq8TIh
rr0dZ8aUGTnhFCtvK5oRC0sA2v0cDxzMT79kDj3Lg5NPU9I9JVwTilPZ1kLH6Sjo
EbiV6W/7MdK5jOXeaewb32bAmozHHKmWPIGNHNDdjhwrlpQabkFttWc4/Jj2n+yI
wehkp3f0AY5HM4+CPlrsp33UPfNzvuHUjXU+M5pDsYXAfLQarrbO8BYdVLfSDUtY
JrZhhFfvn+0JHsz2pj3ok5NsIq2Ypr4RLfYEzYxKgGVx04RSWcS9sYUVA7tMjds2
9Mr31zWEDUrJyuH7jttBjA088ga4xUc/nnirK/qVaXRpS/LLxSxJ5tkesAETefRb
K3yuPvZPqYS/1LLxWn4/bPx8jzjgdP7zNb6MVQn0S0BL1UuCRv9hILnG7XbH6cul
roPd9w2GZxfAgAuTsAzMcf7MGdYEnzqebpDa+VN0yYaPS37SkeXGmlmnU8W/MdgQ
K7FLymogZFvyQAG22+enuN2RZcNUN1uqvrCoBlb0x7g=
`protect END_PROTECTED
