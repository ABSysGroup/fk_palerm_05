`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hvbTfN55k9eV3UqRfSbuDz1tg/suGEDa8XyOW7L2x7EGgXOxRS/P0gguCWN+F6Wu
sXk2xmgzCnKx7XvmdJ3YgSQ3NVuNOacAWWq11BPKOgZI/bOrlkpSriLKMkr1/Jp8
BTxpW0u/7jNj629+DMJleSotkmKM0tF1efLWb23WX6yQAcBpd84i31XbYaANTkKs
rY/bkjRcdD7ZEjWp8/kYRG+U9x0zXxYuoZwfh8Km6fy2s5qfPvYT4ThcivGAV32F
TBrN3SfYfkQQ6ll12Vy2CU3s0fkqJu/DLkGH2j7hzIOXvV/9mGuOIBeE3N/pttk9
ObDwjrGW1ymahPuSpNAKEuOCyug02Ml645nn7ISozLtz/ewSOzyZ0alrLSZwNeso
+LL2eJdjlN+Neor0cCeHvnpr48HofXCFfz45IPLKxkpUi5DNQ9m4YnbF6VQXpYc0
ukgE2HSw+nODRAe+f9y5QB7nuiKjibgVCqR+8W6TjhlnWdBxCmU6o+6k3j47Pl6d
msdxFkYr+0JGFU7KQvaIpuFlkBS7E4nf7D6KzI7kZHYVUoRzz6Zn1HuREOmVhKAb
/+HbzswnQeA1eGYf9TH1IWcU+zVSCXmjJZoMNUCe7wObGssof+hz0mQG4XNk8tSI
47/vWu6A6Bzwt/eWzomkn/Hxiwm7/fi0HJ6BXHsQWx7/pHg8SfTpa6o6yCGyLhKk
tcJpOsh0jkwBuc3CgvfdF236GEZF1xmFal8AUmgdIeLp+kh3uO8flj7VC+BHzH1X
mJ4i7iUvuMDH8iGU1SaZASthbj/mORRcn3V6wFQflBxkDKYKY42NxMjYqepMjfJd
5/RzkV+hi3w+a2OH9f+TDYB5pPI2W8xFkG19KhlYuVaiNQi3RpVqCPkXn05lRbyj
gNLmNnPYYGdNmWgF30OfwbNY1uTVIu3/C3QxcQvVdFDPf2jMlK1yOQ1BRetmKnzs
T6jkI6N7HyXCCpnj5UoEnnghxbdAQ8lv8byCuOUBvapSoAMrQ4z9/cfW5P8fROyt
AGIxNSN2c7EaWXsn0CMckGSnYdVwvGSyKvsLkb+BC0xgK4D9AA2DZUWXIfJjx/wn
38Qz9tVibaCiFNh87pGcSFZ+soHNpxy2hviC0Kj5AveBzFoCcVL0xCj++ehIQVdz
Mji7Dph2k2yIMSppcSogAr6VQ904Zu02MVqiXcIqbtZ2HzTKf7HffAF10Hd2RJni
V5JCA+9GtKGBNi1PTlHSh9I6aCm1q5VrQ7QidIo+Ihv65LQ4ObijmViPp9tT75Ic
LCdrXDYeaZMUTqaM2RyOLdKIoxJ8FmpXgnhL+5IBTOG4+0T1OlU7CPkyr5KERxm6
sqA/LOU3HWmw3I+MhFEHSHFtroHfG7nlb49SIBkAoPmhpYzhwELKAJxP5gZ9568G
fHjn5iUD1vzUKsZccjvUb3kNVLDoyd61JH7k0CsvCdE=
`protect END_PROTECTED
