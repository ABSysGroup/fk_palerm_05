`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H5tyCPKF52bAnY4jjMp3goxALB4Pv1lNHagMqvI+oA/n9mmT+7kXUPj1tIlaSS4d
spLlfDGEn8w+zcaaGjOXkEQT/YtjznY1iR/815lgZaJOWGHnYZCpeW+fuZ0GaVLc
QbormJLxs2sBRLhgIV0Ukayo6X9N4PJk3KM6eK+Xt0in6p62Zrqu/na2JvJl/4pE
URA7Z8xwGiCiKAKgQ/l+hLfd8YdNm5UtUBuuQL2IJqc9oMtL2cPoVUjTdQixltHZ
HLCTme/LBd/hEmcnu3S4WLPQ/FL9+IuprZ0myT8aq6gGlvbuuok57hOuYwSgzIf7
kLvhXShBWU1NwxyZdg5sBg2HhoRxOBPwMU2ANaysqlfDj1ScaBxetU8FQ0It60sn
52hU5IAo7klmOKC7J43AoPJ37lnKbST2qZHfK+2cRUqMmk9Q2GBxsxjm+z5rOxE5
OvmvsdFS+z4lsLQBQzgkItOzJbHCN3yMFkEaGLi9FJd4vC9Wheey+5SE7AydAPbw
a6RU93wuiPykh4OyeEcn5wvrr+9TE731UGAkBZnHeXeAe62CqKb4zsWewVmOWFrT
Y2sHjBQWxclYU2QayTKV2gE35OA2JkbG1c/a04G43gRU5flsDyJfI0qXx9N3axDS
u+fJlIOnPkmTKKwP6tFp1w==
`protect END_PROTECTED
