`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9jtbSbo5TWajay0F0NQtRhZj5I8Y0OeM2G2EBDqdgtMaKFrvzpVSpBdKunQ5qgoX
q/3s3dVtcLnVVlReOytfyPkH+pzBZyk9tDma49Rg2n9/R2hCOlKJVPijaz+633c2
57PLo4Pj3cTuaNH7xhNejorDZs3TqKroLptl6iDo35nfsVjDo+xpMg/p029l/7VT
16uyaDY3l/0KMOl8QBebiGFucIQv1ZTT2Om8uGwNj1C0hKj+FezQYqNy+9xVpx3c
oxMZVmdQBIJHndys/QCqE9xzYI3eNHfa4t1tmRTc1BhXPZEPYEUjlqWb3DV47c26
`protect END_PROTECTED
