`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iYykH5YizNZl1+KFXf/TYwg3hiFyZNuMLIguQl1APDIMfWahbNb5zgWCbikQCSvR
H5GfkMhHeRtZVp6XELtn78V/LGPRG54usTHgwM6/5x0PHPIRL5KJRwfSmaxMF/na
po7xE07wHNDmA9hzZ8sNV3iIVL/ErfIi0oxrAVo9+cqLeNoeXL40nmWh1fOF58LI
7oPuWTqWcVBkc7riQl4EQORTA34G6a1JlqywgGDyEcLxAoBwYARfkstW6wBaRSd1
a2jkgWLMpDkna5wvD1R2ZjqU4zukuYjReqBhwMyd3K484VEUCePIgNY91e+kRyhs
2zZFRJDytgyJPwiQBmNAG3lg/6uP0pSZECxiL4iFhqZNkJJg5y4gT5A9WbSPYS3M
ok715d/Qe6VqCHwcUIpy2O21MvwkYpeR7hW+8uW5gugUjMPBCrZScjmbMojvCpL8
l8TI7RDi7ozHyI+DlyEtcMPPySf1nW1rHgsQiYZVhMTOgg7QH8hn1ZsjG6Byu+S8
rKsnkmW6ENkEDqDsA0+Le75Q4CxJtbz6kFpOZwqCYcI=
`protect END_PROTECTED
