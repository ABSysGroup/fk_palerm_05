`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TV6fsXWk9WbWW7bBzxc2uVuGxy0lqu0Km8gZoPUj2VeLBhgfdLOpU3JOgJgNXjaE
JI8PGt+UPQ1kYOAIN9DOAzqHPUIwte+gDp+MCqd9sp7ZMh2BriOtabmKgPGwmjbG
ETwfNzXfu7R5QOLhd78GLqTveSUMFJRC57s+tDAuAecuo9keHfYah67q3kljplDY
VTs2nrjDFtBOuvq2wvvYACMEqnS2uCjGGe5mJbDKy+LSfdzYcjWVclw05Xxt5cAI
pLitRudVCzV9qOhaA7Z/GRcov4/Ay4At86u+TZ+4mALTNuAGGblXjNahZHXDEfxs
E4SyhSyEw5aBBxwEwMJXucPgGiTLcO0fyfLYwU5jyMXFlHw/YjPDyYk79y4LB0L+
hhuWK+pCxeW8knx22EeKle1xWuZhTWoHiYWyEQm1tcWbhSNS0vtZZZkBL8kwL/hA
RTlj9zgwOwRI/hdQv8kJUJBTxcvwMQawOz+GSzjK3D2Ueg8sPFg2xk7l6IIOUBeW
NhPqfAQS1RyWanohcysSGOZsOek1NgZvErqBLhp7P3S9zxvb7NMJaN+kaPIyOpod
Rs0KrTWS/PGGIJc3Is2kKs/53RBoBe3ycG9GJz9bpDKi1/6K2dTY/CbuRKYoQZEP
qa3arVDIUi9lCUmXSEO3AMPm8UGhf3zsYC0C3vysw1Z2wzLuXo6RH5eI7I9KhCmH
elmfmUMkRwOvImLRHl4kJy6YtUZbIS1m734Q5bcfXiFpXYskIgN5q5zkl7iqXOhh
iZTx9CW6FleyOcecfJrNKFYCeJsqsfa4OvkEZ5KcBNcexJeMbRtNUDLur5L8taId
bQQBu9peiGOUN+d7zlwvw/Z8AMZ6QGOSpDVB1aWy29IO/exvQJQUdUIE2vJsZxPJ
9CWftD1Vyz98Kg2pS8fTILOIUjfArUBEwBEyFP6KwsGiWut2tAsdC2hzrej3XNsq
vXv/h/JyO3GkiYaV1jJexICUCHsjMb4PWbrMIzr3O35VQU0wvd5uo4DzaWDAB0hm
`protect END_PROTECTED
