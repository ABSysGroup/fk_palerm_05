`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ysGPoE4LrJWt0mvh/Yn5WbsfN6Sz8IibNTE+ukb4l6iSL0gTX1W/laArdRrppDKO
YCKE0pMZH8I+fyQv/i5sUOddTaDkxPAWJZp8gBcHJgFMuEpo3tfhahR8dPgBpLzk
aIGwFh9N8cvhzpGoB2Pvm703sJS3oS0yGvVBIMRD8zywAR5WJHUN9WFrjzkydYzI
Of7LKNwxRm2rq68iLT99YfOoXv5s281jYBJYIcf5aklr25nYo7FRE0v2/0xCAKrU
iu/uEhGU5SlvWBIVbGqJ8stOc+QrE0AWyJAey4t3r9U6cDE1d1KTa0jwU42wags5
16KBwlzxekpyXi7OZ0fuEnBh8JCxsc5O0BqpIAIV/DvbbYiZPtlo9kQtWcLrfACf
WX7sENaO4tQG/bDR7cNXg3X95QdGlxCTsRPpYR4KCf8AUiaAf9AhqUVEm542bqRv
3Bp9o32Jl3uwGWYpSCG3tV5cpSOLDv8ewFbECEGlI37KZycX8MY1sWUR+7SMAQK3
yG7hE8V1yq5qoeVEyUIZnPN7k5J2lvW99D6cl/pM4pIOGDmEvjW+2PM9oF4O2r9o
pG1784vAp3ss1h1yBV4Tr7tQsEYYY7C0yc+oQpYaIvBLi/IlL1sj7W4YfPn40ehm
7RLHF3BvuNHNLivLz3aUrJnCF8sPXACUlWmohtek+DqLF+WH2mycFy+A8sYpEr2S
2i3DpOKJ6xuB9dZnUBSgTo/1Ki5FOBFJ4tlqi+NDXEn7eDjtHQPr4f0Ob66XiJlv
Sz7EikdRUcayI73Nw3HZD0G8Sqxkwn1QvmFZRtS3DhzNywRcycseE8WxGLO/JbQK
9bBze7M5CK/i2Ty17uPYlahpRus/CjLAgEVAnN6gQ28Czsl1T/1+lV3hVyyEwsVg
UCmmGTzry0e6LPaiQ4JFZm+MIXK/C47S440GAJIQnpoB3mRV0OE1A0m9defSLj95
`protect END_PROTECTED
