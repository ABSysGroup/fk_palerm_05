`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
01JeFrdUxK3msex0AtG0x2kKu6cs+XD8K5kIS9qrSSO9CpjRgVXeJeY8L8XvJSGU
REuctAfvNA42XiUHfVLjzTtJNKBPPrilcAjs9sMHZl+om4qSX+jW6jUotRaPFO5E
l5yrv/X2fX2NLJeWesUWjs1vJwlZgNuAMqkbPQwcAN841bdN9Q/zyqkO93LHLIDe
mRqOh4P9azSbN41/o8nEzQKUppHMVpFZ//eSn0ZSIaE/KZCR7MNV1ol0Gq1Q5vFn
lsnLfkHO11RTRcgrSsY8JNyBcIfw40AL0G+oEvBwVelfHsaWkVQjlUodWIMnX1GK
8AF2PPg4iECBhwEn4GvFvmexLgjn8+vNzn85VkQ6ZZnSGKaynmxnwVwuP9lZC6L9
an8NtNH2dDqlOgQ/jfIzXtyMrk+m/CGghUcvKoTc4Zkc7+x1M3BAnU/bPPQzRyXW
k+xpjZsnweD95MRQygwKJI08am8GGISJfW1uYYAdwPpgvu5iyDrxCypphW/Yv2UG
y/FQWlkQwclAjKZ+q9HEIsVO7QGnD2/CB5RcOurUVBHn8ROSgL2LX+kxmfzkkIVh
cCMGYHzCSkJcg+xQAAW2SJ4F6eobT04BOZ6JGzjbHGFq/KlLQXREV7PAhZZzWUtx
fZ6kxXmuk/KcUr+PefY6y/M6cIFqzikFlDX0N8Ano8KZ1t6x/2cOZVDoNAJsiBXQ
7BkP77y1LzX5xHWOTgXPXeYk+xeqW+Ab5hshylIoAXPY2ABYE/auyhhkJEWMoRj/
DmtTwGF1FdomrZFAbMG9dSDERGvhtb0t2rqSaGJwX8RmtKm3HqKAl4wZE//wliFJ
EpGGnvckH+USZks1WB8vAWqxtSTcSwUGPlFOyMbshlOtAYJvPXhr79N/YWlh1jG0
Neo5MWvLB068PPqtVS7CEYkFAfnOeK+aIiVD/8jOSRU=
`protect END_PROTECTED
