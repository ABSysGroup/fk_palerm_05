`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+b3K1iTDUFiQMaA+inBNDbtIy7NPQXRkE8sP08460YEoNTzh8kbKMBnUl3KN6tC4
PVDRYxTufTH/nktFYLb4XW/7KY5IRcFK6xBZZCT+IjvUrf1qvDoQG+oAyHUA59Pw
5fqfi5idYZ59D7PxIvNW1TnOhGt2YKT7qBJR7db1T/5eM6+RPAkdqOmlnGdcCqYo
KEkQRXwtSTn6mOmgbxSOgQyyDjiQ36Xuw4HgOcwAwpoyYxAxHaewe0/e03Xjti5d
Qkx63vuLbQFarpqQeYiXsRd4GNALH4+x96qU5RoSmV/fw/AJ1n4dAedaggS1F8ZS
PMTBapBNNmDXlMkYI+RltKXKwc09/8WI+UFW3uglTealjzaXCnCbRFeZZ43nAbDs
3ic0VBPmxKuifxiLr+sEVhj4u4LYU9ilwfo0P0hxOfD0qnFGEeuY9PSPceknujcq
DYyemKCjG+c7Q25dICR+cU9VA8AvCT3rkvpJMdj5rAWunGCSbNuG45qFBzl0Raj1
G0h+R+FZkEPJSaym3bT6QfFh1N0xubN2Eii3vYti1cqfsOVBYR/vWmYkFeUfD5W9
7e2kHmHV/zoeEzC7lEajl1/It4EZruuY2UizS8uVR6Ij13gTz1vSLIJ0B6umclkk
28ydtRvDQ/Sgq7/1lijPDPHZWFzCN93Nym6S1OwWO0o+ntkDkoJ8zzR6gCQQgyIg
ypxq3mGFRyKDVhtpuuZqqkdM/dIMKdxVE+1hcLASNs+qAI+4K5ckzVzRIs1A1e+B
vLnfB4mzLpJAs9RMcHRttD4zm1WCJ7nOqEBw2RJEBqdqBVkWpuOclCftr/pJ+FUO
yVmxZdMVo5tVqw5m0YAPGydTJjJ6ZXYD9AKKuLzemHHKMhfBwnbsFZew2vVZln8F
AH418H1/qd2LbJV5SQGpdmm+z65VNQ1EkAP4wZDPjzocYPKTjW9IaS8isDERG4Kd
7Mbrg5hEzGff8rOhjR0PN1Gev19KhhXVErOQI9HMbb4rSf3Z5LD3EUYcTStGczcA
PfNfDDTFpqqE90pYR+ZRhkB8EXC5y29E78e7BdkXFOwjV858fDGPa1LQ8YceylZ4
+gsMBaQr6Dv2F34o8Ee4LxDrNZDn2Kc2b7h1WHaPdCRuO/3nB9NERltPFSwZuk3U
YFeTdI6+8ShO19gJ//Hc8Mnm2nucec3DrEr919G9nSWM4n7FXLzm//V19tcTRkGi
Fh1grdLUEYK9z60ql5l3VBjLLKfsIQbXCjK7ea+7E62/Gm8lwI49OQHmsd2KZGXf
TlHEzRrgcvRSqEJ/uznnG5cP3bFqcvVX+1bLDgA+ew+u7XSWm6n/kGpcknvM8pOR
mnbr9QHgTvBtZEOUM689MUhp0fZNMQWdiVt/LWJD1TDtqtQIYjp2u1iU+qElZOcy
0M8370iJracqZb0MXsI6TcNafjh1hGM2dvDni0c/0JXauBhZ0sLMrmtAvG/eKO0l
z1HCn0M7vhkBF7JZiVhrW2tJ66a50OceOW7med6XXY2vICRArV+JWVnl0/9EqV6P
aAva4vGM7A6x0RzgW0EyAapngH9cwkmeYXxiTYT8XpwOZkytJhJ+/j56DKQl6L/M
KADXX0kB3lr98RkHmbFDdfXbGD7/Gi3un+azwxF9UQlcL1xua0CHvzTWJ4+b2U7l
WADrc2S0xOSx3wICHZFn04SyuU8VMCqvHFu95nNMEkyWI5ddayxKWC+obh5YtcQ1
iCRVyvKLgDOHOwu4Qk7Hp5WajGsUYQ1lHz2lWNwXz+SCIB0v3uSpMizLFflEdZls
88E/MVurUXWS8S5SCpKs6nbCOv8jMqjsF1qIL/VfmuCjVo+LguS8FjP1IJzlK7kZ
9MFzHzCUsQn9OnoFjoKYZ4jFFPQIF/CzhIiwzkdZulZWu7L2llsuWK6fWI6T8D9X
aXwxBSa6m6+0ApBb84RwTONCfnbZaWY7nVbQad3xEDhHnHr0ubF6Z3KvXNUuNGDZ
itXkEdI+hw4BhApBKILKQEmlCgYt7MDCgeVVRzplMOOZAd4yfNZPOTPxftSIGBa6
brFEHs218ENPVSSxT/ngDUnnJFtCCdBxQK8Jx9Az9EeEocr6U2zlG+ob/sbbwCgH
ey6UL19mF0BLpbsdV0eSASqFMiszEOn5+JcGmhpG2Wa3Ek8D1pZBdbbZikoj/5i5
PceuewA/CfAuLS8Ss7re+XbYLXx/zg4sfMMQgRzhi55+XAb0m1OJbARG5Xe4JF7e
L1HCHEM+xLv2MgdJGfg97wPZKtmFzTktLOmELGFLn2BL7IkK7liRtP6teZd7eP9Q
8eGcVBkhFzhO3fWRPgHbg6127dQ8upe8ymKv9xj8v7QOhB7vMNEEtCflOErISSN4
NVbzpX2J3oeQTBWXutEWD1c/XkpuzJ0UvKHL1sana+OoCLmgCBPGPd60Z1K6dD8h
tN13/nH1hEEubUwHKFfiurWbZSH4XfS+1+VsKeihJXNet7G94dz/hYgB2Shhrmro
Q8PTxR3OZkWYVAel8fNGM0M9F9gaOaa6fGwc9WDBDpzkL8ldU+TsPv+NiCn0YDJU
y0nt2jbgayP9Gve4KyUnuqF1JDG/CFlPyPffR+ZmUqUp9ZdLTWYiPIBy7itC1i/W
K/a5qlBs2stReI1t+RmNvCUDWoAAaTMyDlSJLJAJ/r06O7Cm/ebFdQDb3ubfqvFq
0TFdN6osyrFcbKqTR8TOyusbRkl8DdJHujpnAf31ZQ9Q/He+Yp5EF45ZEPEQ1bJP
YzwC4887yPX5PJMDC2P1koMTp2bWgx1XILHTenDHYDCcPKTRRHag1b28uWCsCa3r
19gMZPsn54oVooidpoHM+3/F3xcqZTF15/+41ahiDisMeMp9r1xRenlfZ9pwEJvm
J1CAJ91Ip+pO9dP4xz+jMLb1/H2c8dU2EpoMPWcthWHhzgHqMfjb805a6/LKPifn
2G7MqWpeI2VknrcKXrZobOvtfy5a2WPAYG+qxQFvXCz4cvctkr1RgrgoN0D1oj72
FhYon3ctLViDSn1Tvugq5vnHPd4jWtvbjN2nT3jLERzMiagG9b7cjXzIfym18J4Q
HrpZMjQPAiB+5aGfBnS/7lfhDi6SH6/wq+3b98HQ7cb+ROUEc4ZkzrGlZMhk1azz
biEwY+6nyfoGPZ4l45TDi7cMl146sGWVrfb9D7A0Um/op0h2y0L8jOqzeIdHgFJg
iAxcBoM2llsLx9l1rY3G4nDkEEJqjWW+GdOKb9bn9hlFpF/TcZ9YgoZj8Mm8BoJp
8tY8RgjkGm5WoOr0xe5ef8MNQ0bzDKrN0659XH1q5KMEe3apyFKfL7isZM1MWuBR
JW26+SkoVZY1QrYE7PLjYrK/lBtqenMilMTccItl5SRlh0rC/Kl5CRjyLR7BFujC
6YkeH4nx1hRrH/pxFDUVVOcuLs7i3te4BtnAebvUpnl9DixGTccxENVttXZEaq7f
4J/nGqkjJN3MdvCPPTtM2/ptQIZR+9sagLCy3mHLiYB7SO+V4b7HJ0xA10Pq8Vlr
/tpmsIMSHAwAnUmfdAANNHVqEhWUO6FyQ3okCTlgURj2RcJNFTNtnEt4TCuzVIsa
4Cp/lYYX8nceiefus6x6KspVp3Z8R6Iia4/SWMboO3Ps01rrMgjxW+VbVq3nkShm
g+ok/jJSaYITGRi9yFGKz9aie1Ltj+D5PpmYIt1m4khamxbG0cJrN/C4AjvqE1JI
3r/vPpeT5/RKg7dYCa82CUEkUbCPYSAFj+JznA8f+FlKqmsPr0Vdhm6SKorrDPMy
zy4grv4SjlFI7MgyDxlb6PCqYrtSDSWj+0YH6DXPv0lNtepBkrGcWlvZta7unhDa
l0nWqeeI6r1NxyT/+PRaQrHI63mDbnB4GyeginzCoj43nlIrfy9bKN/3Rj7HGasS
y+LTN/lsBI+VsvG6YjSUQ6slkupLdMuCUrijvTsBkGviJmgjoTV1IehzVYh42xtv
J149NryuMt3M9f2Ue9XWmKF3o/EbSuy3c0PCniva2K7Rt43H8rIiPCunJvM8iY0X
lLjLqlv+V5GnMCg9mB6aerkVaWY3LvOqDXz17Up9h3Tr9arfT8UpHwegxs8HQjsr
UqPp2KrH6h97jB/XOvO7xtqWGZ4HOSq0+a1P1n/YxrCv3krTpInW2Sl/n+Z4T3rl
Fr9zKETQUwvLgDeYe+SfnOU7JepghjMh+ojkarBJPxnxo5dfqKD3cVg0zVH1735l
qz1My+uLyR0JVVwRu1id6BdlQZyeEFVBmiYVkxpi/ue3norpIv8VWbtP2nlLAgxe
hWozwG6i+/9VBGT2fra53VQyS1UcTBdipCYKWXP8gojLS0NuoZ+mztN0ifeMt78R
YyKtRhxWnXZdu2EKcKKjlsx6xiypnb/T+B9nX32+aMr7qFxlhMObzGlI12BM/Dan
8/DjlP/z1GyThpj/BSYzV4WoPqS3OEwrHL3gusVcwFtafbVRIlsVIQyXcynE7euZ
BzN/Xj7IsB8H5viTXPc2d/r6lAUDufLwOTZp1+hCHuGpRjmOfBJE8uF1rINFBTHL
Lb8JHCRfxDebmj/nM/4yqvy7HKETWY+97hKS40VUykXT1xPW+Q02+7T9FXh/uxqO
dfKFBgUMxNK9ZBcwk3VQF9pYvt12eSX4NJwbqcYFF3y2eG2q11dOLuAfflylWOWc
93QTuT0tXngh/Btn/narwjfHt/sQZC5wJFE9xOeuihXycX1T4cMde3xRAeje7P+e
Zfm6tEI0d9lW70dqc3DLC6ycZNtVAu00uP9u/luzFVTw0rU7wHd16Geo9Wx2QBp4
H6emGKHM6yV36mdIYWXM7olqjyzgtB8NLepi5esHJyCZq2SSwd9j8FXoaQiD0rCz
3FeN/cX5AVbgLWgdkExVgL4MvCR2zfcJmm2k5mmWX2WURJLJTjRJd+p/P+o7mqHx
4FnINyIgLb1jb8AY4y9hy0yOkhdclf5tVmJehM1yGYmZNdV2TggvuoCHFyhQMchr
ZStMPNxnZX/ngbJ4IGyRZ9mhB9iD9ktZqpqglc8lUlBZco7/VcylsZRcjEl3bgeI
j8MY5cEgk3kmBkIWfXuJ3zL1FZSa4cPKYdaunMS34E8vh+e7fFA/11ZmnuNdR7wR
pEY2LKmrcorzpRwxB27j69bK+ABRwKf9e9QE1BWqmNYdHJ+yGefGGuwH9qnL5I7R
bsK2WfV4x+jtWndBbvTp5N/fBcKJBy2gN1i9S8Y6moPzl3hDvBfAXB1FuR4c48Mm
nuhAQheyauCJfpdmu/JO8ceHc8Xoe6+Q8WU8JDYmeFPo0F6omD9+uy+jSA2eEKrV
0jt1WO23VLbv+xUgS01U2qxa9C6Z3Qlj/gqnd7BLVJmYuqWsRF0n9sVKPyeeqWcy
JmmpRGZvn6nGhQgXp4PcJzOKQlRZbQhsOSD/TyOqRzQP9LxvRxSLDA7S+S1sIJQS
GKQ/1p86VFSFuJfNTnXT7CVOcNpngab+06T5BZK1eL2HMLLNhM+wMqCFqSi7byrM
GNK29RqlfeRbUmhqJHMmnHkYvkLj0WSlyUk8mSESSRm2yW+nfI3TW4ZzUCMNmSmj
eGeTkmipJRrnMkdz1pBfbISKwY1xcAh5154xjAn4OBiUvBDwWC1DseBbZb19gYYC
Ygqjs3TwP1jC+vHqJHzb3onUZU7Q9hFgXoMhdFO8SfDKvV+szarUAmQZP8N9i2HZ
gMQA+oKDhXGQu5/kA4DlA6sqLgktk3Ko3lmjO1znq2GT2cT51ldn0l6BXWQZi5bc
3sPNMFxIPCXK4UEjwuO6zpbUUW2TNbYPuHtHZRqCOvee+woMlQgWiORFAb/719ZG
Pv21oZonEgTNUDWritzp3vo2mStR6NB8kqg4ap1MPARmsX6Me7yhGsztEMyqT6yZ
wH38/URkl7fnEPlLzESDV5EuLEtSgKK/76BjTq8y8Eux3tSeHaXjpfLnqjg4VE/m
Wfsffw8ST0XMJ8j8A5xj44zqAszkLyPZxkOTB72GUlOBJyewB5NFS1fw5tHe2HMb
fatXrXB+sRhHKD848FnLd9xY6AVGYZSHAYJKxpIg5Sjmiji4fvm0I2IvgcpD7gL/
XhAwV/pwgdJW68Q6GRA5DsBCjJgDKsA3QM3LWuby7Yg7SMWl7eivtatylwPZDIT4
PyIvSuLb1TtjDgre1H9C5vExKP3wIYqbgzt3geFuEWErFzuUJmqaZ0Z1lNsfxhlk
cvggH1buhqh77dJLhCTdiKd9ikBi4LzNffvASE6aNmBA9T4T6cvhdC0K+zI4gQUE
8CGSbWcWlTGW9ZZ6BI64Q2vWa+tLAxum9zSjUzJVMXpYfdGHJkm3e4nBy66tewOW
1Z2rQMrbywvkIruswgOQ2gT4uCgbM1fsQIE1UjXDIBZ3dSKhJRq/XIvKGQA0b4gV
6O8h9wuz6Td5DFCtZwHAQdmM4eZ2cvcZlS31NAkBv89gYmXZuuwW+A+wWxxZ1XBP
KXAkeHu3ZorJ8xc+rSgKgOsvBzKglKC81kjG2Pu3PBT8XOLaTgBW+URqElmgJo6c
axGlIEEla7UWqmyw9MQGZmY31ia06O+c3LR56sU8e3JqzDuZwUZ07M9bucK9ojSs
me0sZtYa19nmksQ1Nlqg86qGJQp1U2yfnzsSy1jfpkfzsAn+BBbxnvEK6IAqZ255
8SlRxal7Khk2g4IaRscsu9zE443rx9aDdZ/xhX1c7gCfQ7A2jZ1sEE1krP8NMp0+
sOnzyvaQP4/kSQU+LW1R1JL8wJIGzVD4EmuMHrW6c6XDVf637HI2wbp6YbsYe0n/
y4BFa6LVjliReeNxeTJxbEKa4DcmuucaUQiIHWrRNCFdPQFFBeeLRpaxxbPNp5q6
3zNj4JFwi19fc+3xcJsNd9gGF0xtbFmMOhcHlU4wf2k0Hn+ZU0qagp8hogUYekVi
yMJwDacLoEG66tjnfB0lM+R2ehi2LDyGnIxcroseUfwarknyz7rDW9RuB1x/8G2+
cM1alnK5T08ILQnJoOnMCfCUzz8+EVh0uOsWI4MuPMB+IxsiGjC3aMFxu00uhgk3
2HoTmoU+gL2PipVH7SKF3mpB5Ma/xy4Ymtd/1JdMsf6gBwZrURjAIhQcgt4COEzz
1YFD4m4rYpZosxveKUfEeAM1KOcBt0JSCaKo29lEjNefHCfZYtT/raOEz0oyH6ys
8xGtrN28Lj7pGSbDcYrU3JMGLYpcZs3bl4FEoHsSBTh9nWWiSmB4wCHS7KLb1kpI
jFm7A3RqfFfZxynVMqtPmw2DxDE4UOgT+KAbvl8oLt1dsmIZ/SC6t+ev+Esmjent
/wYDrjKTlgS9mPIaBFIY0pWw+uPvq+ndztdXuj6v+Ht1L69d/HJ/lLlDR3taDTUi
KQlBqcISC3xUH6+NOILnNul1/AeufoQ0bnWDE08RxrYuHMHk2gizuv9x4AeqB+WD
Aq7LDcQnjPwvcjqkgxIuGHt/WetOhald2t2nXoLCrycuJfb361FroYN/+mQ0hiqO
R1dG3ZHv6jsdYRPau8w4ISolHUQK4vZiJv5DTA7wny2mI9ZnHdKIj14y2eH1BiKK
OfIeqzUZ3M3sh0z8ipROdrSwXSl0WW51RYjoQgXzmh4BFD5GjjnDw2LmkMsdGrO5
FXBwVxYU/1Ga5IlcnXUyYybYwb0Kqa4Ekc2Po654BVSkxwW3eCPQ1bL9MqSAXuS5
lyeOIImcjwhOeutSw1aWl9XPj0XpOk17Sfxf+CUVfNWge0oYcaf0K/DWkPUOc5yF
k7R++BAnSQpGataLsiKlx4AlkrhOEGmIubLukWCKC0XAUWf8GdqeVWYpS90YghXV
dZwiY5MVUk4VIhjUYyyBdwzix1EPC3FQWu5Kkb2ZHeSsTy+nOMP+lMvXtjAu9ZTe
uJgD//P+5fEkCf7fnTOgoQMRfMnpxu7MFEDXFodGIst3a9+uzLLEMsSyPTj9RwbU
INY+dzhCnoQSmRfuNNH2OhQLemzwh+Mj0cenkppdfvKdLF7033WTheqM114drhYn
dOp+lTv2ioxiyXcPa3xJqWfxXr9LZu05KPQ899d6/IYI5+BJxA8BE6GkpwySbPIH
niI3B4L1OcMt7EZ8uVxVjhHo1a2zFWFN52s6krwOTbLGsk6hnfgkajlnCvalVIoJ
/RXHaUeD4B3JWvqAOQjE4pgHCwMTuaFvD+TE2Jame53xHAQPVGi83oEx3s4/ybzj
ON2uByyWUbMVbDi/p938LDRO3FK7xi0IgDICFrg95mIGFmG598Eni+Suyq/fiz8H
p6NRx5lLZQyfnLVvhRuCTekqCg6JSc7pN6Iu9B8wtBk2gSlnzhAIQt3moWxr+6js
9jg4SKm0+a9HzWXUqcGQhe+Q+YQOVREFs7jhBt9zqeknAaiCksiMhmoC4mKzQO/B
NlHNmJvgtbU4Hfha3obBFs6eCNFDw1oTr9L3uLGlFU/AY7eIMhBwbUFsd4o3rL0u
c7gaSG9g5p/rfxM/5idXK+LBPEpQ2LqCGg9zuKbOyb1oGD8ocQfJKPS7CJIt+h/f
d1aA6Y85h9hEXLxlqbJWb4Dy2591mbHHGWYf87sj2NoD7WgYmmxA8QmfyEqTFtny
i5dt9IGjTrFwg23GxgCZkauKsRX1aBbIBHeZKhyAMtKhvvz2DxpSJJjptmSXtUu9
n4VsKite0rvlCZZv49DJKpJ5OtKyCUiXMInnibOq7E3iJhKGVMnXKchuS/1QfCIr
5d4AauIEAJAa+dLmosQObIqScs/NOMRHoD8dKnrBfYMIufSzvSAv5aZ7rks5hbOV
Yg02+J0Gnm772ad4Ub/qlGmdkNK/V2LMH0CIysmxMH7a4tLCitBIdUoNF8+guHdw
Pg4dCO5Tvvgt/1vGQEHb0J3243bMcVYgOiXqWp2t2gBDRdU2eqYM6b4o39Q/d/m9
gEnPhn3Tjh/7zhPp11tVuotdiyfFyzLEgzx126mc9jfZK/3gGDejmuERtoNtL7cp
i7JpT+DxUDikJlGSUT69bzoSWki3KdBV56piVmb7uQpNJm7jbMfbQZhFWh3Q662f
RkHyPFTNU8dLW3S1QGNCUCCSsbdAA40YPJNlzMJI4limbgez54cCEZcfiBIHdTIK
I2T43euHjAshywZ88fnr4vDiMQyQs9E3s2xU19dMxfjUGJAia+2BZR6It1Avkcl6
w+cHsNgGa1s8XlnIkq9lGWwI3ZTvD3CjzWalc95a6syXnkV0ZDyoHuC0nEbki+3n
ifIeePe6rVENDsFu5+DMoUqEto7a3cDSqKvP19SLGirlicoX1A/v4OLc0qPtJ6Yg
cHN7UYalUf1NNQ63F3Er4oYqBNTIXzH/ZG7ZTfX6kg0Xt3TIByEg1cXXyIvmnl/9
5ZVP2VUuqZHsSJDeYOq7S4w44kTfu7yml8n/tP+XL1aT3/aPVTuePJ4T0Rnjj44/
TOBeY0jajqRUu4VBqxWTKnHXN75PIb0k8ExZ35hDZ/+smFYV/m1jga2On99L+D1q
k7AdXiqKR6ASe/1/mvPC0RGGKbpnQcmu9P0+0nDUg8EMStbzHNjcOpXCMzpL26De
dWZmI2z9Q46viOpG7uuNfhruVi1lhnF+NWJ40njErHGAPgkGZLO/QzH377/AJXYu
x9gbzkROvKzYCXCY++zRQv3zmtCIYs1UlpUzTb6ssZxVSnMChvIVFFy+XeH/Q1a2
vXdkmNAbT4yT4vWuJ8wNXEfOKQ1NsHPJRRVnKWfkQN4deDuuBuramEep/DhzsXml
myjqNatl0rxEfxAjOF2JiQOF4V9psh79E+iaTGsFBnS782c0fuUB4ifd9YDrA+E9
IB1NiOGhQnsy0U7NHmUjxDcMeribYtGYIhzuLZrpgMoUe1h6EGeJ0H4qqiXx/6RY
MctCR4FAI3CgNC3dbjdRH7xBtV7JpgkyM86x1sp4QGEGuj3lyx6FTXdRRnujeqQ5
myS+w/oVRwDOUMoOU+ih0DF4ualFVaPHCdUg6AYUMBpoU+534J+SqaKa9Nt5Mr7W
iVmyUJ63sran9dNWxlLOT8Il9zdDzE8VfpfctEHVC/C6aNBlTBRDetN6K/dN7Jo3
qHjKI5O2pI50OMDhKaEZPSdywGYvC86lP+MSXGv/ayPCBLcFzmDWqpnTazNm2JtC
IhYvQUWeI/a1E/8Vw7IpB8VZuFI9txhScfCEbMNv/BFujPXNjo1A9SWee3+vMmyJ
L3YRauv0gmu+n1EyYqcNlVL6vhM57chAZjhTsgm5EOu56NCt0bY/c0FK+vnUZSbk
iIBo9YcCuobQEGgSnJqx+awMpI7FAII9UJqF6UYE2GujTm5Eh6pNlzkyfAPaQzQy
`protect END_PROTECTED
