`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6yvIKRvHxHaO0q6unjcLfY6kZCrQ572aXl05dbsMTrZ04Jixwo49UTrOzeFQdDH1
KzKTzPFZWOTY4uelXpqfJe8WFFzbbvagE9djOj7JQ+FTnMERKZCnH2kUJVI4si49
2CoqyBBY9uW4Uup0AFM+axxxeQ8XyVBbBnT6MJShrMIyP4Xnnwn6JwxFc0dJ8I9z
pUeAXDSVlhLRLHTJOHg3D4G+oUx1Ap2tw+19yMk5HCR9ZnxOVWmiWI7sIzpSbErQ
WK31gfuwpiNFOCCGK0jrFmF/D4X0BazspNZ11CJpSFrZK0uIH8Fagie+oV/i9EOf
R0ijTFkQMOAzIinfkfxsfpTHuQVworeK95ALxREVYdUu8TY0h649mXy4LsmWHRS6
MXrD3vaKqzIUhBabgtSU03Djy5w3WoxtHwD+Rsfyo0k=
`protect END_PROTECTED
