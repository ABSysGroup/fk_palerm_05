`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6OEAmLFdHJXjxtY7HsRBB4Mmc9QiOVrC7D7XDL01L80EpR/ZA2+tpS8YZrs5IZGw
NjsQJ3uuXIlsuzGEWCupLzDCh7JEGcBlGQeYWYnX46GfAlSW4Ar5NUGo13/oR8vh
3VeSuPmAfkVgAO9JUT5VKxNr5FuHmiGWQTxH1Z8CtUH2/Ki6gcSPYsbZMN2T42hl
BPKpSYwEQfX0KJNpSTIBdxzBsM51rqs/YAbmG1Hbu5WYzKOhQigSh5sQsqJxz8Em
DUT8bBUmtUKbVcPWEzroWA==
`protect END_PROTECTED
