`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zAxX7up4KXLxp5nxgobqQUyrGQCiCj3Mbntx8PhbeXeozg0PIUR+SirHJvKGCeUt
g8EzLKTNGddhKY35FEM6XSKkxrTr8dpCfKNqsIRYYRjbv46F3hEqI2j6INkTvPzy
4tE1TCr88wZs+ZiyNRUGaeTFMzM8tivwJ5tV7rpz9XyfR/3IavV41Ye8vL2jHAvx
7CIkDh8b5YF5JLyt7xSD0AGH0KJ96Gbmiyhu6CmhJpx7LrDZsDzMQb67JLw7xDQc
neTQ+W5+V2eOepxRwK6HioFJxuqeVPrUov6juDZo+iyTxxiiPTVezKttMOzRSjup
NlcecPjIdT3NaCtorRjBh3fhY4T+bNJZ8WJcxSbyLUYeh0mbUl5B0kqsuEWYzFY+
IUOY+RAGaXb43vIJAraAspssGC5Y1Twon/0N8mlvMM1ffiTfNxqRRp4AZKW5xMZn
WAGbD7ZSsfkLTP1YvbtLZeKUWG2gA0m/ZXqDQiL7knGluTMSctcsTSEYsZJR7nti
SPE9FseVhgc6qB3LvPui8w34u3aK6BOXnvodaLJaONjPmLpJiwoCm5QoKRRiEoR7
XQMnx9Ld36ljHjEtcJd/xsucPsEe79uBsSIwx1SUB26rgh4mqwPxEehQHiyZ86mb
3xQAtSuCjS9dQipCnDvioxvhg5mXniGXVYpESpWlgy08NXFHKW/NHftnnF9e8O/p
XHvVmLR18+6j4N9+3OPxA5sx4AB4RUz1mCKiWwLfMCcXB3rqQ8U7IHVO+GQk2/kY
ks98xaijj8zlAqt+MLRlx1n5UhbpLvjlphedOl1FRXLD58o9txNZE3/jdy0+Sj+W
pMY6Fe1uSMvo+JvMCBk+/n9m3hhmCgYz4sWAJMtYBcW2hXrzsr6TKpUyvK/nwXES
MmaahdjymUXXbg4TSrmMgJn34BeyFsthQMCBFZZlcIhr2q2huMO1oLiI6tv9Zfkk
ChMnuJBIkbSAaLAGSCK/lqlo4+8GsilA1srs7uLeluv0XqCZ6Qu5Snu/dvbSroZJ
E7tN+0v/3k4KGO2DuWLzQumTQlxbzo/KH2+2ywPDOyT83FSlt9Jook6lByyVTPzK
7uD0+qEWigbCuOf8QeJr4wv8MzRjK0F8nAs5upPkGPx6YA4tHWt2bHfgHLQsMR2M
aBn5zBS/VYPAmkQ61b4tmhOapzArfFEIgWV9cJBxwuFPsFY0MSLvE/t5MSupbCTD
h1WWZXpp10MtzF2RMoMCF3heBryfliHsemp1bD3vTssSlIR8pXIXQgeO/P1hbznQ
3RbxArZfJFcYDbORcBnHBtgvAu8hV1VH0wJBxwmc/Sv0EiBrHYIgymhnGlgze8x1
23BbiBr4pwdCVoniqQE2xqq4y7sw8PEGcb0SdPxvG5rE/40ofUTRztv4OJl0Oc/r
fvAalQ7l2oxPpj8LEjjZNf5XypPFwaobfExkJykx/gH/VeUEgJyl/yE1iTEpdwry
QaUGxG7Cnn1COjA5pA8x9Y8J5i8ff7iBXvlVvl0rE4Xb0K/F/CFaGIidRG11ODXa
Xv/K65QtZwGfh9OzvLzn7L33AvHWfE0/iLCBIvAVxFQlSuJ3lnROBskqrFOZ85ed
KYHZcPxVUA108I3dlATU3hr/zFshwrZMR/4Ic06aFRUvWcES1b1ZYaXgerF8+mNz
0SLLWaPAY+4vaeZ0srFqnvcnYspYj36Bb8EmJNo6/ka0G6fmk34AUgpkl7KM8VMG
qFFp9jBeGyaWXFClingGPccSMU5azpMF6OGcZwYPex0iHJIZnVEI+d9wWNm2QtqC
xo2aXwf3RWI9gY3Uhg2EaWqtqP/VFL+L1UNx9OowUmtmJegs1IYIbHybVxBRfDiO
G/7fssGPfMj78Sr7Eb2mrSv9KTlHdZ1dGFLRkX9B90RmBi+xC9S1eT7u3vXUjJ64
lzZEgVtCHkEigAWhiuN4yIGZ9xEjc/zoYMNf/aFYJmyyLawd6CXISv6KCbxtWdmB
G8PdRVjZFBv9lVygLxCeHu25a5kZ8EuPzmPQVre56Jclkzdzfa6SY/njLiLJhaqC
A1b9SOCdWuc8Zc2fSLzWLNYP1u8urQ+u+alNRfzRiDjQa+RZBx0PXtI59LaPtSpY
P1zItyxFay6xgj0zcYY4QxJ+Bt4xAvIppqgxe7sCd+qrl9RSGg/Hcu2ysC/eTMAk
7VPbPpXEZ1HxndXk4VSRFAuyFl2H+Y+g5tdf19vQdweCnQwJQJl18c3iHALOPjVO
mf4iXnFDc+ju0KWcfPGmqY/ks+Qxpd5Nj+ziOwuGYV0nEi84g8aPQUZOeiLj07Fn
x40G/u3ogHisGrcPw+HU2lkbjSHR6kMvTfuYdbX+u05R1+eTceoKi9r9/OKitR0Q
Ezlqvr2/28vwHFL2NzqsqNOkpuaMNgEo0mLwp2MjmxCWptSbjnr4ia5KRlYTmYTZ
0eNev7oMlW2GYs6vGWyr0bjl7P5Y4ej5Lq2S7nvuOEwhMqIBbtslATnF99jeQnvP
4M6Dn9fKAN6pTw/t2LS73HdQ2Dgj3eLqzBrhLCeFPehMGarRZp8uffzhQ908o3U4
P0FCIgtG95ww80guGE8NCABTYBWkeR2jpz0YtKY4ixW7JwtcgK76a27NlMr2TSVQ
H2nB81VGnb2sPqckiWQtOmpJvkGaAEaAFsi14TFU+ZdIGf/RDuUP5wKgKm2qcVHQ
uuFX+aNqriIdSmwd7DdSZ583lCcczIXw1P5cQfF3jsul7u519+kjldqCMmT/ovq+
TWVyDC0f0rygN3jOE9Tml+VS5qLUDuPEBwVzvC6Hwe+Zttc+Vw4AwPEBaCF3L2Gw
Uyu0APPfzIbimQ2gTW/F7wVBmkcz06yzsjWIrBDGNbopLbIH8DXWiEOev7A845B3
bic7M0HdgMqBxNp4hvIzL2Uq9MgpfcVTiSomEmmPW+whKnTBNLL0q6brClc2nqLS
5odJiQOcsG363A/L3iS+VGlZyeiIJ3arQb9xxUNIJ4RQ76LehQSthKxKUUQNe8ST
Dhqf3BdJD06NpF+w+PmvmHkNEhEv4U+WZIe1x73/fDd6NEi1+L25hyvk2kgexMC6
c3A538vX/lcDRDB6vXDi3MU+7Y0XTadp2T4Nkb3GSonZEt46nri6QNlFevrHJMAL
fL/0nGz/xLnNloVCqnW+TJBzRpU1FZeUKQOA6+oAsj5Hgf/K9DXS+cAXj8qsNvxi
xBG9IDMSRGq7umoC9GooCuImCixcsGv4i0hziNE/IF/l4xrZQpDXKsF33Fif1SCQ
nTYO89mI/0zalIBZE67OjMdPegui3PnHMifjQYpC/Lyob7eWwrTYJDG3Vdo4RNfC
1m/Ldl2nsgdVa786G3vOKer7uYNkfrzv+jRwr12YX+B5+3t3a0Dxhc0EDHqs81yr
gVeX6xcuAGyOTa9wVEdpN6feUKHxSwMvQr/RltDNu6T6EBDDlaYbGMhJJAiXRE1H
dxdxO2V9/3gR1dXOwSSlCyFVlGV6Eef/ioddC+fkHRTaR8FzWhfK/FB22fO6ifwS
pe/4NhGtsSJYW1ycBBMN/z2F225KEipO0iR2L/kTNvSjVQNP/SrcPqMz2mb47ZNs
YyQHMM4XOLwm2Jc4s53gjF74XiNYukN63maU0aJlMr/fXJYfZI6P5OPgc2LG3xRb
wDlAmcKzfypMBvWCbn8No0SeZuK89o+/2gUXklav/cWvYhGf603E/GYXzUZmu5Th
ludyWQNgYNhub+2GF0hI3sfc70empQVdD1tc3cRRsy//89touAR5foCFm0G8XYUs
en+GmtqYokN27E7LxtBDxKny+ynkaKgPw3Njbj7a9Y4UemPBwZ5wVjUcgS93nP4L
IN/80UeWoc7wYyJxZM6+aODZOjhsRIOVtHmlms3HqIX2USaPpanp2OjZx4pHPJic
Rr7EbEorXaD495BQXX8bTnQUtnvyCdBrNcitAxcWz/MrpPNVxsNWn5F2LKNntfzi
e0rtmbVyHCX+I9V4YOFIoYqL1ZAQNfY3jtFZYHYmoB72NsrlqFOSzGQIVDVNN5/I
80loFIT7z/4xXDXGak24Gm6KI1VnLne/dQIVeffPUDZ5wpPGvtiXufw+EXhV2BBs
i5rjNFOj+Haf0nQKp1f10P4Zx9XuHwhTnx0S3H6Svg3X2rG6ROQVoY4uazwcgdHu
vhpXj1d9AgrxsKQbru7/UolEqk+f5ACZtv//33bihvfsw8VEqmGgYRfIKqfDlfJN
TGqrlWBr4gC71govrWiFxlaBkdbQcTZXnj9h7ho6F9I0dUIfP9iyTjw8nhsgog3o
OePkYiq7aPwr36mrfGm6bwBznnuIYTjgYSyRGO+Ok2KJ9683j/aEroCo+Gvpr38S
h8ECXMCzyvj9FE00plQcyHkZeHJS48tmZ041Q3KmGZTKU/PtEnBkPpAyZ/KPSx2N
c92Htb57R8wf8a6OwOrkq1oxzFskPkbD9FKfmeJvNVfLk32S7Re1+y/sjpM/VaDA
3dCtDWq1QTVum/dRC2xGmwaWTv8hIb7ExlisRv0ddAestm6E1m6sCI1BEKLRwAVC
UfHBTa48xUUj+gTgoEpoxiXBnfdeSu5v7kX9Lx4cVO6dsGe9lorbKfZa3WQ3NjBx
MWksDleU3pvk3nKtApzmo0BOvJEOZMuuh8kLM+cdZsF22/C8xkztM1P0+gsitD5n
oLOEAcfPyCDoDvTLG8miimEeRyB7oRe+jH6k3trkm3c5TGuJ9+BgSPoCJWSkY2+E
d2BraD8Ao4aAY0gCWYw5/FbNm8xFRNXqVyGODg+5y9Q0+IwGG3oEYv8wdx2KPFSB
8tcWQhofsHgIpiwFRJiOSQ5O/ASoOOkolHgT+EHzEynWHo0VrOXcS5Pm8fUhUtDW
AOKKOB+Y9knrHRO3P1Zn9VyVmyJODn1bhVYfo5dpodi5qK686Yvqo5JtvZNxlcrG
3RNJ5TC1qEYSlKoAh8GmTg==
`protect END_PROTECTED
