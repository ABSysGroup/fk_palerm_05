`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2H1aA1XvPrk4Oa0vxXUvy2nofiAlkouvfU+naWuyJ7Hx/rl/cz57qm5UOzfx1KX+
Ol0KLFhOAQkQAuwQkKNjETWNVkWihGS5HRdMQtwdGYhwceLyo3IQAEo5ZoAKGxVN
kWhjjvt660jYp3b2ZGZG6bksf7q6xvNGNyqd9VPAeWt7gHwGT+Hv0ipU5GzMqU6r
kXWoa6eb+z6jsNVjlY/EGnGVT8CsSD9r4K52B9/zVH/pLivkWZdmzBVMxZwTCV4C
M9PRYOlVgCsk3MAMkeew3hGxh49sNSP6mjjKoUeKzgbNZGXpUODpGDTMkfYWOv4K
Ta00hIH30UmNCQ7ePZCfX0nxdnOgB7+2o3tbsWMXwvDYz3ai3yya7l2tJ6EcRh6Y
QK7ANxT7l1UnRPIWu5Y1qdcXmDBfFG9d1HM7j8FjWux05/ChiH+mVomtqQZKxacs
eOagkxC4RpWQcCU9njblGPAhOzZ7FCh47K3gl96xfxOMqURgKI51vEvd9AEd3/bl
UXhzYd8gsz0naxle2+kM6R04h0Wm+Rn4wTJAYDZb6r8gtH8Xt/3wLq3cHzhwTLjz
wjgX8rKKBh20c5Bp+TYZNSoYFIMHUbmd1Y0dmcVf+KZ5nnDXxO9iIwYN89O4W+NW
0lTmQeQzgE4Fewwi89JlbGJTtvOPKkIgCQgj+Nwww8dAHAO59jhYfegWW/3qpiXl
79g7mvQSRUDCg7f+Uq2bW0fue+Xa9umPrEJXyNI1aTETq73AfUFEW5V7/yl6eYf3
0/Iaks9Ug/nk0BKvkYYur6/DQLoN3I0rKsDgX0dwxvDFbn+M3BTVo+k6iPtJLmYs
NLFbRrAmFyHlU/Nnf3c+/Qxab8P5J5JSap9D4Lqzr78dwIxWIlajZh2wDk+sL5Kh
6LoW+4R0LH0PUHK978pWI5v3HRAw8AB0VJhS96xS/aq+MaX6GqNmoGiO8keYrrYF
x8eJmxlDRSFHPLBogcLW0Tsz9t3Vgs7X5gN6/EDZyl9dRcaEVf1yh0rJs3nwjJ7X
c3wfJs9Hywzbt4DNYlxB4/CGZsB8Q5PB4l40XcsADS7yW6hWDQ1mBZa15GQSVSqH
Nq3DQOMTSAmMI0ZDLOT1ZmQVlgfIi7GNF9Wt7JIZDLLMkAxz8TrPizo3R9kqbbiC
rJydv4nn7xtJrxZQoGwGFIJxFSWQ6hmTH4LYVGLCPDeT+H4sqj2ei9e+ASG2A7KM
VXT4BdyqHg3GPi+ndgccprSy5e9tf665pQzWXMyN2oYPw8CzZ3UyqErivlmiEvb4
musfhJ7LuUmwpRvSMRoSDaZ0Dy0MJ3nnFfmIttBdrD4lMgFFAwiHzeMbTeJ12PJg
FexhI6HjZVpGPa0JsPZLF2lufqXMqEjGyV7m24j4JFOo2zhoeMBs6TQrFGmQ3VXl
WWzY1+g6oz6s9WnTQM7xskxIwOzqzihp3OizHeYgiEpE7xHVShbORuADAusJscAr
Hcta7opigcMDCwOJkLaKjondaWdgcEeAxtv9mbNVtp6Er8J+7pmNqeK2rl7btUh2
3X7dUoU9kN+7IIClCEmFoc3BPjEhUb+EikU1fQ/Y6HTZsZ5NhhlHbATPSBPzrny1
3sc46K+cYylHxjvigFkq0q6B4iwBR2k8HvZICxmfN9Y63hxxOGD1j+v67LQRD3pl
9fR8M3fjd416o8X1MvTMCfqgGXiHqjxeTknTOwj/ODrnqrDuILzvzOfBnyuLvfcb
dq7wyLi5p7YM+gC13Gx2+eEfgb1vqk1sJyPDz+ygQJ4daLHJ61xJPHtrvlF4c/Wo
LLB96FIZOzL3GzbGecHDt9q/vY5b6VotBl5tsIplL0hCARaOggDpBpxv7bdUaE8Z
+dqR7AowqXXsXS2ghky7xZ9X3z5IHRLCj9JCPNzxaa4pjnzb+3K2okSfc508BeuE
qPN2pQZd2V8chKRrLGZHsh00Jc2jzg1ZuiyihmPP9H6nACUDmg7pFz+iXZ0mgM0t
W1PRyiy3UhPUxX5rSFicVTCKCAE63jGOYY7R62ZusEYNriJRRD9jgFGIqkjqYq1h
9bgK4VxRhv0GS5r0uNUIHIwuhAr+LygINCIK5+9cXLGXQTTuVSFwodaGuIl99ZZ2
eD4dzpcn4V/tGsAUEr2kH3bVbGeQvswxlNRY0HzTuCVX3tzEYaTu/DBSn5BP4xDM
mBldFF5mTj7zDjgj3tup3JNlShmQlASq4tS8hbIEm951iub+wAUPltp991i8JwqV
Lj7laRB6tt7fH6A24YtvMw4VIW98qaVa+FAScajo3QZyEFMEXCuw30p6SKzHm3g3
o3qWdkjeVZG2rkHeNhbsmmdgAcovYax9DxnQYH90Yg76RMcQPR6+W8PHGyt/5lzW
/YuOX8FXmhyHr5BgxXaTPOBGLDKqoK73Rw2wa/404fbbkpPpadYtnD1RMcnYz8yA
Ay2zZnoBdUB58fTktnDnpDJHWtke6rl/rrfgrwudcDP8yQ51GOXmvzlRnnfNQ04y
yyDqfrIHohdtcweuRq6Ahyo9MEtqdVt/lqXkfjznK7esK3dKZTc3KdBxRVm10fsf
eVjAw2SWzIARRsCLephyQsb3aJCXZC7btICa2n6CpWu0/psrIG1Rbu7lrXWwjQA6
1w3Pmp14KPhltB+Z20OdYWSodjL2WV+cx66OovRVM9cEFFsPLXbR9wU7mycRsLRC
XDYtt3ZiLC/XVunylpCTo8TG7XpnoDixGqUkLl1LwjQHHVoDfC9E5hHhWi3ze5su
H2taxddes2rq3TjYU6aINxeX+Ypb3r19rwdPtamFDxa2h1cxyGX+lL8Aa9zAeiCk
5UObRGhT5cW3NjpxE2P5jTXQmPDCfsoPHs0JRfY7tabkXfcQHJSwjaXI/BI9r0Xa
L/iQhjK6VYxZlIQxhDgfOK+0b79c/YsLULQZZHxpO8s6LgrTotN/syIhP2+Y9K0E
3roXsHAwniOBQfap8r/OmyufpG+jivNNNP18dhYPc/MW8pCnr6+pqo67f0/n+FZt
1LK4FFdHTpKGd2X0iBU8glT/UM7N4HKVh0aO1rO9RMiZONMdtfqT84SeGjduXsZ8
Tza+gWR1Ejf4U/3gQVIxMKo8MsokgRLgwp4RRWi943h8ewW14nmSYNwmE2CQMRA0
xxdkkvudDeNW0vfAKsAgLn2YaYCFbljOuYkYt6dv8Sx7GQn6UAR6fs9gCHnb79vq
`protect END_PROTECTED
