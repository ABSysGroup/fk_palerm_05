`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kD/MX2Ehs0VAFTypKLfepaPwi/E+k3V8rp13g9M85mWM/7qBl8YcwdcNIJmFmd43
zgvOhocggHFW1wx8zEP1/kBwaW8wjoRNDUU/cBO8Kh1qFElgnkUg6z2ngLtDaXiX
w47MIbADsQ5MVl/GKagy+rDUfPnXZez9Vioj5D3yS8hJrlavv5Bw9Tl0duWYFEIK
KAjn8wRTgG1f0DuNeWQ/EqH1cw22KxgUBOzJoNZeiarcKEeW8AUNsmvfsTSeVTdM
yKnrZi70ZgeqrFEuC44caQwoNyBFrBaBqyHnAXygOg0f/zqqC65kjmWYAJhbiuUN
EkoqPVs1mMXIVhuSL60zGOZuRwtc5PdGGPGPRryex1F+GIw2Z6ay6sjj4sEutUy8
VTkyTulJILPKBwTHxDY25+CH68Vsx3QHZPR22prKeehIJ8zoFjzXk5k/4Xk3DukD
v4zFZ4UzRVwnvNc3ZTNeryeoiCjGlV5AAyUIR6mh5JdIr5grMQx5oA4hcMaQ32VN
ehoA6q0y6iY3Q1QyoeuP/qq7bxiOAPxB2La6VQwC5Fmo8PKfXtjBemC4+gy/MWF6
EVIr0Bt+3oV9le/9vlmos2qOffEripOXlVK/iFHEcghr53+fZwdL3BGE68P5hHQ5
w0y89X/xxxsGn0PgDkvoPSUu+4aQuyDNH8vZcZU8jRaI90D/2PDYVOJx518krKBx
fSsyTE7+xh59LLWQkPKleJU2E8zY0qLXnZx4X+RcWA2YdLDzFLoZFhOp/kipDKDj
zij/iVscnwL5KwaWHVOClx8G1zMPkICeH7ng6ethjjNyXPvawGEpIaZYMfepfmKZ
pFzim3r5XqxrvsQYZY2j6Gb8Tt5NjsnZRY+ZOqpgOoqYM3L0yrhUnItKpgFx55Sg
PvgYxWKDAldEYOSToKoE5klZKD/00BpKnhpgmbPREGU1Kq34z7U8NnsJCOqFzGW+
hw3psWQSFdDS5N+7K6IjJ6Jr93eYjbRkHVh/dEks3H3lL2wLF9hOFMo8pIpC2JhF
nohLVzqB7tcJA+mBfDsMLg==
`protect END_PROTECTED
