`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1r7pHWhNI+XIo18te0YLs9NOUKsc3JV1zIdXMPobPH9meVakRt+dyvxT2gzbZtwU
6uZAsmrhmWDQQxFWN9dWVuH/3jb+yiXnnFRfkmLCW8Z8fUtLK4B+yeM7BgNrnh4x
USqDTSX32KA3mUtLIMU5jaUyZW/h2NogFv4HGzG9mR4uARLKUGzaBMRG3Q548HGP
6wn+Rohm9lVETpyT84YXTMsCsPPjQ+X0xhipjtb5/TrSSJlxohUIRJTYjR9RLzoI
VlIStyGE0V3A37w4W1XIFfM/xK/Mr8pE3AKMl3GAQ9yp/1Y8Ac9RwzatosprIRc7
jTYQSwhMOqFFGcXC5eBsr1JIyvtiVHbR8cY122vo5CQQl0q1R6bJk5p1+jgqXiPt
NvknN+B70OMiRGNBhybxMGgvCf0ZxS2jHDDDGdrM6W6XCtlGMTRFS8Amb0aLinlr
DJc+fNS9hiR2U6NeKPSJlQV03kLtT+yE4S+HY9R7qnUI219ccEUdm0zcwa3HzRPs
oAdz2L2zNd1EzKPq91ZH/FCogB3li7S+nAkDqSg09WMU6+RfaRh4c4mCKG6GBUwZ
8HuB+v/6yrOSq6MJZnnO1d+K3egQVBQJjUZxOdxfiHCItYMDIYKMQDW6ejESim6+
LZbDp6AY17ol0nAFYi6IPG84N0eT3d95X4JgSMIlkGIk/bHznRWYJJUQvpETt9yR
jPtmTW2VqPpNytFvrGMEZbXewSQT3WOGxOO9i2cdUy3XIhgdcnhWsyIjj7Ih0B62
Wi8JjJquXLJ1LSP9jdjxg1SuTXxVJjxVDXUrKCmk9sF6eNa8rAPEbGKcX20+zV20
x4xaT7z7RnALY/8WjQp1+rfl3mdzWyRoTfldBglg2n/r2MBUqeNjgcSQJPVASWhb
ZqJmeESagvrLpM/umJ2f2XcOyTjF3z17/s+zbg2aTT3KmXjav9GNQYt+WAmmUSW9
h8kVo97oEZUCbVynw20fNXbmx12gldsQkpF8MCoNgus=
`protect END_PROTECTED
