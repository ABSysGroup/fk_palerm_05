`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+iZDxmmAN0V1Jm9hHM/Goj/Cm76jTuGkvRAwHttBsSAtgLzrj3ilxVcU45arV6Zv
7IfxLo1NJY24l6pEz3+OboPqdH/1LgQmy5hOWawGGn/sH5eP69HxQqcHqpYFLIH4
KuyQgcEYwq647CuLoV30ntAvG+skaVg4xYvXQNGxsytsUogefJAgwfeCMxm8WhwW
a4OLR9y2DvK7wS+SiRAIknFEgQ6Vl2U0Pz3iSJIpGoJ4tgTHHiL5SlltEhRD4MSp
XKNfIueFYP1oPIr3d3a1nP8n6haQszukd0UXfaSuZAhjOArV500g1+e5q5aXZCg5
uTRfdncymKbK0U00xdSjx7Vmdci0uVabxPMv3ikc/gEt97BoNwXaSwS+9v33Uj+B
rZC9bVq/S9LvMwzJcJZJ7bWtBr4cgU46pKzWo1s5JJiWdX1tNvPF9e+qzo6WraEL
0PEo16o9bp+B9FXufPtQtDMLnTiVUHowoQb1Wa26Vmk/uKBGVkiAjRV4tZfSjwh7
i8kk6XXld1lnW7fUDNatM3l0s2c5KNgddbQuwVOCjsDYDaqG5Q+/6QsY+VE1PU8f
ivZCHsplDq5hK27dAWSNeLxjpqr+k3GX4htKmOD+zjXrUqLRVRLjWoSKeXQCd3UO
pLN1dLEeZUpk9w7vbFbaVKgA1jT5QWUxQjETc1M39R4qeiKoHkBY6VRHJ4RMh4zT
m1ETTXpk/VluAml0cWczZxGSCK+bUSiS7lAP/iVZF7mFYGtsdbP4Ddg2NkaExzxQ
URAm64qMzjRoM9G4fESRZkdgbZ4arraP8F++AjsTTKU=
`protect END_PROTECTED
