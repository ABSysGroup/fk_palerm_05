`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Mz50pMwShbo1xHwdRi1A6hai1VrAngpQHnt+IPSF6tp0aL6llN90euJLpjM0tIX
lwAnrYXXzAWiNAmEe5+Tr1XMUSb2ooFyT7dRjmO/JrCjzTYSKELYqxX50iPEfTHf
WhA0+MPDFbX+/O0Ty1TojukfhluwcIwHi6HmO7S7dLMK0BuO8gWE5oNMBppm1dJS
2g060dTGGqf7WLBtWMmNd9qU2stx/LXN7fuEG4j+I28CH/LNrOcs1GglDVlqvRyy
yaWKzyzfWeYbylcOEuPDa1m3oqzaN2RPFZwoiihMMgFPXFKxH2ihQGPQOtr0M19c
RMSCffvgwd33mTeezLj456U0Jp07GdVDHj2B4j8GppX+V3ijJG/jgsOoFSnTMSOP
UqYgMy+d8vU//Qa1xNwSRbBzOeQYzciydhWbeKJFm28DlNwTk11L+AePaiNbehrs
3TINwwBYXOtJCa2qEMy/F+wkwL82TlOtU0K+cZs6zdXAFQx72kujRUNXK3mUYOk+
UYAVw2M34SzM34UaQpdvJgj0h77KwTMYzguy6GwV0C5uG7mhwJhuhfMqKilv740o
552CwhOFDzpyU25obw5apoDaS/ZoqzZ9ZB3yz0TetHwBdB5l4Em7oi49LkkhcDBV
knYbE+uIGzYzE7d5QiM5ZVzornefxBO5OBfS1Ue9VL8u20hEimuW19Zi/rZA6hMQ
tgCM/gjls86FzstEvqcsYA==
`protect END_PROTECTED
