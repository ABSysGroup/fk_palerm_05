`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8DbXFyBsZcj1kutrYWQphQpb6Y3SrO9ioFILRhV9TrLzf2xiPm6ie1VRg4vDb319
sGhmlfzRB1gBwkHI/sg6CjpXXg5/btRs5OyWDVFFCeyK4V8nYRZKzbt9CDoGwyua
709r13ROVM+SgUM/GIG/Pg1mPawO/HWXZ0SrAwLLChTfJf2ai1pSpElFHdz6HUdZ
C+VVs3r1Ic8aJ5UkXMnlBbIiCO6qr+ZKF2CMSXM0H2WoPQTtuxdnD87yPWj+Czae
drmatUv1Sc7LbfvES1sPi+Cv0m4dliKBAY71+gHYNnVdzcldbsol3vDa9kV+xb3F
NSBKdG72cBeUgISh+8SNVYZ+VduzPFZnqMF2jbxF4b3QTJfwVI7a67/Z7idOtaWF
+i7lIZFsok3CB8QBuWot9mMxh/9jQ3wRyL7LpiXA8o088zy0Ikn36wpOeIba9E7h
HirZbLsjXGvtZaC83Q/gdyhu1yscpX1t4WcMcI1JX+Dj3qn0f9qR1lzAZI4+xnih
P5nwh3P8GQsga1JkcYyWDA==
`protect END_PROTECTED
