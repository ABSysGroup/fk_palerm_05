`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gXiCPker3s0pVGbsW/Y5LyUbN84y0lFFxNj3FBGiWByDK4uYRmWHFE5o5ZJPbBnq
76QdyFw8DVfweoZlhH2bQkyFNKiUXeSOXnPp/yV9vCP+zkfBpzg4lWp/LDsBUdPM
J7IXHq5M1C2/wuntYzRl1tcrI7eBQApSRjPXn/wbZeb2KacIUwM9KSdkWoCMcIFk
vERjsSJFnb+WZWlbbwGYm7BqZXlEb+xcID3R3rrG7aUA2XvYd109GHEQlMIJcHoA
qv7ZFQ0cCh/+HPDoPIUfYPx1K0TOtbtLBCmQqJRKRE9BkolfF0W6Uo/7c/eZ1chk
judh9e7rSEAA+7pTsevl0N8XrMIWdR8XmriRMHOENGKIi9BW5DnydWYfseoRVd8O
i6mub2nVKB1IJSJ2/hVzZXmqlZiWya2CD2MEig2wyXY0m+t22hQZbM/dQu0YC3II
SEt0mxN4SdR7wpZoSdhdQ//JH+cgFWQqGR+TsUFwXcUClgYU2Xh4eidniJ11Nrug
+oy/q1fbihjgxkmjpCAkMznxSHTwEZfRmUw5sRtg4Nyc6vjJv86cm4aydxubmUd8
oJAiisLokKx7Ty5t52ib1RLaXDUUVJnDEkXddFPSXZyyhkZNcVLe1JM65SwgPQhQ
75y58pheQydA5OSaOa9nZueiWFfFDVMuqr0492Fk9oxDFl7vUsLNy6bS9J1h2prA
aypUYMxhNr7GIjOZ0Jq4WXqjZ360lfpO2bZaSyKf00g5OGB+YQKM1oFZrrBqWtMv
9jbEub7BdBjzturBsUq9ZBDqXCBp9m91Oj/xF55XZJjsCZXyQQynTm1XEk1ic6fv
OvHOxo24L5gZxORpmxgPoot9bD9P+hpSVwvdQmGBojzwFrzDdgiWp6pPib3pL4pH
j0cF21n6ZSXTjCmZVx25Mwxmxvhu2R1vQBCMomjmCv6ERyXL9XrwfO1Ojhba5iKr
rNgNb3l1ZWki9WxoTbcBK0PYil21zWcxgeAV58R88Xai3xhoiR3EQUz2wIlQ5tgn
eTZtm1mSxoYREU0WpSUn9x/p8IufStHKYF0p8AuDfmvyR9s2ZCWuC9m3dKw8V8C1
/jNxPno1Q5MKOmeR5XsROKJarGsNQO6ke9/pcdfO048brO1AmLN6tFyilTQWU8Xd
9E+f48geJ4qxMJUPu2g8jRgft7xHQHYtq4GhqzekRJD2aQh+WGGLrvqDYbhxZnIi
kaUxjJSVXkHM7GUbCPFNVQloKVdwJ7YUQYVGLJfs6wnjt7SOPtjXPeI4FZ+PRz2d
lHQXDegXJidwUT5yzFwpOvB8dLU6ZXgbFSigl3jFFOlJHnam79FOtzXtE+SI3qI1
ZGA90nvqvGn8I3JchuskuwXCg6O9Syxtm01dysWZuGkcQqMsoXHMy4cIjRepMg00
kBh0XvoiWQyZJntwOp7yOLqbHIJJP4qOBvuXKtt1PHY=
`protect END_PROTECTED
