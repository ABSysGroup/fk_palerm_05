`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bZG+SjLkpTpCQuSTVt6jkErcFHq/k+vJiSTZ9ttLHW/fqgi6SxE2YUlT/XueG4Jp
E+6ZjLQFe1yIs5/w+KA1zCWfIzQd6Ab7o3CawEn3hsUqCWaxF2f36N2Yo95uebDF
O721WaJ56+jLzP+LMF9sfLBTlKcyjyglLfLnBfdEo/lAG23VbOXp11O1r0zemEhc
WBHkshZWaw7oUzPBwxdjGRKUIkvTCWm3y69OVDqCcn6r57SY0oU9AedKKNRALRmd
aMHrirvvGBRHGXHxu7FwOGIZ96FktQB87grRfmJaB2EF4aVkjDLnJe6Tlh1Cxtxh
ZNJjspM/B4lWJfPua7ccXh81IliAK920b34Vr7UtV3dyCTvgxjsUmUz8+1/mhTud
Nr2l2YT8jKcQNgwByZbwwAw2ic9mKx5jmDK3gzMF7LpTDn3Dc9EDqkOAJ9qMTp3H
7lzICCEcS5J46sZBXFVccP97c53w7nMWcCWSCQyYcHqM7YKJbLK2qxfBkytfKnmS
duXWeCoEZkrwloRjdj1dATkFTK2vI9Ji5rz5NrEcii3H0Z6MkhrvCHzD3Tg6Ydlw
f2tFTswaE2RWej2nxvRSpBCnddiimGjhCvDMkpngB/kI7OfgU4gthf2K7fHE3X4h
ayX51B43BYqYUIvpmrQgZAgUoC7BC9wZ4ngORqhRvY3ao78FNKkougmBWFhroCd2
1xida7HCVDwjYEVNcsV7JlXolUzjYG69JiTVBNg+v7JbofG9Qh0yXFsD+f5r2AjB
NHPMGREsl0067OkcGtDf5vUq2KeTWEoOyg46rrjvmJpACNjuuao2J67BWMSKDrkA
aEFqb35cYXGXoVqCbUaqABEhtn599ulmJLi6lcUrJ8+kfEsCfRf9N7wnHlwLZ0fy
`protect END_PROTECTED
