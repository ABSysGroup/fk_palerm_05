`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qQV/R/qS0XqVRGL8jymlBFce3SGc1u/DF+jAdJgGNUyg5yphh5iTcd/6GafKMNRk
N/h6xAtS+eWJ3jmobCq9Vshrl9jP8PQnYBjvC2vjcNGZ9KLSN7mCpdTVZ0uVz5WC
qFsLKKzlo0TP9YP1bz8s5bYhkUmCPElPAjtc8NDcNoE+kDgnZ4H9Waub4wbZN/uF
zo6CAC+hDwa7+jpIwCv/zqj0Ktx0lZc64Lmd0ivewwEI5Lnc2fa1T6sSrvAA9UBy
Y7+CoLpzIm30y+L1gGMCxYQQ7poeikf7k5xE8FnU00OKxuKdm6dyZWhLLHIZiz6J
8szP41iHGJDODzbAySxiAZkb5QLHM7Toh8Gtg4Sq8lJqpZ89JchkniT3mmo4H79D
GkyrGZx8NV4KzOMWkkeH2hNKSBIQ/KosIPp53/VYtdSBRi+gOWJDfbkeblr+MVMJ
3qNqIZwyWLJ7dbnphuO2n6XLlzVD6KNhlbZ0iRhpohnbOwziPH0k9sFdjiM0ZQH+
8Vjzm0np/L2q4VmREVxgBFgJ8vEIkRH6JtxbnJQAY2ssTtDyBPQCg7JpyCrxUirp
HxRCUwouRngG7s7uQQC0luNA3xWt5Dmh0Bnn4+CJ+9ClfYBsopRXdR0DGApTBkEE
wrFCIKs8izkOrPLspxTwTKerhy7c3BnceqGnI0jy0eFdx0ZUCRL+MZgfHO8GUV/a
YRoiwvOPjFFmEWa100vymUvyMsxFN02E7ozd0fuLHefN0WmcLt1Zi6Ntalgaari2
bKsT/JPzkuZ6rDxb+wvbzBFaB3H3a1FCeFXwYKsEdQK2ckgJ4blhK4QS04/Gx961
lW7FEjvyNZj9QQMYZbPAf78u/9s/jDkuV8S25gqHxIwH1HiO4wTfSVVffIfweh6G
423xFSeFEVZVfJvRUjig2cwF+fwRkKKWgqQNswCPKUaauqb6Bs9/R/ChSrRbZgqT
MU/CbPmsmqZzfQo01wYVnpiKCPrARzspN4xc5NiGBYYNT+ykiQXBRZRVK3pwdM1B
SzcBt6NXwZBUs0ggX2v91wx8VDppjY1xkd2dUD7s3AG/RzB0tKb8hF2jS6gLyw0Z
bEbrrUt2dfR8SmfRayBOWyi3IE0UxN2rfDUHYDs8wg19Cwa/28Los37XvMqO5LcQ
`protect END_PROTECTED
