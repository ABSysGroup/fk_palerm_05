`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
URyUiWDahzeDRPKcS85WIU2aBcQqsv/SoLhl2D725pCSVPugl0+78djsNGGQb3d9
VzoDK6lb8dcEO2JLySbzYi2xpZxkbtaRGgxmXAwHxF3QGf2CddcFqRcFMdb8+5TB
UgJXpuvJ9WyMQP3QzXet8sxVmj9i64Kx/upf9Eh/qhNneF35jEa8NueY/zuFMKPF
zEZBrHe2O/EVUGEa1VVj7AsOTO9AzboQ6TKCthYUT5mmLll7QeHqjfMkWpRq67Hl
lfPVHZjDd/yVxOdJjiyDf7C+pJZqtnxSjb705Y2P13/Z9Ig8vXQQ2Mxd1h0iOo3E
UHyjvykF3NwkrIhBmLfzn8y7rk+wKVzs0uJyeoDt+AJQqpDr+nHwTgUsns8OFuQE
z0ernBG9Gwdq3vGjSECfBSfW/EeqtIbYYJuq4qGPI3/F/djHacytx+dGsb64Iyhm
1N0h+qpspyE+lfjF+rfnIiuNZLbSP11Qy6QJxnR6vQU=
`protect END_PROTECTED
