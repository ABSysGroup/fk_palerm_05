`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LkI5NpEWTzf1b4UUB2qWN64D9QVsYphWX9/4i1AubT50uTGnXH7vXUlIydZW0WnD
vaGjALJ8NeM4JOAtRDvHBDhHUTZGO0e0MvoTa0rtkdWDUeFefyraL1zpCDhaOMLZ
tX5dTtFzLeSv3ScfrBrKw5r99XfvoIbEr1aOgq8bnGle0v4rXlV/Xa3/Zs4NbzxC
viPZN53SMVsIYB+TfKmZ8+Q7Nc7ngKkH6UpgzsJR4bluYkVCJ7k5Toj/A/Ovc8JU
ujUvT9L/jQhxuljC63NL9s2GkcwEvHWwVdg6B82g5NKBgH6XHyUT1A1Ir/EDw+pN
UEhEaV7e8ASL9YKu2H37Lw==
`protect END_PROTECTED
