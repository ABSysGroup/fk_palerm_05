`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Qos+postoZzGAjNkGVsCqok10eLki4pVRm5xUhUZ0X6U8Tj+8NcDuAj30NISq6P
GoF7pCglo7PDH+1iEgZMmrxPRv4MXzZyZcehwLvJo4GD6NZHCcGwa0pW7AR/ONnV
UG6n4S9gmQuh3za42kCLGIBVi0teMIpWdBj+CnqnK6A4FofPUuFlONyTOfyR+h/6
CFzJaVcGFnkQVcltdb5XAaAsvHsI4O7WTFc4Rrr3D7p7A717U2OcOpGdW5fiWylG
`protect END_PROTECTED
