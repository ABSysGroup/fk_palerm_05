`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N6qqDZqYVpQI/1YMQNlMPD6JT3u2tP6y+mZNXjyYuO2ViAKPWjlMxPl24/Lh4UkI
al2JamrJK0aWQVltYvJEauLJOYjuxxyyXB24nFW1Fjz+R/yqnWwOWPVavj68zZac
X8jAHZHcDiDueM3KQTa2owWwtRUnqYnWAhtiv+LVF0ZNx2OORD+YDk1/qui79ZQm
Z32eLjlV3dhjhRV5iTnTOEiaHHrbtb1VgcsaMadMEwmJ/WSk3yXSMZwKTDyPjT53
ARBQqj+7sAyDLQmVCrDtWPysi0gNoFFwPbO6CS3dXO41AMdH3n3hi4AvXqFRhROf
pA/8z2mo5Nspl+1wk+pwfyc7yPLCe7+5t4vcW/BRU8EQaI9DraQ1Mfl+qhLSAwMm
nZbRy8YJ5WbnFF8kahGC6Rp5ZhMyMhodubkP5wqAkFzWWVIFKBpqWfRhKleH1baE
2kUsVr9su/rE8G6iZrS8oNRDc8ign4ZgRzmCDJBLyBOh0L7nyBfbujcwVVwdBM+j
LwuJCuv+UvAXABLk8JqzPiVozO3rKdgXZt96xsBKgsApm/aYBE/cHK1pC0alMEL1
yxNd8v9hCG1VXV+OrTKSOji7RmsD2gy2Gw4Xg8PLRSXXQu9Thl+faF3JjU3zjFJv
IHF+nSz8PvAcrUb5xfKrqeQybBtv4oCkjwk4+z7xv4Db+EvqGKu7zkP9LX3wZMwy
i6sRji1pq2Lv65U1EXUxVg==
`protect END_PROTECTED
