`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PZ8JOLAtXtqQi7gqul3nLBPlDcy+MIY1QUKUN0QgvgLaLRd42G592Ms/GvDF9+PF
+DV/hvGIfzpRd7tujtuf2zvlk2y3jp0aGbD01hDtkznH/aiX8RHhVWHbcw35rU7U
8Lj3w0ois+zeHC+ebEvgKWXa0Han/uo/pFGkyQhCUBYjYaxY+DzspRAAXH9J1lRR
7hZbjCs3yzGgSi/o17NLn+IzHamHoinWepjlEdwo5odHkpc8RiSeWibu3Ak3zxxV
DHQhdtHKgqurrOXf+NLyXiNsXded3V6XPCebHRAM7yaQ+0k96RY8cdSLVSgKqijw
aOT4FchntiB0aOsMyLnrk5Fa7APwGZjU4XsRCD/mmrHD2zRZLBWgd9MwfDePlwWn
rsOYlPOETDeKGKN1TFG5mknVS4W1jCI/pwe57WhCO90cVFGvCQwSIddyRutev7GN
RIP5bDNaY8sPxPpBEVrXkb3VIv5fTZB1BwO/st1L39X0OKdvOYq1WZzHtzm+FSxF
pDVvH/9Y1TruBo9mAw9Tqa9p15EjMCs53gL3UPBS78A++aqUUCl8pBz1hwwtPF8p
PZvMm0gSXO7q8c7/2o/K6um+UxOABgk74GjlNs9baHTPPScwd7/daMxNhL4gS+It
hO96ae7/Z9inW44rPklWMgYixKZbd1k0cM009GgHF/LJG0hOBHraVKQG1EZEMRga
CzYIB8z8afCMd9nDe+062LcoltS6OG9QWdMTg+THjwBOPjl0/1OloaFO1VgJAJmZ
3Ly5gJ9WxtkfqJ/oKd4kn/8M+j5DabNre7/mRWqjDntisZCcYTl3IQVQ9mmyQBwr
R3NSXUD0K4pFXgwjvwkTiLoYbM3sjmbvgD/prm5edu3+Bju69iRMzcjSrVXBch55
JEG0L1bGsROCpyRe/ULYYg==
`protect END_PROTECTED
