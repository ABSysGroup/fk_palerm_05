`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/t2EfhJe2EgPZQMdVML4JcCnQeH6NIMAO3EUD3qQ883MyZLxWg4fCOC2z8xml7Da
DTTs86Lg96Js5U51PcAkoSFQO8fqLlJI6+xpmb0TYP3bLNJtG+sWdU7Vqrknl6c6
bzqC1yl/aWFgTvMZtnAK/NQXsHVENg8vvH+VhznJwKPX66xEYTW7k0dBC/84iBxo
u7KfFJHv/f8rQIkSY34sg3/ugma7b+n6vrISqIDjZR1cAEBuSmszaSUjZ8T6ZjwG
LQCsxDoVaR2yHcJna25THU6zVqtbvalSB4BxXBb655srq7hTcyTpDPmTSQ1La43S
/AiiOi+Aom6Z9qceMe4EQApqRTAvQPEc+JVsqoa3eHmhQWoGPVKjTaG9nZjFcmFm
ytOu/yGADMXUlQCa9CnHn83udGpoXMBx6SCfRh2tyvvV4vomPBHs1rev1AEtBPwv
VISywxkrGH4W6uZdeaiSiT9O5es4I91xDPFZ8tDHHqG2LweyPik7uEkwQ1Y4Lq+n
W9NGsui2STGp654iG/Fo2YVf9MES7udGQaE5h90TQIeQl55gRqTweJ4xzRaoDFpm
UcsrnDd5YPhIvOBGLNQ407zP4olvUUJPQ9LaExH5ztumNn7xLrA95szQ+7lnIQzE
Bu6ZQUBk4/UtontR6z05umKVBPoRXO70mgMNciKTou3XatMea990lHsh4kj+9jP7
sZPSqLHR1YLIUvw+U1NQvoszg0QSbnOJnFzT+TZmptFi4fKrAPGS2HU2BWSgO5ZN
uk30C8ncj+HVAGwUKY4Mk4bqDXcIm+EQhRL9e4yQOemgDQ+olPspB0oZRnE7lLzS
5vOtecaY9Uwh8UrWmSOXiJ9iPMHa/k8QPd4GjfNyqD/lLOXBnEceQmrAiaoChp0t
03hB0nZplZp8s5Z5mfaUwoCflrjWhwCySXCAOnVIIE+LYB5IfGWR/DaykOPRNWAU
Y/BsdxfQnHS9kc/du2oidvEmCsP3Kl4E+NnznRNZasgmVud4sRQMJTOI0ZBaEfi5
Q5IfvJAmb9KZIToO06jSopqYH0haL/FJpvwPGzSlJVCP4EmkS/yHiGa6QR/fhnCK
Tj/tWEhoJ7xkGmHnrwgROaHUnObhVm5/kwaixmJlKKISim7ATpcasQEFfrV9eXc5
dte+u0xH8ni6s2KNpuy0AICAdT8w/URD0zu5bxCPqqTrbn+hp5SvOtpbIpe/JDv4
gfdEXYoxwLChhvO47Ku9arAlKzYZTSNddGoyQxFVo1e1x/mmxTbtvPeVXoU/cxhM
jwmLXJnBCKulnKz//uQb0R/6ZHNcum7WOm1HEfnCVL9J2UyH9MR3oNccJq5yL9UY
ETcBTPsLpYOIpKXUfG6//QQ29W+GSwJlHWz1KN4wJE+SisO1mVsksAcD8As0xgki
ApAGI4ZSQxQoS8SdJ7FKDcK4s/DLximbuHMOEzmSWdW74S+KjD3AKgypWdF7a20E
t0zzagd4msjAAd3AceRk8P1y2qZNLF2S5vQe6qo4GwnhqXh8MOo9dYPSbIZi6pbY
IEaGERVioFMCar799hIPcfsG2f3rAFf4XzjgGnAHWtyNIHDCtyR8Bh68ynL66KiM
6/aQcUfWZpNUs9I+KsCzVbhNYE8oBSxjbgUimcxAIr4DKHoLadIJQ5OOQ9UO5TfX
JtWQQOTVMIy112i986XOnovuuV2NW5W9lDqUR1eaARL7cVdxu53mf4QK90Dr7LFx
Z0L5sAn0Q9hAlQqhm2839gT7mVe056apJtigEYRKS1jGNAWcDsk4Vqcn+z4z+nLo
5UG2ykrsK8tmt6uZqssQtv9b/a6xSSFDSnXWRzSgUFu55uCfVm1rOSbhLmmQgsFx
hO6/wKxLvJv2xZDL6YSvwwknbNPAtY/qycospD+GIP3C0bwD2an7XGkPTOrY6XFg
k1sw+VnUeu9t6mcCRGFFEItAdkNET315IDmf86qwOC4KGNg6+NbXj57Nb/LtQmzR
jcwolr3sAsiiygwkGKZ+iKAg91s9ROmiFIhnv5VrpImV5BXbzbEAb6lnHjIwsa46
ej5BbiG6F7g9g5ClL93DH9Tl+C/gWc08dj4mp0apPTzRRFDufPVstOEX8Zvn+Ilo
huHLjK1NpMbmxvjmv75zjbD0RFGanaa/p6eUOI1MfT8bVEGW+jfa5hWC0KLtdYC3
RGtfDWJ2gOKid2bgrYFo6NsJjp+/Z2FT54Di475R3JJwyfY5E4Sk7r9fw0GZE+5W
FAk7Zkf27mlGNLYpcDVHQaYufvSSCcuWfdBgGrW17e0kSH2zgJpF2kt9HIA9xOdG
LK3/kj4UBvA7XA4LQS1m/PE2AjHkX4cQyZz/KTUSWE8yflmg9Cf1AeBpg8tLZtHv
qQGER2UC3YTKY7epl01C0urB0qHtBS4J7olaZvofIaicVxtnU3qL1Ca+kCa2gK1D
0m6jRsucyhd7ZEseBP8rLb7VpTlTc/Uj1T7RPajeDgu4w/H9/Htt/o7KIWYvqP8Q
XwH4hQsrF71tzk3FJpUv6iu+NHOGzakP5y/AyajyzY1930X2a4ZgzuX6Nco5NfJf
wuvBbkChf/ptSvrpqRhX14FqGC78RjBmW51muRitzefu+Lt1oc2bAbrhSkJmkwHm
yu5OkBIOJyXLwJDravbNYaBy1OZK2S/HYlT5YQvmmiOogUY4ofwSSa1FCBz/vnj0
wCZb3MR8CQuGfISC7BHIhND/+3jLCErbEKwUXGkO9DA9c8fjeyQa0CT+CgTUMdt3
WsKrUVDzqhVpHRqmBtbk2KVyCZsg96rBFKVi1vcJeSBWE4RnqvHN6qLGpQrN1BJL
ahXN7b4N9T1W98vvFW0+Nvc2Z9AXzSgnVY39g657p7ydHiWUHxxBFIATpFSiwyOa
uyDKiBRbzU1sJYsAH2DOmBfOOtHO25QE+rvB9JcMyOmfZ+gr09nxuf/qybOg+T5P
Sa10uerxI1mHa9ztJx6WVvUI7pJjzy7Tq9qX0pRFdXDGzW+nyKvwTHYr93Wyc441
C4veTwwUp4RsDPXIXG7mD6byTE4Ak5XGoQi7G4ycL9Bq6X0CBLmwaEHY+ERfbnIx
Ayw5PJjsY7RmDb+XbUmZ0B54h0tFULpAOdZ2ZQDQRYSfpMY+m8l8NUxDLutPH58B
/vOnfqi99w00SGsm0Ih4mCF/QxRlDX/XPYDLqsy4qdvpl+5MtemwN8x1H/j8zglT
5oP4k8yo1X4Xy7DG9ZmE7ndAN4AAwwmMoEWIhDh05trYTygNeYfYOMb0JHvRbizt
uTiS01H/ewLYci/ekq05sU5Agz0BpvfbU6efszMIm8ULpx+KIxqrXhNeLMiAP4gr
/GTTRdjXq4D1qcxthkRi7amJ86yxLnXdbaSjVRpLZ++FjgqyQ6OfZAY1pwq8G2E9
QH1YFWCXEIgYfo6Z58t2o2X4l1sx1RDKOalyZs+z1wmVlIhrKa4m8vwZ9KYBcc0s
rX0L+gWe87gFlTE0XrI7LMfmVOtRMMCAE0lOMeTb1Gjp8QMaBW23SFwTl379iKUs
6t7xXV+EHQU4bpE5TKb04KHjof1gNTe9PWXG+jMbER3Tv4VTjxeocqLPAuYokws4
HRtskb7nrdTVAFe1AmkNs9vrtsmx1vZhiPItX0JsqyPJMikgrWUw0J0Ee/r+Jquq
i2SFdiMh7UKnqVmVjgWhdAqpXEymphehY/oZSMdegALobx+g9RUVL4pLECVB/knY
L4hPI0C0vEGieTTdOxA4Pja2yUAHRSDtayh8Jts/LnUbbRkg2y+RzHK/HbXIvuXI
kedl61l4MJNIFoFNuuUfl2atVDD7N2aEo8ykA6OtN2RVqYSADmX3rvOpxgufUma4
ADtfYvV32YT3PFdAn4YR4pq2zFCTokMGilkiuWpTIe22aPO7GoUbdG6OFwSinbVG
JPubjuvoIYUaB7IcgMLaMjPVN60TmecEgnZR08hRDYQS9J1SaFC2uZbQ7o7/FRLj
rQ5cDodSMO7/XFzn5iH0d70ZTlNXkFHQWQ3qGOesS++n0Rx3mU6xQCkltzdISuH2
rxiK64azq/Y47nQ6Cd4dR0BbyKexK/Po5kP/4I48hz/Ti4cMpY5ZcJtKgVNSkoVN
0bntYNISDTEke8C0/EmNtAoEY6iWB9yLwW0tFSvNc5sCsEDvh+RCF901Aqcqt6/T
Pld4E5UXC3foDs7jF00s5VCvN0YSCpg6PtuWarzHOL/UpBBysuhHD/FldnLRN8XH
QJkuvLGZCRreMVPkQPlncodJV0yQBJMDQ7wIXRCjEzU00kQzgFr4cD7FcuDDftJE
1eX0jlJknyii0o3SzBFtleAHnJ3rnppjKw51S9Yf/0Q9yL94atRmgyzcIw4hxbRP
M0z4+HDjM9op+/TrIxd0SlUGiT2GHHulEAeeKSyW1Lwm/CsHc/bjB2j6l7bll+BG
VnN0lxtNVxBvVjGfmal/G/PVJjlaNj2XLS2Z5teZmsx2qGQzVTWFEPIGObEZELdg
D/FeOTel/RIPjPtqLT3rlA6mVmqm4cqQRI96I6irNIl95/wJT2RaBRHGGiYLHH79
84t3qqvgkNx1t+FBxGN1gd9YbSXEcP4mD22MAIF3wrZv/hqyqbyoiX6/p8pO8Mo2
s208mbBkwHHkf1ddiqxXxkwpgXdefMzPCb3tPxekcLcm8wEJxsLpHGyP4Q8SxAUT
8flfVk8uaK8JVQEJjuLhyB2Lam5nGXaHytBlCUpuxM7qKcRdp+fWkV28dHNMvUzO
aq9eJZovQQNjGUwYxyvAlSo/r5fpxZnUiomwVtLzBRGMxklCXEAEsB0UISQd4W4m
LBxdWyJ4W5Q93clpnarz8Nfj6aXlKlW0tUQdSCdpR0ErpqN41T2x8iYaPrIXsH3h
FHLwm3HwOLEweRTZlIxtsYwYMNmiqbZg4tWNfKQb5fif3Y+CkLwWDJ4QethVeuQ7
oW295quh6cSLuOLxXQX8MWhd9CiJVAI3NZiMvy0PxK4Qo5011lJ8AMc9OHFNrzMY
Ur1RjIcW3Sm9ti1UtpovVsbNVxNEk15vkxFlIvzGYhDrzUnB8r5NkwMp/PFeTRuZ
MkRgRu8IOxULTR2u9IKsCRPsPI7raPOioHNdqD9j3J59WPw6G+hVqyv7Nr0LM01U
8Lw08TfsHOFEFz2C6VioZm+VadNW7+KoGK5C8BCqTfP7drLxVRbw+lBNjydY7MaR
+4WsmZZ372PunKaohvzlsggLuq/Kxf2FNWDfCXHwavjqzAkyMmt6iMBCmwYZCLfF
l9iKZbv4qRHPTXKcQ8MUFt8wzWRSTJ5KawzUobdX54s+teMr4vxfhdtOCVIfl3uA
DAY2S7TXX69G6ycTkPlRpSQPLdAbpGOq/zyR2lb2+6MywQN2sFV5qzuoV6fr76Eq
YN7idt8YII+SJyRLyX3cSs3+2QorXrKgyzbRTpFg0YEb2StIjohV0rKTwwdU/QCy
TwEbWtu1gdR49QqpGfUEeFQEy0DNqyqbAo/xXp26UL56v9kUaXsl72MajiU9ympw
sU0Ovp7NQT+kyYmsC1+vXLAuLJpYjLbsNyeTuLT0ZCFYzYzpgX+3X5Y5m6087biK
eFcx2r/13r3cv/xGn9l1ohqURqi2/vnCLnYAeIp2Ewo45ZVRmhfFHKfBHZAL044b
euye7iLqOQjc8uLXZ5ub6/pu9kCYJ9oONSvE5T5p2Yykqq3E4MVJGIm0W9aatjZx
Hnz4lahe+8AWUVEIrbC0OvdCJO3fIk0h30VGcJwjwzMGD+LjCeYGlbT+y3Tum+Ve
OR6/8g99hFy6Hm9zbxGqaTDfcg42dNbNy8FKygTuZb+VNLar+ZQSfA1W8sfcGqOG
zKcQV+GH528pCL20PhqZ3rU+8Rpe3YWXzx7YJsDVPBREd5vP4E1oFotROBYwnSoa
qNbHCEy9FGJyEb1GaqYDjrxOrgVno6NY/GJY0vmrejoBTE9rExnBMxns4AYFqorX
Qb52rMKvvcNNjq+UkbxMkMducA1h2xrT9/uLg+cevQezNRESVgDyqx4PxYzp3jN4
3Vn4caeIYlBU+tzHhe3BAkGOROT2Q39VkmeFfXzbb6xoS6R6i/O3fj20n4wtXNqs
Je7Vi1T55wPYkItqsZPJ5OFB17s1/cqgNQm/4mZx5lU92zMGJBfCNW/Uz47BwzPq
Mnb6LGYlCNLEb4FDkl+8JTVvC4GnuPU7pgKSLBqWQ+xNZHJi/POUOK0fUrtMmdB8
4UBU1Q7FqhecZ1Y8sW3JrVGqV2AQRI0AIOdFUBiXvT5rXNvkhSzMPW6u/b6vx0vk
il+a2HYnuFt74HH/ej9F/h/gugNpJHhvwn4R1Wu+YnG3+Q4uw6POa8gqDotF0Q0/
v8tI1yprFvNiqSchVJrALpl9RVAjp3DXRqxHI9PVDatxvTE1+orZ15t//zJy8FAN
/lkgLvFqpLlOlaGcbA+94pvlNAyznexj0j4z/KnavJo7ZZSXIu9SsnMbhd1z9aru
DHKBg87pgH6DZ/9gbItrYncSNRq38rkJ4VN28i8AjbfWZXVE9okujuwGFm0oCsvz
sRykaavnAuXBBdhjbzqk0w3uTe6OLOEtdEovJu3sIxN0VK2fJmXLM9Ig6ksMIoOT
c9NtzMr3wIVSDRPjH8/Iy88M6Jsag3xa6g4IBwGi42Pu1Ecsw/7o8LRx5lXs2x+7
0jmj/9HBKsq8mVTTqUz6xM5dqruzs07prBok76wQzBi2Us4jIBsdzbHIfbNtbC1J
8133BwVCClRnx0aEnnJk9iFCset1oI2mXygccmjVVD93WAFibDuPqCM7y63iKvpU
GNNPJ9Qjx+en+1QLDJdbq9YS4H9xHAVZJGwrS6kGF4szVZ8IHA3GNmmbC3fT5qAS
0j7w+IViYwr6nyuK94jqyRh6sOVYeWuqJytY7QAJvzjHrKJoMay/nJeEAm8xl4iS
9cvxvKY5b3/VDRID0QsEAcU1fMs4Fv+m4st4g6k0+lf5EJGq9A+0rsv+WEM+9m/t
6ibosa4TL5DCqpDfhku+uaOLOkwaLWIy/7XmAmRAC1cM3JTr79k0ulh6+YoPwUD2
pMIQkdGYgyQmtHNKsH5BJ6zT9dIs4f7ICu4DIVEJfXxOpHcnG76IYJnW7b9sFgbU
lmAwQWTKgCWgzW76csGuPorshMxdnYsZs+8tLUufoeZdfqot5TMsFGHl2tTVMJeu
4zx9iqzwmRTSpUcQmzdPvAWz6v7EIEp1oxGa+f0tf/rLtQn8OK2gZAyFaik1LQgM
RvL7jmIaE8k1y7evvelGD2T8u/N7bxmcDq9y2MvCTz9+fnyZLsZeoyjT2RqnpJ3A
rgjpvarW7yabpJLMMGGNnOyW78J0NWW2pT/bb7ZFh7PdPGnxgNr9Ut+pDdl7QpvQ
uFwIvPPV0g4StWWgtCG4We90VKkDYKOMzjHl3wBSmOJzYIm4Ai1BAFdYLb7Y044O
LS0228B6jSIG37d/UT5Ijw9hdE4Ewil8c3dJfqGjnZGWdwCGy+nNhFAuSXhq1rnE
46pugzroGi/5vF0lz4+WOMLjSCBEwavjBTQvtnqTkOKQG2YvKqR9LF4dWqOLDrd5
+ZuCfHvJ+UuvQBACcl2Ki5lCZ0mkqv962THoXG65cHh1MwmgUWgH/y1EBC7FpTm1
KsiNO45TAfp8ASdBdvuKotxoOT5lW7fMcKRVrjLB3YQPF0iSC8uGzDhfQR1Wij4l
+2CtinfuR6+HadTBbfls3rKSLOP5o6GJsBSP7/qy+AN+Qhu1kIglnqiiKfjKqu08
9Da+ql64xF52IJAfE4sbSWppjM+OsZWwDzh3Ne2OEG/dP/wdtLyYzX+iL7N9QFNM
19F3pJq7JRq84Yfifl4KlqJRkcWPR6dIOI+9F5qhBlN5UwcBCP/syh2j1522as1W
wqGWeRC4c3dV8bEgyTNGTXpaAI45hbzXJYRvVTMnQsrqm+iJWOT6wmIqoVR6jtxP
a6f6maDjAC6gv06J8s9fUJE2smKzFQyxklaEIADNB/yzOHER8yEL/Iy7zp1Ggsin
CEH1Es8Ugpbw99Xfa+aarweld0BuuZ5BQK0fwM7cA9fZ35pEMl2lMotwVhxRBGYx
DEW4+SvUVOI0Xzrcny1nvQ9KqIUzprD9/QR7ap1F09rVi2/Aio9dgPm26rYcb4ON
mDRXXk0zcNAHE3zPOgGW+jWI1xG8fGztXQdGeasnJvOTM7BB7lOXB7+bXq02PQ4U
TVouSstCbtmLU9ibNzW3rjYBYjCx38zAt77HEe91rt49iWNnmlc+FXboDT3/PZmR
393YSjShQXkIQAXqrifQjUqaiHMdFzqZeoWB0J2K5hVzXg+K3wk1VTDR3Iw7LG6z
a2QNekAzcOLGeBm6cpcygBnQV63cI3n62v4UnxgFi0l+RA1R37aToiOwOeM4AJLh
fqgE1GPt8MM9uIXXKisicM0a8OEJpvMrbj8WDwtd3Mn1cT3Xt6uKiyJvKJxvFk2z
aBIBcOICWUrNr9ExkhBc1vTGsDa3sljvWfVwPKhP/gvgmRWhMBE2WRCtdPl8MiXy
VKbMGkBeRgOL1pttb/5lZjE/ycpzKpaP3EfpeXFu8eaDW9uo64gXH2cRDcEoUy/T
CCxyr7vYHkaxQ2+MvBxoEzOeBdtSnjTrwCqAos9T2Ej1nkJKtFkRTzZyU0WAxRe8
pFCG9EeLdj8e7vT/j0vxfD75gxsPZweIc0pG/12/+mOoN1il0VJgRbP6AEzZp4dN
aiHoTmPt4SNWiWuOl7up0fCdV2GU/9qfrPi+o486guftwMArpKSDW406bbdwNLO1
5qEnHbyPPWtzRo6RkG43gLrJ3CYQ/Ab/s//zhTac/511hSd9yhtD8MAyuO2urZlW
qLzVa5oAg0CbrM8iUeW/dtziCDOgDn4d7lvQaswfpNWxJcVSVfZ3/rXC5W9QuXVw
KNG960zoB1s5ltmcpL7Db2wQ2bLNUApdpqFSLUnNEatb28R+R+tT8jgfP8kRaO1c
0oLMJY3HOVHiYWLqb8DYPNj++WTqbqXN34enmdxu2z8/Io8L0rB10So7PbuyqtLd
0ekMhA6RO6GWWVOotdr34nJIiz+jHmY3wqxGAMiecOFAImwbBy4GbFbayoQAUr/m
GS7dgQCHfqQz/TB3ih+Etn0Z/isx1Vkx6anW5SkVf+H5YsS4HruCN3Nz1g54U0VB
f2kdGxbHZHw/DEhjXPKJvNRtAYg0B+mjYSi8xiVEXLV+6GbcQwOycs1zhMqouXAg
DSFU5oKElRvj2v7g2fClb5kE2G7HTeFCKB1tL+pYL81C/iecUbJhZgtQfcfSGKQZ
DQLSPxJw+Z9L6kRbwgn/3DAR7lyreEfWXHITQFiJVhoYf5j9sU94dV8I7fPkC6Jo
JGJg71ZJutmuQLQLjWdW8e+3UukYF9mmG/WvS+ffrhwcNDU/ihM/ZIZvu9CU7We4
ngHpgOfF42yxolyJbHom1JScgNNdPHjOMkPVEpUXACRMXRoIWNXh0fWIQw+V7fhY
Fe6q37VqRBCPJupfv1/T4BkO+sZ7GIzq0Ut97+w7f1NTG2zB48VxI1x7dN9VUWwN
lR0CNEOv+3aiQakSQ733IvT+xf/3pBus0SucpjHhM6rNh91Oalq7vEPv/1rVXM9+
vBDAbK7XmyMoBZ4niZ7A5ggQtDNQ1vQwbd9L6aKRBilWgZUuV1BMoaVQUiQnfx3l
S4XSBY3k8UkAUdwhzI2TJZmlZJ9BLZIt0oL3wR5JhwaTuzE/B3XtLPDJolxdQv2t
7yupmAcpCE5p7PrkgWHA7Qe6yICP8Jh1hbygS6iWZEZcFV8Qx1fgzndSBuDzbNE3
J0aUNyomxgw5Cdx4iOLUTH1k2OkhmVhcc2xIAnwqbPeJi9Ob1cXptYeXYTKwVvfD
52k57ChAv7Y3qfdDNwyvr7JdgOgXnpJ3tUorgFcqJEBoYiDPp98YddV9ARrZ9eb3
i6E5BN2OKLXDEbaBkdcTaHAEz7zqLCtUMzySHg3U+QvJkaa9QaVcQZcgOxGVrsIS
LIZUX0k9pe9vCs23U+r5+DNJp42QbgIHG3dNhDh6RyT+HrrDnN8zcpAzPAOfvxM0
h3QLckq1KW7KZqyZGECnogUZ3sKNBUlF6LMsoOPhRvK8Gq/1rTaByReH7p3lfBwD
h+NMRsuk2SGUgycgFI2kLoA/hvFVGVlo1GM5chyMzHapJpSmON9Qxdn5+bDoSJFu
INoJcgnvKd51cntKigC3OkDkTlXDfSHqfVGYvM/RntQIiPunleTxgKhB8P9b/RVa
Jl6X8R7r/cf415fngg9IHBNh0so8kd+8WqopeLKEM9ni+XJZNZectuOWcw/DcM+c
NAQVRil6dVTCWjBx9TgLR8sHUuk4rSow5fYmY57E+1/XV7jGGKTSTE4ICvm1PAZs
sRaV2IZk0DjP9PCcPhBBlLEDjw73QsoTFF3Q6QdoOhxwNmOUl6B2iW1zE6BT0HKh
F70ESBaKJXuNnh/YYLkQXsuFy8svWGIr4j0zQOfKUrRR4b982hDreoY4+XLrxbCU
NatINVc7/KTm2QTomiJkcbah/J2wO/D5KnTG4Y/32ANizhfAEHRBKWP7w9XtZivm
PayMKswiQ7SvIgdz9zDmuTIlOlLuKr8Y6glPlPb8xpmOXApqZwKYaDuG3xFlifvH
RAotsUEDIUBdqO4ssmE9cdVXMbBPCdSOKUM26qtN3L//jSvb4yobNulOy+WjzFKV
GtEvL+1EEq5RMP98NAqUjokaKyQSscIWCaAd766Sm5BlTz18oZe2NLp+j4a0geTw
NSk1Ex5w3UHJ2JhWa0Fd/3/eaMEC5OOG8nNhudWr3F+VTSE7pg7M/+m7OKK3XKm1
oejXP1bIFAZWFG/h11o5CuXj9O6NqSk5j5l0BzQL3dT9WMOlwjDLwNccoPLF6gxb
Lg0uk79jEFkVSD1MYOYOH0MMQKsxO80SkYNFVDiNO5LxmRAtmeVYqBrjLtPE4PX1
tl6IuwbomLwx1LiZCiQCDbWHxWrQfVaU52jiv8JQ+KqB1to4uwPzLkpVx0zT+g9P
K1tmUyksb9bJVwDow29QxsakreDt9bf2nLKp8muIh0zG+YsLplEvCU4HzU8b/vbp
ZXIAxesErkgkH3ab/YOrjEoRmv7Ux7+83y3x5xQRmchTTddQOl0+jkITR7LhFW7Q
DIl2b7BysSBOKGHJWzP3pkDkX2x8pEAZdX7MZqfQY+bJBCS7dmLjrmZ5HfErxdWr
XfdRCSQxDP0ddmbhr+v9gEeFTxpijs9PCmOj13MaNzPQAwwEZqeqzYnJD+FnSWwo
rO86XrUOe+zwG7pYlDzXdmAXwkJE2K80L+ThzjftShdFGLrJRbx/2DtEWzQUKX5a
FcRXErsPnMQ3muT9J0AieTS4DdLf5gmF3RN4TrsGOdhbRNrrWLsyMpvRKVUneohT
9AmlXe7YidqNDF3eIBxUdMltkwmC+8Yyhsv1N4arge3fVWNxGXfDxjfx6VNw95ZL
Zy/XFHeyDPR6J5aU1G5k4bGyAYfQxbcEgnXDo/G6i4bNOWuk0N/sgz5byFVKXlfi
/0kRcBbUxsdpAMZD7yUVHBm+eMZyLtYrVWCPdBszVVDF4647wMZ4rW+3iXWbMjza
m/UFvlutoJWLpSQkBJSZAN0uJF7PzKISow9LR2uETrslgned7mN2VfK6owQjxmlD
NCm+pOaK2Rd2MsJ1f2VvVbEZUjcxhzSFIySc7BguabQyI/1tTJm75i/1kfnu/lmV
9X4oyAWiy7j42MXHdlLO3w8zZzB3iiA4Zojr5oj8IMQcSHXic1QdR8KB4IWYR8Kl
gdCeELjhH6/IjaRDmAdcuwtlw4vQrthcNhngkaCjMLfuPC58HcZXO+F46/nlV5YA
LoBlneuWyIyxu67yydSr03F/q6lRtfoWv3sTa+jvq8h4o1EhNqq5IfcTVlDtrpsC
KTEdG/jQ/E7EOXRcqfJdDXRDjHW2+Z1tX7Cj3MyIay5wgymzAsnBhwKGNG6d+CSl
Ufmp9s5p/sve4OK86IkT0cGPY1ZdSsg0jkUmcbxc3Gi/sl476NKfNOHUEKR2ZuDZ
Gbb61N42ypvIZboOz0nayZZ1hYb7G9yoV75TlrjRC3IjX/C2noJkRArFv50YaDnN
jB4rlZA6PRNmbK+9Lgp6a4EMWebHJQDk17g8FmagzRTQ6WiF/JhUVsBc1rOwSNe7
fYcLJHZgBDWCXBb78eGYakgavDNxeHB8+pdzgBeBXSoHR7VOmc99JAQLnGA5W3iV
zTbLwYzvW/8I4q0bA8t9AxyxVbLwctTDuka9OhS6oDYKYtPgPKCWjwshOYFqrclV
mMpUHv2faoTrktp1DTs1RdraL9h/slwxgUf9GhSxaZBrxhFpu0Z01+0am6+uyvjj
YdL4OYin8LNMRwIGNRgigmhL03nLX6VQ35yTLs8YnXcxh4HWnOiyI8HAKaVSGiWy
dXxvJjp99t1joGNg8lmK2CXcMDHYD8Oxsue1aFHJf/U1x5kd5gYwANcQ1T/zsRmp
LJDSgwKFE+rEhhp8AWxCv1se2gPeG6nS2NF+eyi7YWqarLof9o4c+bi26rNOTeXY
3XlmtgxtdLIzFf7w3jefa18qevTnnP1SMlell7z0DR96QFIdN54sZjvrKdoyFYP5
NWNz9PDCywDxaVj7UNAf6RgKeXK1cZ0mo+2B/7TRQJox3iBmf+1AaOEpsD34kOU6
rg50DTGytdvyjeTk2ZU7rfKvRv028PEKCBPdxm4KQpcSLQOz+FHkCSu8wjJTVFT4
h6v4d2TvTBCie2tfM9EOnGobeNULaHg/P/XYOlppNI6mGILr4IO8Uvkj+8RV9xhY
d8cYnSNyxyGW41gw7fSTlSBMnwgTIulSISgtEHpqkhhPAGLrBHzJ+0MZf/d4E7jg
ZxgjhxaHhE6PRVNeWf/gMN6Ej/Yc2a9VPbPREdxLFidrhPZ6yZ9sRYE0aDwnJQsi
UFUkqBDWEbjyDKdzhIX6hSkrj99dMBNbn9phMF6kKF88wEphDsri0iyjRIwHQx4X
8A+0y3rIwzntZc870KwjwT200IATZFNTiwu8XcxpyNQbXLYn/0Je1D0OTzK//Te+
SMKT5uFU1w60M8GG3OypG5v0G9NYx5g8S4pmE9+w5WRg2Zq2Y27xVVWs5wh+G/Xg
eq5yC2NkrkGW7NIU9GHawCFKQGgyTJcUh+Dpg7Z+qcx3dM5ufQbXcBigRRO8VVmM
qbDJH2zZZBgXUBRE1vTtmtNtEO8Ga7jevWJNjPEaH0STQl8TCKZpAzAIiqP+y9EB
m2txoNte9nkYOpwnr/vYPq+ykiy0ZuMbLoOUslMfNU5x4xBvNXDSFrFNBff8ZvdZ
j9RJQF6ZIiR0J+UF6JucrCQaV9hB4QLeP9JdAq8V+77IjomkZIWeE5Ss0azbKE1P
M/8BBdAnD8O99tkX2b13LHBUAbVcHs9NLh12sYtJDTRdT5eC3TdZZ4O6avWM+/Tn
b7JLHkeZ8DMe8xrYZbOjH8QUR4cL+Lrla9MrmQpb+vVWPJS2Nq2dCgnHcEDAZwtI
nfdD6CsVWBsCq9myXxUBjuUNVT4na8IdpuTarEJLF7E05o7ZzKhrIqMCQ4IvllMx
F1DU4+Wrnl10ldy2JMzwR36P5TpWw6X6BRthkxs+rIaIqP+exBt0PWfIFiRREULj
bC67NfbLcP+I16aibOtJEg==
`protect END_PROTECTED
