`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mPLhrfFHsG/yVnyQILyUm12cFbfxdJtp+dGU1ILW/BphmMKXwT2Uh8pr2LLDx926
sAXJYJqSI1Pm1TcDOXwSDo+glkEfwRJtacnYOnAI/LvROOF6Fj+rN0Yqe+EZiTX/
JWQsScN+gDK+Nnd/gcedS0y1qLbS2gdD+TnRhyYvDQdExCPfVVoPmPUjEKEeliQ5
ja5ayxwXezLc+geV4jw7Q/lGdrQt2zDQ21n+iUdUebgDzbf6I0ptRbmMxh23eHPb
h6yuXlJC6J70H7s4kaOTJHgGbM8aFBpQ7VW67rVSqIajmnuPABjYhdburyTuq+6V
CBJ2a5aIGVx/VfwVDgDb/SCVdwHwjzq+xpFAZjMcv33HmemMZud5QsG8ZQUdb0L/
e3EHvEtsgYxJqFdc3RmQPrYmLOrjjyPhYpFrJMebhKLMfv5rnpnqySRoa8l8MBEC
SAQo5i8ZNAwz03kme6+wAq+Zj5RqDcVfV0LLYW03z29HEvwzEXw7NNgZd/B2ukw2
`protect END_PROTECTED
