`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7mO4JIR6Ur8nsLd6DL+cLPiqIPvmOOZD7r1m+n/tNim5T915no2lKV5TgCR0lCj3
S1bp80/LoYJFqG7pZReYDGjgO/UKSy4V7zfP63EQ+EIYVNmivUWSg2QYRGVct4vK
FAf2vehpHTW7rezNMB9l6rnQo1D6snI+yJfHQpa7LccU7x0Ci29QNa5awx2uo6bZ
PP2dYC/+EOSkZOMDIWf6U/QIXemVu5I3r18JuRaNZcbwQNfOkON1qqZIsKHB9DnD
2Ruffx+D5ngP7DZVEDMNY2R4kn8rlaJrj6KhG73Vm2PF0HovUA57AfDaB7UDS9pp
iYz1aZ2s/N/H4qB8s7nxQ82mHd3JojuYa/P7gdTpO9ogKQEZFq1GzBQZkwZZtqEH
/KDbtdF7RmhQlA4voaDZSKOFxPdCdMKKqfF23dzU5J4rsssnt6ZPyprmsLGY9vr/
Hvn1K9CrwJHxdHWSfwUh2o6vzTrOYZkRxNdh6L9aN/LA5oNdVN+ASvvK3COWeZWJ
uBnXAzlMmeZKcf40FgA+6vLOGuRF5mtrxtmFkFx66wt1+Jj8jbpytqD9p6F17f3n
ayxwfesZoqXhkodqzF5WHW3t8qKYUQAJl5DY4hoS6mdA/RCw9KyPkEnoZ0phn3sJ
6xdcDuKtOLi9GXKSVVHxwd1EycGlbkYbbRsPVgePwM6SJlUuUoNhkJBk1YdzJV+F
IvhVYUPwKi4NQXnBrG3/VLpJC4QIRmuS4o0fb5TIP9Cq1Kn7cQN8qKq45r57S+gq
PVv1OXEj6eFx0AQOI+ZqjjH9pX/ODBdYMBgDnDGOcZ6qZBmh741iatgAaHrg69u0
4FrsIjuZVaRdXXb+dC73GXbpIm7piBRJFzsr5czYymaFyy5GkeHJWd7CQp6LDu6K
oRLf27W4RdNEctbEdrZERh3x8HIL8oC/HJv+hzGJtnjDb2RUGKj1hPSYJle+sEyC
uSxlubV2vL/OIcGFaWWjqVm3Sk0Uvi/ipoUi3yHyPyNPgXigEZqlRLrGe+iRu1Tb
0Ih+uuTM/JfK3wvczT8+0ZgzHIwD1T4WRYTjKBxDAH58M0lBd1dugZoMSZ9sN4AO
cXI7UxOfJjUZx1fG8FtQxw==
`protect END_PROTECTED
