`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h/RDIYpgPuOe0Vu0Go+JVOE3jNxYx0I/EGo7+MTLr074GotKuRkn3qRRj5TTgiqY
+OOJGNbS1wuL4icadmU14yYTRqM897ZPRYLMrolbtyZ8oZNmEHt+AoVbuivu5YMr
THE7SRFSQIOd2uONmwOYVYS31+wClBGj5v2hOZD9ikEjBpcWsfIsOsxTGhmerhbP
0PHptOgcoRK3Oo7baHCpGZMJuz66lB3UZeM8fu1xbhc+O0MtOb4dAz0qUls9L/xL
2H39Ty24wtWH8wefWzQe2+WtjjrAIdARdQXup/VF3OPLqPSZQaluCxv5tgV9QQTb
uYXkfeW0ZpDYy6CcxOWZkzEcSZdSFDsTnFsWaR65rPxkaW+uSh8iwzV96KdKdteg
eMFjsXcR1KDeB8YVvcWyrTDRREHdT41OnEhfTZWk/VOK5tEvq5reNC7894cNn8oN
9K7Q3XcDCpkCx3WdXs862vh5kt/SAO8it4Z3gO3D4qRSYf3shsHJu28SirxIMhzP
kaWNq1j6ZJQVVzUcHwnX4QjyYFJnZ3BcAiLEHQ6cDMOtkyyzITDDFF3hA5h9UEXU
0qrOQdQbUmTJ1Q621SiDTQ==
`protect END_PROTECTED
