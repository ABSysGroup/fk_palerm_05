`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uWNEKdZEMrbpREYKZJ2k4EZOv8KldHD9Dc5tIU+RYLVvCZIJoTH6M3ZHRxwwRGxJ
2ulqyXNAJw/CWFYfbxpVqRR/ewlng7/2YaIltumh8ProThtceatq0h5VbB3z0Ek5
EfYm/ZiEl8Q/bc793rS8BBEwp6jaIInYKWJozsxieC+EA5mmGwq/W7TvmX7lFhDp
TatyB4+AycVn0BaVv+6NzF1zZBxVsLLFSEGXjHk/pGu9ICEkZv95LfOADSMKbBdU
rvpPnswX9Xc9NdlrSFoYflqBgpoXraao7bIr2Pi6zROqBnx2Ex/U+K4FVmN/fGgL
MgpcXNd4hEF0w7fctczsv19WT+y7KQJ2GoY/fIha3ev7jpUqpLhiJ5Koi7iB298X
/9HuedH1K9gikZs30CYJxytbz642/+2SIxg7jOkFC2G6V+Pw4iPvAxUoZi78BwI5
wQfM+YmCyPORavrXMGTIlaAa7PdQmp6viW+KEOf4qvbn2BYlfEO8UOT1EgpxPW9D
7R+K8/r5DP0n7OeSCwv+VJsnS9/fKm5BuStv5t9vokg=
`protect END_PROTECTED
