`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P8B6BTCxMEez9gXqVgUcb0iULc+Cc4ep0f7p58rkEZTo+4PUY9eivwsl6nUSPk4V
YW0BXMCVMII66sRFZQiTGxWHKjXe1GdfRiEHC2pVh/6aoTL9YQH+FK5aBYi0J3t9
IKKCXHtkax/0NEDHTlDyn7Qx8uCKxqzJ/XKIr294KBXrlXaIf3qqfU7lLlVNCQBR
vKeUQi7VklSVzLTBSv61vG9shrYc9xE6xgNregYLUopMmKOpWtoeeQp9uhYtQTLY
czH7gVmK8HNtOob/sYlvIVg/upNIcaz0piv9jEB5jY3F+uLr6gWaWVwa0gqHiSUz
G/ad+Z3/V4XWKJMtA9KlIPxZGr7j95seBmZi5o4Iu3U0ZfsTqOrKqEudj8/GnsH4
DAjRAk9LxAQxKwoAs5UK5NBtcSTmfJ7jVDgC9p1KhKCKFEckbWpTcKCZjs8PhUOx
UcYhyaMaUFfHnIgY5LBjOFs2xBxg6nTvYSwMDrgTfc0DtHemAu1eqvTkidzPvLga
oa92lHRCQvdtr5LXNtu87pDMoHtEyi+O8s28NXbzHKxDpVHWLLIciCB94wmKgs48
AdhDe50HxU5cgWuu0USPDjeeTMJ9TEdEQf8q5IOzNqADFQHcPvdPz3goVxkpT0j9
MJ7MrA0l1dxJ55WwwKcGUiS/lw9/6DmOpZAXU9vS1PLR7FwAl1o4W7wPBqm3c5SX
dscjf2VibPp/gSMGDGQScD8fsqubE2lkJFR+bX3d+y784MrQJF4RiywFEVIvwJIa
iKxii5wZhE8NKBwVCSrkovxvb8IN6wf+D3cy70KixlDIW/gmd1z7U7pmwPdSffOx
KuUg0geQKRUSclpRCdf0aUuj0ulspok0AilEVPDTwhHGzbgHPmI+nRVpvqZngfjz
dZHhjtYhkaED01tE8vOVv5Cff32ULB7jwMQvsLqEfsZw9HnB1Ir8Jgj/Sc/ByEp+
`protect END_PROTECTED
