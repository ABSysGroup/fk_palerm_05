`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H4Gsbr8vU8ljqeQo2etlCmroaCAaKLXLYAlkWIPSIpKrDQMErxwNhSBwm8wQWj6A
NcMVkgYeCX8AS9fYUFnLffNDs2IAE+bJQfApICEZ9qAfOiFqDjK/3le7Xpq/yd06
BKBWz2mtQQbnuiARBRN2CeQ4xDAwNh/qH5DskcZ3qpe/BBc+6gLxO7IEmhvwJJAe
tcein38nHWyqemshazTNSt0nq58TweuHi+TLc1nDOmetKR1k9viPTH0MWs7gaZlq
BNjbuE0GVDTIBpRUjxnt4wfySSDyg6ixMVbtDIrn9a6ylxfqis1Sb9KMm/HoKGkf
/M8rYIDzKhS77M0Ai3cqRnegt0eIhZwD4oPIzp2iZkIfxUdu9SXDScB81ZfWqwG4
zAuCpI5fbuuR1kZ8KpTQxCv7ZK6n7wcPpbIM9fRMkq2BhqJWgYHJoHwuI+puFTnJ
CKznRxu95yCgfNHv3g3goG7xWD/9nnFbdoJEj7hD27i5irCNc0cq238SQZ2DymPp
naz93h+MKbTq6R/RB0kWo5UAP9xgsYjCWAfQMuqY6hA3aO2J3jic3k2kQCXJNCe+
gqT6VAmbkDKpX//rcXkxNPidfRcnxFMgcotPvVBhCKLs9Fxec6lbwK/yLnE2UuaH
n1JmIxOf2fQEu1VYBrcs0vVvdqLzCbVAcN7wsre0bEwZTfsBIVlpS1sevVXh/PPw
Uj7c78kOqhBADHm/qzsQGa0tRzmI0PqFoagmdgXhhE8ebsc51Lp9Ad6E/EqJifAh
TkIhRopyYfY4v4sZzdifqE+8y7M2w6NXa0nsL3/F5akRupYbfT8Ans/IcMKx1Di7
rN8fhudOgl2+xckvnp5dH1X3JYmoWe7crxZjR12bMfwEZ1EVnbsli9FBg8mpusDx
qgne5yst+sRCKd8H6F/1bLsyZFSMcea22U/0ZUg5wma5OjAnmnZYsx6VYL7PjN5Q
T01UU9dDrpu4/8rqf1rHhiEk5KmUVOB4Rfl6k9OI2SIf5qZzx1oBIBVzb7+sHisN
MqO9Y7vq7ScwaHAppsXnx4VebTaCdO2hSKQU5kt3SOeAwsMeZQY4EoUA95rm7IWg
IRlDwyurHgvl+Z6js2/ByqV8Vy8TsHvJKwMDdmpvExw9HKGjO5MthXQ7v8yqKoPo
sgtgwqCTrhydFkUd9j7UB09lpWKGhpw05hrd5pNBjMLZoqCU0zFI53b++tUCeW3k
i/14OY3KnhKc6d0mbCsWHSBBsCh5L/lcX2sOtOnrsbwgBlc+5yw7rijdTXGDW8rZ
31V2TISqCsoVvQz+J5KikR2xCPfm5jMeOlePq8UQd/wHtxOeefaM5JA03+BLBXEd
CMBW1AlGLioLl/3MWiuFhOECa+XCKPddZ2V6W9m/qhOgngW6HmEcbvinVpa2zVx5
AJwUaC2Q1u9e0z3opS44zQKb2QqgZyDmFT4F68qo4kBoWZUF81nhkCpoZsHb/spl
Ce7tmfOkV5nFaHGEpul+abs+S47mvgJq96NX+XSXwamK7mBUE6zKHRfX8DnYYKBX
tpkvxhGfGu3XZTBGoviucOKTTHt17zpZE6SXv5BykORti+t34uEpaJQ3Hx/ptnTa
ljZKC/DpqNTo91tznUyqtAq98CluzVT0+F83LCJVpnwaoPPfFSxgI6UbhoBTOW3G
VL3wLh6nCntbSUkwAwKdigoUQq/Fy5utsQeSFKxyW9YnZ1iMJfnHVzU9x+5H1dzh
pEH5i6H7349nYI5ouX3cI0tDvorkXQIVRmNf1LdqMeXgiAMNZqPkrkjy8CZBSVCW
rU6DNHj6ES4UPJdTwsx397QdJuSBr2H0kKyvlSaEOn7IiVWfDq4efhwDtMFr/HeU
CALKlxpxoK59/HWwpF5CPIZg5UGhLtyi5ILhmwd93iSbWKqWgzEif/Y8pBvKQqDK
Y41Tj2nhLxGHPDy+64jVOSr1BqzvKBOoOvf0SNbGyjc6T11ycNHKbJu/ngHO9Ivo
2c0Sg2D5llq2PRmaVO4/T2szlmpzd3p869l8p/9cp1XIZB/wmZ8OoMeDVgpjdFGi
O2IERnOPllk9b6etL0wLjSrzxNbXvg5lb0pzdKxnfmTFYgJUktCzEUD0dgQ6KnKF
PdklP/VpU0YBQZ6Dj6KIFUCZNVfkNqAapTFdpl7tQJ5KIG7HN3ElY0QCs6MBhN6B
AbcJiwfORzi1SelP12DV6yrD3GR/omTkNyT4dWUNup/IDbwhwdOchgLdJ0XVDhoX
NWdxAherrr6/20n7dh/cnMpqldIqOeiiKdSE/c7Uyt83zOe/XhIBGPWnfnokvj6E
BKYfYgOGr4KXzcyr3lFbe2E5t/mPoiVfxV7YLwKhK0cU9XOGov1X+j3hU6ZVOgvM
YIwDkH/RxWipd0STLlQjuQLqanwxDcuG6HwhjYYZQaIojBnDFOuFoaCyvc+iPWJf
GZDBARv3Ru2C3zXsjMmGgWeS+E+pdigbgxHgOE9CQdnNALXVHgdHGC5xXiHjAg4k
7vP88BBymjIbvygRdupQ67VW40GKyIewMicL6Ita6dOI4t83u2MgwSad9CRKBolg
A5+r+KLt7QCgJifH2XtzHgGE/xyYybTcKBEnGOqCuqq+mvOVgPOpd/5SaSkr9pYz
E1i9xYOuYVV3rIKt769dnvyVhiAApW9wiWass6Z0Totub7YfHxcYvCh+9JubdiNT
pO2cRUFqpPM3GTY+gKfpfvzsx+V4RE7QyT1BrvsfJ1rQCWFruHwEy+0XR5Qa1Xi1
sP8bNNxMxn9XmmFchFWLusUqjbGGAb/hTGurvRJDzbKWgZWa+8N1fm2+65nNH07r
MLo7/3k2LFXAcNw1yEkb/FNh7FGbWqiPX2QUOdm4jF7j6cbY5lILoui6YiAxHdbg
8PkMLBYKE+AXyDGzrQ7HPqwfM4RSkO6J7WU8s1MH1M0PczuSWg0MGexVpEDcEUcZ
12HIgH5rE8/esxSk9vX+UkV94I14m0tqvJTd7fNhtmfwT6koWz0jsHIJyAVlDjX/
ubkbHo7jd7DXQ8JMeBKk0jQBg/mS2MBZndN4UWIpKEB1KU/QAMxPXmdnmcqlcXZX
1oiFHxfx1Svdzvaru2usi/ltkFHSajWJ9rA8UpaBWPBeKglHkCP00bsRWGMmeD+1
6jBeXU8wyIzSMMx/hgtU5ueal8mupqVfSczK7zfa+aPPwRuo75A8vlSIWL4vx/3I
HJj0fhpNCsEuZkVG5Hj7CgNHFJYV1DfAbcKgDcvFsBW2UVGgNZDpFxKKPm2eBzX6
ze00XMOfw9xtuMtMgInipaDOKeEqZsMcVkcR1WeXLEsw1qvhm/1Ngf8PxZpZKAaz
GiiZHv/IDcO3SgKu/uxzL3neLbco1HFMejT73cKNm7ylyEp9eUQvkHB3Iinr1sME
tP9ejtcLrY99Qhsy/HTcwucgfDQOrQ097cB4dBK7cavzqZC4mXm8Fv0YpXvbdd8y
MOlOmL91dnkdc3hGhT16tx3AY+xNs8LW6Z4GTsq3curCJWtPHeUkGfEpl0tz7B3X
cJODKIj3MTc6yuhodtKMYptOObY5VT8E3s3FecJfJycSsJwVBcpXstErMYy5je1P
H15XVXuKJn7zDgBgQzUVW9M5slgGrz6cmBfQl5fL7VgTkXfmnAT/ogGbPoBH1UmL
J+ZiMpXdDWQWEVZ+2oVzRbIRUyO7ra73mqX9bINAK29KZkHJ/AgCRHZa6Id9Je6N
L0hBshvyxBpMvE6iBjj1wPOYJoGppuwSbSY3e3QHI00G5TP1mm4A0eC5u/FS8AQr
rTO2kQW/y/1eDQ0v1fD/C4m4/7pGw3alOOmT/ux+moEhIUecVHFjexHtE5X9eX2r
oIrFTHnEiOEcY5MATeGP3mUa01G2y2tm6giseFOvn5eKE0W8f0tQ1YviLblHYkD4
njNvyovcqcG2qEE9OPp9Yp1kSbZZJOJyDAEUdVDpDXyx63B5kvCtFXj2PR52kedv
azCIQAc/dkQwlLzltaeHUND4Ek0UZ/GQqstXABDz9hfRKjKNVTW8E2cvaiNhrS3N
pw4pO2LmMlYooyl5GWgV+sZVWzZjlG1tfCDRSdR55t4oowiY+LOtMxggts3KL8Sd
kJfkZCG33ijDU6c5Mte8TyYqaNLLB3cK/2TMnX+xMXHZWCJyGJT0LVGXdkzFyD1p
iwjjrsoJ8QOxzkF7D9gUnR92VZ+u8q/vO7XbrJp69Df1HoOitBbagzGrb9GW41Ij
9BXX8BCX4NY4xlny6s+ZydPtUqbvrQ88taIvZYUIlnJEf8L6NCrDqYn+DciVZHrf
z6uWmLo7CkoIFaNNerfNDhVq5Vt94D2CyRs7Qsqs8wScgrR6Ez7t1I+MBS5k39iQ
GGS5jNQQX7jmHDYXXB1mzXGFiiwdJGWG0Q7R8e2Q27C0OHcu8DV75kRwYhGASFoE
06Vf8EsNtGHsXS94fNEUHbF8IBJWe2TtLlmnyDSHM56k3drme6Gn8j7chGquvafs
9LS6THVA7n6UInS1+0IczcL4GFVCrD5JHQqQ2gP96aNLunqEAZ9T1B0QgHm0nN1c
YSSuJrQdk8jt6th2uqilNzzV7lhjqAb5UH4cdVM3E2x1WWJahIgjUypNDrAe0PF5
0p21BGwV88/jRC7WKMccIFogcNV/ENznui4Y8Un+qAJnJFXH9Vj7lsVhsxK19O98
CbCFeJb8rtNLPXiggB/t1vo7UWANTH0n7FL68dbuKSCD56bovx6mRyvUHPoWG6K9
E9Q6n8UqY95ra/f4FzNYaCredsmW1uyZTCe9XlXquXGx1K0AR/ieTryVzxW3kguT
6a8kjpHLNShTkvbkTCMnpJZIDeDW/zrwv14jXNu9I8QGtwH4lCBXGPoJSI2xtLTD
KxSICJi7HQ0cJvVlyag/kiAGDQpRqPUd7UaNNykX40htJN/nsR7zQJkCbzSWisAo
OZQfudAvw4vJ2i0IRmIKFB1O9oHr3TOzPSarayELbE3oE8SVNLDQ2RGJTnMNVGNl
nNIMb/d/yWPDGt/33Gh5cEcPq3Phn6KDjXem4oNZGeicH38JEPfcyyforA42zJGx
1wgb8jnsiDWjq29XVTyl4w==
`protect END_PROTECTED
