`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EC75LAD18dNjb7dlkHqT+xKO6zZaxWVBT28ubYz6riwse3BIPrJqCbRMNMKpcRGL
1KqiVVqPgCdUoKNhjoohzjwGIaWb2wzxuoOfgZv61gESTOgFrrgOK0BArdmxpRoZ
WV6P+ggTD5FMG5smUWtcR8UaVtY/o/cCotBMzgb2+kuArS/6X0JUoXizu3fOB2QW
yjRj8p/czmCSF+mhJnZkttGOBI+e+lUxCpgwELaSaDU9YQt8egekw7LX28Po+OSF
vYYDjcYdNsttbUUcFUQSKXPfBYqGbBDbmwNCX8p5bMXvuQAE8PigUxGK5J0cT/3B
sPsLpHqocuxGsYZ9aNh8mw==
`protect END_PROTECTED
