`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xKd6P0bH/k4a1uFHlMmFlYViXoQX2ZgZH2HCFKMFe0XnX+jkRfiJuvKucrZLaXly
eopnT7d80SE7weHyrV7LzBdmBNi3ncxLE6K/4Oi+GrblUdMNxWkfLGGGKHd0IGdN
+nlu/3ptBKd+fuJrIqLXkztNcAT4a3dBrmVqEte8kRoe0eaKhVMtbE3m9a/1Smyc
6Xxpl1oyxDrWXUWl51SM9UCys9yirKmrWzZ+eTNPcL3F07kGTeCb8qRNi7XssW9n
WAY62KMLcrdMqKB/uvKiNlvLkbF1M4HRNDHy5v+lRkxkQHbnJCVhB9uLsuPLuaJ+
THACPsl2a9Igf54x6E3IUPG5z+xcuNfluAkzcDb+z2jsJCVbtfyLa2m6vDXVseZ4
7aV8e4w/FHXX+Oa4uEdiIyjtjx7FXh6gJZv5xJJG97v262mUdy3A/PovNjqVds3B
6cr2Jx2DRpWA7dvPkTXUzV/mhCJ3yYF2PiPM7AYDbeeycpMtOHv3u6oU4ad5S4+P
OclVEGmHQ2o7RbHmgiWP9nioTC/7B08KcgPcV/lpd4JCax6S5v3BiS5L4qrY8lBD
9J/AtBB1jdiUWuvvyXy3yEVsZPrGJurU4I2YOpiX4U2Jsv7k7UMkt78Uo+5NBYlb
ioCvlzNXD+wTeRaz1CRsp8OuFRg355LlrrJzKozQExioc+1EcDfo5lRIVgmG+teL
x5UbTTWHR7xGsdRsljNvTjmC8StTR5Ejrgl9zKQZYbqffLmGRCfNgvQ1VGW1jt0d
IhR/uB0gZJ9Pu/hZIyCjAp1EYQtGmW6l15pibURg9XcS6uvWei1o0ypcu3z/2YZy
ieOl8t0i41UADBdYFDRQY1aU2s60e3hCALXtdvIo2x6QrhsJEMEYiieaW7Ww5sE6
LR2s2PoVwDj1w1LWOhcfyQ==
`protect END_PROTECTED
