`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TibTUX1OAd8euPrbNmu633l+oKYrBiaDnylFj2KAsoNoPF2pF8NUYtwTO3ncJsZn
8x7sZvM/EmPakJIG0b627OsNv8VXgMcIeggNANjG1OUpkArblMZo6/YIXliPLSdd
25Y3yZxiKq9zGeJV8lIdAD+6D/mxgEhVyImORFZfWehEwoP6yoHCPGq0hC/Msd4l
coU0oYr8OOW6qcZnCJ2fao1fauByrN7YKZw2L5HYIofUN1asEhKRFLJusvnhDFKi
sr2k7D6Ll7kMREdNSzVROQ==
`protect END_PROTECTED
