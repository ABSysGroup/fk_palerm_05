`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jW1daq/hBAUez2ebRaVwpiAD9FnwQgxp6JBGT22pMjkns6vb7IxplxhCxAbnIGRi
h114tjv4yvHzWWZem8e++dVIlJUhiea3noY/xiC0OxWnPo4bwJSw7y8yOvr22Iwk
jf7SGKGmH52ULfm4LWVMnR56rfXaxqrXPZXGAu9mlIrjVueZ6JNFhwnm4sRUeGeW
wcI3fpIlAMOJ16xe7IHCM4T5zOAL8Bhx8Wep4RefshCS3gE6bhgwSoN/xxyyjFM7
D5g09Hyp9qDQIyNQGcPwCFi2yAtvutn81QPCv36upTRs8uGnh5NREaOQR+G5AklY
JMyQ47vcRoPYW2gx55e2PsVJ5ERdFvRSn+SPx13Cxz3nAGN2oyyC/csUi6+Z18vI
7neaCZVokPQRYdTmy/qfqHyXGxXrY7abohT9RfAxVDw239TjiWa8bEqnLg92mJhx
gIx7sVzBvsQjxaZjfqjcxkP/TVEL+9AC6MWoET9XXYLnARKgP63LXjmLGINm8hKg
QvQowPoqX3FLxnIn7BxSPDQb1+bV6qCZVjKoOv88g8+PdccKSVVFCgNLBCnAe+Fu
cO7zdvm1rJAbVMWEia4z4HYxh1G7k4ws7LMKXQDQ4Po+Zn9DvpQz9M9ixsXGk/Cm
PyDPlpW1RdfoZTS3NHAaBDc6WmjfqvBv25qqezhpBqUPkq2LUrAgge7CZsFtcEeB
0Eodb+aNIFTZxBl39D1KRl9nTqJJiROIkHDjnIRg3qJQG/AJcpYOJZCXV5xz3/LF
EE20MYs7aU96hMtGvmM8KMML6pwmank3YlI0wzaWFtplZj9yCt3BRuHrfAFjclNg
lyWEczCt05qEcPu0AuctxCTYuIeMNoL8Bhx0fXtcmL3nq+LGDiwbYf8X+bXb/1bw
xNfgVy9oEDVju5AdVJ1RcOIBv86KTjX29MUSdtq8FlXEJrFwbeWRND8p0NUJazJr
PT0yngsj/7p2Z2JzmUiUfniM2ttN9W5gLv0fmwRR75QDoXnZ4IBXY2U1ZHQ/T6hN
mYFwQu75/kJhyKbt3MTE4FmZ6cln/PV4AZShDU1eXr7umYsZvykhBipXrqv2+1eR
hvywWo7dN8hGT+H/eHrstyIwtGohfCN9Ak2eKZd29FBgGWQc8vCfAHtfaniq3NpM
A3IWx4dorfyNtL/tTZHKvBVAz0x2+l46/WA7Hv8NSW05S4kNrBCgPgFhTe/BA1Er
ruenGSHKG23RIbj1qThCYQIuKbf/vLECnWdXrnNF8YIYlCbThOFpl/u+8TZwKX4F
bgDrX9HbEI3P1Toeg+s9A1bC5KTiBML3B8+uoOsHN5/H5UrN9HFFRPaiO+sW/kyt
CxoSvvTJuCENVEwD/nIIE9klne2l2tZw1BDF5QN7z2BtwWzQY7WJzwcM2uYSPZBz
IqrCObVjB/y8gV3IngclfXdu8qy8COTAVSKJUffpPS8iT6azGFzKiy/bdtzUd9Gg
zsGpLG/7ohw0DbafZ/gJQe3Egm6S2Th2fb4YWgSl+sanD3hEb/f3J5GtYU9KkZ8s
JHoPmoFuOYPn79IiL39wUClt33u+2xiYqddWA3yRogId43K63p5p+B/cSndwi/hP
b4h2YH8Vo7l9P67peLyXYF4dGxrao+FnZJONRKUuEjw+TiyIJf3+ius+g+sQ3fND
GcJ5rmp3Rqx6eUU9LNk2dX8NNRaIR6jDosqoaTSiNT1ftuZqEvyWTfby80kbyuMI
+XRWjwKiJHQXGyNQ86o5mWJRd3sCTSJ3DwTZwOk6r4s6BCwHSHy2H9x1Z8tXCQWG
xGEGzYu1FXW99qLHBPZ+qO+HElKL67tJXGaYErVSyhngR84NAoHOLtIk5GoEzyXH
SzOAi5/i49gDEWHa1E2TfFHLeDi2L2gd96wpCWG5nuM5BkxTUNU0Y/bcXz9Z3Knq
gzp3CGpr5dvLTaWB8KR/F4lZkHomDBMy/0yc2BGzAvvSLIbQBzjSBuMnbsFsuSw0
l50fI9YI1z3H7TkmS4PnZ5a1TNU7Z5guXoShOuw2V5slJoE0nkGRZBDXNYQEvbsC
kt+EgB/3lxc8R/zY02eMyVF9p7WEyPmU3juXDrhRaRXCR6ohwV633gaKgin9O8gj
k++EXtwOoqfntU8l2+EreDUTkR+sRl3s5ubg4RGjyxaE5qo6gEeL0zcQXYb8W9Cq
qZ2rF+w+iDbQ0L0f0YmrXRtarSfmyM/dnoxRLeRyz9q6UfXj/c7c19QtTZlMGdmW
QSvxop35jb4x2v/k9hJaJCKxa960bjyUI5WOxrn0sM6PfyrrQfiYJPYCC2PD8hON
RO4w9N4Utmvdku+MMFqXT++E3INOD0VEszTTRilJ27rs8twbd0XmpnsoC/CNY1NP
breRXL2ihANsn9LFdZolsTsJjWkW9DFPYudQG7Qzci42d/oSpdabw40uSOamVGbi
zxmtMlx7ZwgOCmnvDRKlFgl/h+iYI/R9ytA9tI0duFqZZ9owgFT06BxUKK/VYnOf
vAgamdOif+SKA+iEKRgR8iMzrgfSgDtyBIbsvMuuDqEY5dLo0yCKgStAUEEOM6t6
PiOxZ0PGukUD9XblxnvKlAx20RpLszqtWrHymPhZ2PmSd36BcihzWfN5aE17xkwN
JPQcxEmRG+5dW8DvBNl/78IMLv/rJOM/od9+nsICvE8zMG4srnkyCHV6teLTLe3O
GuKa0NjlI3TwBDkYZTgBvw==
`protect END_PROTECTED
