`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ylz1pJp/qPZtaRsGGftGRBpYXkjSWaUgtjiLstCk07ORCAUwkRdSzG+9QxnN5ZS8
0v1eXf0ncUh9dcNvRXJJhgkY0xo6cjEDiC8ePxbeydF1GYtp/FYmwvSb5D0gmYei
QZmtpA0MY0ttzNgJvoJ9U6IGMA7Ra/sWhKVF0X6hGg4NBGWmSnk86VOvXVFQ+Qi2
VgUAdBPeb+M66SvhCX+SkB6Tee+fb5mmBP8haMrP4VEO3tSqD4e/29PKUutDnt5R
`protect END_PROTECTED
