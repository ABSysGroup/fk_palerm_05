`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uUXOUHZiPUoyqsW2rFdtZnsV2CAf8cyxUKd2Bal+Nkd9CIbnMbBr4/nlApH6L/RB
2ut7v3nS2ElcMDjzUMfJwCyAACe3kA/hDxWVLx0zRjozwZmb3ukJ9dflzQasgwTi
wwTVKcUTEZoXFYRUueFNTspxzNjhtmjveR5rRBuonIF2F7BU1onXSH2WOlXnxTqj
C2Z18AEnEf0ihGx324RvpoJ1fCyvBdyRsvGQ1FZVmnvJ2sRToozKOAYfxpeyXY7z
2MfEC84lkgb9qAFZ0fnunus8Ciw9Nz65LdwtOmzRmh005hj3jjcc8hNK6tSjiGE3
DQGLoFyIDEUjAukL0VoJp/tIdXck89wiEurb0Kv0Vy7Jv4JJ3QVj64lbOEjhNXri
YlabKankbjlK8k5VGVSalTnjHMhr6mhOmGv1gICq+9/6aqJQwziQRyo2p/G2Qg2l
kUAZ1oK4zQtmfKyV1UiY5WfCWLgffbMDTkyJrPfsE/GBZyHhvOVT4nVEWSXfXask
mAa0srIuO0Q2395yrmH7I0x3FTPguyMynzw2J8bFbLvHgOW3cUSNWVX9ZKS1MN8J
GKne/diw15jeM6Kb6vC4HarBmyb5x6Y3MtT7fjZXLfhOVJTmN31eLnWTJlxusjL+
GpAuHYf0nFd0oYClQtDx7oQecJhsbOcQxYoyGXBOkYkEAz5ac2BetjWziDeXLpVO
pEH1uGirmFBlkPqdU8rE3m4q8fxG0R2qPKX8iCzmY76yXVedOLJUnL8QYCfRv92s
fR/9ONdJIvjzQal2FCpHFGLpcNMa8sA3jIwb/fgw/6AsBZF0X3xOcPGtTUjsSMZO
0LIe0mTOtKuRqbu3MC1pZRrsToJHw8u9/hG+Ia+qjSkCp217xMH3SRDdDFWNKsCy
OumqKd/m2NOH4MKcMT32dz2dyzDRQzggkB4E3Sss9dHSXv4YpMcwE8M/Zi+9Zhhn
gCBCXLtecNCLbNLfpd76xIAUClq9ArX0JPXBK2+Da9NZmKg9HoIlKu0ZzL2fFIg9
iBb+YuXXCBRbU/6fhsDIhjmC3E3y9fAueZxJDUHiAwdchlsKl+e1HUawd/IGcpFs
UFuCIVkdpBbijjweZ2lixOEik/CxPkGxpcwpYOxx4B/UG9Z0KMuAxHBYNh72C4DN
cHWKO5l63ZlwPnUCS3fn2EpHuJDaMgUXszpSvLP5qDT2BJyBoU08TmVN7hYwdIPw
6+O5mUN64B2ocJiI1JteiGSrbESzxur5b/eihuP70ct5+Wdxsx1fX5963Ngy/3Vs
iHXsZGCrP3qvhiw9zE48h0kKIBj/MIPBLCz/qdufiSsATig7ehEGub/rdmpg38kc
B+YgfYrH0ynE9qa0Mi2ZXocZ8yxh28zwI6FjOiixeWaPQP1UEQhat9PfjHYjbNfo
ndPeOFh8NUY4DecngQybNRbbqHaD47aqoiR+eQwfvWY5g7A7BWmF0tr6IZbG5mOo
5IB40wd/WXIJNRANRZMgOvwB4ejxZjCn9MXc/JwKJTHhtypIogmo7m/OagZbfA5q
UHEjHGfSqvUrQh8QM8q32ZgV6wFhsilTOIlNMcr2QC46TuA0ArqlaLezTBfdZTZn
YJTWLM8GWgSARXEW9cOd+B4p92l+cVBRv+5D3DWks9yC0EIhINpl0Ik0LZkUzWOe
/DXq2Zg1iwyim+EFNRBL8+8LLYgrWj+zoB7vbRTPW7EEVLgAef/DLrpDTqMtoThf
X4HSx5V2BbaDkcxmDkDZkY/z6kIR3RHdEJKeGNAkkwe4w98puxEiD2LjOsGLNteN
7lXnvZB7w27T3IceifsDDN1sM56PA+Cop2JsjsRmxmOTzq9hc3VMboSym4wd/a5U
`protect END_PROTECTED
