`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wTZlF3da9uwhLtxnECGJBrXGh9VcjGWV/x1J+n3TLj6OOOnTmJzQcdzYp+9unS7Q
dby9X5AqocgzTx3a6QuRWMYzd9D7GXDj6BW7NR/IPw/FXMtIZYlWwEZIGs82SemW
DIKPNUD7h/QgIxxv3VFVukFY2GpOBokqIIempq+t1jXtxoivFb6tTxe/qUo3d6fC
dilY5l7Y5cdMwobV6AdEf8UoZbutRn3l3T5hiOwkvR3DP9x6TaEzpuQk1RTVfQcc
2ptae4zBX9axcfSjXdXhK5igDAStNbY6wpT1qbKrsM+gf14FlwaqWndnx/IhurGW
C01LwRJSWwZiKMKwrjw+beVXamgqua/xFVMW6GYCLlbQeD7gdKTS9jDvq2xQP40a
37MxY6VisRzSrLJe8VEvzKjspj5l+Dxqu1if5gGbkEimjPS8NbJzOcljre4WsrL/
wzfxSrQr4qMR/EOK83y1SHsFM7enxVxvaetoLV3qv8tRgsgxknybTIZVH5gZI+tL
kCck0gNlF6MTybEvQxXugC942wqtPant3zITmIARdeFy1GfJGwE/XBxLt2pMpjzW
Qoa3kb77cwYOol2hLxfW9QodwEK6AtNOQiTptDaKDlIR6NGaOsbICrXL3w2OAB3c
G+gaV5X14zz7ayNlcYgHEX8FEWpzsE1ECsVVMhtb3LQ2wv4HVdAlTqzpBSkL08tF
sGkADT+YULpJso2ZUxq0zg==
`protect END_PROTECTED
