`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XpnQ8s2yQguik2AJj6P+4Yo396YpDLHtAZhTu0Cki2okTwi3bv0meYXHvY8299kp
bZlD50ex84UOJP//nn8+srEsFOyhfnp85kP3D3N+tQbHp7fbMAGC4piGwJdpGe/y
4C57+g3fxpLAi3udjrSAdhirh5UAChG7r037LopHdeDmz70A30qzSNjKJdybF3Rz
HKoKoS1x3Pf5liEt7Tko1A1ZqmsbamerrEhU88X9UfHu6gXAFhzSMvSHZrQhLy7i
XGrb9UmLrE50dQRdRP5/rdoR+XdGXa4nlffy4sl0Fj/kFP5mtbLMc4nUiJ120Imy
bZf4x4T3fFxrfwi5bqMnHGiOFgq9sTDyOKg2Q0nznvRQDZObKrBC7MKg1DfWqMtU
vXzLa++5tbDCA3erF+m6Ua18RjoZESZa76q61qHYZ5bl0BW6NXpv958ozt3/KuVV
Pg6MNE1ptVjCrSJ7gsJmXtZhloNIrwAGkqy7B3g3ict1zQqkcwKsaekPWV4KHQDK
VkebXGdtnbMrtIhkSSeDJ/DosFvDiNVGoCdAef+qu4Xrp1VEZPd5uZmNMLaHe2Ai
sudQIxr2JlRcymNyMCPXJfb8txPysHoufT7V6xg5UQmtf75NvOMb32yW+DQ2NLyp
IXrf1/B6xO7Vqq/SHRaWq0is98BEOj25YdTfUxLHsvQcIH7KWfJDny82tjuoQLGM
rW3e97+Aam+h7PJ3TAPOaEhuG6gQw/gY06hvW5YzHgEyKMYa7hb3DQZ95pWxDvbi
AUjXL0LhLKIKBvG+rz8hkzpkniro7eaNfJGpAs9Bmu72O/3zg1ozOI7WVqqoFj42
4Y/PTd6hl9hRm57wwU3fEnXXEVCVV8aI5XZsQZXu0+7+gHES9DLsF8HtmfayuZR/
hLA7c2fW0ttluIcAwxZ3QLle1CqklemaV84ye0rJ9PjfwRhfynqL5RD4ZbA+4I5S
jH4zWrOmJbh2geiEAtUHYm/3gow32Wg/63P2AV+RRSS3jdqEhJYk+s97NuJQIxdC
hTQ0pq0FyKajVJnq0A0wnXoqdY0x/ioVVIxcXA0YmbIslls6ONi7F5lpJQbduZDA
VN7cF7EtA58k3i2b+/RnDWz6h0C11BeW8UgRQUwcW23nOH5psY7/aTQ+3LV9phrn
EvYBvpyghLzhZBKuL+5RgaBbJNTMO4Cm5MgobjZtnMMaO2Ddvt3GwOyTJm83wCzN
j9csebJaHNBGrnHHIZgPIwSnq23d+M9MVNZpaeRmHXvjP5p0KjsSiOHSTmoAyqzm
7wKPInhM2//SxwnywopbDpgSHajJoSvCjTXVh9tijGhUBIXOW/1dJUxTkXnxi2nO
RBvC+JyNMC4APxc/EegVDXSlHO5mcRqtVaL/pO7xq8QtVJU4ZG/MTHZ7Cu9GgLJZ
HKq3Xf0NDQ3ZiloXM95HBeTAGW7c8ApGDS4NmsaaNtmADYSdiUPmPnIQV1AK7lup
IaiOu5vlhglzUTJzBaOeQjom1Px4YoTLeKhovx8/GimY6TovgvtsKfcBeI3mnjp6
r21ehb3pIB01xaRpqmXfkyye7k+JMa5iFXPWtgoflcg9fOm903TwAm1ONd+jVZOG
qh0VL44wxYE6LwjEhtGy6VpnOr2P1rpZGqH0NGpM5sd9eBOptVnV4rAb7guUy0Dw
K+t/E58eT65wzmz3zZ5bwP0Uq+4oi3J0+WXvEHO/2LouQBB8LXPYQ73C7RgXGZ84
aoKUGvzadhqhy4TGAVELzFrQ5zs/FOucNcY68p/WKjDZg+yDVb1PwWkWIrJr8qo5
xte9mtQ4bI9nXFbbFJ7ru9FrpvvU9pPMH2GPgAMDU2S+FMjaHrKieBgRqRm+5vZI
nyAuu9LnajCOiT7oyZ01nh6pWtGeNGIQ6dCgPdP0I/0IYm7gKHKRHesJ4oNndLoX
ArsnJaZv3V3dGTneYEjtsPfSTqS18blGbCibP9JkwAzEE9E9xUSvlYzbXYcd6gb2
e/KLQqOrHULP5iCNepmblQ==
`protect END_PROTECTED
