`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4yTbNFD1fUTKfGU5HoYzc95o422Tp7hCmwSxNkjmtUNV5ldIlJCSnJ0vgO+6zdtp
2tQKIl8NbhZoS4NSuEdE23ChrPLvsBvzIhPpvhmybJJaMisl3Ozsy4m2ygQzDRPV
mqp2TOZeZkA7JQ7qMUoJsHRNF0WnasAvs3iooH5begyT3n3MCCawuoUDu7+ZDZpv
ikkwNStdaa1EKaNPG+NIgE3EkexfHKGoi1BmNDWGdQruSdIKB6gTQFLCGv2ZTW4D
ZGvBapzJnWl96CO4VPOxkPJPeUf7JUTlmvPpRr6bcYQIxm4ydmd4ZUxO7jcX+c8S
pNxW93L6fTUGB68jDHN0vA==
`protect END_PROTECTED
