`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VKjzOGwIqx4Q32sEeM2Zo4VfAPHQrcSxTCR0hqXGJk8ZxHpyXDwskK0dOIb4ZSZb
hLzsePRRyDu0Keb0q7Je4z8cwSsCcMRPiI2WyP8CXB/8IeJfkBt0uGdI3iIT//7l
42joNoYWNOErm/WpUSEidoXztVxnZwX3+Dw9C+2GksBKWmkZs+TLSjYXwb+i+E6o
yMDrK/G4GcrXUSJoDDHp+qlLce+gUKSfZnQmEKV4j6yLiusGTW+f1c+Wia+2/HDo
htyraLqUAOLgs8raF3NGlOQoNz9ph8Vsem9/qQNsEqA3mmthDCODYCn09lQUQaKC
NO4NeJ3Oujh6f6Z5VNFa3Q==
`protect END_PROTECTED
