`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7wnFL+NZvp37Km2pc02cUIlNaLhWuJ+nCNUd9cwFeF22bjj63kSCIsLvBlEy7bbZ
bmd7wCu1ZQx1C9XE9UddsSkT0iTtpJcxwzpZQmD9o55+LxOtFpYLK71Wuiq61t6k
A6wVGDCmud0tzW9rc1ZhbnnKdypdxm8AesPqEl/vhiUKzNqCUewdI+kejJ9fMZNu
Mby9B6irE7Fg8bAsCavGyQQ9CovikQxbmW0VuPlfzMjoAtWcPov/yB53vu04fWRI
IQeu9Ef5Gumy5vpema6Lu5EbnwaTColTcw0dWoru8USh8M06COF9VwHdq9cv1vJP
ycYGgY9n+1OEtLKS8IwJIrFc+syAV4lVYy0HkMi0rNhIoEePK1X6TIcM5B8ULqIU
3uF6Ez0AnhsXHIno4uC58qDXDxWiEQZ4ugTuLkRACyy5+i4que42GQA/SjCdiM/g
`protect END_PROTECTED
