`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8126JE29ruuVvgrUTaXsQR4iTog2OYLCUrDPHd5QykeivZ3Ay46DaAhl7jmLAHtv
RVcVISwwaAM5h12vG2d/p5XzQNkhUjZZKA3gSaZYouT8RUqAcRB55U553j6NfBpS
kTHu2ShXATd2EeAh2qnyXG7yt0dL+Aoo7P0QZWJKsN0MWSzYUKKaovhepxE6t3nG
YYF9cPAOT4Gsy7PXP/oVyc7lNIIxbySdIzXDtVn675vKs+iknJDCDPDjqG+S5Xco
FF4drtxzBmizzAcxSGaLtDKW0yd5klVLqzQCqMVNoDkVkhIBmPX68SbCbYbUI/9J
QuoxYgPktCDWvtnFt7fRhHA7CHIGAI5VErM8Hzfp+hlpiIaXCyVKVfXoCDcoCbyq
4A5tdZbzegp9czZ+JjunAUkWCsVQhu3sMPHuoYlUvUwyDELAd+xSbK8ljY/VWgQp
IprXACkdRxny8Q+h7ayS79B1T4JYMoapG9JcQhQ2JgLt8vggDhBsntmeQ/yLldQm
/xavCOPo7FtOOMXALqrJw6PPfVTU/bpEUQPV6f8IeDFoLeOXQoRUF/XsdTTxan3K
6/4joJ0hQXsTEHNcAA8NmWTGNHIg9ZvNl9zrX9fISlU47SMAVmBOgNxQ3vNXNKgN
pU9IGD3+VXwNqMBOz1N9vUWDvvnNQ1pQhz97F4NmL6xZaqHFLmda8mKJ8TbYJBcv
IspPruCu7lhpcBnHyp0VDMAoZirC0Hki3B1FNL56d1IgkZnBRREJ7DrWnJDCrGnn
jEd9POtVO6y2szbTyLJ6zM92dk8yWDLbfgI6M5MeO0oDpRWhqKxnMsCKUXCrjR9P
qBbq48x7AnaBvbuSIGvzRqYiQlEqw6nQs1qOjICHN50ydallzw9NhOubtmv4Z6P2
4TCw1qyOqb05UNRMo+j5uwxb2BlmvO5tEpSab/zM0n7VfLH2l7+Ksu5EThRAEa2b
4ehMBO07tNsFbhbPvaHVvOrBezypYErA2gKNRYbEKLJIIwqQFLMoV4ztXYkO7eNS
gipLoJt6aGF7PZcA5ne+6sw09OIOvAJSy92l61K1caS81AMG8XsJ0Ow03UXeDzw+
LovXl+Hx/UPujOU1N0FDy1KrSM4hSxI7RQA08z19mjze/CAfxlU/fm5QNyhYsZqL
JOr5S8znM/8G3rGgzGsrnzfZMyZiWORePnhgSIqfBersh/UkAEjrbTyvI3TsLbY8
GsnVC4rALj4DvWjRqJLBBHec1h0ok6RH284INKXc98Bb3ucdrZ7EQKoUbBBFhTmk
kwxS270hbzNZ4be8sIeZJe5L87m2UdZIIXZ9+vymIl3w12e6w4QT9/wiFlmtfbsI
ebmrX44qk5d3EgpvzMRQ6gIKaKVVB4MAG7VYfDsJEfyDIez+GVK4/D+wRPU5A+PV
Tk8npeVhV6gvxW6HVwnb3vTmAbVgv2TIPTYdCHH0Szlr90mpxqtOC18r6bUbgbrf
FFWYOvfI0ZYJlpAvNT9AY2Ck/C1rbokJ7/h+lUv2IEFk5oypJUBf3kEt2A4O4KiF
XJpc5GDYo3g2+NW+C+edElV1ztEcV6BjIWRNv3myOXWOGGwX+PbrbPQo47MUZukl
jCinqyB6hFX0kdZvCf4Pj+tszfUzN4Kor8bCv5TxldyhnOkO2E/yqp/ZXRU2lhMF
j0waay4yOCQtEWn1TGabzdo88fNcMP+WO5wf67cNF0cBmc4tjOkQmgdE2P97bZvz
id0R/tvUeiHv8wYr8w+TLjY3A8lGQP1SwVlAfndbKUkK2/w6bNQ+XJfqBzJqFW4c
z0n2mmMemY7o+cEqi7Rd48SPfJwC+UJ8v0CQQk3Ait/+0+sktkAEYgVAlbXdFTdV
iQ+HjhBWT4OeJwHRFunKCkw6hmFOyqlVZkIMm/Fy2tSzcK+hP8yGQIgBhN3yzR8j
rsZVpy+UrF2zq+Ov/EVE4mac0KknIhO3AKFLK5KPDDd8CyXOZDsXCq19h3JSUCJc
qzmio0hXZ338gasdZ3NZlm/NnaaLGHDzGknE8XYK9g20Uzu3lQmbg0PwFJufRnM+
n0mxyrDBSc7vtcsY8EdKVxTV3qCp1akjIGSG2xoYA3FmpSYVijgO1ddza49CinVL
xxNycRaxD29EvD3pHH0GfBW1INkxFp1NdP+9wznGkgpqiIBuQQ+UkFz/SVAvKhl0
cEgjQaV574tJymBY+4aNnDZqvi9XI91AnzQHD6MJK66X/xLsGB4kCZlA+gGaUmQl
OyrGGAFvcIpkDccnIMPa+stXnciZ8pa9o64QqYCYvdDJ/v47xh2hg2we/NF6vC3b
gsqNFPSWGQ8KYfmaD6mAvzJ2pjpuXd6M4LKmF3KrnaoS1fh1vQt4hFYI2A1LI2KV
UH8LMAJlQRlXl6YpxoZehRLaLU/Jj02VggJ2HrUKoy3gFoX2AHfFnDe1dx4yoNiy
PqO/2tHvg9zyxM9Q6fWFtuKz7NvfrQA3hVsEaXgh12o9/eeDgfXtUHIn8J84OAHV
Uk3pRTKzFOK4TjO8W+4cUVu6Hr0yj3CpbKGgvE6k8l/Rnjmhkn8eZmLgrXC3s+MX
aAFAt0xZD8FUSXyDroCAxeQ5FzTekfAe+fYP97pTLx074ZTe2G6nEG0DbQ4J0l0M
oPFCpmlaxl9gMmwj5kSkLdFW7K9t8RQ1JDMWUvYu7epS12yb8JnBwPNQzQFQpd23
RoU/xOU3/xInchnI4TNnbCRhyOWLqV89jOPfJLQdegrusdCU/ftXMoYvvN1n1Qmh
6ce+qseXUALSP7mIcgfi9tjzkh9dPvESWXq+TT9PQwzcvHInUuX6rWRjaX+/edHm
j0OCmtVrlL821w4AZfn/yllYHxiu2bHf5haBv9OYSAw2V80ObbrevKvE6p55pf8L
3Kb13DxSBBnPb6Utdf/BFllZAhFQ02V+Lh7YWan1IAgugbxZ9cy+jrWsC9SDMXNK
FGJySa1MAHcdmoLBkpP5tjOB+d9FSqXxNKSVeQ/R00hReqvYLisKT3+taNbD9Ndc
CW+R2Gu7q/HR1/Y4i4lTeMNODDo/wbt1VPptL2HFblr7DNBTlqz7JzlhfiItHsW7
WQQ8kj2oydVYcA0cjPY6w5TOLPFN17fzooR919FpDU61cF4W5PLZct5djGXvL/gk
VKea3eNahDF0yZ5+L4rWHCzVD/3HPCPsE+9kwm/f/+bALt7XXyvb7AmW2SmXrvEL
J02qTTPf8pgQFKVk8xy/taF2/F/bQvtL5ppT6p5KfnUazB+2XHLHRtGJHYc/xnhO
vcYXR3kS+winJKlR8H90OWPfYi7w2j3aWwdWPabhO9SrXYAQZzEx+1WO8woxbShq
X11vEjzpkP5A6Sw/knO9DNwNoPMda7KPfoauDO78KlJCwTBMErZbC1m/9EOY1iA1
gJ7FNysx92nLa6CZkTC97Bd/b3b8IRNyHothWIWyBtiWX4mRpyZhRFX95nKGlVCK
mBFjd0iJ0FZbX7mQ7mb+asFwSJOAX92n3bWIlR1xlZiV9PKncWV5yDaOJBpcvp3w
mIm9jldFPeAXKTrPpFPtqu1fLKfGT4fhadGi+88E5oV50bb8lG9u9ev/dwrBIaF/
IQLkIFXQvStUfaKA0dPvSDlqKE2Dg6w0SJI+bM9KS3bWyIPp056Vnz8vmdHb94/J
bWq9vsNwUdxCZN1kFtxJI4iOCNOx7mTVdNwYamrjhCwlRjQd9OAp6RTFaatIWXPH
jhDT3jYue0LHHQo1NXTWxTmwh4oFPLsqDgxEQLSMCJRsTZvhZqEl3tKnPN6rZiR9
DQVvsP42cDvtyy+bldrIsd/m9YufC0mzN06IuzZMpaLMAfmUr+VDAeDvpOFRTJvj
3XWBJc0l26RSsLmnk9QE9WYwGRnak/TNO5UOJPCBTYgvYnlWDO/ZKo5eY3IE0Rwi
teWs2oKvq1XdYsClkAor7WIj0OvhUq6MqcoX8nKgYcgVO1nFBJb4mQgEeGDrnTyr
ZgkvxqHGssVkpXMARBIFLaUfG3X5OlcZKjFdUQTfrtqwNJ6PcG281WvYx7V7mV+X
5Bi/POA0Azx95fpMSLL2MbkMjZ03DE2iS65gW2gRuEX4aIe5RU+6lhWnxJ7E4Tfg
7dhgJLSwe88oPfqCt2oZwGsCSbMeEI5ED98i27HfflP00141hQQdJInrsJt44Z8G
KyS18gzs4gKtYe6OPpJtTR/bl54jw0keKzHaQkUt7Et3T0ZZcT7r2ECeKlMD9aL0
1sB31szSnOztwmyB5VZl7GApCbo9YyhmQaU7UyrDEiBafWNc0GLp879YX5Y7zmCc
s/j7+UKhGekktpbmlKSSPPTfnyYTeis5DVZNT7uH3T4H4NxO0l8eymZpuv+KidA/
oHQLjgzXcEHLK97o58qautGYWzc70nTwDilYXj+eYuND+DuAFWJA5BU7SwPLEseo
kP6HMIxFqC8K6FTmb4sxLEsH2J12VBo82ESJOUP703OEoafrgFqX97a7ryJ/K/2S
Io/AS7owoRDjhN0WrGThb06TqrsCweh7ffvrPAFh+3BenBRxMr/cCenk6Tqr4tJu
a5Qj3mab99EF7kmKGwkPexRPxdIojdoaCjNRdHDWclZFizaNnwM9n77DeMmhSzk1
S5pkkEkXFu/fcnWgOq3l6fmTKs3DEmg0tQw1Ti4jdebpvcvbj48K9Ejc3eGWwVYb
+EN6onMYUQxYIQuo4x5GNXZ5w/cgJ9vwvZeNmEngaQBk0JRwBpId57NgVOyAhCC0
70izXvgG7Z1SbsmOr2Z811wVdKd3b+zQnY7Dv1Sm0KqIXQI5iOWGUb6UXLJmQzJq
SXn5qUwXb1QnVHz58GP1QvBQI5WMg7qs4Ua3IWm2IuZG+pBhsKT4tP4ipmpJDbXz
C7CS7HmwzeJKqQWxU1C8ya+vpvoPI4G9LlKLYe6bSvY7i2MtmDmraLQlmggfO8TZ
ZzTFWl1xHAlJt+DL4xRmRxi1qrJ5Tqs7dwXoZaRg/87OaLmjcEX6NbLAnjNIEnNf
wpU96CXWBfwDZERNPX9cDkdWqybCjEw7WOtBdL5qG0bazsz1aXGg/kVsMcXhb8q2
7y7Z5FD+DcX710vAh9NiMYe0ttlQV/DyfxfyEK5X4MNgBARH99mRhAnFXqWfVyPR
jtmU3S5dRyJaNjZPb5puPaaF2jmOsiAZ8khz5SI117MyZu/+6R/axctups4eJt3p
YQnabt1LpTP7ETVbuv5b1VLqwNXwmw3GnMQ5xzBAO60e6+03v1WEeAWP9dRFP2xS
X/k8Rgb+11YdVbBuLUBBEgPDXWlc+cviyGKWpPH7WJH0Jx3n3v4UWWdzgmPpnV9U
/oFDDGzYr52P9bXB2QIKkK7Msp0Y87IyNUJLpWNlATPP+BH/N8+qlv9xfKJDKvCO
dREszlHW8v1mVYJcA929xiSKt+cDBRZFUNRV1mL9cOkqvmssRTbYXv+aT9BD3tcs
rB5N3PRmZjvgz6gAQR0if7fbWoxNY/92AIi33zrxK8bCS77TexeSZ6rUoVgucKzg
m7WqWqoKFLaVE5pZqRLBs5CUeDbvyLbz0MUxbE8bFI03gqn3Ox9fxxWeJKSaJVRk
SLmVBaDkgmZOz0CMW+w/OYCioukYNuqJ/FD6BhSwEdvicqLvTjzhvBHkzFqQ0f8c
0iD0VIeLBTTwTArcAfCEy+GuDhkBtK9vpXHasS1QHus/iqO4SJ8z8ib5p4IvMq/d
6jgBpQYrBQFm1EbspOCqCBehAAjqJmyxTgnDQWDtvX3S0KMU6M0Fk1SyeBE/PCzq
IAZs99J/iv7Q2l0kcdfNQmGfJVokNfZX/Frf9TNQgX54UyA1S6dE07HR+YWC3zFX
5qyS4f45yKdCWoR38R70s74M9X+zcLdLm8ZYBRjtEh5IJ8goSZapFzn2YSL1SRst
6w6TuewjRDMVyFM0Fxi2zI3k3XtwDBuOE4xNAm+/Dv1pdwzkndhftDUx7SzmEQkd
1W/9xAoTmXtaxjEA3Lpysqc66V28aB4zLzkFxAvLvVQ/pr6bU7FWK4b8OpCH7g0r
SX+adVH719Cm6qJTUZ/xGK/bD3lichgc6x20OAzef4LO2ZygbUy3U5r5yH9HHR1P
TmApXXiJxa26SYYrBZwLpD7+1ynAWqWVLR5g+k3MG86dr+DHNwZNk4VS0Ch5tU3u
vpuDxEzj5EYbzUqhJuXj3xhHsl7ouHrIRoVWNAGhItW7+S7x+jY5JSt0oGnXz3Lp
u35bCPHL940m7y30zl5sGCBVA/V+fGeXyZGwpU/W3vMwk6hRkrgDka7Dqg8ZjOJB
4ywxXuLibhr+uHrO+m4HxDrs5Z/Nv4S+d7fyTPB4TrkZb2hhdWzX0vcsT5GQ5mHu
f8UTwVRThPEfbup7whOSnqYzVwCaU5nxZ9nPTFsAVzrwCw9PMcFWXEFH8LHNcZMe
lbk8V/1eGOpXzqIRXMmCSJ3L4tRQgM4A52jgMCYQIN8SoJl7QpRYjOUpGfg7NYiI
kxdGhhxKhGxB7e26XKGVzs58Jm/k+r2KXD1mHutOler4ntX7chCk83DlyAe3EyLp
P6JNWzjlPbgF2yr7AmLArR2lKHUBwmYkGvsGPU6myHubO03QYU6E6xaWRKgiQM/+
YlKslzXXp8GT3eBUn9uMqqmLBlydznEfjtK5TDcFF+pw7wL1Et+pwwinxdwQIOQE
2O40IEyO1oXWRp5+ycbXVe9xhmOfETW/wA79GPbYxp8JlnPKUTOegZKjnL034ku2
V385e0KwIaMOMflfLcu4kwR63DDA/lKbGR6QwNCk4rWHtcxNcfd85FGDvvE/Dttr
sj3dZh+RdDxXS7mUY4sVDlRD0rPRq7NEH7wPl98KvOmOs67kPAetet7FOl5QLhah
qWdaa3SCFtES5BHnbFyMlDXszwmQzwtL3TgV5xi9CK8rCtm0zqZeg9JZPyR34Ceq
/U3TaypUfKzK7svWCQ1znZyZXM+CLyw0quPvNG/oxEeszYc12pbYRgHSJZayO2is
d/iEtfXYWNhueZcRjiMD4BGUIvM1dpNWRWMWUlAxPwoNL6gIai2HaCvoXGmHTZE+
8idZSz7WLtE0w+XtS3+yVIbA8vdIMFrFIJb90qz6Xw+QJWMydd2WYSr8/bX+3cwA
DDaeuLdKG0C40O979aHB87ghjmHz8eEUMV1hJWvl8aqqXHcKoMM7o0mfllqZAsz4
qu+Zge6zYzu5mIG8Q1tZM9QBELbGWDhWnoqXB+bIDyb7T8XD74E2szzp6cdRXpTp
Rrxo9hot8zZO86HKWPxlvDbHvSs3YZ5cdBEVIMnu2XxbTGyNww0MF6jIxIZIz+6w
lIPgnV1iK0KoNZyIk6u9LrUUg3yFBdzwHA0gOw2s9+1y+mHFquvDtxv/rNN6VNcM
8F0vNv39ZuzY5u6xthJb1mq498Sdmm5eOGNjuazYhXHb1srH0NvU2B9HYi50gh+m
woRRkWIZZtz7AMgAIzbZXPoV3OEjMX1MLxk0CzBjk4s1RgzfQbYOxf/ugaj25QRz
KzeohegETMrU82X86jNew772+lBMTFzg3fbSJe/7kjB4OOrU5wam2HYqovvoF/zm
Bf9v2OYnEKyk1+ut1bxzPLgxsc848/uC0867s/48C3lQmeU/hsYm8Qz1XXavOV0V
uPi39vtWbwkYIGRqluUvc3nsnOymWYN9XtxRrNi5TcnREQIttl1I9S5cKg6YoQB5
oF+b9MNbJMGyeYbuULl5HsZEH7EoVgKrh1BlXsEzeR0hBNNTEiVxqOWCwWHEc/dp
gc/Bs5JHlTHzqEXlI0XZLTEsyEtExjD/t++mBqSyvwYPOKZM+/wnYufhmp/I81Xi
/0PFfTDzLTfNAy4U7mxXmvsUZvI8Hu3DoHmtL3DNv5/VC28VPr4JXgG6JdAmiSea
+miJikxePw4Mr/3ShBraTjIa/Oir9cxCGAcW0Qt4nzNjtChZ8QMvz6g6nvdMoXC8
ssbVtENYJ1inJ5I/uU0XN4smvsj4wAnK1UH795b+1S5XCziLCEHu2MwmpFl2wA0s
OjMTJIeReBUh/qbklSwkppBo8KSradOXiRC7rjyD4IhzGT76A73y4m1TipNkOZ1V
C+AuiBHmby6uxJBoCe6WCF7+nwuGzFgMMwshno063ScOcdVUBBnWiG06MuTXUGWB
Dd3DQtkiqOnqa3dHP53N2gwlfjDpHCz1zLtWAGnCp9rPENxwfZpjvrip/6mGkPMp
3BMsZIJz8WrxrVxE9QLp+wdR4LNagKSAW59oAGjngucs10iehPD0RgMBzyl8qKtj
SwxBh7sNohDwwVXPXwmb2M6iABnB4po+v6bF2Kbp/+JeK4V+MGfqfovN2ipJ8Lxe
7ZxbY15Xjc77lsxhChajtt4PnikegEOa1gGRUHmSEP295B65wcXeLC8UypsAo5To
pNStajbzRfL+0Z5dPn3tQpVTtqHrPSFSbmlhUeOnjBiOklO4JZdQtYotWZCRG001
6Ev5gmZZ5ZUzIez/nLVn/2UlOs7DqEi0sX7qFmW9+r+y09bX5FJPTTFyAS4O6j2D
OMnkBAn74q0HrX736IkigUN0MEfJtIVuJY0V8DKUKmk86Q49b2YmiL8XYjLFTo8U
d1RzZe4uKsVCWt5jRLpqcYyzN3QXMy3iJmokZoGyhoRF+CwueyxhVR1KmR4a1hR6
RVS/2k1lFFFxDbTmVX/DucooyGA3BytmIV7wnbzXae8eMYr/UbyWug9iaNkepW78
NPUiwmzrQDhZ9L+FGEHi5RTXDr9ZHHCLarQ8Ba/Z5TwKBNPePXsn07jOk/9nOKA0
mUln+AHYepys9sf87VvoTzdB/KreVD6bXd2KNlay7G9Q1cexXX8a/wgypkbBs9rf
CSr5zXMhKOiFIKNMghBitXD+kPbkj3BPVr37EMYEW5jm8K6cwfERdgYM+zTTBAZp
YpkVtGJQTXHC2Gfl4XcNHCd57zjJ6q8JUJk+6BmIB7UjJ0TgXMoaNvHMnNWp3FAD
ArujAyu0tFOs9ZRC7dlFHXUDMEGC5A9KIltLHc+fooRFf06kmx6uVZr3GE9zTb51
qhB7mOg3HmbU69EyaLtRADAgK01yKvXIm7UPrS+IH+AnGkH8VY3zJ/Mn/teotuYn
QSPOkKfB7ERcC83s3+/Me+9knuBGBGEH0wYmUEsIUM4J1BgWBmPbrxhCTgI5kA6v
tj7Fh2wlzgm8Q5krdMpC/0O4dAPwX4OXJIG7Zr05VlbhMcMaTsOyjfV1RUlcEeSr
D3AfCY9YE1E7Nd0xNyv6SyAuF0VtU1iyil2XNtIOFNIx3hPHFLFAVOGgD7xzfkw4
c8UjDOL0NGxP9Y2GBPJdgOd6+TK7Gzv62MymtNa4EH0mC1sXfSG2QuiTGfG6wWgt
rAuByHzlzxWiDBE5EDn68pxjFZfWOISq6Ert+mTXtD0Q2t6wjCH+t+if1w/ucP/i
SjSqhu2rgA0ZUXiYsi1TVVj3Kfv+P0HfelM5adMh2CXGA0qZ15T1SRZSqW834va1
XTAq0ACEhjXfMv91A1/DNRlNqU4lCg2ku0tOtowSpqNZOO4QBqg9Rs8c/3x2cCVM
sI4uCGHdXLWOwlpyUuDKYI5lkiSodeBbncIW8l7rylo+YWsnDFm/m9UlZ2bxMXpF
GEhATKICPLke1FMbsEH8goRZDF2KMreA0JTM/Vd5fy7aUROip8k0OL2u8PZFpGTC
sY0p+rLw2a5PCpg+CuBoq0qlEzrCSE2odm9ASk2IzMQEUc/K6llM6H4gyItraTDn
YliWoz8wR3V7jnU/68UvNlOZgbYCJ6LWtAIqQ5cdsntX8JUBdi261PqlwfG72e9+
bXBt+zArJ7OVjM+uwYdF62DKeP52pew3DcnuJwRYCEc+q0chhNnduSvWaKi26Yoy
79xJ2m/3EpWR7d7ayVtPwgFqy1ORbtNT1OdN1RIFrQNj8d+lbYXyxmlptLm3vBIt
INN+H2aOQqLberKdrSXJRPYI17B4+kluibLj+VrDVoeYRRwSnWhj3qJ1m21grA2v
Rsx+yCr1MgES676wKYjOKZZFqiFk/YhObeuvAH/DvcCxV+lS2At1BZhksDUrpRDY
hx8VXUqBkGreiaITBaA9gfzasRBt2rHRynCsuN5H9z9LpuGyXj/xsF6fHWC7LYJa
6YXrIFmZcqt99IsjcvfqSRHtbTb8h/CyeI+MvKWxT8NW3lkoHoiqoSSknZknZdUn
87jlKcY1LonxI+Zh74+H07jVk2Iqpr9WLzSJ6D70Cx1c3YNhygVGjbRdV9BuXLh/
4MwmbVguUp9+9ZA4MvvSljZ6LgaMbT5Ul3xa/UZGK9lHqH8i1ZTJwtboCQzNiF+2
XJjK4r1Xlz6RIUH9EsA4zqjfIcejZLO+nYcbUkdvLZHkNeFWM+6M/jLuOemPIEy1
/qgUoQ7WEq9vJO02xdsIweqBtdBtgLj93VPd8RDwTeflWNY34iYPfBGxXtauEPa+
bBBvqM35G/FR4cC1d22dk34TXtTWirlvgRz7lr/zJLEjbOkq5JnKDRb/ifiFy6X9
kjQKlMEenF21EUcdUJyla+KeR6yaGXrLoTwF2Q/uAc8QP2YH7gRfYjg9WNfgUkhJ
IGkuyD1o5ymBRRLUvLVuNrsnYnSHEEJP78SLauzjFrpPE6L4LkPcIOk9tWMMi22i
auyw3+NP19Lh8hfkGFOSqHmIbNSCHU6qQvH+2jeLGXKpvQOKnBAb+9qdCeWpsyaW
PJWUQiBa4Lnl1sYis//mWmDitO/DuNtDZTJBiflhuTa1lwk/9sxbKPnpYeo14dJT
V1BmLaoAiUI+9o4BeCPgO/pC9vhvUMkaxjtAVGhGnlZubj0HrbFapw5HEF3mURsi
cZwtOTreM7Rcw0KQE1l+aV+A4Gcsq8LvVNIbAVgECieSLrDwak+bTzBGTHR/w804
UDs4uUyMkR4WBBXzM1gckIIyHqvMYidLKnxbMSU+6AwublhXfL/cyWdp6rALBLw7
MH+zb52Xcwau60zGv0Gr009fs9pvaiPyjeNdhL6NrhMt+Jbh8eNmQxHVxCV7i3CV
kPQ/lnC0w6kh0bzKAroi9FtNNdirIBLHZP7s58IEba7xPe0byeW4MJF5st3oVoc1
NwMCRC8lQmoMneRb4+6znoGbtgtUZHxySL+G4ubkv+KlwE2B+pRKX6XuXaYWKIVR
IreWagqqcXnUMBbM9PQ85+NpV3u4t69GpxS+aG5WRZwCNl3oXfgAUAXLXRlooEZ4
Ujf8j092zLOque0xEszRTp5UV7NOLDYcgkOnISnedL5Qj5JRObeiD5k8MLNOCneI
VAffDQJRJu4bK9fcYzOglVWv7XGzGhBQ6oKwAsopOU0g8mGaWI7HQ/GP6fF9yQUJ
E+qvWJLI/7DJ6443IyzfcJVYlA6Zld5XYfHW3/0HcXsAGiIOesoWc5OBOPbeuMk3
P/rM900baELhYa4FU1VkIjStOKq284Vzy6bNHNkV09a7UgPEWbL1KwsOYQd2wFlr
Ao9p80agmTPG4zh9Xek6+92t8n8mp0XpkB7cVAuT/d1e3ahh9s73OZngApTdcasd
DgkLT7il0oKuXH2aPPnSmAsMOA/CiMHAeYILXlTeKqo+x89Hk2oru/FwqBeMeeTL
kix8+YUXXMhg4MCrscbiOdLV0rKSq6ovp1gkyqv8UPqgfVopiMDaCK3uyHust46t
YyZ5ldLxDo6j/Fr0OcBvNLSKdC1s3JdXzkWY+xl1meibmD/9hL0hWa4MhMNqPwP5
ZVGQU05PKMtd1SHJxFeh+C9RnXQd7gLwfo15lAwJ0LDYM8/nqC50n51iBf0038FA
CZgede/UJWZgAMB9L2Cj28wYf+WHGpgKIc2978YMtZNEoZaTcF8yajJirLxx7IPs
2gPBAGv+vXh7ExyDvYfso1Ap9vH9siIGqFTsY7cnfX+GcMpmdSlXfSPnQKyNM0x1
zZodI0Ho6RX1lKmZJDZzY3ZNYhruVtQPj0qqwwWygl8KkbqbsJrZ/5vy+uB7aHOC
x4pOo2NM3mjHPZC3NTYIeREahM/aBw3aztvqumzXg/vOEkvdjSRAUT2j36S8m2Tm
I0JnANN0oA7OF+xeui0FO0LSp5dVnXDHwjkRaT1lILlMPercnJDAlxQlHgDXKuhd
jx2WpeB8gK169DnYnVbnnxQ6KS4wiP8tKTHbTyT8n0lffvC+CiQRkNXOpt+qW8Qn
hQnC5M8ubwUmdVBDZfscz0frn5KSMVZIVNjGpAbEu+D6BP6iNf70GUO+6PXmaEMp
9jH6NZR1SuihnzOvau7Ya9nACs7H+wO2e/X+eFhqVvM02LuHpK24lbok2OImR8ZV
nE1MGXoxiPMFF1Mk6DgOzSWPBo+sjDm7L81FrUTNGGQlL3cRqr7JbXv+ntgGsK65
WrcS0EdEL/tPOScBuqRxW3gGvOghZCxZUnWAOUIxJ8XkAuM6LMwGxUaG7V4pK2oo
AM6ZhKMFr2wrSv2JI5KoEZoLJI4G5IbH3ydaDj0Ctqk8Bu5lflX01goMgJ2qLMip
ncVcE2Ws8QSgD8GfkRNYhGS33IJEFucGysqL8pmq+Z8dmQgLnxko+t+EJvxAu4uV
CvAwoDC/kbzz6Gu+IwvC00b3tFcDM+pdlYiQlZ1zIYwsd6DCfHGyce9D/leUuAhh
ZJs7sSiJDQSIG8IXqAjpQjsWry//h1YhAkXqKBYw5F7+6fb17G8HBlWA0pzaHZfj
8wLWl9/oQjwqvSeRB3ZN8W9xsdhxRnyKvmbAAS/d4UglaEzo/BfB78pPoW7LY9yS
ddWVe9Kn3iIOahZa3ejQ9nbkzohZpqCzCtiiUDf7fiy2wLiMxnpi/B/yQua8dP0+
/FZ/BSrv7aNztnfRT/zctEoX5eWmXYw9fyWNs+kZQqApDWH70fMiORmy5PfkacHm
wyUMxcsyNJdr5eBJLRiJ2uHlKepeIrfVRlyEFLvG6FQkxqoiGgcMZgLnElHGAQ1I
M578Af2C9tlUkrap5tbHo8vlpnBJy3SwiR6IWb3rF2bNdpg0PjG+yAAXybTqlDvP
J2oLyi+PTAinxNgo3CmiOWudFbS/Dbo+LbgyIf+XX8j1FDm01fvFWhFBe9zDAK/u
bkK0Q46Y8HWoGpLaH5MgWvo3OmIvJ7zYuw5Oz25vNuHqp6Jd9bKX/QytoVXev0fl
fOzz65CFzmoCW4I5+MB27zusJ4F/XhcEdq3fhpLJTz2fpDSOWpspsn1xQ028yQpc
F2dqWgQ6ivVFMkpxCDL4AYNkdK+L9f+9TS4PjfysYLJaVVXY16E4+K/1ntWa3kfT
lP1bQ37bUMpVzR2Nd/xvIG30s2/IaPsxKNLxB258n/FCStd9x5ujlxuSkxPoKsYh
atwFc4w4hbJfmhFZLhAYpzHycb+xhdOqa2e9kaq8ACKp59MX1M7F1+iv33SXsslR
PZMK2GJaUBSF383ziNyTjEKKBSsjr3gzP386lvBF6oR/0f3ixLRWqrkz7pZ0wZuH
/eRoBoP/7IYvuMoX5sKKwdQl56F4B9PF4QfMc+eSN00ySSUprOYbUFLH4+rilUv+
pyHYvXGXT7Iqv7/7Ck0ZWKmN8W6wLnXtwUhrenngpmpDCiZqCrlX6IB6/8d/5J3M
6WHWVQ+gnxao8vFZWUHmfrrQWUkShxm3ItRTHDHQXQm9czhTFQfblLbpZZYRNl7d
jOanoNEN1kopsrxRg/+s7QVDDWyiGmkIg6uJEHsSQ+vq3EIJWuk5OTmP3ev1i4kS
EAcLVYDXCVFowPiLYbQUIJ+k7jX+Gpt0rSjjQfG/ZqYZHYI5GehljBgzE3Y6FYPX
3vZKAJqnFWA8OZK3P461wBks6TwNzHNdBH7b4AsRqVRwTRJ2wPrgr8lwHaOmAa20
LisWvDgts0hZqrWVmNxik/bC08ulkWxCU4xrPMqV98qAyWYEKAQXkokLT16jF4MX
zizEgk768QJ0M9NXrkJvAPaU4hv3mrbhwWYB0MGuRoS6CASH56/8MQ7DJ+Zc4T4g
oAbT7AItpwMilks81qeIKxws624Se6KtSFAw5lB4pM68NIVmJBLX8/BKphPO3COF
obznonW+beGGseggBv3+ERsdrdJS395Tc49ZLDJxPyiEVdXBB6QNWiKSIx3S3+l7
yujeOThyeyL6bWTwfsgDOD23kawKhn+NA4uSeXfvs7BiM0y2Vob31oezIF3MPyCi
TwSbO5fd6Su8kp3PtblctGWYmcw6nT6hiBA9oP2jGnXa4BLJcnnlfv9v2oW6FUP2
Pgkg/N+Y9LOcZFHj3fKwPr//1VP174JmAl9z3LAJ6pDOuu3m5kUVZ7VuD17MZ9r2
+IRqG2lV2YlGesK9q8wzSw+Qpzc4KCRXHozOhsm0mwZYUxXZtWaBDFhwz1p+1tla
UpsWqQZg1GAMY9U8dP0fkT7rVR/O1efTkWOaJMjysZQ1Qo+vY02G2GOl5dW/vDQt
6LMnjB6SPS4MFmo5g7yOA5JgdlLPHrLiGDlRsNeK6bfAKuCC4fwehC1mvNks5vEL
NBMbLB2XGyObQEP85ZKTd78qKZMloSXDU79gHIrK+dR95vhOvFsfz/MZNyBtoIG1
s3MmNz/1GEXJUNJy1gMCCQvna4Ns5D9JVE6KjZvSInR3RMAWu0ppwfiBzJzN29za
xCLnLs1nZ6WqjpzX0IRTS2tp4KAG2ENysfK5xvOr4Gaollmxs4Gg/p4JBiEM3L/0
sy4mkPu8a4rB351JOLMbdLE2W3X7wJF82boj+ZFiR0rpGmsqIgqeZMTEGBWUASxF
muOBRzCap+bDra9H7kS4RWZadHnQZr3YAKAlt0cD6sIkg4y1h6W0c4bxaLH2VqQE
GLebfbLKQtx6KGeM5/ODFkPYRuiVpNMoHNlDbo/RI+fZHmW9hlVwJ2UAwoaGNAtX
wvOg8n11jjTyHKilV1LnTHnoA47iA3/2zGo4HsaaZx97YKQbSAE9/8Q149BCQoiO
cHeeRW65WDUPTef5F53+681jMXWR47KeyhfoLy49a9uMaL1AT+8qT0y82uZbUVnf
uEoPcU0rpphD1I70dyIvIqsnAWyxnZvxAQxCsR7uu09NQBwX/dzijSCE8lWA6Dh8
U2V1vBBYuUo0HqtmFSEpKN4CloaVp4m2llFUTefrHLJd2tHGc3mUQ6xY5023VNYt
Nj2vvsfFLykaEYxwsT6xM8O36I80RfMp4zFawdo5B1bjduwXA8K7ERjtRjB/zHrV
4E0WrguqiuSkdtrQl0BDSxI1ZrwJHQaEukJoUpX3N13qih3zo8/gPWit51JNFBMI
oOwDPgvVm06WVAhUnvYpK3bP39izTy+/n8dKIFxky04V447vgX6/jxVJr0hE9B0s
K8pprw36qtvrNmA75O9r3aLme0vElbLRqLGWlSJ5H4jQEmY9wz0Ax6oTspS54Wv1
`protect END_PROTECTED
