`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d3dBQYtk3fZCssISr658FA5RdZ31yLbKqphDOXjcIARFUV82u4qokB8J7HfzD+Nj
tRbgR8G1mJ/rmzy4z2W+hcFngTYVOJ6lA7UPTFeaocADO1i7gMMK6Z78Xdke9ZfQ
3enHetnNEDnZRKgb5WOx/922N8FLunsfO549bCCkVXW9nymQfwuQdLuRcYnqLNgk
I3ByJzyMdQDqz/MKRpZWCoqh2LX7dwW9UMJg7kLgfD1hOLEXrO/kU8NiM1g6kbtK
aUgfunjqIkFf4VQOfXHLcu7wjWXEb80tbgoqnxPMCP8=
`protect END_PROTECTED
