`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mKo1HxqQv3Vsr6ciZmdMs0URXRO+Z29n+zY80DuGK+uAbkyXk+xKeaBY53ILEoZv
OAG+99CCuyp596hj0FkFaamkAkPCw/T5ff2uozQlcnFDHFcKVlC5m3IugL4+9E7l
39VgKB4mX2RFN/7rJKcRoEYIjQwU1QxqyeE79/mQdr1L8vldk5XrDyzbvSmwU+gn
VMOAjVHVnUYnUPGDa44KTAu0zRWSiyfSxajAL5SvjJRcUS9atwaDf+M28adIS+Hs
jAJuAAtSEl02wBK+GX5MXBh7tPCLVaiVGmETGvAljlsi01UZ6djUkm36XMUBBpYH
QG6NPO/4uvxaRUoZavGiEyf28c+kIiVIdG1bzWnY5oYh59ecSTqlN0NQm/EuRnw5
5H7zcyDDJbCWA1qbZZuQjm3B2JzYOsVwswNSCNvji027FXmA+cMwbn2rSxU/20u+
W83C9zXTeoxGfNH5RM4cdiU5W73Te61eiCswEri8YSlFMMCOOj/4A354nnSvJRoQ
grZ/VRAxB4VpptoNuOIyKT14237joJM0ea6lQ5FfZXoB4rLM7vYG1V0cvhHAETi/
AbKgWrzC/t47/MQgtvR6EhvkE9LOGX7Fb4oGKWPiNuaRA40HRG/mO3O7dgro0Uxm
VizHpDukDl2Ejg76Yb7yS25IKfoI6oa7K794I4q3Us9MYHwlsVC/6exmnK4wnL3C
dtxUeGwWFP7MQeHP/iEUrVrBhis+qCNOTBZIZ6Lr+CwMsPV7QWEMbbjCO5x1p60I
5j4TpWTKiNR2razmjK19bSa8LIVSLi6SBQs9DXP7ZolqhPl4Gq9z9JiFDL3NC/tZ
ofQp8U/nd4nwSSWixdabGSVUU3rGVzPfFBD4cUkvzAfNhiNCTpZ80HrYnBYVkbyL
v4gQbGGg5NTyPLSdb/53enFJrgkA/azh4Ie+LexFpQUAFrlLkLC7HHbHeIsf2NIC
7E+oZpptjlnD/auFCtA/2YRn1bCo45qH/CntpDw42vh9uYpj3IrHQt4tPGz3HtjO
w0kpjaxmtxPxIKx0yeYNHlBQR286E8Ib6Mc4gC4VX6BEBTzmTJ5MNBC/+aefTl50
pxk+ed6UcILPFUssBK2nN+j+LWgqPob/eIcDN6QAGV9t/O9VvP7cIVteURxDhwB3
D+9h1eZFnE7N59JUe7k/XaGXHNrLxHDSP5Q6vYHx9sRx56dwyju8AjUOaYS7nIQj
kCm/KqH5VGQkowk74KrQOXw2NGxLn5VPPS/mROMoEhxCvpZs4Eqkj1uwFx/OqXms
C2+H1T8ZQznvSoxH4EbN2dMdMQzN2dmj/ufX6aIF5u7DZ2ngmI1O03376eElVCC8
xSuHH6AZAFZ2wiUxTvSKkVPhwOgtuGcH8+4180DvKuRVtNSLjEp3ghnSCNbqtZI0
ArEt/H5Ip4ybuKKZ9T2Xe1ZCbjHs3fa0YujZElPLBuX83T9mp9sCLNbgxhHEAsKa
q5BGnTUDMTCSuThjHEOXxN2w92+Hzyz+Sd5IyGcplCHpkt4LieWghMIgRr4KxIRn
sqgjsPOR10b3ohqJ1T2RgmO8qVrqYP0tOQnos0z7ZvDbxe1OToqGsJvq9D3ZZzQc
k9Itsfpv3kvBafoZnXdhNuibH9PNRw9VqeUILg0AS0KpImasSpmT4jFIDozOliHy
U6xkEaa1k/aO0iJSksjAkA==
`protect END_PROTECTED
