`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9ueDpSV4XuVB4cIGiAUWu3zzdzC02W93qj5+pdh3nyt1b2c4u1Ew1B7tJE0+dkWn
qwWzAc47+iQWDIuNCItdSN74Kzjdp8PT5i2/8nJ3z1cy9i5SUmdZHTPw3gI2xUBV
rbgs5fhEItK1BeiVTSLWIXOBGQgkstai4wyHXmqHGDVKlyhN6DJdGwQwljku2CNX
WxL1gf2aSMPN1cNBGV/7qnyHJ+e9Xfd0MvFkPN2cSkm7vscZV2FrB5wTXAPxQ2mo
`protect END_PROTECTED
