`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MoI8YM69XVJ7nREHl0/DdIzMk6r/xs/yIPVcAclhqsTJ2XO0UClnDgqEQwW7FW3j
6ps9uJe5QOhdqbamq1STssxcJVxNI+TaqWIAF5pvWZ6IR44BElyYrwvzIOFtKVm/
bcv9ECUGwpf/5ZUCUd2ZQ7NuM0vCBtXaoOFVdubpOoBPnHOVxShODElTLQZhYW6B
UMSaAStyKpBhIg6+TaoLCdM3QzNyqx/spsZ/6gTadbRkDJ7SrHpgHE62aAIU/RxJ
32bjcK813kjYAHcQNOeU7MJaXuW02TVyYuNITJHcv2MovEfewsNamQoYPgFdbhAf
qJs0QkkYnSRBQBA+hhj9GKcE0cbw79n+cwTgDcMVH+Ya9JKgknYLeyp9T5EF+gjB
ioM6mC9PvbchUUn3djBslw5gDNctcVsFMiGW0hNhIQepSh5QpchUZjsZ60nVmLnR
XdW/hBwBezhF2VGr0vFYbsBrhPfgjrhXTvHvV/lprTvLSPE8ST63s9SQbfw6qCdV
p8CkwAxz8D8IiKZ509lBHZ4IaMibyTjHKJkyEsmgmzU2lbe0cK5OXAbuYg9LIqzp
FTpkt0tSYCCQbFAiHIL9Sj9Q68rqN14n/I4y9hN/m4PZBgRFNn/IavxveCP0TNo6
meKKqkS/fEXm+YbXh92sRcvav3SZ5+HzJ278sfGTTUmSvqZ0u9GUaZWNr7rCuyuU
hsrS8H0c/Xvl3z7K5g0oS7k5IRLAMIoiufQIHQnHy06Y7pYty2GQYLQM+3wC41aC
cGlCvr2R9WEm1j5KSblGDg==
`protect END_PROTECTED
