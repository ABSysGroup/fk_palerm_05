`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R4950+mMZXzl2zKkRzXVIGoAmN069HptJ0vI1Ogc4TbJ1duMMm3KWmZFGJ+2/Dbo
voewjqqO2/jb5MqVtSpZ98HbQKo18KW/PvzjJFQ/n3L/EZiGd58xY8/dN3Pp4JGU
6SNjdDR+GN+/SKMTucT7hDelL6v89+CtrpBTtoHc8xTXD4b3BmaF9y8vBqtu6MTm
ZyS7Y/o5DQmKoSxhvcCGKW6U5t+S0zoyonHJnl4vNN6cqUvNbXDU3ttF5gX6E3En
rqa4wpMEyly3huPP7sTXJ/IdzmON+R4V2q7o1fv7KMMutdTIPN+//s5n9Ol1rlnT
GjIcF89w600V7VvNteVSn/yrCBEdlEJJGE06B8zVHFmUCnwU6arf01+yUNLrwQSU
/PSbcAtaXWBJi2b3niNSuSHkiY9A6qBRSk7Fo7DFCcNCYV/hKL1C452tcASm8E/w
mGOOqJsL5qyguGpgKgROlFkWnwbZ/nuuhx0QckWz28f19KZT4dq6SoV5Pna58msV
s4pk1pUCtwFCR23deas/g2i1yKvIKRM8hUsvGW8s3ksDFa7latocuYOI+QZ7WSca
FQX0+3tLeMK3athEGMIXokpisBMDVEqwLLRO362CEgKwsCkAY3VoflsAngzBmvfT
DP8ZufftLYwkNZCH1+RlYgMbkPzdgqat4XGhqbJcqng=
`protect END_PROTECTED
