`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l7iUsoO6CFOjVcq5fyAxsV++pFRIfklTByXuv1KTfZglh0SKgsK6nrsweO7xQN5o
jKeCkgB+HQotderXzNp1Tys73gnpzer7ZA7WvPDUzx4jsd/clVZwbVZoA8n/yDxd
bjzqtmgQXtdFtamlqAWFncw+JfORJCEJDIzDlJ6m5x41xNql69N2VUsCetZQxMU3
/NQptSNQQj6hHKWKDEC/ih/ZP1GLWUcO68JRoaFTipGuM8PTpyvJ9ggvXgHt7oWj
Q4HZHJi+GkuqK7ucNrDITX00GNLewIOX0KnQ1Ls3K2mofma+t7E2GSlRDE+2hRaI
u6lSu4/wE3WvP1poXBEwhnX+FVU0WliTRV98rzhZTo+ahzc32ApdcLEyi6fC18u1
L0F/zMVaFEP+pGkxEli2nWsg1V1z98kuIuFUXyIE+GHJgWG1VnCmLyvhK2TyLTmJ
oCmaTQQo1kyDyuhcmOu1RrFW6x0Wff6NiPXJDrWqHpFaDefjEUvpZJL3UrSgvGq7
gFSYXHIpGoQOc52/ix4Fk9KDrDKUGWfpr8wzT0dhY4XfbC+8tEsvwnAiFIy2Gfs7
g1eMGYB0bsq4RlK+wzpxOUyKcb3t5RuRK79iDfJdx8q33F5/zGJ4zzk8iu6LHucV
XkgYpAZWGu0GdbU9QRC5VqOLzxM3jgH5HJLUJF4dVc174nhT3Nl34MmouxUuTwXX
7Ly64gKvvk+sbvosM6oOL6NbDjsdv7G3r5WUtUuizBmqB9M292lhtv33jEwGsoBa
/dxw2wNe1iZkJChnIpqzV9JOE+yBB7bUh9redmhfMTicJDAKl+5Rc8k2gPpb3XM8
JLXkL/emQq8xgZt+yrzX3aCjYfGSgTqKaLo7vSGK02rLtDSFBBjj923D4srF+HYN
63cu0d9Va0FI6unecNTl/vqgMDthBW21CSy8aW2ss5Hvh2FuuvGVDIeK+tD+m8PG
EqGsA/mZINmvQnNN2hSUBLxB5tT35pVMD5+I6/I8JH16gsaYiq8pThGf7pBZ9wwj
Ky41ON256uitiQKe9UqBr5xU/nA0F40fIrCY2JyEPzM=
`protect END_PROTECTED
