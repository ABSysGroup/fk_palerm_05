`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g1QJ2PDPRvu1nBTspEh/4+mQ4PJdFeObQKydpELQ+ZvEhoR47K1P3oamPE4bhqyk
xqtYeUTtHH2tzHqZELhweHrpEkE+LnDoYOlDh8BcR5sY8YhsMVI3WN3cAPawYcoK
/7/r725Pw/x9a2Rg4kcGpj9k2DLQS+EcTHtGQvmC3n8D6zx/kvnGBTsUOaJouWIK
0VOiODhGzSoMjsiD9rmFciKGV2ci1E/IjzBvdYWdabN3Mf1F87CY7Z4z73pFsgYB
bVzA//uydrl0k5JqdhNmXT4WS6oNaWYLajNncs/sMkOfWPIPYbq8egXW5f5dXft2
NF3pCj4AUGa3N74TTKXT5tYxHC8KW4Vlz/VlEb9yWxW0MJNYubHePHGGhbK27Ovf
umaNcx+yq7k2oKhtKZEgD8i5Wk17t39COImJ48hMoigr7+lB4okH8K7j/sBYP0qN
5iYs27iuqWnnmTyx71H/BfES49Hdk1CPUMIKEnXxhsskPGxDxkVwAVk3/2zaCDMN
MFdhr6osSG6aTCp4kn3PwOIOh6fVPho3PXJSetCRvdpV0d8Pb+F/ZSxjI2ejRDrB
vUQ036k+VNL0fQ1mjuhGEhPZwnfGSsePmtOPnrP71eEoAegWv6bvrurLr9ZOqEBb
ZfUH+ctz61tdGiO5I9QvdWd7kpJrO+ybEqGgwYCRUad7ytsoK0GrMtan9WLMaUvO
AUS7tZn5JJLg3UT/f9y7QptQFeZIs8kBmmA/iAHkiyvrQd4jeh4AfC2DnGrWzwYV
6ePKaCCz6RAD6Md0heKnDh/o/AH3bo9AEaP9qbnK1x+nj0j2B44h9vuK3ibJ9dDf
rq/i6evHPobJGIocTQmUSe5lPB8+tFgSXTjdW8h+fHR1UW+YY3BxxdPncbSr1myy
9XlWg7g+RL1aiQDcUaTxzw1oEbhMJKMxlGrcFD72wuRSIZ/duzL+3dijftRvz5lH
izSynmO4upl9xC2RqGlHheIPjxTATJDY+u+PisdPnGnr7k2NzgVxykVsMpRfbOJU
Lkfcg7g/D5Q+81qQFL2PIP+lOhzjUR/uqak7WDqC/RUYEKGQCxOwBUuTE6wXh4F7
Ms8thH+PTY1ztjRrD8zj7tkVfiCgiprI501cdP0LtU96753twe/XL8K26wBvfMqn
2JJ29pzN692vbG43pk6+p89wq2oR9oXyHJPmXtqy8sse0YgJwRk/ySMjPpNXpC4F
H90fde/3BYcfKo+o1/Wf+geZ5Rz03bEDSoG7fKwJyFpwDRZK+Chb5yvx8xMh9wc0
QZjZijmQ+Q+ITEz8the4Wa5S6UCCFbrus1N1qBcG2qrLn4Qt7+cN5Zd9/kRXKcmh
CKCjLQuQnES1UDw3DffYcyVYBX5YZGv1sciCWquK44y34iU7oPxs7d5mfVKJFQLZ
jO/+TlrcynyHD8TIoGtWUfHIwgIPyQbXFNlYnOXdQGE5jowh3pY2kfom3paxAoeS
tMCnQ9rNb6pQBqWiVGRgnjzMCkWegd0Yf/zm0iJakZSIPu3OHXhLxvW6CQM8ARqn
e/YJLfiwM4xg/MsWKPocOLUigQ0GQfIKGEJnvdDChyXAgq9oHXUSHT7Pz5hbH+Gh
UyWc41Kj7lVev4B5ey8MPqOTuhjy9e3w1VJ6rN6l1rdsS4RjjlgB4RoOMKN0gZMK
naKdv66OulQ7bg+8mCv2tGs2vmtsLcwx5bTPnEULqTY9/V88OV/UqtEXhZD/psop
RUvc2Lje1pwoCEwAXnbaRRRb9cbTij+A/trHCRFuVVdIbH+F1mBPLO3//5LBMUqv
97H1mwd+3CeQJXCsbjcCXvemQiUvgdnvX7QFQFi0/aoxe/8SSf2ZFUGeRXgAFM8T
LzXa8YWEQRIORLt/P+pTjcwBXf1aAJXv8yPNOT/ozjsCgfqfyLgxEW2u+G+g6JCf
FFzsd3cWwE6y5jp1IgfaWx0Psnp+wf+KCyf+COnr1Zzq5L8ItCCpFKsLT7VKQQWD
oXmCuWPiCnD6EDjA8TXtNGCP6a0Fwhdt+ad9KOsTdLr4cd7AWHLvKOt9wq7cai+h
onE13S3AOoApYzysKVxiEs+fwaisSyqGlSDu6hTStC+Ld4684K1+MQTXjFC4wr/M
TigdOegnoeyLrRseCuJhe4y/W4PuExMEnEDOovqhU+QajJj+rRGDrBoS7a/NUnZi
k7R8Ai70Q/QFX+s0xyuyzKschkKq/QUC981Tm3EQsKMOc3iNJl8b8itGadXPQN0z
APA+nVGlU36m4UVnsWgMljLi19+zTeDBSILczQYuBOHXhFwoWjoEydTPkcdjOywJ
fNuTvr2xU15DLwyj9fz0Yi86KfBSdFIR0TwbDW3mC7/43pQdEHGQf3pLwFH9AOXm
6T/z8dZ04aaeMeFOc+TRo7GlZOMqygz+B6Thp/b3/Tox7mYN2DlVzjKdLsL9MLyf
hq5yLZ3igwfLAEGxNP1SUoei2tBps53hRvBXZ1rHCGxa+bVvpahkmaAaxww9U5rC
KwOfAJZjdZnB+O8+XF2G+7Fbm4jTOUMyB1z0I0ZHGrOCb3akhjDNt93+pDqoHzd1
2ao31uzpKfd22q99bSsNXcFehWU7lRN0ewsmaEvk3V9G1BsiHswaZbhKEjgPg2bL
6qX1Bc01z+atDH38woilaZorMSfZlJsug0SlptTYS+WD2D1S4ncUteg/c6IaJh4E
PWLFbi8aS0J/GGmsMXm7hhrhttI4O2Kj5+QcLoYx/8pbfQOHECYFnPkk5VuEnl2S
+JJbGri9qPK9G33G2oIUnNkO+9mlnMOANlvJjP4A7W4SBzKGPqmRy+Qgmi/eQ5P2
15a/r2NFauT5gtNPluDxPMVfQlKwVEoTxJbmQekNhgfI8ZBPxpzkySewFFTv/KLq
vXW+ah46rrIVaDKCvVZklLdjyVURcCJa6oo0K0fXgYyySN5SNe2JZe7U4+oqT8lB
847FE3kpqXkHsJsz+yL8uJHqdvo40s4kC11FhsUQJmspSH5uFIE/kMcEgxFy35DZ
6JRkvv7GF4hhDmMzrcY07zcOvZ9gZf/1plArBPHOjqNBVVKbc2VlrlnQfnAktsI9
NtDMHUwsXBlT9GS6S5EKXg2ZmaYyOaErtI54Ny3GxXIgBKFmMJh+s8jpoqnZniuG
fSpBYrBQDzljGEJVyg5y/wPVUtXXtb3IY67g4rLQ9NCBB0WXNt/MrR4iEIh97pe1
AE0ED1AZmm17TVBPjhG06wQV5uE3sIZiUjlj1dJiWrcg4HdHwDRqB1asHlH+eUj4
2M0Aoe2Bo5A6tuiHPtIQFPoPelt8pcxDkqL9c6INnvHaPlQQ5IjXMaO3gBiwgSHa
lQeA0A0Au78gyCn2avShqNyOiKE4BI+JM3k54Bx9P653N+NsHe5qPpD2BK2ZhMrG
qzYgt9rliM95xg3HLAb5zGLMI0ArZWO8HIrqSXmx34oblbgitGVebAIAMm/soc0f
C/MeTaT4nEFreJSzpLQ6aWbF/nmYhh/BX2W2YszTx6JNlIlYfTJzZTr7H6WBjodP
BAfxRwPihFu5N/MhAdI24UmoHZvtJ2qI8T47iY5dPnjG10+Ya6LZlALuGJcP6Her
A8cwTtmGgbh3enOxGIWktoOTX9CDpsc+Vaj+/r2BIywNSnSwm6TcoH6pxlaOKbME
IS2qyKdxviaGy7lT8o1qL/W68EIDBh7vdhXub6A+ojJfVi2WlOnXiMa6ec8nYm7d
Obpm5zGG280Yv1Rr7Cqj2irOdEoNx/1lbP+Yce+Q+Ni1lJqRhW//vXv/1fYvz8Co
Oop3fOehzzyHmuxUzsMt4XGWrk+u3LCPa/kK1CKlRaWfk7lL6QWOu0kZosPpYlzG
YIgaDy5F35BwsxGLY4ChWR0eOPjN2SDS1r07p2KSwQ7ZBwcXXViSxfH34vh6eOCb
NCnXEtyROnJmNnv4Yp4UiNqKiXwbJqggERopdPJX21loO9gHb0W7p4alSJnpWQBe
oBVIPDJqUeEm1elplYtI6sFWXKhiEkg6KLj59gri2ZZ6iPkxgqI/dxkZ8uSu9c7z
g9MV69Ggbm+qUoZYnDrVfKP1qeICCI1ic3O+JOSZYJV/VEtaD5HCv5gdOmJD5QKs
piDxXR586meBbySAzMZb4GWMFqDv3OVQrnoHOKqxrm+22knSyQyY6xfg45LF+KPH
QWLUEo3p4AhyV4RCjkoxpSjaFhTwiloy3onPI/QHRvjbc1HTXcY/FTuaAWx345yy
In4dGeLcmylhDBaiSbpimtV6xkj59xI2/Ngtiyn2gZmZc3ntRR2XR7BRdoqZ8vva
xidMZfrV0OoqlbYybY9WuyAJgYFHjRLxSUe7PekEirT9BP2uQD7zsTKrIXup/CRd
9ZGwwq5mTr5bHAwGoH9byBSXFmwE5cxU3f29CEsh1sjhwpiMgMbldvDDVwafnQI3
xR+raob39gdcG/lxd1Klev0bx5N4kLb7/Q1jsAKOGxWQUDxH1JQqddLV7X71VcgW
f+v0axAY34/P4Fgx40CR1VM2pkf8lwgm7af3yi5ZiCwLXV5vAJENu1MjDbNl0gst
dsup6fVgW4lWgSRcHnKBVtnrw4oQruFid3zBI85UojpUbf6Q7vkKqF7uAulQk5X+
Pk2zjHRMUgpa1HD2DH07h56A9nZ6hr7MLN6TSUV7+JtZj7tkJ9o2VVDNxePEfo/J
IpMlEYt+Ae4xEpW0vH02j9Nbk0NFr30g+LuXNPjPLd64SjW2q1HuG+ioHpR9OB+H
UY3FUZT+8aROPX50+ETvFP9hARNL84LsrUKqVMldSSK5x7NctC/TOMxvy9hRYOHW
z/9LhNa+Lnhq3nhujZqXuHJe5Ef0onsfP+IZSxXbxlUzVHwu1BwP/Li93ZeCJuJQ
3hY7Ab7WXhmxd2K7zIrLpSHLohxDo259UpoNWNO/s3pyCW9XRbpLIRtk4ETTOwwv
LctgYYdLkRVUGcKV41v2CWejzP4bGxSogeE/dhHDbZYDAJ63R/O9ZjeueL1pNYai
OT3rUOq3DjMj8FuHHdiDT8+60Wd12zawcEFIYoauFQ0IA6dfsKRJcOqT/Ip1ZwxS
CTqgac5I3TbqssXWiA5JRStFmGjBErlVIQFzVoQVSntLdygRx7KThu1jD/5uvNU3
PQsE15s0tLVqY/f3Tp8yHDtaELmXRuXaGdPTxJPziuGi9SaJmZznaZLGLWEcQKdw
UBj1kYqSsKGQyTwERhoa29d8iV4cTqrO4geAxyRrfdV2HuNqGY9ro8zXqUMsau5c
FGa1uK11MIZUAvZKyTEBp74hiJA9aOe3LWXDsod/d8LGoSkCGe8jp4yeoELsODFU
t//88J2mLoS0HZR44VywMpD/Ax7ShEsFSMf0VRFmnbMr8K6Y5dVO7dXAzfOpPRPL
XCceJhuqt3OHfdQHjbGTaI8NQBJqlHmRp3vBKCcAZqtzBFSQ86DxdYiEiySzOn1d
Ez/g1sGVt+w9c8WKhGtp5KtbwFwrD0EAnZEwKszkgfP6cTbCNpwKFksr0KOLBIks
kWRik9BaItZpEZ/NOX0ixRhMcBlBFII069Ql4NGFFqvZ3NPXuihJ4W4KSbkDaMab
8GjKta2DWDFgHDYVSTzVaQDHJUZBOv1ox05IfQGL5phCmVd7Qc1KPRQ+DrglNOPs
kvsN5+TYaUb0V0eCmHJSGncdcZljMUqqYrUOmf6Tt91LWcx4VbGTHVstoDgkwyjP
l64Dx5BZMFHGZu2X/ei689WfCYFHeILSE2KkbH+WtRf4abQPSBJm9Wrtd1ulicgd
hEYe6ccaC0ahtPzjmYsFgUIkPv/laYF/pMaCo8lgtd6Z67HNkkvzTuBgEkzVjTOB
yBtjwU6pL6LdPyQugOfQ5j++q/XVtgYYzNKc/pfgrNihOVPW/+d6GAhSCdaiyXMS
tR7KRj2utVlrsq5JGm+I3ccfWSiWIQVUSWTn5H2SGlZvjljOCTID62LQYP0pKuwj
kSxG6fj6P46mwJlPjAwsQe95N572TYf0pQMQJZH0tSKy8DkzfBAkL94jIE6q8IRY
cfOj8ho3UivhmD2DQzv0NU6pHH1n0JPxPwJaxQb9LfQkVh7BMxfkEBcbz8Me6HHp
axjhLxqwXkUlOo/AsGMivkRQcNG5jwreMI7gke9Ew4daM/kD7QimtnZSai6d6dbV
cEUQbA7d/NY/hUL3W4dLSlkzN4IQvISEjaKFKeedMFOOOW1KNyJDo9DhId8xW3Rd
M+nyd9zB2YaBjGUE0oMhJt9tIvgwshGlzDr7YlC1P/mNeAq/GAHrNqzzELi2fwRC
ciiPierRriEKys3rNtvUTbm1YQiepjKz/D5KYvKuf0ykoQrdzgS5EQtDGGJyq24U
hHRDYADerpOiBXTbwaokrCzmiDXDboST0HBjzlCheVF3qnFRloftIUEjeRx/Qov8
MzOSTp9/c89lvp7WiYlIdY5zhDD7XMc/fjg4rFEF4NDl+sCIXkIew39ycM+4HtHG
T1lYVYuGY3WaZsN0VDnnfUvHGuQQ6HEF3YeVQQRBc40/wYnpcfi+FtE/ARaguqSO
g3f39A/5xEUQJ7eWOhEfulmUSjDR/EujqktrsORmoOGwRQgx1+EdqCa7HIV+/DJt
dGTVFevyJKXZ6Q8CKlkrIxIBejkY4bk3z3pB+D/GCR/SjsexEL40geIp5QtwjKPY
ztpachTlE0GvSr/5TMzflISApCJ8n3MqM8Wm5EYjN9Gyd2oN0wCziFv7tetmbAKQ
/ka4H5Y7NEGL6/2m5ACFAxXrDQgps3DEmbbn664WoQAmxbABpv8iWZwhi2nuXQ0T
nVxHQIucWE9G5dtgXblXYRYpjLE07QI8q52RvGGwfH/gWbTz/S6DqoYMOeBYra12
OtFyaBekyxAtUC0WXmlWFXa5IRANJZh4Ckc1NEpo+QoSvz2nKgrzulIJZvPMZCDP
1fpyu8TaLH4Unk/hgTehHfhBVvYBYxDTS+/IUpQO/wfrOH52jmdvWI6VEink0uGW
U8+ho/PJ7xBC6tZ2AcosxGNqXsv002rjg3Pbq0EbDCUMWzQ3l7Kjty1MDmiSOmk1
ItOJ6L4vC9eWBbJnI7gVZS1G7y+80kDiUWtu5qHJhDrACaXk+JLhuuVaT6IwSBTU
r+m9zLnP1Ivf/rjL+DxLNXWfKqwYHTpGVqK9tO7fs+0hwc/OgxCIaTGUDx3mZMTb
qp5joxysodTgZPHqaMn9iUFYGU7Vb2Go5LrWpX3tASmTpGAIw3N7sRK3bjjcbpj2
vjbRS7a+J5H7fka3uwXVN+z+L5px/BkbnGuwFmEQ7BXnoSZ+K3rINrZkbel5Jybd
SDJFvCAje9xBZi0UEvgSQzmPBlB0Jymj9OUHy7EdbtNnWp9N/E3oQ6rAwS6kQNvU
Z6Gf9Tk8po3izqRlJBTK06b+UIJHUOV6tCi/A2mCOOYFkpWfHjRDWyTxlfpr0DrR
TMd43G81yjviuCQf9Y0yW9eRYeplAknKy1cg2Da4TSgOpU0t7npQMaoo3iHtGSEb
y5b3KT0CQv5A2kwsxfwsDf2uXsfE5VGQiHxEUcTBxMVtTwaCoF7Hf0kmP3CKEb9z
hMHGt8penWxi6WhTAq8P4/LUzWpGrFBMnRI8pE+hGYPoT2P/cZ76cfDkbsrQbjCP
lWt6RxZIxsWkfDnaVF+u67KuI+F/mopqXWctGv9Dc/Gxpm20L+fFbpqDVlq10VT/
W5CGy/Rzvkl3svSfwXmRAIQKopRqzTxV4A7UBukhaiw8RYHwfy8s4VQEegaTm9UQ
xiY87+tN8yc+H+gqEDZpbodYvNCphBhiMZeYq8TiBMGhXmtLjryZTALvAgrcwu/g
zN7uw6U1002AuSah7K61psl1wmkd6z6wV8s9s/Q7crwMb0QuhlCNdjUPhfq4ZDKt
TnTL0Uv3Hcr5sgYyiZcaSULXJkFis/EjC0Ra1jcSAyaClJAkkWwUtLxhySworJsv
y+1L5dsX1n+2AvajjCNWUq7o0a61w0qsArJ9rqIPHuOCwYdQVPejPPTNer3RLl9Q
RBycLn3D2rXKjRRRcibevBRXTvJq58ru17HdseE0/YOD+9KjQ2FDOt3TM6JA7/f7
5v3qHugw4vEBMDSUWiRWll2JDzd20y0jzObwbzBvlhJz2xQ+kbOFqFnU1Q/Gof1f
TIpom7YSodYBOKr4QSwCT6yPmuzkUasfGRUV1RWIe5LKY4USPlhv+PHRv+/YvosF
pVuU2nlU8pPea42okpI0W/HlViNWQUbb8v4vpL89N/lo39FpLknmTMfhj18qvIa3
Z5jaial3AICUeg3GCRE7SXb6nylUV8eS+umRhpMguGeW2D6UzZb6M1ZqcZqpARFY
Gnbog2UlptFbSOpcIGSRittmSR3xGFjUiZd7560nZ5N2qF8XxlSeqhjobu6BWdRZ
nsqjSeeG2YJPx6fq36SaT/ib86TTwOK/clxpwSxLtnWORJ93UDmQSFwE1V5hJA9O
6BWmVoq35dgkK6qUfpPex97p1qHxIl5gJesE6gyRiRflUfprWWUjb9g0284Vuo4P
9cihGJWHBb1Bm18qikr/fauvmFcEC+/vhHU9XHUk7uOX3F91wTlu+sfEGWKudGxc
wUdvqLE5qHr4TWAeRiC5FdVsul8as+dVayu6UBkmqEazTJLNaqGOpB5mWD4PsOlt
mPLJ6WRdZVgJmoiVA13HoHEhAKXYhq/QdMt7KX3Tf6ZFaJ7uvKBx7J/jcXo/uXS8
jI0vGPBaaOdRMdIcyuUjOVBHt0oxPpnVq0L0xGsPUmsbuHnUE2LEmXuYZg2ar7XO
pgVGNFO7MvlpEvb8fLjMdt2BdmxT1jABvm/HKSpA4umDK0F/9P6RVfzbgOdIpU8q
CFSmh1qeaQWVw99r6ZfaYhYItPdAPDczTcF5kdJUOKdRClUZfvQVoSZ9iIUptc7s
z+XdLGPydmkhiqyyAvw9lTaziyIhYMGBlfKIAOFMG0J/uefhZ74f6yzX3PhKlHFd
fOWt6MnPMKRtUzZPChF7+jh2S/esoqKY8A+X7SKWexiqkdfUdgp4moTpdPybIbRX
kpnCErFzRhRpmbvjEUZ+Ot0fSYB9u1Wmun7e5Lh3vOqT45dzhbDjb/sax4IJNRxc
VIkOSvf0jz78uGAfeOYGfRP8A7nGXBiPnWA95F7JoDF3ZJU0but7XqX8+LL57FTb
KO+Jz2k9a4FCAly3aIU6DXjp8leoM/0l0WbxNp2leex/kUC/if5UxkbvXKnZDadh
3G9/tvXOrgjScJZ4vKpPE2ZnToOD14jtUccVPx242HpzuhTBv8OvhxSvW/3sUmil
WaPQ1hzX3dA1uDfM2MegYSoSKCyPECXemtRsh2h+4uVmp2TjT8Bxo7xVPOXHWcue
2VzxGIW2M/Zo4sIY/G7Dy8xPrtmb/RyeTYntje3fei5eatYW3GjLQGP756T7Jd+M
aPt25YaJCwW02Y5nOhrrV1aAG4n9GqmSGONlkz2Dq1v/LctiRlaSOvUSXnMO79XN
K1/IN1v0ZVg9j4OSMeCerwofoo4jjRooSpRGoHcUcWbWcHOHKK0TPQZFmW70ZoEc
sQBAnGkuxbFu9OipBS6pGQJzpT/H8iz5g6YRB2Mo27iPpjv9fruGmT7f/KLqN95L
zR2TCr0aR9vuIGxLOWFihVSLvaxPWZc75TKF6VL1aBJtAo/Bo+yp3eJ9yOsaImBN
SpS2dkKuoO2xldWnnGaqQ1tMTZo7uQuqJ+AQjQg/LMF7Wo2Ts40IQu+++zbaXmey
/2Q1qQWfug5XRpmw+Pl1zjbtJXViLSLaLqqqfLWzUJftHW52MpfSTCVJbkcGkMKf
PeObG94u3fOMFQ9Nk8FPZ3v8r+S1wdfBUGrUG/gxn3mlKD63vOpE3HGAyfMrnhj7
Qzzmqlf9bUM+tr/xcgPkIKTBCqPpbwkS6bJf8rD1FnFplq4uIKp2lHKHhxQUkvTD
pmxtP9zw1qK7h1cN8bcaE7zdF+VJoUlIZnj9XCWkGt1gy49t3eda1zzlckWJPqJU
UwwpBuCTHOMVdcO7t0aINxxpBNKrkd6RY8kmH4sdqOfc3cY50klIk4y5055Uu4xB
vRclD1Ls8DuZKf1AKPfpUE2t+uOU2pg1eUEIuPh2NAbpduycxUvIUsYqLHBzvpLt
WtpxXGiq8GMic6l7Zo3ZQsGLpY0eAgv/ltvSc+I8WSQ0eEioREVRQljY0slAR7Bn
EI+5HSB2Q3wRwpiBoxRidOLumxL7irDFQiqDQk67bvN/4Ld6vmGSh6lUim/7u36+
wUD+aVl6nNnd83hYwA9jUwZ0AEtvdeZlPknKr7Ffgedq5q3buXYJwb8bzkIkdwkH
M9HErL1gYvLIwPrlr0hRcMdX5zNe7mOe/sLo/YfqJqzjnZ9FgfE2bM9vtcAQr0Fn
/fkWYKkkL55B+6bJKFX/at0lfpjIr6m7nT/RqJ0GynOB0Uit371+w6zoKZhVb+zC
6Lc4v2ICtCI/P8nV2lw9G2D6C3UMZEJ6DIw42xnUbNsWYQZgfO93tVsCTO2bQpdz
D1ZT1HX6EDkJRAF3ApWnS9fgsJSRhqpIOEUFIXjtoFVgmjxak+J+PKaTxeslM0iL
z7thnomdGDk6ip4knjfK9Y9tUOQbcSLhrzsOQLcYm50VZFV3ebSaDmGnouzxzPCA
bDAWoH6MfdT4lmbjEjLMUu6a52BN09iiu7JXtqHbEeg8y/4lJIqNRrhdLlcysfs6
lq4ofV+DBe1iQxIn+qsC3cX8ReK/eKhJsuXNA0c5pIAZqch0lYXLl9RdNiN2HnMY
pFhxroj8BLcLG08YiqrM9VLkE9hVjP+Ui1ltWEipjYzxBjubM7e8uCBLRz90xcfy
332O4pC0MnajRy6/FIpGLTgeVtFlAifMWrhb3gUw8VskdKBWqEPgc6X4/RsOCLUC
NwaYXiijzeoPz4moVFmIagWpXqCLwr594In/+ThPqeIDgxv4yF5dsmqJ4hm+S6wH
Kkg7hODlcjZ1xGXU8fHk1JMErWb9hbdYIwLplqN2/Jv6sjbWNwQejTBlaD0cZLzY
kKAa+1CTRmG0nI31BMW7Bg0A148s6RNFbMMXJfE3sIbD0hxoNb9SsuRu3yLNUK5N
pZ9nsSDOFAj/N7clcwZYkwcTZB/N0TPHbZOkMPhOf/qZyw8M+VLeSbC8y/YSypW1
qSoIlpk2VU/6wt7Md8ri9entHImoW94bs1EK3bHifhYIFo6XRwaYvon5y15cak8I
GJgIxk1T9ZSdHOX33NcXzvufnwS98bL1+ME7MqbZ4dnCpZeilI/zGtLlKAxQ95Dj
6BNqfjTQAydOu4sRBtiZQIqOjemBCs6mTNK0V8UESxabbX0osYQX9oLDlYvXcwDg
qnGfQ5EJHZVdd1xJUCqSUsQbVXNYs4/EAW9mrPB3TeDQowZAOs8fsXwM97ZqqlDd
rvKGG/hKoNIThWGC6VqPwMiZTB8muR43ABN83e9wk1Q5Vqqv/ZYye986+02vHPKX
DIT1WyGSwPp7FBHIni4U4tM9aScMlO5EzXXsr5Bujry1PgsGYnQ3+LWx1acHqgRV
4BSyPBqTy4J5IHHdpLD9s0wkxEG1nx6eaXuDI0KA5g9M5aHQDUeG3gZy9H0WRvw8
EmEH8hr1I+/wJENhhybCw9KUpB8BhssJTD+tbD/gnGo8Yh5Luk8RzM5j/YxFEvak
+ONu4jWS+IyqESTYTYd1zfGIvEDiXi0wUkFORuJMZ7aINmCvydprNWJvxO6RRAxX
D1pExJ+vD9kXalTZM6jX+AuBRF8d4eOXBa98VP/zZmGWWWbZnzRhRQDuemXtHu3e
BnyC+kbMNNEJfAAe6YQQhDF3E9yTrd6CV1x5nvXaT17YsvcUBQS5PE5hiBmYme8N
5tFNhiOGAIY08r2XdBgKlGSads9cSTHrpJpW4QH5TIacvM0OXuZ5bGjn+kb7dfnT
f93qws7TX7yxSRVPukRgxQdj9mpqgpsbJPfAAH1aqr286UXYdxCXpEgCRwr/yc+v
lnJjjCE32EPAN7RBqNydxy5mVcFXqsauO1sCSPiGq9qku4ID64LNekUQDIqCqoa+
2bq4m3gzvUv0TD3sEMbWZBsCxNZZnGBHdyN/sJDUiHEohDgWPGgJs39cxwPmlPll
yUA94Nxn2QtLUPgixki9yhXOOrdc1MRFC3Upn8+xdT93EEmqEomqmaxZHMPLhdfB
2h2dcuetyHFUzZCl8/v5aeZtcxqrwzuAYWxtuG9fo//Yatr6DhsXhlM/iSLpqzgm
R/dp3ElB12rkah4fg7eemZO/pWnGr6vre81IRynffvLCdcjh6w4eQyGF1NVofN1z
uZEpWur25U8KljZhkHrfsXXlBa6/PGP54El2irrr42oacHnxrwZ4p5qkG0dqOv7P
XFV2y2KUBfVuAEpTzgDQMMwrnXAKhihvZLpybMZCZ1BRCeSKF46WhUhSXXEf29M/
QI6FVqxK6kw9eL9xZYhg+n8nFKoFlpIcsrvZkGVigi6Oc5LlGOIRVwJUOMgABwIx
K3OeUYXIh3mAoQ36/zCXlRUHJ3UwmiBbGeHW8ytKOxerg0ZRsU2fJ40AXBkJOVWG
77hcUDBJ6zrmTFpLioB/2pksR1ceoA1vqHNgjJs7DEueWfvHjJDcGy4qtbFd9J+Q
lFjKQSnRu2xLsbl3oHQVTKk79VXa4Y8Ng47WYNjjzsQfMcTZD7j1L38lsrQPjvKN
9n6sjJXdjc8W29IaLTZoQuwGWzY+s2Bg+pVsjG+LYDJz5fgFQQyPu17e+o9jC3en
E+M6A77aI0/H4fkfB7WGx0hEqYmeA03euHlcrBsBiBB7XeNSkIiJFLrPGpmggkmP
kICD5J6gNP6qJ1yZGwZRwnj5WYUClIof+VKh0DWl831lFoZ2+uE0ks8gA4VDuiPr
hhArSeMRsXQ/J5P5sr9TKM0INuVCr19nGkC7ouzikgTckvJ6yMFzE5811ZDgNIQ+
RvEpldxGHe66Govj4bzhUdtbggVukHiPg62mAdTVKKrPWJjUJpr3avTtcvEuFB59
cdcVFurHwzOj0hAOXeH50/bBS662jaMf+CrETTJdibZ36xSqC35dKt+gIorMGQ3s
3L51CHGGfBzq1H4c7Zo8CH1U3mV3pOwD8U/V+fpbyjnsUsILCTM2pvHid6mZtvSV
GQRc0rkrjXjzCdnKngl1BOsUFvouBs9A5M8VdO4YqLb1U8dF3SpoY8oyk7xSLX91
vaH1/xzjdgeK5Qpvrxbegx9AdkkphMAXrl1+Yjr9tHmm5V1jYy2vmrkdsO08rjK7
ff4AVUuBOu4qUjmvF8CE+15+XsMBFWCarE24LPreTIXEkw4x39S+d/cBT3bRcB7E
6VmflOANrN6vg9jS5cYk4KuoWi4HKnBxmwVyZE3pCQS+vIRqLPzX6ov7IsyZkpge
JkuYQ9dj1vOeFeHPYWn95X1ZJhY4Aby0XTh2uysDxj6TSYxO4q1g9wZeJXF7Vfun
asGKa/OWfn0CZFsCIdttccEJvridl0+NKO7mzjBhcXW48I7ToFi2Xs29ARpTAuxn
czbG17usT9jjtGL9tM+guX/PWpoz9DiunNuc63NayrFU21SRmGKBvEA7b80U2vIe
A+4EczcmlkZoy4c8f+mRRqrHpMMoSw4LCkBhk+3Qm47tzu9bh1FsrN3REitS961S
p5P4gDXD+7/nWvO+IpYuUecG71X6Mr1MGHUnIToQwGVkBHuGUfz6krl4AX0ZZNBw
kMwhHUn7+br+0oQSRG+SBPnaP9r7bBrR9/r1g7q1Sw0vjRSVuozwNdZo2/AVRfTg
5kXlQQjkVTdYjNPC0YRc7nDBQoUHtIgNHRuHmdiHvSvfczX6IzYjJ8/rS96mga5a
7pi1BtiOFpbRMsjENCy97/zZ+dKF6Z1cAC5kJ05zsLw06GT683hhxn1LJjGksTnR
r2ffw3kp+FoksaV6JCsrbUN5/h3pXxa6OrFL7NB35FLvU8K6d3KU8oNmTofSbrgQ
hhk6S/lgjmr01vw+/rX9ToRz0mVLCnrX+5zTLtw4cxS2kaTvsErf6K5MDuMQcFCc
bxkSW+JcmeyUy8XhcIgALzsRpqcrfLzzV3RcM8TrjDwzNPcxpcphsoS2q/h+RknG
cjJODjy7yWXl0k5mdL14nkcHJOUqsE6EzfBKgK9Dah2/bLiyJA0Hn74aMsF4+APR
rDCrJjNwz1O4Kx96t88FTk6Tbb8f6yjjKhzwEizg6ANsdOoNDXdHi5t3jgxHn8Nr
Kpoc/5gdT/vyHOwFQMwGdGyg/0q/UCivj6o4TZvEy6qLw3wM7XFmSlAKoUfZCUY4
tTMdx6sVPdug0onsJb4XlXXUdaxoRmgE0dTFncU+Rfm7SBLWnMd7Ty0v/H9WXYDV
vGzu4mkqtUBt9nBx8KneVW2HHL0h+EHPHZJeV1FVSZXjRl9kVnc21BzUbKYuWFd9
7KCQsLWPtnK1uFCN9gnL1YJtiLQ+qhsRzSSL7GaJVSc1l4Yqv4ubxRQFSWTa7+An
IiVCwi5QzXQ4oJp9bCuiT70l08V7cvUzd1N9hCyahHTfy6SSz2xPHsrBqCNPs9Ei
Tk/pdyAzwPOKqqtKu8hLDCVYA0Bnvhx/IUB6ubxdl9E3mvkQLC9VM07VCPykRFjY
MbvfKCkE6LNjFevLVAcm1qvdKF7Jp+G1JzfR7tbiQ4ike1+ncQx5hnSBLZwzniEn
rU+KlnNFxioKdxdb2m6e9Z9ZfaEnFaonS0T2NY7wm9Ajam6yQLh4A5XELFcDO1yG
Wy2qkloM6yYllrGajYgiLJob6u2ttB+Pxf+w+jzDAsb3NzjfLzKEU1ZihupWa+ci
OxiDe6nL4Frl/ucVYoaz2KR3OckLPKvfVHZBYtnrICKm4vuqiR5i5xc2cIzwwIqk
euzyvTFVmO2PrQprmpU3Q29Ozq6VqUkzx9vhBC/UFZwQ6njfeRhEJrQ9EM/5wZVM
0GL3PDDEV3C9y7krOneZrlGqAj3h4fX9ewyJTQYjBcMBMGn7ivNL3vJUC2DpuIuE
jDSUeuNRaYKc1k5EzXktFiGKNYYtUESWpupQzugZ+qL8zpYUERsGEItzh2HxduI3
dTmWggy+lu5XiS2Pt2Jxk7X0v5sh4C4fzohNUCtr5W2IK3yh/GxQ5EUHvxYK6+Fb
QQiech2z/zjlPavp4n48ONGJi1fyOp44XRvy/FRetxJpHJ4NGxaVGYxVM90ja+ZU
c9BgIl2jzDXn9kzJuwN9uQz9nrZ3L/zXyeP3nVYT0mJozSxw4S1hNAUb0CZ2G5g8
A9NEnN5xW+fRY/mWl8B38VG+vk9ZQyxj6KmSwMdbfKPZTJGSWW1R51HOgQhNhuj8
OrNoSD1x7gbrijU8UOugMcCnQ7co5/Gk8dG7AcMuAhYRf3KpTbo9JiisuzzNXZth
A5kXewQfpCIErhA0er1w3ZM8N6Jh+j+IxMmr917RjaAJpqYEUTwEHGGnEjUow2k6
3gTR1bdQQne4i4AoWr08L8v51GvcDIg5PHW5ainrA8eV/AFXaki8aSk8dOi1UTVI
tGzmtuFGWOhOdthbNwkdDxnBoHb2CIzBofhMwx6RWzpZQOddV/E7yE2q6SucA8qO
Ddf7hQQeOQfXQgZfn2mcJbqQchAzyEOMFT6A50+iisG8AsMbIu8pq6bP/TEGdOnZ
/gwOP/V+Ldmq+G0xYi5SonVeUThVg/0wYEUcUfYEjBEqaVImFUaOrBVqXoE9cQIf
c8dD+nke4OIY2tXXOB+/ukZ/KI39l4OPOJZgwn5YoBJdO6lcWXPrAjQ+xcalFepH
FVtxnS3k+EvQ14eVbYr/QwE3xR9aI16JW2qnUngXiyHTxpnfjc5Qc4GdRXiJaUt9
jk/K9DvC5rDLvrPmYiehot0JIhWSP/pX1Vn7hNvAfR0tye0M8zAIrzvcAbI3lmIt
41G7EjmUP3pGkXxoeEh9/lUDHl+dYNnBDRfPUR4M8khcuxcO5izvQpPsbvAPsKda
UHtezWv5cD5U2kTQH10UTWb7Jab/J1Z1fiJV/yjayAmolvELdEIzD+KoN97KUoyI
XJp/cxINigyCIAfm+jP7+3xs7HygemYeml9STJQO8sKvnT6scxUT8nzTaNaW/xbK
xIqXAsW9VLgUrl65RwxCeYM2++pSTIMdNWjtatt9CWwkALyLw5YCB1tXSBVYWfWQ
Kb1tUwsCPMKzVZWz7vPN/mcfDgDShnDQrexv2VHa6NffP1UMm2aDvsj2oEpOfh7E
A0UqH7LWq5kHXEK7Rn4ZsYEWs9rvCfycslTr9RBBsMWTvEDKL736mSUMY/n0ipzb
CNfE7a2lKDougnmpUYCaJH9PjPZ7Xp4xjD0o1cDrqNPm1p7/dzPw198fTIgkFNw7
vp8libwE2xKk0q0LFWGliw5cCZ/f2TOjNitcgI5Vx7ZRzO3VCu+L1a6b43EWalLA
h3WaoWdQ9ENS7kQQAx9CicgwcJrQ7ra4f4n6Hb/szCpdYcJQ9j47wHe2DhaT6pbw
PNccC76bc8rB22jy6VBH7ABKYSMIPcFWaRnGEuOjG7Mu1Z7n6WNzF4FHrG9QnQCP
P0wvfSdZeh4L6K+ODutu962baVPb2S1ZBVDrVSLFsiqi/vLfluVOBJMZByb1tSB7
/lfe3sDwpaDzg4LMA33x+ZorgkHYvXFF7af/2K4+EzTOSSzPePO88JLQ+McMlUF+
BB2nI0gzDnU3AqcAOYWfkjkVzyFkvJgED70RoKogf+zhweefOzoxg0MWbxhD3ajm
zcZkO7W7tDIEOGoKmL95d+mmUvEVNYxoUmhwvUWc0Oek0X/VQkcXSRne+wCdeSCm
eC3AMXall4jZ00eaVZIONKBPFXa89FNnbNSBWetOZnmEtr1ZAUi9cytD1a+GXfw1
cz4cvPdO2b70BTSqoSNDMyxfpq2w2yT3g4/plBYB8ZirhSoylPNjlPRjcZf/crJ0
nqtP2rL6ucTil5ioI42kdKT+B2o14rU6aXnRLyTDEmRtwX7TlL474//LD9yzP0NJ
GjtQZHrGjp5iW9VegLke5IQx7Zz2/CRPE6z5eWXUYtWYDHLs4tt/RZi4g48nKGec
56auj8/xCsFuv0g8Pz2vzGvK6oFH8GmZJ+sCClHKPBjDtcOX32LtirK3dDtppfcg
TJx9PN/94pYL6CnuMQBCMcvAA3orSDyPzqEmY3b3ktK6/85sgusDNZ2woNqMR2mh
p1wEFxJ3Wm7Yd2PWxAdXh78cs0YM5zut7z6nkoKe3KbGESI5noKvvHuEgUXrwCKt
Jx/CvEGo3om18l+Ayji6hXlr22QNClhR/MW2s4oDZI40PvPspJOZ1u0noe042dIv
FSwfQUczo/LSUm+gj7cBKYgLbJEx4HI18EkVv1V7gvJ5oce1RbngDfBl7B7qpbXG
rFfGC0bLiOW0OdP9NoIhldi2NI46vK2UDJYELTZVRPrDqGvD0xS9/b/OUndnTO4n
fYWXooXy9rvCdnLOmo1foSZyLtJDwdm+iflkk7jIGpoJ/drhs/2tGYDheMyC6ZHt
Wp6uzv900Mttof3Q1ATnv2F/o3sT2Q42hS12eud0CaOSFxxIeqcxqRfx7yda5EE9
+fAh08Ima6WeALbJM/lTdREr7SYB+0NXTm2+KtdyvT5FzjrJ/V1eK+WMRZEnSXwD
RNM6X1P0kzhuWRQ5QekB159I/zjMpavbsip9ZjpCdcz0FpJnxVvPOKxvH3nFxAlo
Ikbq2YwQEX5XeTC2aEuCN4a2Hg1B+lnT3q3sMMO2+YA3/nNe3JuD4FjuK8I4xzY6
KB+jntc317U58WW4dqzVshxYIGspGEs/xkLGx4yOOYC8O8XM5pQi8ipOCEiIJgAL
QLZ8i+2Dp2sN9qfLZBh60sap7+dZmDBNzXVh6B2gk2AY422W5t5TJuScDagx9A5e
MfQhCs/iS9ekz8n36s+2YMRlqfyDpjl0Tmhi7iup6r+op5sCM3ginJtUEQBvnrjl
yit66zAmtth4zFz+V+wKGpQYA8vN/noC2M6qdf2W2r5nF45I7jEGHMZCwWLKa4oZ
6ounPChCruORAFiPOTOv60HyU9aIjznTSzey4ZCbu9SonNANwZjdQ+U5dbzyJXli
20s+/Xddf/iyWd7PV5Nu6xHarqtTXA7BI7X8WesnSyVaSEpeE5NK7OJP/DTVO/3e
0WLh7koBuFuMW9BXQlDbJMA83pcyTmuj4fGUaWw0vHcsuc3IYX98Q6MqlLveDgVo
CsgN8gt3n7Z+iaOjeziFew5n1GQalftm+dMHOTdXwv6cpj2f8ssuBQtNvABtwjUH
SeXVpG/Bgyn2sUikcu+s4Z53qzeu4smVd99ydcUfwkjlX6lLkQBOW/J5oAyrSG4v
LQtddxMPEmm9+Qa8Px64LiSxneZhNN6xrj1i87HhT7YaDsNuulzPSraowgRKb3ec
dVg6U2TWNwbo/m5BA5xzoMpkeGlcGsDYxe7XfJfzo0IC+BQVc1UabUXcPF5Qwc18
yD9hpkCmlr2DwbhL7iZWhreR9XjZd0/0okas5MrP/Tod8+VPceycMnaGCpLZiOeR
PmcnADX47g0CeXGsZRI5wAamQwQZPmIyv+8SpF6WEQkocc6d4nrRYyWqDbbnAN/r
Zq8y1XlJp3LWSnNXVC3o9u+rwLzReC7QKUqyR42R95ph3/9X9KFLnyJL/qSnOnCf
mtpi+SihN44pvCyrun9ozwNdC7cJpPGf9q4oi8xnIyKqpaMW9ebktSUaQ3WKj+mU
edUVr325MTBVUJBti5xIMjuGQoyfdIbB/CRgZo+5KcCuZ9AHQMae85BQqIb1z18L
8jzE6Ut+ZSX/BZICdjQEvzNtp+Gahr059e76M6VMNYxuC9cpUzfTm9Vk2TfujJxQ
KGQUNwtqkTALctlq3aPOIglyNZo6i0LK0BZQmpxjshCryu0uaGU6bJBSaeMBUu36
PmSX/2b2bXx4+aZ01Qc/5wPSPSMGkx2EYRWHVRJc+peKc3SEfRYgt+b2/v1CxBN2
Ug/QYk5dybWPUj4TanvwGpTHYMfWtLXRDVT1BXs1vm7LxEsoIVw3lvAKEzdnV/Dc
cs9z3Cd4R4bdBaQQYHG8eQ/uhUjAQeDNT+yl1wLIxqZpdjj8zO/dDlgGyXvHT+i7
FcoHZoR4C5+0cVzUyUeLmq0wdiGZnnfzQSEVS2wUsRmzkfdupFiDTqdlBMC3N04L
m6AY1dQY/RNIfn2lHW4Ic6NeWPM8d7+H1YjaE+lDgsQqDwJaI7Vrkf78djNNoKrN
9j4ZTRlCy7bknZGg0cLwImuXYPSkR1vrRJTv2B8s5PZHUhcaEBMhJc70XpzOGKYU
YfYJ9f2WhIOi7gwCxDZN6s6Z5fxKxeTrFKAx+efiyie+EH4FhVUvbj6DFSdDZ3ww
aHWskD/rEqowI1y9NEp4QsTHFk0VBLMT7yL67vMHRbQ0hT07szUGi7MNme2expNq
A+Z/kCQkEUMGAyDBZ1OCv30szNe5xGoV6j0MLbwPsjsVVn0f7whuCjeLWoGD1bsv
+ODs/MmmgDjF3FsktZnu+46kxlQX3ubl2dRNrY4oMZ2SHqvLcYgc/QNtSlMx847z
PTDcMn9sGoEDLX7TBBCAkFT+Vrsb2Xum5F8XUoeBqhWzWtjKE4BFX0kE93am3UNS
ExAWOoCRjHw6a+0SJ3RuQC53loi0ecezTkn43q1pFb5OgnxK7srW+o+EbG5QWGuC
93BK5TgnrDOnATC67GNSBJtJ1Q5RaUP8apb9daYYX8WtQ/vHOPWrl7rsmZEwls02
ZMeCvQtwxdiMEfSgh7jaRO2x4EhfCFuxjcLbDtmBxeWKT5gnNCTzmCTWhkTFL85g
lsx8UAzrsvhdPw7rhHQGYQOHk0UiEYqVriFgiGAreg5VLCEKJ2G18dysup5udicR
RXCYOoXfSg5CCvKio3cWNFfpdvqELqiMOHahQN/B0uRAIxKsTo6v80VMq4PmVW3Z
Jc43bFtjwY+XZOLk8hQvpfwV/zgCTtXw06Pby2VWa4HBgR1kVhXGMfJTyHEDy2uE
jklZW6FgQg9puasHmGAqwJJrB+9CfqBn9WtMS9vYtBTQfMHy5JA5mhtSq7Dk49nv
OIkHDeSkntohORmP0eURyTPwqMN8mtYY/qG7Zm8egRVDpBnkhl57u6O3GdfGSCzi
60Mvzj7rzH1vl4I8J4ktYvSw73J3arp1r9tNVJrYT/ec68eoCPReIQVIkvr0f1P4
XCylssr0j2Uzq+yAO8tUKoEyja2/ImL3c2o4I/TJyTAUYzQnlvEZZhCxAjhE8Ia3
SnnmNdZXPLbQLL+iu8rSRSftlOltASnhii0iAa442ruVDHrrYJ+7ywIGI7qbjb/Y
AZKIp2nT8Jn3ogNUh7WYA+WZmv2bG4fH/Ga65096ydJFaTVff3+3rQRyuB1ymE9i
KJwrt4Nl0Av3B/vuOAsJztLpHSi63mR1Ws7P0P9X6T+eZARyd6Qd0GYRGWy8f6/p
DYVWKQcBNF9TqrW5KQN0l+e+qw7Vl3xYShC3I0Br2BV2h87yfKJ/8YelVCmXyAvW
FV27yimRqu5n1Vxy8qaiYFFily8tlbU8wjGcEKfuKvhKYM6XmEK2lBWIiDxM8mFA
OLRNybcveYUCS3vmDUA34LzjqSVSUCd19p8nrb0wpCmRUWX+Q+ZOT1l5nISMdDsB
YE2ie0Cce/8yOwvpm0B7ll+0HEmbmDAYCvbB5PyKQph+D+U8akI6AmZyfufZ+ld5
bcgaheErgAaFc4lJVpEeyc6dSLWjvgOAUaaKYON1gVLPQV0nZE0F7Idte1c8bJj9
fNGwsYTN9xJj/6Ba5F0UEQMqaRMLupK57jxHvriBkOdqC13TmuyUEtLOEWCdIAf3
x2iJakK1XeSUSfJZEQmgU1sJj+DIGabr/lpy7rG6VmMtVevBs/9t61brw9EHgvhg
j/5uAS7L3ZtOmdiOg4pZQzaDaFtuxW+p022NnCj4d4Nx2CqqeC9Qc5So8elxtudR
mm0rAg5A3NDXILqs95Otk62QF5Vb7y8Sdcq539pxd+KUEfTMAKUpNuuCNczKYRlU
Ayh935+kJtQU3hCEAkHMlSkOIzPOTf5WMU9K3qvErh+qrrIBsXIdTXXD/mOTZL2g
1cEK5tpgg+HGQQqRtt42kGBVKJdxltpUZp4J5hnmxnQ6Nw2rtolmkVAPEUSGiuoq
IVz760I9BCAIB4IlVqn4dwzeY1Xr1h8xm27OgZo0IEtV2V9518wmb4ox6lF9w1I6
iPHYrASFPgRIR1Cn/1nWPxXQXnbvtSDelCl8V7ZsF7VruINqini/xuEsbi5XDSIh
29HNtlhAeL2sIvaYdNAIX/tzD9cb7Hu+tNpqJblW9rS0HCE6puuySL/MdlyAms2E
sOCx0UKzV1SPftsgVEicQQqGF0EUioi8aw6E0Rq9HGTxftHDWf0Y17uUkMBB/48X
pp5nE6QcQe8jUbK7wC5NiqOKVPJJtFTvNPNE6aTUSnhxvO+ljD1gzUabXRn/M5G2
HIkVSH8CySSjDVfkRb7VzTLqkdsNgc9qKXgWcFi9D3rVq3i6W/nGBNaDIiSMoqnc
luISwGPTESiXaFwhfE/mma+i2HfuKRZyEvl7zRt1AsKVJQLzep4YFXRssFERJhfX
BEfPEJLVDmOvra5Mp8LgpcFCsTW6Ny4MH+jD469thwnUTqEKQjvPKAlA615CKu9K
SsB/PqfmpmyKkrnrcnGl4ozYFXh8MzJI7kmJJf4+fORvjsBxsRNMyKMqc+Sd5+9G
lomapYYCh+qN6AkXaoY/ueCYdou9auriSyfOQXL1iVhmJCKGqY3WEUwJWTY8dsZH
EO/iO7q/3OcxBV2Vu7SzAJ5Sz4F1X0gp0iddMU4X91EA7HZm+fbeQRdb65m4S1hS
Nw9tb9ujNWtDLDE/DTUDhZqgeiRIteGq2KUZKDnR2k3Yw5/4vGiKJRwilf+yWFcS
d1lwhmVSkqzY08RbAE+mEHog+Ogt/Oaqi0exP+17uRyyglxifNVMYurKnIELIi6g
b2F4sLzqG8cU4QcIODF6a+cb2jxYnRKycAV50TNLdxzELO9jGageNuQqTzWn9Ngw
ZTjDbqAcK90fzey8T5bgObrIDe9NXvxYuIYElYb2qhYuGRSbG9ZLI91B5KesGYWS
4rV/kIuFcIrRd9zIMgqahoDKUnpmuikBILKAs8ExWgJPHeplrLeMqxHCOZKG+h7h
TsUu/cdWDhggbCdS//CdUgSsfYXdm3UGuLMiVEY6EHgPn9tV6aLFuKuZk+/0avbe
HxEjUxQqPBLuEFqtoeA1zJS68CxrknrX8TbU/BNSr/sv034bRP+LYG7pjwc1Dfmq
blkkFEsSV9kHiOIb7ZCT540n/1WLBcPRLT7FDcVlkPHRANrJ9xlGUqFiX3dpfP0q
a8ZWzy3VRgQGVNYVn6ZxY5/Wh9NkrUDmEt/v1TA2PdSI/e+2XDeLY6xNstK3W+hQ
+IUMQXtaD6ODEm1WxfcWPT2Du5tnmSWIwIZEjKPwNpSAK9cMuEucV3Ozc+D4/pZ9
9GIf1I3oHIM3ts+0sS5/3guK/c2W8qt/5iBQZJL5vK3/sJPNBN5SfI9Sz2JU8/+T
DEQHhXQ0RonfZdk6WEQ3YyPUJAqPHBwP/acul05+9EP1RwRVjMtGG4HzJagM7lYW
V+OSYaf2bwqRElbhlL1dSgJ3KWlPEn8F1Dpi0CrDQjYoyGdWnt+Y7jhmhxhVKuRh
cnIPwserMI+W3/Dx7+l9Xr9/oYn8zZgSPNBrTqg8maGUMU3kUwE+6XbN+hHZeZTF
i54LmJIfB9b4K0SGvwub9jdgQJ3/G1iVHwZfySYektuXiyHgD0udiDArBBRigRwI
MCrHXOw4FnLBOsnPoO4/E7ntQHhhfGMRiHcOI2nQHY9d2VsLQQ+sBiwx70/+HoN+
L5mof55kZ2hIjpBSOu6hpuMNfIvlaOGhurAwnuVTd+iUZ/DymwirAvSirQkP0x4E
QLVjXoy6gisSPGrqxewfnmIE6qmDxsT1L1qMCxY1tjDnJPkE3/Kg0Jq6ohRuKv9x
ryf6P2IvmQNzpVLn2aQhCZJxU+46zHcy+YaqC+sX+YzkU/iLpaHYgjNjZFdTiY8S
Y2AQuRgEjZK6UJkHZDgurbcsWtOT2uTKkkcnlz3Lz1dYfP7LZxFFrV/zGw9Nqufx
fgLeYy/ug4U3dX4gaDs/isaj7r7diUCLI8NezTNVfip4SKmfABLEOjzbKhWd7w5z
7fFGH5Ozlf6g/jYqhSDv/zRYU5KeG3USRv1mvmZeuJkhcAVQWSlswyflTAdKiu+U
/ffQPTMFv1tNbVRcrxeXSxueH7thL7dfRXOoHPdbiv1Mu88qM2a2JTqK5QWvEp5z
lRivgobk7GwCl9tuzSBw3gLI5IfOFJHlCbtjU6JwWu08I/vSTklfp7xBM/FBAdbz
U6O9BC2F40N5ukr4VyS/ng58Oy8GKN8P/uEjbED6OvbyE/DZc/1uudvIqvCGuoGp
Fn5B3eqCYx+U8YHMSePx3Xv6e1Z0vTcHpC0Xt1hZQ0vmg8cGa6eMRNcZba/GxxxC
cRSUn3N4Ld1UCkb2dQm1ShXtGzI7tEk9ZgZN6a2q2ytFZCdxR+acXMtC5yoXFrWV
uO4tFTb2Db8M1Vh7gpn0ZmRXJzQt0ydVQnunRKqZHCOlLX6UWkIGCucBGln38p9y
nhScKnhNvmhqUzb9w1zokIh0h+z1Tk9eH/XPwD5Yk5fgztNTJSMGFmPrvhcCtACS
JFOwUVSrWtn55lmo8MYLVFVVgiAAZTchmdMZldRb0o5ZiHUpcH5yIAhF3JFhPZhi
9VuUNElMZysdyQkuXYrK0kYydy31PNNh4LNFGps7Cw6f8EUh489dJIDwjqU2tciY
sDTGqCT3hRHfWFitqWoU0g5Lf1So+TdSpNrBT1P1d4UgWvcE/6J+vU3QLMzEUWj3
XCateVBD/WzlfAL/SRlACzvFLEy0HYeR8+XJ0QliWOZLtHE2BswgYB3b/rglGbfD
pb5BArk8d25Yc/T9HJv6lEwLLP3FWhRmFbZ+oTN7y+BPgrxkk2OsVtys1oe6Gued
iN2SGe87WDIQtAaov4vP0K17YlNs71I6ongpS+btYuV9n/Fh0CcSCQ8PYdJzh2eS
MB4RHPxKQpmhcH3TH31iew9Ry1KvV8msJYihA5o117Kt/uDEjCxrq8l8otao6Qz7
tZ7sKg/R9HRM+bMu0DyqImN+zbEpb4ebwJsQPRGCXDl3LoDn1lMEuBGam6BHY+Pk
GT8O2pR8XStaAoo04cnHX3D0u7gqRrrEhMMInJt5kO9HTFe1I8LdlMABsNKXPgtf
GCxoL4hSxKufqC6jeh1fqnCYoxE9mlhLJiPVScT0tjg4uUDMTf7CpjKrKKVAxqQn
yUyzQGmHaumkyIGmsUgY5lW8UufEOGSsKYSTb4vZ9LPOvm/Ndoe1K/ZdOqK2uEz9
VFbjNcZ/1CsPI/qKfIFpnpyhN69B/+kEyhce6BXGdWQFrL40088/QxxH6w+5yvfz
IK+o3yEuLQHZsmG/aFZuCdMXOLsArCbbn19RMkh/QrZ/G4ScnwNrYL9EUgxwSWJ0
/Kar5kpgEVkBrvQyX5GKPVBoHNcMjQIm6QBasyqUI8zI4+Z7QTK9XpXWd9D6BvRq
GwJcMafDJZgVfQrFI++Ta5EDUQ8xX/9JGYVH93wVpsmG8NPntBCTfod/SMBhcycj
OrHeDPJjcw+dOVpS0cYD/Eu6neuR9Xx5DRONsS8X43Q1Cqb+2pcuBZqhH+uux5z8
yoUPriVK8IGQ3YNXuZXF8ExziocI7qFUqgOmJVGEkSgBFrJ7N6UFgsBGEFkz08Xe
HwNHaGiYAzwFEWKPJM26y+LCOxCsl7F9Kjr1O2QFetpEbuld7HqDV4QiOsc6CMY7
p2GmdhLezzsVR9tm+sVsaZkXAp4W+64xM5gmaLrDi9ljZ69HtODrV6oDyo0gFOPn
TcekaSRfB5JZ6lGTZ8zzQPEnLpnYhLCB7q4kwGokerSzL4sNU676DMilORwTqeus
auzzORMWmj70tS7VD/r8eMJ3q6TmbekFsUW4aN5jKi+0jkv9F92bgJ6r6A6lAYYc
PHhYOm+/b+JJ/FJyxTi9eZNxeAHXkwpDKZ3YPD4v3r9MLHsLYW67KghKK+uwBVjj
mmDr3CufN8M5JU/iEuBq6cAm3TP79/W3KOnEUeirkxh5c6tyOyMuIxAXuYKbf3rE
GwNcrvOsB1+rjdIqMUiLy6ps4B6ssF4lZayyMy5KvZSUSzkAgANWPyCvk4cMBXhB
HyXlhi+Oh7SjANBAA7xcEN1m5vSX8dElDgv8DuiYlJX2frnXXayiSmzLc7dHLUiC
7P1PCtxV0+hA1USMpYDXxUZuVg2q4WDbTnpWVdOOaIry/8FsqwX6/J3Tv6KIBezy
MNV4c0J3/fAyz6VTL5Yeyrg/StbJbGJvpaZgsPrak4LDUwrLSnyQGgwNITTBlTTS
wKQAoKD6n2QoHjvsviUUKTWFSC+UfQm+Z11Hc/oRzYFytcy61DN9BM51wDgwlzvG
XHcPU/HZPpIewdDl/kzAvy1Sdhcl8aSv8DYrxKtS9PMO6muybWDUByrJYYi94KAE
Rtec+FiAlPq150XBsj9QUeFP9US2d3FZS0b4zbONlspNYwsMZpHC5wdBiHycqKR2
ISAhQ25PbEIBOwEg3bHippria4PWGzXV4R/1Xex1TwTgF6tPaYRxym0Qu/ZZVo4y
xZbMeATIGVFyk7YYNj7rcC8VArvHzQOeqnEjcsi/7fscy7JSN0HtNdMesFWaBleT
tKJXH9sYFjqVHrwYK1BMf5A8kRaT9oSzYb4CC8wj5+q9RaMduL/Gict/QwHe/iiW
dJhGBRhU/5ULOtN8Mt6/Gkr/byeCYOF+Y1cAfmXR/tOjngE5kPqTGnL/cFs7HtSR
8JUiCbpL9moN/m9krtrLKWqa1z/DxBkDflXJSXhYEgt4fCHkxP+chFO6gmA2jbl6
GmrMjoi7NzKa856p5b9sXgGy0e6ddNy3h/OikkbDPqnRiipj0mGMZZagqwUiSkyr
JTdtlbAr/xFGbS8HHHUS02NR8tbFCkWMvMTkyW+mIgB+8vfT+MzcA5kkgcqUjHT6
bsWLs/GAOahdzbOgmcTu1KBcMtkR1kJ+CgvVxuEP1Knz7UO6VIw9W7a37ocVCisc
iz2sp/cbV51cSMZmdfOtLYB92qERvr7FK8mYz9tpeNnJl3xA8NoUN1ORa1AOXtGP
Tkuae2e4HTPvmlpcrAQIxtRI6OsT9KQLbvBS3XerXpYY2pMyCCsnfGqacbk/95Yu
tt0q4G158y9NXlMd7qyqaa+AgP4LL0K8hfYNTaQVfH9SDKqwa+uAdS7jdl3nlTbd
HfoMC/U91Ulta+tcVODzKOG9rjMrlqpeJV+29SgolXX4S08noVKMlJvqga+aHSg4
uebWSrqOLxxKaHyl5by0hGTd/dESZaCQDJf6P8ZUM8gCQ/PO5vJS0U77cLM1m4U9
aUgDBbwNs4mfjneSSXO129ecGorZOJA6fhWhFY45HGSmBmEUaLs6pTkR8G7bTxUS
+tDVpLvu0quL2OD0h4+xQluXngEKEAx18l/FzOL21Kxgq6/0OXmAwxB9bikmggoR
zAd155/pRTvZcsdEKyKl1ep+b0911pjsxJRbYYWIMS2BrukDgzZenx2ITdPjuVFA
XQq56d8r3QnL/JK8QAxzM6OsDWnWAT8Jm6CbHlIKq4mSeOT2ohLZx+HL7cydvi8s
O0vWuKHiSBbylh33JqQaeIdTVEPBZqVjmG4Pp644YEeZ89Trs9c2/6sChWQPrh5w
ONBS8iML5PS3FXOXjRu1jW6/+kv6lvboH3qj610q5CAXUWc2QCwYERMBhojCL2ih
FPILGxTmZMRylBCHemvbEZBTQuB/BlQKqkECvWLZ/Dyo1BvCukTs8/eOT/G+rULF
UJF49dyuQYAScVU80P9Rsc5UfrDqb6jKJNaIWdjO8oxi7Nkfyh6vSs7e9eWvtB9W
JV50/6CA1dlLpudz2p8AgxnuF7uRbg1iJx/lBkjidQU9q4ZHy+ZiX2zwzRTDg/82
oH9CnR1jNnAGigbIR9JTr2ZCdOhXoLfIqeup3z05OmnTS56dBiaLPqgL9UZn0QmM
a1DJT1oTAcOnWvjjPlT30/j47kRAUlRH6mxH6xDBqC+K91YJRqz1LTsMBfEQ7lLx
aO51C0139hW29Da7kRjfdhw/jLAIcezQTJPtzkoHnictV05WYFMDuNxxVUi/2uIv
k/kzJgoSXmxJXrmh0ELmx+ef7d/2Pr2yUiEk4R+E8jLJVVdwNg4N68nQvqXv3tWF
GQApStJc5EtMK3OiZyprOkgoIVoScqY/wqx+joZBKT5/DCXcSj3M7QIeVo2vLwAI
hcJgx/5zjo4ixiaWSYqYLevq47FZLw0coBJVxHE6uUtFwN1IecbI9l9Ql661yYlp
y6s22nmA+WPexbDmnjDQTZtR2t8qzaeTfYTSmBxoAo0KZ2n79mDEI+1H/7P+GeIf
xmu5oN4Pgk3LONToFyfhxhyUEeKVtMLNW1mYxHs/C4ptUI8a3i/bm3TCKi5IAbF2
VzfLQtSFizG6tCIp9xtxeHU3aVUf2Lp7O78Mj3nFZ2WMRHBgSE07Hy48JYqjIyaW
iCZz6JMLJXAWlpYTJGsxzszfimzRZ3LL4Nm5FiiDEEVheOkAZ/HxpZz2mfLn5Qaw
qnXvCxLSSijFM3iMNM2ObwU1TlUfg/aPaZghSUcPG4N/rX3ZQZxnQP3tvB254pp0
IpeJBwAzG5TLG+SiS0haWNly36pm//rRbkDKRbCKurA5juvLtyMHQevyWlXwBMnr
uOmY+CL3JV3sKDDMsWKMK35RBf5q4ju2YcR3IZ4axJGt9Bee00nUAikHPlWQnpeG
CNtBbcBqp+Yq/bRBhIAh3YAB30WMQbf3j8FVJPFn/fHXkkC0p7W6C2DmPtd55Ko2
e+p3cQNlmgQAKQKGeQ7Mn3Uvi4vyRW1Lr1dXrXo89T3R5QvHDtaFs/rN5znnzDvL
aFt/16CHiV63ODcmAfkvOPcoQJ3yiVmFSR4LEUk3Aw+LFli0+BhHDcsJLl4BZ3S1
fiVIYmA2FGZ93ocX0lCQkcTc2Q6UkN69hZHYH+7B1QU1GPXP7E81Yk9VjcbOoAm+
Ty0QDWcRo5DsA6uYkgyIa7J5F/IyKBXnc9QBkV1cyPS5vFa1auoEUcJ2A3lwPVeg
87/sJLvyj+/Lm56rLbJKPwTQVOJjH+ZQX8aC1Afb7TPhdOA1bAc14v57efTsykmk
tVvrMeHQ+DseSmC5Yqn9JqYu8Z6E8Ur5tD860XKSfQ6oNcVQ7HZybhM+gz7bCBTQ
ZpdcdT2OSUEng1BrFxEv5fZQgzmAMk+DucHz0hEnkJ/COMxQPG19MjyDo/C+Bjyl
4UiVryP+ZnCqcZp+gsTJe/RZLsJJA+qysJPfIosJlH0/qio2hckma6gUCKVhgivR
QTHBXgArxWvNljOy+vZpFdyGRWqxfyT/exWGuu92HDmVsV1xltpbEpABDFWZgidi
flxM62SNk9mwBLBEHVA/3AL/DsFKdT5jq9Fv9DLcGaxqhF0Uecf6PkiT1b1lU1Qj
6V0/LQG5xBwKcgi4yJFYijxrcEpkoQ0c+vfT9yea6/7SoA3aH0DgyfG3K+WpGf17
A/1Y6JdMkI6A59qDedXKBK2ggfetKs+xTotAodYZX3C6RDfYUj9x3cl/7nmBo0Cr
+RGnA6eye7FHm2X8hsif5TKq+bzI0an0RKeWGMkMbgteroLyPlJBdNcIvkcrvTUg
3gknBgEO0OMNf2g9I7qNSMuWAcUmmY3BL8Bt0KDj2Dq1/Y+//b/ebkUqwVzLkHEL
qmyNlVRp3UusMq6wFpBNr5zU2vUyScbcJ/FYCCypQJlDIRfHJ5gjsRU20kWglVVw
ErzNSCyltLc69doULxCM4E2Kr8ksjBxUMXBtWjWYZBZ0nRqsRFsBGnMyn4xor9js
GXkW7emk0tuoS5jp5RMp5vEgpRZFxfUaMIDtQ9L35WPXj/4+MbW+H3KLWotX3Mj4
mSXaPVeikXSdwPD0N3/3q1Yq8SrbSbVnelKPmaW8GorMaKL9Ymz3G10ZSmfXBZQx
ex91NHCoRgWb4amMvcj1fWaaDbPRURWxDcVTFvjhia2g6oLM/2bIR39l2hzSLrol
4ESbGPFwAEgZIEWcaRUfAFeuGh8tfJksbZMMRKXyD57yY3anp0UH1rV0+y/zuonw
ZEwtavSLM0Q1PVSa+HPxLGJ4YThIRtXUMCJkoLJTRP2k9d6joynh5xNK4R+ek+7R
GFDLYwN2we92uqDevnPfg115gELM83Nb1lSLocyuehh2TbXGFVXEUJDOzSTFz0YE
xOIWXOg1iGjeiw9bQxSeHNgekMnjytZuuC66S4AEXV2unFhF0lgqfgo8H8UsN848
Y59MvHTXVEy7N9Y4u6uARGFt/zB6N9RbkDzaYKl8slcUgg8NB1EPVk7ou5Cm7hkd
tdWpc3h2Ubr+OZwLyX0XyfBnh+knnQ3Sr71HV4+Ike2t/vJAqKSh6KWPGE/mvMf6
LmoLo7goaEXwOCX5R1QgpCUyBC5e+TI2H89W3Came+ECsP9ZxEQdRBwvN8AgQ3vP
UCvDVqf/MT3Jhn5PZiPqOnAgJloXD22oakhEz4gO16GqiCas4GN4AWbJHr3FLGlh
0Z5Zd4Pwoq0So8lkm8w7WHjXaAcj3YIewCXrEk20LeIYwZ/f6tOWHjoLA+FjvvtZ
N09R7hSIJL2o0q+yq2uqoLT2SzYGV7bjMgVKJpA/5p7U6APPSI7ZjgtpXSrSUZqI
H1mzkI2L0xFWv3cqvgFlKeT30WG0u+U2Kp7ivJoyDzbv8VkG43/jn9LHJuP9Kous
qH6YxyVQDA0BjvSEBCfu6iAiBfY1rXqYs1bUZRhK09TzEVQetgGSHDPaHYz4nTvw
dFnnTYJTGklf3uJQ1+AHkgVem7DHxnIyDOp7zi/YCV9h/rINOga1NSKXsiztnM/a
PqXb1O7OtkHZFqmBpMXB11pJ5/ZcCz3JApFelCyKU99n4UFvHvXQl6yGmFb1O9XV
WYk4e6oRy5sg8d4NsTRHiz+vTLxL2SfrH3AUnrod7jhmr7gpOyo7Q0kDefXv2ew/
vU4mbYtFna71qper0Aw0Uok6TsjMwBDCOrBhSNXwRoy/EnRo7/ELfs3F2Zp1ZI9u
3Ei30XycD0GiH08gUAKvE32stamqG1CJKR54mvRInyQW2+WBqOuMqEtQQuZfgsbm
PTWFHogfovX/7uBnvao6rms4CIF0ieNgws72dzYVax0AkTv1ezboUnSIzr+CuTg5
ve11LeoaQiS1xU94qcGCY6Ovbxb3Yxw57pI1KJSrWR8T0x05Vh64wiFCEgT8MVjf
qUL998pjlMxrg6G+xnhAwo1qxLbFa/kvhvFOM/VMenN6S5zeRs2lVeb/JaDmn1Q5
Clp2sVj2GL8N1aNzuYbqwoC04aInEkcEtvNwP3Py4NkkUVIbzigwQX0+zdHrjzVh
Pb7GHwckTczJY/nLOf1pewZxyfXgJ6ytch05rudmOr1jN6E+gXPOqUYOBF4SxPOa
RmP4Hkw/fQmZaReYXzNrA8ZPfeCK/bN/oe/J2sKYVMMSlOWzb076NEQ/yBOXNbq1
XL54+6Kx7iCkSI1ofo/P2HHidEF0vCi/Uhi77aPx4GBxhsAmnMWNr/4rW+ujkRML
PMVhFh4TiNeYFjmJExnSvAEWieuGjJ+0Me6YCIIOrnlk7JkNElm+aKx84UckeOD3
/+teITbwP3FLWuWX2FpxlXzkPqb6odDeNOxineRnNHbeyTJSkiGidQF6u7c/dxAa
9xqyWN+c5DEC0gRS0F8mN3Dteknzdz+zpodSjCA99WtFr90UtXwT8as49Upos/zR
zmeV5cVMh3Kh7PNTyquKBqqzOYu+S0zd6wAre02yGapyCjuUAxB7uaWf3FJ/KVeY
sWorZ3X0YqNdjzJWvwqWwwAcJzd1Gw0K/jOLvazo1ozLrHO4Th/GFI1zGRBMuVye
X3BS619qdLGqEisNOEL1RMPFB6CoksVs1bB3j2W3ZSsVlshs9MuVnZxBsB2H/JMd
M8ITqWw0Gs7cU2FjSJquWRfQr1WYk76ykP+vaFFaSUYFZC7iLj1g1FGaScZkfbKp
Zuqt76+9P2kCEz3JVmT9G6FgV00+nO4l2MTP1aNkdLfvhviMN43sW71Gws7gghNH
GAcA+m2a99wxvIKglh+wtRK3bKVZS4u5APbomeK1DdbXVMi5koCHDsrEzdPCSVym
4PqSWYGZSBYShEtG8K3xYURZk1d9MpmfSjC9CZ6qVLE1OC9E2wLl7asLEJqNa4KV
o4pFZaELJncCf2XhsmUQf66RNYRJhEmTqcv2Mxa7MukYkqh5q85O5IXXOrxR9eEn
N26ZNpcUR1NeFBBjVwx1/9mVQpXaEhIFTF+jVOKnoGewOWYGOj7xi05srr9CvtYI
VCKOLBC4D184Sb+gTMDcrCowRo00hV2QlBVPKk/FmxdNJWOVzqLDODy6R2Gx9Y3J
KXkKGPvt3UnVGxwOkUIKpg0iZIPecQhnH4+RwwbOU1hnv/r8UrJzzy9P090m/Fa4
Dsc7U6TL+2HlIHOVu6JrSa/SU6ZIjhIt+10eY1FIBrQBblAt6WfVTFY6W6aFlC63
5FKD5D1N0qnhtZKJw1DCGi9A9epOFKaYZIa8//C6hUGMN+mlfWuaw7LnyEykCaQq
NOTwK/10+Inh5PONcLiNxKMGlCfKNMNZFmKAW3TPpipQGplcDlPCch8hK0u11TdL
e5SNQmk90Hthy7wvitg+oP9dtyzwE4V3FAz9EpRTT2ZtlcWT0MHsbikA7wN21FHG
NbFRrbPIsOxxLs/Pc55rmCW6Gceu73RpYOQhjznTe8l2Tqv6CcTsnCegn7ckPKZ7
lgPThYvmGDxzvB9nuUsw6tnhCdt84/CwHRKIYE/RrRMtto0kRkTugW4aEJT1CUup
haP7vcujq4Lpa1rqYEjQOYC/TlT9KZDxb1Idw52Vm+b7Pf5Gq5qYx8gFE4BQDMhN
MbPyc6EALG6dITYsBGBuFpM3vTL7jx0QPYvKm3ySUhSr0sLfI+dPhKCqUXYqUB5K
YzDqQCTRciPxRelf+LSoFb+DkKTX/O1hsjvqTV01j4YD9cSJNRkWZxQX/Bl9EG3n
LvlNL1wGUPs8UEnwqcFpFw/aig3hlq11dhnQf+VUiI6TH4mZUk9CnquTBAzNqFAe
7OfU3rdId5wMWn/4x6Bsyo3pi4A5MCfjaF4JuHQ8ZNFMXmFR8a/6WjXdX0qOcTIa
oPXd2c2hikmZXaMnPZwSakIhWjrKgy/qKEEzXTA9VmUufmhFWHQOYer4qJoSqQF8
QXQKLv9aSwcEu98/u/m3SMCIHjbDSLuPu7Q+kmsBjIjy51DBTc4UsuAfFSF7bpJ4
Oh6Gf5sjtxGDaR54n6sOrTqzQibGPWT3ryZJ6u3/WTCW3wN+ImuBmwtwo6jr1K/2
R87jfM4hlnGUxUYUl5yUDzRZoLimhVyVHWn6Mf1C/pvYV6hVkJaBAtAHZ6klNlac
ie5eREgmcdVXK4KyIUazqUu31xcrW3E2ktO2LR0+6T0bN8QhIJ9NGvNnkwh3aP5f
Uv7WpB4YkHxC2okWl2aeKKxMh0FZEmLvV2r0E6FJ+1VNBsTc0y46QipHbow3sHN9
S5VwlAKEwTJEzSNn5ayiJs9XmSSnJhNorTj9DwEe4CeiQfG0hxXyZt4EZBS0OnHF
EkRbQJ+YTvmM4JeIygP1B367+ARpdfQeMy6YT56j3l3hEydIgjrd3BHjrDX4SCsp
HTyg0xfPs7f47uyE4zmCCMwCUN2xLige6gHUxN2CBIUcL3ceYWvUzHG6dS4X3WCs
GWVWxnzzZFMmlA9jcGQF7czJGMVTXMGP3EJES+2gh7uZct5gNh3k6iQqkSE/DVr6
S4yHAWcs2C8xnwyMdY6Wy1uyfg9GfHMXkOG01IhEALdhodO33jiUObOkKbe7uHP8
XfLRqPaXI5qEOYuPKsXrS49rGAI7VaGInbbudM9e+2UWFIH5tmaiZZdaULkIHz9e
S1apc4zxED/afaFzY0WG23CChl5+DJu+MnWQ8hLNsQ2JW+j0ZGuazwSDAIDx1S/+
vyLW+TiqVPfalc1Z10D27+iIAXc90wY9xBEGNR36y8XLRvrnoT1K6Kuzj4JOyVms
0g5FCWIJWIbJuTYTPXYehTDEWl3pduLRjWKBEVIHrj6ttI0Wr3Tp21p1FKYlRyW9
Y151hesq88mkJ/7IBOKY93ftA5kWne9PtFNAisXmn+LcY5LiRzgtbEyPwFTL2nwh
gPWpRPkjqRa7YtabuvSCW0Xc5+lVES3EVzujTsy3tLv0bF8SxMyN0LQmeFhDiFRZ
Yg8CVM46WUy4mdKLEmWkBTF+UITSjQhFx/MKGjuZ/acYa+nh+7zJwxqgZRiMF8zH
vWo5X45Gb+HttktUyUVfL+HSfhugkOaI7aMJXZFuEVaAC02Arm51sjb8S83vWi8A
TSFe1our3a62NPwbzLoNDn0O02A/EC4Ki0txtjebtEdC5xnzHixppnR8a0IsN100
6uthq2ulwAzp4wpDy3PTdxfP/a+KY8uxcVdhulWtQ1gspWmHfmfHMx/MgJnHJXBi
tBhJ6WwPQjaPj0faU1q/y10q1AM02YVHjL6ZeJ4we7x9iIQtMdoJBZGDospFJ9N6
dPPNtNNKfPLuGdG6+8BK34lZ+u7pEP/v4gfUnsFJnywChZIQjuaKKU+6QKRDzkbA
4ZThecGx/e8svOHP957II0Vrpf2eqMHy1Xo/LtCbsbIIMyQhS1UZ3izkCJ9ZpmuT
59v/c4mSn8LMbZ1aHZj+Uw5poBHkQbJsORqUXZDFXgbYb3ivwBBgmgsLhodCs7k3
dxAe+aA1fXGNT+xj9mvl81wCJBzYWTag5JI+sNPiNU23uQ8StIP6I7r3yuE0zQH1
K6bFdl010S37O7o1eLOemwCzRsJkqz+PPG5gpumLycihFEqW5Qtl9ES7GYa25Lrg
h0BUufyd11ICQoq0pzOtpkWFDSMIAjsJGG2eOIKORMgyGYM8vFBQqCG7fTw7DNji
41kKserGJncoUlgNkm/TMqIgb8mRU5oJ8Dl3LRLKJplwPr17RARTkz9w+Dwv8DjG
Xq9fKwpUWYTPzomU2b5ESZERUzPrM4SvrjeAxnKlvyvekWRNE6gaW9Bh71tLAHii
AfpJ34GdVWYwkyycs0dVWNaCUMIpCs7lGUI8eTYEtKvZdtVgiU+R7iYNcn9NVofS
kUJVKtML03yp9fB54F/LvMmI7UmjBaf5zI59xiOBpoJI3e02Wvn25e7MRrbGLshl
A18lGwh+//fLSKd9Ibxr42Hlh5ZjTw0xRLYR9r67JhscbNR1GHbnl6CyIdIDgO9d
kP+1NsLf0MYcQqHj7MREA/RzPeuYEckhHTGxgNCa1G4ezeGXiYQUTDsXjX7rXSLG
DDW6e/M5SHFX5PUAA+PqEMHnE4Lz/6GIIPE33rOVGa9s0wPFI8beFtM2m42f0RIF
Dzhn47xtwtSCQdb2s6A9ARFD8wrRvMpJz7yEY/LPa+SvSTBi/Qc/wOPELAWnb5DP
DjApCWJLzdyepQPuicwCunLwT7oaQqZ4CFqQvGSWxkQqK+PSseBH0Qg2TG96HCjm
hMR71RSkAbSeOn0dqzmjiydF+Rfv3H/oCU5Yddchx4LPxUS+4xMvMMSOnPMgfeoI
9lgN0g+Ebxq4l8JfkytetdMNQHXKlD8CoODnJesAwyVn3K7IGbO5JobmB5SFpMP6
mMPJLDK7jVkzPKO7WsqWtVRcm9QwjcO10AjJNNtHz4tLe31nk08ePIVCbjRCEVKs
4x/T0Ms2Toj4FvHIusFFtu3kzA1sQaYPz7XFC3CRLRorWOKVTGNafUV0eDvfsOGg
NFapFGoUNEGjkFmu0fNoU5uyww8qxhSJzn3pduLnjq1pNRAgDwqso1n81YyLoDJT
v00EJa9+QsIuZGH0CnfETtbiwkXgFAwSwMjmf5IL1FnKeGeug/xLWhjgJlZDLdOo
keSbOEAJYDlXDFnd+x+OGZYMr7mpJZ7IVck1PIHCHF01pvkY4Av7+ieFIMfeWB0O
oGnYWYFpq7RfFKEjNm843VbR25bXVtxzIJWbkQ/8aAUU9LNw+sjLSO1IEkafy2nF
jEaSEp+7A7pWH7HKGSjoXmc8+/EGKLBD1o3kjuhPScSmf/TSevzjmbH8jvMtcsxF
3H5py3w6xkERNNrPSn8oDH+9mngRR7vWjKC5NgO9v/w93xy44kEAuZteKopodCNh
Y04mF6hY+JXlgpmoQWtQywWvN743hGbLg6mnCq/f75ldpfi0pPnYoqQS6TFX9Cki
f/hA6ilKXaLq+zUHh6fmAP/GPy4+tXVdvQm4axjpC5UQwu5a4LSKNh6F+llh0vpY
Ei3A+QrIaEKJLVVNnB02zwnu6P5bsCUwzBR3ksBZS2y8FcPFTQTa+u1YXpfhQpb8
5Dtmp+FHB1w+o+pxayB3ohDk3Kj/Dt2th5kM11iszUruYZaV584vtv/qPSohW9Xb
VVB10G4rAIWEqDDoytt/OGdd1kt/xvxmdbe5xyEBbWEeeLKi4GSi9FlyRPFFVnOa
0WR1jlLa8aMzPPeDkmom7fmGNdQ9tDbORTwhIhGMrqBC8//u4DIDgSl5FltPpSI3
AYNCIk9Z9DE2qfXQfFYovNjt9R4X5CFTHDBQ1oHAnMbJXlugLNq4L/wE9hXSveru
Ypz2vsc1xAivJX6/QBtvzstQAp22+Ai6Ae9jhML00Dfg8DIuY9SUSAxXJ0nzaFbD
v2ZbH6XwxlONfAHo68xbeH0+3MitvWjvf6tvYIFT1bzyvk9Wri8oKx8oziewZoKm
XO7IV3UZe1xlHV+3r8wf4JZjGdzOe27yOi9fVSQZ9zZUoHzD3CbQQdCHGOwNjksb
fIyRszdQE/lfxMMLMhRQBmSRm49v5tr5CzpR2CqWM7Z5gm6Q2SpBUqkb7jVwyHjJ
Bw56+y4Y8ll3WdckjULmDwDGZwZAfDA5Ji0At7jw/KfKaK3kzysxrrsb+2ZAIrmi
yUnBFTzL2hBax3UA1e9YQTvMOY9tVJUvADxz3RUQLH0rCVL+Wm6aUoOyGOpRt2RM
zmTMk8v+0Dv/CaZ5a5aDdPq4kmJmA3bT+Plp/F/dgc5WwwDoB5Y9hqMNOtPMcQUx
OmqRfnNK7y9FWeE9YY/xBN0HsjiFOLtvrPZmwym/wNrqftTOUGz2N2JFWwBYpC6L
/BwohI1oJH/xojQKv6/fXlyARz02HI+uHj9CeCpv/wprdYqTLLwUn8NvlFFS+b0m
FC9i724hkt8EwTidb+fzYcAmYc2z42/SQS0QujRe8EivIm6cohwLu7gGPW0k2tlI
utOWdNioO5zU+bTNLEWLQxnjn1yc0KLZstyHgTcSkeXITLGXnYs2uWwDfl/cmJsk
5sO+VnKq7Hlhb6KhHILNZiR6ZWgIOSFu9sRwGCVw/JNQUngbOo+LIAj+LBxogUWg
8TIWanKu7uj+why0ezC1q1n6Yr6zdrcAYmTJdzZ5VkddOXmCKqcH6u+22YA5dJQP
/iIQep21MN45O7RYpRXJ2PEI3rcmmYMmR5Lp996S8frUpAAxKeZ9det67kSj3lXB
hIUNaJ+nsAdAlnntPfdzXg7DSIiQ0U36gRghJ9LFdJg6tDNVLFCooRFKl623/9zo
XILm118o2YVUrgJ+2P+GkYsprb4XXCFIllBTBoupF7sXta3C+qRezC9ZZnde9fuw
I+WSApvA3G98hjp3A4h37v8UocCKf9VzJny2avPqGLPXugL5JB+R7jybdWE08VqF
RCy5SNhupO57QQH+RZiNf5CZx5zN+6lElzpeW9dnjiQR7puYtS/MBOkapGkuMOnV
oyc+XCjOJTKXbWB0XrtT0rii2rwBbNYbjLUjKj8bNOsblWWW6qq6BhqZMXe/Pfus
ujoehEtl6t5PKc07LcBAEBMSyt3jd/MoffbDxtXfuh5zxPYr9rHQzmXbZpz0uZwL
Ne06cMX781IztQ3B8zjQBxdiew6inrxLc6meXNsJ0nkZI/2oBfnScg7rZ1AyIorb
/oAk87kNDNTgT0twpLv0UiUYyigtTuvKxAiH+jLeQO9mQ7pFKTmWTo1j8ueEms35
JWsDWQ337/OkCTU9zF7x/u8BKYhwtDd7iVskimjX25gZpMUyIcgvpClRqGaNb5do
9h00yxnZQ66eZvY/Oa5Bk8eWoYEjvQq/Hc2DoDHIBOcTEX61k91Mnr5OffpUku+E
WW8t04hzc/HDofSdsxXAlXga2a42DnuRUp1DDW6M3EhOB3GWEpKo0xNbKS/gc6dN
+X+MG2HB8Uc0GE1PVJZVPGEHf4WV0gIVheyJjYEWAubTrpESUkfUA9lzRx69Yaf2
bwQVI0MDc9pqAxL/LK87C2f8HQIjAoHHvYjoRMk+dDn6CYH7KYz/96Kmo6fRcd7R
9cOUC+zgxoNSXKUbokpN9WNuFDtesEyzCWxbfnLBfB4vjKqv82u6IG2u2oW7Un6w
IDBGaXHxCtfqtB5IdHPgCDKT/K8ExkOfKWS8cVqvjCj9OLDF5ENkGnS7udJhGTpX
DtWzfmRURr10oQFGMpmd9y81FmMq++MfiqnKJaBnehMGldTb24A8pj6m9rWmnE7x
K3mJbXHupKs50mROz7IWdNskGQSpz7Sbw1xocPOhqlmDW8JlXZZkh2XYT2792zPr
hl9ucvK/4JVQFV6uSe8alTJ1t4bF98rRg00tIVHNPaprS7EJzjgZnlikGMPKJYVR
w2fCYCDbJViFH+mXVCUvcZTsyajQG6Ydna4V8ySHQaXPDgr/ypAUasyYuCoSxBdB
FDGAPUnu1V/tVy1cmr0HKOtGFgGH/XLlVDdyJU0wC3pPd7HmeXFWUjQKyqK2BNsV
IISyMk3LR5NiuE0dBgFp8uQyxw4oqSpIAFBZTUD0INOSoWpBu8x/qu6o222tNcwk
NqyUjTn8jCymOHnEQtnwq9hprbtZKvF2a7XKwbDkbpyqNBnCScpLwQ/+np7TSb6T
weVVL+qxMxEdm5NIhy9YaWYgOxW48Ihq3Ncj/cKPVXtoRyF9QN+wdvGmWE1c0j0y
+ibISHPBUCqpav2Br+qsjeDmzZWaxLsHJfpO6NoD1kHRB+8bhCvyolQqC7fzRhaM
PC2dmmdZXPB88bxXEcWW4/Wjz9VZ9ugTRvGunoecz0pgFOAe/OKo1x0Hkz525Yxy
Zt4O3xfDMUcw2Y6ViyaALD564hzlhy7c1PjetOKCZdoEK8h+/vhY6UVQkRQfuORb
gU6bO1bt3YjRMfKO99GVotqC/z6rX4vqVDOXvZPHdxhysoas0sJ+l1fRkiiQ3FXE
k2CAjpfYGNQcylETYcTPQ3BIjvaUSsbxD3UbtPFPBglyU/cDKcmNd9TwsXBzEUAi
+ybyNiSBjeJAj8fVN6sUuJYYyzI8LDZEd4NyGZXH9Cc6KGp+cRPUC3iUtXZycwNe
hkuFUQlemsou9jrumbb4kVkaSnJuQunngV8qmvB7DNso9bpXWZ8czphBEyQq3Rh1
bs+ACekMsHvQ/O/Tw5dmeeKbr2C2zmVPOlS2h/nisY5Ro38pwNZbWyG4jzt3+UY1
V6Dr4D0MQ5mpBMYwp53pmuhWluKiTpbDnMMcb2SNYWBJH109XdN7Wl+9VuZiBheo
Vdirhnsi7UoFyE6LPjwGN5yZMfZAtGF74nweXZVnXzYh08PBHYmZCjTssYBOFBYE
rC0DW7q4h5hNU96VK/e0koJgqb1WnNxNVnC34Mod1EXZ79k1wZciFl4UJyE+u9Iv
B4nn8G4m5pySaKz45Gno1PnH9jK+Z4VqKsgwcF6B+Y/BnoEgP2b42Agg7PetY8pI
F61F94tfN3dgs+rhjF12uLVJ2imBhAgaLCZAahchZ5lpKxV2jqjnjpEBH7x4PG3b
k3xAUX953mHr29b7ypghAGUSVH4hq0ysZcFY3pAfx+kNc2fB+2pUXiC6NpcLbVnw
1Mt8Y5svs0uQnz/O3sYtBcVlNPXo6fAaSJqASIXmtGHGMw3B8L6LLmbFEwLkb3dN
kju+uo9M4UvZ0QhIWudmWHYOeRjvHVroV3bUyDrR0fAjZbWQnKH7FomCIBpdkAmX
MNzbnlbexhvtlVicuWsNaps9GQY4+hZcDlBezSo72V4Yg210fas1gnDlDsiBi29u
mkQHRbFbtzZ46PfZEPQjV4E+n4rkNbjzQ9cGhRc0u+Pkac1csFu4TB77YyG709b9
pdu3Q/Z7JRE94p1UZjXcIR+leRwSaCOev/FCYjFH5l0WQCWO3/GwH6/zX4Xmyc24
mLNClawD26ZGvSR/8GIDEy8PyjIbdFqwDOlylgirwQS3HhPZ91RBeANqtfKcO1Hn
923bBZxgcIyN1mZgbp3ALJS0HVd77aDLmRA5GWyPZPg/oyLTA9Brrnw9/XUwXrpz
c8R8KHdS5/eNgWaQzklCV1kLbqqS9MnbUlT/xpYMR4JZk6Dmwmy6V/BS2bo1FmMa
Y9iHJ6+06EH7EbidIVaXBohet4/5BqkMMjiQ+EHbjwC+cacHsVjmiFQvXYsmDQoh
EzFfYmXM8MKGlq6jHqfE3S3WX0hEhArsbOlteUJW7FsB2GZbNrkJVbf9qW5i+1Ld
+UcLRr7B24BFBSAxyRvsHPeon86qmZTfcx8KP9S4cFto18NWXMDedlY09DDf5RY0
apkRcXjrbqdoiUw7iP0FHHP2h3LvALbY5BHcNT9J0Jlgm0Sx2tPhepRVO5BhhRHA
AYsZ8n6fvGRMDFijO5zLHTlgHASFDfoaaoszXJdhb7GRgNxf25i6+YyDrkM4kzu/
cqZMwu+uOmGqG5jZ4BCg1Zacu1d/8njG/shBKqVwdh6Anz8Qmoah4PyBzG1rCv66
8r2p/WQiNRirXsETuvgz5zUt0toDIIwmzf83ehnLXFzC6Kno8s2x9RZLKJSAhR9q
UTbP7ndfbKehRvp0m8R8R+6UBhKreeWrzl0mT/HbS2ETvRJCW6mGYLjtBQ8J0ZSV
uwH1UAK81psRGrOaPYVUgwVjDzLmyKzPbMiyyVoT1vJOlfWTFHX4NKhgfaEQqj0M
+gX3rm+JDkRZQt7TgTptSwwYgmGvF5bC+4RPH+LSp6tRCCoTMRa2HI7SQbyprPL2
lGNFlxXUmgihndIpID5HKyeLAoJsd5pBffgAtNmSyEkFuKY7OnjaNIOxfbsbHzr5
XnCxp9efD5k2IoXN8iYffsldg2vwwoH70v/Ti/+0/6XXZGoD+0iJOMTj4beFpU1B
zZkl9WdCUp21X2Laea2kR5tV8IgSbKO8gmPZQgSk6WgsMA0VbEgo3W70ipU008ex
a4Shi3R6CfRDJm95xMtBY50A8r2meF+4fP8DCt1PEjaSKqdAsVIVlG3punx/O6M5
p+Yey0v51qXM4c7N+q101NSZDU02xzZ5V563e6e+/yVcbJ3iWFG4U22GAmwHAd/8
DbdqoRoY6Zsl9SUMxgCDF3wTNeY4osRjT06nOxWvW530peMqfw6PenQvS0bftRaV
yvFaXJK+izoWTxE2k0Gt//dfkpvByeaR00REa9d2x6/Sm82wvRZepi8XlgywOXs5
3GjrsK9HVjUmDVQsXfAkrkn5HvquIrydOJKjicoaomraqTa0JWkNwNwKAC8VikFk
MN73QSE+vliXvK7s0qWTDFh5vrIAo4MgJ0o6MAz1lmWP6nWFGi3B3CjvlH69RT/x
PSLlsSRqGGa6fJ1hmqRSw++PBG7HoUv//mpppQvj13ukx6X0ux7OjWSeHoW30nBZ
5dh5Uc/ieYYj9yielzFgce0W0G5wMPQXUjL4umjkesOHk9J4G7Nf9Ql1GuVpgjCh
6uD3XMLiyDES0Q4FpsjtlbZXyIwuTwnUiIOT1IvhhPu10BTxQPsnJ464awyrbUw3
uMQXU290AcVGB1Nmme275bh6DkGsLHJmWLNXJSn9QxNPra9pXi+7c+gy8E3HnkQQ
XXWZwr6KZE+HKweah6gjcv9ybFuFPjObZXaONav0gFs1bCl7HeuDnQYcy62cWvGz
58kuRIJuDLfLNwLR1MgDGO6SEu4uH0YPMVQjQehDRlbEJWcJEUujZaWAn7OvFZb9
s0jJZcb1ZP+qBPMnFlNX6JBVrOwLU+UF5bwZEHTGoiNUrZZIVVRqOUeZqGRVzexb
8smtD+i2Bzb1BWR6KksVFFEUz+069Sdk1q/BFO2/ZqNWyfo1YXsgpVJMMfA7+fQY
CZh1brzYT7dfak9CyzDdiccRxg0KNPT0kIFIZoz179TL1TZ2M0nSOg0GpOrwWfgz
s6yYWyx/JkITc475zZD6T2wBFUU4fvZLeGno86hZq3rsvKMptWLry3SsabAFHUmr
RcIA5b8PCnzH3ckJamqPDotRsuYWRLfRkOAULtK4GIVI4wvo90PxQFd/WELjIleo
Egd+hQWnfQJm4JBUmJECMoASBakZbyel0Qe4DE2YTlSz0CGoVaPsc9SlRKO+SDJm
IO3Vhb14fu7dgK2tMLdoJUxbEgx/rx5ODGl/iYVmT38v6pj7ilxAEe24A5L6V4vM
Xiv2FhjxZ4woZyOZj5pRLG75j0k35PWugBvXj5PB4io0+12KeU8C9UvLS/RHjgj0
k2wu0VtEdaCNrflYq0tCzox9+o8g58/xpyRBs+7ePgT5Xlli0E29CiNqzCOCf8yq
FyROEkLSujkVTmoXsjODx0lS4WWAH/Ec+5HYNbmngnY1JLtGtroLgwkToCJcFy3W
FChLRgMP5g/tiFO+xrdATKss/jW56XaAT3W0X+Tjg5vWKRipTpEFye1kGZhAb4Qn
A7UWOOXzAi9oYlDg+0uaw5EnfBYsn8+/4TUdEpiQil1T7lJSEqDJgpQRwoq3qxTx
hfbxScTHhaWk77Vnw/+bgW8OJ2ud9KiQbLhTuXMAYN28u+xD1Aik/LWPDc5M/f6i
x3d0FmYm+/SjhQVdboD6VOFmFI9fuo8uQx+1VaqrLnQKVo0oXd/8vlBz46k48s3B
OJJc9RD2q/6qdQcz043Co3k8gBKqI3fVEa9mxLa0ry3HpLePEl0JXpQM9MIbMgB+
zkugi3H2lXqEA81GEfg8MyGkRGvMjFwJ2Md40DhsGWZKjUQwotOlzmPASxTxGzQ3
h34yriFpjgeTa12/1w6k5s/6eHkUqwaUUqalfwcQu0+yP4iWhR+0FldkJJdYFyDd
DmIsjdBQCEsxVl7xb/JiXqvW+atFLPj70UjjTQ8DBrUUUQdKDdSaXvsnn5hcKC0q
yIiC80r1WylFQbUPfsmc08Jlh7XlFaWmsy1PWdhfllnNOoh997PMkV4fXUmHUJs7
TWwNSNv6PrEQmn5mVjbvZ31H5b5xe/T0MudPosff6MYcsbUp4rAP1w9UGXnuqhJs
r9914X2wSczOeZ8NnUHHTUf4bQ/rk63A1OviII4elxvArkjAhfzkn83UwDPPy6vl
y1sXwM+T+LJjKWe9g0LHGEiyFvHK4imXGvQh2XWfIX2gONf4mE6dEXzcsz0dHKQB
NBQ5ZRosBdNSJoLs5pbj0RRPM6gM0Me9YHI0fLGejh7GiMeYJ/OerIvjmWwyacCK
dUmQ+cfL4E8JPgyd7b1S1PAvGLoZQGdv5tEsBuBKQcChMUrfMXWGunTb4OP8qp7J
UYicO35z69kIQF8EsqljvVsmHDv9xdMWhpEvTERXFgdZSdHzbGY2sIFPpUWkuNMj
cnzcDDAGhvtxfNcI2Na0W3FAqQ9rABYEDCmvbvoitc8anL4TExznHPXNdm/t651+
noDT48G1XRPe8Exod4PReKh8kxigD6PLeCQ0nJvnA8DCnfWuLc7X1BecpFXyrNgJ
nCrk7yfMCCqHgWJph+A7Ulkl2hY8tFBrRHcmVEGyx3xF7VXrNQtcz7lkw1oJzzPE
XeaqEUVr07/yxnIIxw7NTYv8apE16WbD5CwLH5Z8/TMN/5ZcQapKlMuiI9Yahoxx
rcd+9UUJqWIuci3K8b5DJUiyHgEydiKvFfeq65zErvOyM3+5bZKK8QvKzmaCn5fc
1+iSY7+bJJAePHmISqzfWTHYorQZdiOsX5BwvCqXgIOJuSTVrY9c4NqcRFx/twan
gvx43p1pu0EqyEC/3xb0eb9HUa1f4ODvtyiYww0n+yTdiad7ILbs0ae7zZ3oViZU
9idQyv1wb7ze81RgbV54W8CS55Uxt5cBQ69G5s4Vg+zDnHgRM6qSLA4QsIB2n0Ei
dwQ/aVo7xXhOJFv88176oREPcixhuPD7Aig1mPaEhKhvcSODvMKn5ohEvcU5EKXS
i+F1pD4+CbuhALPLeDyxs7ccvLAZvYBX1+bElvBtFeRgZdKYJXoSMEop6ZuJA1r5
KIAXyZ71IrfKireTmID0ucv0NmZx+TZj0v3ILI4MyHDU8kqDOqQlnfxYrBUqypWS
DGShIixkxBDaQOYZj9Y5NoeQEzrc5qURjkF/d4EqcYtUlNoQR2BeBb3DBgAtrV3u
6PgszQ76A7v/dtOj1NzbIWgbGbZH7uST7oQwn7RwAJrTc4KmrY498d48S38vjyHM
4ZC5Le2gUCqdwCY5zNGehU0MerugzxufpDuLMgQca61TN8s5lm2V811PHEv5oB0R
otna7cqQ8bhhDY/ZRNb5IJf0ugzei5UWOC1vaZzvnqtG3iUgjfYZYMGDXyWP2Qdk
GKMsyLVp57zy2HgsHVPPrivnXd5Pd1fdTUbpmQ/RaIyD0EWbcAnfsoq17h6q31uO
AN8CHdL5hypMIOl9JL5nIdwK1+JHBxa+q5Rc0CMTG9b1V2spiJaZzB6xm0cWnLjA
r7qN0bsXDRRNP64KrEyg9ItRL3xMr98wj/PKDaEFuJ0swbSgztX5A9oQfnG0ngBU
vyMk7RqqezrJxFv5PwfmKcFhdgDAV+VgE5isa6An/1kMSqJMQM+U5h5yokWut0c2
qu7OFhHYBxKYS+DtQxUFm2p85I5il7CeKH1+tPgg1h3mrLZfOwO8LfNjRy5HzlVw
29NG8oLetasr1SWDF85rHaxYkwMQ+x5pU+in4b4w76JWDB9bGmvjaKJYQnaI9rBk
StQ9rf8b6BjGXtaS7NWAj9dzVj9yO/f5OCw1pM3tW9zzFshcYfOCuji8IpZYfoop
t4XyyPbBZSJ/TOKwLS6jp/C4to1x/6wzKEnLb5/UHXJwJRoPtOO9SNOX48dzq5HO
5zQtCLdLtfw0okfa3Oe+p598G+bg04XhDme8saYDU3ROf5XLsnE0ji72airEdoXM
Ic/k3wudp1Mamz0GyLz9loTF0ywFATj6AM3qtLlPRIZCsj5Ql0p+1rOEmyFcyca+
KarGsSG4FoTe0lgdV8EA800WYYnuuD4rcp4eaKCv8+F/GrLQJK/Qtb/PpZG+IDAJ
qynLwYjJgZFMuPKyknjgjR10qbX43bfpnLLp/wcoGiGJjuUBGhI0diWRhR87HzU5
EWVjjVQTPkYNG3Ut/e8vEH93fPj3IH4qkUF5TUsCUdGVgjA6d+zeruxhaMd/vhiL
Eigra+dnrD4XF1BBRvdm22L41pPhF6wmLUnzwQNcDZSZ6FAEyqMo3+yzbl7WBI3O
ZVExnnjTQCkAcVgdntvnLrP7LlGbmTEHgGSXyPqMY8rWlHoBRX1MNu3pPUyASl5d
AiObPsRkqR0WtZk3TzOkHJBgVWPkuWIkoATU40A9W5SS8mA/rWeCPjBTjVtG0Voy
kOI1z72gHY/ueFu54cSeZp24m2a1dpyotGyD7Stfju5I7kECeag5kZYbymb2UyVG
7x1Ugn21jJ0U8Rsb8G0Pgkk+1DiIya4xwK281s/ILnBGFAnUkkY3Oh+ZAQulKsv3
g+M7+yutf2MWszCY4D2BsANgfGNkgYKl+JZRm1I+x1X7qwJ8RCrVrbplQonH4P7S
ANcb9F3IbzicA2juesyoj2eeiloEx/dZpgP5yWDDd1q4SJXDXRaY7Z3123vMCCVh
0lGA7UbACspm/D4tSSxdgR6mpMLQ0Arh1ACBdk/3aeNqg2agqlcFS8xRBFUNazgY
DoXyBrVfZCtRlTaH/y0i5/MjZS3dekxg5llpERYYyQB82WtNdj7jYI+mie3nkjTa
oy44JgN+t+ht/MGiSk5F69IGquRWecd9ZyDNW9wgWHsrB1kOlOROu4o93/MsaNJB
OaL9cH3S7K1Ghz/3sE3tjBlOYdqJYsnV4i9c0X8I8X6KhAaBPQhnLhbhm3OQrFlf
iDsSKxOH2gm3YbuQSKwZBomP8JX6nbcP2r/OJJWtpMBwBBDOqF28IaawnKOBgOLX
u6yujLP6DGaCq12GGZpNDrSh9kvD5iTJuPZuxr2Zx6m9abHgeQXueYUX3u7gaZiF
1yuzA4kbIRhKRIRVoZxr3b+6gPXEOJabRXWiRwdGbvuKF8M0tLHqlDeErnOTSKjd
aat6Zcs13cnA2RI3DwcDiMvLhlN1U7WHJUiVyyKVDgwrxbidfuT7hxA0pPCivKZ7
TU8bgigAgLB7h3OGR+q9qgTBU/Dig0dEBkF1X7NaBv74lx29C9mjk2NCBddu7xBE
lFhHv39RA9j1I8v+5XLaq93NKSbpmtFuAYX6qCHHoHzC+SKU5Sn4wsAtBCaPjeXg
9moWxvrZrdv45ire1vwEUYlLyiX9QNOvJNPviIpMS36nlNeRMvsFK4drDR6PPhlS
eqMHGUI5HVqrkKgrv3yO7OKECnQxbL2NB6XLoma912ehlbqk2vtBFOawB7AnponQ
9dI8RMJBSJHKs0Ns72NJzkeu2a9trANnylvSZ99kp8yd4FezJsKTVDicq+E7NiU2
WrId0+gmWs4GJa0zivRWIC89e2bjRw4Nv5Aboulfu67NlvbJTh5Ndw7HVKE8HaXN
8fReqt5H49y6dhAn37U2f1a0Abl6NJ5eD5kVeTiRVdnkrMG+vsONxTFBVAKGkf9Y
e/MDgELoMU/SmP/CAisLAWEbRELKytUY35xZ4sVmdgwZkVO07oVz11MB2qiAyOvW
EVQlRKjZl7fzwig01+BWA1fKYlkq8qw6VIyu/G9GPPBHNP63MX9iicF0hqxE8D9B
2A7kvsFwVAfLvSQKLPCA//8KK5+ce3bWOp4g2rEjFLCiaRd4eb0zM/QaHw4ZtghQ
/NhTRSB1Kf+hVrxMnQf7PfOawQkN+RDetViDjv6kVfZUstKzi8l55OharNx3suhP
Pxr60qtHUSvxcX1IapsQRQzm5z2Cn4gpS9gGbyBvyMyjIJNwpoQ0y2cRTGSCuFqI
xQ3xJs7FycdfXSKgkdg05lMP80U/T2T88Xq3VWZvLiSG0J66lJl2z1EWKIxr8hPp
jZpJ6hXgk0pzQi16K+Kf5mmR9cGF2c9KdLEUF4dFdMTt/6zkZ8t4brYKT+2ZfGy7
VqAKX1ePeGts+YttQKV+9k7zXqm21OO4i7JdEQBzUbf9ZJk4tzxyAJ2NGIVkwyga
yuWXWi8hH6jU6Gp9YTc/c1bsedU5IIrIzbvcTNHDAHEC0GpRO+jSd7YrzUbsKk2D
W4HRwnKd1olNX7pb5y7IaLocn/XFL79Eq8ZLja3WVv0i8JVMSsvszKSLlcAcvLzz
vSqsEBJQze2D5ksxSJ5ZgXOgIMG5i6khMyyEqfBmF03bvGdsc7epU3p1GMr5N/Fc
pa45Dzgc8ebFovLgZRPWla9XI6GCi4XwpRZFcLobe/paVs/oQUSGFNKPnciDm3iu
N/wZtFxeR0vNiAtI2JbAFHZA3cJt196b7mKv9nvqDvzKROkLiLB7TpjzGbvXB9PS
bQI+0l3if0P8QYT6w3A74yAS5aQy4au2H1Vw8qOaiuly+Rfe5pQmaLvx7mY3yUSv
HsLX5lgLIZtmLHTVvQ4UkGztU8Y/Sm5Jojm/yFYtUswIU/DjeNFqrMn4SVaXnfU8
mlzBie45MCF7wFKhgWqB6K8p4hfjOACYO/faABslxzkqNVfWkNUu5gm4bw8/bfuD
pKKwH8CDYw7peFicE7LqzxG7W7qIkvgm+OF/EkXtTB62vnGy/Q9DtVVrXCoqucG7
/CnaSBvq8xLSPKi1wsK7zJP2GN62tqTYRz2g6xw0rTMYOLl5dY3M/k0QI7pvk2or
WHIlUx+XQMrqEKrnkRIhgFLYbaBViFr3DhssDCzpR40hR5PVEERZVsBgj5M9+1ip
FgCfVFjKyqlnzkbRvkU3oLz8KDmSpdoUxRDtmQBIVFAd/sxnu+JoKKFrll3oMMW6
3S4i4PnF1XQ5JnT0fGzanL936Pu3+IqUoIjkyVO9gC4XLq/D32BRhefuklmEdmFQ
8wqvE9Tyk2FxJmTjikUhLj+FM6xYuvhdC2I46aIy1V6nIZFmWGJ52NXCY3L5c6BU
5eKdDqul6tKIv+kdZ9bony4KZalK1z0Cu77fV9dEF30LiGkz/af2c53zm+sfP/gx
l5Jm9zSaNiMRLsOvqX5qBCwhaBvUPLjwDOnW6rYCSH4/Zp+GLZlzwZZkfXXDwiGi
KZemTZsBDnpjy2nQYyscu8ibGvh5ItHllqk0THJ+9ipXrrfqyNJCy6A+Vgy8hs+o
qiM4giF9iVpxSP5baz77ATQ6juTwR5Jm1QgmhuRBEJt0fGDXEGrFzGTkjtLtmSq3
G4Ig/FFM3mSdparfGWDEf9vwcQ+0DHYEwvVEgxQb1RiOdbwUVNIKFRn8x5Z35lrM
sHH2fOPaon8SXT7bNYUdtWUdRSpzKl43efA8+aAa5E+BWm9nAv4x/Q9pFFxPQQYW
xOy2XFCbEKSFvt/E8cH3WzcuGumvRT7GTYW/qJtMPWkHHoPcg9+ggYp8lrTISdUF
e/sqT35oDrHbiYGAuhib1TQEWPytwUXxW+JIvmUT7Lob7y21Q95mkaphsYK0u8VN
lrvDu20ZrFyWBcVyIcE3Or3Tt2/9J77z2wLbt6FFEp8duMdTt/m8802BbuQ6Vb4a
IF8BHISY637iJoeYWbZIJ1KTAqqHJiFV22imHfHP0EBo7od0BwfRbRn0XBSkbzJX
plJtcdvLd3LT1mMJlm9fRSntCk2OIJXjPjhM0nf6DAQ7ERBFwbVEIHLaeOHrV+Be
`protect END_PROTECTED
