`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mPf01rgLsscO4GqOhO6vR4DqQ/ImlwReI/U7N17MhtyBdd0+5dUkUu9pu0JmbKD2
PXM/edLVQ895mylY98mVIs4OZPZm7UovgU/6cw4wTsz9OpGBuj8Id6ovuRLN6KNj
gc7u+VuuikV2BXVuLZueJU6NsDwpWZ0GGu8tolEqvYKWDCaW6uk1AC+TyE4tf0lq
TolResgorFfY6xzG0xap1f9tjqD9jiPiQnSlbZuoBIxnRgRTrRqsXhGVDi5DYiH+
yjntTkGOAOhj7+tPmsl64Wr70w3IpiztMUs/2HpEm7ErSUcrD/4xZnJ6VDrxTne/
bIEM5QhMBVoJjmiHq4WRmSMZBm3DGndwZ2lBqnC4bqPoEwY+Nnh9/0mdaD5hE/aj
o+oN5W8OVP03Z55kj/zFmV5kJhFvQlN96nh7+7FJJF0gnnLZ74MSh53zVqqBOHg6
Nh8Di+HCbC8M0wiFpsoXi0guhUDV/Trjg1c0IHY4n+wEoLXWDMky4yoeox1MbK+i
BjhrU427tHTMOnNIVfk1u2ClCL4bgSI0w0iayysyBLdNmNTrMSZBdyWRI1iYiz1X
mJ4T84HidUTuTb/eiS5KJS2xeky7hxU2djwS8pomYGV66gd+uD4gR+6eEl1tPrxg
eS9ob5FfWQRiw9m4noKKpuz9FzzThrm4XE+1s9jwuYtpnq0arf8FTWn3VbAK2uSQ
z1JtiOOuriQ0Ab6znYph0FhYZBiEP6+Ppu9cm8QITcqpJuBTofLoNZK32RbxtzeF
WJ5jSsS7zSboBtcZsmXdlD4RGd9fQdbHorqRRz1w1qX2GHUQ3lqr2Q24yyk7MBkh
EfGBoYlZKxwgcxMK8pf9/fzVrJ3j9f2fU3+EZpPQ2cLwLHVJ+3DFJGFuwUlFKDqV
msfY8kRFDkqMHGoZSvsm5u4IfA84/eyi/ptopA/mM5D5KvibglgEiVgVJlzvxS8O
`protect END_PROTECTED
