`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nxx6pZzDVWj3YA67POEUuYi9q1Co5LYW3Wp/GJUdmMU8EcbYUFIAgRNUvR+7oNjB
979lbW42C4mMF8TQgoAdqD7MXHzmH4mhh5xzhhyXGqqkMt4grblgSxO6KLqp+saa
Mfm8T9/WCJ0wNW86KkHBSchrU4Xc5oRIGG6j3EMbr5S/aGrE44cqacKewKjV+GMB
eT3nyiLskKkOld5WAQbmGi8nkx+Iw+scT1D2+zxXOGmjviBICw/mBH/X3VJ5wRBu
TDbaJT8LmktUkcq239d++DbnKyGJ+WEFTqkT5C/zqJ6ZJPNQjyubqoKw18xxt1Z3
FeUvt2exEFGyavIsajPmjv1cvxsWf08OBBeZZimeOlO/LavHk+UAMZFlXCOuOEM4
0cIOIPAOuXWWR0ELViv1FRNDGnaeiwvPT/vHgGF/2WuKoEFXmKdh5fCy1NuUdXpF
8GhMUfYN2f0HRqH/6TF7nGryDSb4OANHKXFkOn0SBnxfZIbLvocYyhodG0Ohnwty
SwzFmWb3wjgNfHGJXtn3rWvaoqNAofc/Mi8sXe8Ewdm3iVrYYmS5MKtHXYQzbm7+
mQxsdyZ4awhje0CAkelTKQZe2bsn5m/QOloI2zicmNGh0ngmFsIcahgLWFCNG9Gv
Rif+zqR5RjhUJrX1jK1iy8rZ6IvER1GGUvGr+hnU9tjPWs1O5JAwHJrv8+URGftS
fSfOGSeg+1HvcUxgDyJmHsDcKQajOAVNJ70v6dfRSX0=
`protect END_PROTECTED
