`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Npnj778gIDIBTCLEp1KFpPmpVgD6yxXhLx0qFM3/lALBcvlF43Henqlh8XPGHaqv
MmnyZJqmS4D8mIRlNAwjvCAwoblrNw7i66uOd2RufmocDNdI6uo6vYHP2vnxXkOt
j9P55WXs05lDejNb9XfG2G4zCIn7r9R22BO8WRqorjN53a1YJqpkcury1bxLiU/B
g5K6pZxDBWp9f5zOa0fnHdS7r5qJJdlboh51FCJ8fFXf0QFX02GGN+WiJAamZE1V
1Yt9cdUuE2YEXiGBaYWmGYP8scaEh1457oGlv5z1ZueKQPqgQPocjKyMt0ZRvM0i
uO419GJIujav5tE7Y0BSdhfp7glqAa0ZhQNsUnnMOHr7QLVB+nMYPAs2rk2SS78b
7DsTuzy54Dp5YSUiSjJpEu/8g6CXlxSIIYru7niZzrReNXjZ748yxEKfrumL7SFs
TkGDdTaqb9ThJ2EZ7G84lol5v+uLGkuNxIXd6/IIOIEAnUrmCjsVKKjI/jIN7N2A
NhdZiF8QUbb4uFNcLMzLB/G/brstYpmf7ustuSTsFaoRomIomfkDo4Iil7TtYe83
ARlx83XHdPrkGJpAtTwoD/c4OXS4njLTyTDcL6IzTVUy3OyTZzNH7LNh7yCzr5MT
RbUZtRhpZ/i4zT/+4m2U8vJ2Qlyhjd3w9SmyqoYwjsQwBpsIXw2KIm29X8XUvs8N
tegroCzbeuVU5l+QCS+Y/faC5mDCMK1/xenOuuxAvUdc92Z/S//dOckAthDtIey2
22ASk9eE7tvXyF+pEDPzC69uJjTZM9+kwnhroZdhAvuoy1TjNFDIWwvIo3HOW5+7
TLbrtr977Z0WRbRNx9++cTgW1LVNK9Of0ttxHRXJxeTik2nzXymg72c0ewud7yfJ
UCKVr0czjWOCgRL+Yvo0D/u7KOWveZDnlo5bLYCbnoUicAJ3RYML65u5LEQQtukp
jsgTBBEOXS2jRpuOYD9YeZZmK79X1Mdp3LqnD2UcPZDejKnsBIBBUsG0mz2s3fGW
ZgBoeeltdourjEEQktgh5F1Yp53ZeYY77xHuHYjGJ+Piwd7iF8/9MBgJtDCNb03q
iWddupXvM+b4pw5cNYoTILWz+rSjg7UYhwpDvPvHHpdmckSnDWQKCU4qFLSfCxLB
hdpy6vrcoYZgUYxyfqMDMOKlh8L4vdBxonhSm5MEbPWiC4O9NQI/qnow0OqUNwA7
31msEH1oT6DVpDNTPq2i1XvSCiceKytT4TLBLYBxm0qx4ooENXDxs1pkAd++sI4/
ZjeynHW86LAp53X+M/LtviI5fzvMtELybLzz8O3bRi0iSIWRqciQvFmbCxkDvL8I
2676UaiH2twScNBjOrFfwIztvIggkZBf32MS9RMTW6kDkKP2JcuCkPfhjlGDM51A
e6jOB1mCKmY0fFVGLVs3M0tqXqky5dqjkI5ftvKAJDgS3y1UIAeTEEJEjuf8UaXz
Qk0uV2u5rqlb2iL7HuPf+S7Toaf75uPqaEnhupgSHA5ELJvukxmT0PMQw7Pf72kH
mrWrb3pkp7DzXcwlKfIVc0S6gPLWMViTWWg3QOU8XX+zQ7W8LgevHSBHHcTqbgcx
04BsaNjbj+YKpyzRyRgyFl4sFnPKSuXY5e/GXXJB083dM2Dcdp35e//Xzzalc3uh
aqh5NcT6TbeQoxwNVvM7rc4MrXnepyYMbnDkYnQDphFNweZAo+hvdOeIsgDLbvPO
/JwZpMlHfcj1kKuNIJ+dqsSJlpvJTK54laoxFFbmmyedmDf7qfF2FwL1Fi7ggF3w
2YPPJBTZnVmTn3o6aqXlGkzaaldFCp5oaouWf4pCZS4bR6q+FP04a9YXJMG8ysn4
heVOpsEw8xnIE4FUEPnQBHG2qmG9vgYV6KBs/NwqT6ONAwMqORtoJYIbbQ6BrIDH
buF3UZgnOAu7IO3HkUmFMECyoHPgNq/7OO+ELFXCTswc1xiCCLHpvX5o/aacRySC
YFpVUNdIM77mNPHMsYSQJq/0ZtZpWdQX13ZJvi827ue137CjN16DgN17iU9jeg+g
aEE+FyTFJj3WZqj2htoOxZ3IJkCacA758g9LojIWRSxJIeaGrt1GD4FuT1bCN8xp
x8S/odjBGCu8dgimggj0+YqNA45EyJ0+LAVvUdrjrd7MXLKqiG9MCqRpM5GrLZMG
CPlS1X9KtogYYMO/xoFNNgF8luC46qlsqhBQplqbFerLNoRYC0xRbq32zSn28u3K
FHWe8v9D4q/F4x3sFsPNgHllUAkvpDTvPIFbUcRftGX5fwriUy50NabNU1hiZQBs
V9Z0UxYsXvClLKK+wBrsz6qYVENUZl3Bu/PkZlkQ/h4qRooL4yfjgcx23UKt7Rsb
J6hFs5tQ9KEW/7bARruso1twJlnjpIQvwli6ZCswiW+NXrFsSmMosj+JqIOapeVz
2dqUdggdX+ja1f2btwB9rqoRq/xI30jKqJRX6R6sd7rfgKU1GWaVir49qHHb/9+J
bVbjwOTSNaYi6ja9jx4n65daA24pZB2OnF2kp8sX8ZD25ELrR7hmlIeRs+BrWD2O
OZzjTYhdTll+QEv/iK+Q+t4hfLURMFW7jD/BSJkxL2CoAs34bICM8NAI4ZJPqUnz
D/pL83otYrYF6cNmLbm8XAEA90bBG3E+vMZqiYMAMtE0Fn/UwyWBb6CppL75L7sx
BtV3NmuvqQSFOsJS7Awi7I6Dk6ylLId9x93u346f6EDEmFPDilhkgtKsLhp+56Ob
wbrWKgFMi49EnVjaW3wxV0mYLq/dPY1IK5zemdPfa6O2M+1ubtHERXCdiYEA41j5
YQTXWwe61kEi1qjt1JwiVPM6KdphOxO8QQzC1V5cuBHs7pcg+Bgf04Gvsb/ZlWI7
AvanXZf69425rSB/49LumIvPM034He87SoW2ijVt4XZdf02+TrqpxQuxvSDQ+5pd
`protect END_PROTECTED
