`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1WkxNE3iWXyI+15FB+1nkPiozaGXNnYJg7Dy/IpIa/56YjWofureZ4/S6sVCkQJP
YzDDvuNLVBwpFQv7Xv1m7diCgILVuIBCGRJoQz7vKmSm7URQ/Ze/9fRDbhvrIYNE
2bjriyfas02hZWZKoylsOd+p8p26rkKT3W+mIejBCoxn0BYJkHuGRQickAgo3N8C
UIO+jwWxpOp6uOEcKavS8uWV6r8rtb9m8WItOuP+WBEqPgSg9fBv1ZJIq7UxZxpl
atlmBzdYnRNpX5YHTf0xThM7zwzsY49oCMI+yA3iop53owdL6Svv1rYdtsKVOrsk
EswqOmTFLouBD/fg+Et//WPI+wJem+9UHJx3LTF65t1ltLZCFrh8TmLQZuFZRLAY
4ysBfZvTJIbTdmG+6f9mphXfO41r1FsyKKXu5bSn67r+7OLwI5AKWI+vZcgae1Zn
`protect END_PROTECTED
