`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
csShx8womdT02ddxOVNSIfo+p49SGwMGZby09mLsp3zD78zya5mNurysGuXtmqAK
8EIxZR3EyLS3RnDPKiPrWsW34pLvAvdkQGkwydzo4Ag+GLhQJ0lf5sVJ2eBRikoJ
lM2jSk2wPDp2cN3Pj0Sm0PqEz35YPnHpkYByFk3f3hru8CshCBJJz0L0nNXTHYUY
MjxzKoLWKXStIEgfoa97aA/5GUEO0k7uckFXtLMi7j2f5V6mGrVsxWRB5YAOfUTZ
+raho4fJNryB5AuQ3eJok6c83DVdVmPdied74fCsGZVviqRzf1HbTq4DMeeaMlXY
51db9TmOQxaJDqRUe8roaH9rBns0YzTTgbF9ovpPfCwpTT2dZNixT/gi7qyGf8dj
21SpMXcCCyOet5T++hUx+LY0WC7adzYfm30uVLyL49S8JbSiA4y9/RsvimYVRLQB
GjdAWoGyMryCiPWez2h67Jl2AZYhLxUUGXWfjpdKgytYO1nDV5Erlh4mNCJnjL0E
ZGEd7tNt3bb2BmWzSHLTxFJSXM+6HM3LH/aUCCuCBfW5OVLETZvJ6wNal62UW8Sn
Z7tDlrv9Kte4nq+nLXjBQ5HL5gnA/4Q+k9I2IVHFkXhCj9dtJ7msaD+TlQT21ken
89bPdnrhXQRoQ39dEIcxOlBD30jKojduKsacIbnL/XW0mrn9h3EgcVXwJgsfVQW7
rZy5Jy/b5Z+3/WS9urQIPEFQAOrkCnHXV/BRB3twIOvcTZbNThgOqcGBuE6Qw5Af
Uivg0SuRnt8Am64+LnFblSpi0YSUohi0UVgIzfR2TPhYoZY+RNZM5RL66WC0wgoS
T1EBzA2+RB5aM6C6yDMTxaKqUN4/VWTZ8cDW+jUxPeszPlYu0VFlLdcsdE2Tasva
qWwpMFIXrFzWoZCQWZNpl1VOeCOgkgzNSsoCneU7tZnYr8xeWbgknOC/BzCkoUKz
00xGeq598qNpSJwI5Y9u2BKatKPyQiASLvMX7NIOaXC/VTXmKprcM6Qa0W2zMrrR
uRvAyHg3Xo2g1T6JdgnsuU6VoyqaR+xiB6f/QwxbPVpojrG2V/sEridFaXrBuqjM
SN0SgyxmVCa29yPZ8wvcqKYrj8s6HQjfHPEciUv0qSIX0DmoGeMHwo5CqZYMyO+c
rEvD+jY0eQwsBOftwJnPbweHSDrZ80oHrAfVV2NiWIk4pvgv4LXpkInSHg+zCwcZ
iAhOC7KvS8+MlrH1/9EyyKppmGndlixIyc6S0fmxZJWi15veGYXVRCDoFBmr/pIZ
BH8ShjzWy1qxoOYHMgIaWx/3+3uAYNwWv2MJHLLy2AQ2M/P2ughY1QoJKpIscS/k
Zqzm3bqvi2tzFi60CHQo4kvB1+WF0qpnoIfGqanrX9XbAF6THLOqa3sW7BG0uEJp
Lz7nIVv4UluDv8J0G4KH1joDHE2jZTI6ml+JHsU2royjpGHfv4ck15KdeHVGjYe3
`protect END_PROTECTED
