`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fmzzzSEW92aYmkElmtlc/7Qoosvuk7e/JaaTgp7Ojj2ddy3INjR6Hw1vVfaokCy4
uVMtGqPsUjr0OYjfxGRUWfZUXC09v+9hzCbQCfvDDISPXGexKsqpcLPhVq3gCzVb
k5Wb48JcbORu3AsrGGgy8czBNCZR6IvSlvkLqlf3FA9dqEXYiep3pKsXEK0F7mqV
DxWzpDtZVZsk4wlcp8eqgbl1mq9Eix1acRG0fLh747tDavjNwz9VT//2Rs4aDMlh
GTooq4kuNWzVHt6JF1v4qXKlpHxHJ/Wf7KwE+lTki+Jei/htJW3RRk4hosCjfGCc
m6jhGP0meOjrgWfx1qQb/c4BbIWGMMv5iORPwl60E46G6CI4lKF87xlLrgUyG6rv
Vl8xvv+i9wZPwGk8X/DgIg==
`protect END_PROTECTED
