`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OlU97YNKZw7M6tTg4aJh9Gbkwh+PL2U2azONo5/8aNJ2I5CuUVaNYbiVVvNufhfR
HicPAjUcY1cRsK6CKEfplhzemkmKuGG6RhU0Ppvs3+JRFmsGvougwHlYZXGmWxqg
4yaSZY0ayB9MvTDRDIs95XVN1m6bZYBNBNZvtkKueffsbMidmumFUI0kB4+RBHt5
gn2Wg05nbM3L0wAJnd2RvCBVbLV81g6YdJ56cMKe7ZzqPdtR/87gWOYgSYq7ReaP
zwZDwF009eVu7Uxl3RUuU6ieYk7Jr0wcgzHUPEQEwus2NRNLMxzNZsHP3pZLOcDf
m7PK5OXTFSURHWCVrD7U1fZbPnUd0l+mDQgE3O0fd72VHkGAWjWof0clJYjc7Wqw
bPwK1h4edItF6MYDj3BzstDip3aGGA601KK+ouV5PSqHnxNu30pwZjrHWYary+wx
+JdwPycDKUPPuzgaKEoNhnAShadsaO341s6ipJsutVGcLRhtzHd8KFyWGCBtVPDF
ExoSh/VyS4E2bHVd5zAMM2GM4K8uW2iwwYwuqpKYsyd/OTdBtpQszLFZ3F7jIII1
djkw7X8Y3IxGRlWhINXmdAe+YcZCSd6jYdnb/b1rHuIXyHvcd9+rcN2WU/uJvqpT
nOgvZaMQDZlfO4XwmVnICH8W+qdTY5cJ+p+ZkgHLVNggIQGJmeJrCPCDxwHNhrmT
7d8lZmaSpMTaVMr3XkSvZKRfbQAW4s0IpwJ3oE7lNFjElMWrNcFJ2sa4DDaxChBj
HDfcAPlkElrgdFGNZZgGhbv3gGFY14T/NV1eGvFGIHp34byQWtO2nk4m9ygwAgoT
RNexgypQV1slkKby8V2Hw6AfCyASAaHB+UiQcxv3ldpPhqKIQBJrQ/fItnCBjJVd
vplBfqCwfImQqcif0TE/O1dGNVl2nymOa6goONe6QrRCYQcUPVVWOqWArnKBNHEP
t5XiRbvFSzUEPJDrwSuRKOW6EQrp0d0GvB43y2ylhOOrQy6kwB1CcYCDZ5W4L/rn
QYyfOt8JRbiRjGUplh46slSj9L8TAjM87VuIjtnzXtgwFUcKsm9stalAkcdhP6AR
oahulaJN6qOKaPtZN8/KuiRsU8XiaZeoLNw8y9RnJG9BzctMPhoAQlbB+iLPX5lf
QNi3HI8O+Ak2NPDjJTy+w9Ta5KmxGjnfepJ2cCF9u21Y8Pd9OBM2EnbfUcvax/Kx
cEQnNXy5zGgFthaZIjB6g7Y67tPdyVKLripseaMot2HuhtOt0uCZQSP3BUfMYAsA
GQPGseq/gze+JWFvzuAXhS2PmynrZiK4HXCQZspX+DZzTvwKsWLqAbFS9jcUgbPM
aokoO7SsEIwwWYkIkbmjKBDEv8ESs3Ij07hMpjDw+hyl2md1Yu/ZXjHKBftD4ogo
ZQVSUyuqrGLtKEPSTXPV56GC9GccXR20YkrF14E+sO8NDkB2lH+QZ4ndspo1SXvg
iF5g1LaHMJoH/NNvxFyQ6WbED8i46WkXHZWHd1CKC5EGW/RCMiEvpTsItkMX7KF2
vr9fMvuvgSgrD5OLK5eC5XCl6MR9HbXhG+70dMPsbMPsSyUqOMTsG9bkWvDnsAi5
sv6xcTbFdtuJx49SQSRVRsHMdJIYvGHjbz5fYc2Odp1Q7AcOwJ+2Mq1TFlCetetP
5G1ucwMcJ88riAD54y8eCJRTxNP1I3cwmje7l1awBj8d5KHG+CMzN5TpNTCBJdwV
X1OOLMjKCes5fYlz0gsJd7a2z+qSAsWu5WSd1QEoJ4NHWbZ2s6LD8WPGZl999B7N
gRDooaL2U0dLpLJZa9BzVBt9i28rfMXV2JpGcyKlH+rob+rR8+cmHZMTO3oNrqzD
tj1G9CR2aVn1/gBVY3+yWlLkuN6VSEWhQAG28iFJuDHyfRoXNxKjlklQ/n/kZ/kQ
aVZQfwjDMRiKzA0zpArM1ktcUoP73HQjUyohkTasKGW3/QVSUhf0SWFnEQWtg59T
Ba/PJCFe0uxrCQoXSzGBy/JTrjCmbicZz0PreFl613/3BwxKSHyH3LpKFPZqspsN
gJI67ESdR00bhezgp7QepeOe9J6gOYt8HbMcqWvQ9o3AAIvGJAxzHWRDqUbYF3me
LryC8wW+IdKTXVFaAnh/sAJI2NreSyAtQ4eKcW6w/Hcx3jtI4zwYM8ccnoDhZf1j
U8G6b9OZC/JU5eCK38nQYYP5DE/GQXibOuDKFDBxZccgIWBV9QJYHxbFZEf5XhjT
v4vxlcZqX+yAddVV18xAleIbb5W7cmPBM/in7o5j1v4dXpjfEqCEcW3LoPNFIBql
cJO13GpTJ/85ySNOmFS+LS0k9yfJIhZPGDpuRcPoSLVtFKwAIoGNO2sCfgFH8xmt
6T96MOvaN5h9fLiu4+gMjHicUc1UzeVLsT6QnfowSVpYRzGSu9xDhfd84GvXVhRr
0yoSXgqilLVllqRpDxCw3jKDqDef6V5b2DydW+bSSOdKtZp0cH5ziLKBQ2A9YiRF
7pnwMr53UnH4/Uxfb2gD7P59UgGq1jvY8CSPCg/lu00uf+Z9M1VbEfTzeAM/XWaG
E7rV6Okxk3/fBmf/ycHtn8T0GVZ+z1pCj4x7+9V8pELCcxBwl1yS22U8czsCh7Cu
aelJzpp1ghIDl324sVMGjJUom5NcJ25ziyPYwNokRSWPXAO3bdownZ3W7uduFWWN
ZvprI1S7t32BlimhgE2LxUVhJaboiy2cNdoiiNfOKo0bdd1OyHcODjXOff0EKR+t
xUSA371A1kJM61DW+a7bMBjtlh32UcfvTHxyrgsIBXPjNr/4emh0FG8MKm8bR2wI
D/ZnvKp9qxBLvB0jTQ7GSQIs3RygNXmUeqQnwR+TJmnXU5US7IPOWAzecysEcXgr
JxNyRYza/tP3iHKBXCgcCIcvbMUwgRcBx8j0Fsr3DeWG5RvZCqxDIqlictB4Eecv
Reb9OTcqa74LQHxA2ZoVjqvse7j57+AlZmWBCF8IowBejf5kTVU4bT7PwFIq7IK8
lu1NUu0LVGqV/h6tDm68UIOHiHnBcQaBruV+9UtPRH2hzkwq+GmjKjo6mikqa/u5
jF8jvE212GgTIWfGdnJet7Z5YvI1GugIznlWHQ0Q38I8G8l4H6zrrCMZnH1wZwIN
TTNiQlo6zzT1D3s9WxYrpdqkNnTiLHyrN0Wh6ZTA1bK0NTM3C1jRulSwh2WfITJ+
hvczbahYxsmo9ijbB4mHVfyC5sjNFZ8iNTqBibJ/+M9GfAd20vTsLUrGgpB/K4H0
RU/30gKr1q40R1UWkKQZSOJERsbvwkWUqhbV97bviQnsbT3TrdYvujkP6RMwDfa7
1X9rTNUAZgcSEH+owTxyKCCYSL1j1uvU8BgGMJg3+PFbT3AqWMrkeKcmGU9Svb2X
oMnzRKaRQX8fjVq/s1qBodp1j16MfM3MSzmMfJb/cBS5H9g5Xd5pRjU6c6GdwLkm
tZf8tOwag/hP08HEI46f0BxH9piqO8F6E/hiIzZS5kpfPqLMUyN3ccNaHbF19yzW
beWLbsUDRnmdj5FUK2nsGnwIDweO8w5yPuoYt3kcX3lJuQm05i1unlApq5WR6L0s
++TFARhZNVCE0r8+2v1FiQ==
`protect END_PROTECTED
