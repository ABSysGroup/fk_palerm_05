`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
31fAAyvY2sh9nL7Ls4scd1DNS5hoyYbecV8xb9a0/ACKBQw+T3my6c8rl5wRSPUb
owMJCMbYZNyTzKpXvMQS7XoDsZwfs7ntNijVq2kG6kVnpqOthHBRtySUV4qAelNL
zvdBLlwMq5g2pXtt8xkHtXmWZPBgiV/5I27aALS/LUKztX4VL8hVH2o3jKyuFz7w
OXsaVVZYSpkqJ5GGpw4LTziydWOdNmKnB+5JLvh9+GanWT4+XABYsOo3Jk9LdVlm
C9G7RvVh/dV0z/ygrpAdvy6ay/xLqbfpaZLUSM1oSEwrCZJGsza//kuz/N3OdNa4
2SuhEudrV8jw7kpR9MVO1GQ0Z3ZeARHtDyrd/Ou5NmeW/gEwcrQgOWRbajNbInUw
quxZTIe6I4+jOTtq3WtYYYBTkhs0MK+CD5++fAVxyWu2uMeuPLX+4cLlMlhtDNAk
c2ywYMk9hcI7aoICnAlQbz9A1eQTMscCwtokCXYMe3GKV2doduaLkjtt9KTzfeIB
gDF+Mtqg80H0dWt05tE4AvaIAnvBR3ME+TW7qYdngZD4Sb5q/yTt1hYMLNFtCrhQ
NZUvJzYi0Cp3fM3ytT/Jh0y0EsT6LKokC34hcX2vboKF7zErjF0zfJBdt9NBTsJX
lX8H5osDSCN9guXW2i4iBqxi+Fz1k32RVFdPyrzA/RVqkwLVagcTA3SGNtV0dm2k
36MzIHkKRc0Eno9i06osRo8mMz5u/MnkGJDRMWM9YqpkUT/UR0mzc5+8NnsyadRO
HCe4BWt1U1sYDb1Ux9t3ELGkbPI9jnNVvm1IXBaTrPyIFnyYafLweu7pTC82bEV4
S9imnqYOmNVEMY9qVtLu0FJiiC57l8Tldeu86A7e2h+BVwi9Ifgr5sPrnP/top+x
pAtgO16JyFBjfydFIpGqQl1q2yYcufTyZwNDzZVoDLR7HY/Ed/yyg5yhl6mse6CR
Yw7eJoq7w/0UUfhEiKqvFynVaLa2TYxP/t9oKPyP1ZhwaaxWoUzZOlVC6EIiFCQq
+u9JGqxCBWyt6ZzBZI7I4bQjo4SrrAkYwDyswte9ZuJ37ADxyI2mIqOEq5Jipj0v
snGxe4lJ507rywwzhEPuBjvYkIDETALV0pOmhzTjZDLOMFvukI5G+RH4BwI0RA3b
opWb5xowydyjsxW55hU9Og==
`protect END_PROTECTED
