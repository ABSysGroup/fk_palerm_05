`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
brggw+7n7ZY0Ogsqg6LQnvWlwC5EZ4kvAAM4chvp3N1KAnPfC6Dn4ObEsKQPO4Zw
ps1VGJf3or/YDmSgOrDW+3y5eUDOlrLnO4SaSUCz9rlJwBWtjPqACp8VMVsCc2Mw
l7OoWEdop81NMvLuwUZ27mysRUjCdgU3L9P9ZuBPgZ5HSjOg5dOpbo8wczlT+GZV
PYrEu4hTxGAR7ge6UR5MposPui7WsYMJunwoECnHhbAgU3sD37miz0kbZhouf1E5
ynftbkT8sYetCauOX/nxDWQqUAC7PQ9njweRf5BmzZj9Ig/Qin2AB56YM1Tth2GK
xAeKqQ0ES/aeR5WqSM8SxICI/c8U8guTOXyltIQVfSV1GDrKp9Gjup7O3gg8fB2O
vPkRtweHPVQKs6e/pdBl5S3B9EoKjl8EkUpqABrmMwPnX8sKOhv+uD+RkzT/MnOQ
lVmz1+V9paarZy6+Edz7JjsW0Np8d35SIpLGKJHl3zhtD/uH/egBdL9JNbAOeQZv
SJD8xufllkZECHyBxk8ksIfIeBKKOxgVRd9RyJqDzj5mZ2V6RViFZ9JGAQZumjI3
gvBnfQqUapja2bYFRMYyojS7gO2OtIwgaY5QcmijDLEXLlhWfB8ueVYxEBRFbC/3
`protect END_PROTECTED
