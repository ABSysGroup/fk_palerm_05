`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9iB/waijUiXMFDtKzjo47xHdpu87HuYwNZSZwooFiaURPLTp3eF1Q4zYawAKqrM1
3H83os5Ic6ItfGBME9EgiGGIWjlEE5b2sthW2Nh9gLnSEbV9g4IEwJNQkww/B+7c
Ntv0jX1ZUFzeldLbBNsnsPx60H/Q4NfhxE4qwcWGhSRgRep/8SXFdoZ6ZxEj/v6k
4n2+eTbrCiXPYsXEY+xI0Vl4/tUTOQrVjh1pOoszAGS3RO3s0pFo2Sw53+77VvC0
p2T/hrV2IKHjZUeYbUcCehMtMYevIzxDd/nNfeu7JTwc8b1H8BkLQmujkPWAH6n1
hFV6DU/c/vos0wgBRji2/64QBkmrwnSJGjWCrRIfACqJV36dqrZSElXs8ufgC6V0
`protect END_PROTECTED
