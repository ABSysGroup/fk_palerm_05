`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U/0mjewLil+fJhG3fXf9rben+/BvBqBjwx0ElD2xG5MFOafIGuZJ5a6CSfHJrhSl
q3CzlbkleIMikDnxgsQsWjOgLQlKDZzKO+6s9tsdrEo9UMCigHDujo0CfKn3U42L
hp0mXUQOLGQrs0Urs1NZGtelhi6H71OxJoUwkQo+oYzy/gL8gfz68DVz0B5ewlqj
rIu0C+LwKnbvXLrR4ZG1PDTFCBstw3IyCjmvvCrYsaBXM3/NpFfjwvWorpZ0TmzC
uNC9lKjGnqoKTscRDP3l3IKdRr9zgkD+2WYOSEcRo9WzhbxUW68lOXf068Q9MMBB
PZq4BpngvAXGKT3j3AYGL969mKPqKcPdARy/275BuMHioOLA0sHl5URZeBMDT9R2
eWqKd/NBouxL+DHdvSvymBZ4Z1t8TS5QZ6g+pH7+gdW+GYLgfNvr4JyU1ZkMcEOk
DMIQAVdHRF2za5Kn41ApRlOakXhJC5Lb703X9yTNEffLkyDTVUml7Om+Ge+ou1zQ
iQ9YoVkEpIQ4gVa1de1wcErQoYXjIHfFi248GwbEcnULIATSzC+937fvlt87mgWx
ZvqEVYApsbZYNW6MkWxJP/ts5o0DvL8VZIFNKCM7G5Xuh2zg14fKnZJdhgys1GYD
PxSYzIMzPd/gDhqcuEx+0PC+kMqwP1zmgXnHeY2ORSKHoS4UR46GPUK3ErkN3S4v
A3nht5CF46KdmgHP7pe4ApyYOJOqa3TH1All6CFMGN5DssVVHgApWoLZ7dtllKBt
mzwKNr6ILYeRjWqF0FTHC1FonIWuCeZoRH4Bv7md5LCoVrdwOommYBe8GtZcjP78
zMyYtMa+NjmZF5c2YGpzYtfc6yZNSuUv3y2VrfEflWA95Qv03QU83JpZ9/OiItvL
jkex09bFXSD65GbuJgpTRguFIiY+uYHQPuFverb81V+QeMpg9FC80dIQYA1kBYMm
mka/YwbipH0nMGlyXIKq3rduymqrUs0zK1t3kjHsVqWFkTpqxwMiiKLqzgNomUpi
l9lt/0619n3P9DMchKUDDVPpur1zld8I3hOt5ii6gkRBolf7zPQC7OJqOIxzqwYE
+xCGdaMc1nqQEdK1dFErGuN/q+89TLoBp3UxDENVoSvqPEDm/GN3XgW9SfcAAgyQ
gq+IDn03hRpKHEa6p4vhhdtCsk2LB0vN3b+SlUGkmvblHlZQYjXproQiLzFnT+/o
Zm5I6zwTrV9UKXeAh0VdIc37U6dD8hkSlzsxvHjZW74osEQg9NHyBDKMk7Yq05DQ
1XxBS6H8Ig/i0LhHkpOK2JU7HJP84Q68zjOQ1I4FM3Y5HSQ7ule9p1xJ65jkM6yR
gKgPwg47YQMgw+N+g5IRwgeLpDfiEUZU535loxFJyPLUdNkVPz//HZTL6HX0lL7s
dveORzAQDM9Qq2thv2p4j8Moegqa2S0ZzxCQIkJVFOVBCqevzV/nvbw5Z+zL3/yT
+exAwurGOZ2RRBZOY6mbfnbRl9QSpFwyHLvjLnPuYe5HLFjX0ZipOkm1JTthqC3D
AUoTRPp31uVhqmibDd/oEWyyredZTkUGQYuuwuksxcVMlhVCARJXVfHuZXlSXVlk
lOFO1BkxS4wA32Hh8MGuxkYWC3poNxBi1fl9vGENg60C4xq+W8rkZKZtf9WSDJMx
qqCFd6H1dkWlvFGwwOmJAEHh8QG66ZOwY7IsIv5e0bu/fmf5UNBgUESKS33JyTeN
AhVu5NRzE+mD0MmvWUTktYG1zO0P0nA/RAchQW2ZsUuy3XiWTf8WhfbE0zz3LqJ9
sY0K6LDsKbdkIoZKobKMrFPuEYvAcB4rQQ3l2Su2TqmlrrJoilfFDuBSV7V8E2r5
si+BuKt+TPbZR+SGXG2VA5wFVLd2mspErE5LucxuoXzlVJ5NL3YlF2Q2G2yNYN1Y
oENNOVVg9rGwpR+gmEnHzL9aCD8THJQaqQLC/t83eh0+QN0SgdTEpZl9nHyuPSiZ
2Oou/4y2sHVvpacTqA301VVv2aSPtSq4oX+kOmdE/XdZ+zb1yJlbg35UZCEoaMCM
ckQdPPjHCyCFyllX1XO83kniBkf4udiTBdbYpVe9dX9oBtNheNWieQgBt+Dk01W6
lv1Kk1x71T/fgXaRngIuK+ijbEk0/YgKj7P5ViOrjo0t+reF7hzElA0OrqQwaYhf
sHlACTO3LS/5TJ9e9DtdcVfl0+EavoAdCitrWZCwpoEWknkw5EYQ3RgNxKmnrZZO
47vM0QmyT+PKHgs0VkmEdWL14e4Rq8eNf46gGqzRFsmPShcLeFrySVRk1cm55a4v
IYeorvYyhu2vmQZz8neN2RK5OHdPf93GCXS/V8ekp2+nsVru/w1oQr9xH6QBHTuN
+wm08/BmfDX81j+kY5Q78WmFHtVs0MExBD7MlHVm73obJ/qev6Mze3qEaTC0vS5K
GEzzhpN8KE2ZikdMz9uDqTWEtL0JLMviu+s8pltuhS4wFLRp0Is+NOmSXsj+xz+x
klNFjzron8pYWXl+7fxymg==
`protect END_PROTECTED
