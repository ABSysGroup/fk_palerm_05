`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wbHRUnsZ7xagMDIyHEv4f68PKd2EvD7pOWvSnY5+p3LXKjgeIHsGl2GGNGckhKjp
bLFUESf6HICTT/6fq9qiWAjX1JjFCjwIO8TEvXL756nTivtZbzSJvG6RifRYN7BY
RnldWhhYElm2/IRaYr+3wDuG8NUagJe2Wsuzk6UZlvG1saBmg55QG37N4k3fwTbb
j60hRSQ0mZVFKTaVEUNIir3IXpMZ1sRYMlKAo55JZNgjGkKJCGkBKah6rUcgleIE
hY3xdJNvYJHj3XYfetXFKoV5ILVZbzqodky8OCMAndkyudUYKmcoeQoNe7LwJT3K
`protect END_PROTECTED
