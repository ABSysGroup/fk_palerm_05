`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2AqsEnM5rHrufF5JQ2byPIpU7FzOweg2ZU3eS732HorJmECQ2DNtGp3wMDpimaRT
OWQsQC3xFGcXmcr8jH5bOwkHZnRoc5gIma/3uR1tA+w1BbCWgj3iRyein82Bap5w
0NNRi3s0b+wHTzGJc9JojWzHW2raRRj+2nxpR2CB6wXvqRj5RWcEaDP+HKkv8BgO
9KgPloSWpM9k2yFrXAnKpOXMmEi8kP4QfzJ7FlAELls5zp48rFajhFIZvhb1isXi
xlCAQ7t4PveoSkybzgyA8PUGVHJ2JLWfhaXxulB1ZaEsu7o9/UcC61+ryXZdgnZI
M6IjqS8kuRt9TqkDo/L9hw==
`protect END_PROTECTED
