`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RNF8drlyzLBwC054WA28ohgqbeViU9uCH5JpnNxGo137yKuunGTkaUvsPhyzajsU
0KOIRXQT6u6q098ZtwBFxPc2EPTb9oQ2farOVAn6RET0cu4m3lvpq3I0SeY+nUI6
jNNhS9H1yrbdZAgCVB+qyKcRrDL8QA1wYOToYEzWUa8DMIr1iHiWTPiGAsX3nsL1
0GY5++BdUg+NDEpTWt2Dy2L+1JFIjOw/qrHJvH+rJjFu+Ltr4hSx3l+8t3EB0duq
z05klL9TXyqrxO21S5eOS174wXu8tEOFc+j+0KuNpXgTjhhQbmbC03ndzG+C3EeF
iSQvMDLqPiM7MH3O2QVaXWI50f2hkQhxhVlZJpBSgQzEWp9K3wlFkxr8cMbXX2kz
NzEQmUFT9SsDCfvD5WEdRyLatpBFSp93luCRYtYXQ+8A+lMYR3XhmFK3vLG8UxKi
AsXYU3qXkpWVu0bugf+RNs+nAdyrKrWNRf0hMnRwxKtOKv3/0Bv8TZVJgjLkLPT5
rDgoBsahJA2udyJZp7mIswHYs5PpSvGXm5I+Zd9aMIs0oYg0ONtGYee0PYN6zW3k
QZ9tsJQA+kw7pAUE+zgdhhjNXtMK5KE9MCIVVBLVjXx8Soy7I21ZYTvqeKPKXWSI
Xc5Y0MChLtoIeb0s3MjAz58UJ5yGBTRSqutNdL9ndm/fwnT9ZXi2D2ydWw2M/n4B
bdD40UnxQ6U0PE314tzriknDxtVZTYj/dLro5CtZ8XGrELGad10rZjX2kWG8Zllw
l6Atg4d0IjyYEsItgnJgEcsOjNxh7tBBbNMVJpnFm13oeIE65ZJDH3M2+KTUKAm2
XC4o6oYB4UlBvI2pgTxz8NmWn3g60bEAI9cMojegopWTqhUJIGTZfJHUs/m16Zi9
`protect END_PROTECTED
