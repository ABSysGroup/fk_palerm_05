`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BDMeKo+t5zkWHtPsHxmsiSSmZ1fCyCloBdz4YgI5gHoY2egZh0MhWNFAL622Ua6o
fEsnfB1risJgoeqeyuvzDnqWuq0l6WIbILysfAXS/WFsT90WVBtt1bgprsmvJI1J
P7WSCrN8q+91w2uEr97Ni5Kv8uFUNEnvYEUiT4sHIft3ig9t20KDRPKNhohYghvq
hAHVGjHiq2q2IWAZf/EX6cNAOVF0SVxmZ9Tgs1GNqMjL/B022aiXqMJ9HWCNd4iy
tMhlCsvyrkx7Xk+zJOx2D9E1hlJ7eApkgC0pEeiGzXZgNhg1JzNB03mCPrxDSl2h
yD9ygfCYhvK4ZcDpDBtygm0+4HRKLuPk6JqJzLi85nBdHJRqazXAqrwW4JdLscO9
apH310K3sVYdx7JsxafWjg1ZGgUrQUnNuJzDBGrMfl+Uif3peW+hi7Iue/aJRq5P
jin3GWnDfWZpQ5Onb+DUpqWQkZv8N8u+aDaehUHH/aukY71PqPF3yOzNjX6B48by
WlrDD3dv2whPOeVPVln9OKobRJPtbDpsKRgoTVrnoqW6DAtYGh00aIZJmxnZU4tF
HDHPhnV4bQZnL3wT71PHoqUZkZCbHvS8NiS0Ud3BM3syn54rBF2eBy8lkcL/XdOG
0jFuT3Yiduws1wVs7NJUkwffQ72W+6Vgp5pBCp0qOqTYb9gANa/ijl7kiQALoARp
XWBDwIX+KzZkNn7jdIt5TQ==
`protect END_PROTECTED
