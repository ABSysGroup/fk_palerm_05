`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lJMvdlh4yfwqii8EZTNAghtA1WCNDlodv/Z51EmjlC9tahpDy3gU0W70MaLgrRrF
LMfrkjHPSCvPW5UyTWPdC3DkwSL+0kItMl3DBcmjn2Dvlkw77YmbIbHWjentbbh6
jbUgaQ3cVvtxUGOf8icOJdjjMa921hW/ehlNkAkLPJ7Q0LYR9D4qEraC760HdcLQ
KguyipFbhE4ozHUFFVS49nLUgPfKP5ScyToU3zTIdDS4WdRpNlPfI3dia5TH89r1
5n5LKJjpbC6MZiJ9J2FTC3tDUoZhDVLZ1gXJ8ZziTo9blbOBPBF58NrtZKVLG2kT
seUtlD3vCOhpeEPHZa1POGF/OIEQPJSm4w1S5fEULavM7lpdTwgKnV3JGaR+sNul
d1eTlRnPM7BksgSAmth9aQiRr+XukgtB3cTfizw7IqvBVl+J+8OI7QP1MWoYuBbe
g1oohkdTa6mEiRs8V4k7HB4fN8PVZAIwRtLYkGgEWOu0cqtoUbaVENzJh0mE9L3x
/Jlj6W1PVoE7ki7bQ65h+oHuuMNVZ7x7WRmpMZ0Lxec=
`protect END_PROTECTED
