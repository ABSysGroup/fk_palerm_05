`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v4mGr+LIb0vw1mCby3bR7/uL5NEWiLIW7GdkkppIurC972NbEUFAav125WnDitlf
UORS8JkVB3xWr+4oZoNoG0WXbVtf9I2Iu6yEUdy/b7z6pUSv9Yonlv+cmFBLH+vd
NYTVrx2HjR4bQX2tZYGu5uH1zmkmSP7YA1vZYPMQMoY9kgOeq8a+88m03ugZDX2F
LP5ru3Wpjaew42Nk6ChOYNhKbfKMLWwkOhj0QVimvw+6sP1mJMfqHwvTOd4MDygb
PSDR2hVG9BL14n6HdYYOnfM0g/iE1pCdHp23vJrij25g+rAXrGJV35XrLwHbAz78
FuYp+iXVKTQnBYnSKnI9Y4dL0zGHI0h/K8AD+3eyEP/hEuVbZxzdm1MyaypVlFfs
X9DkrAdpLQP+y5AWvtNcrkvxA3Lp3DJF4yIjSzkbjDeJdHee+4NCPLT5xiyvcSPw
r6q0b38RszAHfx9upwxxrncq+GN5ZcM+HZb3Rmd8xm3Yv6wldYjB4fXNF/DC9kpA
gYkNEFV2BQH0aQxb/zXXVmCnk61xGMO4eNF7O5iO3XoXr4CFFporsKGNjLmxbFmT
kbVLpa86jmDzgXxVSN/86nDcslmyAlFYm0+SYeZ/QJLeznq6W8eE89/UZ0C5KMAV
aWhUqOqnldqt6qx2QlqwyyiHKo+kyfDAiEYHgaTGjj2E8/Y+4Q4PoWH9xLXRGYE4
bWwG1+eEfmmhupFR3JQq/Qob8tZymF7SBoqany2yiBr7JnbIk0HzR2b02Zuze9gG
XK1MNuSUCzNBk3WomCjj5CI2sM7fPxVSsdLt5+tL6qhGCo3KAX3S4c6rbs7A1Tll
r2mGmFeaUtDPxD4DdaHmQs5QywxjS+rb8qN0AD5X1YVjripOIXkdIh9gZ5kSCQxu
dFcALfEtcW8ofs+wRYfG+bucw545D2BKpXZ5Utxj6YnFwT8KM+D96nZ4g1y7LyuA
`protect END_PROTECTED
