`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zCYisNDaZEaxZt4quP85+eHnIm+pC0gpF2FLR4MDHSDfuk57oxv3EOCAqa14d5Rp
lEzaAlb1xz1DPkDTtdfoPKBB3t79Oc4Qi6XSOGmMQHy7mM9LBtXa5Kkmr4aYQ1pJ
7gmx0A+Ycig+4oTh7xSZgAGiAxgT6qgsCYfOMHr4cLgwWJiDkdrR7bPizohZpgaR
qYsqRZ5Co4r6bc80OuQPZ9hPe1/rjDwLyzI/EnH6wK3vEN1xKDbU6jVWeigTTqG8
c7Sdg5ddTaNMV9ZJKkLIcFk2jPuP2aV0QiSCzTUURPMJsoSoV3PxJbvmjMb+S6vH
0cs6/t7XlJ+M9fpT5AE3hVDN/vXzoxHQPCGGMHm3CYeit3GAB0A1xCO6yKSnrT1K
`protect END_PROTECTED
