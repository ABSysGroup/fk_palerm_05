`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H2ZuLdU/h8dJa/V9sQUcFjcylVhfhiI3xEs4mrjII2VCAGilsF97VrLzsJo/iZ49
L5nT5oqVUnYiAhFDhoLuDgu7nMZIMaroBG63NLO6IpwOinJ+qHDbYFkVcUUsFJ8o
zvudIhz03K1RrfVPgpNQSYaPDa1IdAmmOY4FfSBL3R8frGM98HekzpALruLw7Tgf
nGZM3LzDZ0o5eJc0ZSJvYX/3FHMi5wpQoxglJbQ8U/eYa8xBYaaWAEJ6EVFzpAsF
iZ82IqKAtPLpZPH2AfCFwgYhs2/EZvJfRSoiOsmSgZL5+mtB0EPtdHGCCcUaoton
+c6LEqQCo7uDVq61BWFDgJDY1tXnIAQ/et/4eTn+dUWKyMFlwiVF3OZ5LLQv+FLI
3Y50r0V+XxxC+yj3uXXcydf+wfB/L8hLOifZeMu45zDQ3l/dpKA5mMphuzXaPuHi
jkHF/8IJMJ/AEL0mrFVzxUWWrB7GEjN0HuBEraQwTs+KP/aQQM2/5UHcSZPUoVkj
kgvR+lTDQ+2uUN8/X//f8xs9pf5BLHyWNCveJ8hRwKOChj2QojTN/11dyY3Fr1Ld
1ucR5IrTayZhzVquWFpLYGMm/yaEvkjA0M6Uc7SDPxmEyL6fY/6Jl4HYtZysLNLj
EVsOuz7aMaj0yXJx29oho3Uz/ABGd+1DOTD9NDF6dYrrRambK5d+HWacSp6UblO2
LCNDHe7z9EAT+jiVahP/YqmmDImaujm02sdVlBPRe5cku9Hs2ni6lT47aoUhb4tx
Fys99ZSFsckIgUpFomqyFg==
`protect END_PROTECTED
