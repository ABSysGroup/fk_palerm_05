`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C1McIclqgf1QmiGStVxmrN0FZCWRSDE4ZjgI1eSFNCJ+GRxovF5rBqK2SxFVyVbv
2xLawDU0xdFXHPQEuLlBDjtT8U8nPaYlhZ7Xf42SKmEOI79iAa7d/4YApp0/k/3O
VI7QGbej8K1zGbKgz1B5DHwiIV2Tu1lYLuu0lwE3/GSMRRP0LzHcc54Ro2DNsHfV
X5ZuvoapaMzHx5s2e8JgkYZYME8VmWp5B/j44/8i7ic8uCM7URrevFNutgl9VxJ7
c7LxYvCTKTgh1jyY8a9dUcRT9ZnyiiFNHMcOAvAoyLUju4RdPBK6ba4A9X3LkaFz
DoyU7x0EisSyk/CmhvTbwQK5CIm8hls6Kmb9xt90cxWT2F8TWMz+n7OViHLEhhNQ
QYSAK94iY2cNyM+xeFT1C8kTMh+yjQErfjk/xezP5FXZPNTvA0Q31AR/xAsMbqMK
vp2rTkQB2ecb2+9/CkM0are7U6uaJz+2X01Iv35Q6VVKnnntZGZHLrPkv3Q3JFEk
xKExw/mC5g3D6JMg9s8QpPgO9UkEmezuCTylmnWiBXSJFUXO4UjDleR685axv7gM
BvohyuRJPHpdT/8gNshp7cby+rFAT7fwwTMp5pRW7xzUx0HWyesH2Eyn8FEqa4Uc
R+b8RzB0Zjak9zUsCaTtkjX6QVjfrfh3lEDlI3Nswg4wHp5zBl+IaY2SlaUzz9AX
LopsqpGcZy3nSlD3MaHEQkePZiFRQ4EPYSHP4O3QI4I1bVcxOdKYCU2R4RQp9k+8
8rH1vGO2XPGxTzjLeqffmas6Kbga7iibEdKxC/MC5UfLFoyKPkbF5LX2YUHzSXJA
wEm5oewzZ7ID+N/3f7yb8iqIdfSYVdRvin8R2oNAC+uC+jqVxCRfCRbWJmUDXYSg
ww1rRAsZTcZEjOaMFvHWIxEdZaAGWWYLQp6ZeR7Qw9XLuR6YThzSE0Cbpxm8IL2f
`protect END_PROTECTED
