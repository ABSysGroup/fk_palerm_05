`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
09NPLt0jZ7/tgedJgyAD83r5M6pwhQXWLzdeY1VHuPL3vU+v226+g3MJxeD6so4x
cWO32yd6yJQrLNSxjW2632m94cz7rIb1eOPa0hIptayr+wmNkR/gITlLpnZIswyZ
UxpzBrMYYArLp5G7xsYanYBI+VazjmIVoE2HwR85/a1D2SXmzfui207FSZEPFlmO
/N+J7AsE0mwLTEINHGQlaRzd6DVTWwX4NKR0p2+tKFY8ZgVs/WNocep7zkX/NeCh
MwXC2yGhYNzE1vwO2Md6uBcKPgWxrRmSeCJp1OghwrtQ0rgzwIyQkDlfDHjSzPla
BVNvwLQhezh2LnDM6Wf4twV6WdtbZiYQy0u6O9udKvmRhbxxyegiPO5rc7bF8P0j
jLYybAKe/ixMrTDybHB5FKFJ+cSbsTOGGP/FUnFd6FvS4lJ5AE3ILo3QtCs4AGR9
PGPHTN835n4eanVXFLH/TIaqDnoYLbA5Slnkfp8Riu1QWNLAZU8G87x40YSO+Qyy
Dng9kIrcSvqLs93u7Ilzg2tQHaNleXhRNyaeCXRbeAPBsvOaPFwuUX3aohJ8avw7
e2yy3L09LedDWONxJqIUX3KsinVHK8VSHosanutQFvU+12KebSW/7O7aoD6kyWDz
VYSwLXyk9WgSYjrbC5KrB1dYNFlZmPW5gGeDZjdx/BtSTXleh/aWFStzSB8Z7vYt
xv3UIluCQra9CbcJwXCkWhILPN70dVpI0hooStc5+Yhb+Q3FUGlX4IMbmZUkxd5t
PdILk+pe1cqM+eyLQ5A8OkGzVcOIu5NvQX8giDZkOZh5xg026tvtpqOHxR/i9hZ8
1P0+VMhgvSbnJkwf2XHCGms0YrJk0Cg+6PZ8YNcj4nCqPvPmXE9eUjHI5kIxcXlK
nFH9Rc4Gczz45LxbvGqzhsui/RMVj0U5q0s9W0SAzKIJ7vuvrRRSckbZV8/+dG7O
5hJj1LbXlMRZ9qB7d0o3gv3dyCfcqWDGMCNjeJo2eey8V63eWwOlehn6xOF3Hqae
aXk9t6XOoabRvUsv8Gty3kw1TiXSG4PSL6ogJTza3/fUzu4Is446CwsSK8RZF+Vi
4QlQ5ZmJtj58rRsXl7E15TCE56Lbtlz19exPLGuNK9jWMKQn/r5MPEaL7Qp/uNCX
g3Jeh6guPJ2StBUvavJDejDc9XqfXiVrswi/3LjbFxX8mSmlKfosuT67RewAMBFU
xNs/SMzGqgmyxlDFfnazsqaXCSR60M/nfg5zCh3qeX2sqddiSWQns9GqYq1gFnic
pw6E4PYeoft910qBv+xv7ocNeEwB0c+8zgCp1V2M4sw6yJ0uSVp64t5tPMggdH+o
3VqA08gFFOUSLrr8+nR7WaX0NtMRhbNBzgpA5hi6lN0pUl2eQlHrzhJYFBppUMRf
IM0zdvWqMl5M6mujaVKSVXTzUDpQVgVXGMzPgDD9h7s34DmOxHi0wopdX4VZPdaN
DXIQhqKs6Oy52OxVfelenxVX9p3PBU+jGANw95FsixGNWgYltnYwGJcCZUeFH1zA
VM+PJE7H7s1LY+pG4Hw1kHeWxpN7r0pvREjdKI2m961UgHmGP1ihAUby7Wkfiss5
jVbo+mAaQ2maGZy/qIrVRWcRjNwSV+bDTnIIIST4Kq14oryV5ECYwLIUdM0QDB4D
3MH1nDT9xxenQKixBhlJxnq+XPeeraX147NQZsoPmwiJitRVLZJceZ2JYd7WoADP
aiKOQyEbb9pu0OIvRJe2dIyKnOoLs2x9NzXisU8edABPlTaVxXT3CwWfPHL+de40
Yg/TLlL3x4atfZELzc3lUJ8yhqKRbjDxT8iMVG4pYEVASi2dBnf03s+FqwUmsXJ8
`protect END_PROTECTED
