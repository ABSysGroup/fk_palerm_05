`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eJZIkvbtpihX4WyTdrjtwbILMkx/pdbW2Yo+K3BzApMNXeAT30YoHI+feyHbnwdC
SUnUmugsNcAa+qnwFQt+QXgkR/stYcVtqP6HjINkvVBYTVUmt5g+ZpWvjaxsKpt2
16Wfxtvd0CIIVcjjzlNTF+mws1v849RRvBa4GxmcZbNhl6IpQOB9EsixK5i/1Xqd
F7ez1uU6xt2tBP80bk1GTzXIkO2df2IiCmgBBDU1Y8KPSPuUKQbrMzvdlSiGB2RT
/alfA7fczYbHYz/CcrO9VEZB2l03Rtnwj/c4jtdPBg4=
`protect END_PROTECTED
