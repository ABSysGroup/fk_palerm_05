`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Il7mZpBNXLnpt15PPD0rpq9muByP3XOF4w/xlxQ0FLfZIFp7ckZ92isCgtXt3nXO
osGkSqPxZt2cOMBGFKhmAQoXLtSYS7e+g/xotG6loJfOqggsetgZ+3Ne034wdZ2m
XWxWsKbWMe3yB0kW8RAo7O+EY0I7U4w4HeKtG07oHzO5aI1GWmf+0pjKGCyshlXV
YBgceqyNUTV9jBEehapU01InAbXkXV3oaGwoMHnDty61FKlWxkCGqlqrJ+jaQno/
2B5veY5ol4LUalVRBQcQHMoAdIwDk8nQs1l1kdjdUkvBiFYHkkQuu6Y0OhwaGVIZ
H7wuhZe5HkIsZXOSTu89y+55m3B9NmYYXz1eCMKTkfQyUhQXWYe0mNVfzkLpRG5t
xpdWwf5zDrwLmBd+r87Npg+PyXj+6YMXD8zHOk8elULJD4Y1GKwroRRHA8XumSAP
wgIecX1RTDs+JMiPfVS+mYJWF8YWnajxQhXsFddMMZGtY2fXlQPFGgNOmyJS2miU
DkwebL80tzewNAsC23sbplak+94ors8ag1vSMLZtiOFzXnhxk6GlPYhw8tiFPDNE
2sX6RFoupPIDZ2RHlb9TR9Lz2KaMDhX2Ckrdl2fDWLHrk4dh0iTcEkD/AzXV/MQl
i6JY7xF8xBULgGP6LEcpAbX1JAk/PoHYKLcWDJqv1z67LZJuKxdPjcJNCjyw7RqA
iFOoByYOVWbaAhyvmtoaryMCUoi47oQ9VPs4kAzwh4SzqLHQLjocLVmZoYNlaOPI
G+gJHwi4bgoGt+oyyiGg8IEd4qeMeCfYdbdzKWsofR4XboHq49k/f+NaNY55acFt
4Q9p8nYmg0zsMppd1qcw9A==
`protect END_PROTECTED
