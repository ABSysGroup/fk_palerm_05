`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y2QcF+3UXwTp51MHYCrAIVP2HFeOMrIxGXYHn/7tMMzZ28cBH9SDExkTb7ftAjO7
B3T3Gn4G/ENGMsFXBLwX8o0j5MzZW5TPikyKqsbtAY4UqQf1dVPxHGrgxqeHwA6Z
Ak33DgtY8DdLWQMQ0ybf9jdQPq7rR2AxpmGDR439ZZVIiA5WbF2wwVj3qLsgo325
bPVU8Qy76R41FkoK88mxqEA9xDr6DBeJp4mP3gdBny2vKxkzNLDY0t5YD5n6ZHqk
wRmYX1Wh9KK8B1wI7R27ATmLn6XJS1zFuA03T7+IPOEOZygF4dzTqnydxf6FuqWt
F80AG5WfK7BjzPMKu33MHgesDGXXfEkHp/99ug+2u4BXoCjqezXn5Ilah48IJk0D
G/DmXPpKo7NedlUlTHL1p0sSOAL5O/kRlnUAbsWy2jlaBUjhOfUEdQZidg4k/trh
k1Ph7u4xtrhP+E4C7B1SPO9aNUCRT5s1RzfdBvHYLvs+3u0Kk4zGqmYSFYLCgcvL
VwLwbZDsBkQOCH+HGTp9RmbrWNW788WhCru4B2RE3CMJb+pcj+m5ztcHxAI5zeLc
gQhdq5w2KQ6xO6hF1kXtat8ApTH/jrUNo0MRNuJxsQ4=
`protect END_PROTECTED
