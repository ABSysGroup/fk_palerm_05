`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
17cojcHkJQXBoU7pUsYCUZM70rAon/L5CcGjccQbZFpgDWpoqKS6IHOus7JuqmLD
esVnS7vQ7vDLQRuOYnjfi85+8Yw3eNV7wA+Q2Eo4b7mdIVU/GXoqtfQf8ME4jEet
e7llAR6dsA0O5hxhpaN/4tLhdzZMIknPYndp15P/1Qf2Dd9/ECLt3v+JKcWPObZE
VsuvPL9LH4IaZil+M9nnacJSE+RPjuPVTuXw3wZzeNyRFoTrUsUcRmHpB8Zhbfud
F9LnypCbvXEWMCK+V3n7ZRrkh63hYKIoPkQKSh1xkur5DAX0bdiIPLSNP7S0orBz
bZEwYviBQfYFGvhy33ZXpzH+akAubTyBscUP58vXp60rL7233KhGe2L0vKGHFiOb
D04JAoD00IL8rXE6fu2FPq5ifc/S2Eb7iN/lf+qwLdsEmPBpByztvnqN6XjLXFai
shldSuhrX7IUVHjgw3XSVaquX09M+TQDNKgvKDKIvjblZhdR3mev9yoLjr/NtZXV
r30yq3pFvKD8TklGK7MDU2JN2o8/QQL2MJDo50kfPSoNmiqzaqvrqHE0aGjck8wc
+tIm8Rj8QSUGQSupdHmSS37kRsGx7sgfjhbk0BqH/rXpJUkMUFxmqEFsWxyRY4vl
EqWsI21cgUbrys57rtLxI95pAdJ7C232KJdF8hkjeKLLDF8jw+JwqBaaaDoS638t
UgbNTJWgwabBDK87V4YrBHFBWYKuYev2U8IHRRTlRL1MM4Mcb41baSHkt2ZKF3FN
343RHt2a6FwOBsiD+FibuuCgzXTMokjaSgjKPJ8zLCcD4Zq2nuG4UXHhDFT4byX5
zxYNMaPDie29wrCSeeTmx9CmVSGVxCrVooBEvG0zEyNZ/B/AmMuT+1IepgHZy8BO
Gsj4T3cPFgPRaXuZ+IBPvzyaVy0K+tut49rI1Owh6aH2oLBNHmbJHObgmbCqW+eE
JTVhpam6+TYEctwb9twrw4dDhfCauiuUsl6G6R4kkkPJny7vaOL9fghGR5zqiCgd
KZHf7OnCH/+KXwDbhzGPKcdjwJ46STXDdwjIZ5dWIwOk+Sj69426erLf2UNALEyn
kiYvAXLdlSevJ5c71rDPEr35Ep2T1W7Pa9TyCknhWqlSj/CSctxUG8jU/tvidXTf
wBSlpFRD/2h7XBdvZsUXnuvvdz4mZRJHlXXBZyAeQclGor5sJ59Wfy+sLp5pjZlJ
fkIPgLaGBOC56t+90Jp9gS6+4PbZCzEQARoxX0z5dAHav/9ye3Kr1p6ohY8/Ebub
xd+lBRGsTr1uzg268ZbViD5iD8oGUM9uqM/gh1hqfpfUCOIdpaNdCBLS0xj5Z1in
1KHEexLHfiwj+0y0S+62hbmg4F25+AZz9ZeCegmxmd2IYtgZa1Lzrxd+SWyeZTHu
4oEykSIm2bI5EKwx4bJcmCd5L/ozWGgkFdXwglUjcp94GN8gUX1tasl5l5fgVIwq
146B8OJuTAy8lONrnH0IwT8Q0veoEd80Raw01xeRzLn4KzApEgeH9Ddas6tk4cE6
x5S3JbL+8vr1Ba2P0ASazcAUPQmYVDUVVB08Av6IvIdP0QDaxfVeUp+pyXgOpmwE
GU5rYy03y2F1epRzlu/EOiOSh0T0V4tUr+89iu2nWHW8vCwpOtp4trE+mo2PHPxM
47B+AcAsKdC8EJSGkyzuLlR8sOkVlt1sDMyXBhQwRCg5QwYX/K9sWCnAVB6KuQ66
/ZirO4UOA26GFERtvyESWEMFzXABbt3ZNcYJRR44jEMnlMg3S6lzzMf+cG6eXfBJ
RWZYBu8Rbx92fyGlTze+xvuInlw9/tDeKw+R6E3DhSNGQiml3U+WK1frRZafLkFv
UeJVRw2oidB5urOVyTpPveybyMFs6ZmJqgqiYiZLHGsdtH9ynITK8zN2oHKg8Fwd
0yxt/sZxYRjmZmOkciCJ9CsA3e/3y5YGyZggABz36dlMMQZvL+/fnWScGu11Ycmj
jXC3sU+oJh83DSRH/PuT1s6DdmL8gjmOeWw3rFcNIesQEjZZpLpADlU5Hc5nuTpb
LRCIV/DvVVQVbM0Q+TTG/m0wTWmV5OpCKAnUlTq4a1B1jKHwnnddI6ld1zZL+s9f
KYqdyJJTNJg9gweRMWhZqPiLAB6SHE0LwNuqXMqRw22/A33NorNpU2CFM9/Idh6n
MT6cvo5Ohgnz7HJuLXBS01s7svvKsiNI6+gWuZBRxwMk0xwtEDC5+7zmSKILkAkh
i6QUq9z5J8NY/bEcxT+Sq2Ece0VC3hsL/VG3zzx58HaBtNaI1BxEQ/X6WhSVxo+o
43IWe/TXiFntZndIie00DGNvPc/FI4gErT3Z8yeZ44vUNWmJK2/9wqj/QeQzRDTR
3P1sViYFHLbE7xaB1RKGPdt3WjwZ7zAZ8iJzJhtR6KA=
`protect END_PROTECTED
