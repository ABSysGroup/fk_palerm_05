`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HP7Cj/YaCOWItllOk1an48KXRqgCaU55IxYXEyGZeq9VgcWlgJz6BUKuMgwEYzr3
j1tapctaFqj2KCCErSyGWueZCAGL35yZLJdQzC7N3dKzF2DmDJavzGhsR57or+Ka
oxEyvv9AIvOQ9iYMi7IiGhUJuGlBCSrsukGs0mPwsFjEXamqxndtKDgtJjqVrrCY
Uq06LyzizlnEn96LzUrXyHe5YSpUlyzPZXEZOClAxHhfd0QHqfX4dTEsnJHSn8Wp
B+WqfGSL33+GHyysgU74gixY3iDTGtMTKc1u0fAXln3rVPDFV0i8e1QEwTdK9jY9
z/pLU6Bp9TZHtTgWj9NDqk7QZzq0J7FEvcw+XfWG6N39Nia2E0YsDAJaMoMUAbFo
JUwq+lNNArikz9Y58BpLm16vJhr548ncRkJajdGMa1JuxC9GX75gV+7xEa7UwE26
lO1kbIkoluu616+LrNyD+lR9Ro2TIQ29u+Pdw4Az6Hf+3KwJejlNvHN6lPK7+HiB
YuFZDpdQXXlVgN2NpMd9suU9tjSnBmqlihqzIBA/iwH806868EluQeoGH/4aM1C6
BXb1fk0t1fKPo1v3kfUYC4haVgC0aGqHk93h4jcRxNJdRDPRNq2VAg2nkpqnv+TJ
/sD401IbVU0JUQltb4XMCopvv+3486eO+zIXFxTVGyZRJ8IAUUDUbslFhx7ad8yz
xjlBxewqMdf9ZIgsiflXlQEzeRhkmoFsi42amBM7X8o=
`protect END_PROTECTED
