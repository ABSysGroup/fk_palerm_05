`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pZ9m2C7hWlwOGsKtuB9NVxuhMrtaEEY/VhWEgnA1T6wvqmE+jvAou4grDYt9gScr
bzglKv9TWlRV2VoljdO0ucTm07uk0zcdDSBQqC05lG6E+d890u7P68CcNQUkw9o/
jvi31rC8atyH9IlWJbxc/BNdm4EQhEFeHWqHdqfxXXJzIrHNEpCMPlwYW+BhFWM8
z77JrNc+u0btV17rhdStoGCpeFO1B8C7Eg7nh9RdLZRBE8klSj7OSwxgiqjYUncw
HYVZ91AmkJyru7wm/s8VnJ9ItH5+1vfRn87TuseF1GBoecTKFDIglxDho3k0n9SI
2OzUp8X7yVV/2iHOHIbOXD94j+3s+JexxdPy/gJm+GJD+RRiREa/roeabnA4Da+0
EygbloibPl5mHHeflvwtG4anC+hragi8sfzMbNdh0rZVSVSyhWLftiHMieDHn5X5
8FVRNEGRJjJysIV/bDfXWHTZS/u+2u+9ae/U/q6sf5xiHCTNo8uyH9WeqU1GrdWX
D0NFHqrIQdxDJty7167W9hfbKOYOQF8R9F9850MJFspSRzdeI0SEEG+v0rtvJl4Y
bAYKpCcw48sVLrlzlZHdRNLrFHjsPKdsPIf9opM+hFrIn4PYY7+tqav3AzDP6JNm
5nAOVMjJpoJzcf++D0/RIIjQT3qOgrDPnUgjKbNNzmr6vCvJYesCIiTwOdpsQ+8n
mrnAoXHHyFPOca56cUh9tMLZr2oThGAGnI7rgeJQ0f+uFz7xBu4on+lkigsTf/kq
MZWYVTVRHWx0moChrbVIzwGS/drNaWZdiAzCLwLlObxa7Qxtw8LwwxVDiutX7iZM
p/w5U/OxEhWbCkhR+naPk8qE/wJExz+2ElIoeazlXXASFEIjeLk4W7DhwOTDa9Mk
oRQqveq4kxByUIyok+hYSbT4QW6wVwBzIsborJVqrYr3ULs2XrFURPV7XT6PcZgX
gv47ulycXBnRTrPuGVgWGQZKdow8kelgd7BBnaEm+07lwmEovtutp6nG9ukwtY2c
PLhwYLp1DvxWYteJhSMqw7E44KcCHjhKkHEvy8eN7/CvEfLGYiCVCMZ2y80tZLd2
HMfiopROUBIRDBr3LUjObxC06wmWuEDnaNGr+9zd0RtYLySlLkrAUo7SbMFkq9yg
SJtt76dmojrQSJ4uq0ftIHvK35yMPsw+741hTBoJ0Rbco4Z3qWVWoLK2isG0OBub
vNlw7FY9Cz8w3qTdbyOhWwo3ZzENPfrzKoVXWsqZwsjVJ4R006Ivc/BpKokdQOyW
BmbxulqR0BRHy8zwWC+/K7b+FXUSL0nrjaVd0OLazAF8CBa/MP/ozqlP3FZ3QS0y
VW6Iq3BQb2UTJ7GLUUzuxrmJ9kaa1JmZB1DRzS+spM2ntDv9SI1NDyBHYuhhhkKB
bZYmagTqVhDrnTeM7fwbIcvD6JD/BIMz0ZM0R9OWX+swl/TYbr29fCNRphUxzgLU
nKCl9bR1Mmh4hDaySNFnNepr/pbVML7eiAdr3RkN0OwztbUiPnEVZpIH+syeD9LN
IM1GPCwkCRlnV+jf9Xnr0PXDmdT/wmigl7QnbbeoCCOIfrRWCNszYI/yMlCJbXx8
NWA03D1SnVmuQmkwFw60TrN0m49BASwQzA/taUeXyvQ3hrL6VDuX86mowYB+63vs
m6LsXnCT9THI0v/yKAi1ay9ht5kgk+Dm2vSRXJLG0YZbcCHGIVbCoPT+6vIxPC64
UJ3C0GBeUh1fmetZ1476laO3Lp3qg0tSk0CYbkTbrgyyC8eK0IipfnBzCVpiNf3W
9X43Bq6lw/uv0dO+RSpzFAYLPnlMHvG/hw+jU+lF4Vp913BahDSzq4M70VHsKGzk
bB0GrThkVWBh9UTIvw3errHB44lC8umGn0kX3zw2FGLNKhWlhFYzR8RejiGVxzzM
O1bDqSdQT6tVjGJt8j0m0j6V1s7d2YsPFE1NpUjItj0IRvRI8zcDR5JG0T/MmCei
r02mj/0K9jb6R0HknPcZNp0vtFH/CYFsfWRqTdsBCkEQvct0lPtGe+8TovEoR2tn
dYXbcwk6PzDP0tNMMeastXydOVvwrXUBEIhoc7me/Rwpif40CvY+F1o6BflwW3rV
3Wvy9AIQqOwhJEJswyWtFJWV6rVqy+YlEB0mwua5FO3sbdSO0fbPxFt3YacpLnNm
Yfh/YkKEUrhqVylcuMjlIwtOqphDXBzHcMu0w/nIWNCVLCwbFOtc9ZYx4B2hkBXd
ihFspDApXD6ip610gIYTdq0qhY3LoIUt5f4mbQcsfTYqKMdlASR9Rq41ekpuoo3F
jZd1HnKXnnqCcDIwHQyzHuGBgeuuvLhPluywDH9YB0C+CF7F5v9Jb+klarjBOFnT
Aq0Q4QGXKSs+x/Ry/8ixfqQtq5Toi5sFrzV6e1lSytHm3xWkpgdBbgG0Bcg/i2FH
+XWC+q1heRAOnieDSCrSRXqhUDrRM7fQ7aVlcu7ncsPLnErZgfaFddHrIlbOCk5G
8NPMILOUav4XuD49h7mPmb6bHkSR9AecvlRN5pITa/GmnYGOYsC16lJqoJ9/jHvA
Y2GpKGK4hCPiOZrsjvGAmmKLOPFtpycUmEIsezfpGP9kxHoG6ZP/3rt8bzXWF3ej
9gwCorrOCOorn6/W8uwfPGYO0RZ+N1xZ1iyKvZ2I4L9jMIKH7H7ma9ZHMRsj+o1c
HAir1N8UKDXB0PLWO9U8BDVs+lE77VukAq3jWjltGqiKZefNrCX8RTpiIKPMKQ0/
kFkCAV2khuPDiM7RqnxhFp4/QzYtFEziJRZk0M5bHyYAogctRw5rMnMYA7SvuBoi
+U2wb3qX/zLyY8tNZeGBSq4CUlMLjj2Q/3h7x+J+Tm68hjqyp5dIN50m0oH1NtH6
ZIf5RIHGAP1nbew/QV9S3THIt94iXtYBkF7cRDXOZ+eHZTxPj9ZGO05095lbY1GF
cdxk3J0Vw5DDKuGLA842NIo1eJJVjEAOWwi60tchvLfgx8eF91BWl43wEv+74YbH
273wOu9LjApP/jy76XUtYyk/o03Y68TqDVoWHWJnKMO2usmBxvtJH0kbm7C+9it2
G+RDlrdRvT2ghjlNFBmi+irgDsSlrxCEbAMXqhrPprW9l19CSnoGlGDO4TEJTYFD
B0lafQJyB122NF14KuEmkLVekUfqIAAUH0kjLh578ffBlY32wqGjjMCfiwHoFovX
Vd8iI7qM54L3hZAD08lFOc/daE9eXbHPOSmBO7QBsv0UumPBHHxzcg6z9XmQm1E9
aPuQ+O/o2bGNBfVMdLw7vcqvd9ib3PZCu7nLNTHSHf+WQsjkAsL+YOSIjnrngCU+
Dxc3UIyg+DnZttYskpYTXfpvrFxgeehmEpN3gIJMP6jgvRvGd6J6BeHzQt2nGwYV
t1QZ1fRXJD6BWf91AMA3NXJjalUWno6EW3wrRHmzQKPrbGFf2xNil7XFEXj5P/cG
Jv88BHMI7AeImbNCtkSoNpua5pkE+8lFT1WSHMDuHxKy8ARx6VEAPh3/TPkFdRKq
JihckdqtzFtRYPi8NzB3gVvyb177ymSmK+xUNc70/a0IvXmfEqGyqud4M63mOGaj
kvc2DqvSGUUZ5SLWS4skqtEQF8oMtTHnZY+hGuB17M/V0MYqkZGzDb3ZrXg3YTJM
KZL7SILFh69OM10zwqRcHHeGlJmmxHVOnyc11xperC8HkHcLNhvF7hldo+uPXCFt
zBQ4CBLEMiNjwoGVkLX9mttVBgkuY6ZEK0UfcEGLuLkHEVaIbvRZq1Z/w+cPwEgH
JDm+Zjbd1CnP0yYzLLYVeFk2Sj53lHVoKyVKFTT1pVXhDO9oV2joWYCg8Ff27Dgg
VxnBhtLQN6JkENMuMwfcVwb1aNMQqinI26XgSjup0PA6SynsKIKihm4Pf4gjVMMp
oY+jkwSn/WUf8KnRIbsHotdkI5Q3N3x80m0NINTqcCFiNMtNMIxTMeqC+oC6F552
5xifY6d03tv27JZhgZw4HNck6Ix9WkjcFOtKndmhMXXA91WWLtIStWkIzcjzvN/Z
XMTCk0IYC4gu99fqDyAqcPRc6oM4gPeRT1VNTqH3XQYiqoh/4iwZOEqwCACJhzjQ
S2sxBkVJsItR5IuHfuXDg4tTRa5uSP8ZL2DPGlWiiV1A4F9oW1kr9qUtQFrn2sjG
sdNUo+sZc9iM5cnLQSCxcDa9Ra3BiP3pwdxfK68tmMN0suFAg9ExuCypvMsggyiy
cnmBFRiomXTWsh7PDDq6lfaqHvMr5QWzGyEoIaqBn91ckXzyGkazf+YAIDsZ/8dj
SSbMQf6lK9hNvHgA6Eyv0fsU+clfPptO7i6K59QW8rOezuoHlQs52CbBAG5XOQRM
JSgrcleqj3ikT9OUsPsY0NM8Xwdj+T7CHuRhwITxm5GezoSSKWlYV8aMr2ysjb/W
OkwTZTnjr5joD7DOhAbyuk2nzEbWRSr+0icMe3m0r1y7g/Bg678k0Ic9TX6liPHP
2LaqoCjHfGKKlt2HY3W/8fvvAUPH6zQUjFn9m2STIQkEpgzZ7cbNz82nzZdtlsq+
rNLr5MyEguZ91VjnNvNhMjLe5VEx3PntIsxteDBfVdqgppPoXScWwFlseS9Elqvs
k6TBIhB/sjuxV88S2U3ewT0Ehu3lxV14wdB0D2WdbBVyLBAxFQ+AGFUnCOiNWa5R
`protect END_PROTECTED
