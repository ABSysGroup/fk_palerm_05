`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1JfNm6QbNihQDoRaPKtrZcvU67VuQXDSHnFi2XPD65WKn9DKm8j48KSfgVvC3IXi
gfotyp4eVaBPrfRfDmQWKmXqdgjpqYf689Dya75TjusyN1MgIYKMqWIU1MM38k4p
BLvIryGPUMFit/ie75DQ0gYWwzkg5au4L24H5zJkR492+czia+YdrYgoX7pWx1pV
OtbFFAWATmy/z9gd8NwHBvLu5WNNcVQSbbv0+AQ30JtROuK1XP7hxg97Gy3ZV+DT
+6pD6p8m5E9Y97zmUYheAHjtVj7qrZiVthe9Pn15whLtL+6vkGcEQxd/tpDkwhgQ
l4CWhMjksFxynHJGtvWKQUReuM21RgfeTG+Qlj/wlE7smKMfMFk/at+CxjM9j9Hp
GZEtVYlqsatpZH0Gl2t99e6hdXsG1zmW4ivTjfPWRCR0GtdLQqUqzjS5bt+oQK0D
yc12v5sBwAj8u7m3ObS4dKJ00QDLG9+u8Yuwhv7faJyLCpSTOKq/YW8R1oh8HWbi
XK/frr3O81Orpe8S5dnlnxaEzwRkM0WE4TB+oW+1lI9dlHE3pN9mkf/Nkn5TBhcg
r8K6xC8Tl5aFj/bjc7QeRoEiJR9WA91q+Je87WGpudCpduS0bWkjwnXwe6txMP0A
792EyD9viLZRTTFrFCgFOVZndL9H00OXg5d1evWk4zQ13GrV1gY5OUSex0PvYF3L
yxPPsddEBpKT2io7VuO+6PnGtAXJt9NOhidx0ilsYdrvYBVVcvleXM+7ACX4iZ3C
bzTnCeLA1494Rfvy7myrmMm7R+moOM3RAPgjDWaLgWVMI96R98RBS/kwzWOZM7t8
vhQxDYnjT1pnyXJNuapxlX9FUxKkd7NzRKZCl3vZYPYl8J3gwEwrq8nFyF5u/mmi
y/om/IBXlj38BTLtyeTpHufK9VD/jZ9GN4ebwr+SzfHQuST9KBvN2FoWg40zP2QQ
2caIOjDYc/2Wz99oTj+GGNgOVVn7P1BFe5Zf+pEoBmkkY9QW55mLjOEXkx801rkY
llbi2JchmiNC2sI09PFa0ATqDbuclreUBvmyunrUzI2BsyAX3IcjdAD2DfltRnvp
rDAhNF1s7oMsqffITeKDGxTIfIQCEj1Sx6B9dxZE0CNHbegxQHzEphQKRIYrGhXR
oICNbsd5Hkp5xaXlWfreVufV+/trRgXI4rW8FZqh7CC7MQjI6MSYnnTg82Lu1Jrt
/PBQbPSFG4Uy3wpqK7VnIoWb4UdO4FPtYGpiAkymzLz6yMZZhLWB8LLX6w6iRAVf
wAZUnB4hJrtEs6KZsdSCOrmkzmMOrJncE7lEuxVEEOtyxMLqvENQNEBQaVIqGj0s
P/3YoyA3Shk/gDNlVZoTwgdBXW42cbjdOzXTk5ncaQJ+X+mhvAp+Fi+xhg2SOwVH
fRHCspau7KFiOFXeCS6RK/Uw4nlpOzMNPcyzRG1l2yq+8Ut19/aTBX0DUdokw9Z1
srfRa2HREKspqgUXj/4HcYCsQ9oZV7UY0Nab/Y+BeQOh3pDMH7bKcQJdpUTptJXg
j2BGQkLAEA42HImR5Q9C+7YZOgAHJ7kxdl1fXwgQhOMzw/klCJgYwb5gwKnMwlCX
lo1nt5+GEU3KddnyXz7V1wULCxUaK+JEUgkrneBfWv8O0fa5eBs6nnJETx7Ktiih
lNP7LSA5lIHY+zvqMXQmjg==
`protect END_PROTECTED
