`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DUiqgUIg6dZPp1R69I/ALN6obmniZuIp8ld01aAB0VlQR9U/HIXHSpPL53C7L7jy
/ESE4uwI9LhvnL2lWQ4EGGxhe3Ztj9RTrwy7Ot8A3obrR1tmmskfHZFNQP2JlGYA
Tm4V26ZFmeN/cKdj6a75m2e6IFSx1hlYP0e/SKPxjF79NM90AyudrPviMMFXZmHe
We9KG3V1puUFsGJGwW1EWR1XzyHZlz2wvVrMf/FaibBEMnc5ueubULEF0llvJ3Kk
0+oa+JL74Ft/0VVf63nJtJ1ZEnZh9SoPjlBblYYsX+M5WnzW+jHEvMc3H80lXRBt
Iw9lnIACSlMXlDB1/g8WJ6hhu2sEISWoCcNAnlFSwn0pT+nzPIP5MkpkrBy/O/F0
jN5kc5IzJNoVp3V4Tvoe2A+46Qbcj8J+NmG3SeRI0mSfBeN31MXWnCvgYNm6AUGV
+VBhsfDqQWmFdPRcrf8odIuE7W1342rmRixctSw+hdtBPrk9x/YSJdAVech3HnAY
wVtYRF1JGwrBWgGMnSKEcFUL+cpxgDKC9CQhMofDg0RYgeEh6cPy8R70IJXaXHJz
dBCduII7dJwKAs6Dhig2rgwYrUtJM9tby+GqI8yqVMcCod/+pHCXYnlWL1/p/9d+
wNzXLH3JGFNccnvaOTY3yWl3ozcuLvSNpvU9QAV6Fcg=
`protect END_PROTECTED
