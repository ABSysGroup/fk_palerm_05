`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7an3yYRHdkndFSWj6joRIn6rq9/6U59c8smVBPe0XVkQ3y0vPT82yybJTC6qycTd
yh9WPuMnAyDiOhzNxpwO8/yJKWiESj4MW1zf+Dxz0TVhH6uJsPFfcN0Jqubj27cM
f81nK0UETbAuN+EOOe39SArsj5uHNT53EAsscxIDOXwReAjLM74QSIkKCbiG1O+h
/3bxIA0wGEEam2D6bBZHjWkK0+4bzGi4RZ2aViNGUXJE2Ulj36kKVSBQg3z1p3hz
ST/c7x2C1wzqN3kMx0LpY1zO7h4rGSvh3xAOfwRTGNbX6+Ul4YxvqDPShB5dPLdG
M65qaTKGJJ9GfVKU1gRZdlSclDiWfQC9FNuqAU2TtNrlbgJE/kmECOTxb+WwP9Cg
AQTUMgqMly2YdZZhHBm+3RNl7P3w0SLEO8dgKIjSOgqa2eafmrGz1PVyJnaQ1OqM
FRr84JNknvq+KddZ42GgZB2r3H2OiMGCOKu8XKh1lDChX9awzNDs8W0f9rCuJMyM
+6umY0HjRdqaBEhcWkDiFwf3yU/6eplp9PCMkQeNdrYlQ5qMskyjrUKGFfKcoqzi
goi9T+qUsLFuaF0WZFDyqcODEiukjWwE4ZxRWcGVz1mbVn+sGev2eyqLvGfRNx1d
X1h46ASZj7YHshGNfL6blzGPlk/plhdPR/P0dmDtTik8J8FRdk08WKIlHtKTsdeh
mXvrjoLWL7bnCLmKM+GaPkxP4S08g1FGKZ8tf+DtiWh6zurkTGoAUmu4LYoEIGu1
efsXgXhwCeCpNBQeUpJEa0QUie/LIMnLUYJiOjdxxCnZ76Rl+dSKpXURlAmPAbJ0
RTOR+VJpYg7haV3I7MyFa50kbA4jXXliOPZAvcYFwYg/xsWFHDsv2GgM8xIyMqGJ
wVCujAaDBQy2oI0VPyHaGHd7Ed8TAlpfpB8QsZ6RkLRetDwqPHwJMcrH7QD03dmx
Txe/dNLeToO/lgYv5F3MnGrm3zGr8K+Vvz+0pIuLd1PJ+4RjRejoM+Edz+VO+Yx9
sWpH1eAAsTIOzLooSGU+FrNBytnEIAcIxEA8CsJ6v2NZB8Uc1pkrrjQQyr0R031b
jqk28pwHpEh3PXfCknEY+YZGdmWxAzqazvQViDK4LYQqm9/LZvOrXjKERo5r1qEZ
3xdpdIy+Q3xwtSdyf4S4o3nLK1tAiWAIeZxS+tIoGSWonfM04NoqDazn+FpcuiPk
NJT18EmWNtOrojvvB9lnJESE9e1/Yfhxi97SsDinav49Q0gGV3A20SSlghZqE/Ge
1eHINfvmyiGGrasKMQ9cwxflGv6BkJ2NcBMj1k29fpqEhxrivVLuOEiEbP4wQ+x9
dvyr6KJY3fcl9Vr7aRPnENPyzqEcz9TS9Jvt2vPBXt62TS4x++HuUy8stwLjghzC
QRBU7X2O1QdmoKq2/HAyTuT2Qo1XopwaeNPWintS1+VCxO87vCrZyiute49fFnUp
ctfQeGMaAr0rZsesRMud0Xuy1j5xsAYPLD8qI8wKTx/8a9ry2Ooura5rS+zNHIZJ
XwpCaP5pF2C6F+KUrHioMNrx/Cer5UKLKTiouqj/VvrILrokWWiFEvP0/kTwahUc
8TkUtL51hjMzZZHOtyJotRT5uD9cEe9kIs8b/nFysNLRWCiazfNjnpn+PswAAJoI
gP8B/cX5EYtWGM1cOO3re6iJGDBdYpmwY4L0j6rNYWHJh5hRSGQxODYw/2hpmux7
h1QRTcefdDwT+6oZ4uzTpU8PdMV6ko9g0xOhHt0hXH7VdVXV5PYLyZN9IuDN1+wx
dyLeMEKKDu80tzEyBaJ0XL0epaRzujQArZPSxvdGLU1rBmdSeTKkvylZIjUSYQq5
jDFkaRbbOpl3ovHwpgnanRqrs7o/6bgEFQ1wprSZt0mytAZaBAPbsQn6KQ7aEBrb
im1gVletUTXQYibRUIPDPvQ96nFc45HNzhuP6zrIgSg2BznIsR9Mg/7GB08zdZ9y
cCkPTPtsTTTf+jG5wK21lG4D3SsCU+QmhCBuQDtNlJFZa5BVqUJ+SZOuToruNl5b
OgZuOOFMLLL1TxA93IYEAejx6wpy0/VDmd5jWefDvO7FjSaex6TDtmdqtGE3XmaF
9Rw1vmQ2LDSDZvCohQlyWn+y3ZxZA2YrzHx3HJQW3y8=
`protect END_PROTECTED
