`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bYLdHBR0rggC8UwkXsHafV9E9NKR9pobN7C0JXWb7OX/sSd2Ah/oB0kYFTlr2ggS
B8P91ddwmwb1olcFdi6UQvf4EDBFTVFij5bvBocy9+mGSge/eQGDVMXgCXJPyIIv
zGFUZukLY/fjSzCrwZKifdqyUPafPeg6n1rX9sv79t/K9H5pN87qP73ITUuW7/Ar
Q4Qbt5iXfxBMU7QDkvb5UDrqYQyxPXnwo7/boZ3c19h3TbYYW4nt6403I07oSTGT
bg0AvGw5oBQ2tMmWJi7LndEqSMA73MIdcseDf2wMCkiKZofijmv3RRa7T9/h8RlB
AQXKn+9DcIIRAekvTZVvr/lXTCyD8a4OaIwHBrPFM3pKh7NHwByzHhOM33pEoknm
Z38ACjPRTDXUrzXRvO+4VCyqDoetfsi00SkKmD9bzGw=
`protect END_PROTECTED
