`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aLh2phP4uHUjh0BsrnEh40OoKfGtNWwCE6d5TLgaZKvg5k/n9jnXfZDgtEyhT6uq
CQNDS2QkF999UL7j8gtB+oFfoUO21OgpkZkFeBz+eSmYcB/LDXPG1d25pm76Qto5
edv937E+SJFRw1B3a1ewrVSX0ESsWuvdyGxyrzS4GzVKEytio7RPrsYbukWlUQGT
zjuoxJmDlC3rwQCuT7xjpeeWkQg3aj8nG1jX4rB9xdoHhSBD4gPE8OemQl8Cjlqz
oLXpPHqOyr9MStrJU/KJW7jbPRavHlBPhwp/Rmt1AyesBF8VC10DWWQIF879NfuS
x1JaMFiglfICL3fypcLYijokML9GoDKPphsuosA2l8w+R+JmIdRn7WlO1CXayzDg
lXdtLL2XGXi5WXyOZB1S3R1qhi5/Y+XFOp9mwr5DohbWf9TaNpaSer7Xq5UFsQO6
Wc6H64a0yzJun6zePdMg83mfWSZQaXTqyc9/gXhA2dGl56fwvzaEZwJixcszhk5r
3Oedhi/vcN8q0VislXSjxgMAfVqVzIVxi4m/ecp2kl0njAvE17nSOExncRLpTtCT
9CKhIGXCTLLtSjB7OiB8vyYxHKqp0xsUASgffeLxat14EFej3CUbazXmmdc2nr9Q
jlG2M7sWdXZAfBMRF2EgK5dtI0zfiIfjKtHzTqpx+A8eYuMjKzayn3ow6UBWviI+
Dfa6Ssbr6+57WXwwlNXL7pIix+S76m97JlXQoDJcrYiaRjMdLUs/sJXGjIDFjSb0
MQOUvK/Hm4YCZI78jbqlpYsNB/LI5XGMqbN0afETZ2kTcSOR2nqelbgwPuap+Pvx
rw3+N/gIZjyLONmotBx+8RV39hjqliQPt2TTkOEIb9o0YiHicJrtVjjUCg0UqvQo
5uBw1tX6r9A1pfOaU/WNR5XMVrguKh2SYBo3zMoIbwmAq7QUV8h9lxGeTeHNO5eR
tC4y/ACtjJNvhrGqr0TK5nI0M+H4RqmDFGGyxaSjWl1Jd3VnS71KLn45EPJo5pau
6oDomcDk6ma3nMn1LDfmla0jdIkhvJXHWMhxa6lxd/xFMSyZG7OBr/6Fxx3K9Vbd
Tb43zD2qetHZVS64MAAJF8sQqetzWhZIEGvAhcMlVB7S+f1on3D60DFuKkVW0TT9
r9/DUdCg1fr0tyK/c6dSrj4BvMYyUgJTnDBziP+3iBYA3Zs9KzGBKh+2BuUBOgqI
f6Ipexbzi/BWjYTVNwovQK1VUdByLgcaew1iaOXovI92JaVxZKbFZArO2T5XpUET
opoNV0neHwgKsZdupwxJTP7LZ1M2rDOXBbAvKLxTyMTkTcHE4tJH8Dnp+Hw+cKWr
qKOH+fkNpzQURCZWRmlEFk21FDlD1qqPdojEC6EJFzWDerWgJZcD/PXqDj3BpnZQ
E0fR/7QAvAua2c78vgOOR3uY3qeneSeJZOmAH6eEIu7haEPOEipvjX4o9dr0e0kd
Wt6/D2QyuwdLrLy88T47DEZTFBWCo4Ot3+7NuTdiRThYKQlPoqQFctedddVRGaHI
mTaimCNG3ugy2f56L0vJFN61r4C48hgjFPx+T58ZvUcAO1HmeCXqwyK10mK7sxUP
R7b9RQwEawaedqnx45raYMKuSXNkMFIJ6rj9LybGnbfrNpqk0fvtHY9OfGBhftri
/wQmOO+r1Dvis0JRnJ+mcUeLd0dxuEnt3pb5qmCjQzWkIZiRq8Fr9L76X+LngaUi
tC7RAUwe7RZsaaU4L+iF4x24d9jOI9tZJDMkBLHBUPqzxlaC/dWcfFuUtWIIP9OT
IfKN2GzOLTSjHUK1WIeZJEnGyzJwN4+wBme1z8gyQV5mrqiyXvf2jiruBLzyUHRx
ME+b52PWYf3fNaBEFWnpU2XBEvdhE0A4OuIOQPr9bZqgj5z6CxVFhTxWzF+Q9cYH
JcUjXoePGO1DeVZL9Uo72XkrtDdgdfDOZSTJSXlkm+gnlRXYSOWOO8BHHDJ/4DIz
KWqwx3sCNscmr/Nrp30j5Fb5Myry7RbPYY4L6F8N+0ZIZy7sjpWduwIrOZBSt02G
n8epXumFhp4XDSVlpIHEjL8fPxbiONQ8WzTtEClh/eotYMD36HsUHM8InPRX+Lk2
FPNISE1JOr45VZpQX3gNyizFdCh2YP6T4M6dbuszS+0=
`protect END_PROTECTED
