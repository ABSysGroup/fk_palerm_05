`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FgqLY2IXkm1GyO36HKwO2atxhSrpgbU1qXA/2OtjCnlt+dufevyiaQ8F8qO/qpn3
j0QfJ5UIPNU3+jq4AvKVARIp8/JHMfm+tjxbzbQ97ADzrBwPoqLALJKFlMHhitQ/
JwLDe6eSFkeGhWCfsTKnnlqCT/QQEAYPxdxCzPYriXMzWo3cT2RJ5kcIY/hAhx1L
xDUZ9K+jfJJ9AS+9KzDOc+FbIvbSbvoM8wToAWeNekhuuF6LVCfnLYYtASbbLtQI
/zVcI6ponY39WHGQsGDJ7TZZt6AnYeVA4heJ8t2rAvhinkkchjSCw/q9iTlUJH/i
eVU9dHkSXpNWszVRhEw0sR0+Vk+LD13Oq3KKY3wgye9YmeYR3DRqgoQyrzYLUFOr
2AkqRRdU00xXT9T9X6Zxxh7tabnt3cwK4vG4nosH2HWjd2owmHLt0OHQ5+hKzeFY
RV0gnquA4tIkT/i3725rcqUuqGIpOxLDdy+f1aafNtkrI5RuIF7N02TnzJuEJZM7
Wmy1B0PosahFWJ5jUOyyf+sTej4DwdQFgnW+fW6cMrGYRkV2C/snYy7X9w2ryQyn
ib1wlfDMTMARJQg3fQzozwRxMjDi4ihGfJwJwZceaxZd54I22+gD6NhjzLUcICFe
hZWoz/F9aEU7ZCkx31iz88jUBcczLWTDhMg5ugSocgkZ7gP3do8TZmzCYuEABN/D
fLFMs4OoJqhDtJCugzoJSqxQTMBuR5my2T7pYFo9IgWl+QQuyYqQrX1+GIzO9FvV
oq6gL2b5XMW5nb3BY9fm8t57kBqw99ywf1WuhHktpY0oVPcfwPb+byn4CcMqYAzb
LdX+J6cbznBzQK+l+u4vZg9hlqpS8iY4XKbAp10tOh2LN1U+aA0DKYK+NtOS6VU5
OaiqYqKTb8AbDPy/HCHXoESzox1uFN4pctPy5AaestQJLGJq6usriDkuCMqy4YiP
`protect END_PROTECTED
