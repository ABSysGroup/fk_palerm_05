`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CBn8B2RP6cll6LE4Keg6bpTKB+MNKp4mY0ysz9780F1atllE70tlLm/tWr8gWOMk
O/p60hf78v8c9zWNOrpfQh2zDshxdiZHiqV2zrpdymfbdxTEYRjtHeKNwYwI1pW3
/60efJXkopDd0sv0lD7qVDS2wgP/SyAy9Sr3Pg+nYrhLm8ghjkiiXj7UDUZ8Bi9N
RR584k9BN0+cns2G7pxUCh2fxpstRdPQGQ38NjoAdSyeMQOzlMj/jJxxekiSHB8f
3SW8qMJqghB+wZbgf82XlEuC/G0qZtMOsLXjYpMijs5iUF4kS54kE0iluHq1+Y5f
eezjWsCokxKoXPM8ED84M7S9yV7bybLvwr3sRMzOJpXyub4TKsk4fN2sms3jm//m
2at6S1ItI4vkBVNSiYLicdluNuingbAJTs5f2GQbQNl2uKgbZSNktqCxAWakLa02
z19DMWiHAw1y+HmmTu5au2AKPwKj3wV0zNuOk9w/enf3qF5SfMQhPN+xNc99BELh
g/l5XGMwUM8Bedk46jhfWcwbJNcpPoKeIPw2S5EL9N6Wdt1CvxC2e8EY/uY+PKtF
VeJKKnr7IlFEFTEKObTZP98nFf2SqQB0bKpgLzeXRiKja3vhmk8ULU9jdDDjLPYi
/uCQoFI8bnUnm0Bnz7cz02gHhwJBZB5MFQCVibuaUkieOM0KWySkf7ibuIa8XIXx
I+0wwZnXwtU1vYztSMJSt1YBsr2++iUGluyn9CZ+zYVo1lhKvxd9P+chIo3iL5U9
Ln5zOI2YuBesCQHn2hgZO0lCsIOQ3Dpl8H4lTSdxGfR6xeaEYCRgYJ3qgW5BpHyF
MyTVs4TLukjkLx43vS2BPnXwtmmsXT/1UGmoyNS9x2ten6oGVgDxQ+Y8TSgF+KJC
gz3m7d3PeX3QQqPku3L+DDsqrXKAxkw2vyaopYBnoIEsJ6diJjGYF9uBaquOJ3g+
glAHwsT2nGVaOLPb8PprTdeHljydvJcjT4TSitWdUipjQEEHFOCAsj8TDgm/MFJW
j8krLzZoR7rsVesTwaJKnu9aT56N0lPjlGOWysRCtJgcdn2q/4fjr5C7k0Ni4qaw
cT98dW1+tQ5gKMkVbWxuq6htaSMzGpCZDkqoXTW77B5IVzX4lb3N+WN+9g6N8cJC
tMFipF2a/Hzi93ANPSO+60mOLsByCEViFPAkKqHD7V7HLLW1AVrZ2yeVsMcNY9pW
fCzd3hyjqYX4cuWWBaFiRiXHcBPK4cYMLXVt3+qzu6T58eC30s3hlb2w7L4ycIBI
`protect END_PROTECTED
