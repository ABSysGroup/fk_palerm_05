`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6LY1Nq44wtHlLBO/yDDura+jfWhypO6PhGNNdrzp5uV0S3x0jrrQq3Uyhfx8OiFS
ZuGTSRZch39TQT1oUQ5H3ug6qCNGUpptwa1soGobGr7I93vncxb7IQyu6KR+E9/L
qmDdIjBWOGn5jRFm4wEav3bupVa+GZp7Eo6fuvJemDhMKkD09XZsklyFxe1BxwBs
uq6j2lPuIYLR2NuFWgBu2WZsaUWK+I6ROhd/488wP6iOEba4riT12AcKf1XBlXY6
arfr0X9HgpZuw4zYE/pU5y1LXoeG5kPNkTUP6xJEfMc17s5qNy0UbKbxvnHjIULk
4H07okuOtVn1e4tWupXieVEU7v8hacko6tlw59AMQBQ2YoSrdjMdeJMk601N/Fps
wXKPPxU0SztTsHxjekenYEh2p6/X8TFFEW7h+UPT3D6nWCS2XLe6/rZz0ZZRPWku
ijp9dmWXZ6GLD1AEzMaxmgsJlLQMR78Nd43f95UedzeYlQ/LUa25MFm39PZkTv1s
gAgTmnG8RbV/sHeZafT+iNPlQk0JOuPXi+aolHRqpSUXYG5PHXKcgEF5lkkCmI1f
+PJ+5x8nTSMeaM2W7/fXJCHiaToms8Zl9ppT7up85xmkbbkTZfNVFY1QzptULJau
Xdv9Qzu0Z7LVwfvtuExoQHAg6Ft6CmZBhb1FXn4LB0xOkZZ5/zq/A6evlP/T8hpa
Qtotd4RhMmcz4JpNiDI1o6BUFS7e4cAHF+GzaoVOgNZGBU2XguaMlHzBFhDrx6Zu
1E1xBqdOP+3GATVyNcylPg==
`protect END_PROTECTED
