`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kw1GcD9Zb9seKw+KeTwT9yNp4lzuhyd/DWgscYXiRAsK8mcCgv7K/gETIkFqx7k4
emGP7EIjT3grkdtPfYGJLjVy/hBChdPSs/G5mFXGyY6U/+jsPxfhxSqwk5X4vUpa
kNJiv1PnUwzV4PZ3RiCiT3rtbY6LZlmHJ1cgm1xKCHSZvKnBLZpXSS+674KdKgUI
QcjQc3YzWP5p1gpRR9Bsjcb0vbYGOTMs6Y+hh27UqJPDL0UCO4DKVtAwUU2WPjeD
Bk+nH/H4upBqoCCOUsAOPNcIxIK6WyVDWo0kqs7iIj+BwNyMgUjM2VcviaaICaUT
VsFOe6m+xCJozQBOmyRa9qvBrM742IXBy5NA3B/PlIcHPkM+JPGE/89scd+FLKEP
`protect END_PROTECTED
