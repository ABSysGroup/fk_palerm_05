`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GKmdiDiXlNLcwExu5RGKCze121akwn6VxijknfV69dymj6zR/S75jYr3fArs+xGJ
M9gXH/wGkPQ7J9T3xFZ6iphy/clgWX+8Xm7z0E/MXmja0z832hK64CrOUpiJL3R1
VPrsilloT5sPo2rP85QkTY8qoqgS3flgXdf6Cm5t7ptKG3b74gi1HA3ekaBmjkmw
dOY00HHzq2Kkt6eiUogU1OSq8tCHUDyMBgZkIajV7pXFlywblFhAln/uWuMWadvb
SA/Hllth161ujU1Qg2VF/gydqz1DKLXmotXeotaDkS9qt6f0aHptnFl/n9l40CNx
+HOlpC88VD7zNmj+8zeN/w==
`protect END_PROTECTED
