`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Vej2apC9FYE7mDZkVvEVUpSSUngbuRpB91//726F01gAr8cIw7QRyHjm87kcElS
aXXa9qYMBZ3AdhyGAMIydnGBBqOpHrrxCgR9HxhOK5hqlyEDW1DtLtQgqf3d1R89
h8YS4+9en4HOyKPRYoqvmTvBKNv29ith1XXyqFw4GkfpXqbf7nciO5EvtQNYhKw2
Lve4EZNxihobZxLjtozB0Liy1WT8l/4/4zT7WjYcM2xRfOw/lVeUn8bH3ll+BauA
kc6vcb2whxF2507ewImMkvkIHfPoOi9uiuGkHSR8Po5bnxg4XZ+tVuEZlv3y8260
nCWOPOi8Ei+/4D3tY8apVekIQ6wzo5YzpIa4SmCwakMwYOtT61bv3Qb42urfEt7C
c7HcgKD6TUEBdNnbMoFengvPa2pZOpgS468Wh3Z4YQcFoNYQAukIkTdSOvIZVMI5
t2oDYTsJuzmMb1EqJHdhr2twbHxq6yDjVD4+7A6W+T++qHbOPp3y6Ec5kkDuxd4h
rLqDXBkx6OLZWqoNRefR/LUguYTq1bSmukTceSAp9hKXzRR1EcqPf05vy3eE6kwA
epJSFz4np8Wsf3zZf17I3rMr+/G+OPLMnT25KpaDMmeY4B/NpJUpTM2wO5SNdisH
9Nsd6aWB6o0b1S4g7sGqAA==
`protect END_PROTECTED
