`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w9p1VFvx7FyczDYr05Lq5A+UbTStsr+mBozssO/w1R0TJXcTUmXz75KMrAMnfmtY
illgrXZ1XyraaOsb6M4B9ndinQG1dDfyr0zPx8IptnG4uRD8xOOwcPb1b/j3IGxx
5SXGRRS4dQ0mn3Tqy6pmR0Vf4RhHUDql0GtgeOKyWWXvP94aaKS551JXNQCYlW66
wT2OcAOkEwpc3LxoVZ7NAak2uHnHUVIAs4ztrxBbfqBYVSypsHEB/bEESUg6WIhl
wbUQfoMVHdcHDFa4SEoYP6ffEPItEc0rbPihFQ6xYiNUlM0FIxz8tGiByzPa1gXz
Ry5qXgW9PHKU8/md+dBfA7UsH9O6kLG6pWfsle02zpuWPhUlYY/BGYldUGYMB6Xo
ULDEDIKj9Y/mq5ZcmJolCQqE++qWX0i43dYknabtS7QM3CiRp/727XEmaSobH5aq
vRrx35E6XRajQzegebkuHtKAHQA2i8zRYprIc8+8MOkmjlAFANeMJ1VHyFvC0JJD
3BZAqXXCDUBX9vK9pI/OVrYDegujHah3JYWpdRqOlLzjUErwBDJRWp2oTgO3V1dx
CTv0DPhD7y295uMrl5kmSpuBbfexrqyv89v36zDAUdRFW5PUAMs0WouvmlyiTJSn
0y5jZworD7SjK7DcCKyB3WnjkCieDREowAbiCVvCnaJRNCmBppUnfcrhGmKgZogi
PZy2YEU7Xqjb6b1yPX5CQsDFUHEN3qAoea5GhsWqbvTF8QNLU9wI2S4i4bF5fKcs
akTimhyGJQBs+6W1PaMMGXV23YdWQFVNTLWZZ8wE2gfpR3IdVbaMiYdZH1Rq8Qnd
jrK08TrhuSoKkqwQE5FT1+z3YY0Tjg29hw9JeFgkpt2gjaGplZVdXmB9d+Mi6i9i
22fc3tgJz25Q9SLMkeO2Hwb4Tl/BQgQgbW9tzjJzWgQZhnqTTrBRlecTA3V0lQYR
ds5F5vwE/lTVnxVvBJ/SAKBSWdp0BeM1vgdVk+KKK8dqldirY19lr5w4hC6qH+U0
x2Ya7kqvY/N06pY4pvxHh/QWgYFWBN7G2psbovgia7n2P5JLgAT2yiGxFMP4xLfM
0a0Dzx+RvAQ1UhwwT7uPjHgdthUlQ3n4KajqRTakPsXuX/17ly3TvDU9lq8qRbQn
Ek4YL8hmUPzpntHrppFOWd0EgNq7yOBtAcUtUm0Ft2Kx8Gh7Kr2cYg3UBjBRUz84
wByCBEIvvBzPvd8nYPSdV69e4WyNsqBw1+exgMUnXVDieQY2znGpURbJg4sjsRhL
0xvuZM8ivaNZbQONrXvgBogtW3ZH6WnhExtrmrl03wyk1vl4QRY2faTd4wigB91K
Sep0huHp1R3w45lJ55oitClS6m82h46EzH+Q2Op62QZTc2KD7itVwhtSecXxPRaa
M81M9Hr/vU2vAPS6r/ugUdNw/SIeFTqwnzFiBwyiEEQrEO0XL3OSun86qPbEddeh
h3S7PKH4HJjK87U4RjCROtd6MdLxOfNupt9j9s1EhtkMqLzkQfRWj0eLIaNY43Ix
A9HoJCL3KrbqDwvnXDibEQws66SeQQnGdLIKQKP+37Y1WucqkzrWAS6Gs8tXDJ4E
n2qik3ua20sAWLRFEcU6O9TdKPvuoXVrM1yWmHAd/gL70pjkvt3lGlRoEo3Kiy5e
xJSJkryMZ7O7RtfDPok+Q76APpBjj8jZXG3Jmp8e1/1YtLuGuB/DsDtKsUWbx3fm
C4CmITXaLrRNMl64HCFIgM9BmNvku+JlM1pbbA7X96iCOXNvwoszOQJFsIFugzv8
DuNH1OsLHek0P0nSESxEUf1+Q2lq6ReNaf2K68fKgU3/492UkCFUWkU5ZLAS34Jc
Es2OwrEu4H3fseZebiBHLA==
`protect END_PROTECTED
