`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uhRT20BG4jR/ssl+7Gr23aeRz8CY7p8OShBXIvNpxBxKwNrJhvSwJZhEXG+tEdpW
GFpaq7Fh/9FHBKrS9ABTBlDR+O+DgQIj7o+KLfBL+jsqIwq8NmMfgYNJYU60YOA+
34nMAFpw5dnLFwCoKWvGjmL44m6t8GmXhBkBVOW+1LqRXxFgw3KWktgfYDQ2VF6i
iyfszqFRl0Gp8WDtKaMXAIcmPdUO6TPT/2ctdLhxTz1s+mWordMXQlavTfaySQFw
r9Y3aeVAMHvIe3ieoaAa41G42EUBHWRc6rGoeeB8Npy+PBpvRMsiswLkFdNkOF0g
/OpTtJa2NK0ol1TSGLff4C4cBpfORmcddwshg48nOgcbKekY1RebFiUth1ff5zS/
+CQtFWE9oGA3EKjk3FymQrUem4AMy5paRoHDlmxt/z6cuRvjEBghVsZQF8p6KF8L
2bAwcyYaVcRlBOqZI+8YSkWSvpJbAeG6NGsR2bOPae1ELCoFmvr6lKOLgpVYt8zZ
X73+K7pAR3Uao9LKaYvFRFn4fJ5CGA+YyOydzXpkFITl0i4uOyS255asdWczQuf6
lriOqrWgwASgGtatLN3zKp0JRB9U7MTjN5iDiIan6fIQVYgrZ0w/Q1KWKGz6Tdur
PZ5WTcaJG8YCk6tPkqTvn4fDU81NkhdhzGAhilf8UThaWraJT8rqieaDdnzUhVaG
hkK14ai23OhBcInBa1RCWb1Hgh9H7jzbZqKQ8CfzChMqZR1Ck0UDxDgSpIil2aCK
0WOYohHRqz4sHwexCsRfuv9lV5YH/zhsdkItRh8+5CJ/JKat0QMzww0Twhv+2Sn2
raawRq6OuKGebKXsQ8W5dgVlQt7OtlbQrVZzRh2H1RiWAcB9wasPRjDmDn2v1r7c
lXTGaqnkivklmFBUDO3DuGeXqxBwaSnmV+fZKxLAIOY=
`protect END_PROTECTED
