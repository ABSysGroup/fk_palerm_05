`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/w/Lc5VP4zAIXWBGTVCzZ56e0rqzQuNZTRACrH4OtcFjDHjipUXvGGgZbpT83Dhe
mqEuTIsfVB7MmvuwytxLlDFqgFKh5rmjWp/IWSAPfvci1GVQAjFQFYAzMvwgSKmY
dNb+QKIZALta55q3qXKwyE7GMDG0gwadIw96Cm0/zw244f1B/0CR6vXABLDiKIpX
uWJoVX4RH4q6DegNM/XsxeLHvloL0ajkJ7ipGrunVkcPKz2gIyAqmabzA4Yq9eLS
ClmWKFEoQ6aK9xVEQnHWlZFV/WPMo7icihWGw+fGYC8CTbaq6u2xN010mzzKYHCB
J9l63gSRS+1WNXP2xnPacFR4q3UFD8i7nr0pe0lBCXswgs6WWqZrN6s5gHCzD5IO
OT2fSYA6NAyyaX+9a6R/2K5cmemNRsDYzfQPw2r1LDgzsA+j26w2leJ9HonrkM08
oue4X6QgIqLXw/uvt7ZrLcy4623+nuiFbVSTz5cekBiNh0mhvxEJASCy/x2brjka
eM8LSYJhCoSfHet11uXTZ2zdAi4WbtRZ1nGz9qPIItocBVWrypWvTO6iLgVyzZzK
8OUllsioJeLYNiMX8RjhHzgKWz/08G9ioYbEG1QNj95SNMhTqDCoUBvp6e3hd3t+
/MlpIvzZje0WWISQXvdKE0Wptf4rO7l9tn+pPTmaUB5VAda1hbGh63iyAfot0TP+
NZ9EUFxukUxO5RW3pA9eLzd87+LImXEtO7FrRsuuvp6JukQNsS2u9FGZ1fznP2vh
TBwNMnNqvT2P4N6BbQuLJ1n7KUCrwmLDXEMs9KZWn7/OuvMnNnAAbXLI0wjCoPXI
zJKR5mWB1GyPsYZ5Jy67qm0oUt81JotUQ/SCi/s0MnhhX5op/NOXjRWBqK7a25B9
tL+rmXd0+Vsm9OdJWhXCZr0e7OIXKOKLcBmGZ0LBMnDuUI3Hbw8yApMxQAj35IuO
4upOlqj7xKx/H9+RwEqrlvJkeR9NqFAIbi8zS1zGAmo4+00KVqQoYJ6btq7deShq
SmsYc3tcLOOmWmuFrX8Rt/z4b8FbqeCt2nfF7OaF535z5nPDtf9N4WFnzjWx5zse
RYjG8iO0r1McJrej2+l/GFw8NtHJgiq2CLxzpT+2ytHH4wxhmBB7JbHFsYjjlldG
Pue3Gk+I9yO7wNsQ+294gk7lSHyxZs7E8klJrrhyxqW7Few0LsGxSw20qxUVNX7k
HI4YiA0sw2QPoC43Emare8k1xR4uBK0rMR9CEmxOv0AEcv1pT79UhC1baio+f+ST
Gjq7omqOpDY02vbqB3b1k+rGVcgg0Y0MFqQ+JLr6nINT5ULA4mznX2uEXBKBuPYh
IHRn8BmtgVUYDOzqUPOdj3hnwUvXLWvpXkKbjky/9E4JV05l28mdLO02d9u5mqD9
DCJL6RJRd0yvJCzWYh+IIwzO62LlcZOvqxSlCF35hH0Br3QT8bCQEk0HLnjxNOgV
IBoLPMvncIv2FeWXOfxe6KSpAb9wbkmB5DX7LpY4RTWc/CLB2BwPKE2x384druWc
GAzp/4ED8FGhznbuaC3iC7w3kUlr2UiUhQJGGCgVnvask+615yVp562TXP6SMQ4E
htXiKek6kTUXvkyUC3onk2l8gDc+zsf68wrq7xDnVvjCUcdZ9WPa+rzP92iWJOk2
C35pRthhR8t1AI8+g6bjoYMmRYZZJ8JMJOt/1lhfvAjXHzWgHHg5iifd5cxpFJq9
RobEFB3u7YjgwFgURWgcPP8eVrG6KNXcIjlxGVc+okNXCsNJ2LWfSX1Vp2xEdKYA
qkZcYW7jUbyoL92CQWPzYBjS7DrtZ45NB+kcQ/QYcho7tCP1tmwyuInaT2hlXH3p
LutdNld5ZiFPsBaNdElPjFnMA0OuPRLSb5PTRT8ItEBroVhgFVV5+qOPns1Ah8c/
ySpfNebeYASt5gyY4uUNHAQlu0zR9esEo7AA9u8Yf1Dxfnk2srm1Xuv1kk55DOXd
ogUg9ut+PbZHnF1r+ndCQFcZS96cK7AspToiY36aF9kj+z+a1hUgkU3zK35V8F5E
zCmimgPkSNOwoF/PoaVSFHMdht90uQXkhFsDlqI6edyBGEF35nAZf/A/YzaK9nBs
mvXjgUL9Yo9yuK3LUmAYFxKgc3v7rKnIvY38aYtFzyXTyuF/qD0RYE4S+FtA+9I3
`protect END_PROTECTED
