`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7y1FW4/GQlhHieI2El0MD6IlJSbrv4fjyiYUCOt/63UuowShXSwHfL+qde8wPjSV
h8RRVEw9MCz2RQVL1+hlJ9XDN7l3FDFxRwDmA5LdIEp3TKYG/TFGdtYzhLvttNzI
GGxuAKxXyLXGUvqmZQ8gYsKmIWMiDAslnAVIYUyvZ9iKbAdoxUQV5LJF7fQKR8jD
bmLLqWzxc7kViTNaGtJASP4y+B++1I+lR/31Km7rH5WtkHrkNjS1t/C8H1V1uH8R
Ini8PHatPwiMluFu4ub9Fc8YsIuEV3DaEG52E8sdc4Q=
`protect END_PROTECTED
