`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pDzYgVDmYUnCVpk9G2gXyLpl5DQ0CZ7/OTd07GAow0R+dGQZ2t96RL/E/zSd4bMm
xeFtLvDmti/heWPqv0l0cru05Mmjc9I1BXxzojQa/Ssdk/wzrw4AoL5R8iDGhE0R
fon3IIz64eVRw1yIqm69ydjifocFf46QfCbrGH8+wftPpoBqa1hmnzV5eM+haPHf
UKAOrzz3iyZS/12ePuUs0Q==
`protect END_PROTECTED
