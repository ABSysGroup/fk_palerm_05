`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NZL0FJR81WCkf8V6rAVyURgxrkOOIDUk2zm5uByh/hYFPN3rzY2K1vVNxsbtKnwC
BVFW3FS7a6qBzta11dmy5FrUD1+z01eX6UevM3zr+cLBMIZaIPbBf6NCzajeKCo8
+vmhpc13YNO4PjDK/17pjuZXeGDK3cf7C95uaVquwKxf4TEj2s1d4DJpCdTNGcxP
p5NqHp+3QI4v2yNpXyFggTUIoyVTUkf6YmOu2zEU0RsthsLNkLWlm7BOI/qxHSR6
phB1xY3dddtsPuEbxSYVrVlmY0E3eS/Nx86Xri9dC9oxiiFU6BP8pWTfvLgYS6T4
Ur8uX+Z3jGNuLOHC1EasoVYbO/UaMFmsJ1iWfzpfVsUJ46iS25C0FsHjbZKzxBzw
5nrj3yijktDVnbq9zgXJM3xjyHX0NoChnVvZQkpvGzouXcVZhT6pVpYCtCdyaxV0
jjdwTxdOdAOXFN9x5RhhbvbGreUJ5/ljzRKt+RQhUqOSd3LpFTcWaSPoUJiNGpix
iG9Agi0DklqE6WvLk9lK2Ah/eN97vLR6jM8FYm4mNhAblKHG5lNvCwRFCvSMxv8z
mtsxojQ1nvADB8ExtAkwVgY6uZGkGp1dqPl1ny9sowz2yJWiwK5qE4LwUKVpEGQb
XI4tU0brKWBs+d8e02ifYyqWJQwjhtzmMrcVvZkrO1T8c7GYkPvx3YD+HdIauBL7
pgSufxFL4cPtEGPdgr1DwMm8Xke3SGHd2JaXHg5RYf03Wj+3coK8fNbWriFucR29
qZ7dMq5jG5GVMETkM1Sf4dPHSzHvlk5T8Fv2+raeQWe7HjV5Sn/kZEoVDnTAq6hC
kVkLv6OLAoISDd+VO33aW/MtDvRt2bx3xhfBisBWbwyIyE5I7Sj9pi7o0RnPmzwV
oygSGTz4B4Qlgarv0krLUChrZnj8T92cQBjsMk3efv5O8PTBd2GZAmwp6jtre5qq
UIWHawNRCL4y0Omx7XaCncVR2qFu1xLvD5ghbbKOzfGSIvwLkoKLhhbR2FWZtQks
8sS84VRgwIcVkGFkYKTZ+RxuqNqz6crpsRSIZDNDClnv6iFZ7GkGz+3La9/FXJS2
TJwT4vqocwiDv24ms4qpTasUc6+lTSwkIalKrYL9e97xg54d76DEIM2IiIWKa4+u
pMXm5S4+sQ7C/RzzeZ/VLNZKhsNJWTKHJCDpTQhuRB8HQYANgi8lOK7uwAUs0jDO
/FHbmZDEX39f5rZJqasYGTcSKhKJcs1sqauz4xab+qewDTS5BhG7A7kVSQN36qo/
5tUaM/PIedwY0xXS5eD+z5MyY82qpIrG8xlZw5mm1QAgGTwyv8SRokcEbNmqIDeP
eJePmap3imilwhu1Yhi+0yYeLsu/GKLKdFwUCHWPFzyjlCXHFVx9P/KGN/t0Y8MV
Ck+tT7grxtYkQzod3PIITsJd67SnVL6UU4zoGygHjhVhx9z1hYaFmzSAQbqni39R
wzDbqUoHYh+AtBdFYJDT0ZfDttruN4RXs2ovfaRvVous0oYX36DvBaT+KOrK4DNt
+2tckz1zqRpirLlzwbkBYeNjL03Nu6WMPuKCzwMSe9Xq3GU6NhJkqH7zVgpfY7xG
nPBdXFnvaBC9UsB684iKG2P6zqmFB/kPvM+15fyrusaVDgMjWavxAeff5JD/VVcP
FnY0Y1/6Q1VB8H43wNtiAAJY7GOLc+dpG6XCNpWA0xH93V5XgC1fOfDaCtvqrc0f
XPWz3+Zgj+PWOU6qtJBCys9fP0tchZ/xBMmeYvLeY2IQ5vlyg4hJvB9++lOXj9BQ
vPb/wYu+K2mDgzguFU9Hj6kVYhl5ndIOKuRqK2sz1+AkDNMH/RhF7jRrS39fOos1
cY07401didUqT9CG9Ez0Buy0EO+WfZoXTSL0cmfPmbbjcUVPuWFkcHjG3skFbIRb
426gRwajcMrAZxDPha05XNNAFwNDJkuHeyUb3SvQ+6XvTaKbTjQTeVomHG2cc2Uk
iMOBUm5OLid/bSwmqCxmmfDCSEC4C7Z7lJhmE1jv3Jy9LKetO655JxMzGUHu02Ou
YRZGjPfykE0z9dGapQMCOywtgkqZ5pfcYBodjtxEuGiZgCbYhYOAU4UMkhQpRXPH
1ZIsAdDIcfQRYiRgf6SGAdOeKunFubGOg28+1rVB86/DKAhWpMsQ+0f40aZoPO6R
BLr+4vv8mIJ3lg5fbjzBHLP6HruCWVjLZczJBgy9L4YohRFWzdoou0qW6pn0Jkmy
pHlg2JYrgdY0DEy7xBcZ1fkC8/AnAWG0kc24EblmzV3UJFU+PN1dvjVBMMKbyHHp
1OPz0SX/an4DbGSNOaIdqJQAvEZp3hqB1Azo5j/fSndcloa7rizzaeprY/ZAS9GM
Aovlj3AAkBvQ2hgCFF0qMysAudzLaqNVtWgwVBqmQlpGIvimVHEkom0GqqsqRaSY
9fr1d2clDN27fvZ0NvIlN7q7xnkwAMJ5WF15Wo0rsCzGO8EX/o6mNGyIDJjxnsZm
kmJvDuIfz0src4EUPIP02becVFqE/gXQgUh7xDuQcejlskhRwADd2bWBdQi5to+Z
8yu1oagLkODHvg/Tk9wsVDwvkqr++PrZRsPR4dQ8vlTA/1SkV9OTMAO+7OrQniHp
XgHgk4iGQ1zCakk2YB75FomlHP68hRoYMYuLe4YyslNJz3CnRDLgeOuiJIohAdcp
uvWNU/9gXGuhUi2DtGmMS5GTZm+NFIYW8qE/lItrktik8guq/T3QVEAP+ir5upDy
D8jTgsnvKcSfGnYFC4HlBIQfcNhelgEMGnrJF+y8Y3aT4uBA56CeT4HHmiGqWTdy
gSIy4LXmNLL/FosMlJPxaqLeJkhCBKZI4MGjXurGqdbWjxxuqLpiEUeyK8SuhFnA
YlUeqlmtMGf7PkfLlQt7rwVmDVRbg846YxuJS6pi+BkOpaJvWXA5glO/bFdOGbxH
/uOXLQrm4tcpCxS+2U9XbIxgyT5YIDVBas4sEKBtMkj0my5/6GMxpSa6gLjfeium
XkD2T/YUc8IjqKOYlDJHlyYYbVJdOPkejHLL9r8hDnWokFxyAutcVhrxLdI0r1FD
tjUnto4FLdX46EdKUyvb77GZlLX4FffKAZ4DNO9D8qsneQSZtL10KTKlxAatFpAQ
bjnGPc+VopKB/bcrZfHc+os3kVVLZw22M/eV0mwDxhpgmDHOkrZ/Pzg4pQdJn+a+
Q+O543+l7+v44CK39v7R1X5bhXMSJobdKVsPJHEO+myfyE+jgE0fQ1dwziqa5fG3
76jZ2th07fOIS6ODirSB+rXrorTJ+aOr/wfhTaRELH5O3l+u9Woemo4aUQWSicy6
kfDSAqH6fbmxcU8K61P36SvWQwY7GHIkw+HbZC3iqVW8Z13TDFpkGdXtS7bWj8L3
vMmHIRUwVIh/8Vsbb6HfFoUz1UdZ7i8W+DE7QJN+msbqz7w9/c2ieCiyWBlEyUJx
nM9ldkWjEIVYZF1xHjKQz3AMK/NhSjI4B3cfSk4asUQz7hckn6Yj+/E3jgZjHzDz
HOS+MrHZfCI/fTnwPLsE4A5Qd73aKWyvxJDsJiNBRvcg0pFAAmteVXVhG0KP72Yp
ckhnELDKmjW+CfGrwXO3xiw/RwPSDSyn7N2xilpegjlcqNv/cW/W73W6NjxlOjp2
k3AtLzuuxcsb3wim1X2heSnRIJC+iWCnSrZD2uWt5K2QR2zgUF+PdvvS+HATJXWj
OgxkAqmTvcBxU6FN6dEJc24uT4aawOJq68ciNQaEmzkf9M7bmibvnjmQPbyUKzL4
vDvs3AzFvmDl0Gg1B/xPqHQ32Im/J2w2rbUnityq7swnm+KDEG87rUxaDrPtcxl0
dB1+q3aOu9C2sobhHEATqFDcLqJJDv0t0cfcL/BbPJnT3G3ophOFBRCnr69izJog
33/2o3V6ohSoYSTKl2t/kgoeFKxoOHpO8Fcvmok11RrmgVVhJZ9+WobKYyjHhKJa
7aIZXVZwpJ8Rodp63XgHCfvUk6LsAyytTBjfyQ5X4cP9Y7IGkbMAg2Ig05irLaJ4
9Ih9eWm6XqbuwlDfqBHeaImrj/8oIHBst7y5CkcJ2us6Q4LwLprkDk6gXhZ0+h8x
4BdRBNxC5nT4PykGTI2+Urrdy5mzOkIhTg5PF5ICf+pw2MOEWGCDIMYX2InGcm8N
4d2Kido+LGoWHMukYyh1AXJnZHgzNYhhd1k6ylhtUZl1DcTyZDC8wK4cHSqd6IvK
7H/uj0k80xuadMkaifKZyJWiawZnAFRVDZbHijKop/0QvFofZ8crreuM1CsOvB8f
jF5cDkmZkXqGrCz4oom3YB3EgYoljJ8ZAfZmz4yHq3Ez2eRoOQcDOsnoMvXFCPRB
uRQv3tLxmjX/XUU5jAwDP5ZAeAJH8j2re4o740Z2Xmd30v92uPbX6oKUWMSYSNY3
BT1NiN3e55WITNhvcFpicSpJNIiFNOg6hcqqaFWPDTOD9sjNz7Sz5lwUosdyL0zQ
lUqOnU2Tsu//x/z3E/sW7vPu6OzE8pSKtmMQECYETbuJTGIY5LBdzXbMyZcZnxUj
s/gRCKHtfQprJVgIPmhuCDjBdtFb+XC/30uGde0WykB5FW3rvZMEojEKqpsS7W0y
9h4TxKzycLjESHDxG98Y1OIwfAUk8Daf4f2DBni1WWdwdxSqZT0cHcyPc9jp51GY
Fj2wxJQzSive+EBozRaAgVRjwiXoc5sDZE6KbqdDOP7/eGVWGjZZmYtWe/tJv8QQ
Fr1fIvHjBu1BxHZ5iO1T27mtA8VeEPU2u41SuM8atGXTvg/CtcqZRxlthgrvycX1
z6J+zMJncre7EAJZyoh0XzpkNQ2c3/fkRasE4AHigjKXrt9gX9ftzUFzLYXcI9gm
BhU7Rkk/G5L15oxa1yVJ/BGXRD1Xlh70HfM1tWlPeE0MfTGl397e4Lvdz+qmg8lb
sMZ0jJuvngOdQuKkKM7lmYNDlEYaDmkTfahynnpKeDoZ9V72xPEhrlljRGSum+w6
y5Q551lOoil31CT7FdhHpmJ6svS4D21T9MRz+pab2uVPG5m4FtbTulNrqtbbH06I
fgb630azATykntOwQwQU/dxpv9c7/2WOh+AnsMKuBEmI/7sBIQSsgTNotOnhTacE
6lKWw6DsunCudHKcywvdWBjGZDPFXulcDfzIyzoQQrLN/Wqf1i7Y/AlEKMPRrvT8
aa0vkX3my8y2Fjzhcw1N0Ca/z2bJLxZjor9RK2tsfD1FGkuns93fadp7Ad28ENh2
fzGatorwZ8kNYG8bhCRtf2tbzgAAhEAj9yzPN7u/0dJdY2TP1ybuu+y0AVuI8jeM
bjigblZX44MaiFub2g8tPBspQipUqWIZROGU25eJnkCuXsxNTcAAsT/tjGSsDVCH
DaUfWlaVwXh1fAsxClFnsLoVWKyD1W7GjS/BgIt+DD9b8ThVK282QU6Ev2V7CfYp
+NidS3QMttKozvEwvLJLWey0L9EVVTvwCUGEfitFY91SiZ0X2UEeNjnyf13AqMKY
N2rXfjesa3aKKNR/Q2cRqMbCBthTNJ8/95KecbPkwgylYyNDvACOAcDS8BoxuMzW
Pfw6TnzYj99vQej2Dfl4XWTUz06kWNXoexagYtgBPO0bLC2Kq0KrEH/wef7W1GFO
wvF0RKD6tYSAkxHLZSkjPdDmGwVSpDZsoi9aZ0t1geSsQiL7/R5qFouB0m+ppxdv
6V+4qs7bf99uT6EyLMVglbGjeK+mmCC++oz3rzeM9pUBm8JGOulzVsp3L4y4U4zB
2DnXROwGBs3vgK7SPIqRu5jIh5rMSFoHEzHHppk4odaLH0eSqGqSwO9yjlQEiORj
TofOni8FL3hzNwv/l2ON9Yl85xwHWpCJDS1k9cwSFqp3kdX3RiXq5bs4ZXwDzbbL
59ihxL1kcvgpGYmzJIE0GwisYsAaJi+NIE57KlEwzo9gsJ7gBUGFTdqCd+SC3MWc
9p/zc+7QjN9c+W8xWhIG9nTQ6TatR8wi2f/SZI/pRceCI/SxulB5Gf1RE8BKyDJE
EtKYYgv71/pSxS5GuOImpwI98Leg4t95DSrlbAXSIKjUWk+blToD7Ro24IGBQFmU
LbBN0YpD08v8MaiN+MT1h1LCfKGVkgO59ZcgQsjQzuQTuiX5vDruqFvUv0h9spTQ
yNq5hmnHFvQdLVAhR1qdlbLYOL7Qe1t2MZnuXNQpyMMT7mWLXzIOZyVGTo/uBzH7
8gpd39HnfAhOHlQEAr3sdiz7oxjqyQ1NklIadAjP7JAgQkCUvmzKQeQ9Yh0TETxC
LoiR9L4vY2jtq2UWUJpPwEVl/LDzheKRD9n2mExueKM4dCQ9AQB+RzqmJgI/WZyN
E3ueWinM3FQ/pMn2HZSd/2dI8MmHeSHL/oLjcxOY1BLuksgkr5xmyuvTo68ntgyp
qIpdmygKWKkpZLqxKB740UWgegPXYU8iSkRMtxrU1BBQYg37B90yYBoQrzoMtL+6
y/VP9PFirSkrro278IL1ahxJppmCu9g2FaL6dJjOHORZ1LbxbteqJn0kDpwXKfpp
GaW/7En8Foz+qOT9gE5NTaHxJPgMScI1UY+Bh1/LP7yHba4SuqALtT7QhtzGALxl
Jev/oSbrX3vmYO13ZnUPWJHD3lrXBJf0Dgf2QJd1+qF8sAy5NRwDhqytREjY3vY+
FaAkwto1pdzfdcCBXzV36sljKbmS2lNOWeNTjt1pmHDwMaPJJCPqxQGqezTqvMLo
OtHHjGYPwPxVbYtqvDt9ddX/JUoCBkRROU0vEXLMkkAUEunyx9OQyWZFyU/f/d9B
z+vRn/ICyDGrw0RpaDNxxyd56H2eo/jjfOZJUtSOT4o0Ap5aQTpACDDQc9VhXvLR
17lahYNcXtshZLIvIWnB90ww8ZBVbe96XeV6m2ddvVcWLnaPDBHwEVo3fbK7vFr2
Xp2l5p6IObex7bq0AvvoMYJ/k6g1jcQvSxOenEwUlBI3nKi8UFcYoZ7aO1HJfDkp
P0IwEk79cIxTLU68aaAoellRLFYumIVEXPDKl00PkF3PjD7DR9S1f+lDPoAhqIc+
MaD6AQviWX7fanm9+XD1Xtq/rUWgvqWqrC0kk+g81e1WEqw3OXLierBk43tZc0mb
4NUYezeZbf/WBv5WXGrYzlPCm79ZgbWEIfJm+YLdhnZs+4e0g82dyPMCpLrzRzxK
GzBT/+zwiBB6fbNuHUxZWT91OMARTcm2opLl98I6Tnyeu4fcoKEuzt5+YD5BJslF
uC+kemeAgVKoC9kcdb0oYESmyR+X2/7o9xRTTLZi3qeN/9wyzkeCT/FQM3Ks7id6
dnEFuen5vBQE2c3y8EYCrNTFayA4ABdHF+xgQmdeBtZNEebSPfMtOswMJgOX8Dnq
oeNXgj3ymQKWioYLMu2oeA==
`protect END_PROTECTED
