`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2aex3RvCpuh5uCrlRRfjqNOKbzey9acgxXp/FWgbGfLGp9pfA+TzTYzHHVxPls0d
LIDqcWMIPb6L6RDRcN7IIhSRhG58Pf+ZeZD/QR0wprri+8elpN/dkTwtSpDYmEhm
bp5BiIMKczN2LewIt8HqCCQXfuFT5rj/82ii44LfoROP5Socrv0Wgg/53QLY2/LI
qXSAT7tD4svLGgT4Bis0ojJVWI/yKbvnVoxpzQ+daTsR6b6VVYUXCvEU5td5A7Pn
x2F4qO6/0ZcLmsxFC6MU4lUIdrvbEiB43t1m+jVOAkWiRp4jyryZWFnXJcvDB1AP
L/s99NZgUEDLxtQJ5BnK3nIEqA2zCtPOnpasW/3HOP5V+hPJ/52AyBmLiR6CYeb5
+jppjdBeQY3ge7BE1eh7GwxKzOZq9YsVjrkYFckukJ5SIT41VVFYJTjeIVfAsmGh
MSFZqie4H8cTUDCJ/2dO3EGwdPTeJkdWo1n3KyDfO6rYUpS9REgVSjBebrePuYu4
MHePfRw/KSzMEgIMNeagPjDn4XIdYZEIUtz66oVOy2yCMSRRZ0eV4Ka0LnzHV12P
K2uYdykErZ6m6vNrn1tR9pXwdTCABi7BaPG+FjMbVW/APXir02KpAsgd6XRm0TQY
o5R9D8dklmr9/Kq38WhAoE1PocVih/b3STnlNCjpimZB4Jk3gAoAjsN7opQrqfNd
+NMYUH2q7hzBiQVxThkBFga3ikq9KOjGppuwwgcn+fg0g8NaDccaz5BPUvq52ov/
BIY8d5xZrbKHgfoqnPlPYBLgBr0YVxqd8CgzOwKpVzmcHV23jJA4a+rMfN80F0Cy
3Ux5xK3V1XLDjag8sUMrub0IPfwRyXykPJcKhM01KkEabVbCth8eowuovuu3V5LY
V+ylhry7SLkMgZoh0jcMXJVZ8KwAbjAZLtSS7i5tmlsWy5A+u1aJ00BvRV8k/u2a
Tv543TgO0p1B2/ln0af7anJ9KQWCATuX/NVJD21LLuLi9GYaxBFYtn0UfNgleP9A
CHTDjI/cr7X/Tio5WujwiovO3ODJSBINS8lDx/j9f8FIWsj0utZDndsf++W2c44D
eFyCvgRUaxWjLVoqWlQovcPnZc0utm7fGrRN6s/qBPc+yUHfR6fX+ARHDoqx5S5N
rffs155J/1Un6c1D9MQxBPQOu6Sltg0JNgsC/UsSsZssJ6SZdpYU0QsGknvYxLhW
4udjgydC/WgcvkowEQRqOy2sIYTQAJEQA3v31uF1uV7tXYPjcNega2P7BhRvKbUz
KfyzbXJte1eDmZcurXm7/n7IevVEO2lub7bkl7WfENc/5ZaxfTRIOk1hoK/3IDDj
H/crNH/2tYsUqklFqfyE2j3kHbptcakEsXtfskh60LbMoV8dOXLizRPmngq0F3iS
qV+8unrlT2KiqGBOnfg8trsEZHZreDlkHrDZ3KYlgLR+VLR33ceilhbxsYYhVw7V
WlHtC2Sv6UzOt7yOj1Kjf6XbOrhV24Qj09eaHcCxQRkgkuPA9lTIHlFPjrhAWWqH
dWelCT3Ine6a0gZSsCuHKqNy4gXp73XrSSZp8xgao9MEjhQ2ZNAmiht0TFoe70oa
B17GeOAW6m1GmBrNR6Zcp3n5XMAspfdx/kQhqoEDJY4yCrOhY1WmX4Lj4tAFFgaf
Dd61OeqFSAQhMwLmijf7YpoxAkSxyd4g7fKku7BSMCsFATCAzu8HxZsDDglKgPdC
L3S4r9W/d3KIcBjPwSGArmmh2Y97zTIq0tQrPpguxXPryjE8hxhNWxW6KP2dVa+G
64GmtbyQJ00zImGiVHBdt0dcxoNB2Y2TD45vCVCK99UPrQTjSKlDNjC4Vu2+3kns
k1cN8/86BSAd8DR2xGNtest6DpzlrZENERPva1yGYag3p9ouF/T/W5/9oOKL6LYv
POsylh/XZRf4IAyYtu+R59XV2K0aKvBGqm03OMgM+OnU51PO3v63t6aRduemICXz
fM4df8s1bkbVZDgwzupH56flN6ur5r8EeXuYmhf+PSoMEpgFy+rFeibb/bUwIxzO
ULaMhZ6eBjYdU9riA1GHHmSGazGSewuNCQgSIhGu6dXGfALWYM7tRbkmBg3k963O
WlWZt/EqJomnMQmShOl+FdMAq6RGOhm5KWYwqcoJxr8=
`protect END_PROTECTED
