`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lS2zYddvGWv3lY/dXZ+FHyIuugq8GltDu61R3+8tHyUJ/d6r70OlR2dcrT4PIIl+
VNQJQ1p4MJJSKb3LlaUg73ie95aqjRjrV7cEn0Y08sMrBMcEJ60XcoVYIHO3deh6
hjwbVCPI9EXwn7aGWGk9CCuwyXm8km0NfDqQAb3/GlYTdQSVthrvmGGExCoxw0pY
Gq6kq+fUMOdspL7uESnuPKnjkiW7RAIutYagBfGEoKMycZfW/6/5oj6LlNkoA8Cs
jTDvelfmhIqnjP1U50glN29b1Jk3xCejZTiUH55orXr+JaoIs0tH0YWcadq42+5s
JIvEhjEziRE+Y/2DMvBcQ/zPuRtI9MaQ2y42EkN34sW6pygiL1AUmHQD/KYflvyj
oSQCFcbDbWST70y1u05emIbl6RhQjpLNk6g64rv68wQqgC9+UMBMSthjxG8JH8e3
ZUQxuyQC10isEeZaBleG/WZYiqMdBvupwiMui+YW4Hm49blGVvXYXXnJPP5aWJuc
1s4ADRf7dCpN1ioQVnWBO7CvD9P9cc08viejICOj7Yr1FyMDUVnNXLLuo6XbKsHL
yyBSETxtz3Z3tG15sramPt84V1ShExFbXoqo6CSLLRAjh0UBlbKVB64VaPk2e9NP
`protect END_PROTECTED
