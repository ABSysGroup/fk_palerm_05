`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uXkIwurLAtxpL/jE9wan/pW6wbdyqOC+86cG5zYpMkWaGjSw3fFIDt9MKNZwpBbo
6fEVaQe1vKHp1h4o/HF+RupE4rjrdrnpFsLZslFITiPioq8CjJVE9Epqc3foAkjE
ZTgMnwBh3O2RcjyH+C8iG8mVAh8WE0jUtTiFsuaTOOdemJpabEA2/jcjGQKfGmkp
klLvjOWyIKoCw+kxzFWB8Mzz3muVtJdkIJef+ntW0kywS8sTOKW//SM/MCjaVQNi
/orquA/gkGazDDJVmp5v5ySqJ7rh9W+LrSdiwl3YdxD7yoZbb6iA1C+FCMbGhlyT
kICTHh0RLcIqxCxfggicLsnGV1x/I6IyXQCygBrfXoSIkD4hgD3ecxmNMnqj4UTN
pmo46ltagUum6fcNluv+cneq1unP+FiI/r5V9s0eh8MqHGdMZHKWgBkElW7CIcCD
gNu/FZPrhGfxw0Lxm+HLk2/yzF7mQtUpg7c1z/ew/2XIgNxbMQYhZ6apjvRhdUvU
7Fa2HP+KiO/9euuhRmCOmKehw+BzM7FGHTUMQTUJrsatasnBgjeQNAVNMyx87cH+
woG75ANqrwwIhP3/7CGUF4XFjNwwPAH8wWuASFVcn7DHjJCRw2oZKJQd36mrvwEC
Xuyx2m4NTXJdDOZZv8HMegSaCGS3ydBxdVkIeeWZ7+d/mNKuo4f/H9seDJ3+O+ya
yCuf9H2uGa50rAxoaBBrlWMMd9M5+EaSOUV3fiDVVO6ojVZHuUEU3t0WJpdiHAL+
l/2lDhNTin8/eEHSwwVj6VLg0n5Z1BtMKfK1dbrVm44LwVAeme6gE0HmD/QjXHjA
uh663QSZFq0C6ZnbG2OKT95e4hPZucO5vp4UpIopOleoNq81sM7k1lrzozr/tmwR
oqmWLG1hyuFidX8a7jv1wDpbz8SZ/tK/X1vlbeEKHEP00ir71LBB9boQCZFajLqQ
ZLIsBDdzrtF2bgCrtwqjhZTvtebx7wPErRSXVVFIXQHd1a9ABhvgTd6+ymnPVs3k
hNtPkIs0Ui5SuKtuzFe/HDHPibRCqpVvFAS//92W38Cm7YCDuFlaINGgs4ev38RD
D3fwwNgvsz9/kb3zTDQiigLDMaLgeHApKg3yhkeAsjPe2neBa8BaydNBfuQQaf2M
E/P0xACheyZuxhFDaZOI9KqZC/YOy/mDLvpY7gX/KaIt3MZ6ucJKTvSn/rkgjonC
wWUiVb75mZxE30oBLRhYZ0KU621t9ftkkjoOMiTn0fZik1poxv9rgq4RCCnHorWh
fyCQssGzxXCw8NkHgOvoCQ==
`protect END_PROTECTED
