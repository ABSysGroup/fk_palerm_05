`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2qboz7UJquaj5tcPg5Rb8hGjtRsh9bSeO0HMI8FWaXkln44fMPNht0o4I6CDX8jh
cwnTqMn8QFT+IrEw7oWjyjcKJsjuilK0Hf+kNol9pvur681JJbhQi1YqUEbbkBNh
7t+mu0pzX5Lsj/wwtNL7cI9Gw3CckHoOxJNABgu6YDwUinBEYOAOZh7Kj2rihX2p
VHqtJGJmltltWNCGdowmAST0Bw3pbPDf2h2ZH+O/TnnuXaPGj2Cw10s/qZ0P2fWx
lA0hqbo1MInDawYpOPFBVKfpF/pDKVeQNnzOtN4nmIdMpRr7i73yV6lYdqwmo5Sx
pgn4M6D5Wh6AkVDrA+M2u5a+fnvJUnGMNnbSNbljpO+QFkfaJIN8yr02krxYAXZb
pCYtx5palG8ocCJE3UlVgPIijcOY5iWaW8qk/K/L/apM2s1wYMkwKiIp7Ia5r6Zl
uOTW2f+02m5bnNCTQzmxek60M+0OBZCHdtMFiMDofMcZ7Jd1Vfc+/gY4zwqXYBM6
NpmdOhR3sbWipjy2iAiM2tEt10zKFrLgbIp3SAaf551qcczSuAeQsbnzRKy42tuY
Tr20JRylpunYcjsKtZysl4rUO2vB9iMvw/c/yGmpQUoJ6jtVQ4XaDa2doRAp6I8y
mJvq/7n8Oz9jQ6P6Fno+B7uOAj2HouWNkN+6wtMFt9q0R01oxBHe6xGC+nEGh2C9
DZbqVwW0qJeT1yE5J0rWeZLYZOEyk5rv00XQyyEz6AJDr1V6RSEII+fIZMnQMSod
w+2vBjG7PK5H1+ktJVZsTtm2DMP42zXYb03FxBhHSpc=
`protect END_PROTECTED
