`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tGf0l3oiPpDCMdrJPwC/FxDNAW01X9zmvVsOtIai+dquIACS/WpfcaqfhqJOi91o
tsM1MHK0xNYzZSyH9rVhM7H7yRHHpswsCp2NI6KrkEs5hA2wQUbeLWRZTswoR8IZ
UOk4LePnGNRjejC1/8MeNn4yzqjzM3pyszQNvgt6fRriQEDAwB48HU7ND45wt78X
YZ22behJsBQmkzyzQrvF6aH5nxX9OYl7t/xL4Xk6Spux+Lze2qCmmwMfxRTUtyFQ
TJ4rXFhJ9nMSot9k1RR3ABRwOhxKkPNG2lbSbQdZKndcDmIR/WVSO39ZQSDBsnra
988WkfSSp7hmCGfCi9vyVEdhH8kJFpjRvPWOG/WO0tjVKVmIEz3FbxcC4JyvaHcf
L/y3A1vcn7SMux57TKLEOarYJSDKdwu2ez8IWLwiAj4Er3lWHaj7W+cJKNerMEIJ
CzoztUh20PNekO4Ff7aKRBudZD+xtMQEWYDxUd6olPNTqYUgQQfGjWx+tyU4IzSi
1sCrYhVUpRTE2d9kgy9Gi7xivpn1MZGcYub/FTRFREh8TzqLNB4u74GPXl+X1vGR
BFTneo14pSqyabqEcKb/6QJgdCSaWKw2YV8EIYcYQi3DKHN/2iplIWicJpd4G7Us
HIXF4lWEmYr2GlvQZFznF0MV1qIOyuEiI861GOEa/0LwDv8PZYPiSIWgd7V/Ia9/
EFerjHmA43GfBJddQ23/xEk2tpuWhO47j/1MWhkuHc5K4H8LOUdTF1W4d8YfVeTb
`protect END_PROTECTED
