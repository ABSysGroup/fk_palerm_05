`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EsHcrg3RibhlBiBqJr8dp1yhdGOlJxxKLVlmd/Jm68bay9y4OMFGy6PCRVhLgP3q
1qQeOrCNxuTZzHGLnF68Wd1mlrS7aYF+YjFQohWafIWsaqWk/xZr9I28R4hV2S9d
PDr4UktECzDjOGz85ZNJCEDkVkBx/lwgcnz1o1KMeDQ9Zz593ak1vjjrZ3ZTrL2q
3HDEusJ3+W3saeVMZUXvbTAkgDMWrBwkWuzMPQn4o8o/X285WedMiAQEaskYPdOZ
99lQ0PnXsKthd1XLTmWTRsc2zLhBiLvmKkfQZmfyWmx61Pyz9pcYIt469GSWCQfj
Ti8B0opEUAUepEaldyR3GjNtwhQqydIdOTYqJCsC44Bb9pKgUjXjMswjAH07Jivr
EJDFhTExxTMDHNWf3evxB/haMGvvbRkxXN1XYeIb5MNJl88sZr4VPgmrDSg2/Tj5
dk6U8jhLaYOUs+4KWrsjJ4NGSCGfMdydbVCEGuGzwVrQ0SPJ1NhmtGICGma160ZV
d9s6luH6skbT/DebrkjqlXjuHHWW8M3ODMv7Jfd1CWXjjAlDwZYajVXDfz/KR+SY
/O05nd85VO3dumGICFGvtjsszZyC2+J2LTiWbpTBizrEjyBiFvXx6rPDIRqLM5lS
VnBtml6I4CKZsaSx6g8Wr5eTSE/UCkw6eDLtmYnK+i8kGEkA91pYNY6km3+Czjc9
HIbBb/9fC5ELZTKpuoEZhWDs0JNwB0NJwjLHXVavmChjnRqATdFibU/9/UHdyOGV
ePR5zBDxLKmfVezBacSD8+JovT24/63fcBfntt2FDrnxErImJEhWhofN6K4sb3C8
6UuCK9HQXiDiT1EDuZzziT59RHQ0/w2drd6e3mCmpEnKKBREh2gngLA39jgUQ0//
im3CYpSAgF5MKYCP/Z0Uw6+OJ5QTGh1eUdOpPp8WuEU1LD5jAzUozMMmWVnTaP4Y
7pvN37E0nR7THhR5VZ5xL7HL4HWGwpSboECOysPZqUl+GNWaZdZIyC7toWEkmJS8
ly+Qfz/2Vpwnwpsc1+BRinPOvFUMj4ZSWgsxP4/AHoOr2tpuzAc0EEiYawF2SCyM
o3QslbwVHQFp4OuFRqLRkJ0BhjM6UAiYyHDjf9hq1j0QKkrPv2z0v40BSDCQwu0t
MwEayyjYksk4rpouOUCn6UGEHG1N1vtKMCaD+/EEOTOjWZSd+828BiTKip6ywD3l
V84gKkM/ZL062IbjrEH3SfKbmqMkkyG199go98yLLXELTflku6/YKxr7xWIPve3C
6FwYFKrzWVcVvugdEXlrnRG/Uzcar31FaOL/dDVU2aw+8nX1NfcSJZQaCd4/hsZA
R+E94XGRrvBs+GnlJBe53FgK0xUoh6rJODsjYsLpOnNZ9lnUQH20gHmjAX8GpsjF
P5K0Svh/6cqfza0HBR9vs8e3A8QkUB6fwIZqAvex6Q7DxbYFNugXLMV0bz/lAGkh
tX4n7XzAv747QGO2AO0tleWli19o0eGGMIC8h24ifN3uECbNiCrIvH9nmG+gE80k
Pi6bRHBtSykqBmcOt1p+3oDVN0XUh9tIJggC4oeIjP11WU/yx3Ar/TCt4tdDue1u
//LC9e/V5MSRGO8kEG4hyLnfz9GJxYroDPszR4LS22zjMgeTsfLxo1kheIR3usJg
MJmYunu6ZT3wUtBp21XAE9ptW5l2Yk+HKgIbV/WP8Dt3T/o/ypaoQ/35YyGGZLHI
Ai11j+BYJ2Ir49t1CERyQxUQ3+4S5I6fP1ZRYF9zcrAqx/EE/l9ybps5Qj5cshpW
bgYMW6dEFwZoZKllhlXSUBC6tv8quSlJRPsVSCtfhKP+PPr8ENHVbIIYWwNFr6s5
kd1LJmlsMaxXAK8oXfDGzPaiEI/0jZD7DllW+eRET3sTwc9kngkJcZP5qiPQrsFI
E6dIYWq1cRz3+p0DmUVwrid2HqfcuYaJrYQDTk59gpdy3BOKqxqMXNRxKbcx9rzK
qC76zK30UF+gE45w1tXm4dKaPydEiSDOIDmeJ7/bXh4ddPSpNEzjO47ZWfX2z6B/
uOTeGuS4tuO8iWhX+rC1Zf6dy+INEf23vXFLrGI2LQQ1r7H29RatPsvna8nxO2yy
51BTwYFxsNzYkPaBR+EubB5fZK1pFLUIRrvOgR2QhLd45uvSpSaGgur6gZZ8+cG0
EKy6EFLYkSGKUx9skGKjA/Vtu8RnoO0PNIwblhAAHsGfpipxZTJLYNvHfG+MzcR/
oZ3FKMfLkmthzMTMQaURzB0VGmWI4bVXXMOVlm5paMzj/sCE2r/htSE6fOE4WXcZ
L9PnIKW1weo3uxSofHT3MrBnmU+z2mTq2eNt0aO6dd+v9bEiP8QA8p5oYL3JvfJz
PJ25xSGWheNuJg0KC7y1ESRDsqnGP8Iv/d6B2CG9+Z7wzb7HAl5U3aS6kTIlCUyG
SmMzXUiySu2lJJCPZlGknxqIwdyQoheKINeaOL4GoST31bNVFLcpmv6I+tKfNPtx
OEubWIlrPI64lOfrhPxkjxMbzUI+y9URL41OE79XQMcykHG1+UAhvuY2gUEAKFA4
AHnOfvKuzlOmDD7TSAt+wkyQXHqI4yflBG4sbqUpAkY5YZVCtzGXtKS1CJUBVJay
9si1VNGjAG8n+F4ldWh6oBD/0VhVCNOcDEX4EidY4L3pWeeIg9Yg6vxWdzxY+k2f
Pk3PRsx/Suox8iJiTv2NviRxpIJ2ZgLlpkBWmJTNvlwugqp/27o8uCqNjv5BsfMp
L89zFmHlGELmIc9MkFM80kDrbJx/Ak9rM+T4VVPqYUxuMeGZxiExpRblWzck5cbE
RsGE4Wyb4NtVm+ODQngkJJQaTQnhmvL4b90TzoA6TN8CUknWxdSXjyCsh3mmS/fE
/MyaoVZe/PEOi2jTfWkRF7kk0lUZyPTeboRT8s7+VNp99alImk2b96Uh2LspmO0c
BD95Cmxc/aC2ROv8QRJ7ty9nL5YUETlu6no8zeFzX/A3bZZxl7uUfr0gYtF6QkG4
wVYlSAVpF68fufuVAAiIzJunhtuuRxVuUhtkD0dx79H1hBexwUvuvvjpfYwcrRPl
kIMvmVgNDfKbyx/1xse7w4GqS0gU/ipZnrRm21cDkjcjbhR6cZdbFcDjq7P442Mf
MeNqKuI70RQepP9WaCgY7sJ7HgQfCWrnuTDWNqpKWYB7xm2UXvaL4SCOWaQjiNRZ
+aPAiVwjztubFuyogLbGNPh6fBRkqswaBqkpobfBEDbBLfSofWwTNI6Ojo/JB7nt
im+edYQn7+0v6XHhw8qd3Lls5x5KxEyo2zsOM2xOBsRNedzWNJ0Qo+37B/F7eMg8
nT+HG04/jXQ0j55R4GzKys4WwYkHg+5P226ifGFBw4mNVjB3NAvF6pk43zqFoja7
BcvEF6dMOnTXvRc7xMlmmKZaF0LonhFTenaFENWKa2B3NrefQSR13bEL1vtvjSH4
V71DoUR4xG16aWHpJfEL7yr5xt0J/OsMCvjtUXantyTaO59PVeL7ulTrGFHUVseq
7hNPijOgITyTazpyZT3WM51MXC9e5K62s4dXZ29L2TBIi1/bIOlsE1VQhnCmFBaT
gILVsIS/hpPSc0s9bY1Zoc0qpY8LC2t5zcNIx2RPho0OEjGV4r/3jsHWcAEhLq/L
sRCfkJ94eRYv7ahPtCGIWUjmlM6JZFv8hhStnZ4Z7IJqC2ogHABxM3jS/1sIV1z8
fg2BgiRhHzw5AJQmwPY7n2fCGWE7Snb8qlY5mz4Akx7gjqcQ5n1lev8HK5qV6Rym
W5ow9dfi9eOChZSkAVxwfqSBCAm22BRY3q57B3QeAF/UWw0vOO7O3c8ruVKyxLrQ
ke23x/QgYCX+eAdZzwI0QgpSGzIHMzEb/pyqgm8RHD3Kkwir0TlSBbIQAWQoDBOq
f3v+9mAH0SM2ct0AkHYuMU8iJ5onY08AUNpQ3lPzoYR6Od4Za8IaDSD35sB/Pdq4
3lD9kL4vMQw4lJssA6YEjcUT3Zan6PH6tWlKyzZU3x8kjzKQD207+C3kdujMNgb8
SvUIZDgINWH1nt3I5pE6g7e2VVtbyKrbPQuRLuPQxpnA1y45e6zLegg+XCu3n9J6
e4OoXdSEXnkROccjrI9vwIT2KzHUJRDROBv+LyWSAMfO9lMVkmuXhjH/kgQiZUnY
qHOhRn1VkR0ghDnLrLRuNXCPiPYo1InAwY7GfC8V2s/CW6ZlOqd8atYh9lo5MSWa
7FwPmPYva9+ya33aNSMEpO2jtPKaCT+mkHt6HJ/3Ccazhl9OtiSZG199ENwWLJZn
FfDAasd0whiD1NUDHF13T1W1H4JOOq+EB3dEXGs01vJG2RKxTODMH2zHwTyOSY6W
ctTxv8RqcGfKz4NAK1mL8lxQWRPghv+uiRuO5QFL7TZbTfoL5Qq+2dF75ggbcYbE
4PZtop1R4Sxb4tsmStrBJFlrr4nmGTkMbAZIDh3x1Bqm1Lby6TdcG4j/EKeDbYRP
kv7mqq64ktOv1d0macjPIg==
`protect END_PROTECTED
