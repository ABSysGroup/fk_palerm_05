`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iRIdox00GNxWAjTu0go1g7NeGsaHHll94grYB+iL/h1hoKarkOQ3YdFzwFVDae6U
Z2rTfLaudivamYIJ9UsffGmwOAvQtA6CO7ycAfET4+V2odf8ZRl2XPi5LxKe+UzA
mgs/EPSX68HwnzrNtK/9SM3KtszDDgA57rg2R6jG2jD81FHE5LxrOnPmBWdmL+fA
A2OrXHAIQNafQgK45nlpTnxt8p4oyqPCwyiUf0LaPJ3ZncNTJ+tboFIjchadFu8g
CxFfixFHcz90twVJOplPgw==
`protect END_PROTECTED
