`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iWe1947ioBMqPzkewSs4KDAjiBsSJfnf+v+6/HoSxn+GqfxN6IQtmvSxWdz7i5zw
1n0tbmI4poZkVN1KIzhkAYjTO/AyiFekFUZUIy53zaNB4H5x1c36VZvhlYYG9sti
ppEYFGJ6MpBFbHcnkQ6Y+1NjFNtlQEE9/IyjZEvD/8IgLklPNd3el2K2yAJr79ko
niqolJ2Jtq1lLGkPHlQt+EFf/wNdll//bWVssvznzIOrPBEX1BXtknxLvn51pnGS
x54ZUx41LKhk/eEzmPd0LYOi1lQQUCIukoZgLyJ2WCTz+ZF8C+KDt1EN3HqrxBqJ
TOXDze/D8xXoEb83etHT3nXzVMPo0Z5E7QDo5bhyBFP6GrLslOsW3DBQsimkeKCS
92xfWANRfF6GbG1z2BusXErRyAIQs7vvvfV6PxJ9QRw=
`protect END_PROTECTED
