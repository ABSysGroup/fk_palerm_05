`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wFRv2oH1Vv5RJyDmohekTa+yGhCooVTfmibkRmtemfdo2fVuf3ogt41bR9ura59P
4/UfJRDxetCDK4eE8dRbJhdv7ZIo1xM1gDl9pK7o4slUPHoYFviIWQ2WLYarnR7W
AsYUgZdue5mN0iCS5UanHw7q5d1uxHhT3B94fcsd7wwXFu8GeHvbKB/wsoGuqbSN
DPDQF8w0Ehso8SbQHgPEflFVzMcSmeTcVkVKYUz/dO/suOJRgtrQHQK/kYEKmmLA
3l6Pc4CJULRM5lL5svUdqVS079uaqr23nCjMkkoGxrZtUcK7py6JBEp0jKt1hqeM
V6pUwn8ZAizIEaM+kkRFX6Bm9kviUY2ZoMUJ1bZt4w/nIT1gTfYYO/4Kgjzb4E+P
rjOPGOV/0tfvyLFHZfRG8Ta6FY+faUIlXN4c94yhbKltWwb25vaQfKzcoPD7N/jV
S4aPrmByUHcLf17eKHOmQHRAzKDho182kapteFskP71iv7BMXig1Oum0wqYkWDc+
vBOh6zk4QQPZS/SHU21idgUximhmihwHNsz3H01WhNZhgtwHMIQfkuZZY8J8EK8a
Z/WBKXO5mSD4+Kzb6LqiliDDE5QrgRLqSZlRj1sI9K6wq9tLMMB9tndi/g9bKtWM
9oZekG3BKTDNtNrnkkbmPKghQxm0tN2Fg5GwHgVI3bFd9sm8oFMa3F4BSbj6UzIY
DxzSFjmclM3hMwHWYZpxhzPFVsTnXRVMQ33u6vpWNpztvd3F0dnzn2YMQtJg7g+v
0CmrTAt3KMBnme06iCflK03Ny9iJQmSLkAYmhcMvBXf3GhahIGg6TpKJlvPPcrE9
jxGMrdBWBQNk/XRlOJzumqK245zjYHMhYxxhWrbOXGRr4to3CvtOG/YS0HpIUh9s
HSJRJZ/+Kog5rnfvjzXR3cJ5dfhtAot3SgqY93WsgAub2AE35cbAABIdHnguS+X3
`protect END_PROTECTED
