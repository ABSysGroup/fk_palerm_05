`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
34qy5ZdxUd4WirPKfWpRiuZpOmu1hYB0vkU0bOmRsERbVJwiNn1vrKvhZCamgIuU
LftH4U+zIAjv3sx9SZW1qu7SO5Lm13vKXDVg4V0ZXTPo3s0RrGpkCdG/HazoF3MH
OnFDPGSzOZgom+DnnFZkc+p7fgegYNo8Ezo9yiG7war96uzYkDQ5TK7Sc1kBgL5v
tuS23aF1wy3OqhUpmqCE1xDY7vRsDlnsX/dpxZcGQp0dkUtKTi8bK2qphlNsJd6F
LB7C15Fdx9MvW1h8J4xAaw==
`protect END_PROTECTED
