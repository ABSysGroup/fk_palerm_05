`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BBtMxmX6xo/K05ecgD++UPSxP48RiSORiNDBPhVZGwvk1f2FCwBt9yh/oOtubdbf
g5LdWV8woiDeKt6pIpy0Tn+w2j7sReiUfOAA3FNFf5o5yo9qjRlF3RRFBeVzWN2t
HOw+MVdbh9oD2SY9il48WoVRULh7dB/cOAMPHNixQmRK/CqjGmM3fxPwfKSCvb4u
r7xD7dsvdVNcigKjzrQTvMYs6xDmyeXyZ0bBTRwJTLyiAP0l7LZXze95Vk8eW2iC
aZ8P7PT/Y3ClMmOQaR0t3RU99dUubBT95Rh7GXOtquv9YYi1fA0K+X16N8+ScWhQ
njGEqgCE87oub79iyiMMqYf0tqe1SsXbqNwd+KesIale9Q6LhZAJz7exUoYNNCYU
eIN7HTos2Ryky+DTiTC11EJOI9xtBck0LK0lu6ZDG86duh23QFHJILZ+IwanB1Iv
yMhcmy31mRaxO7taxhZqYayFswWHr/ljagym51QFfK1F0kn8GHObei8g9kkFof3i
OG6wEvaK5rjBgi3joqj+xPk8Ou2Ktg+0dfRekiTChw7tw/5zxUenXyOpjqJei63N
o02y/QGFCvpC9S2CXk7PvzM8WDlJLAIlPvTxkjwmMpANxNlZBvsuV2mNdt1+2cmb
Q7rLHwCoyekiUJjaQO5Lz5UasDnVsY8Fz3aUG3r8Yebdjvl+1roxiUbeZO6lZ5Yj
YqdYzRZ1xu6mfitTsoPAPav8k2ZYIxjCRkmnyPPyTBHS0CTwnM2erBunLMThRrdI
21bUla67hzmkbOep88DcVpet7bMbBg9cRQszLoWm5rX9vYfet2FfsgXz59ih3f9l
MI4OV8AAXUwiwyBYR60I31X619XxZj7a5qu3Mh8zwQWn+VCZYZ0B3rbwEQxRSZF5
WnaUf5j8Hbqz05AyfakPhCLu4lzXo+Y2BZ34kKfKT04JS59R150+Yu6gOcqY1yGw
`protect END_PROTECTED
