`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EHrzJAh9w4DErzvncFRjy7M42bFTGCt7SB51mN6feYnB0orLEPXrk/Z9RZZRKtId
2V+5t3EQ8dRP8OG/UwIQwiGfmA+f0Sk3rlZK8ZuqPoMeN0Q/8BD6JLzOGEYWU43H
euWIDwIXbDskxybToNXpgzqbWn5vws4Xc4OlIy5P9YZGT36HJPGQmkZpbYdwj2yy
jRtnfTQKkjHJhMn+9DhQQC9glrHaoeSh+e3utogr92OgXq7LfTxeCqqhzVlpxOWs
kioAbjuWdkrweu56c01ifcl3zlfdMGb0vI5qWCqi8y0+pCw3meKbSUF0If66vPxZ
ack5/O2XtIP1QqwM6QzwnMHnnH2SN5cydUdu4935fKhPIeQ/OYOpFe3oKZE5gQv1
/t4EfK0APSh0VxsvEB0ZvAeDuKflWHJ6ZlQ5pe+cjzieP3KuXwN/eUPeB1D4YX3A
f/L4gfduc+lY+30Sd9PC31AE7FUnncBEsLgJNkd5SFNxNNNSU81hT0ToMomoI4gR
VZA/F7BpNsTNvsRiRQrqZBMXnDmgV84KCCXQ2/hVoSgUQw/Q/dQrd2Vi+B3wRygQ
TkHoeB+x6/pxB0AZCdJ1UTsuZsQIixFKKPZ9fVYbDMtxdq0IZes17wlr8swe2+EW
fDGTOnXIN9dbTdniV31AJtseAsnBkoaI1Mm66CmTKNJ2g29FhmfIR3AvSt3jaT/W
xYsac2H0rEIzyingvL5VoZHlc6TbdAzIyvJcoX2WFbWvmCEq2JyZB6K2hr2Hk+K7
tjJ5MbhZnVPCyhCD218Ibum26dJE/DyuvfMy4UtJOiCWtLBAueWbgYwE3R34MroX
6O+fB7rji685TcwJ/mxgmpULfgdvMbwOEhB0SMg7yTTUYJk7IgIjtXo8OTKiEmNR
Z8h2yQapsIi0k5HPbcxo7wiG+0/alEtAN6utmtth4RcRxNQvxNJgXkdLmbAT8x1Y
NgSnVQb+PM1CjGSc7h327yFyPl0YsAx1xZJEAvw86o40Fx7+H7OhMwhG5wIUJnjs
kFs6J3FXJAzRFNc69kq2XtojNZE20AijCU/Ah5ww4SGc24lof1V5T3fP3jK62OSf
syMegiKvV3QBXSPPucSi1SLV3nvf0zqBILpSPLjK2S3vvQsbEmgrICPFZM1qJpDB
`protect END_PROTECTED
