`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lifuwE5iJvlsCqGEaxJwx6pJDjeRs/nRVfs3ULLHlAeIFe38zKviHYfSAfLWssNu
8gGU43FbR4Ej+o91oXg8b7MUtuetFYcqbZbxTq+DiOHQxLLH06hRimcCD+Z/kX+o
gJe4nmecBQ+VJuadhELzTE2f6yVqiItUniHSVILrUJPsb9/CV7hopL4Mj4xxgnOP
X1ib8m2pJRmiQMBELGjiQdifcJ5Yh8y/K83y7fcsQ/JId7oBPkO4taD1RTvXxAQl
wRd5lJvaQ778QCfrfiE9pNRiYNZ+LZUtuQDcrVBipoRkusnYxKyg2LwUa/9bv+on
HOVIibklRA28nm6FR1sRuw==
`protect END_PROTECTED
