`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DUqXJtphwVvdQ4ywdzIdbkBBQwbq/fUtkCI8czbsE0DF7AuhfTyudMfwKzm1DTGt
HcuU26BjG73JlYJS6/IyTMC1ixhHjixI+EE/CgtAsBrogzCwb7dl8UiaR3F5MzWE
pcCLK4X/aeR5k0M0OukjE2h0kkgMre6ipjb+YQdDJS7trgoPApweDFpPAOSTHC5P
+m6HFmdna123/YdGHMvuhY4OU9uG30IyrKKjzwdlEXdZKesLG/DAUqUbe8I3DZ1+
Q/edy1retQLZPVayuoN1pBYc2U3t3eyFaFp6L/gbgXlGQDSPO9V+xn6fvuRrHCqm
fGKv+2jLGO3aE7orlbzHgCXKJNpxQ7/wNU4pVIm+f47dKEoiLnSwsZtncRAmaKfr
fboWuK9rga1671L5ZMqut+cwdChzF6NJGGRW2jPZzPi51r/do4cmWLh5e0VFBWAd
9bOa1DrpPZHuPkxXl9Ce9BtUDGehyT+dVuxjhmVNG26HsI1h5v20PnIf68WFFVDu
Tq9soOFZ2OxzmlO80G8b+CGiZ+ZxXy9oDtBiTXHT3sdnOSlaQ3v0DWnZWNXFYNRE
3ughC722NEyZGPj8fDYcLNzyTFSzP73ovEGb10Ee6qw=
`protect END_PROTECTED
