`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iW4ykHeCzrQv1YPJQYVkQjA0XKFiBpojtk+CsuXxPFLryS8Aytj3nJ2VszyF1X4B
x19Eqs/vmWTUbuCzz6KTg+6GPWUdU4zv6b4Mav5Cppa6UXWKXxlyXkvY/1o3KIME
SmVeCRNTohoRE5UWc616nrT3OyAtXp8PVAZeMM85SJkFXBccKzsaDA8wCwaLdsqP
/4QfbYJf7gzYJge3//fYtWBIsmJ14cWfwCtXz3n6VigqZSjCyc4iLzy16yjaJN5i
t80jwWou/M0xpLx2oZW85OJyqm3rA9w1pkdnL9zy0DX7amBEYG2j+vhgt3n11Lom
ax7/bQkFHUeWyG4laj9TeWMRzGnU4KZSPIZpRmWqBZpkdfmG+9V2HLbQN7oJLix5
WfN/cAxMbIo5gdc9GUXMtKydvsY3r0ZmHHmN4n61T0Y=
`protect END_PROTECTED
