`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OPrSBCB2JYYA0HuJTMffH6Y8Z6rPPfSN06DAMAI2ST+jzcrl2vBEfw6NUDDQy1eN
de/ZituEbONSqPyajJeXQIcKjUahi/aLLOC4XzKgdR4d83lzREJJb4DUhAClqSwy
MCHI+MCAoVwxj5oOUOrXVXK5AGcPqa8tRYnjlJ1PFmJnfJgAaeP6sDr/0zngsMTb
VgfTuSfr5qBf/sc7MhjeBdowvqrgebcxhEEe9tvu57w6L72zVDrXD1SAFkOGvcUd
yjUR+rxezbDi1kH1mHHQsFur2L/ECS4FOJ1Ny7OvuxEVxAE0ttx1SkcCnWw/a7BD
YI7+gPN4lFIdnsQjV82KEa/BfoLEUmgr0qiwzEmwOvG7M/IWkyP6sCLzHjT5dB4i
jg7RWqrIJXfqFxIhq8tCqfSgo5bBKIwHDFwGPHStM3rC9cVfhluJa0HyuhMhPdQ4
`protect END_PROTECTED
