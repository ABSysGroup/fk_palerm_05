`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6EYsJSLJFCgD75byaUNLSlZmwxpE8guEPcy5ulSqKczKf4TCra6/pqz3BRKsjNA1
/eGSyLGv450LbD8ApLmQxCFB5XSEiZRQj7rQgY4pXHxEekp38QwAJ+2OCDkgn70L
ifZD3scGkLy9P2QiplFm+oK5bDQ8oguxER/DImC5CW0jwVVOtYnVoB4KqwTcUqig
BltczBfBHzJFzsghJ6Gx9gCf2HdgOzS8CZmQ/K2hwn+4r4nL8dxVceFoR9LI8JZk
PqcOBHH9rHIwDTQHYmm34RasE74Zj+JoFmFKqT64nYSyIqAi18znHVydc328hamG
PmwULtqO+rLQeW9XWHkPQ4PM/uN9N08PThGA5m2xDD/qeAs7YigmQ570z3pqeh+j
rbp7Hv/Qr4ZwP6peSz7S4bqiDeNL9i8qN9y0CyiVDrWzE5KwTAIoyyupoRdcRxa5
TYzmmxtzAGeh71clgHrzXJTmCXUM4BLDOhZ9Zz3xKKLEZcp+3Qmg+0UCPfcUCQOa
`protect END_PROTECTED
