`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R69xfsxZnCDS1CxhecIN8O0DoP1NgjXT4jbAzhy9fgqulyIY/EglOyHH8gKeUm6o
dk2dD7+v7HcUdptIqMVtHqVqYy5dHWPw/MjlRBUUQKSc6ExFJ+gHywf1sQRY1t7K
cOHRi1gAPTFLkuu2v5/nLcm/VBB15q7LQoaRvPJ71CT1In6YJqEcYQUVukzYawWM
ZnWvApmQcHDcDmiPE9AS4ISMMHIOLZSMhArudZLe0DwB/pX+HCpxudjsJAOW/FRP
9xDeMFxL/b/0iD8rpyTlxXChpp44xCWUFTmhEHLdLgJE0daL+SpF/VqsOh2r35Ea
syIjgzmAWesBs8A3pThhEQevfqWtNa3+ef2nR5zDCnvkIpUfzyPK7yyBf1V046H2
i3d+W9oZ4ccU2jKQrg99FZBiTHvzycffyFhWpTleHVsCCSLjE8OpDEG0ibHweqEY
eF7wW0REia66JJunmxgZmaDfShNcaXYeUkoBlHZY/ZvO+kv14oqd8pQj0RR9+DP2
ftH99wpyxBOHPDKy+eY+5426/F9IlJVIZQUWvKn5m5FsDhw9gc8N6rtRh75C28zz
4J17e+rIfqxg5pas0TRIAWZtWt22IhubNAzm6K9RWqX+qOZqwJhEGy6qxrt7EG8v
UkjnwfyJijporRp4AfCjMSIi9rvyUmDs0eYjiBnLbEZ5Wojry8I9neGpMnz3nhYz
XyJzGVzLpXIrdXvg+yuXpFyzJ+yAumoun7y83Wt2s6tq1STnjN7fXphm5w+AnU1y
NyLESGjgtO02nkMyMKVYdX1fcyd2T+lLTrsN9hVf3zOI+le8SOiK/Iktt7jEoq6V
No0ebXP5WiGbbB4BrQZpaw==
`protect END_PROTECTED
