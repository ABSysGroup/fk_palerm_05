`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+O3NrH+JQ4aIWGu74LAqefBgpluYNzQ+9bGGp+jHW0qoQJCZoWGuqEN6ocRHnoio
oWGWjsAZE7J1XDCLTrhObYjekyUMVLz03nOyustrBn2lkTQOrippDUw+/16QP3go
Qs9bK3tltOM++fyoPlMjf0unZT/tA/i7yLFRB9Rc7H20sNHdRG+dSKFGw2zDKzFH
hAhdg6L0tBmdUMKlebXDX/D0OJ9bjpjW4wFGVdqvkbCX2dEIZzMRozfy6RlokP6i
m828LgTgWP05YZVW3B4LJw==
`protect END_PROTECTED
