`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XfK9urqdNBBLwb1U0bLHgi7gFrs3wjlbeoT+uQSm1N18mljdx0pbk+CeaE8tTnMz
Bsowg3wXGRuiy5xU3TAKSyW+pTTfH6GDSnmjl9NCf8a7EWH/femMXKxgho/6K5m9
voeBGivEukF/SkVfyvHKvsYzU9JN8AUuFEKZ09knFjcTRZV2t3AgrEaEMo/OuaQg
ph+61CGxhiNUVGT10xFiBBjwyq9XrxdROH6xp89IoLLk7JzjynMQaJrDJB32XQip
AGIKrkUxtHUodjDX6N2XGOPpJRjSVvbu7JXkEOw1MpFhSlx/LHMxD681wirFHr0G
j1ZDZSV5iLo6whm82jGQoQ==
`protect END_PROTECTED
