`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aQIjzzmdsy4/D+csRo12YJbFma+HYiZ3mt3KsdUYwQxhefT4K7ZVQQ015M3Le4qS
ixa+HVSFdRquoz1sjkRhzAuUGyk6xginToPYEm+grBqeVdc7D19wNauYmjZS0hLX
HyLqm7rz42ku7MkysEH7WzABE/J6yAZHV36OpFaSMnP4bCun46E6+KLCYlsuTOJa
A5CnUwEIh6wjPRrnJs8hvW6HBNlvEr8811wLPGJ1q06B2fNAu0vpqfqn6EYFk40L
iHRvcCl9kyd42VO4qV39FQyTs+j9o4WVo4tyfJ2jipjEBaRfIZws3d5JlEmMGhHH
Th4xPDlAXbu1/boF2bfI1/eH3lKnWwraHeGByxR1BwwoyX7sPZEiqQQ1A1oDL82+
BkPAkvExXbi21f23Fgm3pJOQDrdyu0W10jUb0IaXNw4LBCYsl7L9xBOJpTidrvJa
mZqR7/+AowWCy/+AaVHLqDFd+n0APscdbR2Y8R7Zk1BxAGt7ccBNoYIXOEWbWl3B
xrRQMqcoN4HxMtuFFxtQjaOhP7momm7IkMhM8tkYypzmSt3ek31oiRt7KR0LbJ16
3//PNwblF1GM9nHSl2rdSzaoBJydpX7M7WkP0FSDwHee3Vuh9btiYAzbFWI5MPBU
PTqOTiH3MDUaDB8URIIBfw==
`protect END_PROTECTED
