`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jteYp0hKy+Byv7x8jEilvlv1rztVB0wOFDVw1qv15+OHTbrQnk46gP8yVni9xkv0
uUi7DsxcxQW1CJlOfBIC7EeKzkACdC+ATakfT9xE4oaTv02Y0CEY6ZhprvBy+sLj
23NVrv2W4HcQYh6qBkqhfD4V6MieEdBK2zoC7WpjtAQdJYFHCFaOB0noaW4devLI
fBuX2NM4C1qOQAPTwXelw89PwJxRLZbk2AJpYL5Dh774wiJxSiMGXmKv1Nzag0ri
Wmk22TtRLpF9adukc8EyGl8cKhe2VovIcW5TCku9GzZgVqs0VBj73NDyTrapvZpP
zdaKIhvgaOZmEadhuZoAMS2QL7fxUDQVak4Kmh1y84UntpXJto8j6nX+L1ePOX4n
KaxVMdskYjJkQTghDRn4csAWE/yA6w9S2AiZZl00TUoXr0bLqbsgwRZ08cBBIeOu
cV1qFS2hgp96keaDBDdcrPpYA7suFM4BmbuR6EB1egAXcgtrHNZooPIYYgahm7Yc
ZcY/32yfX4Vfvgdl/eTuJ23Rq3Sag9n2Zs+2ULGdkmBUSzzzupUMJ65RhQjDRc0b
woe58LBWXcNdHjW4uxA2sywgf1/QiXeCxPYn3ZqKTkp45rTguMCHpI8fmqvP7UnB
IbrHC+s1zFow7G5baPztzSrpGpwUHFFl/sYt6ZNIH2HoNpR6eQE+QH6ujYWPd/ZD
mgs8PSrlPLWIrIEzxeD5jpYRA/c3+HLCoRVJ+7pABrf1iBQZXIvDXAJzgR2WbBz0
`protect END_PROTECTED
