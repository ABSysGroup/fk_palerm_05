`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DHnJZEXUs57Rd/gOisk8tYTblco3ywcpb44kfUdXKceDT6FOj0vFJyNwjlB1x8nW
yuBX29q7l0ClufgnsA8whGJ2wnbxtqdo+gzCnFkAO3cCR8ZdMhI/fX2wyzxT+lcR
Hyx4I0IvtW+DMOYL34zZYvivX0l0w1HpsPUNsVEenjKJgbnKuy8k+qiirGzWvOTE
EFOpeiMUGZyIAKW/Y42JAHpASjWP/H42kcyRuoT4xNgqlfesSPlkRoubJtuB975J
/0wgQ4WBgHwFz06Nt/88m4LaNEu5ekLSYkvPf40FXkvixXoAaLIUx3gYXNMB2wDG
ESGiTyPY9ojxCASeMyr13cRuFqntBDWgcMxey+oOLbcGa1LZ6FvlntnyOZk9Z65s
AxgaDEteE5pS6uwpf5nOZ8Mb/VL27FxSMYoDLPP9w1Wm9nHPsVys2RuLIlfXomF5
`protect END_PROTECTED
