`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5NhGIQPg7I+uHR9LyrKl4AxGi2hXgWAuE7zKUH7uOdD8AB4MW19++MySQALseFCu
e1GCF54/wIylfsSve0pg6g9lHQCdMB4PGn7vRF6ep7ovoeyr+TD0nba3/kDBtWUk
1z+vgK2+ZL9q2BoA32iY/M0zJVZvMGBm+ezgjEAOfIt4k0R43F6zYpTvEH/c54VS
L/PTjThaAHiYXICSGW+TdylECG44hFqOQ7r7eMmD086rRImmmoFy26XH3Vviuzb4
DGyFle2HQVorVMLcAV1nnhS5xPNRT8fFAfgWibv/j3ONN04M9cxz/uSgnUbGs2o8
8pjqGY/H1n1CdF9BSM8V83PhUNavjriHpxWK0GAMDkryqB0Dg6m8DBNaNshuycva
T7PrQ5EQxA1mvrJ+5oib+c8KUgUackvdxqifTyoI4Tk=
`protect END_PROTECTED
