`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UahXFtOPfEcxD1Ud2osQt9NwHjZlydq4p4QbL/tdNJGq4PVNB1+G7KOLVmrxgF+a
SQdK8FE5VLNKhL1z4XPXa2SG9e+04VQ6tedBEOPx4rzPGdg5gdYRCNzBgaAM190x
iZK3WbmFzVxFM8G7llQQn6XQGfIJGT46ESQsz3tNtfpod95qtJ4gIDMgdJ+lheE+
IMa1UfFMPI4fQDUzdL9N6nLQ6nxxQ+6TToG0QmYgRz6vzbwnFOa/PUCX72Vez1LS
on+Popa/OEi86iJcU1WCrlfGatGyv38jIe0EeTOjsF7c28HtUC+Z55CuzzVl6MEa
e0lQ9JCx9EAEsMdNsnF5Rg==
`protect END_PROTECTED
