`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kjW9KSC4Gsj2aRi+0Q7ezf/nm8Gmlmps9wu7wtS9dXV2kOWMPx2RYt6IgbICHuTV
YZVm1/dmwA7ZGly56Yx+sPFM/kxBqV3/8+aykIx3juFDfzXBhG0vkyUHxecS6YLe
ad/5ehIKcJSMnFbgEB/Mtuy4ITftIDgZRrZpzmGqSHJCCuPimBOOp3rmp3cN/aT+
ueELjuZZVBWHmmmFppFy66FqgX7cRZn3N1BwPhBmYJQY4HcoZdoPSHb9hzAUX/go
B1QNCDUESFUwaHiO3U2P5HMNO0wehqHZiZNhZ5y/itoSnE17RyvAQkMXGxpdM10Q
sA0lkk9+xE2jYfcm0owDoDh8se9MROIBhSw0w5k/P/ShQZbDwrYKeFgbzvth4QoA
NUGdfZhRkV1EbTPs9ZnNyWB4ZkIbFelcBpH1zX6BuXPRiNmawuHTFQMp/IlT3Rgz
9Zzh0tzmjYUjP4VfrsnBhlUCd5mo0JFp8/U6Xc3FAwoHwq15iRLXwsz1fkd8aTS2
AhAnU4oeOQ2EM4GSVD5G0Qt/PmZLqo4EDnbgXz2bW8JIliyiqHr76S+JC451VGze
GE8g7PgJdSqln7vt/mKVaJU9XAaH4Dlua8WpzisfUS3gY6tYPojOgiRiNoKbWXKx
TGLnHvSuT56REds9+rVrSbRRqiZMZFXeBTsiidjkmaCBa4aDKsd/VFxzYJxLYk0d
ctX1MnAhvpeuYU1CGOJJUUkkq+XYQ+yG+Y5Yml3JdSf8hkJziRtQC1TyvjQ/hQE3
GO9qQ5oQpas8xXB921IBFZwD+JUd7BK3x6ONazzlmEVl5jXwfLJ0McZQuQC2gJfT
SpK9iVVkGrL7uKvvUvymtznia9aqbHWuJ2DIcbmWSy4W+4JzXb81v8BPWYmzqioy
aX9edei3fdn9UHmYXOlwm9MfpKoAgN2z438hdfnY280/pVfBio3d9NNnHpmSVwtd
8Hk+whY/OHPidFEqNYp0yS4wFLi0kLZKxWmmAYY96pHXkFKPh0DXQpkGCIQX/D16
k9Bwy+X7o3kJfBKCFJdTMO6Lkgobmxl3BE3AUlNLwzwjtYjTXbZIfcib+1r3ONdq
tnqlYYZ2ESo9aXB4JGviaFpevOS5aVChNBbAEEtTLVIVV4CGHjmhMQ3PDC8YS0Ea
9ZJTcU7mPwoXhe5NVnOI2cjp5c8IVMgjTPJ75HU0wHF1w2zR4XRQ1C60Y/yU6rV5
4Z0pzyUa3JRF9HNZltQSXUzWmHlJxyrS7tuhR7v5Yd9HPNh7Lf1ZC/h4ITRark5L
6VnBSDlycMjEkO7aclrdKJv4yXyw2JcbAC6a4lassUUlLpCFmksQHuXpIHS3xAIi
Er7kNGsYmS4B0Tb8ytFMaZlKyVmM0tscc7oyYCy2IFpYdKeslds7Is5m2uuktmvY
50aQIlfYwdDE7UaUy01powzpTFsOO31aFqMWwVC+IbNYS/ZYZ3rQO12bA0PMkVfX
6dux9IM/W6ZotpBWWysJIWX9QgxaUh/SA+KII6FAUL01QFApqTqaVwhyKIob1VHS
ieMdesa0uW1epRyfqFuEXJpjmowz5UtxONm1tIZQ0dnwrKX/zaloKWPUt8RsmfSU
halcdb5EgMJ81XyiTihdwmr+DGH9++0iB5BhHxd43lm2LadKZbj1uMZJN3lSpdbP
29DYpbK5Ke7TSUeaW/rj6Ctd2ESoS3mwAJfh8HWshgrHPmHm7+Lrb5Aaa3W2n52Q
hEzDlkxSyrqOSHHtoocbHRkZrXFCdm0iS7rSzHoq7yr2968KK6nUTcPiSZjzLwiD
RGNhigJFjwMGaCDVaGouxU6mvVcUcVeqWwKrDozFphjCvtbvwaeQD+DlKcYOInTY
b2SosCPj3izl+77/Qeimh8KhfzQrzV6raUNRnFzyTQsQMnpLCpN6dIsQKNgOccg4
NdZTxEo3Byndjzhmzv8rAc6yB8nCP/TvMT2F9/bV1/JtBbDTSVdy5B0ELED2O+7W
NydXHJRwHbYWAuPInaSqa2/Ql8sH10FJGymwppP32yTwpUFmKsIkFWUwFV8ZoyEa
VtqwIEMJmpml9+GJw11BoOSrCSYdXxRvWPeZzugOoESovCCS7NsiYajQqh7lR6QR
WKro9/0YNIuA8PFwTWcdKG2r4n8IdwuyA1xw5wBjKYyZ0ZIWVyPRZJgxa/x68H4L
z5gnwG0deyTXqk43eFa3NVJkl2dlhrw+P0KsRWciEl6t0TAgNLGFIcBRwNIteB96
Gq+f3ujfPKldEX+lZW/cRrHPsqM6pf96iBVnc8q7LZCMbZZY6dNOzmaXwsGa1BKj
EfLz/HQM8uYRGbKjD8JsxSvaxnjTsF/5jBn+dS791KLav41xcp5rfBESUAKL0ejT
sPH4MjFCukyG0tGqLj05aGOY4j9K7XAa2xGelOlv67cLdQM8zfViMP3ow8ymggxv
qCRV9vVVhLyGB7f1dE5H2QvON5VsdEVe9bHyA0styn09CVolDkU7mgF4xHuGqS8k
Jzql+J0g//SwRm+IW1IUfdNx8IEngZQLa14MWu4QsdgyW2YyEK4LSx2b17kHvSF1
FaX8zA4hOn3ZSCv+mq4WlHw8fuisErAdoSC9HPufFMNexWsbvJRo//Ip8ggJP7AH
bJf6SklePViEGk0ESPwon3hlakbT8lu3jL56QioLgDBshQXVYwyRZzwNTrrr9lg5
zzCb+MJmXBta3Fha4Sm/R/ftn2JGb8I87VfaQtUA5VHyPg0lEvRr9Af70VBfRVJs
b20JnlTVWqoxw8h0DEhhuCJN1IPh2Yg9tD28BjHI1ccXtF5GmZu5uQlYhmXxiCoZ
H3V4/Pltx2nKwpyzaS0yX+Y6B9ZgfjNg+WZYgj1E17IlDKv6VgFrvyzBl/0gpgZ+
6GCVunfTU+m8xlL40Ir5toJy53wRodhZHtGwhg+/VPeG6k8RzBNli3qgYpFJovdN
FEGVyGOCXG1bO9en8lpQ0u5+WmHUHQfZ0OTrHP1Ub93ZHE2l/H0349wu5DGInAeP
KyvY/h6lxQV66ZPxpcrFG/QfvVLj4ZI9w0DGG6+slEBca3U/YKrmLn7cXEZ9ccN0
4SGsRldyzPTA2rnKCbLQvEkTcJiv6Cp6B4hbOcVLV/fWKXBCe+zz97ods6P5qL9I
oEGzQfS882qHITynx/OngSaLg7+zBZhu6x52ol0PrBXRnDzVenO9OwC8UGw8n6Um
vElhtpiPV5FvoOoql2z7x/kYWKeDH2ZqpNqC54SjmqWwMo1lJtJoCg2G6CDRvizZ
nZFYGkluNMi84rJhmtvPL9x9SJ14EHriIFiCjygnukea7Hy1hxG9wEE1c7V6QkEr
N5wQJn/Fqvs0bMucDjuAAmfurar7cuKbGhGOx2iTF941kIf1k0KhhV1Dnr/JhE0L
zCHXKy2wU+w/W6NereEqYfF6L3Q97XZ7do4s5QB/0S9LNFf1V87nrWCHbaHd3Xom
10D69tpFTXwA8Q+9HmJ+m1ZnXRLdciqdXzvQvCBWsRnAfwGTbwsXDbM+QhZmHbVA
cUvTNkBvZcVPMrrIVPNoqyQTv6/yvmWlnnS54sAiOH1sIDNwckvO1L+gTjEYMszH
2aqDLI1IX0b8QXVmoqKXvNGussdLHKg6qiFvg3RtEyRCUXuW3PPnZpSUX88PIRLt
Oun8VPfkJWupy6Emy3wB4B5eBB/D7itXBfJ8aj5ZBASHiZhKGDr2/EO2v+Cd8XFn
CCEO2ZAM0Jxch9y2uMnp8YYx2UYyThPxf05m1+OigaKiDIviLBqnkzbBNrsDR/ug
glKnFD4tuscXhZfwvz5sWPkDv7aGhpsnAxQnpW1tNWf+zFMsWKAcBV1DKshXfbJs
KOgsylCwEBmCP7TyY3c28AWCgdFiINCHsLnMXaDnUuZqd1S5nW7sSACrCgOnPPgI
xCTGHkpUhCIaDfD8qNdntR71JY9rFccOVIB8CGP+mt25E4uUxdFitadOM+p0SYpW
406l3pZzVl2sI1jR9Jn6bohFp0aeWtYbayJzuTa3t/xePpXajkgB0P48iTFurfKj
8E5hE0EObBubPWRVXdSlbZbcwrRoUZ4mpR39jt5EgEigVFu7gDHqHzBiMSjGCygb
mRaPstJJQeDccIAbLT/+6Ocqjol78RT87WlZQwTuxI1hLnv3HadqpG1ypJvQ9XJp
+lXIbxNVqQouXvSO0W3vRlVFffOP/XQlasfLFQmdq3lAm0sgcvfB1cNYmYFaYek0
oL6vDy4sWb/DyT/C4fpw5KaNwjYeiTBgXq7yaOwhlbH0XuEFaUoVcLPReuHank0A
u6i/xqrwVlyVOrJSonqiedWwy4En2AfUAEfo6lIr0Jrc2YMZp2iJNendwOKJ+G1R
0H07Oe5G1ZtVX6VmLwFJjnCUO/imzFhRlBujPATqOt4M6L/jmEisY1Abl10FlT0T
XWr5LtNVV1fiKf8FsXxRxA02SOjKDLbtKwiWZBfD0dX1nK/CkAl4h7lDFH42U4w8
0YRE1odniNkqfDy8tUGLWPJlTY3MD8/aWFZH2n6ZyWS83EB1INYWXOw0p3ySJPcz
R8d0geeAwsU82WMlFB5tOe6hT8BSwMoft7VEbGJ1CN4vEFDBYtDAcFdgGt+VMWa7
zdd9TS4JhOsoSkiWd4a9FUjwUGgZBsAhMafKM83QIECaXCfL4BIIHagfu1jPdZ9v
kFkho7p+Hb/913/qILBfDL1PS9CF+VfA8oTXZBqcoZSHnft+hBxtcWFNeaL6s5qg
+2Dhlp16r3lUDDMYuetCaX6HAKfw82P1aCEoFIO3cqbu1VrqGpI1lHFtK7PI35Ke
1B16KrLWNYgMkAd3T36k8ehLCBZa7zQZpH13FvhZT/rFKRCEbdy2zU5JIkrr81jK
H9I0YUBm47hwqPC64QDn92SzrpS6sohH3ozCBDxbL67rHZIvx8gmyOyMI8ja/kDV
8LlVwe/MuVDyndlBflW+VT2tzK6vuaMzl+mkm35P1BSk0klIlzqoFTolXZkcozmC
GLrZkAbPFc8OxmqKK7do8EHO99HK7xVwkJcdJxM2XMKVG2EYPARWMGrhIgz7q0nA
MfAzrrdkSwQ3XvEHuRoigQWVfVp9X1ddCElGYAFrKKAE//rYBfoquWJRcV9ncm6R
6tRquPKWgYQLc7Fx/kxAWGtJ0TJw6RgwJOEXN5+VOHXrggz9olAE8TqBPtG6RW3J
Y7rvox+TPerO/LEh7W5PlTb0RQhHOc6vURg/92orByxi/OgAQNKkMmJ+Hbu4S3tQ
zTSRLRDBv7a6SV85WEnalj4N9pI5TIiaje9jknpGwbswfrYvQ1TwDuI2DgLhLlYq
p/PElOY/43fK53OLddsqWI2Qg+rH+KHPCKFMRFK04Ql7lXA9ch851TTlMibHBvOb
GCZBb8x7zju65qdYcQZome1QQfofxVL1VGw27Am/zczB8MdfeyZznEZz6MWK2m+X
VA7kiPg9mrXfpbTsXnTsBNXQUDzez6jpyEaObuSrapNdctQCmVQ28lmSNYjV6I4z
mQHEqWfjAFHNlmo5p5LtkLl+b+VWNYv3bGfElkUvXk+4vLhWqaHDpPsN08aNvZK6
24Wvgx9j9znKyPPS4lu/tuRD/oLzYt4NBDxmgFpns0SLlxlkgfcwcVdM9Lkkx1m0
oN/Dwd46wbMv8C4OC+UxY/zAzfzsTVYR+VqC/B1Q8ihBnpJb+jZ4xiRusio2zJWU
C10fhj0n+I7sj3uNTC0BN6HWKOSsQ+Cj8jjbWbUmraE9EqFAYcaBezZGaA/KMCZL
BOo3vmnPrQncbRcEbd4Zr4uCYd1US2lcoBbFMBC9OAI4J+VJR78ossTUBmp+ruPV
jgPecNrGLWGds7J7LzHRCUHLxoeCH1aVUUu2hTSU5d1slvh8M4b9dRKqAyvi6RBY
XTt0rmlx6k/OjSpli0xHR7GiD6Rbx+j+G+yTNpRCp0r2wY5fy4bXglDleQOnpUej
Sjek4ijjLKlqMvD460HvPNLeR40hURgveRdhTcHQA12eXh9OJHKeeLMXH0MvXbu0
7JBlx7XAmdHgh6UHISNBulERZ5Vcfa3Q9MV9pbqtHId+BrjHWMY3vyAwwziZ1hx0
a8H7ZkzsGJ/7xKjBgrvdTJ59M+uZ+1zk3skm3q/7UjaJAPYaNvY6BJcMAJDlPhhC
byOAL+y53ynY9cs2CMbFrmeuWAYgHxZL7Z7SyaHLabwrK/7PJnysbADS84UD1sg1
7fbAtcYUfhZnlW18AVX0Dt6Tuf/mYxBc5GPathjB9k+bGaq0V9vplOcNfOh4AT9k
axEEILrhxjbwtsu1LfX3MQGazxw1bGRbuJ67/IIB75hzJ4Ks/b43aNbdNC5jIPdz
DwLL/WQb/gioP/7gMcR4gg6BoVohFSWwdt7RF/NQBLs6TiwAiyAcR/kPzX0Gyv7c
MULLWCcHANnqNuXGJyVxAfCUEc7IfWaUEF8eWhRlOmAUXxnNulyaH6QNmV6m3wQk
JfHEVVapuKaC1lSAAr6qsqmpWztDycAhPAheRZc/nNszP4fY7Yzd5h4NAQpmMrJK
bnYVDAnJEsG3rDqCK1cEVbz7/HyjmE6rWlgdN/ymKrCNl41wR/H15VnVhIWleZyl
6ZPkHOjVlrj86ZIgaIMv+pC19whs1ZN2gt/K4T9bjP0+PKoGMTcHiw2+1E28rqoz
KEm/j3Q1TSgJu8AElkpwrajbwrjKL/5PeeOqF6U3KNM8he4tADJpMYd7gLDdeloe
jAjEjtfc6vLi6y/q6JCChxeAICZ6mrxtow15XjRMpBSFabIUVrjQWYOeBKiuOai6
AeWAPr1xxUmlyWss+XLM7pYrRHx5nTBGZpuScbzWkkfY3R+VEKZOiJ9523mOgipC
FQifG+j0JRqj4BA4ewUWljJN5v2CBl6JXwr+vZB+G1+S05oIoFgJtDaiqAk8a8x1
Q7qkjdHgqLa9WS5Azn2nHGZLw3RY9W6hc03Jcli3RrGw666wXoxVpaotw4RIqcMs
5chypwUSfn0tpVAB8eSoOOnCb+Z1bfzikdtEtgZtY3K8gfHA3L4sUWlIylvApVtq
SmDhLsDR+nhRDbzEcGjoNO1/zu1xgyHIKGiMBzXuJqpEEntFkDQHWDV9EyluueBA
fTqjwXObWqayk3oAu2B8UmbfkWR9JnrpM9hDaQz4inz6wVumTrNbvB1+nft0H/rU
bVn2+cXoetnWxBlHeSI0RYOPzUuWdc4COvonudnH7GzALiysb7NqV9wOouHC8Rkp
DFHaeWrKtAmI9gJHJIlWv9c9r4WG72iplGONJ9xpFJftHJIiTS2XFr+mCO1UZE/K
kS/Y2J/pBpUgbvs5Qj5YLUK3kUNBD8wmDeJ1+JR6drnM0ad1MtOQfhrCbDuM5xYz
cYek1XHFvc1zOKHV8RVqxeaaldMKdGG2jhiKg0a/Zq27UJ4hvMzg27B4SPkePfrl
2V82J8ExjNcPrBgDp7q/11GRE/ZvGMo0UET/k9YwGfvNCCzPWnrC6KigStKlEzjM
Cp5ygo7xt6zi6q5FXAL5A5NFr093s6bjolKlwvLIAIu1oCoWtKd8Wp/N/g8qZyk1
VoJmd9zOrQztTJ0cZAtVecA4Y9NJCvePgAl86TSmWSk/JsE6V46ZBRkgTHTXe2M8
WhCcD9VklVNK2mg6SuaBOMfrueC729RNWY+gy1KaRQcrxAlOeTvnLRuf6eM172vq
65zSQd3rbQAGbNSJpbbS3Yjbd0Ft5camzEVEwMxmT2LojsdG6BC33AYo8Oh1I9Is
8uOLOZMmcklQ65QJBED94ZOrfDbTXLV9f0FjjvZcfrqnb/KEWUcDv9Fcwqm46V34
DaHXLKQAS27GAA3vFetoltaIbg8QL+mpt+EIS3brrIMSIx5R7/7B1D1hdQ+LBbNT
849j20U9j16wyHNMSbgzis8nETHnStz1NwiI8OM1+L+Y1TZTAuxeZM7JAcQZlmQs
m9GsSL+r/XFMJJDRFWHjATFazK8ayNycARPAuxcbLAR8aAaA+Z815fq8/k3WDmJS
garR9RLh9x4xmrVc0P1YMpYDDProGNHua12qjWUD2EL/oT3+caCJ7QH8SCcLuuWc
RfxOAK8P8i/MaRtpmcANGw41mEniPkQLO4CF8vKc0VlU0AJDbMTAMtef/g/kmbaN
VF19IXKjoOUNgNhiGSOaY7MFiCF5h6F119vbpQc+4XJsDBWLczOe5VUJSOLIpCv6
ioAQkM21gIEfn9HiTZTYhLNFuNl3mLHcQdo+ffHyEiahUxAv338z+55ULwk/0NFl
NzQtK6lpxw1ho0d5CmtQQwe9/DSK8mlgERG+USo5Y1VZy8CuNH48f9kmV79OBeZu
FCHxyjiza1JBNbB8RbOWEpP+acrjDWGgyUT2wKDZ2PxBgY0UUhBnUp0uKO+decX6
2hTLFgJJOraZ1l+XmpE8VPC6VjKtpRv+rAwO+Necg13rRmrYk6Ro/J0w2MyQkaDH
0GckDUW9mfOaSkAsth6SXJBbCudxUEY1ow6O6B9i5r0+4HNiIFw8owDRFO00anWl
ftUz3oU1DKh+NZfgWXODSxCCYQQGoNcV5hiEkobz/DMYmfTjvvId2KfTelqgwt5F
lkehTozjo12TIJLTCIYayf8MW83UyJf+M2NrEA4hde51V2XCJ8ws1m11t4isCk3r
MSKdIcfsTdRTPmNZNH2x7Mk22LUEOjFgdJ5+dE6693S31XU7DUg4N41dp1GBDSMJ
87r0xciJqenCsKaSaz2Se/F0lcYlAaGjT/k2CME4oI6QqOo1n+lHd+W/2nI/RuNe
DcBYjJXgv8I4OLmVyyZOd18HGPnlut02mWS17kljunoEBGEUEjNjEEUUoZg8WQb7
ytrgXKRD2c6yyFr0Eq9bKIIn4+OkDjKctR0Jcp0Hdwll+xng/Vb2QQkxGSdJoZXg
GIq/lrdwV80r3wAKJaWGSRkT9B7QO3BJM6X+5nfSR8vNUdg3RrBjo6pWW/OWvZfq
05V53Q+cdMtXrFgthsHGJj8Pf8v69W/vERLCcDNP04rFnYreP1CgyRvKP2PDY/jy
GiGkP/ItyaQYji86xk+0NgvCppq3CdDHc6p7i7sMcJcSiM3VuVfivb5782XYQHvv
aYttD9Swo8yyiTZwHuohX9qmgyQQppm0bEJ6iAxCG21gVsVA+CinXWIQ+fxjr4xl
SqnC8hNALTYkuwFoaPrs3E4/7i2V3HFcpQ4j9KvO/MDTvcAr4IjL50kcEwigpgPx
Skp+YRJAERaiqJcoirQjSuI+i3IEyQPnfUaOsGbzb5WotWWni3f9PjAd+G9s9Uwj
RvtjP1Daf7l0ORtVQLHrjtmfTicJLbWeEvXncU1AsVG0h8IjkJgqSlJ8OhCBnr/i
r6BQAEisE3qgsAfURqW67rttdbtTKXdL5iVZrnKQ6DPRy+GHlS/MDLy5HZvJtt4X
/1y5PgsEEn7KHSmenzIIj9PZ1Ix2xNp5/gvmTt/fhX/oGdJBkMEaBOW0gt7G4Byh
dYq+0KkErpSLYbQIN6Jxr9IZi5+6koY9bi0P1wYNHz68dhg7CEJgR5ot6FCo7FP7
57kyvvYAcYFsnMIGvE8+XuBS65QAdTHYdwdHOAaz1GQQ4UEvMr2E46XYWhukZ54o
K9giD0yO3/CHk94waajCyeavFiVv3kAOANDsPz2OEOIt6dyXxRicktv1Ef9CvKRA
YcFqAe4jnnygccOdBDUpJb9HtwfjyV0HjAm1PexftkqHI9nwcEtQUtyTGn7zv00f
lyeAz0AYP0cU1XLFbvfS7aTF/KR+9pgRahVAKOHjTsoIvtW9vuB2AgQ9PmxlVgB4
Ne8gwjpFN84Nyp0pKkCmQ49JgVTZyncnXtBQ+MbbFRX6IwOgxmNdBFeZ6A9X6T9j
hELpPidcCC9O/Z+TpQx5XCXXv5zi97Swlmac8rhkfm1OsibozORgTF7CVi5orTzN
hmt6LPTTRydO5wwaNgF3I21X1zRIYYqtbahCDCCO6qhMk066P/xizr5OSfiRE7Ee
dV79hA8wbIWMn/4d7w9FgiwyIkG57FgoOJroAaHy1rwpBVjlFY7QzDLo3tY5OQ1P
th6HVpPkVPZg6RfAw/OkqVfG3kqT2bOQ+an/JwJ+2qFvFm8OSE09eKqWV0nMRVu5
r9ptQKqWeuxgFYtCMVcXyA2WAjOzJ0+eCz1rlmjx2k8=
`protect END_PROTECTED
