`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kl+YU+ABfGykgr/yueLbUS6c8w6PRXcty4yBl7clUjQBiDCgjdYQDRt0gWyQ6KXS
Jc/d1t7WqqjIstDt3iQr0LKj3rfLB4cNfShH4oXNxCYSleXc9uXoibiE6ebRBi1w
5bPIQsxLxKwflhHbzYCaMQ3ZoGgKplcIzTLdYJbgKbyBGsNoszDmvvt26s0G5Rc7
mbzqBd90eu6S76VNEeDuuKV/lokpBF8amFTiLLl5sq1ssdmXYhVCMDzm3v8cBmwV
S6gmNUy4O/WrRJLOfqs1QdKtF6RJwhTMoL9WEpul5PaZ8mHO7BBovZdznMKTzP+A
39avkJMOu39xm5MzD5QGluX6RcBRAZuKDKT6dHMTDFQEcSs/dVbe/LKBeNmLzMCN
1tOeIXv+90YTTINjmUGgs3gW0PxvUsIe/Znwl/MRImrhVEnOU5nkqnxmC5B5c8/m
LCP/EMljhnnKHE4Y0socdV66VI4CFokMc0rmPPX6ZNwDgzAQG3VZqOQkq2d1VVln
24pgGKSG6WqZWqfPoLaOT0hZDjbquqlQfhBMR+Qehbk+dVmyrIJ20IvqWVitjwT0
Z5wkX1ZC3rrnhIbpnpXWCj/91mUdNzxlF56ygXY4hRIP58/OupgzIvYv6vzrrWhY
oiWT9f/aASgN/jznJkYjKQ0IbPGiANjzet1J/q1CBpj3xaZCeDybL3FiNoN0EgQ9
vRyfKqhxOuloBBlvc3H/sNipjOiD6yp+oIKQfTMRNQjMliRFjS8U1XMevp1OQUPc
7XlOvuIA4UzHNlgmRyBQgQ==
`protect END_PROTECTED
