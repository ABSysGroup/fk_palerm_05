`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Okc1tDchxPWQ5aJsogLYWzXroGY+IsJGpue8V+qvZ5cNmE/taXUz57TYBhOfJblN
8g1pJyvexqq8B1XBaPw8WisbofF0PWL2fOGixtGZKfGFklV8zopwAUzbstRqTqjH
FwU3/5yDOpchSwpG3bv37AkCORc8OhtgfeD6zY9znXv5q674OfyESKfAweZ9RCca
ecbvVAgaMz8VSgCnZHkdUP1Rb5x28theOW+X36md1V+pUhtz5kIuHPw+jMYPfDwu
1KeN1YP/s7xnMOQxQGhuQz2Es9CRoXwlUl4PJsYdMixbfgoHT7QfWtw2AUKvHSXU
Ge700EMcWVBpliu0aV+zAYPYM47NeRPGnTGO+gS+JbO0Vyj/gx5rBmxWccgHdAVw
sLJ2d3JRTbTyaHhm9dGMBYDuQU6jl7uRddoIEWZdi6GyAk9/kh7AisDi7Lt7FIDu
jwXVaLk97ifQyIGvlLe+6cLyDRz6ViqYJpig2XfNAbcjGsOXLbeqUWkL6f+qBWX5
yCzdHEYP2Kewy3kx2OqJVoFqvdZquISxOjpwtjh62Ju/9Nf3m+3de+h6ZxSg/RTV
9SJX2xL5hnhjBbOrmOmaBnmX6GG38lbaf267vFhSr8Pv5eByi1RR/gF5/XIZNE8z
00wL7QBjvjpvov8ofUHnzB1SDcRYvNHdp7NL4j+YGh5PxQn04+kRJfyoJ/F83TsC
GZBgWwZ5dZ97HoNJgO2WY8tKaZUOTIqNKmPoJPtSr9sAp80QygTOOfQypSIbOpG7
X2e4oVhrLHl/2YBqFJt5fGaHPbyauzNaiqB5Zjr04vltLMNX8LqhD8fUjXui+gYR
XY4Zc6CPRituou5F5/CUSeTn8G+K2f7XfowlVjmzT2PAPG5GylKDqoU3p4haEQbs
bpok42PiCfMjHvfqgh3Dqb7+sj+OGpk//U3MyZ1SwtAJ/xZqBo6/RqWvFjDcDt5j
m74N0KX8g47XMfzX9Y9P5w==
`protect END_PROTECTED
