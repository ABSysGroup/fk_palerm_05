`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eWnjBbuN0U3LfzJCMEEVV6iPUTvDLZHpGxrQs1QOoQ6mcWurHfIWXvnZ0SVp38Jo
qAzoJ40Dz3h8zUuMJBdegvsEtSV44pirYPVnE+ZTumx8Ux/cF15M4DfIq/f4AZXV
SmLYgFViR03IgGKl9Cvj8YUa1dO8BXLnQRkI4B1OQ2Ero1t8hZj0//O06+v0BxDP
sdr/Dg/UHQLb7sfNES02o6/N/Qy+RCLGoQqWBp/QwME5ljx/tLGqtVhr0JZjwpQi
SBCrJsoTeMJi0rboYQHdZHDy3kcYihnkbiwDZ5hj36jZZgkyFCK3HMqs0ZiBcDxF
7vxMb57hcrGagHtVDL2Jb/25NAl3WI1inCyrs1bhOECBBKUhCAoLRUKN+16tr/y6
IsdOwbBNLXL7Cxg2LJx/r0KAspa0qdJxMnH+ErIzQYuiF2r9nCALRJp+8ZogsX6h
KpRNrvfbHX8MswAKnCi2XIMndvNfBiVAJQghS3TfufXhf5b8Z0Gpt5FhZmH/V2DZ
0A9Gve1g2vMEd1bmq8+Dtm9zk5tsmAq3/a9TyoPnD1k1IOMZGjQPW33yNozhzlZa
UGUmpf2RHGj8tnDC1OcDOF1bup0vPm8kfimjGW42mJwT+VrgSHFFiacg9VFFjiWv
zrdao9IBw4IbiHVMMQfZqrm5H6rFjJujPt041ZprESg=
`protect END_PROTECTED
