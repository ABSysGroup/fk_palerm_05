`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8lhlSLsdORQ23ApQ8YKV/Zezu79XM021hdAJheEBuVQQy2IGj0ubze//9QnF2NTI
2g8s13Oc+f+XvauEcg9jcUpxdbko5vXGlmL1D7ZKkZxHjlMFNxmPA0XB8b5l+9EC
6B+LBC6p6BgMi1SRPGh32t5yP7z6FRFWwp4AecCthAvoihmRCqNEuIJMS6tDcsOQ
gChcvyGO+U13wfKkTEy/Qa2wHC29LcMzhF51VobO7wbUAYicSLvk5XE18HOALYND
QeOrx7F6jXnXl3ocTVUDJX7D20V1HJtAxUmo3xZy15mamgawSoafWhh7xyFsG1Rv
7JLwIZnlg3oMqmrLc0JHJA==
`protect END_PROTECTED
