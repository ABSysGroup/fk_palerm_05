`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DzABAujJAUSJ0NLIVcJmcNGc1fsEfoTvP6YaEaZSicC0LJBqmr+zFFykLs9OuRjF
LKpL4vUD3xg22rZa7J0EySvzjymVhsbCFGhdeCF8EQmbL0ScufQzh9E2zyu3aSPv
/IZQ+EhvqU5gpZX7ER59ajdaqjjPBFf7Cci0gMCO6cMrY5SzOyc5OXeYHPtK8FMo
ds72fAgfzTrzvAo6a0beyi5rI5Y4XxnPFVL2VyxFRrGSotBD2fxDsw89DH1VnKqh
d2uA/7txlY9dkR4/njiY7kElTjGlovlYjtjWoeXE1fErAESXuMqrHSROOXS2Q84r
l31k/x/cp2R871Cul21aHoOVBkRAKK3FdC5TPBa8Skjtg53B/O2pedFPxx2PslwA
fjuG5nDPFHSh6tQJRftChGWnqCwXQzKdU3p3wr2zwbLB3XqMDpihRhwLRs5DOo1h
uO1nxG8NWRHV31GknTaJc5TposoqQx1MhQBcQZ5w4KLLZV7EzBzh8rPeYQwOTIkJ
x3y1OGeSlrJuzloe0kgKTzFVQCI7K+w+XrqASffj2HUzzJA58CVepim9c02kZkyh
4cw6/NzEciax8YbfVb9e64wiRZQnBVMg/NeF/teOSMonI0JlJiX+aDcehlb8qDT5
zOgsJ3EvbaeQfTJZJjgl7m1dql+g1GFH9KMSOGGunqeDXD/L4lEwunQtheckJXMC
nK+ZK4Mbg2aXXQ6zikyOHXN4W1jmfrRwP4oV7I0QSo/PwnAmpVyVWF7UkqNT0ai1
Z8CJakbdk6/oBL62WDLLm2KShrKzeQbeLN1HWGBLFWzpJRUh2MbnhyYILIy76VcC
elrMxLa+mX/3zZQ1gvYZAKyOwT5U5+YAjHrkyuiWqin6wSWg/pjBr/pFON2udtdx
ePKgxG+8CcFWVxsDiyXqjCTvbB//yUmNgIkgZ3j4K60J6O7MV+81H7vvgwUi9apL
wHb+TeN0UN5Q/sz2BGGAhnQHEpe9BMI6A/zdeoJkgCyH2pPzLgwq3nZ4qRXZkcey
n05IO40F1RprawlN2WkdtdCtE2nlYws/BsgieG6zq7u5dhtlZzTt07FPCTa40f1H
Cc0ekcXXrWepMQ0zlZUqdckpKyNfczdKhszQy0nNnbuKWSotfSH7g67Lah+DVSEy
xCZMiU6OAgHidFquMQrTLkEFTHE7lYiFgk0TDAeqVmTkxCAu38PQSr8zir1mIqkj
NfnyF2I7qi/nY06fiNsCmmvvS2qMZtIeRPI2RlzcZnqiroWMfeN360HRg8X+TxQV
CbI5WrwRkOKSr8JsudduWymg/AAo8Dy6URzJlWb2mzM0qth05oFaBhkyDJWZXNRa
MNanu5zlevUAm/y77M233xx7hI7+6JADZK5UkyXFjWstDnnOQt6DPsGDXU2ufd5D
uHLe+OCbMstRIk2gWXCOWPrWNLjWGA8jp+HAX/5MT0A8SO5mc5wqz28Dx2BxyBZ8
ZCseVPoNx6uNWTgciFqAgw94JhMve/ZOAQyOqKPsHMvBrhyP+PGEkBqdouB3klxg
9xLsfwrR+eddmBanIowwUQRKNEU0Ff1uNCopcirS23Kr6pcpLNp6WnHgUoxiZKFs
JYjpQaVe9/1L0RC2Lu1E9fvbiU37hrZAd2DdRgC3tnoSr1W79N+/TejmTOS/xGsh
2u8qpsNhx5QrGmH/mcrwIZ4J1ope5dUdqmHUyrN9rQDnZ9OnFfEQQVTbad15qvPy
suCWLOsUMkuzWSLGbufhdzzZNRkEzl83z81H0UDriIj5Dlhl922E8stUjcsI0ReG
/tfHBRtkgR3jX6Bra8sC/s9LCSVegS+C4Z7oJtsrBNYvgmWIrb9lJ4AFu6YMKmSq
QtaKVe37eM7MNYGetVSf2lETkQ40YAy3n9hxXSBR/wMi/kgzO5N4Sjm3SD3mR3wC
jOZJzn22Q71F4b70TNUub/jzXXRRo8PbAi/xjl15gk7kyZNvDkka1NTYIHr0skI1
wATx56B5dli1Jdc4gOozDkDNiNsAL5/UVSdkY/gFmcOQpb3pPF7yLbS0qYpkxkyI
zIkksn29uViajrLkxtJdnAFfh0C7rT3pcPcD61P7bo4nxM7leuM7PA+JPEF/6mGL
EOSrWxOfXQ4HZr9Kt9bViyqQ4UXvrFDgmxLFCSx3/UvJM88LnQ1ap1jRdx8Zb4Fh
`protect END_PROTECTED
