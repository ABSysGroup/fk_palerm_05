`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q+v0+toG5YVrkb4JrbwCJrWni7NoLiAp0PMt8wL/1Mx5ZbdwEw0OxQnwRM3rQn5X
aB6sU/AGgbE9YseXquGLzhHMqAUUpiLolcEEp1ANNoAHovq9BhOfhZBZU8V2QKLJ
qDsY1xbe/o1F6yHdFdnA2ghe8MRuzCVQZfNz84skIxreIabZxLlkxfzfaXMM7GvG
08DCIlEednnPz6n/jjBfF1D2YIxOb/ksPTe/uMhkQVFNm3YE3PjimfdZi5v7i4a6
OMTuDVQXgAFdLwHfnNDcm/wXhZ5xONmXXKZlWEizzQ9I1I9I4Yv6xIOK8Ker9M0G
g/HP8dT9YZ+WrNZegjuhlu1jZ7WS4x/nqAE1yz1MLTo1ia8Xfn6Nb06p9scHsk+W
m1mKQnh5yiobfKbiFEnYXzoFOdMEpvoqTIq/9C29hkAbG+WhNDLEFw4P4qDN9Mu7
lWVMy57qFkgMbDxdaFkn3TRByS1FD/f06CB4pdhCYKxeagqPvyBmfFQ5xhkBDYh0
EwUUdg1oGuGrJPVjH7xOlgUPuAXWLaebpsv8be5r2DewvbX/JE9NMxV5M5ohSZAV
mYqYHDokuQODzcQFAtN4qJDFJaEz4I4sN6u4Tr8CjS/vpHwsBPwHfAeEkr03nqv6
Wak44ow0YoobWo+XrML23vtv+9UA42rZpqadMluH8LWlE4IN6fr6ebloHoyNZrLv
JykN584VoPUo/sdESL8F6RDQDcOtJULFSA7gVIEHthb6niFxu6NSXujv7XiDeIHv
7yOcnA6dTVi9DVs5jEXCsqLVZ3DKqNuK+vKE/By18dLCwqGZUYCl4tGRyxPMiNFr
L133ziKUJrVAHb0LEF9RXJjfpol4ESM8MhqYhnczUAkRLBajIUrIQ48AQRAOmtZU
g+xCYFXBNK59dsFHGHKPVcvM3l/hFZlb7plvfdSEMfyvymiCo+nSweRpVb7iECkG
CUNAfs/GBBShDsR+cfqFtQ2N/lhsqTmh55oqWMQKeva0+iOX8iObzXRSxYfuFSDq
pW4Du2GI+aewlzu+BZZMx5jnTjLWDNGmCyj6LhRP7y8BKFodNPNrPLfB2mEMYjkS
3vn6eMEVl31MLIC5JsAzAxk6wpd8VR6QbB6F+jpM4+ia+Y0ri5TPAlNpGxdnZNXC
2Eu+bymP9R576UWa+csiqlotH0kSdYLvYpYLDaMwNeJ5Gm0NzFnHQP2puTZdmnPh
kk942tM5BpQ7IZ2Wfcy1AWkP8wJirrIr2XoPFrKIX9/rkkQp/yt7iRnuLlxsDWhK
LV1kJShoBFVuNFntd/DmUZxoPg54E0TSSTa77qxYMa/o+wqXirUl64lViPAA9U/E
+ZpEVYaLeEoNxL7YUzc1w8TKsw+UE7yVZQJqSDFSOuXRM23fnmYvI8BTGSErEVnB
l2JmPPztTlk421kGadHaYTGDm+zebKMMI5NapClHgCzEQprYpahLUApAZx+7muKD
d0vvcVKdGRSdp57ZYRA8pOY1cLGoGADyhhpe9DU4pdkvK8AtUb9AjOR+CNFcH3bY
ePOVmCdzjnn5idwNtyPHUlI6aFVhY6GJc2zGZlL/DXkShKKkS3hzzP51R9FmYlkN
jY2GCcSmbK6E+RwSS9OiQWxBe3/Sn99kLM+JQFgZNUo3L1XoZfTdCjOaFe9Lx6s8
3kzdyip+Subm14UMvVyGQVoHlJihZASMSPcrd9THP2id4CrQq+G+GSnwfSLrzdTH
/rioWBJsQvF3I8SVvKCviybLoFSYJ8BgK5p4VhIoGqhqPCrTR7Dx+NE9NfU3r/Ay
K4GFmuS2Gb0H0EZDSlLeOfwWFiDhhzidcyU1QmNffFokCxYc1gyOAzACvNy3RMu8
bSzroqUF7RBHNjPnJKeQA0ue7d4Sh2eCrj4ceKif+hTiEWFE6dphin/IqytHlV4X
HszhpB6UWcxGW0yiO6WbNswuLSAocKzOqIiIf+AzkxhNTDeYWi7bAhZl5yhyB07y
EPOleGleJODXjj6zgtDQjseDTCgqtahIWV4ITYIzQ0I/YWTJcT03L/9y18z4RQAP
iNz9ff765bAWXK+D+JZW/u9T1QDkYgTou5TaWFoIM61TGy8iLdJUmSJvvz7XSAZ0
3jjECSw+Yn7B/2tH2tGqdLwRW+TQoY4K5S8aQgyx4YhXK/ViRM6GUBnoku+4x0NS
UJt0IKV633uCZ1LY5jjdyjXgcDXB+bzIaHjrjMjvAYvkHB4FNLAILHx4Mw57JNGa
lWJJTgVY2tZIEXF+6tJ0lhvmcbSdjqnV09zwKtcHMCPTSWu+yaEoT+cqNCVrKEgG
CN0IGtWjtgAVPiGDWhO5WIkLFuLFi7M5+m8qTd6FIIsoo2r6v5DYQLqp1NkRsrey
a35qie75VCuRsRhCmw+3vHGkDHkDUVKpv8sWDzQXtg2pJqGY/xU60p0KWM+tofZl
3YxTWMGly+o5N2yoFCpmIE2Y5wNmuQL9n9KG/Qfr2qe6BegVoV4QZ3jU8HPD/aJh
6JphhErfnIiZjvwOkEsTltpAdVe0/lEgsm5AD+N9O1qvxVIiuO+xHZNKB9/Qh7SD
0ftOVW0RSXCQASRXOmNeqD1u2kZgj3hBV5iAZuSddvaT43nlhGZZNcH7Wu+KWuWh
uWEfRfO4lnu2iGMrQDzL+V3d7N6u0RZNTz3ImVXPZif91Mc3B5NUC9f/xLNAS87K
jMhRCRE4ZRbwKzDUyYb0FbeBDdfNMoqgFzBb6xGELOSgSbfhCfbo6YPK0dex5iw7
rTvtMWEp8Qdmyo/dNjkI3lxT0lpX1cOwZzVzVgE9VeGSJc1LmTHJDHJJADD2VAsU
ne4/NBf5KcNwN245rG9Me3jIEngQBqqgezqMPNVR9/HrfCVIJ01e3S0wSC0su0l3
ZfEyMpW7uKtOq/QlPeLKLz7O/ds8bofIZgH36dXnI+0VPDhKAscEbL35cArQCNUn
vHKtvvs4bFTZzIs20tLTv5kKBauWnsfnwJPiqOIZywGLWdWvJ7M0cZZ8Y73v7OoE
iIccrHjI3GkH6m0iYp/6Jo2s2bQD6IK1Ly2X8Y6CkRdKmnATQ2Lao2nWgIECYG2q
9a5o2goBz9+wtfvQ0wVkzy64ULK1TAg+FIJ32XWfoyqXwcvZ120geBTynIc2dhP2
IV/vdnBb3xXDNN4guYvNPPzsX93QN3Av9GtlntuLw90e2bAF0FHvD19YMH3cqcgN
rD/8hfPehXSdAaVg4XjxZWyBFK20zKjGZc80HOLqlatOEVSOaH+4FidWH+PBVIUm
t2ccHmLRzAjYzmPsFkP3it7Z0ktg623IurjJ8Tvqu2y1E2NMoPkr4R75m1tyLHsk
AOCd48HOBAhEOYvIdcH1tVLwwkmozF4waHS39OZYpOLjaxDsrBE5geJ2FEuoe+h5
T6Lu3sRacoynqwb2rGkqn+NWH8kuY55hZjFYi2TkAaAxl704aCNWUSvBfcizIxB0
bucp3NAtBsKg0iS+E+CcxujrT6oZUXV41iq3MrVcZ+RO2k7itkgnhSyXJnGFO5/U
plFAu3WKn9/ATtXUXeI5pTSfWfbvmcE+GhR8ZYSJIHWCMNb0awAt/nby9hZxnSLs
L4il9T62ydGpiUiM+OvRr65tVO0hqMIQXfOYpd19vbN1RpfQAvDkabxBiD+s/yak
crCN291IlENnm80GC7F+FihgukrDZnv3lysp9f4k1YBV9y362I/oYBm7xfMMHVQf
aqmdslXun/XDuZAhPhToEqogUFE2YtEQL4UWFr8nWmFRdIkoy8SCS6tPirgVl5B8
M73DENcGC3VCwxf0We3PhoDlXqEZbmWonXMNkK7WCm2hGS21YyYP6SyFX5DnWZer
Lta1pVv2a8otVVmtzdrFCnKRY+9lYaFmsg57QlSFlI7+bOLSnACgyZD/CFMzM/5/
rtatHz14PvNPRNamtp1u/3p2hKVUoSgqoykzv6gq2VHq12M3tkDHvJePEUvk0xNt
Nklhi5crfpCgK9wWt7OJGM32VJJjDavPTlZMbXfKCOQ8GyV1qsTsmojlIAwRu0gt
n1nzkXJ94Do4f4jVjdl8lmSPGeelCvDfT7Y69lUxCY7RcoGGBW3sdeqw4X2UipY9
v4eoFKQOiEwf8BscpHdC+eEVevesF9kVFPDLupp1FY8cC6L0yf9DyDiWfJf3Y/Wb
FrYhH1/jpinB83Q+EDAwANuo2dMiPzjYnQDRURgBI8bjP8yVJSdy9pwwlDT1YOC+
8HlyarjAARpdgZF3NWoaa9W4C8iRB7WeD/ob75unX1u14w/wVUqOPhcNh0e9ZUga
UA9bmm/MVxYrZrJHja9lQX6KVjEMq9BX4+u0Q4n+ddKSzmwm0IQJActlVqsYOh3P
7nHr9xSXnyu7arzHQL4aM4EFFL9KxN43aL7V00gDeSX7HZburMS+xTcbCAN9gzeO
qb0ZdmQGlI2wLT1q4rFNo1vmYwf3EX1bgR/45wbq7PUsp7/LQ+dwwqfdJgMlS4Eu
PJ8kcPF73mrMZYrlvlyRJhNluNfnKDzP2ilvwuxsAxsvQyU8AiF+HoXNB9zzG+Nn
pu1ibW6aMwfjoQ5gzgQfgfhlDkgpEBgunzJH5UKYR5PSDqjbYAhBtRTmmns38mjA
r3Bd0+oh+ivPQySJJwZRs3AWrM+YSDjf106xUFDGAKqoHENBqQ2TYXhZ4L95WUx1
BjhTUm01Adg+KrBbg4eDUHcSXkltb61J70hScj/lylElTPDtrBIoATgfbCmVweH7
0wGFMmc4fkeFH90iHbK186iFENkq/XPpguwg6xG1XGx+AuuVpaUub/jlnhDnhvOq
GHz6lhO8HnUKUmeGhlXWsyo6rJmSF+aA/dFFuG349b0aTkoYumToEEMMh48UVXGs
czyidP2kQTs0clB5gMmkGcgQwDpj3SCJZiYd4XbiyQA71AYk8oOBibQqWGb1zAyx
+cvQmlMzJPyW3qxY1b2AdmQauFxEWXQrj1gdF2m2Ixqi9SO+tSGIqJf0PVAiIDa8
LtcXy+rc0nAogurSwhQc3chS/Syh6bzTWlQOPpuVqahaM+NE8ErPWayKE7Gw4Sof
UN5u+xnRuKg74IfGjuEeBLV2fxO9fpMnfFJ1LYTTAcWP2XAX0yrHnWi6c7qCCIg8
gG9TgLlDDAvu1q1+8lD0tQAdfLUmvARCYHRR4yJtruC6kG/ejw5BEXfuLFs/Is8y
hWk5z5v0MSdhRKGt0t5CDd74pFRkbE9KWFZRDjql6xsJNeQU1Ig49wu7iSadBsg6
8lsue/hc2SU2qGVeRW3rwCh2kUxD/c05FO43twBQigSLT3/rwafZwRTlORP7Ezns
iJ2BqavCS5SD9Erw5/FI765MRq9FdROh6RzPJbef0M1KKIxv3BHQQMySgVV2k24K
oQDy/V+TsNKR96I4N81vtKCmmgeLAdCduMqNOJTTvH/aKPbv/q2ViK59USItXIaX
/jSrn4swU5x74iP5uPrTPSQNBFgPxmtAv8bdXLpX5yui7P+R4/LbuwWmtbpvaA1/
nIDuR5eS2SHCFHoG0QIoxC7w4EIBrRV9LZwkI8fRYV0DQBrW0x69dDGDvlha054b
duaZkAgRtEi6N2v2WBM+ormb31EWNRqJJ5FxJCZguM7VaM1IQ2ZKGsZYegDvDJAl
WHqrTWBgMCsf5R1Y4i0p8KBLyikjdYfsfWXACk+p8MQ=
`protect END_PROTECTED
