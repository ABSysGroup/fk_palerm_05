`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FsT6HAuwDqvfoIbcOVMWAwssFdkAB+URVYhhfA49OZg9OwZhG1f+ruwa6XS6+96C
HpQa3OUYO6fBdrsW1bPrKQIRtGI205lwBwJWUjgh8Yq8uLfglJTAEnZ6cGo1xHBF
zi7Had5FjnaXWkCz6mSHRWjzmqwTc6Z+BdUPnorbEu03Bd0N6YW0zQIBZD7u9UsR
g+Z9gl92zLMCjBG/PnorBOwm6H05BU54w88x2pMEhR+QYwitK7UIH+U9gvD62I7p
FxDQYUChUIf6s8jPu7LzZVXwpkCP0A7O6QIQd0mDqK6xZPxnVrj3P53otHE1lswQ
E6rrqDEDYSwJEfn7XHCZqJn15D7Z9LZFwUaCtrZyX60AbUr7lDx2u6hYDq2wIjnc
z6OlLqjgn1oTTU+clAXZwj8TTm0b8tPuwdmFRUSjKv8YTtAMIf619bPFXJCY6PnW
F4RBSEHbhm/jES6eupSuMeSnsHCFwLfJ70mA5EPmyautgP3Zj0v7G9F095gvGh2P
fwZmvAKPZT2N1MT+TJAG/lBREHk6Ny9x8F91bDYD73NYkCsXziYdl3fTS3a8UVen
QO6YUerPXVvPE4Lxm3+xqan4At8Cy2wGO2bYaHQSdpSfvjDQ/qvqMi3XkEClMtTq
HCoYa2RSV3wSq2rv00yihHnYuGG+UwH0J2FZaSc9qWP/r7ATBu2GMSL/ctTpWcQc
yaG9DXYYSN4S2coi0K2rkVH6T/dOETW5iJNE5Kl7daXdQ3VAsgp7FrpmIVRNrdMx
Ak3ob88Oz9Fv4njLainZLCyVA6RHiRT5dt8oJqWIHZfuwKpM2pwkbt99saliFzYG
BFXagH2V3ZKcphDrxohSIktaEjQ0vw5eWDFbzKFEdedu9oQq0+XAzbiB39bG1j9i
eARxsIOjx6W1VlGRqUwV9tDlQA/rJMJZ0g128JC/WAjSC4ILPkvNBL4+CR44jGn8
bIaXtJZTWITvAZPHnlHxPvvTEHK9YrmEeTs8mJf+Ehn1j6fAV6B/ZMgRBG7vFSzT
4Fni2gXUr7dLZcZti9r0kUl0SRzmFaT5vJ0s3PsV96MPfbyUAiH3OD89ufmusIBM
NlS74hhJK63dDYb1nldR+yXHcG3WL17r9/lHnle/8mbSIfpMhelN43EUDGc/+7fL
+C6is/r+s7lSSXHE/PwZK3lhAb1faWktrAOtmhlYdAkPADcrWCnfuY6eIIDoaWEA
HRcU5cUjp/hVzoYND9Aw7YgQ7Th7jhKHy73qQoLnaP6y8opQEFXFjBZDKkxxvbPE
X7ZT4TH9TGI3rCPHUZC39KP/SwQh4lKW/SGPFwmHoq6gNi4JHPUejJ/pa0Mw8+Lv
NxHiwRCPPo0ABBDge3Ri7yHIwpvNHdZ7zZj8UexExCRp9PtJ8l0HE4I5o3J7NKao
R9M82V1qtqXOU9oz3qYUGutt4aAukCRgZH7NVN3pY80yAFnISqqD5CYlSc0n6hrw
92l8ZNwAZRC9TI/mBPoUQCsds8SL0FGqVZ7p0fdSheRMtSSYMOFHcu3N73nnsHiZ
Vk3AKD1NwZ1tf/5Burmbhs4zGBKxOtyhdtRtADt5IjVfenLtPT5hSf4KM0ovBGkJ
CWsOR/boUOGq0/xyauMtFU3dnAyu+hwBD40VlSdrPWfADDA364+MJsXULHQ4qGtE
PsWdLAf2pmU1hBDE6qsITS2XD0ZQNN1aQgCJJ9M6N+tIjIehW3AXxsWaPSNs3RNa
BVrITgIsW+0zOsh5a40hyVLjht2lqpRLfek8PBEKDrer+x21j/ZWedrdJ92E4KMh
CWklNoCC/fP/gfjnZnMAgZqbprcp7d65RcIdrZ4IFHqOMMhMH3nnlTNVYgiBcoPv
2uz1iQKtPhagIH0wXp/zf1C2uT0iS4Wc79KVs3LdeJRAJURRzkqOECwUuyrQdQZe
/hSOe+pAufFjZROhbo3xPHnOHjA1YlT5x2N64clGrQel5DlbI3KpSYa7EOfL9W/j
R3Tm2UYndYzNC2k5XDobsOK9icTV2K/vQfqJYrNu7gU9GLrmctfG+9z/2RD2YGdB
Sx5cQejTgFhy8DXeKuE0CokekSzjkX2Eeq4YpWpKvG2OC6Z+dmJsPOOKO97/FPwT
SdTytd4XptGmHuFZe8QuK/dLBtaFl1xoL4ytz+SlJN0=
`protect END_PROTECTED
