`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WtdiiRlgMqr76F4dtlzoyKvZGkHWdsIVQWc5nLXiw+tyYbhvTfvxdEoUX0pcYHcD
vx6JXNQLl3xXgC5Og5woYtm5ivSZwvzU2snce2bEabwRRnWaJ10a3FuhArNPbCtV
64t79YqI39Hd66I+Nurubhjz3WLp3b+m0PgHopdIKhgj++o6z7RqLtaRESsVqkK8
y7wVaYPUs8bkbCZ5rmLy+iRgIqffBQYtfS92w3mLAr/cM6FX1UsMyvB/Va51IA2H
8Q/zdTTuyBRL9SM1hgYR6McO32e4fXgth/hEvGdE3H2BYk3TNu4uccvVeRh6nE47
wG+QOmjcUGAXWXLaaLasljqGrZMMVxjGQZLUQ9BzZDplnH2AGIRTgwLXzwWCMXEx
9rBZEokJJZ8UKyC8o7m7bYPTBLWMfi2ZHz8yi6nbOHIWl6lftWCInSomD0aCuX45
YqjgicpvzYzNn+cVUUiTME0I/dBZxiI5qOYB74FOXlWqAuXX5ysXPm3/c8stRye1
6R/hGZjHej08QTB7P1S61NqtsMc4FfoyoZJoU0ScWyvSPIsV6f/k0Lqhi3jsZn47
Fy7i3ZOm9E801V6aaqd3P5TjeawM30Afg+JE+MbRTyOB+TdieST37sdbo9plCdZH
a+SAu8x/vpzNhubHSlwa5hUVDmdJFjL4YsGv38vl3iYIA2h2EEs8vnsv7zZ/PqIr
QP9OKUjOM/s3BV9msc7xlkY8koU/iiD3Y45BpPXLUdKtiBoW2sHvsR7otdbytcZg
e+pcNU+rMOawJmc0juExczSNL4fghs/vtpSFOXGlb+SlSzGVCugg/kwJH+Tkg9Wo
AYpzbdowFiK3crD1EUAt/iNb1/HadUseGeTLEJWJTYWB1a4ACBjwC3OeiIUSVkdf
I8nvrovERnRZdlODsmThsq34Mi4EG90kU1pSkwOshzENqrzTxOl+DLJ2J7ncPmp0
h4bCeA4Kodld3F0DF4CDt9wI3NylgO1YW3UiDL8IQgx/DXM2+GqHKznvUve1LDYf
rpPcVdpPpJGKUtLPTmZgt7vZe1GPktrxfRhXYmAzhQY0INAIUjUH4yJ1Idlr5ZbI
YWWHfoDYP630VUEkPLFTW1QhD80U8IDGz5M6eeRiCuln5m6Tg7VPsvIMvIBVzyrI
QPntCceJvpY0LPtMZpycS8akmoKpGyuSgy7YSqYfcydFxWw3aWvNWykqTVrfa81f
lsLCtZuTVFUW6D+I+h0Dfqdkv1YNtSxKLUsVy0CTdIQpLa1mCm07uhtRIjptI2up
21cKuCL3PKY62r/8aEFFa6tpxBYRvZ5H6UfnZ8oYRQXYogeCIVXq3MvAIKhGJVps
LC4B1Unpr4FtCA6j5V+Ngl3wzIm8Iq6FO10LBEz38EZ1TqJyKr3zUXd6JRO8gglA
QkUJu30VBnY5WYsfoOY16Py58WZiHwrMoTLJqqhdtD0pLwPmYvAHgnH5qAYeQdhm
Fri3ZgVj6j2fSLWas/CEaU7fJYSuaNcpI3p0BqJAspMg3oy/0NmCxZxGClbUEALU
8b7yi0IFd7NG6Dcta+YMUZNPWEXuRAby3oO4QBxgy//JUUEpOJWAnyJhopnowKfv
nIlNobzv5ZV9aRXLHOK0yCzCOvdVZEGoGUmFsMhM85aQbuiJqjRDEgze9plMiG2K
sQTFs+UUhjBVrdkfEhWMVLB67Lq2pLIOeASFcCCERjcjzsXvhEZaCllCdIcs7hQV
rpa33gVmK+zk2Ji5w6nEmWAFTstOYa67tchKmCoZCYYdnFfcwNeyhLNjNobfefIo
D8PtwqFxjqVYgTebYX4gwOE9wP9zMG26ySrZ/yRH9sIQgF3aMb74gUjl/n4fpZ6z
JIRu1F9/VJRg3Zt+KxlmdHECwz4hxh0RHjjiZDuYf5FanMEmootohXX/i8SDMmzp
RYd9nEqWAR+WF2Cqx/bSdtHwlkKySUpeZssGmxl2ZVs3ySWLVo5M8q2KGzPIqezk
njvYSJjBNuMPAg35+yviCh5KI/Y1JD4XAOhUWhPfRKq1DNAbsHJ4THvjX4MnKHGv
ktjW02fxjop7lyf9tvwM3KWfOWtHrrQXiCT+jRAcg6Ihh1RnWk4zZDA/vQ5kVjBm
wNrE8Ux9qBxD7eyaWEWIgeiIqF/bHk/vnH+T4cT3i+3UpcHP2udQ8W7g7QUE64X1
3KY0zJu4zNkm4aUrxTPVvh/WDJmUgJnLAKWQcKpjkh0Lykj7ID6aEIOKswHcyni+
/bCap5kpsdGwZa4WDtWrG8BaUSvu2xoCHIPRAaG7P3BEJhM3QRcjYQfyQbap2Odb
nR1k/tZreUo+vQTd7LY/fUes4R6YLTThuf4PPsVuWjYm/ycL3AJgPaElDoXKDuc6
VXJKAsOT7Z4jUlVoRLXwvNkhTc3FjKpuDyrLvOQ+XsjC87FF4cnPzOKLsNukqZ5g
Bv/31FUHhVK27tPWMIfAUuikTWRZxDgy3qor6NSt6gy2rbEus+fli9KjDYNwDH4c
Dnf6020HLQGTNX45s5DnFCK4rCTSeQrZsL+q8yGhIj1mmKTa1auFU4GNpk2Vl2cO
nkqzajLVLGhXDA10hAu8qcQcCdVGvLFwu5WU3cegEJ2m21Rf2g7P7YbLMcK9kyki
9wi7JQtfR32pGF8uMmS4tt1lT36JSW5XDXTd9zfzPr7IowhT8FEQSTjvk8v2RTj7
Lzv49vG484Z/2YjvV7TXvqh40uOUyPQeX3Jl3M9VPen7gskqKzTFEvbI1z02BqI6
gI/JBMY54PG7urxaNr3NpGq6osixS6GIaDdRSaQUD+2cAlj2iMeknGjBrvjjnvpA
bdTQPx9lYasr6BUnipafy0rtOYPH26whcPzPZAvfBB8REAnJy/hooRFEpBSk2d1l
pbgwsQtNfOXl4apAuZfTslrUzHQxHEkFFcpM0mhEEe2OFhfQgUjreo1LIDAgqblZ
+wE42QGUiM4W3ebR69jaDG0X0p+vyYK/HZHt2zLmP5/1II8TGG4MNdlmWSeWOtHJ
27im0Lef/7nQNPauUJWe8upfqcrRkd7g+5CrbeOmdQiSdj7IBM8XMu6pLGlHzjDl
ZI3/HJtAOKaRoefL0THJeW7k3TP/3tekmxztjy533PFDwVYfMWJXJ2e/kFzCI24P
`protect END_PROTECTED
