`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zocge9vsFu8JhUtIGG46nAs2bU+pPU4IcBziDANmb5T97KleCJKDYy8iS58uUuPs
Ja7DJnMgAiJ6iZGvB2GBvtGjwEFz4No48HQhWPmy9PC3beOiuv1KAR2t7bq5Z9vL
k/xQqMXhervG4737OjbtwoG2RX8tEPbDLtT2kJNdvHXVT5pGSRro8fX7ZbcSRYSc
HxfxEs3IC4q6MBk9ysejks32QdP1lgnrTm3Up/nrsA+9p4DmoD3esVYM9zHjQsLp
AIybVk13NCXQ/OngU2/dDUNo8+2fOeF3naIU2ZKYi3V4UsFQSysIGOj1lPUgTGaY
fGYW5MTx36OI42oVCKC8JBW3681oo0lyEs4bUKnpPxqZizVUoYo5gV+60pnhokF6
hl3ENYvJvClso9Wd29fstzNzQ3BkiVc7lhpPo76ku1kgWxy8TlLVgFfIAGESASGZ
mMZJdK0aaijt3YFTmgpX5AUxsVtbRKS/EDTtH+7WpvD0NiQcW1uDP+Uem6AP1m6e
ZYknWfimnG2fuwGxDqpIOv98ds0Pxfx7EB5/w1lKZnk/r5YR1SYKZFVxc20voAjC
IVA68D2hvy1qUdgm5xhC+E3SIfHurQZ+cEpM4xq84U9VRw5MXNbAShsXxjWlJZhe
tWDsAFLpiY5If3uiZJfFA28BAGOvxpCnCfUwKVm6Oj+nox3lYb1ay6JlFLQhbMj3
pTi8M2xywD9goXl+gfhMp9r4kyPmAJT3wIdsl5c2hLLI7laUuTC+3XNfXBb6c5fU
mrQrmEPuJ8dguu4vhkzjAK1SgB9JqHk1GlwFZHZxTr7lNNI4fIjLyRWQilL0yf/7
HXDMwOnYMq0yq4tYtPhb9AhO5N2Z9lWcf40V+ieS/NegqvMMozSWNBlUViQzW7q3
bbes3L8G7YcXZiwC8WCcM7l+joR/CzWvTIoubpjZLeAMQP8xcoE3ccwDuuAYQY8A
`protect END_PROTECTED
