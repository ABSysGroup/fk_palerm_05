`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JD5rw0Z79xwMdSptQveCm2ZuABCG7MlO2BxYi8zy85u6sY5ebsY/hhdVe9Z1ACOp
p4taRWP3mQO7zzuBBHKCWymihO0deHHGmVxWSbCK/lXjSTcl8lwDXoWjlL6M0loT
DqUD5S3sSNzRTpgk+rm7+y82kU53i+UnkfUbxNrSuUygoNkFy9o30xoiqznJSdDP
aFxnEbHg/jRYh4MMQGvG1kNnx8NgRWK8h3WC7O2zijm8na+ES/gQZPdyQ4qZSlKz
vRqlnQ0PxRj2HgKXZ1JnzF/EsXrg4iZVKG079i62sH3A9Ki4+w2OnjgouCXDT6v8
1WJi+prbSKmMKfugrrbeT3Rah+DDuqGo+Kygxn3sI1DLeyWmBUqtJkkYkOBlzwTY
Em0NqD2hDPLTxSIyx02NeSpXWS/TS54/YvGgua0/xpUbxBXxu2wmLVbtph0dorWU
U8VzpxA6WB3BMFzhXBv6FgaMKGCNAD/9nXb+KAq5eNqBQAwl69wUKSjP5OsBzpqO
U12d3RTrvtqb42F6D0Pfp6iRMj/6s77mPgrSzN/v+zeJBlg9PSwEo9otR78M3hGp
u0eAlFOrIg/j6o8Xn/4by7jfoNCnI8jQNU0dVvVM8fPE4wT2xj7D/d72LDaBlmKX
/WUdP5H9A2yfAxHeKcM/75o5i1OzIIi1OmBdHfpUT+BJtsQlg7RGbFyIxk/exCnQ
mm+mpOc4UhzP4O8d2eibLQ92UzaBWr5trJp2NunqdGrjMV8uijsZeVu4NBjEmrC2
pn4e8tSvL3rjuKZcKezPbv+yfPlieYibBP+CvAlNIQm3Vf3+KGAFuh0kl/Ncumlj
4L+eYKLVFD9yO2TXhs0d2CA4EFpyH5RdAjPkJpauNGjktXZwzw8QRvzVU1iRxGw/
0TUamY9YJYP4CWUJzMBNHNSJ3jEVWMFh6gAM+eHDB0GesVlPONIu93xpUPAaGqJX
RQe7GRpyOWsplgBYDuTT5Y3kkSabwA8RbQh25lbGpsyvV8HL3WgmQBMD6RayVHbW
DZUBxDNV4yjwRUqeWMJ+vkPIIkGTisK7xmES2/mD9yXxGeEXKAoupmHeDchP6ca4
wjmqnWMvp1EkfM/LvgYzAxLDGMZiUwdiBy8yYC9sCaPe//WYv4hSPGl1NM0Dwanh
GZkzYqYEJHJlxYvroftDoxcO+MB5eoSfaiPM1yENRXFG/yu/5GJjz8u2PHkQ1pFB
rxqIiayWyO/s24JnAyQxAaDwCrYkr03aeJircLZd0JF0wLe81BAfcMy8y8GkW53E
2KcDf5B4NYMgjT8teDlBi8J80cr8ZNYkeFvXZr5Mr/4MtHsh+iSOMOgl22GO8zqh
QS9bgDU60Dg26c6fC7CKwE7WqpUAoaZMAXta9qZBWGHa9aF8yrDIm49C6k1jDe3Y
BbUjArrdHhztQ6nt5lp/vjFH4LiwLKGK5PJE0YM7wNErfl+i0AhFKeXsDKoSr7sJ
UQ1VJdm4IHWMJFfo7gUu7W+GfTREu/SquDoayluP+xUnRL+C54fmZbcSwJBVpvPN
+vNfClw86T7lH8GfM+JQYbK7qJ8e/Nl14YeyH0yKfNoOw5awUyUypdV94TJkVdFv
qfy/le63xHk2VQYJef7COzGR6ZzRC9s/bktcRaXoxsuHL0r5h091i/Bja3ZXGjEK
GxniPE7LGo7z3WVSkd3QXSrCWqzfObYcIU14iCyWHSdl2pYq45/hBwgEbwW4i1W0
croznWpNitM/KiidSZ7jYRwkpHzLP6/WgFLxoyzD9cajRjykWnn/g6qB1N04y2rc
3C7xPVToLGkRTLNG+57ZdiRRAl+BNWxIIl4Vfhbwk1pl4+QsNicbshifC9MdBqIp
DDStGjeUvCC2BdEJitHMz73+qLSC9+b8VANww2bIefGDuTXHxNxhgrwXorvi3qKI
ZzAyWjVEGQa2C1aKPQdiB19xZCWshYWmRTSNulp0QYtAadj040QdJvp+ml135FGT
UAFkky1Boz9ZlaAxwheK3I7tG9QUi3WhaMncGjcasqV2xKHBKaWhT+MRBHBcPieS
WDm4M/HwMmJattvCdmpIICkc0lqCRvLaeo5KLB3yN88CLN87Z45DAlioPDwT70kn
oTGWkshuWO5IjyGxxeyBqXCyEgs7ZZOydzh0KsTJ8O0eijaw0ahNUvcHE9I+E3zW
JD/JIbVseG6e+dTt4aLzHJaO0LVMA7eQdbvLfbWjIMA=
`protect END_PROTECTED
