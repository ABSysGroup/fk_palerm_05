`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kjloICf54HEaQ3cC/foYP6buqUVY9r/A9INKeyUSSfCj5UaIpABGmKHAm0g1H7ot
r/1eht3n+WjbXaLdTtdf34Ld7gxtOSv5UP8viVmW17Z3BkL5xPFMx/87Ay7mk+Jc
lvW+cyJLN/fcuG0udusUuKsTZBAAtEOQKwsIj8p52gCrIxj6dQPN0FLStqY7nGcd
/G3A1VAHmoQr60FUnjXOlNKkPLAoItCmSCJGdEWtgLViz/YgCcAq3S/xjQ1xrWja
X2QJv7uD+Y0UTTyp9Gwj4rkbB3u0c5XWQ36wB9K/rOzu3dY70xjlZ5ZmiM1sZAGn
637ZpcZHsTiPfF5VdMNVrg==
`protect END_PROTECTED
