`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hbYm4/eh1pZ0TRMHjyvWvrA/gek/9kt6Hhn/ajVcqwZ2LdcEKkIkZw2vveeactSp
qWHyXk9nyQVJqeHvoHBkVKpF6+Ay2R2e5KBBrWHwk4oIcPnMDoFu1hRQzeEGIn/P
FiMD2J3WGYBFgWWyY+l62krvtrkvlHsVGhgjLFVFyMVZmO6uvNxaJp3pSylwhvkY
4Ia61c0vakwprP4BdpIJGeYMbemnaPDwr9NBdTIsG3BC5mcUL6IMDkQcNLRlw4ij
0sWTTErkJW1aZhXBqcWvMDfecPs9C99wXZ5rNZF0EY+bodzlyXRRkh+NqTBftCQB
7a/Q7s+w+kwrrOqUQjTM+gDsMqgMCQoRDb5ddT+2MX+BANMUBeNeymM0YKfPukSE
XqvEe+Do5VnS6UJX9ahvYglQumVpdrksQg9PZ3F2hJrGFWK2QJCFWWAWwYmhnTbL
YhiKZfxox5cyInHW1k3PgmPufd4o3yiYasEPBqPCVvs=
`protect END_PROTECTED
