`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D+h0n4wosYuHK+6yJIPI0yjSgsLuzSesuW6nOjaF/jsaPICSI7hfcgg+utwKjZ3C
e2mD/QCN0PP0Z4Q9SiaeXKVkdnJWOJP8MOu02ZYwANGOeJ79hE+dBiQuGtKH1d2P
KRD03rCHGk9zKMaVzRt0jW06AwY+mKMzfYcU6papiLdsOzeKwCWC+18jQu6iOEKl
zamxnz/soDJ3M5ZQfF+3hDHyK3MY7Oenlfn5wh7O2+54ffWAE/yq0YfTOWP7o01G
vjYPZxmRpUZph+qc+8fGjaM1ryFhDp2JUrmtfgtjqiGzAFPeOcoGqd+M1i8ihxMa
h+t/pzZeUQkwD6H6hKCD80D5a1ovc8prTbs6tPNfwFSEBUBB848cEDFwIjVlo22V
DX6ivgrcsao6okfp6K8Xk/JEazICPSLuaBYGow8hwkx2OKfm8lbvaUGmYMdRbnDO
IyP8zDLmOt5gQLGBKcx0Zddceu592zVER9hagW+uuUuTciJeUbn+o8yrDunO8t//
9J0y4U4wyr0Ubsa+Lg/8b2GaIv+zHShIMm+M7MIV6Rbm0yetNFyr6hobpGebdkKI
tSTI2DwoKEJrP41B8jlnqKx/DDCNkRlpvQD74e17pq58A4jOUJJlW9D06NDrdkWz
u4pDTvvztSvqotnsIN/MGw==
`protect END_PROTECTED
