`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q2rmcpWlguj6Y+fCLbgQPP4o0cp8fF1Sn916eVERIVEVpwF2HOW4LxKVbzmXBcRK
WEj+a9u71IUl3sW+rQ/LznR951471UoI/OgTxZYWzt4sEW3/y+Ff8+xLWCYDEDdg
5VBcRQUV9nHIWZnh8o/mpRn7fU4Yhifiu21PLEIp8puYuMjvH9Bm94+v2Jcgz3ol
1ZxVstb/f3WQhW4Zs4Sls62YTGIwOzl6WWmyUlFZL0/jxQ5gBPOicUQxULlqCiI4
`protect END_PROTECTED
