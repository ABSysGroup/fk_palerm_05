`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
57NcPX6cqAL/Kb0hCci/2I5Sd5f1K8xFpqdwwpHjVMXtU5Z7G/h0O1i4xI/g45LW
d2KUMRFe009SRYnSfrnxrwogFIqDrRiezIY6gxbFfRk6FEbDTzPIWkKz8e7A/FBN
1H4yvdmWuoJLuthpUUJZ51b6a+i5GvP6udsA9p3GLIq/m7pNaNuNLeHXhYE6+8QY
6Hy26LuEE6EPgGyTTw0yNNT2m0/6h0QUI57aDnQr0ggjyEg2zF4sTzNVmDOPMt1J
Kp51kXPkuIZZz9oQUn5CM0K94T59SZXOgVuAuT8fjBl57FCC0Z0Sm32VoePyROg+
Emer8cyqM0uubHHAClmxVqtS2TIX4zPuTbwX/xKKYfqbqrra6RKlzGUnRz2ueq0v
f9zfVvHZp2QZluvld4Seo1LbsZ2Sl/tg7ruDEe+30OZIcwNHtUtacLHtrvnp4R64
d8XXg0BpFmURofoPqAlEWz7/QGIHrGi9ZxuvSmMT8pSXPCtKCsnMeE9HHwgTvieh
10YOL/zHJAKf70E+dynWjpCh33rCo3/QUDR8+gvX6mT55aLjXn1YHGOCP1F1RXYI
YS06smQGQ1W2AGdz3GO8pEncKPKjT7klsRuG+UX3RwQ4zw7fpu1IrnKVJ1w57M6C
an7IjBL9Ow+eH+bQLpn5S133nRsbPQKWxlR+it4TQPycSRAm9RBodOTB3TjvlG50
`protect END_PROTECTED
