`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vaj9zl/+k8TsnCXgkYIsWNjZPVRn8XOmbF4IkGRdFX6sJGSPIW9m3aALRQPojeQV
X9qHDWmUXSTJ/zw5sqDOO2r5MlBjl5BcoEDD6xdwxomhVdnthkJjyK08TGqni91b
anaKElceKFA55eN2PxLYD/HhNdKSoSiq5E6QFuVfA2CmXriShN7t+umLmDMzVgbP
awf7cUFpHjmqQY3j47Wd1l33QC/AvX8PQu6pkhgqKAHPfuYdM6T/e3X17xRRHufy
720aDJWOi6LfoVAdcLAXveh6YohS8hGajNPOp0vWUYb/PFD4+7hjdhQqBAKoVdc2
BrjnWsrI/FKQQXQJzMVMK+yD+a7eO67hsBLhcX4O/U0SGAiA8xdHb/netWz+cn8x
hbH4Lohcm66dqruTy57iT/bN0iaedE+dM83z4FNPjbZAVuwCM4+T/NetfOVl/3Ut
OIKyWmTDaItCMXe3Et07VfMnTYnQMkuk2Ltps2cAuQ8GL1lPvuafPnvbMS76Jd6h
ezMi0ZcBOZut+0GjmuvZV9/C1yrsabfV9DcmHZ2u4TI47M/NfPb0VOyJjCrXBWVt
YiHuBlzH5G16gFMRSOfcSwR3XUzuacrIrqnfmkIzfVUlFQoEbGjqrqUJwcAbvB2h
q7xWYEVUzZzRXibKNvE4GgsSycKDgzIkdO7NfmsHnYSSXoK/Qi/sHeENUR8K7H2L
0hQ4bPcXIlmTFhYSVdkJRtP6BsZMwSkI6uenbk/aHOnieP58q/CO8LR4JY/bpHOk
7kN6d5B4Dc6Rdc1V/DwPm3UThCJLG163GbkPzCAOQMtcXsfD99dqrlRaLPCpkqpM
hRskkJQBoHk/qFJgnuyg8B3GD3bO+5bsyF1bIQ1+zwlUiew1os3dpVCl7oEnOjOF
3jw0D+ZT/armOQAqBUwrhe/tuijdEjuOWIcDmSGK6xyp6j8lmQG550cefPK8uegP
SrCIqFeDIevQjYKnte7wn4DVuzlXrR4BeNJmqED7rYgWCjChCpN8aIa7KyCtStEC
BH8vtB5QX2i15lG/MzC/BKdXVdVXFKDn8Z5zfUY7sZV6/MR7leX2MztFCQOmKZtH
a6Qrhqrv8AnOeZPIjri9rKZTLm5vB9bggnK0+jHMCMHCqiT5q71xTa7AdFXezO/Y
pRodpv0jKBADOSjPX2+OPmDvhxW2kd/jjsoIv5YyfJ5jSS/DdfrYgfoxMSVKNyrh
sCOtlGWM0Sak6Ni/ZKB0TtjMv/91g1/avurDnsaQXOCEev+iZsQNMBtnQS626SHi
EdqvE0EoSUnRaDv3v6ofAwuA8SxmHUOgNG7kC3bJ7gtRHd9zonCLQ8FQ27CIYsOa
T/P/U3M2bbP/MgWl3uVC2Y825zFq79YlZOygjPfaUpQeGyJERasnKlwOZpPvDLUM
REVVLJ2bXRKIcZE6KLmEZa+eIOGuxSAT3C55kSNSazztMdcDYpjMouak0ScENGbc
dYcW5NwckA3IyALH32cfdoni/Pa3yQlMl635IyvE4lbqXu5gQGk+okDiyn3T3p/N
bM1RT5U61hufz3lMalMrepF+P7LWedMX+z1jUBaoZdTt4pLohYOOjfAT1NXgSItK
ihRjV/qrx7d8ivd/xkJ6ECUtEA3v19Wkgm8/lyCoDKvho5KufMQx0R5s+jxnb7+p
lGAlx23cKZTSjvjeffyBLRR2nFESXNtKiH74RRgCrVI3KHz6FzW6jtUXR9onMSwZ
/zS+lQkuAKZNF7M+jIMXv4mBz3Ov16gfb5eUTZcbE7rOVmqBfuk6cAOcq9aK9xzL
kSssXDAkJvLqvdKs3po/pwQXZBN4mXWIZLkdfwzvjgcEl3QDAusCzrlC1a7aNV5f
vY56T2DEklGQYwbe4wumtdT8AasnBwsHp6syyFxEtcV5W0r45Vdzd7VHE+iqSa+m
KqeBLG+9vgDJbtTOUsSeXxEEPwzQUTmjdMdIkuUM+cc5liW4mScBA1VDB0PmwBS9
7VxhrmsNoZQw3NbkhEwj4PKXmYkaXvfFu3CMWzsBIDgrPLEvcHwoIA0PaiiJ/LBq
EOkU/8MyGnr7VR1zwzTQPtcgaBYjEOlv/za8I0+82cZnPhZsMoKTd8tmiGLipRe1
wS5ZTgOXYQhRc+AzAlVkfixhV3u3ey9Z+HDF2B+OYyc=
`protect END_PROTECTED
