`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KPLibSIpN5BZg20b0XPbSQ9WA7nYSupMQoe2vkSX5GL4Mmcd7EIb8NNsO5AgrVxI
x7YVi4Gm2c4Y5s1kCwlfsi47w5JFXRUPv6u1HkHjmEpTZMidznlPJByVhNLXUUXP
l1Oazn/COcBuODLsAVU+iIMGcUoHU3Rj7dPTCERidIyKk2RyU3ArSqv6I1T28Vc7
kz94qqmOuACvOJ656uHWE1/+1cRTHsNPM+80g823yihKhtrE/8KV3AIfFTyMnZ6k
7JPtu/mENuDoacQeklkEZrIDypKudnQL0p7U8O/EQ27LHDp0hAIcHG3icnmblL8G
oTgM84CKay5f009XG05nX7JOBaycunffWj/xlxFVKw0zXwaSoOXGlAg0bCH5nqUx
9dSbU+UcK81HmbpzmJSVTQFVY6YEEcxtO5ECtBgDyK3ns8/yoN/3+BRQ7hS9Y9WY
LGKRknPWRR+8ICUW9CGQbIJSvy8sUFX5In+iId8pLOqWuhTd8THkIMwLdhkBXrtv
MddSOVjPqBXL+ny6IzGFfHxRWBIfdnji7X5Fvdf803y3lHkdMih95nvuwHvv9ong
0gIM9b3gEfvRTw00FqCHoPDeN22RtYeRi4XIIoA/uD63G2eonZdU0xkWaFoN6ZAq
ubnElX18p657XOfiHVcU64g1YkKXD6szYqnl4bsPgXA=
`protect END_PROTECTED
