`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o1GZOeMlnmElgqEDvTBHt78GYnzlvyQJF/ZZlWzSoWwVck8X5l59Kl7fY3QdKyQj
e9YnS/ZMHOglXPvm5dwTD+GM7TwNKqohY61Vy6zvYhQW4qIhrv4sC8HVSX0iap3n
M25qWCWNsmXWDitPdFjiaeENQMp72M84iBuZBgbhEY9qtFErEkomMHkgL0YUmSkx
viWfhWz+PkF8IX9IIf6FplqgfT8jGMyXzAKoHGRYFnwZ3Nhm1VLsvcKBaBo8RjEt
sfSRJC5CzDvAL4xXLtkFzXufVFuiom73nFXJ/BBa3H6YpSrri3FCxLJUBDgTOqXh
RsVnKpXuunGr766h4OCtkeJdrq2gUW9q6ezr5WTcH6sUY9FSmFpNI8IOdhZLAVs/
08V1tzv/yngVG6i3HQCwJWm/lWlWaAkKU6nPDjSeaa0+ZJNuP5WqqnkwerTUPLpC
hStp6aWuN4PrEE8V/FYChIasvqLbUF5ICeVZzSDwBBhVoQDiFKYHaEBYTcbx2IA9
/jsIHgscrvsLZp5Fmzbnzc+PGJW1pxXhEIHerHR/mjPT0eihRlSfWo0At5u42++9
nDiRAJk6sdPfMiFZr51nXmjWnjyM0+ik6wsvaTwIQzLbwF5+fmvOD8ugkU267Bdd
jdVCIexDCoeA0w7QEky/jemNVM+ih3OoQjBbDFv7tvYxbweVcUCMTPQ+XU4mQsXN
Gm8oSXpAcceLgj0fVedhqdo9sSHKCBw37+VA1rNP7MovgcOSBPFsGdptHn1MDvgK
A3bT2esd54fpKLE7ov7/nr07GOzZ+V43Zk8bVzQZj3zWRo5VHP61nfWobsZJxdV1
ugkPsZ5fMFgPruKQQqtjrEcXtn29PrfQtiTToyfyBvv7oFx75Hd5u9IxPFTq/rhO
BH+x7uEJKsJQKbZXpZYm7Tfserp4Cz8YATlSt2JfVyBZN8UnGynQVDOgGHqwPFey
RJhqaAeT+g0zRjRMF94BiSGScqE6tDJOdalB5T+ILdeiX654XoUWNUBtBT6A5AOo
4vb7LiEjyQ1NhN+iLUp900jYo7Ot6zdF8v8pzrU9nyi9nBiLs5nI2mwky5mnAUaP
UpWwaff9TtIJEhNfEMLPFcoH14adU3SGctQMXdNHBM/i34ZpbPyeeO50s78KavEv
bv1dPUdXd7wDrUCZJggGMzY0jhhX0QgVxbs9X5pioGFrAs6vK03q45EvBGUhUeU6
fIKwa774qTIUzcMN/IXGRZwpOAVwBVcuH0o8FchnLxtBvBtPPwBoZe+droxTg7++
qMrDDDnrTeKdfLFVC2nBMNGeZvxFQjxpzVm45E7VDR8zCCLejJhtolfZUvn1mFqd
H2/cxGvgrEcGE5RIc5YBFALOnqX5z2qrHQFhJqjbEBl/MxPXJFXs/TKHFItWajaI
9tMvUfDIZLets272ZZLXf3GsoVT4PUFBIj8Fn8pSlBaTrmAxKcOGU1Lk+H8hZxWk
3AVYFRflOwzc5TxirN3jBBRbPzErHT4YFNpwxgaoQAJi7OrKQ+8YtSne4mpc0FfS
Flg6EAI+Iu3TIW6YxOX1EoUZWMarDRXDBMyYqsZKNk89hLMbvWEwK6E0q8FFRoqb
yZmhdtbfKo0JrhjTwV8gm/nYGWl2UeURwadCvhOeiWvy+/9g/rAa3BshQk2wpP9O
o+SzjJ9I40HfvIq1eckrmpeTyP+IPLH1RX9dR6P1dwUKNQSSgAYr5OYiorjRlcgD
s1GpJUL0krE8KXmamrIinfz2aeVq4i9ZNERiGxF/JG7qB47x7lQrGAPKu2eEzfTM
LVYAWvbtLdwLccKw9jUK0OhBetVjQ5T8A7r7YyF56kONbxvGE+2QrrGCcGPc7wR5
D+yw9IdxZzfGcUYXZRDGjfQQiKXfBBMQhIH8lboj+sfbyriuXgXvRfoFz6urbvTW
8rgVvnzdUZR6HZ0xN7pJkJEYOpBB0qfZ6nWan5Dl6IX8QtsUEsp3RkgyuLxCnuLI
ksBzxoMdNnZiIT2PqousLugX4a9LAO5OKcbYA1YattdNq8SRgcxrv6uEfBw+n3rx
DvWYAlJ6r0mr+wLQ4nB8be1zwLAtJDueh0SvBwBDKUPytbQfZ4+gHXXMwl7d43lN
Arx0rizkFzO6sD/YnaNQ8IjubFtbgQP+yr7XEV21B9WAVfmh3u+CaGRMsByqFlUP
RWUJmxKBcSFWnZD9dJ94aLCZjNIf5oRwyaZ/PH6bqlD5ROOP1PGUOJJIiYCzOZCf
eSCiQZpgpWyEMVLJpWnn/rkGpQRDpWxesygMJXeU18tT96R0lNtHwu/PJQK/En6B
23Es0EbxKOk7go5u/IGrZ/9/BA/cpKjNSe8aWpJC+O9HWrvPgFCB6h3wCPP5G8Ja
wBlXAlwjpaxnYWgjythk0fxJ1B0yQikEfTlNoy5gPO4FcKc5W2I6D4ZT/XcnyCCl
3WNq0KjzZ1zSYscY5jc4mmKVfLaRBbjQSRX5DhlJDORy9UKh4c4+bE6s7pDV5zr1
Jtpg4pbQcPYYz9tlBhW4MFXqSgfAKu90a3lKwrJEZj6CT85V+qVKCjYwSGTv6O/t
CRrkxo+rmJ3sYpk16I1vOFGSQ1YwNiW58EXXXY0ejhUq+cwdv0IF6kgLmVI7Ag2/
+K8N3bHTN4iTwTI5aGRwp7dlLVGMSUl03LkoMwcIgE3fWtNQV0SmF2DmWQNq4Gq9
44gn1ti6wwt205M43A4iInKfZrgifsAWbPn7aep4utzflvy12JAXp+ejhNdcHpgu
m3FWrnFMcFAYZsHAGy5p26eBKLtLy29qMWMDXKI6ckaKRaxnQJbXhx8hE4Cazh61
G8ObDXO4LZ//8RwCwgI7SJRbyL4N4fJ2ZaGLvw9o1TKfYIyijyHCl4VCPns/A98r
W4FbVg/JCZgI2cv5nrKm0xVOAJBqVETHo0zVqhU3P+McZYSqfeKVrgVxZVLYGV7o
iQXlRlZn2CTMT4G9TQOwkr64Sc3UJ3XVH65OjWVSg4UXzJnNvmSSL/giuU1xB6BE
K1raF3zfQaTfpMlGe1q8rmJI5iZ06ByXhhseQqzL+rlZMuSPyLqdiZ1e+UapyMXr
xwa9fzIrz5g3xIXPgdV9/r+xWxF+zeNU6RNcM/7MrUSmPnwXyFS1HYS09vVY9U4D
j4zaxvTSl3NFCHMf65SnswIT04MjZR5GTU+0Duk3iVOftqnOA9Zb6d1szeQnp3vN
h4FCBJ3y1c85Je7Vu7xPi/I+QMfShVWTz/snuvrCkIpLyLa5NkzXMU5dY81qswLu
AIetfFqo5BhFBsUk2BIyBuA3HwKkHDwd5dZVR2JkxxnU3h1u4oJEvZ5cXw13IRkv
ggUi15HkkYptY+KpBxDywIPPGTeWZhPZDoNOwgb+s1aZimudxMKqoNklKU1aXyGi
cJjBgAgEPFWNbViy36nTokt1D1AE16BGphqVIEgDMJxYgDsK1vejb9H5XUOdnZ59
0E9m4Git9KfpU757j03HZoi3YrnVc1XLT6n6WZYOYdDCco27oaTFDH8ohAGzbwNs
LrFV8+7P60oXhe1ouSwa/YJjT+jf3ym57FCP4mWRj+TuBybD7mpzX13wYkvgOv7L
UcHRwhrfiHQ0/6I7WzOjIu7ry9OgoT40BLzDGKMhRpkeXe7MU1O/IzooZxN3PnHo
433o2YitcCR/Eyz5gKbQog==
`protect END_PROTECTED
