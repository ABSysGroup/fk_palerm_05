`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kLVsVQrEz3G+LsAnm2oza9iNm+0rYcFo8Ij7nQsOYpdNv47gGeLxWu/tno7JIwZ9
o4f1LXQCvEi0ZTAzxe4zZg94BYLwy3buYAq1c0OjwK63aLhOzVYOYnrOt2h5L2Og
pOz3wD5NIqDLB5/vI9f5LyTC4Cv3bijPAufe33uxTnwXliU4AfYmsaYkByS+6Ty1
i1fIC3Bjl4y7VsZvWZyEHIboD3vW1echlnV7NCi0GIO07GrCwsWhr5hnWBvqzaUY
3tl27aOe9gSA8rUF2pye4lb2Dk8MAbmACCf0zssyK7xXa7/ADwLGMqw47UQ0/Ssq
PL2XDQeZr6atSdguZWyXIZX/l6jYxZqucBs+Ril/evsVH3FbwDspI0HSeXWyu9k4
9DuU7vxkKtEIoilGu9CcOE+O4MbwQVYQuWaef23bvuM5gPdIAi6wd7vwLhc+IDUc
Xlj6kFakVPQN8M+rsBnbnffu2dUMw84Jp5of5VxVwtosTnfXrqEtlGJvFX+2VIEM
uMUE1lVUICMwUFcsxzrl81WDlbi+NB/W0a6qTbXqzmBpIVNnrO0hYW0sFSutt7ie
azGTi0cV3x5/EVqLDppkS250n4yuXsfwV08996sGSvgMoxk0+3qhncmGwYjS/X9z
7f8873qzMGQhxq5FcrhuFd1jj/9th8LSzngnFH4/HE3v0x78cIpXHeSmzUOAcwNw
xPlq3PaNp0OqqBCG5OOK4VypJArFEXfFnMm/rJ/p/7ZpLKC2nuY94yyGGo4dN4DH
/Tse4A0BeA6PdS/Qplz3iaWSnrD0mcO9xxVLTmDhYJDe/DNsw8wfKMs6OHnB/2h1
QdtfdFhhEM6rWn8lXdKF0OYzCRjsYALVKHfJ7M/JVlEAJnUUvNtC1SppGtwL5oYn
M1TVzPrk2x91XBL+tfy++Y07m/T5OR+2URqQcO9JeO3SDMsJo4DSFzVUPxl1G0eD
+obgSFrwZNpCkVcuQUqOsFofW1fHGcsphvQnvCLvvjUAtniayZdIQwHrEnfMtyH/
`protect END_PROTECTED
