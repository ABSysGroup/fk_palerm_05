`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1XOf9Ad9PxPC3MUBrdkDzm6C8FV1g99pZPOsEMIQQNEjJqVfNj+jI5peeY/RBzgF
Ptq+TJQz+OSNe2SbVLX6KG+EDC+aI+1mbzrupNCnqSeJY5Tg/eKK1Ef1SwjWlaBA
pM30bra/fZY1IcoBwG5IHBhwKsY+Tf6A1MbrjY7f45I8bI/QDVLldpaGrccGbJS4
JL7mcoNCm8lS/IcKqOGbjXe90bXyaGB3GPcnsGkxprxeVaJtKyAXkLOKAdzxTuTV
/0v7c4PCL31ypMn9dGNHfxFJ8KcQNeSWr9Vg7oymgdz2eWyn86xgYU7zBEoqIS7U
2JTXDTLi7kXUYxDX+4PJTB5U7ncodi4+P/7yjN0F6Nv0OEQWCTz/A7W7VSconfqy
fNBfWGgzs3+S7UEsMM9elMgWpAGwdHJDC4IW1PzYh7QuhIxJ7KhwPwY614mgtkVQ
I8+0cYpRFpqZ2BJOsjcK9TtPR+e0WmAZtaQFO7NH5x2L/ceIGaYc7WVYqcRlc+Tr
pQ3X47qn99XGUcc+mpwJ2vq7+L/1D9E7hSwPIVyspKa20mgtT+zgp89A2DGJ5nju
LtfEwV71mdFpMjfHyK30lzgMtWC6BlmjRxWKEiC00S+G5wCMmSOHucRTPOIoBM68
rKRtEuXHFRWrxtJOtyHZ7g==
`protect END_PROTECTED
