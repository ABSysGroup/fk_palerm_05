`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VzObLEMA6cOL4/XOgyCSHeiHKJ5TEJCf1N07SGTkp9ufqNPBpgU062eImQwQSjzv
cNHOwgQjVtDnkA3DfKMxWbtwbQQ5HRZGcF/ackJR4GGFb+7XaZ3p5VdXb/CVfpSn
gj5b5aopYZzahGMFx8qbRo5MLhuUPY2qeseL8VYGHQwDeOOffn550Em0FyfEpBE3
9jDm8exzHAP9tpAnUgLZvA/ewOWawtGj36rgnLZRGK9l507OZw2gMUjG1k/lOvSV
tTw/k310DMa3ryEri3rY3bMGdWDZxYbAIrhJ42tzU+x/KNm0zDEVhaiYUhKNbNZV
fhlgGVG83MvH4vENI/z7veCZtJZA19hxUkrVg8Hle38heseHiC1bqcie5V7+3ctV
7Pj/xy3rTwGy4atRYOgY8qZaE+c9dckH/mHPFRj8e0X5GKCZWl9rDRyUUEpu2PSv
5Gjz91UFHj4AZir/xQtautAxNm0UdcR6Aoy1zfbj2uWjucrF+5T/vcPSdPcm9Zn+
dZThuV70Qi59+SxiyDsB2wA+FkhRzHNv9EfysHNSpUp6zGGv+06IcUnfG/SMSZga
sAtxBif8wjCpScrNVMWYtCk34jdBCrKbgsR0Y5ELXxBbxCqfZIpFxOE6nl24mTLM
1JBQ05paYxsbyG/wr+wLzWtgNOydS8pfq8iyIi0KkDuYXXIYuayYMWbE//ZZZdm2
jxGCNtvHbaXlnT+lcRepKJiL4085jWcCQN0V4rl5iUVrNSyMKeBvrYRMXA9CFkCI
2tKbcN9sOvf83mJWmgsXZrWUNQX4Uzg3R0JkRGet0Q3mvt5Q61XNCnJDOxSybX86
sRiiXzUAbRLQs1KiZgYCrjIolqHKZ+TUveiIRImwpbYsNl2AbxaCbLM39Nos8loe
bp7jNJM+ubkOGYXjM5242GX8V5V9xn0nhAgOAhAqtIphBtsOZRlXaZc6s2ip8csY
1swX5KosnvTImdKo7fpfC1AuJ0Zc7QV/VFJgZq0IGf8ReQneFn3QSMqd7If2BdNt
H1+VJaZ1tF8osXMx2pp/UuyFmYdw0M5qYidsP/RjiC1kNe2UjOKe8dH/2lacYwKO
DXWfOkkltK4HzDvUDmg0WJTEivuOejQzIJjU+HZGH4TiwjrhvM0uWNNKHrLOjkf8
61bm9s2pVsCN89sw+zz0rjsh2W08FFZD6XobndYgBZLpkMq6MWCBf9IYQR6lJoCT
JPeNJVBwrVdm8t2+RxzEXYYmP72FhNHouyPPjHnCjzbjwPu+Tv3Fb2DoWROjrsrV
ZJVcxBZ4M6PZ8UsNOb2XyM3JaY6y642mRi+pjlF5BXuXfluqTHjJNnq1R/7pup3A
YVpG+9qVwMXtGvTe96KBR01HgkuWF/5dxrr71oRmCPEOACYp2Lt/AbJkmB3bCJQG
Z76o77eF6YFwIxGF7nUH15idkl9nOsUM2NWeENgjFqJJTlUWmgsKBS5yRlvGHaaK
21GyJBvgtq/se/mILamvoUOen3mvd6qSgZFLe6WPdzTZ7Om5T+KyofxHqMjiuGzy
6G8JB80L5eini3uW414pW44YgKm/ZGoHlebszUpPIHkNTBWjSTp6z76gaPeGuolb
KMuh+AFbvAqUgF8YEqb7KAmKLOdPyW2xchClwjhFeXtFBU+lNnf/Xg5dQdKXUjNW
6RrkRQ6p8XQczr0aG1xuBzcc2S/ZIEgH5PJlyhzIjI4P2DwYmLfWLLUw4RhVjnjO
kad6+pp37OWOBrfnz5pzfk4q/iKnx5xfvZP60KYR8Qe7oRUuH4PItcAff2CXAK9l
JXQwiONDkrrB+/h5/28ODHNi1mPmz/VaUBk0iE0RwPbTnX3QaKFLaXF1W0BprZrw
lMVAtCbKllKlVF9pGDNE4mZjewK3X3h/TIxC/ue2iJO/HR8qUQbTWxnqfwH6NrZG
8Qj7+39XPW9bHsS0TbPBtAWPmey9rDiOgwmst5HTKf5FzSjDKdrN4dJMHRZtzmaF
+L636GcnrzsuneYr4bhXGWB2hpAGJ9T2HALWcTMsh7qJh3c+hN7vpYqy+hpjAl8Y
MkSrnPUy48oxvoZK7UnDS9V/XvwM2KYTpGamDzZaQr/6oSIkY/V0Z59WZcyYMjMV
4kbedicn7F6Pp0fNwlfOrXuiFUjx3sPCH1W5aYb8Dvk1Pe9rrpNVPg6nvsRnBqE5
0AvlkbAZONf6wwThoypui8ax0D6ppch7EmWhrTV5woixKKfivY6H8eLZEwDgW4nk
9ISZDQX8kmOmy9qVHx/VheWclwTPpWpGd+v7SNz3qpoZ3RI2exwPZ9pems2N2EJy
NFIex7fusBzEa/HLC4voCcUMrBuaOlM335DhYb62sCyLDyL9UijX/2SnkY22ALZQ
cMYnZLe2Y+6+3jBAf6NWudgD1BEwJ2DOi/6iX7zmyaf4vNfbkwlItwEwSDm3CYNT
lmwZ+dI5wAvmpOON+MkkvtrQUhqh7T7SIrMV/zLyCp97SA96lm+n/Xx2Xaw1FRSr
Aok1CUxoyNX0FvX5ZDMHAWMp44cKCDkTC2FM1KV0US5Hbo7HR1anHy+6rrhrpKkT
yec752YaGY3W+DPmyCcdW4JpQEtpgUUWj8VJY2nE4EfjBUJOita2sxS0xePmr8EZ
aXB53/Lh0v/ovs4EAZtQ3YYkKqd/jWIzCpXdmGLf11ig/1GYh3/qB9wmEFxy1GDx
PQUEy3+3nkqQNlkAo3Ag6mtK4obNJkzy2DEY7Q7lXpzadywWERmK3hdZMk79sVVo
Xtfip2+mnPzLvJCWPF+KM1XBqvZDvEaco+kY4SJiJcWtljYeuP1DUFgDY/+z3kg0
V2YftpuN6Ll4kvBkMWGR71Y68Is/Pcny8oLFt7jCohkbgT/VrtmKCNPevuKdwZrp
/h/Ls3ujttelLv+tW2MFGr3EJDC/VFiKPLwqAR3qZWz/BK0FTLJYRKjk3R+nW7Vr
t2cslwtNOnwQOzdC5b3Hhy7vPnosW8gaMaeuqhYif9krocd++1FlQdbQCIAjLNQD
a0ciheFZmQfTtePLb6KGZyPLnGOPJJc/eDhn5UkHiD5UCwT5W0v/JfR5O6ZH9h1o
ggRUZjJwESCck9cHq380FeI6U7u4lTAQsGYqG1g+2X6X5vK+pv4af30ls/8KheDc
Uu2aOXm16U41MEx5RMRcjRAwvjsQhlsGWDxkuQ6OZbGNVi1RGtXllpLi1J/okf4E
npt451eiPX8pMMiPSS6A50JKIvCf43L4oNY+N06KB9szxjpQA+Y5czH/C3QBIRzn
ag/DoAOexbDpteUpZ7/rl922blPS1aiSK5G7oMJa4GvF7tOdKwzsSPOlydJIWy32
UJ1Rm3vvhkQS4FJNtVl+Y+iZ2cCl+xlAaBqgrUL2+g+x6qNW/9MloCzK6hrhOPT2
MK/6MYJWgMdTFmbvOwkUjIF9UaSBF8lnzMSlr/GbHpDmgeZs4lUef37XofI1mBkd
dLveuiro35r8nQ1thu42D3BA56eY/DDdunoihs31AVLG63vunHHOdG8G26ucftle
8qQQFbpTzTaVBbtNRYc7SM9eH1vATWoJ0QB136Gmq5VF9l3x11dugj5csaVCU+3C
PN8hOWUN9aqYWbkzR6mVqw1hQVBAS0VjnAuv7aSWEY596VwQdnOqQqDqpo0VSJtP
X9Ve8YnZx2B6DZ2VN82Ux1s43fUbO2pbf+xPb7HsYGdcguUpnxLFWt/a4ofakk5t
/M9oiTilNosASpXxqVoaViTdKefFZ2ibUwKsAW7aLD1qFdfphV9MS8uR3qewGxNr
zzbZYODIAb+8h2Hn8SbXac8J/bSWT1F1w9YdmFBNI1vKvRUJDAaVtGMNMPTChNvu
gtQgcA3uGW3ohh42B/SEhC3YYtsK/kGStHEOZrTqjJOh5CfCOB3XSxYHjG/3HrRi
EMm6HW8ncEUKf8kLPedMqVU9kPoJ7ZcmmVrEtMIApnXAl2ACKIM25tzLpIW/NT9H
6OHm8DDq7qX8MvGmBgDYcPvoAz8FkpfPtj6k4i++qfXbecHaD2RBIkBGo9b6627M
/lVwiy0GyDH0KcW06sBhnmcq/RyX16oDIFb2HAsguS0mqsYE1b0wxAY9yEWSwbFu
xK6nWcb1mXrJgcLfogrYddzzqq4k3GD+Dni3NrCEAfqlYrgNL3B1W5X0M6PXx+nN
LkPBwQxKzrSrxOmVTT+qhzkwdzUGE7YuqbyXE30SNMv3CP+eu6JvOzEBy+i+lxML
Vo8yenzoiCEAoamLvZY48705qMr+a73dPXpR9DWdX/sBSCeqADCfxBzsOqsoLOKF
2r/uX2JjXyIJz4zWDnvOlGCWtLwRJOmJXqE+62eP1Hi+e/SmnBvFqFHmqaVUPq6f
LLw92yJSCD4ii6ETmqidF55B4vPgrSDFvF8W/0+5UHEcTpiC/YzPS4f4otkH+Gse
2+G82qhKMYkPB/r/9VTEiTUL7owskqaA23xXlFLn/w/PLS/pZaO7TG/bQZgPM4lv
B2biZQM13cZ4mvzTCQz897kHP7J2Yabf2dRxHJZsrlG9jd9fpdE9mXosqF1JXJ/q
z/XcTz5V83GpP9vw5o3GYqV2kXjWdqA+PpJQy/KYQ5U8KXNjb1YIrJrUPyK9n5gJ
3w8DWkCPUejUUcP2KYXdn7tkiQ2qkqciH7ZjozXkhXiCZoRYN0ZGv00QKqFTLAU8
Q3OvXa2Pg8M/qXxT/RVOBYg1EUbCgU9wVSRLLezzk0PURTOAO7/B7ezRT8qPauFV
ZAC1Xk+2w8GPCrKIPjozipYdtTmUw/iyzi4/9KbbmOxpzpWznpy6ro6DqfJGtd4o
gfmWpk0tJtdYpXuNStWYvfNnKiwh9n3mbnrfNsN1FQTjwIns58eVQBs0zgLvLcrS
HSLWu62FjRKytly87EyRB/ywDXjIOW+27v2Y1PTgriIPNvjtSOGOlOzGHRCB1L/M
ETo2aPSsTiCBN7D6GERy89ZjtIQ+ha9Tv+jChsg78OKy0tce6M7v9vVojD83O/ra
S8b8wLYJS057ZND7r61m3RuvGtUwdL59eiuvOs2BQivwy+Qo2/U0CSeNpoIlrT8B
yXifYl2PX0w5LB7jiW26j9fXVgzEoqYDoG9xrxL0e4z902225ZcYjTdxcrqH1MCQ
hX/UUKMsYOLgRgGrd51N010yLI7K/OhWfgJszglqL/JQ5NcXWDi2pnGM4waYXMbP
VWNWRuFMOxfRha/LGK8ZrnZWIvsUVHR4+pM5VCqxmd1DNr/K8qiBnYVpacnYiphE
NV/pF+fxZjJx/e1sO3pqX3Xs2DimskbZPxp6qN4eXmiCt9wU5phfs97OuEOrQh2N
6poNbQ79QBZX6wqJ8xxteDBFv9c7pmp/XCh2hoHgSIV8e++BfbTbX7qLKq46NSMi
XjLopsg0H9v7mqV/8vF3alQwCRmWJaN+MC5anihJG2gnM+b1BqpFO0k02eyDBJn3
4shnPzDsx50fmKdRcKjFQVyRR7LDheqVgCXNpT6lZ0FTUkuSTF/L3IVfRxXBR2nj
dPFQOwt2xu3nheBD5bBOfbDEwZ1Xx0J/YVxG2dRTMDGznBfT4E9FIjrtVpIrRDOn
RDEOxK/Hm5eO0xCom1fg4H9HH5CrfPFSI/QT0TmAVtDNBlZ7VdvfpNMXsZnGVSqS
Fw/jwa9bmAkpU3otPLSv3/Irkd6+CJ3alAzmW+9xrPmxBRguRQS5C1646ts0wzqY
d6NKf4Kwx6O6uOR15GQgazH04f25Kuq7sOG7FA5kE68Jqpj1OFeO38PBLwnF8Srq
9Gu5lmwt48WRHSYg0r5aFBR//eiKABM/v9KfV1jwDbTPkwIzlQDCLvXB0mILca/k
ZQkIHIXHNDXTWyiSEVe1tqsdNvB5VywF8iDfE7YqEVJpqK6kNuJ6FhV8kXfPmdT4
thi696exikzeQfGlJhrWrhsl5An4s/AO+KabbrJafQuQpEJOtKhcKursuDYRnhsB
tidPlkknl4LsrgEqaqQgjTChf353AZnMW5vi5SrOg/fooeQ8xEz7Os9S9/ODWx7o
xn4am2G/4hHWnCeiF8dYl3lazEqGbJq12xxbhUe2TvUAOge5u3URjt2rhApmaR2K
yMxcfdGUJuBA5cUN6NAEgi4NGzHCaIjZJ/sjCD2szmZNxqRLTXx7R4QgRlUK7z/w
1t0ihtkfpt2YM+FgI3uWvft2HUjw5Kw601a7aW/Ud412P/45p5K9QcXyccbcJ93z
8q7l5J7Zq1B59tFdT8yAhJ+2WMtVdc15kX6HcIUdMjQbqK/NXrI1io/J8W17D25k
WYdbvAIu2CtB0D45lIMUcgtnzAV1KB3gd7PwoG/6EK6TilAb7UpmRIhs846WjnEl
gGm+Mf842UZIbyh5hvXp5G/UcmxKKOvTkj8c9rTKgqEVa9jt2lCyEjG+MSwpuP6R
f7FMjg1r5aVqze6Fr6ZUAIHiOZ5s5BdWx0rCkHJsyjuQd83jubD2M7dzUa4V3J4E
S7htdjKaEApo6UVZsAR3PBFECqWzBn/r9eZLu1/5PG2wRHkC4zxDfLknWDJhDz0n
nyk6i3TQUp4zWZBam+4NaFWHCaSBmZiBGDi+JjJWkimTgfVas3SG5jsTwBOXWLvP
ul/S+Md8345l7Hmhebecr0K4K858p0uCrr5bju6k6YXNSCS8kmUUGh3sU5nYcuHZ
0Pg5eFj3Lsk3PbKrYvX4YbhradYHBPh7JnP+BKs0YQ5/1TSjjYXXh7pHVnJ0Qq/Y
AQ47ml+fdphDI2zwOUgfR4d7J3RzQ3kTbqkyy9W+whtHBKeeO8vnM9foxgEtVEUW
JF+ZIEWQdO+vRFJiNiM9Xy7sqjhl86hlQNtHNQuvkrcwg/kmlMPLixKx0feBtpqa
JTX3SlXNehrrOhOrw6HtktbAgJVrlAbf9s7x9O4GdeaD0ivLbcR46crNjr8GZsJs
7yl+gI6a4e3vzTdxrbznIlT6vz21jSNTAGHA3dK28e+dtV/zIzPMO6kRZzk0X819
YCpofvMKb/pYcAOl2yyhqLwsvsCAAggC/xV2esLGFvqbD4mfQYYA1Nv3kXFxpDaM
036bLUmuGcW91/VC/tdzt46/1oqVAUSuVdefGQN1kSdMedUvaJ/4+MgOuF2zzRf9
Gd6pRQ2Y4ap3Q1HoDxSUHQ==
`protect END_PROTECTED
