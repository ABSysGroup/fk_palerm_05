`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DiXbcrVTLm6t4iUl820kR2AR4hRsgHEfAIWFJF1v64pjm8qzyMIhiwGMFo/xjMdx
HuzqlOisqNAvuEio2mwbzNr/D58cgxo+04s9JZXFxu2WqONHWd21cmFUhKBlNwpE
ZnFtjiWdy6mbpG8hkDHFpomqfe8DUMlZB4aB/DGdHE+HqLpZmLHzEQ5BASdXp3q3
f5zcLkHnq7jXpQZ8oUaUYjzTgY7p8ghGtWmXidAbnwMpxslGtexzM5qHnsf3r89A
Dq5FgJ1NkjMCetPfi5kA6wUmhxCedXUwT3QJPaY+KKpj4MZLgUDVd0aUBT8u9mvk
oGKL10QVLOxxZddRCYEOQgIsBaVceFGIX8BEWA3/fHEXZA/IoKz9+Nbd2lC2bG3Y
QWZaGBJ4A5S3sXR7eH3Oz1lHr5yv41jUeh67ZktagAvumWMik80tsYEdpuVa86hZ
osAd83k4qDtT6XAwcyrq8putnCKb1OQ0cGFGeMIL9P958N8hhRxFCn7MGFCI/lTs
Wz/V08sHlivoB2cyPMHWdJ2R3aGDJMjwrlyZJHAkdg5cBFXkQDyyZsfYfK0eLQzS
aqzTLiK0OLsqxbY+pXHzZnM6LxNNPoe4e2U1gtd3qUyDjI+NPOQImL5TwIK/lwBg
tj5ShaCbkBmAHNb0G8PfEwROEEps6nf4D1QJoZLRtDYw502fpYBfkyPQA7yOowOT
lSBJ3lxYmiab8JesjwTuH05elox6su4/6ly/lan2rYHKjfUvvFdl4fUtIGIa6nZn
CzGnnPaPFSQug0XVyW1OdwAgxoW+tSW+lbnMoi6XpgN57av3Ejf76lAFG+b4edD2
N+QSBLluMaST7v0NL2x+neXv+RXb9pB/qenoMGfXGuBYd5hxIDZm0slZmDTNvAFS
i8CHAwbvvmKQjQ8wlkuY+A92HBGr8WcD8/j73HI0d8d9Y38dh4FuqXdddb0ZDRNB
rS4VzSA3Cukcfox1UOiMAob9m/rYFzTkTJv9Oyr3+2F+emduCgQp6gsz5eqwyqnG
R7Cf7sCWfCpu8zHnE0xXjNhcGeD+2KSedcXcV7Z7ozmsTib93HffjixkJQ6ZFZWL
K1QJbqPin9rgCtoz/tSxG1TFavFt92QJbS3mLEs68fJ24B6HCaRhrbEPZ6ENJ4s/
0DA63cTOKGdTKXvbmDZfJUc20uBkOq4BIdD9bu6B57DsKyC/cQ2xEjo7T8XYBP8s
PYx4Q6Dz4DIorg7Ej8RtBmNir9AKEBuj4qh2ede3FKwofN2Sohl/Yiv5fhTQZY53
HsqwHrvtplS5jgNli7ZP084qcY35Zu1XF672FTjv8nd1vRdKElpV5F0rp4yWlT/j
7jI3B7TGzqbm1TfCDwFTioutzgSNriAkuPgsD/mji3bs/dQLC+zpamuhF1Cd/pHR
`protect END_PROTECTED
