`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g2UOebG1kP6Q+Lsg43YIqNeESWmLdfOIX1iHluByt+ppKgnfX9METfd5D6I8NvnY
DYkrun5QiF0nhuubKLzhUoaBEUMD8s83cBSeqlxFkQ+UEJmq3A6+i9rO4omD3VPK
dvTaeMfTDd8KZuc5mlAPqyGti1BxYzTbIakvhbrkIyEU37nu/muoCSialauS+uLp
J/89Kd0Pbw7S6lwD465UYEs9YIvRMY/AycqxlRkzv3JgOZp48eSZeoOZi4d6C4xn
ahOxZaYhCArgFZo100H6R8VVQZrUq7hCcUKcYALhNaI4QXFI3Yz8q4DcL4dONA6m
14gIQ9W/Y+U64K9iS1N2URO5KWtVpkrb/wLhQGz7NZGiEk6Rcxh8lzRg8m0xdRVA
bbEDHdzjHc+P7hpJNaJ99OF1wWvUM5IHbIrh/KUwQaKos0cVADXOfsK1isbBZeL6
9XG8U27dJ5k96sXZTgzEL9YL3/QZ5PFXIRBO9//LKtIj3uR7+NxxLztDJlf2+xzM
XJn9ZGTCDFUjrUJP+dl2xj+UHvleuz16DucRiU/4di1ydK0NMbdQbg0TuIVvUoKc
go/DY7T6nzNZ+/Am3Z/LacD3kOmUKhPlQ1fJJjGFSYp4KorLMpVZFQPG+HYdGSSt
YvXbhxqCqWzqZWG3aKzkVWO/9Xtn1zvuCb6r5GGcsmpDIZIETf8N5pFbeipmXdBd
BzTWeTD3E1Zs1CzMhzhZfIBwpXuWkoP3ORM3cybYtirrZzq8uiDsPX4prufpajki
M6eviGR3AML4GE30Xc9K8bUrUN0LAxo3tsDdqyE2vUur99FZD6d++tnJUgFe9tqa
JL2ctTMA4FPDiBPAXX1XGhc/k/rtI2Ydrn4d3/B6DaxyYEGOSqbEDcoAlFN0wTEd
5HXDKNlnth7E5we9hkSkGy6wM+SsqJHcBqz4mOjPrpXVSvvSFghNhnSQ5Dh7ASdf
fo7il9Z1xJe3pBT++XswjdeK6/1zPWo7qPC0PF5b2/LyprAjgc5g4qtYV/3seN+E
OU1m6EtMp99aQcdp7mHMhWeuVFUtyM68QrwGnzyKjQoGTxqGiq7cNqIS5Q/xUCpz
A0wW1oWqWJeInxAGXXFFklmoCSE4OjV/4wILpXQJJ2/JFJ+TApiXqyUzfiIjnXh3
f1FDztWJQ5efm+qs9ACTDJ+ky3KxtkqZx6H7OAFCSa9lhpOH19Nh7PZfDTxz+pOW
mF0rXmP6K9Kda2+vsDN0vAXbeDgRh97THPPGU5KdF/HmKvy/4xn0o7SHR+ZFzS3g
nNuelAexgUZBieqL6P1EZX0VQW7sR0+gGDNwt/6x82HikNLzUvqVIaiGgTc02S9w
L9WXbQd2p9KCa9LFMDrfwIkNmhLZ8QhlbzOYtiJ/wh0BtckZfdrUAOsp/Rndwzni
AzhILrB3FUwML/W4NLg9Ll6I738betygWv0atsOLM+VH3P0wvLrdbAc2YDIiPqli
nk6dYAjv7wD5WywTQ8TV5Z5b1KXpy6X1cSHu3XiS97uMNQhCXE/9uXGN00U85Bc1
JAt8R3gnmvpDlOauZ8+bJAxWTTgf718QzC3+u+owybsI8hmTetdSlc00/9QtSO/6
DotZerGsHNqxUVbAHPAhN+TQhxFJe5io5qvquEjCQZghUBvhD/CdS8qXKEWeFR7a
zkiQdl+wBe665ZXGmBULebJSqNCXjpP5T+b67f+45XO0yetapnbJ6rG4snnsnfUx
YlCpzl8GhXzrcCxg7V9ZMA==
`protect END_PROTECTED
