`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UBbqzwjbek98OAFRpLPRMh6pH6L1zoi0KcbvPSJZa0rs/mT0A0suM02ibIWyp8+8
lIktvXlFq6d8WMmiZUBsy/aKMxbdIIGeJQv1lrqdkRYz8QtMfBRNLn1gMBm5GV5R
wLeHmXc6S9WknmqW8O91ed3ozlAkfNCCTekaTE929+1tULQtVr4XhoIeGNPNElvi
U/IWL6Shnw7d/xZgcj/gPWbNpOy3e7N1lIFFY+IZu9sHZz2UQhQIjDs9TVL/PPfT
i4QT5uGJbYyS63hsNnxYC6TlOUsUrx2B6JXwaR525FqVPt6l7JPk4HS59cJMUpQA
GiRUEnIm4411fzAaFFJaYEP224fZgeyPErfTanYwz9CElvRE5vOdWTdlBy0rN4nm
r5Rz4tXNC6xkXoB9evmMzAk9362f4eTYxgxWUIZuJFgY75ghHtX5QC+dvorMZmWF
uyQq9SC5A1r7Pnl4fsa64EKMiJ0rCMPhmAvnczzo74j6XSxD7M/UYGIpDH531oJj
KXt/VKZhZvqnUa58Ov/r+hoFK54ZlMBbGCPQzz6KZ/UTpsS56j9fIJlLP1WzoWuw
qgi5pga4r0RB39YZrewerGeMPiA1f6jX8fDuNhv8FeSUbw0t+n7MhY5JVRJ4K66Q
0UjhyvqBb05LKdilfKupESMwVJG/ocQVV5cvei1f4tl4PrePK7rwg9t6ELH1a90R
44Yj7v948WHSbVj8g8lA8aPSqPGxcthGUtTjifc81XYWoL/4DOk02ZozKf6e8NSR
8jopfhqaiSkkA8IxjBzZNgcLxFsXSkyNjc+SiUKV/FnHS+j0JFZWd+rBCBInhSuC
NJP9BLNHkowNDj3VaTp5e2U7bsRzdB62ZIk8FwQCmpFuXUewFtEbgfctYi0XNaaQ
pwYjLB24jcIinjF3zrGQuNs00ozhNQE/D1vHEe+BkRNzx1oNJzCs6T4HYAgtnVN8
3YNBwETTEnEhwT2XVulwN0ee78Lvbw7MB+FLcI40Oz7V3Dpf4qK+ZNH/WgWNMZt+
ok8D0Nui+23tc1gHohzDwLgd+7pc7R2IZgcZuosPt/QVa2FDRqNPQL5bLQqKFXqy
ouRe9ibRAKHY+tjJ+578yFpU33bF95O2zvF/LLfL0+hUbCqQpGZFXssfVsVtHTw3
mbwnAIKLooJFf3lmmaRPXIWpxKzyeweQ6DErimZW9Ia0Vg7FHsaaQcezQ+wpuBxj
yKXMuIfqKlVR0Fdy7DQtBUKgrA7BxTyDDX/uFfwLSWeEMtnhDGqlqZK2HNs4mitC
gCKqhJt329BImvYhUM+d2YBudF1RzoLTPm/C8dcQ2sF8rvdAmsT6BOayOilgZDci
BFsru7ZXvLoW5z0PbHoJGnhhDkZ0eNc+KalDC5eGuYM8hVArfUgaXdAU2zKc3NiV
Zf4jHxPxro+XDnJARU3lFJTN51e3O+7piX4Z6F7LKVyEo82bhnHEiDsZqe4xqaTO
9UppdAt6s6zFVAj8eSnTeaVnd+N0wLkBIRqvJsVN8E6V29yobiMI0l9rljpZSyly
oIEQ9QQori8PMdR4HAqCNRMgqUAL/or652YGr7GeurAjWOyCN5wZi646KaFb4xDM
NET+gOpN7agvffOGBqlCj+zOgXcZYZebo7xJW4E9ynNG4JIHL5oEcaL13qWlB+qY
9Q1AOQaxL47U+A6vb8vJSEy+9i/kbW0oaUxSSe5dPK51EpF4U0I2y8OisRk6gShL
K+SKCo2mn4IToMO0ws4RV//LJF2t5BYf8MjY8IooVQIaZHEfYs18Ht5kuxzdwGEp
bxOyrza7YN4ZxyttJTKibEWU0+WGAeCU+FO9LrwTzlws5y8bTrGPDx6JxobKiDvw
9x1jbJ83ejcwU/z5T7S/tNk0ygFrK2PhO2pT3hs9XbDiCyi91t2y5sDVJot9J52d
WjorJiFd//FBukLQZ6+G8Ha+ogyb/iyFdGv/LwKPWKDSVGt4TD2jFb1b2oj33aJC
mgbFVXWtP6ypM3VwiwVIIrxtMJEyKnvIyJTZO/bGxLOBazQn7OPHEAtleAo+7WGa
KZGfiFOr4hKLRE4ANQKSC/Qd+a1r7FQDr9llSr+cmH2xR/HstF8PGM9eMOlo/Jgw
DTWQMjiXw2WicKBxRqS1KLeUvcB2C5awFcRyrTdOmy6a0ekkViE4ulzrydpbQ0NI
e2+ciJGsXww9JNxjdxUMPbgcHdcdcF3LJ8q4bEPfSHub3Z1m638FAFDaIoC5O1ij
pQS6/FHVrbYSYTAd31dmcV0/HpWXieDwCPXhwMmtOvMN3qCWFrWfeGGOtXkYJsB5
PWyL+5HefX43iis7IijD8eQ5uDdNAnyoPZ1Bj6f4KNcr/JN1TblpYWTCVZXRroFk
tqo3jEiRF12uJQpuLue7kNDjGXdv8EVUfRSCf84qHhCm+hK0ti7LJNGnbXICO0Jy
iVWFA2kyN+qCmRVA7CCGFTsiDUe8l4ik3ZRFj1uwJFlHkRDCdzAbnQMpvdC+UoKu
lQ6b0Awx0AOskzcgO/AN+/N040iG9TWqWckPam0xXP4OVODvGDy/hxFC9cYEn9JD
CyimDmgcQgX7YvjjN9C+L1stpcEM0fbWYedyitUgC3IXBUbfiY3uksLKoWet5FCY
NyLomOCzDj8+fDWINch+uOvBAxm0c8IXpkYeimFFGR+Pf4NveUqPKHRxtB2QcdUB
BXf/4nevqZrj1UFGfl0AxcHd368Qr8wB9gB4G5x8gbjcneLzYyQMxMYhWrNhZxOy
iHxMZ2h0qdvGTJaRbyKGjp045NOv91hjFDyzXJlv6p2sJiQ85ji92GGkuxMhSe1O
yZxb6OXgIcyLXyQ5UF2epnczec3erWjNJK4lmoDgITdygfjhz4ZrnH46dcW7m876
GtxPOW14CKO5N6uXMboleLfSUS4Zg2NlFOlhD2CuEJdMeDCqMpjWXzdkzUuN3agg
17PoZaZIFvz956h+GHxV0d1CJRI+fsUD7GxDjiQQI/2ze8d7OiwD63jAVFr8dJ2e
6sk4aV7sZGEAqdGP6TT6itzEKPa6GNuJ5y8PqR9iO/Es9r2cmysnfFuRI3p5kwli
OERMBvBZKF7D8I7I7I72zNdUaFwXxIm7V/Zggf3//tHPWecazWQ/EwlPCqLPaHws
6oQIxHG+J087Ks4bNLn84bes7BRXsWFsCoeDnPc2rXighhnOiAfHdTiQ6b0gTZlh
1oVhY4WKHJmTYekaDVYSzEN7RyBS9BNFz2LkKDjOdToxeCGW4fGd3xWne5HzGQ4b
omV0ervP3Acg1aKDVDHlyQWhLiHjMgoU2S9z3fieVj6IL8Uo0lzBNMhiOiU4hnLk
nMVdkXprwqfad3qQ28j15utuOUlvIwtkB2aRKyAn+T6+Ah1gP7DpOGZUG1htoo5r
sAd1ol7sZs8Bxf/DGFdBJt5t3eSNd8np0I90tqIyn5AkcwVlTNDhVDqpQU19M0ck
MD+I/jo10Y7arkcOwVbiuCMkXfQXGPAkdjam8izy6027a6+xNSF55GZ8DS8VnAWv
N01rvbL5RDqyaTa4GUvjE5HPJEmlKTzdSCds19C0zm/WiQs0PKeRqSHFxD4gR60R
SvkEfQfI5olrOeyHUZ+tJf/XJcPZNbLuYKau2z3XK/VAdZmgieyaCy9su1z3gil4
5wKqwVI5+5DM1Fg7qV9In+QQGojSZ5GMoL2xP7GTGXZWcT6o1kZSrLhhFSZDdAvZ
kVxgmb6UncxEnAqlHsnuVsU34S7XwYEpjFXUxyaeIVx3AVwVBO4d054y5fuR390o
0D6DL9VV/QIZTUbgyQ1i1eJ8wBb9S/PRmxghJay3bGIgT4IwXFXC5EO2wy0vJHjq
fgF9yLn5L+NYwVGi1OMiyCil89jPYci4+pU1BAe+frgELGPHv//1p4+WSMZ3CqJI
2lGPXDlWrT9awpC0773kv+cfnV9oFDKHwJm0MnuYB3zYEU96qtkqJWWSWODgzH91
Kskke2Z4kJwbledHokBRKeOAj6keKWcxcJDeW0g7N9AFZCy5UWtiZOSp1/KUoeyU
0yiwH853TnXEGqKZGoSK94t96Dr8gOgECDsCEIsAlwY3GCx2fnTNYpyy9WPIt2a7
DBIWppRPzZqZj8LuuU6No+2sQjlxbZjAq3kTKxRnUEdinfwhHTb1AmEd927TvSKi
JLKuPjhYmwlt7wt6CjkbDnQtelA4LTp7QUhMEFlsYPbvAPpEWWPmqoZEd/DTduB3
xDXEhevlLLkTX+U8rLG6V1JGUnxx7hH2VmzWlbWMM98QSA/nHvPRUlZm29wXQL95
lt6xELV/is56TMB6KEcA8NitZTbYiqRM+H08tWmkt86Tfvq74ViqlIhZqv1Owq9X
NXEKpBnguwMv609hAVZo8Xq8LSgeOW4w07jVsHWtizkbSM7MRjJEiA/tKozF994j
NdYeW/udUzcag09rCiZztsOyCEnxQZIRnIASsjrolUf9qB1yWabY3Ud3pOiREvDo
C6RjPOXbQ98BpVBZc6/q4Kzq1JbUzNRldjVVpWiiqL7v/NldABfE81o9R8no0L/O
UDYm2BaoflC8NOfiAMDdWI28YKh4kP/dE2RdhS9287jA1qf604fdAkwbCUESja/o
9X3VSicgKORL9tv/dsoPxbaN2BqqvWMs8RYZ5ZYU4maBt7q9Oeiyn2nynYxA4EXX
FCBBltHB0sFa79JBMoxbKfSwcjS4YLwXC7cbo4uLYTapWc/UMjnSF3c/2J6ZP42o
2jI0FmIIntp/fKNJgOxDIH71yH3DMrUARypQjvsKzQTiItgvsSj2qCQg1nS4hFER
L2geO9XXkyjXvHo0PxdGcqLYzjaeQL5KRA7lnqeRjUDxRPSpuaGA5AlQ4CMOxnA/
PDfwDd3zXwMVSDkacdaZEkX7BxYcMYZCcd8NdYwDse724bOw6rp0qXXReDHNwGaP
I8CMyXlqGwDh3Ct8mXQ5cZW1GVQNtTTgKobAUKL8D1razG9aBY2mZqef5Jqr0ZOU
E85+1cOdHPwtYycaGb4/MdzigIv44G1Ig4L37KI+evO2UrxLxTAxjnM/GqYTp5DZ
0AJZcsxE5zsj94bexM+JaU/3LFyj1grpLeijuhH8JvKzMB8jtQ2s0sb1+kVcOc+L
d3OfwRIB/L+JGRWqU9x28wUeMHO+sPJUkKGgVlNvBilkYLVFOWZdoBCve5yi4Jbk
BukeYZ9Yzk++SpURqT5raFqCIdQSRpIGDiWSjBplk7cW0sx5gB05dzxxKjuJJC6I
m+HlEyeHJBzlCBwKqiTeiA3/m/tcZXB1gp9kDKnAAP5ybUeBVR1+6IDbX0kuF2NG
qyGbDJl2Wvh9cX9RQR8mwpV3msKPxq1BstOvzOhiKaiRMSngFZv8JQeBCbSKAem+
BFTmJk/zaqWCtBq3Nh5rqQ==
`protect END_PROTECTED
