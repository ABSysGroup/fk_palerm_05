`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
insh6QKj6m6g3h8XcjealUcJWH26s5lQafWMkkRAqBRSxDRSwhBffHkxY3HBzqg5
4TNpTtT5Q0zz5dbFpcogCh0Uc5wrKUqOMUIk47U6AxRVyjp/GH7olYJts/IXZFz6
aYdt3HSnBbZyv9vK1Qq774qA+5F1H/gTwQrZMQh3CgKku6cd8tpK6B5ocf75qXus
e+QwqdE0AE2qNIhYyKBNakLDuZekp3QOf+vvind5HEj67ysenlCbbOZBVsvxVY9d
cwHZbiJNNSw9UCmqGHUkPhKa5KODbmHvIgdOlBY9scEcdK7DQHS0nM1KnFZ1s3/5
A2UDnkTSrpx+OwBJhIIxOGj8qjwxjFN9aFVLmJfNZe7qLZDfIM8JdJorwut21gzo
1XQP1pRet5AC6ArtnQ1N2pvA7Wo8+8aaZI7RuTNxeigPShwICiJvrPxZvcFDZkJV
gCbTwSWx+tBpvKpIu1Ja8P0Clb+RXMdNfSbnYh5rw/7HDJz2N54r5US5QMG8mKJe
0aD3maGvI9l9J96qYCjPfdVnU0HGeEdZ4KzwEitLaZ3Qv/7rWhykNB8Qa4r41xUZ
LBQWLelXaUlsiu5GNggIuUZhJeASEIgY2ZzDEbaz0W2ByMVciFz1iOx3bh0bD9UO
NCWCJNGLWjl1h7IZODN6L6rbv3LN+YBZY0ZkxkVJ8TJJnFgfe0UEqa/FCzql7dEV
vqtXXxg4io76gQY5lJZv1j7xjAxQfNRFCcUoSLvY+YEl330S9xlMJBlmd3drpnKe
UWffyUaJiUukKNb2Ks4pc80FAoFJGm6MR0nYYIUDvia7tb2GskfD9BOsAtZQvDIN
Bq2RSyhFlTCptQWzsZjlhRM7+SUOUorrMm6h7mBEfCJkk+SYdng6mANoHvoNRMtk
GAClLMprdF9WlSqsFMtM4WHBTO7vPTB35AAN170l4J8bIKzC7xe+M4mSXC8dpuHw
2JNw+VWT9ZZbkRvRUtHZCWo7CWNQA8Km0VHpVv00A6F4LSZVaRvAWrF9hvdyY0cp
CUgA6kaa8DJ/vsMoidBqq6izHqYDC0v6YgCNsYCuvZhJtn5yytSl4bxz5/5GEM+Q
BzlSaTEb1TOxa4UnXCCpqlxZRLBRSIZk+s4gd362vLrjx6XT7IZUFTjQjtZ2XUmA
IUO8+uEu6ptaiRdErfTYEIM3o/EtL8bXKRNC6j8/BVs5+968Q91eynLk5CECZBcO
l5liZEMw0+pdZtlbrl/Mzc4G8OU+3AT7oMlLfe6TcYcwRxdttyfHRMDWT+dfghY9
IFBG0nzvqNl+d7bqOL9063aEEe4bOzbRZtYKuW9PAh+qRH/Zs53e6NxL+1xWNav4
0mBiwJm16+KXqZ2FlS1zYzDQGxa57hTTL8BplIDg1JuGw5oFKvZtA9AsYMdABKBH
/R5ZDJ9SKq22USxf/OpzfyE0+DJqKKGZuCsxgzS4ZQrKs1ji+i4cDa1S3ui8gBDo
N5HxjkUDQvCcgziOkvdvt1Bxp6lMeZ8WzvKSaUii8VjGyhKYEwHuueB658gpoDHL
W8x6dtKQvjGmljWbvR5BXhTysnht+pWuL6EcGjfg6BgbayQRBi4hcA38yVSGdyZZ
+PisusnsxaFaZVU1Ry6Nvbr22qLuj9914s0U72YaTOF34FmDGxe1ux5emrmNfiLu
qjw1T01fN0Z3b2c3StMsIF6trSadXgoEtpULwpRyj6AR3gHNCT1TEDPlS1mTPI7R
irS0k4Q9ScWsMSvRH2WrnG5eIA2uGALpWJ5htTGGG64dcBn/6YFnuF7y1hY0KQp+
spDLGNB8u8R8rpCCgbp37+vVDPvey4LMw8HUpio3iYu3an5ojBDCl7jlXlj7vHtY
EkiJV4PkzxM1174pgKXIgxZ4mdIPvlLXZtqQM8G7gCcBjveP9NsH8cpoVQaOiQoI
PFBriM2yzs1UrF1oWJiP39DP4vnLa7ueKXrxr1QtyW6/NHuHuNXIuSTEnOdK3vLi
w/u66MDnMRqZRrpZqqw4M6zvZXAHstdNtVWLikVvMZxaQyAsUjhMG/vEI9d3KmTx
4FCbmVtVS3Klcs7Jx/PxkrVzhoXgElSKj7MUO4Rxtw48cLkoLk+CIvVP0NShhgXt
ujmoRZg28dlt08dVMaSNT7XOY0vi2SEkmvueYFMAcWoTYn0lv03cixI5ecEUCFRd
RK/n14kOrUsoPOdLjVRccVLbHnXrUMSriwAtBZktWPatp/iocxAPogP+fCkGkb7l
+gt0M03ZWLuUfIYtlnjON58PyWROgtFPaz27GrMIZOoowuOfeHKlqRF19ZHODo2G
bd+sOGkK4kxvjS+QTcL9MiI2Ke78Yv5EHSjkeVf5wvtvmnX8MClPJ6V1XT9nVqcR
KVEstS0JqjVM6DvxVuf449dekU6A27sPmbjHIMKHIxeqgL7rx8mji14lpeUvfUSh
GDpFgcy5rEBz0DBTT7azowNR8Wwt6N8oNlVWt8eTHa8W294P2eYIrgjwPpWHJniy
49gezQXQKZ/VNcEHH/llHHIlHASVkSV//q54Uv0hkzwTw9c/I2plNzq4UUGPliIc
iBDz/emzywFykyAfx/Zg6Q8+ogBe6Df07ZHsVVn17tivgsBdsWQhvDlqa2hN9SMp
qmwFbJlJtghzpsrZyM7KxYb38YooLSdRnlctzKSISuN160TqjbZhy5THucd7X1e7
Cxj17u7WHvxTkNIEoC4ax+M/RhMROYJFKfgrLdRgjvLNizAv5apkmwFof3uF+OlJ
9hhSY8Om7DKNDKZx6AsLRfTQvZSKv0CuEtVEXJ7vIboQ6TT66MGj+HR1fgu4XNgs
SY1OjoYsdgHGUWQ9Jhn7eze4hsBdS4AWgNAin/wwFsVW+SNgKPkLkN+Hh/y+yX/2
mzUkfNYYK8jbXmua0FbduOWXK1XvSD1BHBHnSddhY69IdnmS/N39B5+WjAGtcL2T
0MuTFnjNyfdMBXzqRTdtO5m0z5fD7RWsHrl79BTgYguN8fuTYwU2YjlWy2y++MmJ
Euuq9uJ0N3XSfhgP0E3HIlSyqASMdNXJUs163gG+ecL2FaeL6uVwdzzxVUavSzrL
DoWK3biexEc4wMN9oQgoGj6ESt3qDrss9Yq2PwPS9BSKk7SzTzwQvcbnZZsmc9D6
Q6VASuGLFnVjbcazvFYVeNK0TgH+KooZZBzZpkS5zXAz/HFZfGajDXxk5f0aO1Rk
nDQEToPhTKyH3gzet4Gdi8AQtGwopQ6iee6wNzVf8DLFeuABGnnNqCaeVqA4OCl1
H7Vdli1EX+zjQxKj9pspglV4qdynEjtObWNivLGNDub6UxQ7KwaVX3551eM69JK4
x0ne0Km4wJD9Kog+nxGrxP8Q1ZjlE9MHx5GWQ7tVstcLQgF3oaocE6jpjVUT50yA
cj1Nxp4n648JuZ+gg5bjwGZ/9sYR2u1IfRhdVGTQzwQNnkVSyG3GGELxUYCBEuW/
kUGOYEdqTtmNz8Zlk6eIM86KBPOPf1uEdnit4CYehSo=
`protect END_PROTECTED
