`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pwyWsHnmvIREZZM3U/Boz4LRBxwGXI5QtkdMCvjGZlDtePgwW0YRo1L/+Uqz41JT
pV2h5oY93xHrSyOJm/9t5Nwnkvpbqex2o55GW+DuJQpGaiQ4ErABb6FyMg1ZpmzZ
bLlXFLrQj3zvfeC19pWkqIm0GmwKKzFtdxFyTNUBUljFslCcasqYs4dysV77x8uI
OCThQs8Icejzi9cqX619gcJJLWo7PTcXhUAmFw1jKBqMMTjpQOlODbubsiaUHDP6
FH8upZ/k0/yAcUbJMvUYFpd9o9Zgq1WMyLN2KLLGEjlCci3rm9MvWWi0Xkk3p705
a3wmBumM688oPqoAo+4EUw==
`protect END_PROTECTED
