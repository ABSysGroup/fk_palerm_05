`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fRWTP2xCvDv2XUwvKz1EULy+cPTVWNovD8gTvSOKLHtSg4QY8mmLUZg+4LJF41iy
H8bFLbWqx3mQICafoibHLVbb9qbQZ9Lu53g+R5EkYeKjgnFZvBzXPXzMS8JN6yIH
Ur5jf3q4QivrCHB7peBiTv68N4fY0i3m5ct/ruPjXbsQ538X16qgZSH84cit0Ts7
bUrn+6f7bLp+eZCHlLrN3tZpnqVkIimBx+Tky7way5nksPLAeNTN80KJgB4FYW9m
4XtIFbJfwCTHtxmldgM/W0UGlPC1JuZNdgNgbvBli1vCEtNN4LbgSySwoxD6tM/F
CTBg1bHjxHIvn9lSEz5bQPukb4IecbWgSsnZ54pQVzQXDkXdOsr5vdAIR/9giveO
JVXIN6eHypEFnUbYpJMqd0mLheH5wb/vSx6c5F9LpfeJlkWxAgC3as3Wk8PhIrMe
`protect END_PROTECTED
