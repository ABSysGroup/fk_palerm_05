`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RMRhWJ7FzF3+uTQBKdq8XOLHqU+JBeeGcFoWqgpUlAUMEXBc7sGUyueAyo88ZHdf
w+cm7q64jt4w+FWF9Ulhysta/BT5NiIUVfY9vjzj+1eavsyq1pMZMdDPUvKujqI+
3tUcZfVqVznoYJ4hoIuzy/Ge/fjr+7VDzs92PDOgqMOxBmMTiPqA0I0Z2ONbb6vy
zDhYO43gL2YqB+9IEDefyEgVt0OAKj1yxewazupogAC9G8IqK3IyYBIgmQz6JXad
B5yYCCw91pyFdtCHKri3wcro9jelbsXJ6VHyoborJTnbjdljS0D7R8VZ65O0UE3o
6jVf3T+a+I+dj5Ucup6YX94MrX3vTlMIHEsacQpv6/6XphINz0WEU3zv8MMmh7TX
xBWNQpwGVsntfNCskzlzi/nFHXeCfX9RY3slKieIYwVeLJy0sQLRTV0JoWVxHxu5
mksRdczgU8mk1Zrb3XFWsz3/gY4VXZkFZWINMfQtNKYf1hMQX3s7oBUNr+oIerDx
APrT5vQN5El16287cUKttmG1UwAmLtAofl/HoQFNJdmDlopLBBzhvvMNd45k5i+x
vDBe1T89fVB/mOIVZYyH1iYoEsmibWKA49qLkg7PTpGCEbhr/Y7WS4BvYXocH9kn
dlqq7rZHdQb30CuLQeqHKUv8wEUJNS5GWQhyB1uTFe0TQiELgsWqdf7+jpF4z7U7
4Ov7k2FDsriThy/XOZ3MDGJVdNZ/fRCz0i6fjbT5dR2LdxfQFVio9/vNQwGn4dT6
8Dbg801uheV4bZnMf6TNZg==
`protect END_PROTECTED
