`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jK/r+2rtFAU7o0MFphJWnCBO1jvQhNJzEX1PkMFwY8ZMZOomeVkyZbKB8xo+5oPC
DDskiZKwgxfrsvjfklG8etFaHwzvb3/Xqgdj2K9LtR9jaegak3O3zxxjRoMw0Osd
igDpvKzcJZrr2sFe0qpQj/F/FvnXhU3BMqCqfestKbf0f6Dcz0JSXF1VBCzY9lKo
VGCpyaJswP7mWgunec2ZDxSRFSYAG68ckjOQo5Fm9LL6VQ14CTiX06v50Xehy7Vy
vjUdh/drUC32gdAJFyU1oZPJxvqrRHu9V/ItImmyx+M=
`protect END_PROTECTED
