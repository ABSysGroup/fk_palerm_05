`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N/V+lhkMPrTBwTPtX5JoW8w8JjiEhlw7xV/wqXjgCqAv0W8SEa/qWe3rWGYAKO7L
Y2D1OE41vzK7YIxGY0JQDBr8UM2mg7L/gxS/acNIh2HvCHTa6bVcvs3tMCNEVS8M
dtuAyzhg43/K1ttFatk9EMoj5NS6VUSyfNaiHX7kqhpZa4Vbn3FPEcpYSIolZi7c
wMGu7YvaI4xstnocFIm3X3o7Ohxu62tqPGUeOH8m5/ud1lrGYg7VZ1O2EnnaF3G8
7f0Mh65qqVDxgppI0p2g1gpm0X7zwVKahabLrKcm8QPXUJT2W4i79fS2wOdXY4nS
AXWI6w816Hcg/NrpYrLbHK+kDsmbLsqtGX24Ai4FnNjc7Py42rdImk/1E3nBvx8F
WEiZ1PY9E9l/7LPf0KTz3SSgOZevOiQGf85KLWL9P29iZ7eiFYcL76ZxafuG+L5+
`protect END_PROTECTED
