`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kHqFC4p7EHi/jbmOoknXIBLXzx/81qOk+AmUxKdxwEHwd1Ct3WMZz3kyw/kZy2az
hk4PaKJxQGz5WBOKzsPGD09JnZgrrGlxK17/BHeONMJukEY+WzmVygS0vAu82KWc
AzuZmSNwZuoKGKMTzw2vDiYEneH81qqA0zRDYo+Q+am0yxPQdp+KoNZ0WawmLpF0
wromYeLaRE2MSfuR1s9Uw/j4zVG5ZBs6xH2s+EC+4kDIchJv9eRmQ1z4Nj5Im4r0
x0ZFpk3xQbZ/jcCNLNMOfQ==
`protect END_PROTECTED
