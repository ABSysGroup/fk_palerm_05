`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gmq51n51LmwUVdFbdKxw7B8ynQBjXXB/2M2bZcBcP5Qb+Imsf9zyKv6NU9BuWwog
6E7Ndz2pBOYKLtg2V0vGVNhx7oRAfGCTKnl5Us7E1HsIS98C4RrtrbZQh+ZnV55r
sXKI+i++LuDutwb/Z1OUGgg3DqDEFRcqjcxRxoYc9OY5F+fMu987HmXOf6keB+ha
umRNZIZxJvwgVQ0Y6eeGmyI6gK1NO/ZnmKE40x1pIOjD/aigffgqj+dkRRjmFddz
16ZviZfr5kyTJjF/wIeTtPHjGwnD0+pNqFjwCmkilIPFZu/+BB/M150nWqc0kN8s
J0Utcv5LbNHheqxn/yvsAOHk5QkPDnRTqEEC1lMudW5XPXdUBa0kuAcDNAIdisNb
4lA0Hvk5Kw7IcNoPaUQmwJa04OC2mVy0UOsimiX0QfMkRgbKPx0EEIpphsTaw3Yl
NG86ono8oJwOYUrZplCRsw==
`protect END_PROTECTED
