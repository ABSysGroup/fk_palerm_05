`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w4Nhf/+tcxvBZFULpi9SDN0SAUV005eW//pyAwSqLZMQoKyI5uJriUkdWasU2gX/
dbOgijUkk9PP7wTE0HE3B8Zx67tXIY65ZhbfCYGGzg/eMntOP1tvlkegWILnVKXo
KET3oqv+6HR8S4ae4Ia5bR1SKIKZj5pzIHf259YZYRo0Q/u50KgSTmI50GvlVu+K
EK4VtfYQcFOYamrBEG1fwyUwWvjYBEq4Qcjy58Fb2HLLqY8vPgVfyblw9ENQyWP3
BHl+WxkPEN3TRXdFjuCXA2ecsjJCBoMxUQnPsSoUZeDkSKczzh3p2V02Fh+3p5LV
KfIjVsMiOWeAyzaLcp0E6gmpY/AUG4zWKGc2NqSCi6/nz7ShW04GGgkypWDnnvlf
c/wcNbepdpYVkJaqjkdieZh47vWfDk9apL+/KlKufp5gLS0BQQD8Y/jHIXBWO9ZF
xJkfMpa0A6sMXMPyKzPKwC4EyPvaEVoO3IQe0pCJx1+dheDC4DZ7quhijNqpZTqF
w+X0gtR4naf6M83ZE/i/Pyhi1VJaBg1s3mb8nbGDOSOYnZGJDKecS+JHyIWGuFUc
w1Utua3dirrhYJWBsXhRKGAide72YyDbcghYE8uvInt01ZfhP5FyDeSKOhaRutcK
Ar+4Z4ndrYn5ZLM0x4fm0Kbur5ov+GWGXC7N40CBImUwVUOqmAF8ZsuqOyrUJm7z
/CQDL1Lul9ak8MuKDNEMTJT7axcIi11Pp9G+54cyZRWqUw4iNX9/QhpVZJx0QTRw
SM2RY+tqz36pWufNmNCbHnkyVH/KFSP5+v8h6CTbgkaNAW/sFgM9qlXw1d1X9kC/
7isCcT4/43exia9wo6RA3669WtQt/pAqcAdS82kTbisCwLHJopFKJERYSfLDWyV7
2waYza8vRdgq9d97wto/yxaSD4Q4x30EJ3547N3DtTSyBlUXAMRTKXnA4niudoDx
jKVt8Oiwb6MfQl4xvFq5+q2IMWiBbUxnLYf2q1meEOwsjJImwAUwqeoKPdmyTjhc
+SBpZtMuz9glcESYlCwa+Ob4lvF2fzeocVKhvO7YTXCBVW0j0dvrdJ8gjJtnvGtR
QIAt+fsRBsGl4bxAEN25xh0irHUwTotUpZ6RexScpqMbi6s1hvRKbBrTDGk3QUDt
bCM3y+2wxuXQpg+X9RIdaMnCkhBPaa1zwvjBKmE9mOkzlm1H5SrvVxexpA4yHqrR
RFBOPzYP+qTkDr42AX3AupgDP7wd2TV/ANIMqjcXfpY/IK9e9jp+S4vkNWc2e6VL
9xuTaEMiEg8yNJQi9JUdQ8qlvHnWFpV31cGuPOw4fUV6NdoOaX61YxHOFVtDez7t
kDBYIQlDEln4+sXN+QQi7Yhoo+3tW0+2gIkvgfKowt0dY0ijzMZqh+J8nRh74xeg
Gqvkqq6Etaat7k/2UPr0SpBJUSLJ4Y61m0dhXXa7MoWNSz+dV9xhKoTOqtIwryf9
IWN+HSuFlXHcyWJdTbpTYF/5+P6ZYs0as7dmLXN2IYC0Q0VT0dE7pFcnIJl+aIqs
JwVasT6cTAU1FQlAdTTbSAK13fNgjWLCJ1w61vZcJnYERXPLuhtuCW83hr9uW73r
UmgC5d7Aqxy92Gf7XEjgzdDAjsk/aFUVDCt7EJ+yw4lFfvFPxkHnfMXLFnfetzg0
ke23ivJ5gTGDP/eV7/5yko3Lg0fj41LvNkHiJYquCT3KXwwnLZ2A3G8bKZdcZVFq
nE0i1qFjNO39FW8/d919hMqipDMgzJF300ruhqyJLDMfrkWunjJ+9gSsGMV1EtDo
yhasLoOYDeZIuuqJRenaqozeC+wsPlnySdfvcwU2R3LGOJhJHJoBgUFWtWYncZDb
yhSYpLbvj+4kpWjVYnEL5P5WEdXuQfnfdyWGwb4bZ1K4ywMX1+Pn5r7436KNk/Vo
6miuWxal/BbVDL1voKEkJSNstgYZ5F1yyVTF1MdITPdiPqZQ2XoZCT6fNrqfqS9C
ULCCXh+Bxm/wlpvjPc8I/dXioPrpoKHPAHP3pdkQCRjMswZFlBp2uG3j2f7VdCkA
IuY9SCjxgeOcvQ33HypZXBp6l/vyLZ4bEeoZ5Aft68Lh52RZH9udozOu7AfovA01
iZbuNRReIeiLSd7E1S2nEFKfsGsyQ2TjZCNyxWKXmwLvhbVt3yTGnKN1pI1UgNrU
XKgZqH0rYhvl+hfp8oIf5AZvRICb+l7z0Q+gKcHk/SyEyjX6oh3xZaMgWaJhhbq4
tZCjRX5lr0iVHGP/DepZ6cyRkSNagIBpeXkm7FBJX3Px5ZJ41e1XVdzSXMgAlMlW
eBUpKYIo2zgPyOm3AWOi1LL6wP79PQH7OgbzVlwK7Nk/KWMG98V1DrCDEgEHwhmu
ja4JDnABuzwvsEp+hQY7G2O7A3O9AN46NNPSw3vQ/Z+PYwMNC7V/SXmuzyTeQ7Ll
wOtpA2U8pbg7muOL/AWN5JF8EriB/jkeBMi5EYBjpcAFBAC7wYVzc0wZyYxOTj1q
6l8tALv3MDQNsi5Cmj5ErXtpQgZinL+BaF58orKqB03ygQ67oT8mpCn5iUOskZ8C
PjjVwLiVjtb6XRHDIHW3zf1Wcul2mbr+ShFsA6eo+86EDbfpon7YDcK4BXyGssKf
QT0mb/peMaGQSmFtNgbieT2eDJB1lo+GMOBrUjiqRKJnz7EMlFpra+r+J2fF2CqO
Wwk7H8PR+T2H9vqIcxZezm3j122fO79e62nC0q/xmBoCR4X0yfj2k+wxHD6fIYFg
xHDN8WOKRW9DsTXDHbvAbPMudhbPnrERe/7iMOAMfbFnJ5BDpH92ChAkA5KwX1Ym
s1ZNTfAQkZSaLJpIEPOKIqdvcCfiJF2ZXr2+XzJGLdUMsnCl9cKnoECrcWacrIap
L/jJEoUvA+noOQSFq1qD2rt+xO7A4cToxmPHwj1338+dSg5ccJC/rG9T/zC2oeqC
xSRMNFb02lwZIK/MORRwRGOdSpAY9aQsd2Q1nrtdLMUC9KAIv++tp+iuWJ48GEMT
T5TpiBpSW99/2PtGsPTqw3XJOjlMYvfQ6wC6moP3MWo/66znHXO2BcJWSlXrPq76
hGQFhrhRiGsBjpn+gTSZhh07JBoWLLnkncDYCamYtvSD+ujOIIehFwNMo6dzYnK+
OyuN5UsPXsdWTZpeleXYDAv1hl9T80elzEIdzIkGaj4sb4NRKFFDZcvja7rvvauh
eOFkFaV1CwFQ2yKINxTOv5AOWOLAG3Ciy78H9X5a7CFS4R9cGIvKOy/tuDm0zJj6
rIBsxsJJrZk7ufMYHH1bOWex45JS2WK0yAthBYtENVCOPChRPnYcAjtIDqjImJdN
Nviy+rNqVS5M2Xem6kGbmIF6Jg68K+fTScY8aNY6hUdq8UkE0R9fET5Hs3mUQ0v/
pGoS1Y4YayKRIuB6rKNvmzb8vir6qg2mTiMpcn/GLfrGtqy+gX2xKt0Do5jwyLUJ
1tZkXnTtQhn8vahg/yeL5WsmY19TQlhXnddWLPxnnJwlPLIlB3w67rsg+o/PZfJ5
l5wQPymkPkPnOmrBjyzyzw42tXKxxJ3iyZECHwll274OL6fmpqysEo/TKbj4QbH4
td0hsj4Ey5G1p/21+yMJB8p7mV3nRyxV6twXreFRtRmEey4pstKzmZB0wcAj7ga1
Gf7EZNwhvwkzSc7nhaXICxaa5snWhAbSDPCa9JR8bqWLiwHm4OqH+rWsIMOJJxd1
igx7EEwLnXjipC0AGW59hi8AQuhNXDbyIyP7cQFZii4DkT7Gsqrhludxr6I80PEs
hWx4sWChsoosctavMeuhe2MPknBju/yL3t3KDpDgUesQV/0xvP7AH9Mjgt4+M63v
yacJVcaYE+eVD3nFudAyiq4Wpd3iL2OtVd2rGMQ4BrFTd1A/rID9L7VEa0CjvTbP
NKRSJ7VSBh80u036CiHWTRl5XcUaEDdFhlhoD70/Jt+1+8sQApZ4idnRZHBlyR9e
ip0zXM69AajCa9lYCTMLNsjD0Y8K2rbneCknuqTdvCgw6WbtLrZU/5gSsWIJIvu8
v6O6JxupnIWmsdoo9owTzeCW8o92P0egNMuHwg14azI/qWkNt+IUFJlSkmI/O3sI
8tdxAQtjNkPww/mGGqWW1IL+CoZ0DCZdLE0Mvs/0kZu7bcFmcZzL94YKscYNkQNS
DV5XpcqzgD/B81ubpLXU4VWSfqdXw2eh2kk+UToTZyAEjX+/+t9cY0HJFm+6w+cQ
iMPnY16yY6vfYh5JIv/jyOdDGAhZIi7xV9Fm67OnpkjhwP+JweyeL/26W6j2lKiy
kqK6SMD0BvY84zF1B4x+l4LI3IIRpaPXt+Fn6IORGEznOT2MKoSXeDPBKRjYTn2c
ZMlEUK1C2qbuirI3eL/GhKEUNnRWenvQMvKqQ/RQIrQOVmxoZDU9vNx6ZOcLQ/bW
+MxSVYIwORn8k657P+wqSd4366Sox4ppM0mwtili4oVtqeWYVP5CixcyiavpM7fJ
Iy/H3D2JM25/00qasyWERxfbCqM6WP1RS1A06WHUny43ufBsRXBSO38ZYZRqj0ia
7Snu7z1H8jpa9Wf2mizjiELQzemZ49dVQqYKJgH1OfeAb4GCIERuuI5VW3T6JvYl
0CcwITpi5nYhtG4WUD2gVt6aMM1gtLJ8SMX9OJCSxjcz/dUPJejqjx7l0yziygN8
6JGj62hyPL1swpB1h2g4v0dt4cZ+K9Yuse44/tpx7I1I9cNFjuYkotSZkSdd8Bcj
oK8B6Dhc13EVXsdP+sG1CbwEjS00rUWLZBEh8FTERbRyztUsEtJh42wYGjlAEWnN
qOjWFqyGKI003EdZ3rkKN5YwNIxscpKdO4OTLimyxb2LdH9FbuueCoGoUcio0VxE
XyB/PZkDAN0//rwa81NZoAcIpO1SuKnzuEpxXvi8K92Dcx1xASMMC+pOc0i9V1xR
kZpsIVrFjqjF8y8/2E99IDtVlHHayeXFkaNyRwHRwGJDj/ZwRMMgaFsHu6FVpmc0
LM3T8WZi309AOm0k/QO731C21UGH0zF8+0M2rrW0/QzXACFDovXE3+HaWliTtLaN
ec6O9FO1ma554mP7IDAkBHL56gRGc/srL9fAx0n/n6OvE+XWVgTWwRSRg43U3ATh
sq7f3L8ZIHN+35LCLjgWeBxqGGNrn+SGghH627yku5TTJWJXMiCl+zggnBAfqEfp
72p86S/I2gxNcA2Hgszh6vwm0csqEYYFp7thb9S00evLfeeQsDkreIvLZ3OIEi8A
O9xWH5p2TyfWdVTZY7zqVaYX1cHrgk5mroepyuwnW1QKzpZBYKfNKUlv+jZDJiEo
J8vMTkwjXuqny+uKjojmjNVrxENDYZI3rAJ8pq6HZMNLEmGfjdNGYyomEKhrGkJV
ZJlO+RLnoozClg/ZoGm8ywX6aw9iFwBZV5dBLx0YhkkALZDPsV2yrD3aLrCyqRO3
5is4tdMPVuLwD0leHvu8ISJ3/CV9sgqKwzC+hOHgxPf5gy1UkfvJVBUkpoE6zirp
3wTFR/+BC7Gwg3FJK2mPYD4tFQP1+KILrGx/A641ZABF9V1fLGmitWpoT7Roc08v
K1AZl0v4QFTn+zXSGejKlOF2aO0yCEGTefF8GFip3FAfqZ1YnMXUu6XcukYB7KHJ
HheGdYGa6yrv9RfftZ8QPM5bURIjzfJY3WygDmNQ+x9lsdmRyj4x9IoKajobBQK6
yZrWtuJgZSYuioap0NmbCT3Bos8aliRBA4eiuW1cDh6V78qDIjiDqaNtuVFEHxpP
ADlOmJBozsMFmdL6BJSG9ulFo5/jdsepAdrREiY8dm55po6yozDsR6mfrPujdOlR
5wg0RTkvkR8Q89aaLU/wQoA7a1paLw+uhNSp2pWQFMeCgJkiBgp1hBT8uj1eQ+aE
eSE/7s1EkqFgl3ChLSswmRnr9+FinmFRyrZnZ076dN82z6McTkzQSGVvxbXeTBDZ
1MiZgd8E83tOw4ET22Wi3hubYaWisZc/t/+TAqM+k5EXOyBzLhzB9FMrRZBXgOuP
BTyLOYfqqsZR4Jkpx+lOo9wkLjgKfEjytEYoHkrP4PTztDNj86Th3NR0F7Dg76Jw
xCUhiA7tsyFlYMH9EEQCveEWVgmmKFewvWAN0dQjV64Mckc19jQxUj/HM7eoyiTH
VfViJhPiyICHLSdkbdeRAnIDDEE9HwAxMktJxNYUGID85+66hIKEsdiAR1/pghX8
B8Fvfu1owr1cGyh7lOOXldkI9q+eHV4zJ+jrOaB3WlZnBex1Augyg3hNLxQ6Poat
6wIlOYeN0sAyyyaUPxUBLzlL+8dRkAsTMox2hwfEJ95L3G4o4el/Pto35Qk1uC0z
0VmmkkApRZNaM7TEjc7gQWlWjxDfoSyewlRTsSMtTTLK+TnPdJ1F00mV8xDVoV44
LNJKKqwB8aNAQy017sDvDOudH1S8pw62sq+wPHgVheSqK7b9fn2rFL9wscRW5jUM
J2spv15SWjvRUTpMeRB9LydhVLAbRSrWzos9NSToMh7Co1KMy+V+8BxD6BnIML+U
Ai5yj1s2DofzDTTkS4l8O7CREZHRsfYOdq+9Lf/x4Jjqt9iV1HSNUePgNvL6zWHl
MtFSBIv5fDB8ErC247iV7+01D7Lt6RgzAHb69EUWzUo3M0yWUIqHCyJKXcVYi/ZO
yucaFCOmQKyi+fL525gKj8DSVB4AenvAuZs8pVCZd3drU/r0JjLNk7aI/nvi7QJe
Bu5gJOT6KCx8zi0w41zeDAhtXlkTdOvjEejmo0yDq+QOhfhvAvTRcUeGheHoQVkq
7MN+8eIpVIOTymAb85e7KaNn1r96xHWYWCtPE0vpT6T+VapsvPBmqQ/JZPs1hPqx
59RLDwqRD0hXks5nl61O0Hy6HdS6t6+emKTmkQJD53rTnUUZmwAVi4RmMiQ7b2FD
/cNcmkIFqWfWSS8dUDpTjsocc+7GB0dbUpJjXcmr52y0eHzIyP1EazxYcN2b+5ne
HqEJliKXFYfrhrZM4hBeyYI/7TvV9Z+0wdkZeh5JB5k+mLDfD4FTiaMKvd14Y372
dCbGCHtE5ICklo5fq0WSaE7oUkSYXSEKf3QlhXwywfcYL8XXm9kZhMShPMtYhqqE
OgioV0fDN4PBiJUWCDaxOA==
`protect END_PROTECTED
