`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PZgCVmaflbhmtJVXlpz2r9HD4YgClnL/qlILwMi7kKekQnBOWw/jTZEYDIsyAl5J
4hcHKQQCWhvm8VKI9EubBI2mempFseunCX19lhOmkrsxA9g/iZe51Q5IP/8t6rh9
09WiOTy2X7xgHEK/PmpIKt2ZrB3nxF1C7JXYVTXadfwEsEXgeoR4Ivn7Ybb1iHy0
4rJcPppd8v/ETG+MGg2cGf/0m8uc7tVzWPmkd8hb3eKofBfcjyjAjGtjQtCLudPY
nv7YREMnqZSXiwGlrRmOpt/5kk2PKGqrBTLPh5hrN2SdDNxT5w69LsJMEbVfaw2c
U8xioR6W/fwtUUI1k4aJNQG+DmruvnVkuzMlmcitKx409AXEiOTIbxkBgG2Gdr0b
V5gMwlcEP7FCHRWGfa3i9UwjRf52G3kou0DUHb0JUtbyWKDmvq+m0JSbYGye+zAw
oUJWuzzZlDRjh7IGQrhd1WnOi+RlQbn7+FsmRV6P6RjE25f8AjSb7VIequfVgO6X
J7hXFsTSCqPd1ueMMTMdAmus4uDy7kqMprZLMW3w0FSV9NjZ3DaO/UGPqceYMS42
8zjeTy4pXtLTkjP81NfJmPcvj1AViEcc7ZxhrkoozJrzKOb3H8FRdZKLgi2tC2Ab
Bc9A2l2HuaCVgEaFm1TNAA==
`protect END_PROTECTED
