`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LKcCsCX7GjbSbkhR98g9u9yX3FGnAGfEIVOUdXp3SLRgJZdcLjx1tquSkC9zJRhZ
CBYq78loyYVMTtF1vl3YQkN2AK4bamJ1FSadTpjm3aMrYpn/eomzZp/z0xKx7p9f
0RIVFX/pilefzzSFER7WqF8kRcBpI+xjB9i3MT2E/0ubE1QNt0PyRMNh6PF0fC8F
P++0FkJFzpOCc+uKd9WXSoa5LMxzHZqY93lVI0FKhSEaLyWwqYuw5unJcizmCkVo
AfxZCkl8Smop1F1/y4TwFfce6XCgW40gJxHCgsWoy+d10PuZ/MMVTP94sxzcbP2G
8qieStOw5Gwi53prZwti9/VhmcpuVRdPwZ/8XZHGS8UFDCPKvJrMtYu1/MNhXGVk
CUowVfTNFA1jDJN3ZwLJSjxVuCs3s9MLPnW8mw39byh90akTeaT2o30rVS+1eQ0H
VOX7Te1jOT+9/UctnpmUUPXKZHB6W8Gu92wwbV23ZCmw55ttY9wo/aPIwDyizkDZ
HGdcegfnTImyuW+0wk/e6WR55rt22PWlZdnlvUBEY2WdAwVv6fSelKpxl3R/KCmj
9LGYJuI6kz3Q82g3KwURlIhlvpgh9Ib54UAytuJedI1tBEkNR4zvuhLgbdHxIdbC
79hDLBMnwhOrzUCLbXPiVK95EbglfsBYTI7S4OtvZIJ9a2KzQEudcqMMIBjJ/6nS
xeTF6L838iDaKXdGFn5RFiAMFdMBfBG7GiEBHDR2DNZp9+g3nghEdDtldvuwyLTW
JOqUL+N/3k8JZykEUsrnVuCwd92ceWZNu86kQAQNKhWDV7SkR3LMhqyHpCEF+ERO
2ujFxEx4YVuafWRqB61SZxyycPMx0WHeoLe6DXJPrWsle3W9cKRjxKoBslSqFk2v
Kvwc9ee3WjbSL11NOeB9YEldqHvg1zHUTLhxoaW3to2tyRGZeppXezo8dIMxWu/a
3zaIkqfdRjnBxci1hU4F8RUmjMVSRVS01PheIiGcyVgSEttBnSU3yXuB9IMoGQRF
/d0vgwb4C5BBak0VwrhpvUH50+Gzx3LcwlDeF9TpY7UKepc9acPQebyx4ToNL0AE
0A2pEQxAqP8fH+9n5fjyroE4T7Qv3L0Ros2U9b+l3KPolH9XrPadLE4IAJIJTsxj
JYBDb4vIq/K/Pp6siDwofm0L08BiJ7ZX+Z0Lx88hOTfd6syw2soyh++XBwMZnGEK
3z9Y0P6w6oBYo8fAhlPfnNm9HrHj6PxHzMEZvR4bYumH6T6DdO/kQf/seyK0xDjt
k/LpFxeNvqyn9VbugNa2JRY9jbOdCutQ52Tv2RCfCFqHWjq3FG9JLPEnDHfT8KcI
Sy5497mEtCadprmK7z1imb2p6UKqBiPj7LjSJ0SseNv6okW8U2TlwWdG1uSek6Vm
JfWhhrDWw5eNqrwrPLEXhBTmAHPuJAONGq/mb7GBuQ5GIPPB4Y4Dydv1RrRj8NEm
6clUg+Xxb8Y3kOepOCdCpRltDUwJcSkl8lsKQMgiuPL87uim1ftMP0Cu8RgZL+gP
KyO4ginFkdBGdP+Iqg1kPMqnIJ73W+BRrIbZySd0vNPqwny6PVqeZYXidd7nRnXd
VrQsD0wLUGAd2KF6wGVdSwxh0swfS1X1X58AmmRGONeu1YFBKgGKzpvs4YNrAupf
KlyheVAFfBvZ39KmqnylndYliSc/8l1zQFC+imlmNmv+U2beRfXJCsmLidx+UKwS
T/ldEL9JxCansVF5C6Z7CbwiXFO8rodKGzID/KQLihhMN+nYHmAr3IvhuWlDe32f
Xs5gxxr3zpjzDV4hGlP/n1Jg6CdWdZBk7lCX1q/k/O7fgbb1k+R5iQs2f+xOd8HB
NpyvOOs4/UC7Gvu+/zQKp3BXFyeVL62zxYd9sgZTnX6DYLQWmwAvundWfPYxecix
QGja/qPC4nWx8vgjIXZEWJ25unjI+OisdJ2AsEEl/C3wKYJmVoMGq1XnG8Aq5/vc
7xxntE0E0tRSVvFIDKRqvaxmgl15a8oHF71VD7zABXxbiReokOc3zxfJ/7DIaK+G
ktn8tepASTeHmTInhkqHPdIZycqHk4VMYAbKwdyvopjJ3ovJpJzxwcQZ7HvFlo7G
C7PQkIj6LZoGa7Jw9e/h18/CiGcMMPg1eADrGHFhyWPzgsYCXjEygIrKFMcD8wPz
1TyE+vXbK0KNT5C7cLCsPLlJYCfDVU0gmbXTTs/Af1k7etgsXor7DwR2DGwu/Ed6
HWs2WHJYjNZ9hcFlhslbJQuFgXPYoT2yqvL6AnHVQphLix/JBwAsq/RaTPdqFp4L
qgtcGbd6Z0uEiwvbYZ6yIOzqS1w6dSNS0CNlZB+LnfZA1hhIWEeU5TLNCtTiEwBv
ISMgqfPXJjrMT/OOQZWjh99SI+4DdBSlaSxU4T2xgIxSfcIe3opDTHYWa2SkaL2L
VtJI6JzKGjTOa70GCxak0oFqVjSbvzz6h292UcCDGWdYCOMX3FL29CRUMrzbh0hZ
Q2HJKrDXMnWfGJ0i6pieFEpodqbt00wHnIBPiOeLtUfSNQJp1yZHMy+/xAXZhPG/
LrjMQkIRd3ryXOQKBYJGcg2GWYLIZjJ4jjYXphJZZ62bDzjgVJdl8s5CqfZ6ENQl
flRDcTFhUeu7cLBj4W5fExTbRlkj2XvsFxQbWey/3aMSXb9dtAfwRgX+f1j/GNhV
pr/ezqCkJeJlKFz2pmGCd1SmgJFFMKQp5U7JDDVvfe+m38/DCMYBrdxLo5mRHoFb
//zuvqsE31RHQbz9/NNXUCL5yrZHJIWG+akYrC8WK49sNVdawn1WjksdLYOJcNUR
he2F+6s3JYnl8CjulIrqgzMxsaFnhhXWuM8a586jqS1addRU8HhGei1PP26uFvT0
/OZz4PKOztMVWDJ93zmKDGpzBWS/xTtiWe8mvFaOujpTVtCvb3lL0WnT8/4AiYx/
PWcA9ZY4O6l88lXfU9hy2gFcev6mI8SfBnez1p9XLlbwCbdeiPe4bcjtLeXt3rIe
VXUSw7PcO+CwUM4OAsTrIQNDGGhHb4tmyj17R3HftmGjmAqPlUem72Vivm1fgWav
HXbVjdY7Ctnwzwn5FtdJ609eMUwCkRorTaf0DorjCWqXAfkqOu0EYKkRGsr+UqjF
JkKFyD1PASgvQ8NGw9eLF+oHaIG739I6Td3DJtie5gMia1jxL0YHGPMy9ts5vNks
F8Q8ifn3SURBtTvEL8R2SEwjeKcVNjD6jhqYEapBMA4ZUGBwjTqCfa04iJk2his3
qqw+YS3KzgDyLeFTrJB8OQDu7iwzPhNMZXoTWjn4irflIdbN8sxd0vEGsiLAprnT
dvviPCAYT+fQ0gaBeLn8yTlRfgbDEvlycOUx6jXSOLaAsn183sLwK4LetULgNy58
z73Lp8xSFhC8zfJzyfGNcrAKnDc7qkOpAE3kCq6nX3bwaP0k7iVqHwAsIuvam3ew
MyIWiJtN6TIpUPXoj6Jq2/ou5cS9cP6kf6mJNG84y3kaqHpoNPbxQiXA8ccsfBaL
ysdX9g9DacN9LjXo4MmJL/HVpmJ41ebUWHdvN0AID7cbfTZzsisgme6vD9zwQ2Mz
k+l0RnvExGAq10pk7yrFLg/xYA9a9U7v6NOgwFjmwNxk1BryEe53WfhfwU/nMrgo
wOq+77jz5Zmi3QN39CHwVLI3sz/dYu+Am9LLOLBpb/vk5/RZJuyAR64X0CaYDXVX
XCOYZKTYyUUPKKlOiRYvWzAad+5XixHHH6yWTPDWMEV9cE4TQlWdgbeQTLvjbsUg
t541oFagdoHpQ6K089PXrbOWxfCFkB8kMtmjwQQmw0J99WdsEd7IfzlPLd+fJ5Kl
DVp+32c/E/rwMDv9KUlofPMr6mj0Md6LwjIOo8LJ2uFeLelkjdnooYpxSjrBsWSl
JJU6y/yyXyHtdltRlWovk0TwgnkVFC2Yin2hTQnByWmWSZZuz4hHow3yHIZUVJq5
8o2Y0fsTyHukrfCCUG+uKYhw6wKtAtXTD3uc4bk3FDxkVdWVSHdyQ+QDVhvyfe6k
DzcXIgt6atII1OQmhm0gem6eEhmqTdYhj9wRyRhhrjW+ue+n9vRv3ypgaEHyWHS+
YCJEHOcQS2XvYmvnfcHvo+KX5cu37xTNpD9d72p0Xmym5Ff4igOo3FddIS+Hnkdj
FHNsJODGFxoZlsmP5qluQDLB0T2eBt9mPT/AbBHGtMW14krp4LNm1V2oJMEoOQxT
zdIOobeqctzUj/RLROprsC5tVBbvcoyYYw87TD9ViIOeJkRqm+9DykS4VZtGDRxQ
9hr6dqBRAgshVq97pujoyjXpwoyoiWUZ2CAgiaYi93W6+xdg+EesbeAQQmyE+FqJ
w6uyidScUMY38kZ9vFGJYsTlzszONfl2+7cX8ZYsdlAAz1Q4j9yzKR00RTFyvR2g
QfR4DIAnXNC2rrm2dJY/7WE1C1mpo7fucIrTsMQ19jhkpBvWFfAaemkilf1xFq9j
vpKQPlbjeHpOhRjw/bbZOgFq35S7TZpYKKOA3TQXHhT+EXbgv9OHHZ2ShAguTUQc
PyN0Ov9LjoWTOIDTRXUrG5xZ1slx8SD3TjNNMkEpZeLe5maUaKEoC/5LPTjYNWVS
Ieldtgv+fbM9Dtk0fMyqNSjvCuAbb/0xhgxqzQe6nF0vnsYz0DfnrhrP3T9xaUql
8rPm53WPEHW9oDXBlS8yyR1UAifhFfnUk6VYaNd8T3DQy5RZG5Y6BMAAE14GdydI
7XteyD7rC+zTFZVsvxKJeXbxvOwNRzKypuaZdY1K73ZzPKNHaGspzhK4q00JZjGO
Guh2Zh4zj/TxeD8rgEcEdP8TPFCoMq1Qbn7iZRJGuCoj+yGe0Nma0KHGR5FH1l8o
wMT2aMq5MBFPvrtfjIlIn7WWbc17lGsN9RTb3ZOXaYNLJGkUFggNn2W7gARybaVB
5xB41FXK7qWetiPExFcBoJ10CaSokOy2PZJrnzEjxnP8vP9pHACthCu/3a1cSdvr
wou91/pk1+3Cfj/yO19e0SCCu9GV1Sh/4pGSJ4mmVC8xb7SnA/xiGpCwU1DOqR1E
7R+Z4lx0q4sKkB0ub3xSaAqbjv2mQJxS0XqPw2EHMPcW6aPun7qlMQ8BB+jvKmWC
cwY5L7xsEBCvDlk8ViKtPOOBYU7SKOgxnHfl1pYz3fYdey0vnxrStX2AInrg0Bey
L0cFcfQ4g1z8cSPaLufEOvAwoQJEHI6un+B0+BSFIIbvqUdliMHQI2SwakoO0Le1
Q6ip5ELXQs7CjJwVlxhoaJqz4pr8FfiUQxkdDO7bI48NBuLwvpVVd+o8XEGFm9qs
bvfeWsJF8/NmEhLznHZqAzmNKCztgGkZIhnj0FvXfdX8qOGQJoIMPyPifQDwX77B
bwMoPeFxr0e/Rcsga9HqdZPiZHX4t2JrV3hi3GGp5hECHZNO8rs80hDf6J6jOqGd
J0bMWtG5ii1XqdLX83XiuYt/9t4SaKxw94g32j62dL26h7tpQs/ORnpDNV/w3kwp
5htjX4GLzEVlvAhbA2NoQC7uiHuPt1LbmpgDBFRNef3MX6m+h0M1bnOFCQMPYcJx
1VPn5Nut60yJ3sUNQ1nu//ORTP/3dEkJDSxLW7oaf/LWnnNuK7ovdXIP7f7JcLsS
1OiQFImwOXeGuTKDNlGpc+oU8BQet7cNlQ6skukGUfE07aoiX7LGH0rfbQsOJwaB
X/KzVprOafb9JfR7Zp2XORNIpHbttm0xQ43wLF/NGrYIHT7Q8ep03RP1FJKre/4/
HwcN6tbroSmWyqB6Ig8B1+dZ6kD0k48CCsbIBkOMnn28Zac3CeSk+v93uD/3XIl+
A+RmnSKFRa4ssJHilCptYawDkWIaWnrjhG8IoEWTWllczSecDuBA8lI75ElfRMBR
K0nrfJxFnI3lbD60yPbfG+XAyDwCsQG65k8mrMCgKWxz8GYAcw2emlpVhJiKWh/u
/Haj3aL/syjyco01qvo586dxcP/OsMcQ+awOLwDee4cEbxiOKYIG+8sQqklHFLLG
3ydNA3AsdmfkjKigS+rIYAzQOlLMxyQwMoxibB+Wd7XL2OTgCPRnmz/TD+kbqirK
CqZAsgZDnm4r3GVbK9tllgZvP1V59sLtVW8P1BB91mmiavhblFZ+NlTEQcp2U9iY
T7KBg8ExaAWGm2tDDJknJR4BvdXLlQqs/rfP1veqkrfdAGLWoEqNVPAqs5Zx1GLC
xuy6mgG56VuUbQqOt4ndrAWdHZkg3CiImhkNkgUdwjwI2h77vxuQvoieKW73WqP4
7L5mJavwuokc/Ej/s3A8MKAdUWgL3Y+W+2rTc6K+E+EnSJVpKw/uXO/uEhoMBwRO
GMERXUumxw7XGaSWg3K5SLH7Zdl1a/wvl+V3WiTQ4Qyi08W+KVjG1eqhgHCyZygl
3bMUuLfMuE7/9gCdlwysKbpai43iuoRm+R7pGgk3XEzTIpNDySWmN2IZQizfCiyI
bF5k4CZaxatXsNQ/oQU+hehVyOYhYkQrlVITk7LtchZqZ4kjbXm6L6uWiXZwetSE
h2x1/01Kju3ua4TKuUli0gD05kDVdcU3TFjnTqT+MsDJ9awDKH3W2CoKHPEAM0L7
2z+dPKeekihRVNkrQzr2IZQd51s5rHaMFsVEq/lYXwV8T47Q6R6oRiENjd748p3t
1GRmmvXqqj1Aa2MR9gT3buKbz12rwqdHMceDyvrH0fV5OLZRpuogcRllBJarAtCi
b9dJ7th/DvSqNjIMFt09HRDLX5rbK0DP+v4w8zSRypHqfvem+yG/U6QSL2jGeM4b
uraZYuXNr3E4jUKm4V8g4T9p2CNQXElwYq8Q7VMeaKtcEr95sx5+K0pdam4HzTTw
kS4/Nmf0GuCrO+qYoXwe0hE1j9bL66IDSz+mZMJ+h3MsBEbADwDdl/Chkdt5wzKw
Q+rtQyWkt9vTr0Mn2pFk96XJ5vmD0pLRVXOGCNmd/Lm4XBkWy0cXMusj04+Kt5TU
ehjTpblx8vdDx+SzgVk2pTus4srqsdU4FMnl8NgS8ArfYIK7ftzW0VhnSkuyasQz
hs6AX7fFfBpKocp9bOEgDl3LU4DOiUb0Ev7+ikrzEXpY5L8ZIuIW7n+xsfdT4gkp
LG6PupcCxs2e136i7WUjufzx7kGku6f0/VY57bm5qtJUjrXV1QdA0UKG3bmzBerX
g5ExGOyM4DYsYut9VrLbEUmKZgVSA4Odw8GdlPPz6mND+dsD9IzvRXTNktHcPGAT
PJxY0WiqmCsCZxREnZ3HI/R0Ku4Mzt4nddYCteFFqcxNV2tUVLpMlUq23Skh6k0V
6ECfXnX6KOHmii8BsFNkQMURoFyxoLnVnGsk5oVnX0SFkV6Zm3N4UV4dtTHASIYQ
HLajxPN8SKZBMSA2jVj79wuK2PbXi1x7yw1RXzPlLCmiJzdfq+I1GjO7nzZNljVf
+/w5l7VgiO/CpaOdYYzLG+RrX+sOPVGnsWvWs2sDxcp2GizE7ObKYX7ucA1ycPuZ
NYvEWqLMO2UqiTcIk09P9Tqoa94SmyiZ/jbUSFZGgQp44Od9HG3gP7JIqvqdUePp
nxFGd5wKJLTcuM7hgA/9X5BfshwgT++zk2idbBHsN7LuRkqHkJro7sLHy0FA5986
zRq5qnbXNV96TKrrIIm2scagsctFCw7rVpcZir95oJIQ3akRDC4P/XGgcaGQzFCE
TD3gJ5/UspsFACTpyE6klFGtqFGZkg8wHeTkPM98xn+DDUjmO6s1AvAkVBTqshgJ
iD2e0Ui/fS7UVU5uHyyRTssGGfWuwia3jRlpJkiikuShBdSpLsCpGRWlOIgQyPjd
NkCkrfVn8D5Uf7+C/i9VPIfvXT0DRMIq5Tj6qegs3ErXLOLu69HCeS+dKDca8VMH
x7z+0UFLxVdlPjF6GTi3pwVoV6zn5o7uzHgqSWU3oUYJN7xiPMH/YxsHeVxcHoba
LIavOEyoaHjquL2vbEpSA3Qxkz61s3SBhzaje4D6ZFvGio8FFNBZtyVD6VXXorsO
YHUjiJfpKaw7zBaT1OLRKU4YIkzjOUN3rIxvLY9E7SJnxiBlTokZvpPK0zER22lQ
KGl9ORbfZdFWlgrXuk3Cq1TVhj4La0pJC9sYhG6P6V3OYE/vkkG4BMprQWDQ9/t2
qDlwuC98X6K6WQ2/NnziA14hH0xW+JZJsgNJ+2x+vKwD522498WMP2bgISTl5H0z
3n1BcqN25MT+ympUPag59GGjymBIcW6gJN/PzZYSM6yXWbVNquaX1uAgRWZb5gjC
t5l0kWQoCMybBLzoxZShmuaVJlbJKNPAaVCB9EtXiMLv3kBYVKT2H+r1oNnLZX+u
Bm/a7ofsHLPx2n0b85D6R/7IgBHyaJbbF+3m9eoKX8aXUbrzgR4Tf5+uhE5IVGa5
ZBygr8xLv/GevIyTfPTk92Bd1sFlZ4r8p1NL4bR/BmM6qNU1JSdrdcSpMBOYYTYk
b+MJHb9wK5YjxGgPclZAc0oq/jEQljqSvb3sWknpneaFgt6fH4oP5q8rduaJ1Tgk
oACcbO2jb/8uZzXOty71a8NxBwBWE5APbaPE3vP5HFTsAbNUwzcZDnm3WmsDnP9X
pHatz1n1kDFg1yOlyQ901uLOhntXL3oi/560l0JJgn8AKdj+DsWZxboXs3oVp/Kx
CdnloAtYy7vVrM/rzYWXfQ9/Bqai1ugZsxNKhkbMvAxlikHLPngsTdDXJ4Rx+xw/
xTJPvW+oNtnYO3YvvNjgQD2l3aixt1EfowMXCWkUdT0UpoJUCLfjiJorxNpPS4g8
ic/jeQwT+7AIyyGQLVhRmlj06H18asYLZ0dbgdLazldKF5+/EmpPzjS0sXgdBwD/
3Vs3N+rXzZvOfEUis24shwnaY2B6jnlIV2ss2MGEBwG7Xl4KGKNsertUiNcQPg8L
bHwjXdY3qSfqZfjX3AhLMcb82y9bQkr2gn/wBbLS2JGA5Wfyf9/qOBb5TdlFQrQV
X9ZSGVwKQZ0mTXGOBAZksh3GkksglRfFx/RLrZZrLdqez54cBJyPNAZfm6pnIvon
pKUbDZ6Ol+7y/4bK4iH/7HS7WJz/bxXqLedqtslMEZ1ZzXDMxdyiX+8mfcTFo0C4
onB6Bqjsa8kloCKpDwDEKCjNf5rGByzpIWyMqlxjqHm9zjcidGvx3WTWdWgc2QM0
RdPageltpxvCHKEvw1LwIv76Sonyr8ZvLRh70cOXsjzIkmDSrQwMFqbyJFi752sG
yf0o4oeeMgKEk12dKPS+lSEfcghWTEZqpvizTDIZTAE+KLqLz0jDFDb8RIIqtptX
jUmn/Moh76VZLdftwad+NJ0dPFtGzJDfm/iFsXuWUIVT9wAnINr8xoK3ZI5EBwRt
O0HgqC+0qg14FubE8o+QTGnmhLCVq84y1DLhfXV8k2BsBD8HTCFEfhxpdKuvgKnY
w+CVnQeVnavnuFFMh6q6QdvYnSjDeDiHcifgJPCwSWWzm+Kn42Ex5pl0vhcyia19
vCrpWqsNm8/OR+sTCRV1WsbJKYW8m0D51bgOShswBavllGVCVPiVJMwpvKUmV64j
W6Yt+AvoVzOXeTWW41afFg5C9okBSRKWxSo+QwKw5HqxMWDODZDDLUfwogp0jbYd
Q+KuTZLKJXykUfL6Rp9XRgB4byx0xNjlUlkm+f4yOXQq+m45JFwMoAbvMZ3htZHC
dKXsu8MKy5I0NGz/EIa+2OB0kepxeS1WyPMvYbQ99gO072up4Iw3i9ihOMDbhx42
7tEyIvQnRZ44I4UpmDFwhkiGiP6cQp0lq9TmmFVQCGm78r1BbmaXSznMgoUphPp6
ozuoMCChxVr+SgpMNDEmV0nBk+54kUDRTuWvKBCMdjp2N8hullyRoOM2QXVTYlWi
EoXOGFQbR+XeZDdhIncf+ZmKDuHRNVRsd5c5+cxVt0RFQDvIjJmSpZoESlvN6NpL
WwDVFgQlmLFiIbU1LpLpRjt9l3rw5cpvNxYCOPRT+1mDmu/w9cP3JzCqppaVJD6x
aR6t6N1E1O8252odHybdlE+o5SjX7GjUgu7NRrrrV+zwe+seNziCnnoDPcShAGPE
H7tnj157LnuqMpv5027RMSvM5yvgPWFbnDzTq2fYkudMv5PlQLFDqAXMesR7uabx
nYyibZMZizrMJfUQPn/aY0ueM6K1iksbMcFcW0TqBXDXeCxRZ8wOjReot9Oh+z3C
vI8U9QXcm5tXghPWwL4tytian8qacmeTcg/BQN/8kgFXjRjRvDdh+k1Gk6+YNq9m
P7vr6ThH0PcE9wEMIyL8kT84qM3wrfKhmCqySKvqEIuTXoDp6rk0LzEgSyzxN8wk
BMNESKsvupRXDLtctweOdWbDFg8yoie8tXGRBJh+AQ2SAwwNcp2SujILsP+5QjxN
VHmFE2Bm31GveFTcFHh5owteGxAVHVUXYYH+rG6JxOOAvvs4SmEjkT9qUdnDe0ql
zlMB1iA8RWE9fD9ZqnRfk0Zl9K+tVdjvpA3Mm4hEGlVUWPd9aSg6eKQaHRqJ/AEn
HNubWgoyEhTiwLe8NkrS6SDaaD3+vlVaREPXg34PXYkcKW1Z2M+kR/BF5Bu8gA60
dWSATHb5Q6FzKbM5wB0KD4v1NpUidJvqY8CmpGE2YODIgea1oXKU0uELNbf4z6Ej
4efmPnRcbPKRRabtPjvKVghfBf1V4oais9tEeda9CiKxQ5d1qVDu2Jbp6zbznfiI
B/mOjdZ9N7Ulj705nvfHJBTV9KikxoBhsMmS1SZsK7g1Teh3YmhrbH9SEdg8GXHl
CK/8AHdRovMNLnGVVv41rWdP8UqP88bNyIegLofMOizj7H6cNxUidRNJzeeqURGX
8FkgOZ8/4rlahAzmmg4N4KhCIKSABsd+TeYIKktb7bNAPfrYAnc8ysjyJXV25zrW
broKbN6ltc4QKETpoAci7fVJDtCqt7irJDj/8ClB8c/V9WPrJfdokB4S85xASVRS
XvF/XJNLuObulE0u3VVGcpKFDQd46uVHPlJ6a1IVxPmvT8dnGg98nVQxF5R/zXE4
OB8Vx08he3TZV/ctfvYqxa/ogykoCki/90ujaHhMNLQ+TLNRhNVlAqBCVtxX6Eoj
5E64CqiPCga3Ny3CfKROVmM1AlfJn6k+2WVM8lqr8a6WUmVNQg2ffjgwLOMcAVq2
99I1VuXAe+2Hb1yL6Wok9sU4WbbBJDdJLjXjM5d6LI5wk/R/TH0XsxsjN0ntoqF/
a5HDdJTkWQC3Pd+Tm+KY7d+mQD3qJSG5yPsKCNIjARBKRoywvzH/sxkL47P9Ro5m
2kmdUrYKwYnYWmlEci2cKyvQuEjqy0pn2OvMUNma8+2eODNutXyUX7UvAY2mG1V8
l7lYFm/OfvuI7HooBo4blVq4RykEMn+F+qXbQKFIlKFswWycc0GgjP/Il/q5dCDY
B3fEbFgXgTH5rklurk21TqvSXxuJU352TrcEoEEruQPBD6rbLgNZu2AT/EyPyyqZ
gZjc9c+8kxqJg/ROkIOz2wC0xS0fjC/rolPuCQ06mLApaFxs83tEhzMpkh+3pWvn
+lIP8FrtQnpZCEVcsg29pOHXZoCRzUbGNIm2v8qvHS5M0ihBgiVr0rsF4hJ6Mf2X
D3wqpDyEasjbtHtkRHwpydvf6BR1FFWjzOrh+3EseBxUDRvfoFMbnqIEJihDoOdN
M1VLvPf58MHyvdRYBonurFWpqjsgEp/Pm3BUxCWRVfOIKhP8ANdgwC3S88nweEm4
ejA6aj0N3iZEehoflSeIP4mPs5BXqBQG7/W16kLGl3JCbq5GP0pVOjxrGLgITihd
gknIFYSRq5Q0SGw/soxdaatnS4aES2ogNHPhIxC8WVY/lXA+Wbfx1pii+AyeQ93g
dm1lxno4I6AVdc1Ti43ZqmF1Ih48RKIaiuBsWy+twOwXD9/T1nGXkalCvNaQP44r
8yuJdmpq8nCaCiO/afXYAhiIRJJQOcN1Mt9jq9lvF7CKCGbSx5+dAYcWcz1hvsXo
6CqbjBQyP/D6b9XX/iYrUHv00wdRJxOZf2KxvrZtGpzDeYZ46uUKZpZru4PdlMS2
/77QZ7yLSumeBaY6sN5dI0+kysX4g92YEwGDWsmgoJCR/ESHA7UE3eomRhm0CrIC
/AViwkSXjtu/iyqp0UK49/My97eW2Op9uj/Huah0q4dYHr5J6uUwOT1bAGGuSvpu
Vckx1qP+8pwtHO0fesGFU/JVhb8b5j8Ht4pt26SDbvyMMhYJZtxdRtOnjJ7T91rU
8/l0seeCV1NYoSEub8CMGPV1GImIZPJFdO9OwctYR2QfMx4MAExRnOkWaRJvV0km
Q3xCIAXk8E4Z80bK/52b3uh2mer2hgXboVeMrarNVmFGbgimvmpuhNtWdYEQvL3T
h0+6yP92We+K5SzCf2h4tNEBRn03UhqXoHV0huVAj/k=
`protect END_PROTECTED
