`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
crGX2IPlThFNpDYXX0Fqje9VA70QXAslduZoicXD2aAYB7Z5XDBBnDCI01jJYZMg
FKlXVUDIlftM7m8xxLlPWHjy8T8yQJKSXcYOaojpj45ihX3m41SrA+bQdjXUEO81
1/6AiU5DSDwYuGgWT/gRGkGnV58vLCEEm4efdJUFNl7GZD9OXAH1IyqaYVF96Pyc
3mg/wQ6PNiuZW5J41Y3sYtkbbQHDy+6F7G+/CbupspSYdCjrb5wEMxLo5vBikB9M
Ar/Pi/R5LGaiZwMtB2PbrXZd7itdnPTvHlkqHPfW6BYMTubN3yXOeJ5EE0qyZIs7
zRL/3V0dyoK2GDbNg9gWbT7D4wcwFHCgl9u8uT1BDMJan4KuWfGelumAqt4aFdCn
/vE/lEdcxkXoRDVXZFxVZAFZIrGP9fBhIcd8tOToQFAKtz9yO/DgJbmuLfc+hJsD
MbMgYXsPTU06pGLFOLPgEydz3uo9M3LLnPeW7d0YQ5PuVJBSHWEYHrDVGNxQvUFV
PSZvKj6mxgvZaYiaarB7JGmyBbQpMZil2rttDWFL0s797q7KmvL7YMpfdGU230rh
WH7+nD7VOKFKCF0Ys8mGdx4mfRdjgwSrZExinqMLJs9E59FoHO0OwE+rwgywwdoi
EX6hTKj0z9lMi5eBT9twScus8migOHe0cMF3qA5E7Sxk4dl9lPTMPc09RScOWVsY
B/xx6okEtyFnD+KmhyZtJNUKI+T4FuJMT5r2UtW+Fk4+5oWeOM8ob2cOet9ZmxR7
KuPH2Cj2lJgSTy54FHu4Jbs3BKpDcf2AFffdjWNElqx/erXMJsdlggDYhbtpny4V
TU2AfBw8u4ZCelg8DCGwmNZL15HY3Z52Xfg0VJ6BSCRGe8e5d8oS8VKcXP0feLbI
s/gIVhm/k6WZWpSxEyOvsfYx/Bx77z3ZhO4o1CvTfyxtRenIAUX7lWHFEpnEh0lB
Sr2HBvcIqAdrPdy8zXX03Gaj58odFVPIhIr9eF2gm36DT3bdo8r4TUe0vNkswzIG
uWlg7p3FTqF1MOhceOZJm8uy4qv/74ZEdOxP1XWdb0RaXbj8HQ8Y7TZ08swxi3uo
jYGiCFt5Y1nj8cGzHJ1wRvyvBsLSPD2cvBT4kWWIa0xgcnv4nSHD5L7BHHDKDQBW
GyQKa6KcO6vwhTaak1dYS1E0rDh+DrnfVWtuE+zuzFpjWnOPaBvRBo6MlsxFbxop
ij7VLiwX0zJ5b0Re1trHXRKSHb9s4LKlXdkQXUFDjYzPe4TKWdNrz8B9ocS9cOO/
aINdY5S1ShIuiU2Ad7P7Fpy6IE1HQm0iAeOnNdrctrrPkJJruU2dRk8+rUCUwbmT
3ZH6NBV/tVwYXaCAkKfSYNd900/RMlcDClZendT42yfhMTEWUtIXk1qjRs0iywCY
KVH/pxiskftoCSIscMg+Cps5cW/3XfW6I0pMSW0X5DHzoh0xt4ZIBsceWLrkhdek
tT4cxzIioDiWYKcCcgqerIcWEuOmrdXXVepO2CKbUxjsFYlxZb/Z3DAj9C24LK3D
b0BNTGKOdhx61Bpby+R3Z7fnnD8mm3OejsTkE6h3UzObIeBmuBwWOYdJqHX+BIC+
wTf9N4f2qAg1KnWhQPgBT4uPGmPClI/afwBkocQKu0zG8QJWbQiSVvTG1WEqZIRR
nAlYiiYjU28cTWIhQjfLd6k5YKFru6ABfWsT1fwz5yqG1Mi3yfg5ERVWHY9QOnd4
i3Iknsf8JWIP4ioQIEZzyluJzcdpGgCbn+5Ml6VzhVCkmsq9CstW385Tf4QO7PYA
tlcMzv+M0ZjMr8FeXbtav6ESF7DNYB7QwBc5I7ZaQk8lIHElBgmkuCtdW84/J8CK
R0V6RkrNQMKvIbwbejVZ2PZPxEGyNbquNO5m2KsfwC6RA2LjZSyk5YcHiHg5EKcY
ur3ezEsbyHVXCPyZxJV6D43gb/DHeZAnKaNCOPjpKcG347w4rjmqPyKsuTpCTea0
4QBtC9RXmIGWmsmetfWPBm8ch03cYatdXJoV5XCy3/3+U4cd9nsmjcnU2sCfcJLF
TpaTSBBmDCbOG59j914YY4PO/iQHQWNMu3w8TQnJJjx7wRnWvczJKUKFrlXVyl9E
KB2J3AYfh9IT1mffFUO+ucAxjy6KHC7KQ+6AQadxQSh94eon9+Q3zEV/8S3ARVXF
LsxpkTeor8nA9HBjm52WdCUrIR6GPaeKek3PGzXzL/gnf7Ws6sYzuMzUn8whwdUI
2mbqGnoDR3yEJOPxvPliesD3i+VcP3kA/XXoqwPg6xFI+12jO+a8JE8q15EcUeNM
MHKwj1mrNHoJnpsfrFdNHIbj1+DqgiSymjpC7RRqHLvNM4jR4f/ZpnxUWN3uU2d6
V7SBrUjbvaIFPZVoetrSPsuzmeAJWYdBwQ5tOKqNsHLYuUOB1GeqaPf/+qn2eT3z
WObYJxLLZDN+Qgvw26afHRgZ8fDfMSMrGvJkYiPfItShQ2CDDNKOpqPq0ovs2+ZC
I8omcV6fz/aJXtPJ7qGjckCxkFh8/SSDb8PFD/g8kioZZj5VYB4pkPQW1uiPlZGO
Cbb9mPpGc1Mn8kniJGP6i0xsQiEvI+05abQ5WQrh0VwOob1uAYjgsdFY4LGdwX2H
rPfDZHA+yVvTTYiSVpstu2ZukaWOyW0XVaBBGnC96z6pRigU6d0KVq+S3URLdaSq
tlMPlRVWTqRcxZ3Kf8XoouYvF5O5FHmnONcZa2f5Xo1G535kzEh/6sFrjbcFAuKH
vi/axfeyNWXmdGbfE5iijpbOkRCvUMdBvt1a0J/LPB3zzXDxO9v/JJS4ZFxL0+CG
F7ef87LDM/18pj1fvdK/xfpYRmoD+YNeaHUefYxtruZrsoDubk9Vw0Wk+Hp0LpHN
Br5GwkJSURSH1c/aKlUxYcnyF/XJLbfw/G13bsJSF3AIIh6lPd+uvFTYdQZ3ik4Q
SbGUm3+kVnFn1Uhnb6Jm3JewFHO79TiRtOlHj9AyaLvlTB7SQuQ0/THKQAw2BRgE
dw+6ZN0ZkQ0DDgN1zmfRxZeCFDit1vz6rW0mpN/Hx2zqaIbu7j2bfADaMuBfx6m9
qayBUoUwgUpY7VgYW778xHHllCh7jE++QGzXhEgxAj/Cdp1v40CzOf4UqPhfv3OF
xZk6dA8HWuCD2IVpTbywjB6LPPyYy3ImepWbQBC5hJjWqlvnO01lpbVCQgJBgT2a
VPN54oQrCFif4XESB3bq+r0kDxP2WvzbLgGTnq5aFgF86ZezDOTb/NItJAvwDj17
FE1kIxmY9ZR3uIuSB0sFicIgvjxU86DCWym2rvJIGyQQOdfISjVHKj4SjHz1KFet
aya70eNfXjGen7KpEDihT2n1JK8SNTq9pqV54tfp3Ac8waGwF/3nBWW5abMYLN3x
3ERTqkC3koao7MJcbXdJVxDPO/zHecM9zOVgdvp5OFWii56VgdMeMssst3gsSyzw
8XdMfE0Nq1IhPyMr2pjrL7UHZsdAB1+euxjd4EBWRf6LNUz7xL7+6Sjx5sbdoPMR
Tq23ZCKxtE96J0Xw8Qll2gz2/k5rkK/+0jAzsoIni4mUWfdpD7gpf8OSvqTO21Bh
aIzPb6jdY4aB82MeqjqKVqIQy4EvvBJVP5uny10/I9BgTH1KZxbVFqJX3tNwIO+L
Tq3Cc1XXsl5+dnnwLLzNF0e9QXRc1SnMTkJbNK/xQfetLtwK1BAcwoEBmNe9mXdP
LbTPAz3lgsPS/PvTeXwBAtgQKtFrd8q+p6LUxL4bqVrw5RtunRtBh3dsw2wIO/X4
1gaFOJ60m2jMq1ORMM4Xl5RZfEih8o1CtFnYjWs/OZeKq8NReINOQrOCRlCcnF/k
K1xlD7BP/wKoVrMKO2DRw3cQPnVoGmec95Yv4wDNDWrR0fXwe0Psaq0/7CVVUSG4
kbOCmihDpBS9RjCqXMf2dSsozhhHLdgsEkcycHtUYcIlAYuHV90mp5y18IrGP/If
skzYMA+PqiOPShl11smOWGIXRxsZW7urj66V8rvDrRZH3FIVnM2yVv08cONCiqm6
Cxj0OW9wzPYYtQEesTqc/UuuGxaFLtMTmvzGbaByj8+NkEZjbgBUi0e4P5SEvSq7
Hm3YTByiSlkpBMW/PMUeO001ginjbl4lvATG2xKiLrXLD+dbCNDo69k1j2rsQ0xL
IKUkz2rrpieFFSmSsD/iySEUlibpmWuVa99UcUswTfip/HB2GkkCN7ktpQQEZ1VR
OHRGFScRlZ4yEJR3983N/llpWeeS/IofaiK69lphHkIB3QkNK9/drsWwM4d37hpK
34OsrCFZYZ8suNK5J8iaqvcXuXlk4L/MSwtz2qcugUqbzInOtjVfPmcbvmJgcLlV
WyJysA5LkFiT7XCpBxJCKEmhCZIyPnUCCK6pTIrC3Gj3G4C6vuuL0/kYciYtZ+pc
BODTP39wAh3xXhf0aJ7p0Y/VZSUwJXZ1vrCHsXn3nicU10JWqfHIToTkVdb7X2Ub
59Mrp+AgF77A8XRJ9ODPE2QaskPmCS5FPwjbk0jtriSACo5BaTlnSo5jtnqP9C2J
N3p+BV30aqjghJHXrJUYqA==
`protect END_PROTECTED
