`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N0Ux7k8O5Z5RnJUMnSxTC9vBbJAajyyMqPU+weB0giBQmadIIZZZVTBzu2TgaSBD
6TYfRawzjtqMVOOZrznKqXvuQ7jKmo6NK1N6OtrFpX4Vstc7OqRk7CC+dcP7udge
gxzN5wU14stxLwjinvQuAIZd2JDXZj/wVWT8Du1chSl++sKnfGiMUFFOOBy7Ribk
DwUID+kPPwLw8GvJIOIRdgn9IqveGMUD6FM6n7bF1L950SRoLrWZk9JNbKO1UT3F
S1IakIvCPxnTu5NDvSHgnRCR2LEOBh0WtWytx6WJ7mbv2BlRgiNNCs3vimeX+jx7
umaXPYdcvYwJfKGIEtD185Dq5NAk3DuuPie8jxjCxi0Cx8BUNT6x5LRSNrJ2qwh0
44QGudPOX0qOQoJjmdTUQCb1X+rqXaet02ImKysmUZHmkljgpOjxIqlN3qpp+eVR
5053Xxkfj0joNHmC68smMj+/arfUmVNm6Np2tQirb11fJe2FRk/OrMrkN4oeI32v
TlPdP7QWurKjJtMt2bTPnIxO2ZzNVXTIYRj4LIrl/fWbDdqsP+haJYBvP+5GsoHQ
gAtLgIPzg9x6cC3zapq1Rl83v3nMIkop/jKG2ha1QMQZdX2iqYftNrs+Btfw2F+J
rFTO9myBtYPJkOJW0lekDvw1Sm05AR3WDCNO1Y1STNJkK5/RqWiDmZbrTlPRIqO3
Nsr6Nwc68+WQXJy4ZhAavYMc5aLVlH1TVak53/LMCkajBe90gXVLi5GAkCQdNDBe
PWy8ByNO/dHxeDozKodEjkXui0xThSKNI2vIFEEy5VWHr+Mqo/0ulMAUNklxUqcm
j741fHJMQZMjkQqf1/YuptVwvDxkJZLFGbEMNUX1vs4DJEHxredP2P9tkiWAvXFh
vf6XCZoRN/fZdXseRFMBe32TwZPLlbajm3WsLQxpwjejkNSgVaowwfvlfPeTi9/V
X22Pvlda1/rKhLeWHXFuk4L/3wL25DtNbGofGwz38KdDySpzqBtFFKmA3YW3wpsa
QrZIV2g4DqHsBBoV1WDkjQ==
`protect END_PROTECTED
