`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SZ9DumsFfyl35h2SIzRIHiQBj1KFHRG740GJfDvSEdiHDVdLHD3tptRxqk8UDzz4
qABlVJv1gFuHQ5Czv7qtakG74tBdsfsLb2eUrcwaG4H6FsYu5+bm917cWn7hnGcq
fhcyrwjw3K2xxBHHUGVKE9QQgLq53J1/LK0w1NkOhYLM0RfY2b5jIur4f7oHmPFc
rLAW5Ik0drM0R9/9u7b/WSxInChPY8Eod/Hx3KRj/W9C7PU0n6eUoEOP5NErX1dC
XRBJbi4ndAJhHv25FgRonLq/hD/2GRVjyQILMF/s8ooNONDmJgWiKmStAb+55Lb2
LAz9uLhdRtqPUJTocIxRawgcrhr6v5jNSIWXbE/n2/QziAIDyJv8GL5N8iYHUd8v
M45dl/RJY+ueoSCa1bHGnNg/X8DhSYCTLGgimLgzSwBnhOH0x9HvEsicG7+7D21s
zvasUghj319nGLBfqTyPXWD/tmlWhLvIWS7g9PCAP8bFWATob4daP1/4yMpSAc7j
7Rc0bTRHLGPj4L7+ZZ23IpSJEUTamsOfHwvC4aZVSjsepeg5eYhyizbe5h2TjZmh
a64XLfMjezx5KpkgbHYEsJBhjdhmMj/5cEch/pdQv88ak0LNBuM5LXQIk76pZatm
`protect END_PROTECTED
