`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
86h7uRqIR6QohimsUfgCoVj7ZU25Hh77wj3AfDkdBujSMlmJRGsiiQjOTw1gtTzK
SFg27dqsKqtW9Mk4IElJqjjvsNTOr4jbdCkibZSdS39mKa6ULO8rGHR3QC2/ggwG
I7yzJXXnX2aVwmbUfMQafkWaeFtrnGu405JdbyCirisasiki3ZknaCCyCdOWbsTL
JjaMiTkc66Gsc16MJNZ33bBxJ2ejjAc9RA4m562WPX3xEEQf3MI4tjGYI/xXpuQ2
U3VHloZBBFXJ/r2OOQemL9ZD90TSrsPAWjhp74iOwRljMcMLl1r4+W61ToXVGTmx
AozNfDRLSmj5drIjg1BnWsdN/tlcVy0Rnx7Ys9DfkwU=
`protect END_PROTECTED
