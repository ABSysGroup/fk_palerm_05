`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m3eMBCK9HvahFXJEBwBXvdYm3kD242Jj1+KTWYUT/YDxLuMpedjTAoARtGBSuLNk
PYJQPOrCOh9PyH18hgZcFnSR/X1j+pcePfpOxmegjioR7Fg26AZ1B08/bk6QpGCt
QplU6Dc2zAwpdIHmLWxrjviTOcpBijN9wvGZZXnH64W7ZLKwWw+cEyemTuQMQ6V2
qQKw3ChRsqtAXkrUA/2ohqENTZPEyiUZ8+oLE3UWvT4aUs8chW0HvNrFIdSWxgK/
lAuWhgVRZFmJRHTOtVgomKcftCO+UlXV5aBDhCo3PQMlXJo0p84Q0VYZ2JtDvPWc
`protect END_PROTECTED
