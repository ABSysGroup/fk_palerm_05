`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tll9Tyg4nP3WSyzzFVfcI0mxbEdibLA7N3+14BfkE8eGzurGiHjbWtym4GsCdxzO
r5csEITZWRLBgjYYx5szcSLEDR34BTxrJWYOan91Q8LYP9jfTZdenVMUNWVHh55G
etfGarvKDBBvoDh5FeuvfxEdIugnLEIGkoADbjTeRK7In4ACu+7/3lVYjeEs9wmf
q9Cquo1LvLthwO0OmkFMlWAv+xSMNaudU8M4nwXopthqLR7RfkjhNom8+zwIDITa
Ix6CcIVRx492gFbh6w9G3DdjxqWJ/frO2c7iUWd2vBkunL5HYHN6JShaEKScdFQg
d2HgSmf3U/KHgZRqYV4wpQI8TPoeJ6QGC9nVFKGVqnoaZeDCZ2VeO1r2fYiCypLd
oyzvv19zHWfNHUy4D9ECCy8KB0+odk9y4yDkIQlzmP+3l5j4lChOsyqPq/gjDT+7
lrTXCxFUxT9Hlfc8jvB0lMRSmiggG8MqYiCnw3RYd84A0z46asnSpSbU48z6Zry1
eA55DfW64FqftybN2+YcBIHpS3ltovmZqI9mVKTbGuzpZ4xsVY6eDv7QuCOjvaSU
JNPUQ0GoPrndd6u8GJmEInWNVIF95zGjTMN9MG9Izs5bN6mqSbjck2Zpb5nyriUe
tR8LaInLRbTsDn78i4+xHiMVJUaldZ6uxUYq5dvgzm7KVBBK0E6kcr3VS/BKqyDN
xyeMp9Q5aoUULPx/KbgxN+gERdrABaBJtrb4jfvoj5DuA8YDnpX5qyvg7XDAlYOa
RU57UiOIAKv1gess4bLu0aunLe7PvJcYyJWCYOTXTdrcMCXP7OLrQ0zKuhOBqI1Z
worocjxXCdjbuXf717cBljZmsNPwaWThVMzekxoVRToqVeu1+ga6ffRt3ddfrvlI
ZhcagfP+hO6Kq6+oQwRLuabuEvF9bDmmIZlQI20Fcj+5OHPZ/HGZ8cEbfxaD18mo
T7iixZ8dr/6JJU4tubZxUFTGhokOmaJ0dMQExt/ZfqalidfG2REy4vpes9R4mwt9
8tM/61qiGjE9omkl50PaqTxN7sDXsn6h1dby5T2mKXMyHbTY9gCcwiAGbKxRKlEd
P1mkmAw/V8HazwP+lz3Qm5nmdRHTRSD0LWrDxvliuw+lIWug+5hq7frpsf+iBpSu
Z4WAYuc3h//0mH7NuPbgt8dne5/YvCsZImIeolbBHgih7+cs7k8vseamIRPBfpNe
STY3xxMU621SKnJEOwLyzkkoDlxd2KCKaGLf+sxkx+9dJEws3+GbKcYv77Phxelo
110RfEZIOtyAojRvegGlnogHYg5ezVQCQliDTasy6jiDdp6SEufMtolX6O10N5u5
7s1Jxl6dwwspdN9UrcGO/a08dq1BOqDSJzBhu/FY/IZtRB1jdaHE6H3t6EjZBvfw
ntCJMkSQ3Q4nvG7zDkwkjRfXGu3mPlfY9Fk/WMtSbq2NeXuUtZUBGVZilEeGuyDW
qxKrHFWim4doHKzkgis01pJrivtYpf0UnU+zH5g03bYRxkv0+ttGK70yvxhA84MS
juthA7M/6hJ3ZnuPFedgC5ucgpiWEU2fIfMg5qYaadXfaf5Ote+1Xj0fZXZO9Vml
yL574otPKB0P+nUFavEwHa/LieniLmhRb1cqo0STIdteXwnmbRCMFNHxj8SHh9AR
zkBba0uUmL62/ig5F8XBf/DBD8DaZuNwXyXYuy4DaMRSmW8WuhwdK1so4VHJIMbD
Ug2EL2da8FoioptZnqwYBr85rCBLpeMUty10SIlGPLzgT5+jRxLgGTVpKVXtiKUs
PWRIEIh0DYLYcwGau2XwoCV57UhymNuqhvKhwNISEfFqpncNVVpT1YDvY5tPmiJl
AFtRPeaplvXxpumgWwJm8HZSCSYG6jaWzqBP0+HrUsC8/0Tye6Kc9QDHR/JUgw9C
MnnOe37KFa7XeldVfWgGeyVvu22eEuwhnubmerS5pnKJygNjwYBldbnhw0mTj6kD
BJUiiyBZTazTXjgiHG1gtzgG6wy4glzQtp9lf8rXiZbN+sP+qKngF8RZJAtq5AFk
1eCY0dIM4xjf6QlDfV5//T5lssZjASk3P6pK3jCBShI/JxUpz94FZ8gNEhekbyTS
z+VksSoxPY1orXTHfkia3/xeio1cWk0182ks6vPqciegPUh3kwdLavCPkctJ919y
+A0KR+qpYqPDdNApig3XQkWJyIKhfMJm5AonIfAh+Iurw/PbNMmUfUQek32rYunB
NpcfpqQi7CstxFaiZR7GP+bU49QYDlSE5tMYAuICQGt6pbYcAuY6aSKz+V6eVx8I
wsRGzLHbZIAAngJGlZxg78vs9Dpv1PtK3GrWmDZh/Xn3EGJbMVToX38A+5G+j29H
KVnMgn9k/o8tj4GxcLXq9bFfOE1o8Jsm34RGB38MVl/Hp0W4cjic6tkfZpe1T+TI
6aG7TB2FGZJsi+8E6QBbLjGdqEQCLHYUBtm3fA+wcfoZEyvl1DpqB0iaICIWe6fx
HPXEbvjMQrI+enVmraiznOwTEo69jmU3HWYGZrvdveY6GawxfBQBVJw43BXjRUO8
c7NCEw+8/vxjOaa90H/WMMGV4EraNW8+LUz0Cuv9uDcqww6gi7MmUKLsoAMkT0Yq
gx+FBuOpSjJrtDN3JZLWuq4EYiTc5jYdbcZ5OfQfy1Tt3LOsQMStAAfNPx/lfW73
2WbUduM+TjqNgNKgychzImW6yEjg2N27wL+KO0mpndij6C/h//9zntm5UZ10yqXb
ofPAmFnmHI1PM7NDXUQMm0oEOrQj+yW7y9LMcdzN/Gno/eYxTxFaXIPaYn04QSBG
cjUezSYEvlS1+iRHGiKxjj5w8FYwIxHjFUHZGYedQcnaIKu1k4Nd5kuppX0NtmrM
wA5MT5+pVXEKKpuCaKiXy47Rl2+7mocZht/gviC+uotmrUmy9BSUHVdXu+SWflKk
fWYVqaQUYkK+13ff1JgEOk3+crUMAEOpE0BTboCyevrE1YX3HFa+LO9m1cScS3pi
E6KWsI+MVFJFJ7/TJBkr8uQCpDUiMNWJBcBukSW7ecUFd4YwzdHnYevPFxD7DEWK
6rJ5qWDw72V5Kpnl6CItbMldzMs0n/yWFhHVa1hcbhmtXO6Px1scXaCcgIY0DeIV
HTB/1nxadlaBaYnQq8CyhXLIomsLl0AxdKvk1xJYbrHbFt1XxVS4Am4QqojS187q
Da2jTHaJzKOGYMS0dMx5JkDHfOWbAxylUlwkp7YBursKHusYSzaue945rBbXIt1K
EBtlh5s2WTvjG2kLKPUHhiFU/PHYU/LdXi7IMBQ2GrLthqxM1rYH+RmEfwkW7X32
rsW+BWj8COguRCuoYcKMcxzyLXaQB9dh0naKfAh868e03LRJK+/0Sx687U12Ovau
4SFRgo9xSgCsHKH2hoy06Dth6peQPCYXQNDSPeTf6up2i4A9RpNbZMVotujDhcvS
V7WOqXT3lLBhB+4GOYloFJAY6iTb0OiLHVSQqTiK8/zhGFuUyafqc3z/S2kqoTPG
mpoEeN0Y8XWeI1vxOpAZa7621IEGFCNnyK0RHafJqt/WnYohiKEkXW5e2pgQCs8l
Yusk1j4N28FI2TsS4+40g89eix2rJQ5Iv6ykgZrZXEg+eci0S457KsR0BJJ0eWdN
DBOMEG2AyDSYMFYEzRb/qi4DT5uG857Ef5eUu4TbFnGvTS2rBGzU/LqbezfqloqY
gw7ZsHlXRcZm83KmMM6t5Q3gY51g0NqF845rCQnLsjVuAjRqppdc3xVIZqTMKSW+
fZM+h5gJSEDCeDDquwJy6Jo+Edj2BVKYHhSawrWjxBfv3nI5y6N58FLABinbw0Qs
HYJUEWAPCH9U9kzkTCQO76vx81nNIwlpoAKEuFRNp6sQX89HONylvRYRYMyF7+kg
gSkFQ3q9SK9vxB8EN/fhgh4QjySk/M0NRceL9ZmTONQjsiZZ5S18onZuGvO02LJ5
jLKL8eceeu87czxjXPTsBXAGDpo3T2y/LdnM6bD6oRS+OSR53eMAjDwSwbHbAllY
A3sVrtqMTHo20G36JUdz3rRTucVNggfIQQ3mtFDL1UtcZBwo4fkrDssyif5h+Pve
gZH1VfiYwUNuCtt7pzJ8RdtyeqFAXIg81ozJ87cRtocA4GpoE6Aubyushsj90Hub
etMtqSbCLklg6ziUA0lw9p2RPlJtPAzkO4xCqMyIDpwgxs7ZqbdNhyNYKDafcmwf
GdHbv9K7QA03XwVKV5OBmalrEYwl+jEOb08iJIIJSb3LgQ12D2AIQAcLgjSp/lNY
/hRmveIoVKQITFADZeqtUMrhdRV5HMcIdDAGwDCMjmsFV83HOTsT6if2X4FT8LRQ
oxZ0qxcbXxKBQefOPrWUNryhgJ39BRqpPbzygTDaOW3XYDNAmZxnqasXqMr1c2/J
eHAUVb/SEkd8u5eutwiFa8KzazOKUug8zRJ9NmLF8FFDNdCyVPQ0TeX56QI5fdzo
5vMuVVK8R/kcNlQea6BO2pdajci6/jXWKtB6hVbPXCtucS2UXZmSj+01PBjwGTkX
qLUGmOT6yBipNoIAmEGb8g==
`protect END_PROTECTED
