`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/DrccfmBRDBvbP0v4bkZmDbqswAXGa7mv78XxYPZbbmLVAxVeowbmC7YgGOj6Cgi
YhiFbaz4GskNrp0Yr/pNNyHSlgWgF3kdL9gslY5ILUnYja6aEnSinwmQfk7eigY3
cN3D+sLcBbEHsMXdqdsKsfNRQjj0D54WTNrChLPFGnAWSphF3Yjxie5p1bx+fRmj
9uxtZd6zr2a4z6L/HDzxx/l0TJF6qMpYApoOFRXSahv5Om/B8OOe+K/O26ThJGa7
Vc8BRFk7/z7XfV4N4y16Pk31IYeoNtP5SP5MXgCCla1i1ocnmS4yBpuxOZHErgMM
yoWUwPebBELvSXDFIfIbODEQOxtC/KllAzML4MTCQ12s1GC5g9G02dtfF1zH6l8H
J2lmQ6JX9k67+z+AAwrMdJ9mJyDfVQ/ovnIG0s18GKQBUZXykE6Kn4ilrErIYlwc
6p1pSVyS4yby2TNaXA+iZObGe1R49K5a6HqhBuCHgNT2i+e1WDc5Epe1RljQEHRy
jhFXbKZFfMxQZW/5xqP7v+K4Jn5OksDaQvIMc0rsjOITQHhiBsfRbDr6vFSW1wn+
KiHzQbNsYBHwS/hQPWccIw6O+tU+/U8frSAg3Hx/cZoCtWR2Gvm3iUEzvf/+KZtY
OI+FgbPvk6YKYdbVIpjhsICpsC0byGNe+OaJBFur+JUeZEV6PrL1nJc2zCVc0wbe
VEfugXjNgWGPCfnpnhcAzQ==
`protect END_PROTECTED
