`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rk8y5xN8DGM8nl1HngxU+v3+wmdenK8eTEaQwiSqPg/+j23FtR4ORhlXdoNXnc5C
u7LNTqtDl/PkCq+bL0wLQqAXovivAVyzQ6nOIhxO5VNs8CPeIs+/T08GBrh17X9X
+d6LAHvh7/A6cXtGOepZsXXzqF6I6ms3cGtKGgiLbvGhyaN/i2aERL4kEn64R9FJ
O3rWiMJiTI+BsX/2hEs3f1gdAGfKHz2xqmyjx6HV+0eux5LsODvnajl/+xs3p/S2
ltJ8vc3WSs/7qZLtoZJV0MF5zrL0/TRZVK1EMIQPxdr7wLTVtqx+O/djtxzRwY66
3CA23FIkt7TlaCPUSIPSx6MElVGRxSYQTpar0CXqH5q92/BhB285mjIf9d27ReCa
uegUhG7RWvzx5lyT1WsrdMcSYNO35ljG8SyKShFd04RDM5Gcj1a7cok5YawxPS9S
D8XbpUIZRK5p3yRb2Olx1/ui9yKtElQKVCUIa5CIfZVyaGj5xbu+1KrTz1zzUKsL
Q5vKmV2y7DaYKNrGuUoxM9rrltXI7/lRMH3bydSp8BZVAXeeSyK0VZs4iWYN1mlF
u1Y72GVohqyxHsuXxtUOlX/Pdyo7bzxN9IJBAqNsLKWUA1M4knn8a/iaO0JIzJPW
nLErRte9NMSxvtJ5vDZBiRPxIHD8rOPtb4oPns1GARua/Dyg128MmEhJZsvujklZ
TJzYmVXzcGYPjzoWuAtd9ZIFLef3PeUiD8lTRKcEdNc4PT4IB662QYSvFB7Hc9IQ
I1z71mBPw6e6TmmcG0O1IkrD8KiJrgvs5m8y4CpcDv9BKRceOtN4ueNBGacPtazl
zawMVJpRjrvWTxyqTAGrUAeuGxVZjWlxlYb+lL/5Kh9M1V/JFCT7nrM/O2iQBhcx
MonSbTbpuWhdn8tWW7kI1NooDsLkC80UUhT0Ksbd1dNFU3y+EhIojtD9OJrNtQqf
h12RnmJXjomIXGWMixtcrOjBIgbdtJzlwCMvtg5qxty7Kvk1morXONxSCKmOmTak
lmdYKZrmHnw4/vcUnE7dx2oteWVlt90hRWi92hAQ0nCEH9XsJNTg556f28ZSR6Pi
AGbJ8IYxSCLlbxe20mWcmIqQ+V/xbwJVZvxJshAvIW78UOqEp4vgy38n+nTk/aVa
w69+P7SMOVIPv3gOT+DMWrjfsanPuGy1GAlSO/zqkeiopK1cUQPUlBIIBos32q7g
xDS7EWw6bCPZKVaA0Ibrwgx7MLWs55bPJgjyqKPF4SEbEApIm1Npcy1vqx1pv9NP
Yyl7oDsAqmsEIj63mQXza7W+IC75dHLs4Xe652KSxTTxgdzl/dCMqP8KIeR6yCTK
s6hash5GgflGsrvSAUpxxBItxmmU5CXtQr/RGjF4elkVNl4gVzi2ZNAC7gEu8n6l
VeWILNhgrjjyHKNlITDpeEYldC4qLsBf+V276f0mzMod318MpZ95Q5/XoD70In2u
kboD0EM50SFxbnf13qy9sbMRiw7YZvebsa1A0GkWoy5XgJQV7OyAsp5hC0dmi8fV
FCxDF4M2KQcP7OkzD3HEbVIqLD9LMl2a2S6Bz0MLHGWYKvyOvc+rgUZ3XCCd1aXA
rd9XEDiKczdLD+HdZEG+EkD3I/c2Eut15lh8bSc6jhWwRvSy4dmt3dJFyzS5LZ15
dV/Vsk8xoLjpkOqnAkvih9A1PT1Pi0REK+u5FEBZA/TqzBrQ3ZiBJwqx8FCdaiou
aIW1tM9ukvOYPHDcjUBg23SKLqrp23Ig/83xS2EmnKswSbgOAazj1Q9JNheJqutB
E6rZ2pUcLJfhzbjUar78E/jd2HZzYZXkvwqOq8D+ANFzGWiquW2V08OEiI6UA/WY
4Dm8AfiCe08HVultRQ06krOhSfzzBKtnEgCqyZvQ35OIgASjNbYCi63ZKun4s2/X
uIF79IzZWuRXBAbo0WupFN/OZN/mcZcVeFKE8MFiZesw4PAwIzoj2lLmbf+qm7/Q
0DxQ8MY0qArBLKnBNy3FKl2RQm7TEW7fbn0lvEtTXbieT8Jcnc//ofjERN/oWDQq
p+4sYXdmKG6Qz3pOMM2aVnmUEbSjyHChHc5atHCUughWpKySoP96GS/2CJnZs/iS
joL122fHVaaRbfMBH0KiQoO+v8k0eoLGN5ZAWx1Z3oh85HhXq9vgcEQmOExu7Ii0
5z970nHSeWHSXk8x/oUF4N3Rh7dtBzyyJ98YNYg7xRpuSm6pue/3hH5FfUtDU7aq
wfNoFeqrDIUMO0yB0Ye3ashagFz4m2lN7wq7QsyJ/lXo6aLYdMiyBwTDs40I/cPi
GgxL/NpMycJHRJ9H3oMKMlYFdHusQ4Hiu13J83HQRyz87NlkofH2HJMWR+/p/ZqS
JiwE5n79GylcNKcFMe6fZo2YA71nZgozEkAOiZf8tJ7WajpySCdTdYJK8YWgUPek
OBrX1KqsS5WuDyTN32OoSvyLjTsFlg1Muum5VhDL9EteDoGK8Ki9oKjCZEa3zAPy
vSB4237nXFct20QCFI5TI5HfXhAMriWPAk5Akjd8BoVynKn9/IBSmKNwBlRWzdy2
0XAySxQz131SaMzg73jCL3Op4v7Q+F1nMVfeTFZZofcd+2mMLrfXkAbY1pQKPym7
mqGxqoGiJlSAVDL2RhPDnZnZCThh+NfiVYhhZAytRS79m7c2Qw9DgujKq0hDV1um
6z9TkWfa0vgizvV4linXGOyH7yIP2EPfbQ6eWoqP4CoaE/hfKPbN4YFKKe0LJd5t
IJBTqAMjGfhyEr3EeHe2TPYUwbSTlUp9OM41IcfviVDFwNT8sA1lJeRGkIb2AAeq
jTPei2BZjEMxzEB19mT733d0CeyCdyvhysgoWC7b71VE4T65bivYRS7xF5Zft84/
PTdb3z42fj2f7mO6mbPIwd6uYgOUWaxvF/wEQVAPqt/CKUBlQY8FMHVqM5eRom6d
SPuJYoUYaHAHW3Saq4jTeGVQIgeZJOy8Q99+4SYBKeVHPH6xIlOBF+jyZbnhpvt8
od508ROHS1Nl01UiuQ3NmBaRz0/x7MN3zeOZv8WzclbmSgNA6Jbe0e/JFUTSc5S1
68QkZW1tps8R5SDRxZDHGdk1xpq1BBx1d4Edc3wmx0IEFP8bEiG7+l+kXV+QDRGr
qILJTNCAz34LAEHtoGjCGnEeQAf8+9ZKg0p2Kv/NC3HG4jduik8rjWNq6hGQpllZ
NEyl4FYORtXHQP5Uyab4gUgYz5NKjEo8TdG1QtnVQbdOvlkB+x5ZEGu+pb2yRaNl
is0nJajqljHH3dHcLz7+uoZIzYFc9LFUMUjUyQnNV2AdlGcs0ddms26Pdd5p7kQf
ZzLEnPRJwAT9yOeRp+lSfYL4zdLZKlx55tao/tNbTGwGO5TBrl0CdHE6U+w1N4Qx
ZVNjiBs+UzpqNQXMJFnUj1kUzE8WYBmBO05qLMCQQeM8rtGWjZiBrAAFrBcmY6X+
AnqKCuMOc8I5GUm+jz5/jG+YvDgNsfbEzL98eAZoB/4l3IJZ1A7Zubnr/cFcg6il
2MBlIJwlPcpZsKcIUs0GN+wrmUGKHXabjxCMncAmLXKlQZ5NghoiP7ADDfHWmedu
h2DlzjejvOt6d5IQnur51AKImwfFHh5AJYQldI2NLAs7hpEhd8hJI61ZZKX6DGeY
bS4RG2QGKQSU2zKeN7/SMth/NZzYVPcNI22o1FVej3DCuKmzl6tib579VofjPKNs
qi5StoU5OCwgUY6CB6pIMSXNqAN5VicXBLj6pZOr+seVST4OuPMr84CHu9OW5xWk
P06PwqtYkHmueBUom2GgCbf6rWoM6A4iOWbAAvuU3GzTxGfAYgfzEO43VWUHJo8K
3rincrkpN5W0wl+oWyOA9e8oEkxnr44IuhidfoSR4odog/PtiU7t3D67reulz0fZ
wgkrXSork+6OfwChBS9kgkfOLOIEacdvZe1dnjYT4bhAU/yk/dm66e6P1NZKxT1V
MlqCskxRVjOV0rXyWpGqpCSSCvl1pXg73B9jkdmlxRyxKs2HrjtLAQ/P7sShbKjN
105IUhiOiYrFQrbOGRpxg5KxaxpAiMoWIfCyUBfMZtVd6466ZZLzWjhutpjD/d0A
uB/QhU6yDd2OkUaWJ1+rYzUYBttb8MUUCU4IkPGDd0oO3ozdNvmYyD1TBN0zbTsx
hiLtkICAjfKzJFSi6Bjycj6KZbWw8jYkVKY55XtQijxqHqU/iBDq2D5caiK5PC2k
Ft+bZKeNNvxiiMa0Vc3i/Fbjasl+l0QMRjIfImyRN5rizqJGtpyDPJ2sg7BW3waz
33fySwH7dG0hVzslhxBfednA8Rp/0td+H9DEpsml7PNkLbUzmPrUq0fIL1x6BYNT
o/2azdxpo+QRyaTfZo2CE0EPwAbJ3LNS2tD5W6MZ0wHnhGvwA1q/hx1BwJyrklSF
bhOxuNnSJsxa8G+fhNxCiqIs5qP7S9vUh5f8DrTGRZgNzqMQ9VzHP8fHVmD9S/2f
Vt1wDjSjwjyYSlRbIf/qNKNFayyJWw9o7l+w4qQ/B9KnKzHWa81eqOKR+B8xzWiZ
XENAofBlZKRmdnF2Vv7w4wecQ5YzZma5XXR8WkHvLnrpERtbEtkY8qD7Erlhq38k
WUqEfEL/xZtNFi9mBA5h/qQpbR0Urs/PvghaISgEQn9OHDJ2dfgv2Vl96F/X4Fvc
ZTarwcQzwvJY716qlmr+x9aws8FM4ublNWsxQJ8iTCP66Vi11r+N6+JGUhuMYI4s
C2sUbG8SMDdX1ZAntUib8lAICvahNKNf8mZvR8TVt96bKReqmCMUQnMOB6iiQQor
IiWOChWC1amCzsIlCj22Fm2UNNuuoUrYmyCH3Wz/zdkdW7qTSA6sNtL3MAcHMzL/
zpMiCAw7+zkxW+MTn4H5wdL+JSlWsdN81P0h3idfj/M3/dfdbgUt9N+GTotfqQtJ
yeXLqtytrkFIWo5/hr2qnPJ3r6q1mNCxgJPJNQQ3yuUC58c+PSRGyWbM4sz/UysI
vN1a75SCmFKgUVIC65hxxugCbjLNgowigNpEVhqk5iOIhDONRiJARylsITl2V9ys
Kn6CB2NJl64Pfn+LyBVcN8H1soHFu1qApLMV+nhoWC/GNTaDgg0+OPiezHk81nnn
G+EukU+ie1SZZ0xDJu3JG2Nij5x5UyBdlnPSizPLKp/st87g7+IwabU5WsIMhZ/T
C7gzf7R/bZhln+PA593uyTIbVjXedM69GpOxKX3RkovONa+KtBLiMkD1qy/J5M8u
lxlu0ZRnfMKlp/unk9FebQfjT5udqENhGwq8h7DOB5N+5pEJFlzrA1+QsTeAJEeP
nLETsp/B0cpk9BsZsarGj8cE0huvuIHlAqNBuZbLYD/8JA+HGxuft06dUwfWGWxc
PRsIl/IccmsyDVtJDs4uOitAbGe+JlSGlEvcUsbNF8rsOgS0w23P1cFtIPew+Htn
FQnWrjyoLjSRea/oqjBCBzaemZW43snu+RXWTb+eYOxKM4QcO48P2JV63EKAhB3j
T+pqpD8fuhP4Pi0IZhCW46Y0faH+KWPU+HSkXuZDhZOgPvjaemkNS3L2L3F5m4bk
WtXbGsv3nPDUpoQCbKKimBu+gXyBm32Cz4KZBa2ZsOQmgdKoSNhRY5uxbEhdlhmw
z7UEn6kJAbCUDp+Tj38EkPpzWbGgQNQDuq1XmvzO/nOz3IdqabO4RkGOz6NiCqSi
QKeNW7WQfp9gaSFKm+n2SjTyzxCugyx8OB7PYev5Suegzh+rgyqyNs/LoZSWUMi8
WC81RGEnMsJorr7UKpO9/cbazSNL8RCKA6ficOw5vw9O0ZSDsFUMcGeDSiy7QPBH
WkjnlmAsRlquE6zR0N8CgB+dJanSF+tnVFo7sZTBq53rM/Mi3w72ZWz3yGQmJAfl
cwJr2kaRF+g1LrL18a76J5tPDSApJPV1/QSUxoguhoy/1M9EcLfvXT3Nhoas1v9U
s21ysaCQr0Yn9QssgitjZcAewaK1vF+rSJhP9fgasQXUFiPKEqmwjVIoWXJoht89
zp7Xt76Cxlxke2DZmPVCZEbqbwhwofcbQrP1+FlmROxeKWHTmRex46wH1CfhU1xg
pp1KNn0SVbmXg113CGmvqaRa5PcUMTHpcT6lAOlFTK4gftiFPHhBMh9IwquoVpwL
KWNI5RnbtuPC/LnRDPfmGxyn2SY/VsyTzMrlgAy++h6e5gv22BOKzCpIuFoYXyv7
+6S2TjbN1zRi6D4QNmrKz/94RZJGvFHh1etbOTOu546GtOypC5RoR65mXGFExSIt
W1Hjap9ydJrs6h/DrAfQ8E9rRinw7nX5u3AYtJv1wlUAIjd/tQbVzVyjAJW1VA6N
v3gTBm0glk1+osX+8Nb1D0P4vqODMEpc3pSThxKPP0J9FudXgO7u7qVJkIkh/fqb
3QiluIyxUrWMwO0/DNpcHzVPx7IJ1C2ojqoERg99wPeDalBqEtqaEDHuVSVwMuvf
woerNGCInUgeX6Lih2rylmUJaHjxo7jQK0A2bPx1etystelQVVm0gAjbfUttOW3I
wIlZOJGZdsgpT3xDjToCrqzDkgwSZ/wAC/wXkmwbrXMB6jCHoGTjr72D0V6ZmERk
+OQixOnSlKVuSfWPJuk2B0R9zEF4349pgpEqfKLUsbKXQ0z5zWhO6ioNJE769m62
cK5eGTMgo6nig5/0txpTwk0aqDChGgXg4/0gNlGXJQ3+SqH4MJ9CzJaCzB6TzcMX
yrCNP2F1JvnpGoVo1FC+DcQWcJ7He8ecyfThasP0JaHmpdqH12Q1cLCXWhgFsfKb
chqQAsxy7i9EBQMgsgjqNk8CLRTiYb60Rr14BdWzY7eqeJARqKgEEBnlKLM/HeJe
qgM/emsf8JE2Bv5sELqcbdLNVgRxwmWcWCwYnam5D9dfvEVcA1JxB/MVAUq4rcM8
M7F8UKuMuAE/YvBNuqF8uIceFJqgwV4S3Ut/fOLXy8HksKhpDDZQC1ugupKtwL/p
7rx3elJpaFt0Iu+xx+LdbwApdyWq5i6SOq+2v1rQ1aWIliBuB6XYP9lY/VNPTO/B
PmsW/JMzDyLWIKFJCNXILU8d/+L0YsYS59fnQTY3NkeD+dwn5SUw9X/PEIwdeztK
N/z7syo9aIu/KGiRPVQ8jM/W9TjwwuhjWXid9+GnjJgZ/AIzJzwzbYbly/vpHJWd
h67AhTYOjGp9d9671o1/JqSKPLBxtclynQa7SbNpafPjTzGMXHpXdOqtSv5HiRXe
JPwUV4+mjDffGEzMYQy0awCvmucVfAS+DQpfX9LLdq3kkoOm5FMlVwAxsYe5TW5Y
ibhvOKgDWSv8fLB6oRq3CiaeMQBhYLP9p4W1XAFBEHps8Z+30t/uMvYm1NP439/u
fXcSdaoGuw/zpjdpjXix6c0hy1Jf5jiUwrmKa9Ka15c+g7PpGos/iLpTw01ZWRTw
Lv9kEH39jDwg/pfiCibCudIN6zMThJYEpJ+vxL65dOt7Ni3N2RRZapaqICurAAeq
BfTvQiy2uCC8hPIaDBkRIcaaiQOfQBp2GaYNlDTIMl08nIMsw0UvOtIFd9s09OAz
JwA7WlBrul2Nha7lTFuVRc6lLA+YY486hh83NG70GGRP0p85rJP99NjruQ4Z6Pm3
R9kbC/xz2bK3d+hJir44pzUb8ipoAHEq7dqyCHzycgVS5Bv/eJHcgw4S+xrVfA0a
s0aeJLd8uY4z4gnq2eOku59C2/P+aIbz37AT4m6+CeL4vJNIMT8/4Fz0g0sXViaO
chX/BwaLXixaQgsV8rBFgIVpliNtoZc9+2UrPxEa0vU3TCzN031L+FMkL8CLEdpJ
5mkYwTUr83eIM8yenekPQx6c64JrCvg7ZD0B/fYKAjOhQ4iq5zq9Hwi3v36PGoI1
lt86xOSZ8R6rSxFYagaRxzpFgs78n8i2mWNqlcUCTeVu//VPsA9Bee5PCXsFyUt6
W6NB8rCE5l81Ahe2pxJkVPG6hR+ByJmPj4KpkBOwn85iQNZvqwVtGbMaZh9Nz/Xo
UoiWyHj+SL5yise2fA0KNbfW/NLzacwxCJnXL2O2aZN8XB4d44ok9kz9YB/lOxC/
vmGN4OF8TQ4LBdlym0ijQwx+d1se38UZquC25242fkKmHMEeKmYLA3fFGaS1+Mzx
lIsMsGN16CYUbp/Pc5AbyhQ67OL3jz+D3R9BQLtjubOjgEKSrgnHXXUXCnBVZ4N+
9gOa2w7/k2dzGjir7Zasb7EQQ5coJTVkUamzzyeOnOVSkzQv5zZBpGTOMccQ1GAq
XTYbPGUhzqvkUEaU4Vl7i6KQNtphHfVWMLf6VbO3kV1u6owimdVC0kahvcclL8Pe
/+3P6dHDMYQBxqlx6JtPqmzgtD3W9+a5Wm2ZVlvIXsP1zwmRW0zPVtL+EruGQSCl
3eqf6EqxFrjsZfCfYofJ01jbp7IjivwkY894UDgbP3ax3zTYDE/m+xkH0CwBky+h
0z5MsapJ0G1TJjONqbPGcBCh63kt4wh6ee7WsPrxC6h0WzzUb4yw/TqPgCGEC+vk
KGGLA/srhXjYq+WsItP+ImYY1+Sb4nw0M0DuTUi1YAGpL2T3VMKmsRL/Rt053kfw
8X7rurArmHhI29fJ0QvbWhm5wZtzEJVtu7NGdt1VdBTZKznZ/Y6A8PlRn3fvRI2k
q+/WWoJAW2zGzNp9hXPYw06b+bRr9leGFz4p5kKVFVB4vz765y00C4ZMZedAPfOm
Mw6vZWm7sAYKhdx30zjsQ+coEmt/p48LnPJKCPi/ARzftwLMayE58gB2L2MHA7dW
yfRBXgSiZrZZlnnIew52crJM203UNzUxlH74oyYONVqvidir4cZwFiLDolnVSGKL
/eThVjEHq5GIBhVb2kHOGyLFGBlbtxkLhiXTUI4+dB6VeMzHN/xkp+W7O0vVpi9Q
VmsPJ+9ppX5c7hB2dxqjlKPSEs+yT2aVLE3fe9knvCeeWNW9L0HMJSvM7BjCofZW
nOXUB5ivwE6xYIZvyExfg/i8LI/fci0LiCwr0IhhGzYJFKni2W/GdUeBu4JwGDv3
tK3XoIyAh8AJbtrua22NnQBxaDVCWkCtgguUu3TI9lvHdlfYLmMCPH4/VHNJ8vqM
6a25+b5v/LC8Y04XUf0WY+14OllxfkxiLE+hKwiBe4UY5wmUuXvmWABtDfzV6z+R
BPTI7px3LiT+vWUsFcsRiqEaAnmLSsh1iNz/lAuFNrSsxSSm9IL9Fn+OGhTqwbG/
dWYTwPLofofuWGFntMGW57H1PUcm1hIZlhRyXaE9cewBl/2vbi578P52PeEggJpi
UMPV0umcaFfAEmkKdVu2bkY0qFYTpEmM1MIlRPnBVnERIp4UbKsB81HKIE/oPXvT
5voxim7X6bRj+c9lBaTw0APau6qSqo4nZFChbI/YWoTPPkwmi+dAVWMcm3MdV04S
VuFwI6tY2ecbwJQiWpjWMUMYVR5YyQ1ZWfV9c6W+2xUaeOMqTY/MzaKVjteXFX8/
Dy8JGf8YdPE4YSGGNzfYSkubNJfiGCXQtNl+s1jIiz8uMfM+eFRyiaxtYKodMvFP
CxPwOQcmN9hsvX/0Mrm/zo8ObCSYnA5x4VV7qVqz9Lts3u76Z4VkopH3U3RENfFV
TxyTiNUypW2gUTJjgapAaVD8N0JgJ+bGotBqa+WxaTT1xRtIVDKWLUMOwwr9rkIS
B1DsOt1HcPppkcbm8ekmB5dLB2Nt2CZ+NZ8Agw52sxM64z8U20Ijz2LTP1TqQj8n
t4OirJOT436JSb4r2ZI950io1k/o8RXp58MwdepW8IToZQYONRDO4QAZ2fgnyJct
+jgzaXmHUV3LQQrqIUa8SwuHjg866byOBzPyrkZqCpJFah3GcjG4BKnNANaQyxYl
0/Xau+mfcObaUhUBGvq6mR79H7dSfTPL8Bqd5MhPwuSKCFVdddlFL23gRs/K02nW
oX1zoTEUVTkFzdmrIIyhCm7bRHEhUwRjGyU/sDSdaOXacKRgd9VbU8uAkCkAO2zP
lN0ge4AQCZwedy43/mHmon2Q4Qr4zCRmPXPptTuMDAUF9cpKOvLs/nIjMce41s5w
zBcQUIfeE9XQh/1xVRqNMaEGtmHpnRGZAuKvzMtPTpRfNd/miD+aPNnOlt16MfRQ
vWyQmd1t7hEAj/1SVl04BLuLBs7NYQ4QAX6XqCnl3DqEPQhABW5OzF9x5F+GBufA
0U9azw2slv0PVmKdqyQ5JAju+ytkHvstyBROYlvXZeOjnho90gWANCyxp2NwS7D2
Zh1PWe9TbSUJG+7fptSgh3XgTrz9t71+fXr934t+CPDd+dlG/GxYsRLHxisdLQfb
Cd8O9cssEScyLFiNvfvT8K4dJolfPtK/btNrIzfBwAHJFwYljYzooskm1Lg6AptH
bF2YB0ZExz4hYYc4+SEmHol5fIZYlrKgDYa+qy9lNkpOY3E6+AD/kpe8Dyjm+bw0
M9xl1IRdM4iA0Xv16jpllkndGX1lvOka8wRX7fdM+0NehdMTQkC0gB2KIN4s7iN/
IwVEduUzInbMc2EpbLpQ7cbuf5IaNtPFmeztlUdaPgZd6JXCbTOuNyyxo/r0l39A
G9yh69DbaIJGXLzLUyetsYSSWS7hADrwpacgTvZkYXwRsxqFmYtRyK1rxGTveqIY
L0Q9kYNGwyCS3X+duTg0SCNr1z0KANYmqTsGMxo3mLyWzjTTYjJlWIWTsOKs5w9C
apbUubFJ66MEqI2e3yVnCI8hn9DiG4jPd/vSKIa3s3Xzlax2M7XqezPUT0k5dqes
ic0fqZmXHVwdTH2Kcn+IRIzpvS8Hx0SSN9BGI2Ejl0ou+0GmoBfpZJ9qyy1vCT8u
4bSrJEWWafTql5w7vFupnY8adCjqZvqT6zrNvuOBtq/C/8hcU1qxUQ3ycxlBWjh+
9GFo6N4+qnYv3th1fK1tNIey1mAJkkxGGUzsyUGH2SryPx/CTW/SyzIe7shXF7+5
hf32qAWwufdHZSFf+X+AFiRyvlexswyDDUqE/Vhl3AAK4izWuK+gJflh1BAzLkAZ
QpxSIhjnTwT/caowBEGrsY8xG74IYF00pObmOb+aKt77WLmaq6KIIQLTj1Ejz+M+
wrvhsAKd+leX7HKXz+Ew/pE5htUWOt2Ibi8DtmAxkhAw0K15G6zBhqD+/M2f/89Q
A6T7dp6Lt9YQgUItmY63glewbPQNwtFmvFcdA1NzDx/oe2HWJtjlj08i7s79H0ZF
LlhWVQpUkuPV2gOEdHvtDdIGVYusxLkUAOvdDx/T+Zs5OtZEibuIuj16Ztu3sXmJ
gWP3Sgizjeiw+tDPqy3yfCPj0/7kSnmwpB+fxpguZdafwYmQBz7covyQbUSUI2I+
CmhrZprPqwv5ar0tlpiaVP3THgng3Lf1zud73ekvLcCBMwBwuCfqvRIekeKkCvfH
R0f+ZGFilf+1usNmHlrFK/GUcgAXzZ3mNdLt5ivyMBwiC+oYhMIhpp/Dp1wlNk3e
8xwnAdEJqcUDDnlL7IG0Wf0G25m0zE1w24+uirQqUJrkpn/JjULrSh0cTwX7i1pM
T+OMRH54iDHR2tmK7JlCcqAlOCKN9WXl82ZlDuyiU7ouN3kq0sweuNw/0pLaJ0Lt
UH3gEH6Ki13IvvBmX8IAi+Di6oF2yi6ZxZIzDMelfqHOQFmVFAkMz57SQZIZM4DU
vZHAqU10xafBgOw4KwE2IgaEYJB3mnIJ7/p/m9oQT7ZT7T7EWPAAgumkJ9ASfA1D
6lWR9jgOwLWg2BcWx1yz5xNkYD2r//uofdNZTQsqSc33Nwez/ulMkQhZW4NZcUOj
JpoqBHigHpWBpHp/OH2mkdZ0Xbl+Q4BkorYOIXXbEnEeyJuFWoJNG6kNlIwHiSTK
csnvjk+vMlpFMJeGC8hzkbVqQFE4G25Rr4NgQYABaX7xyW1C1NdqXwTj1V54i2aG
Ysq5h10WVRduj+6YEdHAg7IouiIs0HgTpHZ+pX3a95YmdYJ39xK6HkS9LBA6Fwkl
iXBBMk+XcukFc9AoYBAlhnFiA63Dchf1tJEUfXLoBx1L31sTr5VM38v68NjvUjyW
W548uhkNCvi27qs+Iksx7p8E3T4T6PU9GHw4ri5bt7vc4q0vq8Zp1NiMA6b3GaZq
5acayRersoh6Gl0QSExzQV/TkEEEZOD6Q5ugazcdk/LGOeqTFtiZ4TK2WsY2HNZ9
FEPiyXzvHJLGcFOjKA1tJ3lvNjFxpFzzQECZRvg/6KLN95yRPeKIMP8Lbl5AlA+G
KYEw8gBfJe27A+10WuP2NvAC3XCiug59oUpcOd04HMffjFlad9WLdp8a+sZRwfW4
8O1a+2a1GRyfKg9eCXZVbEv+F0//QX9boHDvBg3yxgMTdx1fgdEd6JIWb9v9iiDI
xtSqepzqOGpTBIq6nXnE6Z9K2wXmOZH6s0zWgPgyu2dw+H90DJp913+7Wb4DH4TP
yMTjFt7mwTVWltqL9+ljT0LQCLIR7m5QsszFRpV5FKMNELST21+hdTUOYPKtIhwK
wm0sUzw5ba21JdN0Jq60GgvLmHB7Oqv5swxdwri7UdO824iwOrX06c0Ms3HQpqe6
MAjQNVCsIlRWztEN2D/jA0HutjQ+UkvMFqDyzFCDm1nXrjj7sifxy0+t25zmcPm+
cNBOKmucp5vg0RkrATpUSZQKuzFIdmSaJ79NaywvnWNywAA4ztWI5f1epqGf4bE8
Ai1uOY7t18/6raa7O4sf/fyxPyQZ82n8JYDlFzzrSMlxvL0VmuizehSM4Wvioc+6
55NdSLTQhD3LUI4H/3yg89lg+4pakXeGNtp68uRZr18BV8KRGeCPRYtsFW6gzS37
5QqfNodthhONuCDZ+2fGx+cOd5ra5I4xRnmmh5LZBOAaQMIbF8NJJ6phL/yRY5nq
pXPu1cEUI1iVbsl3dZHybjU8aolfrk+VoLX8QGjp/mQYjuzG8u3LhNii4IrmYm63
WFNMj9WyaduNxgrhN5LM5q69Nz6Ma7shanxgFlWH7vyL/a5HQrPBIDXmCSC5CE7F
EC0w8CRE4wF4XETlyuuUVQeERSjfuMNYTvxMiaKkYRpaiBVCtzb+0U82wGQcLo17
qIlKOdZG7Pi5jSceFwwprpeuog1K+76RYusaakGx0IF8fylek7QlZPgEccyvDezs
tq04XPkZeMcikBoK4tIMORVtQP0LQx53PnSIb5Q9gJeIurro6lKAS7HI3JbZ+YQ3
tF9lbohE/0ZM/64LzklMkPxVlUwQIsatQduu1kJCTNZbVP6Km6UK6T3PKKvYTxeq
GNRto0UMNPjsw3NT8pExM2txASV0ghXBZrx9EijjNOJ1XiIOOdg+ls2MMOeEzruM
rl5aFNCdJzR+EwqfCH/FEJjeTjMyDM7KT1C4457hnqW3jv+EZC8RiVtYJ9IcBZ/q
wPMBjRI5gLgzkMRABxjNTAjj/W7l8UuhwK/hXgr7mUYNV+HdsG3J0V40G/EtYV6F
4lruze8ZZYtRw4ycijI0zV0nLYahHyjKT7pguAKtVBZIoG7mV90Nj9YOkwSH50UK
IMkM99KmaYTShVuBsXshHoLPrvhuxOegPX9mjbzCOcZ0TZQi5pUH0BGR6aJddVM7
EjX/7no3mvTwXYFoizEoqmmRi/NicEQZfe71XGLA+gm39CwcFeYBchEndqKJZ3nN
t02s43Fe5cN5KVs/gnb/WMKokaR2T/pKrpVzaUcPmaKVy7PLZcePpQTSsKu40ugA
dz+OLAlQq8DY9mdW2d1ZCwhUwywcCrxiYC9AQ/lEJVStLpOXZJa4Nw9uGmsftD0W
RLnySuU9qZmIqA4CS7lOGBRqKU1iHeeYFZlfd8WjjSo5B4V0o95naCDlvmc0hH4U
5nmunjRGexLrcOqgBNNZerMkdFN2N/iyhkMMIXwDlnf8hQ2UMZdxALuLLjgRBbcj
xuI+BW8Wu1ZoyLiul9qL5CQU3vhUUzKY4qVnEokRxT0IZttKVN5OKVffqQvnUCG6
CnFlUAFHsUs7HaRVnub0EmhRyQKbzfrIHAxEZp1/O+NF1VD73FvmED4Fe3onOPv3
vUwvHffLz1fdLyLkpmxP2uKO9dc0LVb71640OK0wpW/yWqn2GlprEvcLsDtDEz2F
zzcss2qRmPUh1jcG34Mxs1GSJGkty0HKk3Z9vQfxJuSaE7uMj9+avV8/fmVTvH6p
I8/WCw6Guf2eAmXxvuhEFyJuZXOvPQYH/3XzU1ojINcH6kGytr02BwEwxW3tFYYf
Ru0GFPH+aTi3XUzo8iTf9Y+0Q5YQ2tdx3XYi9EOWG23sTMlzejtE9xN3nBfv8rhl
51fzB0bmTE3uzqkko/CNnoJY/NuLSodKVfr5tyYuIdYn1MQi7q/eX1zjAaFtm/66
41J2t3mLRZmfbuvuH0vCWkLyNvHoy7qDgwkm9yIVeGtmxQ6dM8RpokpPdeoNHMam
HNKzcVD3lPGOBDWf14Fu33pzEXjT2DKhIjCtuurPPfc9IxEIVSszFchbY+lbE5D4
fWjnSpSR1XiheXwy1F38pjCRUP2z1vxmYhmSOy9Y5kpMuE+O9pnx3G7tPriKvLsq
vI72XiGSZv6SUSrzW6kLsbb2PtMYMGrnmJ2Ze1oXjEezaLblYeahlEXn/HjY19Qr
Ixf+AWV8py93wOwjCkP7x1hMH9JVJ0xMosaY5IUKPTDG42ENBZ0zOHMUEy7ExliF
WP1Ai/3h9b8yG9BT39BsYglnpGVD9B9QG6CG6V+7aoTMBN6YfkrMMT/H7DJfU6fn
LVlv62McUhFND6yGCco/s+LiqnxkPuhXImp1nCtEABCMdMI8A4Pp424C59FjuX1S
OJw6bUP2p8pzFYmK18EGLi77Qdc+k5zBPXwASEBNXJVAnV/uO18QO8YWHoY5sFWd
uprf33n4+HKQVhu1WdsLIaKTuSdtoKaGlHbed11FsAyOCi0905MOb9J5Hw3VsDsW
gD3qndaD4e16vIqE8Xk0tYrwsF5Fn8gTG34aztQ3+K5X2NixAa3KvrKPialZ+6yg
bt3Njyzp6MNnA7iDJacdidRTrNNwCaAgGW4R4k83cL2l/OQw+pMHfKRF+8lZiBUD
sVAojF122fK71l5Lo8rCg2PecnVC4ft5MY3Q0q36f2knJyL6zvrP+QEAQCxhRzbF
eg7IhzEsbWACsZ8LiMSUvwcAwgLlOVgSkddRip8kX3zstl7hP5cG1WgOn6U4P1Dz
NEj7Wbwd88yy93ujyNcXHQqnbkVVMvl1qMlJpUVm7a0VGb2joS88phq3U+K/UJvs
U1XwjiSSgfzSokE5JkS+tw6cnH5tK2pPyiufyrvse2fYKn+jdEdIx6itWzvZKAY0
Iw5VaPTTEQkmZ33CUBm+qTmoMSJCuNIxVLq/zfzP1qABfkMYFS/f2lgOCqSijRvl
utPZ9O4X4zjjFCa62LqD2fXbP5vtyiUZv8IRD2iOqNyLMHo+rEvuFU+RTG9Jv5CK
9PcrK+bvNmbIv/Fimw3U5CRi+dZUAimU909p5Xs9sedEeeEa1LEVH1hwRVFiJ+z9
lWDqP2drcj5FNC4EwaY6PS1wTed559KwZQ+Yi+vTBEO6x2liVlrHYjtOLj/Cp17X
kKANU/2BftL5hP60NBQND/W8SqIHCx2tuS93FrVYemMrEm/Mu1CGO9X5b+2qmSNH
mqW4Fp+c12ucYstnK565SGwRHRSdhsZy7WsFAaguJ9XI6gIqZxAjnkFQoUsHy66E
vi2gp5ZkM/4Pnn5S0zPTHEaY4TYsh/O6KD1QuDrlZ4oB0IfDrWfCkVdo08ixmT61
xi31p4kqMVBUefz+ve7EHcgGvef1u/hpNfnB+7i4eYicK5ghS4GsbC/SVCu7YHUq
uxc3thvTFKPq8fUBmP1H1uXZE5QMuACKgifLf2AqCwtBCMBiTAowTSRAkS7LHznK
/ZvEmYcXAf6KVmZY3u9oLG+GKEd6ZN+hVaAgR2s1JDQRbxg08deo9i2EvmkY8IsM
rA5YBynD+v7OqKfOUdEnUiWrPRgCxq0NKl6zH1KMutG6JnrffUVlFmmJxhY3Ja42
eZDHczOdLYaQ46Jl7p6SO9hJ+8tEO98LDygt+Cc40d9lIO09C3R4+fBrdXB9xPV7
T1kwTy6A7cyXZsV4GZTUDIOL+u1OznI923NV0ChCMG6TXMvUEflWvUpUkYvDFmdh
HTr8EzWxQBiX/jLvFAraBql/3+rZdn5gy88Hbfy9kHbumCE8U/rr+0JljJppnBe3
tig93p61hDWyiL3HjkmCcwMu95T0nxyvDk0bwwSv6mp9y1AzhzXzl0rVdp0Vx+m9
uQX0XPatUZYerP3Yx74uC2fJEi803ZGUCwHM9oS5yAyW1liBGHpqhZGp/NlyE/Jp
wnu2XJey1pysL1RtGb0raPK9QcA52JMuK2JWvMcUFSgqJzJ8sK69w3emPZYojFQB
hpy5nKRzn+Y9ZrBI4nW7ygGJMO7VUsiBuc+oImsM7exxQEGbazJe06IrNiCp8NyA
twQFe2uSZcq8mdzrHmhhHKbSqydylmEiu8biaojvi9fqjj7utaG+o/QMmL/tHElO
cX5hK6CuI2MHtTbPcAJyO5Mz3yiXqFhrdj9CEfT7EtgBytdisOK8hhSkEzepkWz6
q8LQH0k/BWTZsfl8rxeWVPGPv+1H6p4WI2q+jYQod4uQ6AohOtOYyE2F0EXiEING
ui0Kr1eFkocaVOe7r4YU051cehkDjgPlESCtFxw7pux8bwDwxDg+glN0dXACnVxe
9sHY8Eda02jTa/Rv44QCYmA+njLJPUb6O7dpD7qH1ceLY3nte+ykL22yhlMDTZkH
dUhfjakraiEuXoKKDAnHz8lUL1pLQjCtC8odca1j0zEIk+Kwb5F91Q3wk5xIGrpX
MGDr5JFmrcJ8DnKZDe6uj7v4KiX9mtPVa1Xq7tg31M+pd5s3Hcr542Ef8rQYWt0X
KVoscz507lYQo+7d62bdOjVcFmtUDljJbAvxXfmBjIWbTHEabnQHw8EBWz3+KWSz
0yem0kP0xlK2p+tQy1Kz/I3cadQMWt2h1EPy8/nsjvI=
`protect END_PROTECTED
