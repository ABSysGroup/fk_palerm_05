`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AYmuNkZgCeNIC0y6y2Nj+/HQqaTyVszOjcUKpnt2rWSEDcUHE2ct2p08nbL5bByU
+j06+hhU67b+EbuXZLh0TgI5QSlV5u+9H17BCp7xZ+ma8BdjasuhryxcHXVpZ9ZM
bZs/rXEm4aTEm79PIDQuS+z+jIuQWEPb44rqR8cmsyDZm5flefQf44R//Jt5Zn0F
au29E/8u0fmhZvt1WbFftjoZEXymdcbaBkjIa9VAJKM6LqJwGeQ/5a7NCuqfmDCB
ZMYZQ9ERmd1jp0ueLjOZRCg5r9NaWkb9aQVoNDz/1nR0AkqAT1LSzzjqSJBZBW1s
ed4L0MeKKjC1gBLRTayIWg==
`protect END_PROTECTED
