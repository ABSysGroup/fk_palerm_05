`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3JQGGuom0vNpwkAAjWIMWkE42MbzIO4DxdR6uqQYD+AtN9f7U3v9aBc6+1Gvptd+
T4V20LB0DWmL4NXorVKJ3FRCmQ8UQrnrwmy1d3ijId8+uzA/HkgGgVgOOLX8UHRl
l0SnXhWKXpzDPkDD6fw51nZeAIDWw3kgKrwbAwU8mNAJvzEmyAkYT2RRZBHMx0ZD
ikZ53JhUFitEtHwl6gmHWnb/cGjY3SNAdDzwYHjX0U8lAuI3nv260Wufri6u/1LT
KClleA3MkpwT5n5GjM9v4eiKBVqRQhKjn9uwPFvwWzluNbw5zJApZEz4QBTlhMaq
EdEBOYKVOgWA3+OTPQmFe7XYgmbkyDW87oHNsBlQta35m2aGXEVOU1wnuLpbWnXN
wUmYMcEIDQmdFOakRhF79UCAk6kxg0iN3y8wpNMAAP/hASxLPW6xK0ugmsNrCkRe
ybnJpMBprArViKmCXurAQ4E3yO1O6CpJhhYT+NWKbaZAPDSAQm1khRqDm0DUkrCw
rkl4BHMRHJNASBmXOoQDhFlFXf0qAMVNCGAnvByMH6oKQ6hfXr8gGhoDFVHH3HxR
Ya/QLKIdI2c/MSMCOFbFKg==
`protect END_PROTECTED
