`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A/mLdEIU6n8pThsHGDi3xTTvTHYa3eotXnEYqUBmhC1rWMWsK+A98WPWdy3QUaul
I2RGvZc529STgExnOoHRTbtv6MlVBpKCrPXixHFTrFQfWfODo9feaWS3NMjnLc+T
PfLNe2yYyoERkR/ns2WKBqRf0n1lniZCiGRdqZXW2C270UsOKIaypu072larMxHt
Np5WfPLXh3PoVqNcZ6Irb15uB47qrPLbmZja7gQs+cjKYNraeYTMubU5aNVii2fY
1vamFUqCBHr5xX/f5TKa7ivyrVxoip32CQtR6Y4mSaqFHf9UYzD/eiIQ+exs8qMs
eG8YA5pjRD7y8u09VlP65ruNJwih6+D4yP9daMfz3F8LtmeEPOgD7nbL/Izo+t6M
HnT2AOpd2L5B1cRPIXbQn9MDUmmUtdJ4unAgIWusZmKHfx9aZee4L/vI6cCNMVpX
HbeVFyFsIJoqLr3HNkkATJDpmPVJYtGQcm1hB7W140mAlmqoQlc77RJO6oNDMHD0
lHxyrlC/gNTPbmJfCQhMR2SKWz6CecJ+yBIgfvw+9ealvOIz39cHEiyoJfVQG+Vy
Y64whaJoiubU34BxM/aXVwxDzsNxa+qexpWT5UrgjVBDMaqX66jqujmBxf0Gh1Ab
1NLWzLdiF7ktVYSWiv6hbc9eTDXiBYYeUNLe6oTD7rjNIRQmwWLa4x7W4uD3AcWo
7zivMjcmTAxrQ/vwzzQp67GQ9oyWxYEoGds4Isjlq+eVaugKJLA3kzQTYkIw3+vv
z2ZbYHDjRLVZd/qmhtYcMFdjUE+xUzzNXqxrmNltGOWjDD+Zaspg08uB8p9GnCDq
rViZSDqeCpUufdn4K4PDD/HuLOuNN/desllWV1GPztczlh9s38V1IpqGv8mMZAOn
MEilK9CeVtpqZJ0FhRUPyuV9v4roIdfs+kC7SeBr7qSp9qnPRrRMhM93rMgx97DI
UxwGllbwEerdbI9VQCwgvuhtrZ7KI7kug5/w0UE9N50yhTQaCtg4PPZEg9kwUKCa
eSJqZCQYO7J/tK5Nzu06EKuvMbjkeAVqWlrB5YzV3e6XZw8KZu+Pfrxynt0eoZcT
y9eLVSdDgBXJ7XuiOIerxnras42oKGhin3uPejJc3aHQHuudfT+F39QY9czzIwKK
E4OVE/yMq+Hgi0cq1D++rYyr5xHf65J5qobsrtgWizq2N+XRuNKewpSt/4ut7Gnd
Xxo9I7vp/9qSRb4EuPYqvSK1UWy/8xo93gMvnrcNIq+IRiDWsV0PZVXklsEvyPe2
pD7e7qLPjOjN9mmTYM5R3V8bnb3hhfS8q46FlYMDaGYpImeRKpNCO8mtCuQNWU7F
g1Y7IT2VBvlG9W1G4aSEVdOKzGoOy2p6FIoCTTzTmENEk0cuW3zgCQz/LgldqxtR
4ULo0P6O7kWBBI/7xqQx4c4cuclOr8Jmlldq+dz1/cYwHUhI0+f+yKyb0xBb1E1Q
kbM2O2rGoedak0W9HLGefJaVi+V/V5vwKiHQPvF2nwvkeVIq2aOI52mvs3p//2lC
3MV3GX6+At/vJRRuHHHuusz+Elr06zY74mxVLPg4TDOJqNsWhr7fQlhLDKwNA0hh
n547qwB1bYVTA1DNQvHF6jhHold2OClidYypD8C9uJW8vUwaUSeA6nOnV0GC1SY9
Ul4bucD6+uH0YS3AGj1rsLFdjtquPLlneeleguBwHaa+9H8OeNMuwRqiaVvm7TFf
I2o4CK0GY1ecBWjpoKaAsMwNEadIuWUqBLE6a9+rjz8fJt+CcEZYjIRb1IDjlehR
eXX+IGfI+4hbzagMPLx9jPRNWWFhArkJzcTCVymOTSnCjh3e0hj4DxQby1QDxUHA
bP87wvYz9Lllnv8vh5840F0UsaPGkmfl2oESHr+cqp7zcfyWi5L35PXJt7i76Md0
BMoLjNjS1+xzRfo3hDR+hpTxkNjlDA3T2vU9bVioF0cJouEjz5u3iTKRTzpyVb69
iYfLwbGAwpG839RrAlpKkEzAb5EHHujuVEerz8V5OunwQNhdhLSehUeejHHArClN
X0ZK7zqMgDtwHPLRRBTVSyHEPestZLAA78lyka+VxKeaydtwPGBCMH1T/y/vBbAd
mf2qgqQbTqLsbMkaLWyCF81UBnsleuJ9NsabsZL7ZGRLOlhcSWtwWvzn7GmR6t1A
LAyhSWgKcn0FaIllJb4MvcpV85XlfyzDGNlWYi+XTqYhOS2T/8KmGzGp1+QvtiNJ
9+j/KR3Qx7ie7EBIfTb/8i0oHj+hgZxm1nbrLkFFAYU+c4Fnx6w6SrZlIBCUfwGj
4bElRfvDFqPMg8XdvGtDu6k+fIJdWC7m2n2MJEKQG2g8qMdjnmnvUn87kXWaTx87
QaFP9Vn4F8cZ4tbHchlMqtlpr/e8vwANozpIt0QcmaRt+WxqLDD+fIgnyLXExm2m
DFBoWLpW6biCQpNJW3+THkilnboO5VnI7ymPVGDh9NpzhQ6m0cDqz4MtiqIEAbZh
fagYIDmx6FFnSKEC16Igyrd/XU3Lwlu+w4myCEdwXexxPnCgx64mm6OyZBclsT+6
SAqY/jKhMVF+YpvPsyZj5hdtuLB7uNlPfjqNhEZV3KPVvCEY4l7tg3idcSUAwVPM
8D6LtHXOEwSXPZFR/8RfEHLegUVMZRA7GEDRZHjox0yw0xjsz7/+5hzUArBzYEEr
MV3qud7fj8FE6JHvwdqoo56sRa8osRrj0U97cZICcSqf9695ep9SlNW54FWj+zZo
gQSpm+ZHqlI6/nO9LZxCbo8k8ayKiQ/FcVFQ33TgTdzxn8iWxVlyq2cJ51SQYpRi
mmUt8CStaCANvu431DjJAM7EXCMDMLm4YjG8OLWvC3knENUKJOaVb/2Fe0uPsS4k
8w/281LjsVmtJOZXRaVqTF5kS8y9HIfmBjCUbOlYEopiRbmZUVGJel97s78KWtF2
5dEVYn0M1JYjJQ2H+GlPuLkCYBfoQXg7mAfq7wNjZv7GOZdYShaH7OAfVKdWgMIg
WeH3Eq/hh+EGhXEh+sY4nlyyZDAb104XWfgS3IQjgQK7A4nYaHh5MsN8b2okK6B4
8DK9tv5bVuOZz9SHhWV/RaN9hvZUHxDxk+Maoz7C4Bot+6d2X4os7CVQ/5SgKM+X
D38Q2uafrmgPJgdUQmYpLU4G532jjvHEQAnuIKXzNcRysRYnSj1FS7NSYAVzB8Ws
Q+340752DyVMRvQr3kheF/6cCfSJCGqgvGIC/YMTJDk78xPi+y4cIdXV0awyywzM
e1srxyo9Hnvmr/wQtnQvyKvFXvrYca4vNs60lRkpxy0aOCM011qMPoAiR3/ERKyZ
Vw4+/3bQlbXLDHxSNLJfG5ve4wvbuQxCnBTl9uqBZgPPg/P9pojO45t27O38hy+f
wk1V/OxKDlMgljBKjybBoUGO1BIfUx+qIwreo2Dx/KRZG7UZXx2BYw973dpGd/Uk
GJfLky0Ee+tiRS+5XXNK36gqMFleE9SJZOoZZQdJVmDQjMN3aPdxTQgJY6fl1EPi
qRuIeWUV4AbhtE6ZtiNlMO0rp+gFrEwQPNM6728PSiX69zoesg/1YqjWd88WpecO
YB6rw5vd0OE2THFINK4AsJM1RQAPquGtHxwa44e1ZS40ndVbCV2XJxWDTEAwKJGg
GnlGGizK/psWU6bo3DHXGNRx800xgFiAiX3OhXVJxP4tajtKHIxDPLp7enjIsDJN
otgMP+F9ws1+hwpowREmnapHfL0IjxYSLr9YPhdonyZFeAg4DUAraL/B+fDsATpU
/5I5Ri4WPwfQz0lTlJvZrcpbaX1npKRJPdSprFO/czwnHLRPxddbLjfyE91jN3I4
BROPRiPQ8j9VqtQsmOEgcSn5qH6o92A69+ge0+KnqLwyM5OohTCVTwXgowD/AdTJ
r3aVMeJrj7lblK4Ge8R5P4anOF+wrXfmGAW5kzsvbR26WqIgxWLVA9oUXmJpPmCb
U6jZCZVk5HcgBB5n7/u9WzAyd6x0/vlPbBaiCSycoZcH399NYUjjozXmFG9RluuQ
JsvSYGfSIcmsXJDs406qiW1643qmx7KZSIJAzC1FOF93yahJNZyJbzpDBHvUPy0f
P6nJH2tuNHdLBDbXvb3esqOXLK0OCOsJY7KdcS0xSORbCf3JZMCVu+U15UUN8KxN
h71+o+UmTVJOvZV1N0FmaDjQDZ/nkcupEqkTH9d+OZIW75++DHSePb8YA3ftrPTt
LZpq5xWewGHxZ4WpwLEeP5Eao3SPaJq15QGdarvD+Q3Vqpt8tV2/8MEp9YiNZuGy
sdAkORuW5CgscxjvC1qwjyECgbFbdwPvAesEoXTVNyXSPRF3FQmNWqR4hy72YsyW
lbgvAS+I1rjLnkiemZtlmaUrY2SQL6OoB6hud+y/6jeOQFW3SfNDBgDDX9nlbsDD
fVS7ItsthNZ0becsLxjzkpduhdq1clBqH499OHLVdGpFRbjdazlcWk14uQRONR77
5YMWZVebirWG8APWp3j8oUE8lCjapr0oLNNUpJ9WSDZmIqac9D9PO2jl68ZB9uKL
8xV2OJqoJ6lGU1TTX/z7WlII9ktW5DSJ9tfW96YJ8XW/FwCFD1HM50gBzz9NkEvp
0F4CFlz1OFy2s/3rfvz7SL2ITNdpXrP2MNkn9CcdxQEDeyPbCUYbg71dYPmFTxaS
69sITcxZaA+zAcKrEuMkpXMS8bEoWS0xLuNl1F+gh/aWeDz6lyHwB2c62laBho3C
ktZzDYJl07hRZNpWU1CtHGdwx4TFhEOKYsK/5oENzXZCoJgUbg5ds6uKcL9+q2vZ
`protect END_PROTECTED
