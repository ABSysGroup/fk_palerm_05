`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b7ZRHaYWNxyhMNqjcZSNWQREoUy9wR6jh6+iJ2LT2hj8/57K9fPU4MpXGVgbl4RK
mZ9L3m95H5r+zq6CpBghXoYikLF8+o8K7qtKuJjvMA6xOOIdpxGD6+atOGr2Hjwz
unNoSNY48cyEc+oVoXn4dEZAtJWnp2BQqsDTCVJ1ALnLQoxiibaetwmeApWdM53Q
OoHWPYzQ7olz9rHe6Y4p7VWvwNG0ZRvZ/2HaiM3CyBP8sQ0amAkSFFWxkEpLP4xo
CeFihytfnC/TvnEE0J9/dNB1l+AHe94VlCE5Dkoi79Au0GnbkiLmjmFu8NVo8Eee
n8dEGYgGSAokCRp1dU8W2w9pocb9IBzyIHoNYJpvc2Xf9huNHOLmgQh7EdFaduRA
JBDw934UrGNTwnvDmov2VCijefbjrsxJhm59d4BHlvYGhFdxmiwjQVCa6fSvmrfL
sDdIv6ti4tENkWmVx2mt/xbfSiFNqHWSoyXJV07ZHCnlmY2tVBr6YyyHlEHMzfwb
LUQDR1hxNeqqot+wWEglt99XASntkQTHn+PvLJW/SiEqquhl4xNbVXis/I54hOKv
onpxL61vHv7doE2/5EbyZMMqwzadp7MhWZStsvo1XIku+vzOoU3Fc5zQOi8k6W1o
IJ3fxe666SahxKKci5HtdrA3DxRjNRopecpBt6nvN4o6+KWpVFM7ih3KsaIY2bss
a4dEgDTxxXMGgZfDkn7STx6VZRVGqQLICMZeVFJvkfTuxw+/9q1+9UecNEVakAxL
PnMUbesQleFJw7zYkpq1UA==
`protect END_PROTECTED
