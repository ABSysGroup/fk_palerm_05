`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0m5My5FFASbwMMmqawe1SH3vOBltKH2HYBGwA5KyMDB2V8MPg0UBWP8lP+svduNU
HwuvXOSogWHagmXzHGMetLdLwj1HU5ukkLFvMitkmqvF6BKaQVyVJC+SMSycDjBK
yaQl0FZpXdZAFeoirSCacqtm7NgYJIftF6T+pX7D2NP40ldZhOIQo+E8qyHnVL7a
KDlijzZJAnSzOchHD2oRjWsRt5F7NdSKdanUns8M6KNMC6KZ8nNk0fJonVTz0Mmv
9mcMIz1geRRo38dIIaaB87dPXM6k2SdVnb4e7Acj4zIx8smsYbKrXFDB+BR2rwXW
nfdde4nW1o7TmxIQZY5bzdDG0YO8IsCjq05xgYaPUraIK2eeG0w43wP8W/QgTClb
h5ib54ACqZsm4ftE2QqE9IpvpMp3r2A9qdA4TBnqcE43elXwMbFuwHWfyKZ4zHfs
75VpN6+MI6U/BcpxTj3IftmDXW73anLTF6+CVtGWVNmdspf7gezZeVYC+FRwpMVR
LydlXwOsr8s046GuNrmxFr8GI0/GSxyj/j33FOfokw9JD2pmLpvgHjMj+AtASctw
fKl2EQMcTjDSYA9auWVpSitIKuM/JI5GIKjdGKMUtIGeOO05IQGL6fsKGCz7+eC5
Ur5DW2/rVnfQKz2vWIfsb1amMcp6LnM4P6bU7jRkrW8=
`protect END_PROTECTED
