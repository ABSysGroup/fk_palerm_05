`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Z7H/J7j1lgoEBwDenOXNBphAMmDCu7hfxJW74Hgt0qoEe48j30Y743i5mrE9Pnf
rXTevsQCwEq0o3rBU7pcHiMpQ8kb62gXV6wqip0IiRZLxLdZ1HusjZXw24CiO5UA
QWWvXJaD/7smodAxujlol/3LuNW3gDZWMz3UpFrg7VbWxRJ4V/A58Yud7B4CtMHQ
3LF67DteZyZc+g+/zb1aWORAMWimUkB/EdMn4NccTfhGxbwjv6XZO2TDzsfjShzI
kE+H+nxnwsS0BaQtHLZpkZF7ux2F6hOhVBmlOS/6ycihqT4S3nbYQSYxefwHxB3Y
vKdrRjxNIGiSDbvLUCUoU27CpkMKYu18Q47osKAhUuZtXzxaAtHhx/GNCgTYROqa
4wJexEgfuSaDFm4q5Bl8Vzp7y2AjWuFQev5z4mdNtzFtk0Cx/Vn7swkd3m2miIUo
6UjLDBdJ7HE5u6th2cCgWx8R34LYJUVUXes2Nq80FcwP/azK8EVevvMexzZBY9UV
ncMuChzH3g7GRz9bTLjcsypG3bR5Fkomy6QwZnId0HeHoU1K53LCIDn7iJbN8Uc8
/MlrJgIX84+RzZ/vySU2iM1QGYjIVYZXdGOY4jG16mhZQL9BUl/gVCyW28leBGAC
DMyxpLgvAz1LiHGvhKNsHmOVJBDKlc5dDjTdm9tKhwcmLq46YLeul887EkgDIz1B
FNUPepGlXFkhY+tPSCyuhkVGJEBRD6w/UDKs8Q4ujYpo+hhY1bBfkRR/LwuLV5PO
pZMGD/4rZC605kpe/aNRZuKXySa94An9ujfjtwOFIdYs0RKL5Y5Rb8aNZLUVvTp5
pH77vBsTFtxfdZU5WJwpmTqrzYrr4xsSb/JysnmaN2wbK8/yZhen23MAZPz1IZBG
avsilXhJqa+tRLTo+A08gRZpBRt4mnLRKXeakavBOoeRmxCV2RFW/4L+6+uvuRgf
KNHaGY4uQZYKAz5rtEYuquVDKS0mc99uubHJ8lFIHaa+9JjVAGmHqUuRbYfHKaI+
Jcr5tmmfakY79si1kyUNDFcmS6drqKrb3Wly1jZW7AbL3q/gCox8z5btSCa09ECT
nFEmORuoWQiTb5LK5O1HdWHvDJnXrt/67WAe9pk9kYRLhEaH+NzRsZqVKESWvVqb
Fr59GhO9sadxWBTtfDpxrOhB9rsllhcHN3F7qltucivWqM3gPpJaqi27yl3CtAAp
oz8iTTupyya8UKrg5nddPXTIII5PllSF16qNKbFwlber7KQesCD11A+ysJhX2UNA
xXai7p5wRBfgNotweiBbfM3joq29mzT+DigjSiEo5bEMbbvmqX/YHhdDfgNjrTGf
yYveE4Ev+dBGdq/ko15kS0s3YTskw7Lg39n6tPOdPPis2fqaB/Nj3R8Uea/zOT4D
L8WLCWABcGXv4nw1HynOwd8+dNU0xl+3LkBVbXJ2uD+ZtmLPzx8yq3ZpPSKezhtj
VhEI45FiXohI5LwMUTrPhsQpY/NURFDDcFpvOMq5wwGm/TbcTk37/kp8vL32Gb6z
NYUX/6gPXBhByt5zoKQlOw2CllEzmBlG1dvmVM6lkMfSPS3ryLbo7N2RDAYcxlk8
pJVpvYhrkftN0beiKkG28J5RzPcW/oW7IBwYROebfLHNl4ODzKJhJyizXdn6gmM/
I42ckMrj8F5HMMJGeNjmv924akWcEsuar9P3V5l+sGzBBU0JN46s0F1Cg86b2j1v
1HMBFApHs3l8BC3zukl+aHycXRjE89BCwLMg8MIRj9i9eZQNiVfB6bxklUk77vQn
ItMMBHSaVgbuFUSKv3rwK/sB/KP3T2z7/7BvbBRYTOiEGfSO34npJOu1M3NU5U/a
UYfJyJIQ6uhNbX78Pp/nIyGMJregN7Jm0GmCJKR3E9Ga7pkfcLmdAdzpTgiAMUmv
3RK6VL9ghUk14NApOdxa+RIVJDlhQVS8mI4wuYUHCPzJP+Sh57EjOs7NCh3s9Bqe
paHxVRVPmjMrAKmvBQDw69mwMPzvTJ6PNe3qyqwaSlaxEgIJLFbyYtKBtZGr3cSA
TpRzS5853hoGNLUZlrTqQSaMJaHjV21JWHr0hVbt3CQC6RGNX7CeWO83famOu7NF
kwbYf6ZzTFi4PP9OPbDBsMG9bt7H46yIZBHG1ImooOgWok93nk+AQIgORQXkiOSY
E+cA1TF2O8qa0sh4cqwkwi3R0g5KI/+kdJFuDjRnlIn+8d8KmmZp+FFZ1a7KW6Ep
WuQPUQr3rLUVY8yrYlDUEuPJJLhCyhodE/MyjkvvSZtk332Dy5uf6DRfe3Xf5XEP
T9s9wljbZcJlMl7ElOrrilXY9/BRvgRNfXdKZloiReWcDepe9ibnmh8U3o2JxRaH
dp6wzxV9l8k/1rXFCJiFwZgQI0XFMdbD1z9p+T2gp633GOFhTJy/s9ZVhxdCSvDP
stTVIF8JNhqm21qbDElHD9/zvYLvc4FoAQZ9BQj65HtkqkD1tTJdfHhkR+vIn03n
WdwMTXH7GidMT75lem8QGU2IohHhN4sKiqj43U/iiKeWSpIg68ns3HT49viLVbh+
MRQGlty6eOaFcCmXrP2P2Sa3tdTape2lmvYVDDekmgluPKF7fX1Z80vkzbWLNY1w
3REED48LOQHQw8xxeMbspMi8NLvw/mtteaXheLIvnpP1kRfHna1krskzqrdQIWOY
QWZmALmgGRcRUPc0h9y0Of1dbzXlnrLoxVtz+3lTSMXTxsw4dEwx0kG3LCnfKoSR
Bx24B4gikRisavhdjgUreZNy8l662pm0WV21+VImZNt7+pvs9aylUFXcpwIAa3Aq
TlcXlufsdC2/CKiT2lsixOQETyaU3hjz7G+5KD5fIzpdLTLqaOMMOKdqRu1dda5R
Wpc+kpYCqsfzQB5tV78QkIripPX5Xso86NqDP7ca85t5iEsXq3oEZpXPYq5ZB98i
7xf5h4vYQ6vjGmMjsqhiS/CAgNtqL8dFLa5XKssKIZngGta79bBsEVhPQpylbXsa
lYcEzf0YmwMN2Hj6+mBwRv4VjxzZc7gUk/9pmv2Szwko/pHjfk0ZR/WfkMKjeQ4x
WPW+UDiFYrqWWV5peH35x+4lSuzOQdyU/6WTYXSs/LLT/IxWQIVM1pf20OOqVQsx
4zpMP+Eaaend9yXxyJYYItBt371Pa5dpklCqPhOZDZL/fQlXGcDQ+lFPD774ve8b
WFvfdUX/x2vKn8le5vjXlzs8JXc07wBdpX09zc0tBFd33pgU1ztzdBtFr4NvslF9
AG8+cactHqjzhb/l73hb1DT3812t6T28iyfg/WBPioNgPjdqvJsGzA5dlA4FlksE
MOW5NUoi3VAor43I+iMYrH25lvRF0lOaTD1cxR6YrDeBgPrMeXHsVVOev5uB+0Q2
4M4EjuA0Cpy/1wrn08eTjswe2Jy8+H4ZKNDbO30D+FHuE6QCn95G6FUEB3JyVhYa
jOhFv4N4UQPd7b2wTNSBHwH/vkGPmvUlT1ZiQGVjcyZ6P2fqf0aBl0czkInlm9l1
82YhRnJUZGpfvrAHUnVJ1H0qNbfqT5rwTG3vLSxR48m9Nzp+6pkibAwI6oGyM8WP
vt60CDJFx+9D687c+nzkeOrrNHDvx42ZIddyUnHbV/11GGu+Vr8YKgDOVIcIMQj4
D73SUHUZTIfBWz4V1IqlreDqBfw+6/7hpBKsijqJvz/VENp2fjmprrk9T0wq7zhT
FwxZhj6JzYUUCU29xJ3156DoZy5KYe/m/ArLaIieQ5nACCURZ61ZmJxv41vIE05U
j0RJZa9UwBF/EHhzndryfqO5Pcbreeza0ASt6lcup4vBXPWF+MnZbbOQ3yQO2SzO
1hEnPk+TsE4iAUKA5zSlDolMnXJyFbDUq/Ip52T0Mk1fVcxMFm04gtq3lUfPmTHw
l327CHSXJYhVVR9E3Ar2xLv1JgebWfOxCF66KXKVt86Tuql1s1vOlVtQReuWbd8L
AkYjjhc1kW9qBKh12nKH+ziqwazemvyYVzs7cFxyaY1s83TVWVDHO5ekmBIVDBO+
Uf4js5uH4Iqhwc+JcA58yt82qUIG/LeLEB22MMD/eg78hxiRrWLU3O6wAOcIVRDA
U9B85I/HjOaya+YWoHTA09sChqPeVut2JKtQ5l2Uac4TkGgYM8YnP4neCSO+EfIn
`protect END_PROTECTED
