`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a6cwa8wgX4eAzh8eGs8e09wd0ZbirvgJ4B5dsgWXy2nNSYE0HTrrr4DPQEewUkyD
ivEc5+TmEPpIz4deWAYvDLNzDlYdhXEL/4AY+RB9fpYPKwreKB2jHTSx1P2Kisxg
65IFGlHL3OxCF6Rrhvc3+X9DEyQ9mET66JfteEWDgQozB62GZkbL2sHcyrB06ApO
eDQYWK8yjywiEHSG4jUFuSKootP2rptx2EmsLrVxxJyEVDGeEZwa+WKUyNB+1rs4
j8iYx5yAyaeNLNhBwIAYzs4EHJeQI9+JHew1meiz9HYuLFKgzZCqnmpYOg3CflVz
ZMd2bod7EvwKCQCXYpPjOg==
`protect END_PROTECTED
