`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vSJUWJmcUWcPRPvrr4OzcQx+Ovi9awTtXCAQf7hmVQYcgyyb6fF87oXsOcSLg2lE
0KL4UFSPnF4tgcGt2vHWsL4fWuMxe7vCbMW2MHdPpV+3ImtigK/oGjsNISuX3qvC
KK2qzgRY5+jaMWbMij/QWbewKJzePnYnFB3uyPiunKSshNmLGzhr90AzCh00qrQJ
aBB1ZwuCKoUAk5Bxf6j5g83XolVJXLku16m2g3d0bXWGmjmTDRo36c/Umrtg2Do/
TdQ8rg3HneA3DWqGXbx1S6Z5h61SNdKVJ+rNUo5zR3MeNJR8QETQYPsy49Jrla76
tAuWgZGi8iS4zOSzhxxLJHQD3vdDdhtk8wWN2jvenRlBWIL9sJIcvJH7vNM7gkIL
rYsR0dhKSftwxob+lGYai6gCHXOXKwF84dn+G0Bc1z7/T1rQxqzdmhIIEeAxQhOD
EPNOXfKgivGtXeVQfMia9HA+LRgFN0PFAERz38ZOtqgJmUn4UapYsX9KcjgbYsKn
P8Ha7WRn+Bx4zSu/x3bBaSXVfJ4cyzzH+2gcQMt+NL0kOvqGJwxWEayl2Sn+XqhU
FeaJyfmzRzHB0VfVXer64upZz8pAMlK9WB4gFKrsPZN3aDoRTAy5BLU5a7cjEFdZ
FPf6nY15Z68ZD6djKhBtSdY33Qkd7CfGPX+4E18LFJnjLFYkvhzvBAeyG677DDt0
Vgm+DZf7Ts22fyRh5alH+mPFv3psP4UpCVjMFLN3p0xf1uziZe+jRyBnO3/VKHRo
`protect END_PROTECTED
