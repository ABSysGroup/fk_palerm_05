`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AQrsX76MI2nJ01fZEQkGcwMKsNU4wYRvoiY7W0/E/RTV6curKOZjwFNNezaAft1S
lWLw49tiIFBneqxcwsPQeCWifEirJPGWldWvP78jbRnriBAtgyj6qMW3W/WfQum/
HKEx86ZG1VKsgJ5l9LNQs9sDcyFggOxbiI7ADXuaQOuJF+/oqksNiWg7ha5c2sfq
0MNwtXsmmlR5fT3HO2RumT/PVN1CCYJn6bZLT1voUEfUjfGE4GAHyXCDDkiXRZRg
4iEJBIfsm9PxjcGOCF3JQmar+mnOJev+LD6coIxSQZS75/b3U3ufNZnujaSHFr/I
Z35LrUG2ONZUVIkfcrPW2itDcbEl+mb/rBfUHR7gCCjPhEvzsODaDQpJFfHBPXbl
S+NMWXTQqu/k4mU0K4MGPxaC5w7dHfkWnt1n1yTsKD8qQ8H5Pln+xHhfkitHfLa/
zmTNA9E7rSa5wFhuzaijdmV4+4jiy4DzwtzWgN4JimKPCA12Qs67LrCZs2Fd84b0
R4Egn/MF5Dke44Qy4nueDdyDz34h9ZSQDCHOY16chnl/IPJMd3Ru0QY0/KzcZKSL
ys1BEnEDbOALW25aRiPB3Q+g4NZI+y2RFwqAb317ylIXFB8fl2MhbYgLFzOziQdP
y1PNZiU3BwWo8FNldfqKvH86UeReWqp7+t2jfNuTmTHvpvwrZuerILk2WiceTREZ
5I6WahHq5QddWM+eDFjeZEyq9kPmD2hWcZqb36HEReDpaplyKmRRMXk5q3KeJdIE
U/2WX7MROFEp5wJhDewSDyiucemu4J70W9fNdIvFVfD8+A9Zki4M5XeyuAh3OPd8
0DEFuav0zIgBmL0JY7/deNKgIV8316F+WXn8ylFkKM8W0koOF/bIvMTeHUthCxVe
wuEyItkAGJb5cM52SvVXn2Uld8oCPRSKXwrucWKhEAYVxBTrbrA1W6HvraIz7pXF
vCUWZN4XoARmmv2s/Cr/UybdUdEb6UZuuzQ6r8aMPa0eunVvyxa4WE9twtDeg0Mj
m94azVHv6KbnmXNS6NStj7XIst7jyoAEaKmriIBUmzdowR7Fyl1AxPUXQ9CLYIhW
lXIWpPIQUdousWWzIpK2DlkGZW6J9A9+arj3M+2JI87o+5mA04HacmUit24C/S7r
UBLymf0QBcA2YEud5+VYhTpjWcIwx2OhTKAruxG7xuk3AwkH4vho6XP4Dk0oJG2p
lLWBXB/FqT4mFWWnJ1Ezut6zyg/Za0GkopoV46cd9zB49eLjeUERKCk8Q/eNZTVJ
P7tDIPh48gtoGQyK881pTncZarvrw9zD6/fOwZJznCLvTdSel6DxHZg5MmcWCqCH
8FjlN0PSMY6NRfAIn3p3O4xHjHks5c+DklYax8CcuCiJSO5GKRHSozEzaLQtHaH3
3G9gIEirXGCxEMt2nadYHtufZh7QR44Xc7tzuJwM6viy27H4IY+wIBdigDwxFwed
06alccNpyYaM5klLtGesQ8BbwtL3xqsmjurYnsOAXL4XKeDQi/JMMnhUaBuaIzAz
H10iOGvfrdSnc6EeLhR30k2frrlNLK9mEccULyIZ59wu5sL/FEU6/8DU9CGHnNPy
8KD53n3VNnQMEq6VLM/wr9M5d8e4TNESutww0NLoizLS6qx2oL1iw0Rs3KMQdn3a
vZXYCZ6CdXsIt95v+WUwg11mog5S0VKqumhofWEFv+q9whFmhfh3TXzyVngBv41v
BfcXj8Cq+xSbljQMAG8zuj8berSQWGluKRA2Y5oYHyXliZOmRpa2vcP6OQt2mcXh
RMu2qYiRVHIMh85+8HGp8ixtkfAehZlS1BFMnN/VwCagzOEum6wUHqXcDOsHwdOw
n1qSGqfeJCF5LDieW4YBJ3pbvMpqOJepbd+Bb/fFjm9vYVdQdXu9KidWnn163ojy
4UhF5mUmVI/MaN+By5cdVdbE6eaU68BArFFuXf/sLGUj+mkXU5POBMdymxBHsMW/
nGcG7i70xlkEyTO02/9we4LuLoA4kLKGZC2isODFchQGgGjuUrgfXe5pr4H2gmZ1
DpA+LZkKMHIbpv/ox8MBURn/qiPIfVxb7ycN6f6qQjnbgYlciNOF/leOinn+ktt0
cocdDP8IWAS7H99i/47LBw==
`protect END_PROTECTED
