`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
prUeYi7f8eqs7XMRcu2pKcnGveiqYLKEJUvZfQYPnJAU5IdFUXXSb/EyJeEqaPQo
5a+QdeiSVGpxcIILam04I/eVt0HC0+ycvxtAR4QYjrKpU98g+uet9mYIfL4RyKGp
eZiRqHoFg7zO4Lz+qbZ7NN9fDocSD5726YBqV0hnXupzxfxDgbXyleMU3s/4fUIY
wb1EM1qu0LERuqbFYDG2xTtS5vRGD4B7XE/MOaHPHMkUdN5Hrrfln824hkkWRfDL
a0/W6upYLeK4Bn3GzXAKSavlvCB4zj1/bpWqHbYIcoPxuZag/Mp1b8xKijVHThig
AYNtjEzAZ1vRHsOaYZZUlcjSwDuxpX14l99T7I6NjFGLatelnqimnZlYHxrxyndB
G+vHfbI87Fk19KpjAsjWp19ILOqUXNpGRH4LMig1EZFFgppBmdbLZS/5i8+l33ab
L8CXbeL3D2V742X7RJ2jGw==
`protect END_PROTECTED
