`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pvYW4X6Ht0YLJjVREsgsQgHETJSl98HDEVu7q8Ie7TpYiAnYNN2rZlmq9y/Nw+MT
ycyPdtwIEcfgqm2R1JcE8/yUXMI2LgOJ7UngFuHoZYw+J0Fek4EyroZEjze43k/L
7kBOGV7vFXf2pXL+VVnx3dqCZNDJeVKPW50MxA4ogmxKPKuhhHa+xAZ6YyarD4H0
HmKRJOZWKBWAeI4C+RiKTtxSyI5MT2s2snhSu7wHPlo47/NHuC29YA7jnQ77Dwsm
ph4NvrpdNZw/dgTMCI+NpWiHjoboosM+2epz1Mc3Sd9fgJhujnDMi06H24KMWEdT
waIJ/oftinRUV1WDiA1ZyfVzwoDfr27aaor5syDLhNqbv37LXaiqJkPOnvKOQTSs
FxnFz/BRpyWgTJ8s3NXMPeYxtavC9G9wCOQi23RQBdx9WNYvqDiTKbj7If3glryx
QfWd3ms6ZsvW2wWNrpIIG6mzR/B+f3iHESN7qDJbQoJ7rmYmanZIbWO4W/cYOoLc
0vnz5kvyd1PKLQCbKbrsphDQe3gSWleCoIJ9tdFtzvTNXEd6IjH6M1Fy8PTKA7iV
Yx339L8QcZvTCFZq4nI1ZIcDlVplV4RG9ooQz2IWX64+rxM6ttAJi+P+qR1A1KXv
KJBnZkJQXZr4I5Gy3YZwAevd6Jp7Knxu+tzoEdTXHZGUBTZVI+X/LeigXibnLNkz
EwY7uRE4zqP3NAz03gkBG4yEQuoarCfutl3WQ/BzBhFdFEhEWSN81O3NnKy8W8ON
T34fYom8+Dhvtx0WZmAlcIGwgie3cF4vAx18LHBqBWTMZfKaUIlcnWAwxePEXPMp
oBitchMBfKX7Hh4X3w+bvd2vr9017Ehlac/WOlEqtLXlROU1Yitn7q5UyD2oy1ph
eRyTG+fW+laRPSkLY7bG4UVTHYqw4Z4RzC7pfOLPKqyTFsUuYchmQP2/PdL8/KYG
txItNA6JvSvC9kX9O2c5VjGVPfc2biKQfsZluwDVHbKL17B/qdVYE1rUVOOFN0j1
HrwvkIfA176jO8jY5lX8xUHeS5f5mLiIglT6WBVnOU48zwH1hlBI2f/VNVYFcZmo
cOq8BOPHfInbFBUr4BaKfQX0tvQTpOM+91AobcOLhXBjaPZoYogGcq+IVq472Sfd
uwmyPd4GzCDNPUSJhyVT9BAvNfZpD4v9sZXODmOkAeLyt+QMSbeF6xR3dCDeqitR
dsUB3GtfCqlZLqkUwgvWByjxvafOEDzJ3TXc/u2FDPcrycZ6zotmsbEaiWQb6tFw
hxTVnMskF//a6IAilY7GZLt5RA88u0gPrE+9+Mybj7blZoBLaF76PwnSfwqkervY
E37eVL0KHtl2TpEaGh7rtkLth7rIgiqiTMTSTzDZBamBGelPQur5vrOP7ZFo+FpS
`protect END_PROTECTED
