`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5jclVuJKYvM5XlfJ8zEXVekhasutl9yFMy/rM1Js4bNRoSXz6rirOjHEXhZtAnfs
TNwZ6KzUmovOQW+3r7WV2do8Bqavm/g8xyGhG8zdLYkN1IZYQ1cmL2neO9b83BO7
4/638A9EJwCl6RTy5vAZVfmA21gnfeYysb0gNuPHEKPfgMHgcjOtAjL8uD/PVfnA
NaO3QiQwQQpWc9bvK+76jyt+VcghgczDAZLY02TIgd/ppGONtpK+4ee7dfGbzKAM
qSNW7O8Vwj1V1cazGZGbqvl3tKLYrE4spUhChzP0JYqpC88mJ7OWC1k0uJOqkXl3
hgcn09DfFUo5KwyWD0nMOAYjczunXCvviFGAbd7wR1gi92ic55EqF9G8+pveTzto
GuYAQKbgEEgxbXabh5OVLHwXGouPOLQTvB6U6XqL3fAesvWcAXhdSVTEHqRN9pt3
NHtrW9CtQ3FYiy1OX1V/qA+SlE8MA5bgYIkTVdYLzFn8xajNVSHPFGkc0/MYquUW
KrlV4mDk6EnTb58Kl4vp+pUI2T3l0EU+q56awBEvAUJ9fi1w1XGwPMGOhkBJ1pTo
QgHPWvx2OmWhesp7EWE2P1sVCLOpNiemHR+1ouenSJQIb5Dp06R+AfLByVBjB4ts
ysSZQK3lPxB1jcpoNxqGe/bu45mVDCOgG7xwYJSGRwQPVYLJGBX9dP+iMV8ocoR1
k/ybeaXCX6Q0Xg0XchEkYVlINpFAdpaawvJdxvHi4J9ojLoE3ob97evy5ie6sOTT
eT3QgOKXkoXOgHcu9U25IX7aRKv8Zy+Q/G3cGT3jixIL0MkwH0+ST2k58dy8iC1L
VDiFS18rKIcnTqJW3uIBK5WjCa6q69CpPqT1+2e4zZEmvX+FKF0gS4JVS6Y1Re2q
g59N/U+Wez2KQktAIl7HZ4PL5Y7+44SjR/sy929xqnR/yiMwBrTGBgw0/UDj4mXK
mGVdHzQaQo+pzKIYjfepimaEKGyd/ySjdQksJoH18zwa5D12U2c7p/K09pAik4t+
8Ke74wBO3/kkTVkDcNdtSZYl5yN2jgTVj32813q6WDjbndr9TaygMgXDUhKTJ6vi
hiw+qJ9MyH5NYxcLR0WIjPbakv7uVRUBIRIR9E7kUTCTpAeQga4gvyv9mh2a+P5z
V5kACpNnkQKfcPBWCbtUs1ojjouljev1FIgxADwg9yllnpFpUSbPqjQXoC8ovT/Q
zd+rI2qwPXYldZwNxtL2KktJgHpqt02ZHFNG/dR0Dh1Dz76ybbwISTZ7qBdt0GLS
ii57F+6D0z+2N5yxMeGmb4sw4r8GXO0mwKdYJnmTX9BLR8yHT7Husk88TBzYM7Bz
SCtBc7CxUbBbTngZjQ8ytrNEtfckgd6cEergRuRGFT9LgYGK51rMgVtNAm+JQ0pi
CABqomKUsUZ0NzRbGtZqSivr/zg2V2gCMjxShdL4wIOY2OCbqGQeq1Eszqti1AsR
PxXbgmzPzyx44aEhjwOJYB/Q7YZPG4sbGpmtCOu+X2fTyw8HqCkDR/CcBW+t1IIW
IxAdov4OWv8ZU8vpjQ6p/iUfsxX/kMqVRiNvHBKjvCngCE77keMeVAnzqqsn2ILs
08YP5YQ5q48qq9VIcXd6LQ==
`protect END_PROTECTED
