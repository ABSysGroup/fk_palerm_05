`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
my3xJVOYLUmC6Q6i89C4rcnI1jbqEgK1oj267z/HBy6VvfLVmvNDaQbJQPlM1QDB
ch8+y1WNCN8DGjEOCIsbKlvV+czyYOwqpyg8L9Tji9dMr8kcv4ROI7fhXZid6jIX
lxI3nIB8N0iu9utSDlcOgqoIoBDCEVZCcWhE7Tym3V8nE5JJmuffdtHLJDIsDsYP
+koZ+ibJ9aTcH86NAthdUwoYl3MIrxSGl9j0selkoNKVSdoySRmEnNWCmcjjP/+W
mPmo5LfnEZ6jVBJR20MUdussCgTJbZH8tBjt5jR55zM6UVzWxcvYJ51IWdzka+iu
A5iDPFXha3ZsTCdxsVhiQ8vpY7Fg8MCYf85IJHdBYD3ekJougV3WnwCz6z5kKTO8
wH4LJhEU0bXw1z8Au7wABXof9f2WV5cmPMOlTcOdk1NW9gmjmS8jnNDoBBO+fDn2
gneYEM0GegJ3HrHLMVUoV+IyYGQWmTk5uYfbkbCDNbq1ls1rSVQdqBiAxOrR1KSS
gFwdDSMQqAi0NcFbBveLTjP/IdUQpVsgvIX9GC0eJZE=
`protect END_PROTECTED
