`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cSW0ZEO90GI6ol/sjjYSTFKiID+/3JpFZT9jkSYuagDIIh5gC4nexwlHljs2K6YS
wKM2VS8ETdv3vr+Mq4JQP7MfxRw2VXPlPVsLc0Frh3VP9Bsz7BGNVeJBR1yDPdmD
rWldShePkoFO9o45jQQ5wMe9n4bzY5Kgon4eHRHtV1sB7T/DVxRgDqzCjDZPp5Ec
UUbbuTP4Mu357KdtkKSQGe3qztNKBhmas3e8A6qr39p5MmrHhql9ihKf3I6vHD46
ya4rXEaVx+ggNn6UmP5YIlrvcrKMDeIVl28Zapw8GEkzkXnzSuoe70loLGuYeXHD
1ZhLGBLYEbQCYt0XCBs3hN+229IlEZNVJpts6eymp4+yJ+x02gug0pJit0igwvpy
4VXtCRt5Q5EaOZZy2FjIa1qyX6buQ4HRp2iBjgYlyYzPoEcf0JOUv5YeqcbLVEh1
fE9vXN1/6/2iHZgEj+ZNyCKNG26pWYYkLcJ0t5koA+a0IH+iDjqgmHcMkm1IqrJT
RKtzEju0GkK5BDOAs++SwX4BityZUqdjggVLFfh5Vq31UXhYL7mg0plidukmMXzL
vzHafC6PwYWTb/792hxHybalYtg6DlYGxoGR7KY4xunPMneuMnlhL8B57jOHWbTk
KmX1Xe3HE95/k+U3K4cJDfBnsOefkQCGgPnLxWBnnsiWClmZhbtE10DflECdfE9p
aOkvZVnQ8sD9eo4x3gXgVSrx4+8I7QAjEp5s1gdyZwMGGenRQAgRmRj4mnJTJAf2
FcRA/nBqUEP7PbUfYJf05g==
`protect END_PROTECTED
