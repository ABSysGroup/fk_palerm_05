`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/e81nvvjk+Tdq4+A7HirOz0LZACffyCp0+SNmPot6TQBfc4dY0LyEwkLTTV2i63q
+7+hD40cOAm/Wc0X81RseS/lJQmkCdgypVhLC4OxmnvcQbcWbERjaVtIT58FdTzx
sl6jPleLZjaZnnbNgNz6TUC4tzk+iMDLFxlipV2GdFO47LgZCeGAdEHArgIMR8Mz
znxtiE3t1iBUrYBedUKuhNepk9a9GAla3Zfh7QT/RRCdtaSVxh/eC8zxZ77vJ6qQ
WdOMei4nqdgXgCKB/whPxY9wfgNyUtKKyeEiRktpitIXwDDhP3yiUg2/E3J9KRYb
NUnMoZjQsnXQk0SZ/kWDLyx0ucoqkelw2a+fL6PtMrUjjj7uDNx1bBHz/JrxYDWq
HgZVsbBLcHlhXU/kmqmoG2W8wlU6D96mOfp6Xf8mVjTC/PCHgCEFcZ/2hlGxh63M
1rsp/KllyOPqHZ37QBvTrh8Gkc6PLZBZKk2jac05fcjCi9X5VmRwBzith4rkyVTu
RCxt8MgKMhxfZdrULtMTCZakhRyVI4SQOfxt19uQ372fxaPSzT2e02JlGNJ4YMKb
lxzFmfS8v8ENIFQF1HmhGvDKMsrA9lLvpnhnHzn80a0BjyLBjRFwMTkbjA8uGCBV
DXHzMKWmGotkNPaMEkg7kMMO/UOHH/2k+5AH2ON1aDltfZRSOxNJcNRiR0KNlrKS
+eY1cRfFYjAdhX+2OavaQw==
`protect END_PROTECTED
