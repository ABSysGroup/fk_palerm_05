`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BFKGqquewfH/y18+Ka6Na+XVAF77/zbRtxBOjRF4MOrAHOlFA1xjECvGDC2eT0Hv
ZqVaqpR/aLbRurquK4bhHVfyKq89mU/fSdgedKVEXkHyGU2vWGjtv3AIBccmska/
46P5u11malEZ6iVbuo6GCIbv6JowRU2pPQMdbNE1mo+wnpQ0171cmCoqvRvasR2x
GX4W9WVoG7sQcqrio4J2xoSNyl1R6+5QalnOyqBsH5YvzsHaGETOO/CGRcJnGCeK
w2ucWOBp+vLQl0xt39qNY4qoK/m/fQ39WZcNGQ7TxBYrZG5N/Fm77J5utImiRwRX
G32iCx95piLS0FCOS9TVt4PV3BwnvxrD7httzZPjold1eEZxy5JBjgGFBeWv3vlb
U/2FHmT++MD5/QiD3m++lw==
`protect END_PROTECTED
