`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I2QvsfmI2lVsND3StStcNFzb8V+YPo21PhFztdfg+GkAeEhVxHmw70kefonooiCZ
GRh7SMcwAY2489h/mS+XXP9WQhpGYHo8Eg4Zbt5nlQrv1wrqdEpkMcf4GsWGg0r7
UroF1DZKXF1BrspcvtI/e+jmondAbCVCyouymDbd/vJPhIIw7BemrG53ClAOb4ty
sfB5wWDkU8gXpmK5AssHbHY0PmG0mFhZZ+eHB7BXPaBjQNSYsBItBEay3srx5gkA
pZZR2RbG1U+BlIG1jHiF+HNtfw2fP0XBM3xyPFfuPmsXFafGeA99OLP2XDX8B9SX
gU/LMqy/aiWnZHq2R3x82Q==
`protect END_PROTECTED
