`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wZu+AVtIgPleLGHloOSjKNUTUb9KQB0fUcsJ5plouDmjp8KgKy28b4NPtvuyNLXe
VieBpyLpPM/JCJzvwz/hj/eqU7KPN1aZUVuvYbbMKsjOWlYRJgYzabzBGcM/2yhP
TrGuxn2CZtsVoWlP6SS8e1D0OMcHWpFQUKrQyacEMGstFnJpoWuCVQBEAn/Z5XRK
/P51KjgFRf2Rx8MTJ1E+cFobDOo367Smj9W1vRTxZ/FeDqK5sEyRmAKO7vU/hVho
yrZ/Q2aYQSBZTrC34I8JWdg9duJ2tiaCTR3KBXAWa+R7ouAIjM0QXRbFqyhjVLJU
vbbUgtFpejJTpdb9iH/HQSXF6tcu3f8w2Ey+tIhplBkE/SnbbMaKAQxN6b1VByp6
fw6rS8wdZro659oWT3A9eKCArg+ABDpUxkk+Wv2D+XohtRlFXYDLmyRhv7In2I1P
IMDzXqcMNPWcm7NK1ECF5OSthrwmDGOQ2JI8qNjm70OBTykkj5wJg8GqyXtL8aAQ
8aHiAk85yn5QCL4VsaixJ5tsjUaLFBPD8s/FR/JxykSITnFKzzmUCHyEJjkPEVac
gvAth1jKd7MO6NUE+HVJ78RbIACneolsOEpFTxG9pQQ/PBkOzTpEkFPZv4YhNRfV
BlDHpwGmEyVj9e0adZSGlzLwCZhOm6Z8Zurz/DeX3oTtQK6N33uMRzxdQ6gG2YxN
KSCXo2ScvDCYelxrJPrORlVnzoFm7T6okZgUP+7JTbx702PYpw5DdJGjf3ykJXhU
Kyk+bhW2Wrr7jybwTINr7rohyA5rROf4kG3YEXLOe3ZpjqatJ35lIPG0ljrDeO9g
VsvQyRaXacyOXyYuRiF1cyydLB9gDEcXfYr3ccBUbErAxrgOymTlPcPrGWbm85dq
cwUdMNCBqpHTZYNAS5+VEcVzMmrXrsBvG9jw9Yrl3T0/6/zHB4S+N/oCNlLtGGiP
e169QSTJfBAbRFVgYK3AcvvJBPHHr8CI1yhLy0kZXz+oGhlM1wj+6xMsmLKSYZCa
`protect END_PROTECTED
