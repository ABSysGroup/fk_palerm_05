`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MAz/VoLIo5H2fhMW+eE9vjtfXOLxAoMHDTmC2CyIx+2aNa4oNPOokFckD6H19Zeb
toG6tWXfEsYTe1RpwU1gcnJcXo3xhHsNMwIWlGWkQ8rq3oXKKM3T5HSbt9Egj9g7
8qbkQVg3wFftoySnnEYlUcGrjpV+bgFjFD6AvxY61/9UP+UgWtVoF/cgyTMtc14I
5nCEb5puHulgux1o1Ls1QoUvoeIVMHK1ePMW0IILQfLfiU7XyGylbulOnp9Ca4nn
JJRzRI7NT74hWGcN/6wxEIgwEvzAxCr4hf+vDRZv0E4lRmpIn5hMbkVzgQMzZ2F+
27ZPbgytDnUovn1Es51tqK5zMEKyNh33SWGI6HO7gbedvzgwZ/qwfOz9SCPAKLvn
qzOfBd15SF8ltux0ss0RYWm11V0WDMg2giOOdH8TmtlHmYSJ1pqWA5Znqo1lqxz+
32d0iZFfOTSsEzmTUVzI5ryx1clxEesvnvKoHBkEGOoTg6fYxDIgnfitAlrT/b9Y
meweOsdjTdkZ6yb9JOnwk22VGePXhDb4b3BtBEYIfFdYcY0DSVqtJNSoS+cSKNDx
CeW5OxJzUAFOgd8cFB1RxCfHeb8IaHrozrmxKHZ36oKmXAM51IIBKbAHuQtsxIpb
ERZfznIlG0sBqfHrK3QRpKCG0cym0rtczIBf5/DcAn3RAFyrz3zZsjYj23sxQlGJ
EsyWb2gfOcG0F/PrssySyZN8JVwdRXFKbeIcIdBChlquM4YWDf6eHhVcW7frJ6uq
Ky54Hn7CT3/IdtIxsBrjy8m9N/amukI/wB11s50uF8DwLBWuRVhlM7jD3EMwaDCU
2FZy/BJ3ipwmuXxZ4mc8+epzm+LwyroS91/HfoHoiSf/j1xu1h5SMR3r5euCAoNa
Z1zMnjzJIEzo2+rC9Kczv6S21PBHt6IAoyc9FyH5YGkLjtph8/iQI1E/mtb90tg+
fdR+W4wSF1uRvkAZ5kf4KHPM8EWmFDbMhWZaaytpi7A=
`protect END_PROTECTED
