`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+mWOoATSDuPUzVUq1PNcH5NCSmS0kvx53zq6sUEgdxhzHacU6eIeTeeauhzTSo91
+foX7jE96Lsdd+ORHBOVeFGRt0+UQeS4th6K3pZk7Bp5986gNbPjp8Dnc9h07+YA
x1LELWgv6OksuZ3Mx3hU3M4ZoQS7ukD+5e71qPJ9fL4FKIdCbN3RZNVbn+iQ6kWm
PN57lriG9qAKtQjqDC9fgwISmjvHYwn3mjjb315iEuyegnnemOEGP8f7JMZAmkqy
`protect END_PROTECTED
