`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
duaBTIfDtW3qGD0urrNlhbmvUSgho7bE/Rcx8wUS2gUENAkxSun8iUTMt7/vmoCm
EtNT6FnpphXerK04Wkfn33RKrJ+ZeRKK5s7B2nV4TvJTpwJrETGIAyHZbRVzyeE9
hYJpNEFG9KM8tUL9Z0zVBkfaWETzJOazKobm35kDomUF3weJQ5/uQQ7SEGxUmsif
k08wtM3G0l4m5nVY5Vo8irLqzOYAvzHAjk1dWGNp1mSAbAshZQEYimuYuYnmb6bF
8UM5bzmaI168RkvpHjv5jZXKREmIe9e48fYW8yvgbn7/41HLQrSvZiagtFDMzoIV
zxXcSw2b+kiFTRdD7K1Got+TIRBJ5BhWHjEV+L3JQz5UlTOT1ng93TftrPtqvN80
sxsdXJshWvV+dJMUrD1z2RnUf8c1NLXafI+gefwfUfLfvi9IzTqeD1hAz+aLLpYY
UdkfoxAXT0u2wVj3SLYuYLTBsk9B+O0Rj8NfG5cdWFT9AVMCiPVK8tJEFt+IvWzw
X4KMXl3+bUThWOhCT27rmx+XTy0+J2h08fZWhtezq5XdGwgRbwUpYhcc9Rv6n7eG
do3hAAmXeTzqaK6g5PkQVV4gOX3b4Xuqd7bSzxA4wrmoV9Ugx0RS0wlHq9yh/xuc
dJP050bFFY+i2irBrtxydUFNKFrp8cDxFAXREuN0hDx6rpZhI2P7EBu97tUUNHFF
4LNkQALyDzKo2c6dBiLlYR8jxUwjz2EHxR2wMAjtdNsw0B5kBLnr2colcMWxRTmD
1tj3vZvk98YlvE1hYMGwnuqxHe/x0J6MYy3e92NMeRlNrbq7WlzDj+L5Zi6E22lP
S86ZofB1U0toEpOPIUmp9q8+UudKlsOom/YG3FTOjj2dziOmKQme/06mBxeFDSQL
xh4X3u2Wqitr/KVZvQgbaxU4Wg/7bSxVBR7KRr+TyFj3ppZBqBnX1GuN7UFwWKea
gfET2aF8r95bJA7xWQbkUnhSEJK4rX3/T0RNP1utlG5xP9QdtUdjuy8WUkDKMuHn
kfpNz2s6PFRYl0ZeWMnJ2LnK0jLYXFxjNvz9evQxrU8q6CbbqhwcA7C3CWNRn+7Q
`protect END_PROTECTED
