`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uejggcTuyfs+FXLouDwMyI9EZyAt6WuGlQt9s8BqQG+oZv/6xiVf9qqGTKbwLfqT
C9ZlJSnpPoqhP++1kqDxdLCw96optLZLIiCckgbOdVim6KPQNEERc/ptskD31JOt
5NIHpbVgCs3GvCPemFXJozv+8p5AQB8OWS3leMqVFmW2f9+WzanRc6L93le7dYxt
MWeisHYgqul77j7xONdBh4FQEk/eJ3uRbDvJ6Fv3OHagmtDlZSRd7eCUjcxt2S+R
Yfg4f1sErz9hehGEfAqwDmIlOhVgtGFSbbt9KZ94QeU=
`protect END_PROTECTED
