`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oXkoD7ZFExzPNv+PQSNQBTKJ1ugzqc1WYCdKndHtmSs9iA3vixq+ZrEkTDfZwfzq
GWBeffSowX+6Se9/1T529soKZIcRVgYddSMKW8AOyARChtxWUXnjZJXeYZHjiOXY
SmThjwq8e7lCrPAbmmcd6eo5PhReYhBGz40yIN4PeHRLrYtquXRA5aqdiqnJdnvY
bLuhRNBpni1gDuqTRZiRbPSac8Ku7thuhfHBAG6jVswPO14A/9oigei+2z9wh49X
EQKbxIL77lpWgpdYAJg60yIjT0wLTrJ76JGjSzDnRS9/bSet1g2LidpVvrhQS33E
cE6ezoHNr/crkmLnnu6Ogu9/nqdGUzEOuAPtthGkQyXlwpeDqjFzlwBuc3U6sW14
yz4HxrAjf/S9bMlMkV74dXWUKTACXj5XaM8LgJYGQSAUd0YAkTAiDjPXrTK5duit
+/wCwRFqErLjlGgmM4b46Tf1WjuJZCbyCgNacbS9epw=
`protect END_PROTECTED
