`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NarEhiAiaNzaeki/qye9K0pnUQBtaYQ9N4lQfbrvNfxHUlsz2HG0srRGMI3CqXjW
o8MS86L2NtGcF5rwYXJ6LHdvbwe8h778fDJT8T2tpHGH78O3LWMkdlOgiMQHBGxc
xrz0i3n3YZb/UCNeJeMr7DW2wsz8XBkq6EigiMAzf85F3X0vn6NUVxrG1Q9R9DNV
1Moke2ON+uys3QTmOYeedB0vyjrjuohTJX6tApKcFie6rdHaccFWK3z9qw3Uh/+Z
h7t+UDrU90AMTgTnw/92Jd/CF+A4Rpxtgrf5tdJGypxPSCib/FhgNdOVLGdKeRDN
kLrNqEAk7kAVsIirce9LBt8HPEaZSkmk4xBxoqR9dW/1tTHkb7wFTroxx9JzTMlw
SzAbOORc1olqka099SyWmqu6BT5yaoHykf520Pb1ggzwL/+LRYLHHq4V7tnqH/rS
LoNtB3CNeGjs9V5EDGZ7yJ0XbLaGcNwD+Os9p8yrUfPtWNo81FaSUIqY3TD2hd61
WlPNfLrAKNtEQxGWMvN4SIUqYooYstGXGXnEZH1FtqZt1x45zbi9iaDA7skNSHzg
XlYCIDeyh7LvO6+ptnecUq9ooHbbw5XcijcotTzMtHXDQJjKZoyLpA4fIiStho6u
ejxyJVCLassQLXC97SoAmWCs/Oh+tmayaOq875Se3XRtb/49wS7ijW5BYSpghuLq
GPHcxxjvLJs0qXKv6BFmN1KKl4qdB1XyBKqPHIhqOt96L8XNQ/HLEXNbZr0sLxna
xnoT6oXLt8r9bIPBYhIiiqSAXLFmzjgIwmVEovY31xQQyqevqXShnRu0/+/YFHlP
IbjPtAb11GQnI+huSjRjKs1mKHL5bL0ajKo42ekNi22FoYHq1Yc1rcwW12m0lyB7
s0R+7BinrulJ2HVs8gO2fxyNqkqCq193ODWBKTtX0y42o/7lAGkgEdGKl0nYjhaa
Z+4XwTFTDr+GOhMUBtFAnXf6xvAHc/6gBb+kcMqPj2EOYRNXBezAZY8HckhXGm4U
XgDGEo9KOF5l7EWRmWTVDSl/C4aISgOkGm57vk0eDbp+zhbm/Rct+bWoSpcFuYyO
6g5p0bJSRRoMGfmP0BpNipOwpEhutt9z8VkDX5rBH3WzD22rPHx1pBIgFQKQy88T
xBmmTOa/tuqC+AcOgZnpb23Pd1boDXoAiu0c1c4RlOabmkqRAFqRLw4Tt+wFUWx9
I8l7tgsnmTJbNVg215K7aB8zAggTcFIAFjJd3HiaQySyKiTdZ8jOgtulvc6dljyL
YxfyVd9jjpElovs4yXBPmA==
`protect END_PROTECTED
