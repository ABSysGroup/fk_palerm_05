`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3vMVrp6nlV1uvIWhTNaP5f2uo0+ylWTRapUjUYvRleiExqBDRq3WdxyEVM/ueASz
LA/1c9lWNeDKlLAu0SgFKPgKZQPhFZt30d5qIxNZMOxYEcxtSpNRRL7Hrh/TCevZ
l+NevTEzOIPQB5WoL4UjMy3fxUFlsy02f0NR/v8x5J4QfXCduXuRCD//JRyCLpHq
nbymIOk5xpcE283/g/oZ04m6f8z97s9qm2IXidgir7tvx3OYnV1ElUQVDK5juNPZ
+3BobZbGoSomXCbXVh9dzJfVhZNx1cwxtmWBA4OWDw2TzlWhZNCyKaGObDfaDcaV
p/hIXunT2bTECEosCwZe+WzBeN/+nutt2zCV2wMJrUtXZCmS9/r1CU6Hak4bBS4i
wpG140KYyFqiwSaB+LhaLRWlDOZsyLbQ1QvAXwkwD3cw4wvrnsEx2QbgPJZrvT0g
p38V59EQkWn7WA2bpt0/o90YjqrLMQ8MUs3OpqyTbaEe1uEPp6LnSJBLSRm5fI3f
8EvzB0wQbD3jVnlWhUroqVZtW1u1SnOLrEYgZrUA9oE=
`protect END_PROTECTED
