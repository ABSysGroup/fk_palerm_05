`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dr/NbE3lDZqfyKoLjKMfVKa7XjP5Gvik3Q6DJW7GbubLNSjZ3MVDkWy++f3m6dCJ
xG2G1xJDOZMoKE2dd36SAhxOjTP2o0k3BF1OWpunEX9GIYE25ulB0TPEM8QIChCn
Zth+mEmymfomDyE3xEnZzP38r/6XhTFGg8/Zx0UucFJ2LYx0/oK0nxPrNZVF4LSj
Bf6OTGoy9aCweReKeIxRmKaalIoEQoLLs0Uz9gyOooTxIRU9zWcrtnm/fw/RUhGt
83QnvcPTmnDzpmeP0fM4tA8xWV8f1RGaJwLiMaVmRo/Xa2CmMuvtdKh/nXqyf9jO
yyA92AU7mQgbptzDuJZw3+fueKYn8QkDKkOHHv1wjGg=
`protect END_PROTECTED
