`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wvhxP62jlyLcZCxjT0+aB5Suf8/BkawnZrm+7n0Fg4kLH3FgURHlv7TTkLyRTy6g
S/85LJ5hwHzp63kqXuteeGaJRrryjOe+/8YzKdFPpjbGyXaMeJEz8eV5J/21atJe
mTIvvvOQlcBJfUbuTS4s18oYs+MqQQZLtypitfgLcbiGimSXFoPMpD0JH7h5vOXc
kNvjUbU6GsxxFaefuSRTh5tm2iH4+9Q+jq5LKf/cu+weIPu0gJdSHd/X/udBhMU7
0QWUeKUpVEExgbOqLyFS6+LvrwsZ0yWXCbd7M5qD3PMnciuMjoqelX/TKprWoUBe
cKPWXDFkw8jNLPbKtgnmL5QwPliRRiCPhMMokPt6oXaYv4X/O2hlN407isDd1vn6
Ugixo9JD+pY9QPHxzZ0HTW5rqdUOo7o5OCDh30HOn2R2br+LEC0Mwvol3FaXwXCq
nQWcWJ4br6/R6lqQZWquVg==
`protect END_PROTECTED
