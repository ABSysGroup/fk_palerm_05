`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HAsfHwR6IbHyiwq13i0qOWXrS/2aP03JWQRUv4Fs3xn2ObhMOUSflU6NnfFF1epE
WiyFTzzZ6On9pZeSy4wms6J2Q5rGYPwmiHn1tUctpIi5Lb3stjhUG8w89wNN56DR
FzXgosc7HyWFW7SWeH705v7U4jJlHAvmIqqnPVQ6v0ZOraWYIpirLBpmoBp7Ygvy
+iDmKz17+yQa5bM/AApDrPZA+0JxPvYNQCL/rmMFGjDuTQXxj5/F7dLg86AKXHVN
y1I09Cw3B87HTxBKE5i9o/On34C8fcM7tFSp4xIXXVKAD+XqYPWr1xqluClOvK2K
8RCxWu1SUsLlCsyfPc0CqQTl/eXsn8/x48nfvorSL5GEQ17g5qZNauyHKHAC1iWn
FvAwDvO31HheifV6uMUUPidVxF8mZmX2wFCrFUNWWBctP607QMJVg9YwlbinIW/w
WegugEiAQOJ9J4lhOi56PUU3e42E0wM9e9PJDkzy9fqggoyz5qZ2EEkAY5s5TF5J
ah7lsadduyRtTQ7fasw5fTs4T6LVIFh7wbl7bYSliOVA2t/klwf0LbA0jeDn8QRF
/vrl5z5SCNdIKuAInj1x/eEpjPEhbP2y3wk4aBPuoYzjYMAVWIl0UmEUhdlWBwqu
QFcgo/OKFlVy+8TAVZehAA==
`protect END_PROTECTED
