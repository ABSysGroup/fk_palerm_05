`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HeFdZhAygmu7qxaDu+xY0rWoelYKOHY3ZNVY3iL6agwjRer3DdrEEUQRCrL3X2eO
Zi/KIgrG7Hr6X69tkgiw7z+xR9MrlXc2biK2kLCgqnEb5lCniqc48PBss2X7fDAO
V878uDBG6LdoU8Iro8jlbXwGv8yIXpyAHGV3fogJnmk9FPdqO0FihrFgzVuuldjS
hG6ZZe41+AlcDPwV7590IHCeaxQS+GkUUSbnVlr3b6gDK4tNpFbNAZJZGwWW0aK1
Gd/+IccnNAv1B2ZbHYAbuwxFW6KyJvtkINm5jn18u3RpSy11C4o5DpiEc0R0K7mm
/vvFBBSKXpKJ/XbRb1SOIItp7TAuZdnHlBm9WaSVESYZJbjJiZchCUw7cDdbwi/r
D+p4CiKWLzXooUE0sj4w6lHFvAqfO+Ybp9Hc/QiQQpa1M4dVwmg8WYNk4JqnVouq
i7gkxTYZmEP1gcUHi4QKiHMZw6eH6jvHiC1H8fP5RiUTXTG17/k/2V/rjrplbMS4
V9RJy8eaMYRwfu8R6+QytKMWinNt6HgPk2HhUoXRVayrtmkcM1hDcdQQ0/BKThgU
UBKpCDapbHO43gjDuwtglVmwOvO5sph2jqiyu0NLmUV5GmdtSGtIw60aV82bTwIs
EoqNreGCmfFtMshS5wiRdTHPrMEAtEjY1zUgvGGAZnr6KOTmYEJABdmeDevK7/Xf
kh1Dm9rtv205Ih5+sJz0BGpS8dKsyPlaeANFxUptwo6FicAmBKoHknThA9Bv6QlM
gnbN02AKXHWI4lC9DyR88tBi4bXCA13ibXrbhZ2f91glGu57s6yICj0GOJfejZgY
jRJblvu9mwKh9AXoJjKLlr+YOXZa1pRlXYiDTqxp62npw/hJU6EsN89eFQZ9URoU
K3eDY0N62jA+SGDBsXCgTTRa9wC1rip9ZEEJJkIgZweUviurMNJ9qYAGsRW7Lh37
Y/dTxsldOV5gDDEE7H/Iu+pv44sq9JLHOmQVjenWPpSmE5uX1Wv5WFgKRKuH6RdB
NNCIX8KEoz+cxkwvdOFkIryOVn73bdLFjhfTPFfWnDRus/HBfDZJVTKsJAkjw0Ub
/I/Jer27k/bdz0QNSwTvyJNtdK7jLOFInM/z0pwUY+tsN3ZgV4KdhbSAlw6Yd/3V
HTNeo3B7UOe5H4jZgFn6stthpfofrevvQyEvoAOhaD4Y7Wyd+NQTZLgnNHlu9PlS
vjTXRD7ExtqeZafH6kWARw1kLX/dpwX/yiJVFz7/YJOlip+x64RPvht/8knhzkgz
jyo2zz8QLAKz5huWv7ppHx/myhSohAtE0JsCpJ2oBclEpR2FTuRQUv2R5PqCkqBH
NfsEdy1Nf80ntw9s3EVq30lu1qfuG/L1aO9I2SmxjXp2OCrtVQoCdRVETSIPQ/Tm
wpr39p5fiwqLY3K3rCIuBcJTbYbfLGW1TM7AhBPqU+Mpz/nDik798fHqE2lUS8co
I7+G0Ee/ow9FxQ/vX5H1En/rvKhaRyuVMrK8J7zebGk5KEQWLPCBulM62aNi4COJ
nox5OU5SIOdo6hVqjNo9Bf8Ha8sQDrUkwAD+AlySq1ejaekZAthalF5cR6X93g0a
Lr+FuZxv7j8g+ABPVcmUc3ujmh6/Hc5PevoNQqHN746n6fv2FsFROyvw3sw0Wnnb
uC7PV29uTKjFuaXUxyNvHQ==
`protect END_PROTECTED
