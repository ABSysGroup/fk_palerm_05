`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zbKP588IWwnhsug4b3p8R5eFQJCJIYRF/wGj5MBei1a1ip5u8S1yvuz3m6WlHQ3I
rnVd3A6BqbYPuQYGtUDLKwNc4eH9wPp2UO8quaa/uyD8jR3hY4xuvjB6fF/QgDod
CQ6h0pBvVO+8mka1IVvgmEPmOG1n88/jO0G+hohVoAAYDLVOdbZdJIT6WKLtNBNm
tBetHhFi4mi9z/fDt7SYy+y2BUw+JR+rmy+v5vneVfvjU8xzuXaOSUAM1j6qeQNp
zrdd/l1Oi3ivn1sg5zUecf1l17DkvR33peMdppnGLDFd23SO8g7elj4fPVK6xkaJ
0TZYt/3fpqKimjJ3R1+YQeXMSssyGoWombk9fY18wsISaMUAFkqNyO7g5CAqg+kp
+H+BxAr4GkgROM2UceNf+AGUM+0vbI+j1oNBAK26gEWXwiiRgECkvkWCkueLGPE4
0Wu3Tz2y2EFf24Fbs7wx0UvCwO88K8EthLOv5iEqNZiV9eNOlmPg3Hmux2TyqRue
br2DU1Y9eLZPrjmOLVy37JEssynv5TnxmERHTXFWqOMyLPeGdTNeUJ0evA5GLflI
aCW8Q2iPx/flx1vbC4jg5QID5cVyXrnw+Q0l3v6lbz89cAtLJwSIhHaIuI1CboT2
trg5oKESp0YC1SiEQLG/TQgV5AbcrWgYIveFkLlEvNimZWJwoEWVOZjkVT+aw6sR
8lRTNmJbACKMm9ynPw9YycKmReQ5qEO03AOHkoAS0o7M0szjUVkaJxjVZmJx/PnE
7YWda/pF87isAMr3VvABEkT8aP/tqJ2KQ4A/OjQ1caEUM9XDmYrR6HHOQl7Ndksh
Notqygh45Y7/a76h9ZypwxQKgTSva4I6JYFPSqXXUch3H2L9ftYx4D5igoI6BbiF
EcvHnbgnHQYR15VNd6wnAK7xz8BYjg3lYgHhPRCM2IhtqKAsHprdH3bxXxemm32c
2X+gKKSM9YbtKO4k6B0O0SWil5t2WuGqtvpEe1loq0U462q68jqmfIyW8bKWBnWu
o2Azvg+unr/8cdFhl8+fcxiClmolxl6V9pcNHI5AMg57nfDzw8ZyUnkgb6DuDpPx
VZ+MFz2AUPnE3os9Q4Bj22RPd+XFrecziwmEKOZbRKoS3GjlP9HTkvVtMoextxbW
+3QUF/aTE4wvXx/jxmu5hEqTks2IqRLK19ybmLcSdhKV3XKPzbILaoUpm8ZqmpEC
pctZC0GtlKV0eeYfIHhAZhK863TYp4e0mh8fJRZMzLbvku3bt81EHM7lxARAup2i
Kb5pv2tS7/jTCcMqJyypmtFC7SSFXkFf9bqj1IRKSwgDkcWPdpjVlc8/ACbF5BN8
pdUckwdA6Cz2tfPv+mSgHLeC1k161mH2EX/Q4PRCKdKF4jZQyEJ7wcTLQH3LyOX9
B6KQkcQXlkSH5hZ9RKcDj3UMWfAjnWXJP50kdLhE0vwmW/m3G0g+wKhrimUDP4IQ
HLmIWe41u3irfihQ4sB8/V2DKtWwSv65j7L1rhC/FyQUbTh/ZzupJRi3Mnt+fi1d
/GfQAlKy2AMVUGezikNgb8W2pTpBEyECrxKTPaV8YRAlIgnfwzopQTJ52eOjZMMV
2QK4TED2KWkiLQ/kG5LgVppq1j0ByjKVsSCoYghwJMrGHnTYZ0Vx93ca+5ec03GS
TrkPpOa6S/MzEpAKgPS8j73KRDBD4VnxXqiDGH+bRZuMMvnqmA4HtuZfebG8NFtH
KMbJIXrTS4wkVjfLR6u2neBCF5mumIPWq7HKUwRSTt1wt7sFgRK1gTp/2uWUYHgE
0LXVaFDBroqzUTNOf7c6Hy+pJkHxXhX1Ma5HbrTYwkFMzoCi3QPNnKDeB9rWno56
mS1EjXLer5u5mda3HuKM9R72BzH1ZO1Nm3HQiWYu9Q43C/ug+BKrSW6ocIAQWkmg
ZoA9zY/HhdLOj2sHXCf9/+CNPRWE0KKj+IPMUjYFGWcZnxflWD3QgeX9BP3GEbVg
XM+JA9wNcgTktD3FI28lJrnmKJvHdG/EuAUVyoAaXcZo1cPKSwwKT2SHpXi/kcSP
R723dyty1sbh+5O0ifsr61kDNeWcw4qEa9H3BW0koiimyJQryB7H5jZbA8UOCVsQ
/c1Clz7xCcbfCb9Ckbtgowc/5Eo1QvMWkbOt0YF5pSplvRNtQNBCHuZKpPdwPved
Za+8B89uFu2glUv9NLSHCP9muj8Bk+D/fZ3GsJGfdyF/FHcevViKOs5fbAb6P2mf
u5iGQBvUMHwLmdzY2oQhXCeZX45o2PA4SmsmEiZYKDCe3ZESyl0VxEmAGlPRfLZ6
GZfXh6Pu6Vuju2vcv1cjWoYaFU+yLrWq5SR7MJ9iPNwAY2uefni2Mi61if7FnPqI
E/DttzNDhH2D/mYyl/CJV10DbR+27kLUUaA5Yh4w7cQelElTOsF/PANF610fhsmw
xqC3AYbmBat6/dARjEW39ihLRfZn7GswwceIqeBE2+c=
`protect END_PROTECTED
