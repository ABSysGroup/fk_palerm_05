`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9zqCWST1SjazmdUDOeUkMbgyKtjMB2ZTdEVYJtaUGR7JznMgzKb/TslH0yCv5KwK
fX8F2GUntp6EPyvuvba3ADytL9LxU+NiZ+RN1zhyzCFhIuVTz6++wth5X01JAgNM
KF7wxe0i5orhLRg/xOV1dkyBm+N/VdZzblIO7pMNfXl/jzpwWKTX5V7fBcVGx1ny
2htPWuyZjYHP8BmXkitVN1EAwkYGctHAn5A9X7fKxRF1965+qlRwPwxPO+tnVVUQ
m08b95qZ379JRk96Bl/jXclMzidif7bezKMo8bVYc1RSOH7f0/5CaFhpeVZbnT2g
qYWxCQQCEyUtwdtZr6sCnGk93kun8dgx357rDpTeOOnmdi4FnRB4UjWzIedH+Pce
X8Nz0D7jYLkvqK5GdAAuGd1elG4dozo/5gsQeqqDuESTYBO5ZdH+WYGX/cnWSuHN
nIJh6VcQ0EDJ7ORVwNVq0Xzg65y4KObEUcinavu9aBUT6St1iKEuheZXRLl8e82F
1YRyo44ImRlDdBay8kl8ro1tc8Molw+ayQiq4FhVJv4Ja99umbRQfryUzi0tjjba
b1H4ilvILApL5Q35cWRBgAl+vLgwvD5fTYY4DFPM9xE0nZe3jC38eV/niK9VyC/W
hJjJhTtEY1HRLrhuN/QTeD0VXCQuKZNSBjRXqWXthOGZ05oc+9bcCvH/8AfX2II1
gTdFnXiP5Y50eON9quEhREBL0GWDVtjHdP6t1l8weEuv9W9Pe9xCpPNym6xRy6RI
rnaQC1ocTDUkEthVcInXRwnb68zusOiJHZHzFoPhcXBA2MYOQqzCv+vY7YRPTbiR
146Tc2k5muhO4LU0bZuRU3QE5wqmFwYIvy3oRcuMwYlrKIzy3Ipm+uxh6mj1L+jj
Q/pHkqOBbwVVm+iiRY1zQsQuUoWUTf88ZPYR1j1tbMcKMQpic033TpdLzGeVcMuP
KJjrCuEPjW3BuRNufn7XQg==
`protect END_PROTECTED
