`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2hQAKQHMiT3B6pMF5RwJNp6E0QxaQrBqgWElHKlkxVihpxieA9yYS4RnvR4Ha65H
9d14WMynLQjlc7wbc5n7MNJgWwfFWcGERWCvhOkzqXzIucW348ck8lG0nvsV7qjB
FRi7d7raArFlQX6XBiigDtTA/ZlMKsZffznQH8eVQRu6QOFKKWvsnDUY8Z1yCapg
7TFk27f9HNphLhBAh4U9wANJ8JTaHKzwDDX/PGgF7mQR3zhoPqLCml/wiOqoz4Yb
Y5XAMJFvfQJnOXKXDtTPwIqSvLSdVzhVTqMtqAEtGYhEGozXvMHFA8gdjZqF5Oed
TC4Q73MGLI/FzsgJv7utCf79uAACFC6cPHFExpDMvRnvgRdesRVszqB9EwJDWshA
+IJH7zWvRq3uGys5kVK/g3m7+cpo0Zn4G2T9JKxDdP6bJqt9R7GF2vzaoiiIhiQ0
sbGRLJrPqfygH4rOWBKhVUuBMcgwoHMqsL/JYyt84h1dP5fXhYJ/e6R2wrgqI6UL
Wpv8MnexZiNqgpnUPaZ1y1Z4Ni/Y9nw7FY9j/e73odDAOxKZVXarmxNtE8Sf1s5i
kO5mT1hCsMF7QeIhbP+OIRv6Ix3R/k/MsIN0GrkbkEj94szY+bmS5DCV2w9O+LJ6
aw/MZBDi/0aQci7cUBC6c9A74QM5MQ17wTGEBDwPss2MrOUcMOVYlojq4z5p+G5A
or51j4ZBp45YEoTb+YzjeTg9j7wHGeeDPNtOsy98KVDzZWpT9MssIrvuMfaRDhin
6vohC1jcLAncLcyoR3+fbcfXm4RMP5VBIUhHi+RdQYpMiTNfN2wrVyFix8LP5gKJ
7fnHjY0nEHHmgMQpqPB5NDZlR5VAINpHblKSO+lYV125f1Vgp+tyyrpPhNayB6JN
yZ3nw0rvUIMmKrcsU30rCDKS4bUuFLkneD0RZqYdPnmfofpbgXCVA30+ATJYk2Hp
5Ig2yDiCYMSoBAY5uuSpcTU0Zw5J/rxNLS1+fSHPokaFE/HCZ7Dw+q8lIPajMR8u
J1Ck9cZfS6ZKScU0eiIz4qx4ozPdY4OIzKcGAkaqqY0Jo43vmriuMiYS/YdiB8l/
EHw4CcMgaGXPy7iTWBiIpvsr+ZJq7h+mtPAiV7n1KatOvG1GpLGwJ8xAs6ruR/b4
+WAxUrJPpdq4oKeOrHzTZWRQJ9tLGfLIRAlZv4Xi5qiZoRuZz1iC7m9j58NSOf2l
oMNkPvdzPwTKqgybMxl6PezbpTjdxHGM0oDFUw2TZmaNBsW5aQzTihRW/1UeAhuW
zkdmxXQ1uIFHkB2OtQfUKDcImDkHju0L2u4hNcrSXCsSA+7oo6T46j91U3gVef2S
eJGC29ROcsm8vYZKtRFMqC2HJMime7oCqBjA467H406+duAkyAlH5AEngR3Ip27B
26IjTZYFMY/yQVKmJjZfeTtXLiSQpTLIW178w2l3N7nl/rLJqzEiVylLs0CpN1Cs
EPqgY10VSAZU86+qgvmHPGIE83v+3K+pXrx3l4dcFfrMCJWBOcHsFb6YvGtU8w5J
UqXrm7Vn9HGkm0Gl9i0ic2RHI6IQ2Q3ANKmmEfAGaShE6UBlmKTLx2Xk2w32rMdB
J52IMQwUmTkj62f6EgqDy0J5RRkNG9abDxKuHi5buBNJkeAtbOlFdUNBM3dZKZMH
L+X04OvfBV3mM2srefVNwMal0d7M0Q+Ah2I25//AGVZ1szWdfYiuRdSEXLZ5lSX3
6Ps11p51IKP1q3sd2C2wZX+TlTJuAEKTysHHwzaLc5PCf3ENlwpmsrUtisWm9P5D
q2VwYuHgBQMOER0SEy68ZgdnSFZsnkAXC5AtnpYGIsVCcU2TYXxaJsUOSnCIgWER
K3wgm8nl0Lq8jfY7T3SPWmWxunRygTSy+LZkdNHtZ++42yn6hooVJkyjTlztz/Cy
ljweXvm0mQNJ6vHx/QO71AsuwItSQBAzFI8v6MpeTIpwzNfPWDJrhvHMtqW+BRQT
n4DCgm6m0DY2DKEza2RPGLf0q0hDee8Fkr8Uw2M8DX8bMplIeZj9R3BKz+0O3/dZ
K7zwu+9z3Ddk0pMgcL7f3gdzNVVPkgAm00xxRy4TzjqAgo4aoTSo7+HOHKNdKPL1
dNkCG4OXE1+WLc/lbZ28uoFVykzkX3Hi1hyHJT6xyX5o/PCkciIaxIKSxbI7BN23
5xmYhZdghA+erdTlVFbNOC1bFZaJ1AQoWQiyfunvYQl8e6D7e5cV1hAJsTbkCo0W
MmA19f9Mv+v7QfXtn1HuzpaNdsU06E7Xpc/lIEed3ktRx8eVz03DoWhvKIcBUi+1
5AucKS6uPWxRY37BDzX87FZrflVx7g2YdOmWrxucpGPZbR/HGWHRtOZ0KTEj/wL/
Tb8MDUt+9Oj8mNTLUb93eGIwBZw/H2E7F1WsUTR+ujiDhgAr6FD2TBvwz1ebg/dZ
8P1wYLBoY/c1byOW0lSPDaqKaBkRn1YMMUnSRBguiMBCYeaLyAoS752boAQgQKj2
OYe382u9Z9YS6C/G9JNo4csKTPW/OnQJB7R4ly1x+ZasmDajL1pc7S1e+7nalFUS
PMU2C0jQQped8BfczhTnUJqBHyz6yjlTsI5jSmOcE62dW8AW0wVm1XigVuV6pSem
tRFp9u78G/S1jg9WpmIbsQ43NSYEVS9pYL/i0jV6f8kzf9Pb4mFv/1ScZgfyuTGg
mMZRvewnxLsdGHutXESS2sUn0PLjSlNCm9kSVJxiJzbq+UeLthpy/rZAAGRhGixb
wPABTfoopIzQ4d9dvAvgwfczKLkd4OI7CLCfErldY/OqyopO9WpdSEccyJgtthyC
ZxT+0EOCGBMV25lFIEvfAKEn6CmKM6Wv8LDCKqCAM/yKMIXTn85opAfd/aQZENCH
uGZpVZFJUvf6e/UbrKWBjiDktmZ11WpWcQUOFYUiZcNS9vOgRV3FQwHZcUOcHrEA
JE1m4rDnoRK6WdM3mSlXpbKdq1MntFnEOLehyn1sQa3tz/dK5posEu2yAHvs8R6d
P0zOMYW7ygrjfS5MXFYqwvMnK6W0hKItI4IIXPfN1nVaWbPFxsQ8FXtdWDhBFQJ7
b6PfpHVXtLxCPTVBRDCxnh2FYM+4XZ+Cz61OPCmZV56DZ5EwUhilQMdlcJCUnzVu
L3uQ0v8Qcg+WRaFV37u9oNCK4bc1Bx0DAbMKdk22cr5A9pUlUyoaHYMKJmoQrLo/
uWIFlAZ8bCKr02wVcKil+F1oYwvDsDNxR0PEhUJJ6F8z6PiduMXUZJ7ycmGtoPim
lS4Tk5j1tMOP3vwt5rwqW07xSNpKRT16RWjFmuHQAmn3MBYxmpxD8fn05sMaJxS2
QLjtvZXCDWRwNpvwQQjLATtldqlTmI2vwf0XeAjzDkFJUS/GrtSoGIpoYdzzKCRr
8lEAdz23LXObBaxU9xbciwUtNWJwfhUWp86ddt2pQuZHeLrizT/8PBqjjL05NLEW
WPyFxLGCZh6vzO7MURsg0brChS0StmRwTaSGvbkCXD1+5rnkckE96Bhs2alieUDo
U5/LSYYA8XqbbW7V725kx7c0rcxLbqq/NsHkDWmZxGpxmuIv6w8c09GSgxQ6nS3v
e1kkdRnuqkjWhTULM8lGrnerJLpQ3KDeN8GBzAZwkx6l8AYsGO/1BbVrsdJ0OcP5
+VoLD1Zj1wDPYzvoxDfUTHigPfWuSe/BHtVv6tSrWOAo0zNe3ZuPh7/diQmEvIDl
OMUUUm6DwZYwtcYx65iQE08Ez0r5ULS2+8ughrd3UE+Cq+xENnk0vXcccRqWWEM1
OHUygm1cukRSMgduBvcZ1D/g63Cmx+06s3wUMUP9c0gyMTzmaFxei5l8qZdqJs3X
0zKzGdpPXwj4uSyNGLCmU4L9yLQCYkKSuTaTElLd0W85yCkJWGWfIHJXMvEVcIFL
0St/HuaMiRyOkvuC8dst8FQAcEyULv0Zym7zLo8P3DnSEZCaNAP/NWNXoJhsIzxw
wgVVaUaLhfTDIdgN/AXj9XiYxzt+emPYyudJAV+8vrugm+1HETjllX+eqAYpyANb
BrZIYfVcDmKRjziBU8bpTwWZBlJRUC2xGNClfBfEYG/0Wmn04fajpD8js++hFjbF
vgftVKuaFSVQjzKpXGq0JMFQ9qeczL2z1WYE/ykgondbZNb9G4LyEcXiZpu1er4V
kRpRq9pkiGo/7oorJQ192TBiHRLmxxdcejtEFDmNWLt5Yg2NCTO7gWEREJONe7o5
zfQ91TmQdmOFuLcjU3a0iCx3X+k16PthYRfaM+76NW19mpc7WwILmK5X8NSwNtkN
at4rZIJtGHKL9lYYVxc7D3WCmIrPqpsmeaYJkm0OOc9ouXDgzps9fy2sHwVdSzS2
g8GnYHhz8yOEo7uZqM0l+fWcIkcIcX1l9+DNhcIsVKfyfeZHJu3c9GRCZla60Ha8
f+Ni/cLQ9k6brhdTUFSML4sEB7GnRPcbUc6CGk8XTGhBQ1k8GNBWQCUYAYjAIo7b
sJBuCOJMsrQVTQwnM4JiZUboAweEWbkQ5iIdBhNC3qy9ecIsYH9fVEu2OqYvzJLy
8wUdZSS5pZbyXyJB+1+GL8Hzxdrd+qYkrL5eXmXG5VfKWEsym78kvxVGZzoXdpDa
5JRfPtYzKF1LPWoxadUMw5kJ25Wo+242Th92W17WlyXuV0a/u798r6O6zM7is2EB
6V7xC6JQiwRUkMxJnmIp3X6WSGr0XnAMVKCvfmjY8KgNt3LGeGWMqLS/47gYrbd1
RAud0Auz+oA5CTid4dxPJ3czMgtNqxgZmdJjvdwb9gsqJrkq0mLj1hPdIcf+yR7x
Y3VAKStF/Zqmda9Oy+x6iud8cxC4tKllcZquVWE7fCRQ4kuNStiINpXDTUmpwK84
gqxC4W/V8/NoXJxqH1wbkS9tuHnPcDZfanAvimMCclWDmIEYvFw2mD/EPIRHkuXX
H6RnyB4NbVEORqJzdXfMWe5HE4IepvB0BUUXT9LsuJ6f5/6NFLqwiSfLl4y2VzVG
iRNAdY2o5aUrKee2k14dn3NAVUcWm2NcpJvjJpk+AiRWo3U0J0banZ7q9GrcocNS
0d311f/Gg4K4g3MPuKNPJK3zMIfEAYlA/I1ZIbnmG0A9o4QghEp8QiJrEB+Ax1Hh
qNdeTG2nbNTxkg8VjLjQYCw2mvG8jBEG6zmCDvXPMPDqEXJsmD2PspOOMcOa8g3A
Ewjk5dr4mbWqPZMRw4Gr7rc7MtM2wdkZO7hNqDqC2sqYK1kYt0xboawf/YRbb0oA
AerdiOhziFrRLRDOxtGL5r7YA6QnJ8S2wG0zHTponqNhxW6MNHzxXQLmUWhPcarz
+K+5wcH5g+aFNpIpitJYLr8NH7c7m0d6cpRIj6tDVWxuP7qgmhq0MVtM0wooIJ+c
+tcBquha6B5ha+EjvWkeQmgI1lh7pKOtNuyMS9nWwwdAxfIgvy7LSy9jIS0FSWEb
tBX2qMNj96xFBQaStPM8Nty1NRhc/POlS5n/acOZr/4ZIy5nxp2laZ7EXqBmFfVE
y6olb/OZHxg9cEdP0J4KIRDAVpy/1jLCTuxvSK5e22H0mQf5LkvHs2nJphwETEuD
H6dmzv7wSz198W6BirezZaGUvLwrQZ5ZABeFpCm38l/5/wqw0lrluIkl+O2HjyBC
bl2kzHjwsfKb8qBStnULaH8jyGWB0pdVeH6tFLC3bT3HY04IJKaJien+idzkZKGf
tvdBeutjR3NoWkiRHPl+dhHxyHTB6w/9UHprv9i41h9DE3COw2q2qJIFlRXNHCOQ
6iCH4r7F7PzCN08iCvJn4NuqtEJsSFeq5kfDFnlVNB1TYEw1w9eOHRHIKL1dESnR
GCJGdBCgC4qI2RRG6YOiWQ3LyhFoBxUXIWaXeMNiFnBoeBYxSFUekGADQq3wK6rx
WbkDlCrWeR9A4f0Su4T+dUO6DVfpyVTt2dyNpH9bGkVEOUpkrLa/UC1J8FqhwXAL
iu0Wj3eSyAzxb5uu/214BanMrj09nhBFW0ACTGrOkLPgCMuUKEAfngdNdcwEci1J
hx2Q3PiT5qz/bXCMsb7PoKzoC8kaREeMLn2F69KsPKpMPq0AYUDvip4I8wVoJ9os
n3iP4SbL9wzEt3hEJYuGQOlpij9IooI8hWSME+vGRvqSTAUntj5trDowIbc6+gj6
x3vTghZeLD/+yAaDl/9TK9BhzhyGlgLWV2F0oPSHcKohUk8lm9ZokiJUwTVK8m8n
l7JXMNHPOjw++5025znpCZcktn6OixYJ5x9q5JlBg2lhCqD1lnZHYdsKHyrjyeP9
vIOEVqOYM3IECywDSVQwPgVIcQlTb4D+tnZe+rKVABGpA7MXqo7mG03nNwTNVgbw
DQkHufXq0thgQNfN1vdofs4sHYHc5Yf7ZoXjwyawkB3iD7kgoV6a/bF04ly3p4Q/
pm0luXk3zHCaKo0yWrA2fzjm1LQL5gPFX1qsJqmV4+I=
`protect END_PROTECTED
