`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eN2tahnnDrPaVycudLOo64Ws+13c6SjNdpmScUD6RUi9X+lk7oJKJaBh+Iar52WH
1JfS/g83EXGKZJEWAn6iHaG0ZJCq7g5nUx/aj0PH/5xq5UDq4nTYoGg7cqzbTV/G
bv56yUohDJhawFgiBe6oXSRmP0mJUe9okqQyhCIx3k/t9VlxW1FHhoSbRGKD72ES
TILucYWqheclcJrmrG53DtMfjkDboJ29LVgKVSvsi0jomF3ucUi1bBMpAjhPzp/M
22GWubYwoc+RwLd8uv/HMKkKhBklklh5t6OoYpIOaDyIk0MuVahTe7d8E/coCoWe
NzOUqshGFujfi8vkwihjTkGGQ7ues/B/6eQaV/NCjjorZrQdCi8BCRXu6sOtYbRl
KGB4yvgQ2svsaKukW32e51FqHKMhIQyG8n8MTDLzmY1u09LlacEK2xZSp2VK6dR/
s6U5u27Ey0vLzjDwSYGUzqo59Edq+PqQ3IURX0G3Jui7PeVGECqA9RUHa58my3mx
gzGkKAZROXMbYiXqksB5EEfaVCTNsG4YjPikw3HERr5J3a2TovqZSW8bUJpjwqyr
vz25Jwg/5ZQEca6aXQ9RdMbH06Wxg3BvlID9+mDlAiHkVYoAnfo0frTfoNbho1ym
fHK2apmiJSjxNOZ/BYlkgL5hFB6LZSGnzUVSaWRc6DwrXqI3PWs33iMjTPYk5gy+
n6LQdaOxxb73cdciAiH4Vlu7C+60qws7qLryEWNR5M3LaAbBQx+1OW54RKNY4LA1
njybcGm4TVIkQEC/ABtVN44acVvDIWg6+KTRWJUuPr9B0nbkGpy9TvR6MiunSGFY
My3IDOGL7z5gcXeWi+OIEapSmg9uJUJXgXv1MbvX9HiIcxH+0R4b5YCnJdzeYOk4
38C5ENSpfhqp0FLgSZua/Yzi/ekSuFMtyCGboEzLT1rBZclF5+Bry80DB78bQk6b
dLRIQBSH12V9XEGm6oO9Kv1SpxndZAJ+BTsIFpl8RiigGL6YLF76n+jpK3McRrcP
YHFtvacZws2NFU79oJoRgm8fVa8ft9+b7EkgcstKYLuxyBP5etjGxsu2xbLfsSW6
YXYFMEpcrj9mw2B+xvKP53p4lKZ/mE1NZBJAHygr78bmqErknr6qPnvM/buQoB5p
M0jNpCR9MWBXYJCxSI9sJWPb9LHzehupkvKxE4+zEOPXbMMFeaKmnZR1UIvyk7yT
OdFAsNFzRevtyhMwdJNh6d3JLoHyquJg2xyEunatuWVZ6IGGej2q3w8MRnbtdT4i
HtsF0n7f14+s1qSmAwtvMpyHtnSwdmKdDogmOM+uHJS1ftU8hF7A4FfYZn69J4L3
sBQTDh/r+6+b5OQ0sZYmeHY8MiUOVYMY7qkhqDvcI+30Pg/za93RA4mALFhgk1tq
XSNlJv2UlHYcCbaiOHVeGiRZvwY+NQCLEB5ChpZXfkdb0tdQcn+png16/w21mElO
`protect END_PROTECTED
