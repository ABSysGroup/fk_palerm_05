`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xTBZQ1Dtapyg0FtC4ca7RrYleadSmhRzX1lBNsMULS/gyFIB2be5C/URuCGjaKZZ
nhT9VLJF6BWlopoB0E1apae7tSazoqsDn0DWWBmJo+e6WMUoyNDI4Z1umDNilvVK
WiSyKMLqZ3Zpuyd0xVeojtK/LEk7ND/m5TYjDV99hOmSNACF9/wvdlkk881bwyRq
Id7KC1cEPPoAP5dHsjLRMBVh2ICKP3KAaDY4pnvZ6UKDYSok9+8DnatxHm4KkWx3
q1TC7ZN0obqwvVSpORIjZvGTvXGcnI63M3vF0QSVpqqUJCa2n/kONF55n1BrSLVl
okfpM/J38zaaQLVia6qH9+SOUrxtoQE3vWDD/IowXRnXwiy6LeA9arVydnafdZ5G
vMDTazhIDoWXB1+2veFQZdWCDgiEjmTaghuffiwI+LraRQkIjk+vAa16m2g/45+w
2k4r6ExPoS7Se5bQBHeHtyW5pg1RMzKrbMj4PzNEF6CDgSDwUtICywAoA7Y93HeX
mKC2oKGq7pWcdmfK+AEXrdXi5Pnbkw4NowcbgLgCRaVY26zOdNOgOZ5anU/h0Gnl
LBe+ZCPB3smJng4aYYnunkQc/a/ABbhF7FV63ax8Flddz7VC+/x6/L+MnPblS1i6
cUrsI1w3JBBfz+MkhlPVwSqd85NtmphmH5pY+JgKp8BXFMk25VvaxLp40cUTjYqS
i9nzYQ82SpN4vE43bjMqh4ewF3YxvNf8/1Q1LnSYxxs2DOxTcBrtnN+6XAv4/PIK
liAhYgVzvbHBw1+NuvvSdwxCMW3XAaxR5j0Cqt506myMkTRv42xllWhHYDgIs6Lx
6SKGIq0LEps3rivmAkfflrP2fyudt4pNYyVvGse/oZJHk5g6uk2KgDFEU9zYznA+
+Xtq7VZ32kvRJZamXM3HXnn2nUpVMxr5yR/HdMkTqYcmTf4kATSv5UEVyiTUjB+M
ZHtcmQFqFEcITWeUgCSDBA796pc0eaA+mxI6llLVPZDv7UL0dztrSMxQmzSMP9if
yP0qpyc+1cheYc3UQ3samZVFxf59VxQBtwICqMB3FUWYZjQVy1UHXi2+6iuF7tsL
CeZ0Tz7bLtGVGHhyoO8BKeJ01pOCXPMOGiweOj6f9a//NdMikz206SHMZTiqwwbW
jyGz0YjD79vUGFk8Q7uDNd7Ttw3sFjUrQBS7djIMXFMQsjQmgmn1NS5jad8LOL+H
f0DAfZaTJBjCZLitfjpTrUGPmOqzpqY0LrZ/rJwVdh3ynvYcUsodg6WhJ7vUpXxU
n6aSOwxQ/GSjPeisQyZhCT3MSYpZn43fLcoJUA6+a9HOyr3oo7llaDoRMxLGKbAd
ufADrxpUQxSk7ZpSEfKcV02KwS7YILojmaahrbgapNH/wMtPwjBHCqKi8JfRnYVV
On8yhmn06IyfBqet6xiXx1sYBYGIfA8qoNU0E3Xt+gMkdPblaTuKH9El4Spbq/80
HDJ8wCCaFJ329Vsk61EKX5teA4pGm5UvkhLx3l2g8ImCZO5wd9Ayrp5GGdDs1x2g
SD+Cm/o+wdQ3WtxcpzurlJP6TDvMYihdJghupiz5MazoA4iPc/7EZtyBSX9O4Xwy
JsHMJhsc3/FKCv1pw69GlMfSe0MA5l5+JfLg8s6dfW7XRh5DYoRe0vrmvPNpWbpG
AmyrUC+DG533pxaFiq9e+sznU3GKbxpOMXVf5ZJlKbIu05kYOgTLpZryXE3Qtzw/
VFOFQ8/0N3niZjeG2qtnVlDcbG/lLkvwjs5WlFZc7qoqi1zV/Gv4wZ55oxhd1nZc
BofV4poG+0Uh+B3oY8E49bkk8lm22VF3AJ+9vtF54rqnNZqhpaZGA2f03YwSSqiL
4jDg9D0ISKe3k13D9cS4f2l+8GgVYwsZ7BudOMeR3eeb4zUiES1AydtZvbAZ43KO
JSE/KDZJI4dPR2OrCU4u7kAVpOZmobjaXhVr6USi4wcNeweHk9PD8fG9SO1O8yGp
erwIPR6z6SbfrthCLEM8hgj6LWGEwD02KadyOiFMo1C+6S1YS1CQKAa9Kism9L9c
6OrL4Alm3gl9Gs+QIqpJV8QDSJHAAo2IpkcPZ/gV4wuhoU32RXuBiIwPAfDfSAyj
FBKcyQZ/S3RYEAluXU2ulyN3aYYT3/MxoRnDU/emoUYYiGU5MHJ26MI8aKY1sk5S
Psy46roFxlhmvq/0gwPp5Ab2NuIxH5/xD1dQPLqeZs83dGSkOLZl+dv3pm1tUSo2
99kUREWGC/+dA/1FX+Q06wh5L+DwVurd6rXRKX0jTyXSc5WNOeEdBkMZysLkHLRs
EvG7zMLqGU1XmYwGEI1vwaJ7VjEGMVi/daac0w2xkZrum78SulmAsAscMf+rssSH
r9ewylhrEECrbJ85RTzENhq3rfV2cii7Ck0Bu9KLudfbXSqVAykssKbNcbfThXk7
1/A5pO0U0Y9ZpHvcKazBMxCTIC+/IQ9qCkUJE2Q7Z3LZHeOsp4xKHFSJBTtixGrc
ZqbpmCD4R99v9zU6j4RsXIAGND0UFaykXTr6lt+fP37eS9EylfpM9s2Rz7HUXB9S
590KaWtWRkc+z5mzD0u9sUoGms0QPNVp+ryGkKPJpNOhJGWgtfQyjC8ZxK/753+a
oANg9xEWIekV/U+XXI9KDCBlnEiTEMvDfAVVJ3+jGnIl3z7QJitVNPlua+e1m6t9
vl9vLic5tSW7RMu9OJOS2cYMHh5pSYaHgF/PT1hpoPuA2GBWR1TggUpQVfuW3uac
EC624/W5a2XkKyBkwrR6gfPAvqE7I6Ts7fGHJtsLUxb5Gy+inLdIahKCqDY86xbO
YdwASk3P+APsEKS2G+GS9oajyN7kAaRVDAgoG1lfUU+FWAjXnWEtXZJRa+WOIKrc
jCnWqGnCzPpwS6XkxxdA6r99W8PjwlRQpFGJNvZ5aGcfyOoK70Tr5v8hY8vjOM8n
0gVKMea2mv6P2eby6rI45I1qLsrBApQ3vVpmAjIJ/wd0CzuyRbhPi8fUipSsJs9M
59g9SBZWPxBNKkou93ij/WjD1zgkbnf50ipJEJGalhd3wyMSKAEYai4/PZHwH1ve
vix54fqPuLT1I04aWVy5+zhlk3K87NOTmgYiEGhjtrdtG1T40qo9gZltXJUkNpxn
uNQdPGcH0mM1UH/lHlFheTvSBAj1FiTuT9vwun42GHjfzQFeztCz5H2nawTvSpTL
91nHt1ki3YpKJlz2NA2kRR28IToF4YkLybzrcukPRYuZfkDdfTCkrHOnrEpPLw2h
KV0x2+p+tzUSBGFEWJf6NAkXHU3ieLBXw7khUq26bbHjj4ZNBZtUe7UZEu3MyGvD
0Fipyntp43SR4/eXFjK4AUvb+mpIwXXMOdZtv939zR6JqREhhy1RN7uOffSc5xfa
FnkuKp+oqgo7Cpp9T2cbRp/aLI/BuOH6SH8n085/SuKxlSLzFo4RSqun6FBP79nH
HmlW2t0/dZADNqfE3hroLZZU2qkiHJpjvKcCTMXoX2MfNM3JO+AEchn3hXJURZbB
W/ZFFA8RqC+rmS6dnmUr2xgwh7/r8sFU1yLkU1e2vI6du97K8bhbY14et2QaK5No
FEK19BhNBcIxssrZs1t1b8lwvn7R1R9f2Gx82oFINuo5asFesMYaV5S0mTI9mtWy
ogWMG/jBH6keW2RGUtEzgMpkxFeaoxo2jcoVLOalTHKEtP+n4aU3edaREzITzsuf
5/N3Qj0xrtnsbxZMRnuLMmSr5238cUr+ENTjjKS2ee4gGw7l+Z4izbeGypGjrDab
2yUQpvqqZlllEyKSTgLC9vbRIFa0Gl0jYdL4isuVJG4UYWs5csHqMa8P7XLVCBFw
RgF6jkgzIDXSZlBlBnLNluN81dFEIrpsXh/LStucZL4/FfHPkGcRYklGZRn9ih95
HRrbYG/PP/bBCq9m81OE9TaXoyJAE//RCpYAoAA7JAmplgdZLbcApXpwPq+aH56d
3gHHXS/sWvztI82w8lXBdbPDITn+I35p4S4dCHhnmIy3yV7iZobiWRTbF6iLR/LL
kt7bTAw7JvRt+bVxbLEqslez70z9gGMsnpXgXRICPD6sn2mbP1QhBO38+Vbw9j+G
JvN+AFeCmHQcRL/a7NBTFj72FNIxkRG6/BDb+t5LljR//e99rR+0ROkeYSgO+1vj
pvSHj9h4zj/bCJDyteJqRSuwVGcm+Px7FeiSgJi4fosS2MPSKgn4cKcCtj0JCZBa
IMsGfE55GO/jmZOTm3YfaVBUULM0yuaZUnWQa9b50iRi/F5w4pSokr8CKjTMP8PW
eXUQSaU+KVyvNPutIJ/2WqYm19tbPTIQE/QoF5OrV/GKhLsSwuwB9x0u7F+d/8r6
IseREzFLmOJb0RzH2Q+7+dsFIXspqVFLdaRm9a5VS+OGJZef0hCNGQXU5f/tOQic
WKnGig0PaziiZTGXKlDkaOr4qufXNf1mEff3OIl+9CFQsLAASFRPc8lgppGlBlGy
n5epJJ+H0m2lcIF1g3o4mMYYp9YUCR+pQeBfUSnFekAxIA4Feqzg84itTOfjjDV0
azlV/dr26Co+2zGo/0j+oqhLwVmHoZBOmRWiyEQlWLS8fW8Pp04Vo2Dlf7iqeiUk
574jkY9Kde305ubBUwHmu+zXZD1XU/9RE8SwXNTuBbTjw3FuwevcwXekA+lto+eV
Daki/gakqXhbHDMQWNnDU01BHs/ySxJTzslXH4fHkN56uwcJC+Tq+s0QoIt8RdTj
MhEAHKwavFrAU3TEgkaNFdhj8TfpjhwVLKubw+/umo0oWS4n4HcAmOvTYbycmsDh
NQ+cclXATlrrb3rb1UTKB7j1uAdV6B36bN2FiVL6TzDH1879mxfg6h4JQbvdW8sU
gfDNlLyDrthhy5t3F7MJnnjbbsUPCYoQnVZbk6s9gzu2l06ePL0tmFRUHyfs02fJ
DeT5wo+3ISZQrr2RfZrhGACWnHpqAyEoa+RlDHDKzoFUY5NCvwMOjk+Tv5X7jvkE
bbM950Y+W/qt4Vqcyst2wmGf3LCfXz/IR4/Fzo+kxDYOV/ik0vzxZf7SEEqKig8o
Qmv4D/ck4ABTfsO01nbC6OjcC64miT+ZWrcgpOfy64JkaAgPIIgmgazRleDDZnes
GiWJ/TmvWlNB8jmXDvzk2tpwFpRjhTD+1FwJnKypidTnbgC5pjngmyY6ncF2wg4G
aZMH4xBnnlDuyva203MRG8hCSGBz2r6fsIr0aacHq3Q1fXEdvMO9OLFFr6BnS2UA
KbYeCkvN8evbRVpRwt3Y0MjBrfd7BpFqlDsRbcxuCLGoW3cOM+U+M6KbXIYQ0r0G
m2nqoevbZkUS8tamg4//sQe8/3FY4vgb7htUYs7CjuI96Sw5PppRbIpYAGnytKjs
kgXwPorTeDa7EYMeFfRrj1xZB7DoNMIEdeL/ENKHz4gzCIgEZEHqd4C8Oz+gcvKp
vKfVfcHgZIxh/l/qWoeCgmjalb745bXssDucLg3aITozc/gFqewt716d9XyTefmD
ZO43ta419fBXqTnp9+Gvyh6TQjoiPiAgkjDWagwYysbTVBtCkyfLexb9zQkvUr/B
Pz9/YlytdKWkRLIdR8vALavB+oI/6a5vGh5K17pW334f7/gmHrX0x8kCQKae0++a
X+xZBVBSUoBRdp7AwOAk0PbkcyjR+ijSZsZNMvoz2NV0C6m0zKSWEB4HkPQslzsP
1/2Dm4V0EYYMYNpXOEtjHnX4Jvp6MmGjeMAEJOrQbgHOr4TJ4PSH3cXSbiNH1gQk
oubZb1WY3aI6bzycfKeuhHY8YVUL5W34b9tnbS2s9AtjyTldzY/FORYtLx6IiAKp
xqkH8ke4As/QjvPMMpOE33bXvziVmmIE3oWM+VnxmI1wj3QHky849A1m39FemHpM
7mqXOpzT60AKVSizMahIrk/EluhfiUxZerjFUw+1MPTqRmXmGsSrF/lHILXKzvXk
TNQlZMDuSxdFc6nfNPjQlYHLigHu1KgXgnOx+gvpZ13W9v+tuJy+m9n6HyHB13DM
VshWXiWC56CHMNmlXeV8BZ4Me0P/TShDrA2Gauy6idZjkbw9NyZ+szOb6J9x8BlS
q1E493jDXpSQzOcnjJnLconfjUKtnJEUZGZJI2mg0UtL4fbgfurIkN1Muj4KQN+q
pBN/jHFqzaEPgi+jkITR7oRDM9WprNmgbMTh+pdBpHBD/LaCsowYR8V01QRSH2rd
KQ4GvJaTauZsfEGW2mnaUxuB0q0sNczc+bmjf+FXYVO0O+GaW5QXaQPGkc5LZYzS
oauPmmDAfrAVCPbrfvytOkeHaelIX829sHyjppp8wKiAcv9L4W15TbeHkxs/BRwU
8m7glZ4wmkk4eLNHDHata4XJBtUdMN9B5gAzNSF6UyHlsi9Si1LHBR8MV/OslAYo
U1oydURV9+p53S6igp4psAIKcLYCLAbl5AUTk90qfzVIo9vzfwdCKt9wXp7u/Tao
EbTXnp0GWOJF23MegZ91FRyESY/JvKEShujECVPUf5bgXFVy3519mXY84pk1Zueq
UwS4xmKm3Q/vLp/rDW5TaJY0S7rNbOhMd0amxMzS/efCenh0NSufndGqf2pAyN+l
9Wl7lLJTImPPqcnRyWJTPjMfWu9Pk/aRznMUgjEwRFKscgjQCH4Jg6AjvlM3opSB
VzQeYObj9k8aFOHYhwsKS8gk0Hc5P9r7OVF6V7kPLu6EkppfdeewubLfBVyOXtzw
0UoeImum87MaRy1pcNJEjrjPEKUToqjgwFO9AfR+PXFI2sl3btP2RhRr83zyJFVv
cJNmgA8lksPotTtS3E5Fj2x7bTK4Xh35LaS8IO1FFqKuC8eYkHA8dRE7Bzfxu57Q
t9GhO/hGogmq9rZs7yA7YhFg9R1BHwGRPGZRD4yTZ7qgWVzhmD4mNU0Qp4CJ5GsM
z5iqpSKOhU51/I2/6L5kXF6QSkb1y/X0oMMlW/7Qz/E1XJzCOF785bOlo8xfcnFU
Kzx2zduRtU6KptUZ8vUqYwzHDYB4002kVdA5HB+LLPvqxUWn5EinWhDQTRP0zfqE
rAoTkOPLJ+HBTiqqC7fLVVHkh7+Q1Dbt3ZqDWDm6xwRJFf8tuRyFqdyfu/DUkbh3
F9BE74oarUvINHYSyr/QJ2CGN8R4+jq/Fbi5mmJAco0oiaEBYxV+PKWtQQRl0xrz
eusn9tEvknksNOA78VWZSdEZtO6khKYIHhGe7LD+96SFFvJr/HM1f5678JXuzM4g
iPSYNicKCrUiwxxLOt6RN2kHyCzLU+2SNqDRnRH5t7lFIG29yrlFtrypMEzJObKO
R4ggmpWb5YG8lHBA/6Im68WftL0nFqcUTGBrhKPBbyT6rcf/mVJs/1uXUTjbr1zJ
/3M1mQDnDv/+obFdJF/LQI65SyWAx6eZnFVsXw/Oc++Y1Q8+fJNIkuzIfffJ+EiT
updOkQlihRzGUpjd+HBDrbMZz6pwbFWvL4tIUtpw9GM8Pr+urut23k9SuiBiIN7T
s2ugRCqQ17GCSFU6WS7ytDId8aPFF3XMmyXJikxjGjb+4YndGv5vFoBVm1LrvX+u
oQL8jA4g5UV3EO4jEWa4yHUX97FKyS2rbP+STCW3CQl1COVoeet4lgPt6WD6uVxI
QEaVbawBEc4KgcxEF1Po2AJKAlMDThSyBKuFa6u/zHHF1mGXydtpFOMbQfb52hpd
SCP1nxWBegyr/lqPqdH/6lsciIARCFGSY7gm/kwV5iwr9lDTa38PYvR3v5an8LLT
vG0dh7kna4npxMgBdu7mDR1qN8CdcBsnCWknIRrPTmYrFfga6xn7ar5DN9tCfVDl
4zNP00q7nAqyeWMe+Mr8IkifLKTFS4hCIILi/fHjEBVG5FIp2XFc+r+goGLFhno8
T7KnmFifkB4T+/2vag1fI3ida8JjFIdxBmdCHc3herE5QZFF8pAmlmlIrRbIGt05
f3DROBXapJdBEJuOUBFN9rUKc9lR2yVRPSabKHIpyFsBy7f2DX6Lt4LU7OYPvQGZ
LwpP8JF4X0OdfU6vdZ9Nxc2dI4xgeePFU9YCUIBbdudwDxpJ0RudNsetuhZ9ISUJ
UWsnjA2wYCL5NYk3GJQzA0d34TrdOxrHwu35gifeBMl8Agv/VLyFI1a2dvZopPef
vcIMTuAmmdngjbUZ+hdQWE/v5u29RW/1Rlif42T9tvKapPlKAKh5ZqwgsF/P9e/V
+Z4VvZz7xzzrG3wyJaIBy+Gz62BT1HHpydwZwhPM6RPtK1cmbRGp5OoV9MsKcG4c
jfxeFeNu03lnIgfylx1QYz0UpG84KR5zvNcoYwtWZK4o51pGknmHn7Sw879FHJSc
fOdONnDk/enSUMU8pMRMfCsBW0CwIjUKih3119gdEFE5zjjG1PLTAFXYQDu57Tkc
yP85DOy/hYcpdVUavAECjAv2mNe0gjDhMlrN/6NNxWlgAonkb32UZUTnZgPxntUI
QVgvAy0hkclYEjdiIFy4yx2CoKSt/92Wiu8EGpZ4twkHg9SPpuF1bjx4v73/8sCX
Vps93MbsQhCOJo1Kn1xQeV/1Pp1UBnVDb1uLj0yk+9dlBYJQaBbbwt+9y2+//gC1
02dl5kKHfd3Uai1ad7AZSxiGHvJOihEzxhZDag5fwwg3zupPjHCi28rhRi4gfw/N
sVXRoEf6/wsptmoOk0TmubDiDcJxwehw+rg1CrntMZVVhENc8wIvLU521IiUIiQ9
3FXJtpOKnWJPWMBdoLim8GUa//tD0l50Lxyx1vRh3xVGYifzRQqHej+hoYdGIV2t
GlMtGNtLaeHJYdZjIzKUepKBJpo3tpWw4LGt/1ttfaTY9x7kdJP1KSsZJRZR+tZt
`protect END_PROTECTED
