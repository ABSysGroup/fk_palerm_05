`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
izM2UCUJ/U8ryvpSA3KoDYBBWvn4cm1maOgxh4QZJb1XiD1tHQ1Da8Ujv7LUt3b/
rgXwNrmzzWv9JpHi58f7dHpSYz0MHICDUISG36TSTk0fHgSSUOi5m7SrWrTnysnf
DF6NecYOEZL7n8okHRY2SnzjqMIIPZL2Cr//jnJPnaS9mlUi8fml304F4pY4Ij+2
c8gZRJwfZnCmDu4Zh2AOKMsTeFRm0UT7jAllYDQJvXpiVMxYZaYbEzLS+3Y3ClKp
ie1C2bvS+7gM+dWWgbCdTg==
`protect END_PROTECTED
