`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o2cHIzvzZvUaHbJRITGUj+aETVL+T5yBC+gw2gPI0o7jfpsnAosHoVLUGNs4wU/0
/zei/Bage2545MxOTtVqAfRG4mvnhad5UPAwIXZ0rFRl61R1yVN/MzOQUqBSozNR
ravkHaBQbfgRfY0Gj4sl1LtKvh6fGxcHfbQUd38eZpe1MUwQRD8mVxDBp8Oc6w2N
z9vzouDfwnc8QKVXLx4l7ZMEIuKuzreusNjhgr8NnbU9XKhqZW+ourC/iQCI0/l7
jRiRMEwB1LxplOqF4Ebp9I28lgS6RePxxhtlw3hZ8hzxNe3LQwmezJd0OLgxJ7z2
aNagEbn7dR7xxoP5z3VzOgpeS9xS38Z0qr0S5VfSPknBa7U096MT1cG7xqFIb3RN
c0j1LsAgt67MyQrIee+woxZDjEmILWJvaOmdA2Nf1gqxELYIlbn+P/Gn36VDPLA9
CR8ws59vZ6PaHmNl4y+eIZSGBWIj1p1C17VbMi2R/NcyQfwmedYWFEVnZtTXUMgR
sUkEX9ToZhG1nwMbqaCdJe6FOQdQV+vQiKm+iX00Lq7Y69RNMlgIXj8kCHONUGcw
tjVeQIjQtkCyYzWMVRDcXe+J8hFeF1NsaotJqZaijJbyqCpbGgaGJnY6ATMcLzQb
GI/3mpaD2rN81zAsGonXPiMrCDsLDZaoS+ukQ9Qt7itKbPDBjxS5M8Ftw8qUNr9c
575RgOwRwOko+AaiJtaKC0g2UOA6k5Gl3ZwV2jMgTvX77gDJk8ZXSqrcJ27BgP47
KsmsoHyx5m0avXaSUa7M9FrESlcpO6XV95lm8Xy7YaXW37X6GlT4QyMeGmAJh2Vj
ZQFs1bEdfU/sfLf4ziI0p+UxMuNBtdoUu+AFzaQrtst5pOwwUHTBvb3C5mggZdh7
KIr6/4JO0fLDVCEe170+TKS5sveeJ25KDkxThJKznsBJtA3Z6RVR40Txhuger0Ug
qDYpPHTgkq61Qv853YydayE8oI77++rJP4MctLotJHyTOINN/Lpvue/9FSddyo7x
l8HZvQton0T7+iQZkCEpZsRDailnKgXmoIf/z4k7Q7yo1yf3DHMWyhJ32pnSHJfR
iHUSDO5ZvFjWJWA12SeRt8cvISgrAjTgyogLDSkJJHgHgzoYLZqPLrKTQTNVF2p3
G8KuGYdl/r6uLaL74dw3EnyUzeqzxYE1WTiuhb2TBS/mWjCpKwNN+0YJ7CX66vSb
NPQmvSMNjMJsUh/p4QM2JtQA+rh7oHymimJ3eeS2Rjv7I8w/9xu4mce6Pv9sZfKH
m1/oyp5PB5BP0Lr/kYIUZ2J1WDby5o3f2Xx/pkQvd6KMr0zXFdyJPZSNywuBKNyh
1IegAPcu7pEKQ0ulvnCPhN42tDWixEhJEOYdD2TWBI0s0U3E69VJcyjGWe7v3frV
5ZHDu4pwa2kdl5rNRjqm8ak6Qj3Gn/4Vywci+B190nA33VsAbsJ0qEKSmUrqZN26
+xV7XFqhpKBXsrWy2KBdy+2q9u9KonVf0Eyxtm1qPS5wPlegB7YCuz/beZfv1YNW
dbLeAyuDUoAzC+Y5q7diXcOxG0vqWB/hh1AO/MHLdV/BtNr9y7zcodG+rJpqCFaR
DvjZE+d2jrBeA6si89HDKsvgXOhvRWiNqYTla2s24aVTaRJxz4jbcX9OSHT93ami
5QkzNdT3stlH/CwpesVRHMPKZNHGgXTRKz8RDfkyjcEzRbu/DZudufNWsqE/3a53
CP9h6wMq8Y4mPUfExbVJq9GiBBGh+Nq+VGbWc39X8ISVuCfZcUQ7poyqos89MI6s
eY5OHoaWE2xNTvhCxZBYZ8UY1calQ+VBKTXXT4xPwEVvE4uYiV/DEUQJlAa51brx
4vZJg+KVxfVt8YMIhI5zMZsb03Lxa4+QJa06XGma1OEgj3soWwRekHZGucXBd+Ho
3Y2Q8ySAbIhEXcYHCsu0AKK/oW6xWo7yQEmhBfm5lTi9kJclFmwnjc7qRlrXCtR7
fnH2aVl04lYE8SWl/APRulhiyS0avQ5/zlkplqaDLj9P1RLHBZ3janD7w3UL9Da3
pCKb1RwhYVyGJLJVkeahDi61q1fOYGHRkrxq1A+Bov0Ft1VS0e5U83XYYRjitNKZ
Pa4NNig873un5lSNfhKp2tYQMwD1Dm5NFgcf1ARxbLa9TvIfSX8P++2m/87znd0O
3CJnrbur3l3838GHa71gNCyXu6HeiplPdWkb+KNksQr5Hz8Vkt0kfdJ3CAdmT4Q0
Q896xB0AiFK2DMg0buvy6wBCEcRtEZW13iIId125VqX4bOBfGqzUlOamRZViP+9k
N1+qQOxa5ya37+M8O7S6/fyv9MDfTG8eldoBbdYl/edFKK1PdTJfeM0awm87Puby
jj++d9vIRwhbPkP7uGvX6ilo02cYSc8CUgCt9LAXLx95jOklDX7ZiVvff+ZOAQzX
na3oIMwXujfXBrJ67rVf839+IroIZrwa/nQZiqqcYlPwFTEcxpm/cnaxBBLKQosa
WsjPX98jp/MCzuBfdpxgXlKVG/+Sh+9dcoS+HM7I4Bt9+yxsODy3Pj/EynTMbywX
r607MrEk/3e5C0lKE9KrQPLi90zgztbogAE1ba15JpleRyUab+QAU5u3ljAdGfwY
ctvE7JbIPj1yv9R81jiAZusHOX14zZHAwPWqi1oNKCa+KhrfkoWkVF8zdjlWM1tN
FH6taYZteDubULXI7sWpK0SBV1TQET5VnrC5L11AILVNPnd8RS2gQwM7QK3N2jLl
4wUylP9ZlV0Lz7QDHEV2suO+OePsEyQ3737ESfLOmQuydAk9REH1JUS52swbEUex
Bwd2p/agK6kXwHE4EKUZBTgj472YaqJUE2wyqFC6gLynlfEQRpi7zLIlW/USG3zk
mXUcpM8vH/6K9iMGsJ5h8fOcBftkx8sw3y1dNXuuhfdj0H6fp+5MiXLEuQ33F3X+
ZwHuGnzFAwtwllEQAikTr+UpZcfxKTues6bZnlZabV6/obd5F5UtoU6yqN63LBxB
u+D8aQ9TbKL3BOO8T3goJElNG6ur7t4PSeeywzRxAe/7efIPuvYtAfM9Mo5SUBHJ
1xF5k2trOfXy6xAToCVzOVAW40Afx5iYPjJxifhVzeD7n13iG3bD/o8fzsUvKUUK
Rvl1YuAR+Pi7QbEKbehq2Yiosd0CI5R+SzpH2Y2WcDEy+Gp8ZIB0tqc7FcKu0lBe
tPD5UDHOX40FhxmnIZQLMUMhGu1nqfb3vKw2lgAViEwZv65qJV7Agi9xAROpv+k2
d4C5uBDYsWum82aMAfw763lGYBuDbtiBU8TnLzHY/ElNOyC6ndR7pyUS8FG2IpiC
QWqa/bR4RhSFcRoPA4X1kIRvumsR0lI8iSeP9vnWo0DX6sdzBFiOTu2g+4QWXXlw
Qth0mYEh1et3RGKLp//vUIjJ5vrcVRxCMh9P/fDKt1Y/zyMvscr2sredN8tYVqCx
TRK93u4I35n2hd4r7lxywEy9vi+rOk/mB70D8jSQARLbmLMdlaxJCrzLbOJv8Dm9
lPVzg6Vzmh/RgzoPDqTtez4iFgkppnUWT2+plkj8zviHAH9gu+ddkYzyRLVEETIE
b3BOVMlycb5aTnDwCcd9bIXz44oaNS9Y57XdLiKAG2VwbG3nDLwzkgL7Hu9U9a0o
TZLVM3gIzE+5/3svWV2nW3Fjc6izMsRJZC8WYpf9LM1JyNg9S6Ve3tpE/0GceDrS
JgfKSRWmZKz24Bg+RPiBQUL3fQkxVRMnOXRW7VEWXxU3vaDCMPRGLp2CZH4/bn83
gYSunpeEoMwJ0+S4papjgwqkz2E7CnL2ZwVCt6KZevj12ybu6mU6l8+ViWqvQ4qd
4QkloTn4nmFLq/rl9NWQUkiWR20qyczNSmB7M1JgxTsQmb7uenFMi9zoPkGCRV/C
CKr22P/x1fflHBxttzazz2jemq+9xFsLTbADqbO2Dqotyo9rCJDz/9XYHNpvc2Lp
VJ9NAZjeDETyvGOzwXFi/fdL455/aWCGqEgwNDLdPUCYhH8w4C8STRC/jkb8Nxvg
GCG7U8uMeZI+KxGZPgD2UJa9iOYap3L+wCy3Qfqai0vNxEMVkSFtOtsJ6TYE4ov0
Pz4FBk7ytJF4Tmew4sefieQBL8CMrcmC2gVy+iUjVvsUL7OWl1Yn2OvglTdErmlX
nY/9Yo1FXu/THT2Ydyj6Ey9C89iMOmNi2j2REUYNEWluN05VXK1OPFfbd133W5PN
aIKoEIZB66YViI8pUyM1Pd5UQWLRcHVYUoh0Yq+HTj9kMgXmBJbG46isU3brTBCd
36yVamDId7cKgTipx0ThcIog92lWVIJS9SVKskfWySuGdteaYRRuTg+755VcA5ob
K0ACE8TvgmmAuDzaxBoCSmqFzxEH5aw7SwW+QTP3SGvfg2bX4VtI05BjeKyNrs5K
+pZvnXuDMtNbO02Jugx4FRcv02gTD5u21UR6mxnhDou+IuJ3swTnH4G3pNItaJxi
HvQ1Nzz4q6xCSfYiryb6QvEQqCpLXgX+G53FKWsuoy7gETMQyHy6cAXrdnIyjx5w
x15gz3xY1STb9/F6dWqkv7YzpTAm6cqcfGaLTcxXmu21TNepbTwfbel6CIzLuPuu
jNI+NM+pfqBRv+Xp0xGMbHyTgxzqdCRu8cauJ4vR7v6dRx9qG2zfvwFhi1k4I2u+
tB5D+ts4B0SSBSyUaTacEQntYiPM8qL9HkVVwMUYHlJ+aHHrKVnKQLq7naVCGsnU
ntD2VjgVBtAeqt/V6AUpcrWXoy3V6x7+fZQsdYVx3UY9uN1gHf/oHyVLIi+vT61a
9HjMDsLJC6494gs5Qsl/Bh7fp8Khw8zHmj0vOwJ4O+no1FZAm7Csx3V8S+MYlexW
vtNV4KmWs/a5W8kM2gWaeZ82Ee9JoZcpBTX4VZdlCAS7M4fSXo/VETOwXvyhrMJT
2hMlb6b0snE+XWZV+WoSNEuqQJUSzQPA/Ngd5UHAVOD93erWhv7PKq4dBh/xMp1G
jlyRDiurqKl1viUa74ZAgsbxF9BOQy8wSvVJbK/0K+ECMLkPG1NF4eEfL91NXklv
5nYigEZlAF24q9xt9ESX1UjcKtZt6Yay1Oh8p1taRucttfxDrw7pihp6s0YQb5vh
ir9aHsY+gpw6VFjL/tGsI5dzCcQus+MMkf/X1JT1ujMv+wr7dxS0nyq6MAkIlMSF
U3orUehozqJ2Lc3HkHCOEZq/DvrEsIMrq7jp20fMafeZelDGeRfg3zhlISBbVcQd
ZBKrIZ8m6nQNbDnSGQ+Rzxly985ZdFPwRBFkfyuPqbHwUh1Y13KaTOSjIwy9asRh
Qcs4LfYeGqOLPAG97Y2CGA4iigbMWrEBJbkkjL+yCIuDBb6GkqiqxWg9XNDc3HWy
l/t1twm9N6+fcFif3Ci6AuQYb0Odmb9NFMWvt7LPeZYmQqpbAeB92r7FnZmFq3BU
FUw9Ix87+qfjR7qSTNT4Zsa7mpRiqOBwBhSfQxw+tciFBGOGo5T6rqllaCQKQtW8
lG7pp/75eE5JsMuNtY3pp3LiYr6otxQMC6dDivb0nCFYK4j5XhBnCl1AdJf22VuA
t3kQmxCtIY18r6aY6WHZh1HuHi19bFPMwL6ZOJ3HoCocxyAyE/9zM9DONCT+26c2
Ny7La6HXjBqis+QRceJQNVX7KlGKplJGwMJojH3MhWCxImFuWDbzad50SiDZMHmf
L69ZSR+CgfwBv5cVVkYXXps5JPVmUhrYX4+/6qomjTXeq6bo98KJGoZMgNJm6Br6
6KwvfHJOodhdwwUWPsiyVfo72Y2BDjKOiGQSY1Yhvygxo1/01xkIzohbk5+4xHZ1
H8P/o3LaiYc4UF4T8ZMyh1eNciXq4gh6XghihLMISM4hjsCK/dolMBlAXheVUg7D
frqS9mG5yEyfOAcSb8B9uAWhwk6nuahSvSS4I+zVlvoVSWyMaJABeMhz7wEo/wyt
nabwbExyji3Em9iLghr7rbPo/cVqfzHOtAhwUy84twafh97zosVQgSrmKGcwyqUt
eqCaClwiqFyt9ZN+hKl2ORkReX24gxV0BzEDzpnOdSHjpiKcfDmO9nBr83ah1s48
5yR2kGPbnEhfl3KLss1zI2Yd+h5zcJPMth+igTuqiwYSosRGhXBsDkEPiMAa1yBF
QrlB9YNpq1s1dgZeScKoINghKI9fRsV5BgfZHN6Hqa9MjuOO4nSCOEuw7bC25FlE
lzclQsebuIiKK4iQmUUcl9CNNh9dHxnmvg1DiwHQPWip3HiAqiY4VvsURquo+TMM
8moD28FMIU4VLKQGsrRlLNt5wySJEVxfoyzQkP5rgkuOwZ3R9yO07KHUEAdCby9X
5U7tUeETU3R2LhC+0FkD2uiFF89cX4VAvDtsHmAQe/VyoYWkqh5vQtQV8NvGlbMv
yJdKfCgq6G8MSRqHzh6TvLszul2IywtqQJZN2UNKUHQkwsJ9vK/TyFip4payEX0Q
UT4WonAJar2O7Nab+byx2NGcgCAFRXQidkbHCJyE3lBxK+S3L8ZOfg6eMhoKonR0
faSKWzHH05e9WdQ4j8Ca+CrXqeWVuXIgRvO2rZwkha7zq5JqoMLyM8jf3kURaKZ8
4RXUBcgBh1NEmG0cfdsPtQJz3ZS7kdSMVnKMgZogt7qdVzZ1eAEXvn52q7xSBWEr
IAKuIr8eOvyHSjbJq2nKnMRFjYs7h+jt3RwxVYcaQLWyNOQ3WZUkLg4FtjyusKN6
5W9QHammlzgJSlgkeSyjVhwAt9ApEHjLO3icZvzttoY2taZDA89fk+3iPpRP0sjk
NisVMIZd3A9+8mjz9yfI6qquwX13jT0ODyef31KxFe52HcQbv1DX6g3YKFKIQr/Z
VCQm4A52a+L4PbFyRL8eOhK0q1ekhbX51H8uMrqqldWQvCDO3t5lx1nYCZB8EUSl
9My43oLytb8LEyqWEBna5wad/I8SRs6T31sZpGUIppOzd4KJ2PL9WqsVbq5Xm3Xi
jouqytQnMkGuVWBYXPPvDeTAfiZL8k5Sv17luRUJpreDTq0I7xF51f0nzxJQW1JY
t5aLhRT79BT/RmMM8osbOv9lSJQzB/nNBrtv22GKJjfYaqoA6LfX8uRalT0wGUfG
RhSO1GQUXZercnBrEhnk/xey88EZMl+Z25W1ELpOEw4e5br0WQHrBzlUULwY4Zy1
zILydjrsWV+8GtGqDj3is6F+n+zHWwRSkzLgOayOHymCFNHpZqGR3PgwKqpBzM1z
GLcPvzDeenBAVwTCY414bDX6EecjQCHJiOSZmQFes5ORQxQYs8fsmKsHqbMaaskQ
pgszh7EgEYeZczcl5BnL1H06SitJ2S72+AiIr9HQ3A5ElUSQx+A9jcFyg6/CmEZg
hLBKkWx5hq7eCuRLREjLbXAeOEN66LHocwfhFYrjhjzY6+1alDPp99Ww3Ogy4m4C
1AwBhmoTBONC22/Pn3mW/39tAEXNnUMZCLIq9ueFcx6uXLoNV9PXiXLmj2BlqY4G
TYM9dX4kATKGLzoyQUSNv5sfWzQEKO7ozw5C/tILfbZjr8avak2AjwhTPVUb3x5d
ZgCT156KWHkLOy8HZsabTJZI9dJqnln/EUc1CgWXksvp+DRoXQbi/p20EOD2Iroa
yHkyVR5e0iwIds+8A5s0Jc5T1GpCHvjkyZ+lt/lpZHYa8YiLbpNRj2A5LgTfTyuP
6+qQ0sSMdcKjrGxq66VZHqnGL1jNHwt2MD15Xvd/FPryLiFLvsOkmEKoIr/vbVjC
oG/5Mk5E0jJoRyALY8XMlXmdPMMz+3CNEEA0JrnvAukKpUp1OaEq/D5wQq8vf8Q6
pYh3rg0Fhc/oKs1OA8ul449QbQRavVMvziLGhDNYtpMKKkTnlAD8l2OnDeqeGQoP
jWB1APlSh9aN+SA/otXbIq70Lzgg86XokmzxgK2Gv4WTDOH/4XSqgJy6go6aTZnu
bEJuzq0DuvdSf90e0Uw9Xipptd4opJqxb1YW//Z6I1r7/6KfnugPg6kZI2rayX4x
ZMmQty24ILYriFCswAppFbffGuGbdqOw3kGLi4gaQeyRrrY0PvJxDKbf0AyfvpdX
2PYw4MEnypw4dCmjQ9uPs+8f/BjFtGTmNgqnuBTqZeakH9AY2qm/PUHqpUSmo1W/
dgLjZyltagSrlC9Hs6b771P7irnF/ZfMu1ZpqyHrUI4HYxhyY+9iKAhouTQDI0q8
Zp8OuSL9gQ0rYsC/jKTM6ooSza6x/lKy4hP22uhnKX/FfqBt4qBGdF1gfPwHKqi9
USkbYXufmuD/QKbKl/VVfjnbBXBliJTDQtIi8X3x+8EHNqgTFWFJbZxcXgXJnjhC
lJE2U672FJli32j44839ttE82T/YQ2RxG0B3w8XF7O+1k8zqPcqAO8roogtv3Arv
d6xCmVS5BJUwedEcX5MxGL7t1QKdJ61i8dep1k961Zkha+LrKJa0julzzxGxeI9F
fbgJnf0UOyIol68drOR3l/MvS2V+3Kvn2e6Qot3ootzbnZR4OXEImvE27ZVoB195
S54n6AyBgt/DFfyMlzHmcmIa4IUzOASvPNfx1GkBqVBWBG7wkHOuyceMzNGYZ75D
f4pHrQxwozS7xivOEPkLxwGEcZV/gYtI4XKUfm51EOfcrogQ65AeNZYkXbzO/1LX
wE0QtEqzUm+qrdJTdM8bUtbXtCb4GA87w2Vja11pQXFdp72mJSDyHRN9jy1c+vBM
KE+//6ipVO2ReFkxPrX7qIwgAYGp7R6El1A4XloMDTs4RXBGZHq7KWX/ROngIOeY
tLifRM602dLs4g18f8Iv1YpNM+B0TXIK+Pnbu58yATr7yKrQ2LGV+aPnccFvP7OY
yY69sbj3Gzy/hmilrZAkRurTt7IHGITNTD0O/QnSq47qWK2VTnGp5Yjdq+Z7kH8P
VKnRpy1buZnA9aqNLTkYO9ZS1V48KNS9Uun2rcZmejGKHXWIXSk1728EwjV0CCLK
yBJUp0vfRFSDJSNxVjyz8rk1h7H7g4gaP9GM6PClEua65Z9khywWT195YCqj4huM
JaLhEoRx/u6QRvP9+tKWMCTEb2LdoKjbeeW4ydOnGBBM1PpazzJr2hkcpjTFVSIj
bArdc+SR4TDZqKglCyG+eu8hoVYpbF1Ufv84/PseSGT/dPb9skbcG2djJyCbF7pS
QtzzZR24GvAn5eICfIrIHzQ102chY8hAcMxPZwnucWj/j7HHR6Yb1Zgen29A/r6y
V3CoTlL6U0ny6xcueWr07ebwxKzScw5g/pH7+lJ7fDHysSh5FglouN/1pJXnZDG6
Z68GrL7/k3CiCranMCaLy7ApGdZ13jdq5se/IszvWlAuCZY/34lPxMCdIwjArGjI
fqNiWycTR6sY+uMauXYh/54KdY33UkN+smxz1jCckPy7QYeRS8nRKt2Qkz3KRxJW
Vj9wGsZRuKTywloYuhbpzgBV3D6FIHRFKE+hfxAfEBmnHT57qx5b6Xkcj1JPCDya
a73uni7yXo6ifxhiZvrACyfK8jTY19k1tnYwCxsTTRMh2EFYfmcmXh6ez5zbXwEy
ZU/XAY0jFFuNBt6FpSYtMafQdzLrHObF3cfCFar+WjmTcVaNQT8g8NeRtAm6qTbX
nal4yxLHDLoZpQZsvLTgnCceEZgi1QzwM6RTcyCVgA5OC9/K4hWslHbimWGxQYTB
3c+pcVKSN+ooKjDI8NqtF0PD5Xz9mU8CHo7RD+4/BWG5/6lD5yJjTg870gp0rfIX
JD8nRhDB0/6jEEu0zkvW22jDL0VFn6s4AuXAFm6KAzYzNfNyCuKNGrp3T7jGBgrO
jrNkvlk+ESE+STRm1IJgX+mJuCYo6Cb82TLfFro5xAF360qDyrhbhdKGv7o1dsUm
oJWCajEbgChuZQdUkex2qst+zIu0pswm4BD8qcslG+FKLoRjtHVdWOxojzEoof2N
DO5fu4Ufa4T62LBeHA2HPrD8gh/xmbO9121SjVf6hyOM20z6mtYW98QV/2lZi/E5
FMTBYWFdNUouecmwmjggzX/tbeDMDY+zBKxBOjj4gykH3n5lqlS0B6Lon1odTaLC
/X932NvVLewVSeI6Kb/1fhf6TzyXDfzoInDEVbmaUZvj+gQM/jIQj3sG28smNemp
r730hiUnv3JLwxvY6kpwMr/tyuCeH4fqN2GtXo5XDx22ds2XoABACPGXEd6TSqVN
DbWpaeQ0iVaWz86SWiDa8zdxHztyceawMuPhEsnIrlW1cc2wCGV7m3AtL5lt/Hv+
St2bw5NkTGHpnf52wgLvlk9WSNMYb6ww+sRuUA8g2jtZ5kP9523rZcdgMnboaA87
QqG0gDmQTK9Q/0/s454ymMNxUkMUehj33Mc75IwYSHX1eAof2T1FMFklcBqxuK3O
3POzORjBj3u0Nwoo6Gm0qYX6Nw7WFWtMSxCZtEtLqx1vAzwEoSfO8nd7ubQePHf5
qha/vo2PebaHsjs2Ft3102rFVzHQsHZ7c/fVMSnASnI8N/CyGZudpFc3vAygkEH6
i/qzd3pLgR+LkLi4Eps0Ut0XaYTN3SvfWs8sh1e0kmPh09YbMIciCLTTHhuH/101
l81uMqBIulquxIfWDA8EKyc/yvMjpZ8GjkO19SdUGzzHHxivxAocjJTBGIA+8sYA
wWdYgMhxMR2F1XmKvp9HW3HsRTH9NN80P0CVu/KgIDk2DXb6VEJnnt7hCSHXf672
cZaDOHPQP4WrUd0mpk8WLKkst5DAr6Pj+mq4I4EvwIsOyAORG6ZNsBU7S3CcAVcK
jlq/8kNmnpd7Fi31PuBtARatCGau0BZUk3Nvab4clGfeXalsTbXq4AsSqurip2nw
NYjVmOBek8Doeyom0eKT7yGsxZarSlVAkt/v1pDFzC0LlxK6XlSx9dB1P+e28LON
ltZS3SJmDe5L5gVxjAaA8WqdoDxcbCUftdYkzJGevBsb/LlKI1cy9WIjcxB4M/Uj
G2/ZzubAPi9aEv1897dTNisMSL0rpvaxAWL+mdQsYXRFcz2ycDLf9YoYF8GAWegH
FEk7U+LELmhOuTa9m2Naz2jkDuE4Smn3IuyfdUsPerOb8n2V6kOyYVYHrWaDd3I+
f+AFkWV79rP//M6XxjPQwM9Fjg3WdvcNv1fecJ06ZR2IL8wWjiN5Y2qIStem9YMw
llh+ZzaAZjIme8beZUH5jGdIYqIWUbyyE5ulh93VSa8Y5beYEDg1HKb8iOiO2sRi
DjOLECst5aIEgmXs7eMrv3sktxYM+EwWNgl5qpogMi2upaoB2xpdSaWb8QUOnypV
xbutlM0gWO2t4Inp3j3aOJwlZ39KQlzdvtgDTGNeFNWBVLH4BrC0zJdrDv7kcQ0E
CeJwAHyyvuzvAzhmZ8/wkhCFue80kWffrQMI2uUhy4KhrXlNglM8auvWjwvu+vwP
p91/0FJ8nzb0H8NAd+Rhi/v3WW1wBLuYZPXel7TrLq1aPsUKVy9mNlNbkBlpYU2C
rkRLU6zX+aaSC09+uUQ4SqCIy89THOsPdyMCFJRE1i9uuaQGIsokX0/K1bTyGcww
tPrmnA6VUBlYvvq6QLcoUE/LEBZrp6hUmPhGX1hDnEUOdhKq66B/8jTRRRjIXXQU
JdF1Tx9ozsxf8JrX0WcOSCJbSM4F9SgPcl9HNWZITJiI6HTboQHy/dDIUKOK974J
xipNT1O3705CaOgtWAfmA1IazAzL3MXi0MfvrTFio/VDx/bEGKr23uDbFzFPHfYw
iaBKQaTojEuNmqyikVRlJhDnPNKjpZA2IzOJYRsD980I9Tu8olBpFs5zrU7r4Dwb
T7fRC4Dw6wXYfoJ4ySR9BwS9A0Yf83iLhv3tZET7VyTqEl/X+zE9kjNzW+Q8yoUm
dLg0MN3SZu56ji6XnUjYBqFa7f1DDt2BE81w+BnjyJevYxeiRi9Tsu1CFVtVSWsB
gXdXLrjKImyvYxpsmu/8y/nW8xgiFIbefDK17mDtRSIVH1qUkTbEmHtVp3gSQhDL
09w4OefqLvs+lg6xP71W9QPLpZ44dDsCtK98JFr+/tG083ClwPQl/eK4d2ZwflXT
K1EACsLL0aPoEZiPapv7qtIQYuRgzF/xVEtWbIJpZcpl6lAqMoaNp6MuXy09HzQy
RjV7MjvIu1oR3ePQcOGPeVj+0v3Uye4fmvSiom6GBlmlcSsPegPUkb5W5YmFPclb
2WMjuGKpMdgC+YIa1cOt0l/Ubu+dC3nDBNHd5ZS/nlPHndNm8/kOpgw9z9Lp72Rr
riuMmfLgf7c3VeQerv3xiuQBCIHE5ZpDdLlNRgo/J7CSzoDBXIfakf4kQfw5G2IX
lzbv5IQLUMBoEZturmEIRk13gPwlOcfMYXei9x1ghcHRP2KhSxqjsHbQ+Wzaqn9h
rSePgOrtGWMjBHPzCx44B7Gz/0qQ3PunI5Jc6N1iyd0zpez3xa0SIkHGAeXAsTnA
tj06lMt1YLRqXFr84ib+Je2D0TrZn9AVQLIabxKgWmaiUVyKquliTDR6Cb0tfrl1
zn1zlWAqmmzIIwOSBNo3ovAJdJLSYlHWLftIi0fZwvnTmR1MeQb6wqFXPZ4ZWwWt
iZZyfCyXGca0HOSJAC5mxG0Wtl6x82xHfBxMhSFCgDrBqO+2+1fTIThNZ7dPF26r
TQy4eSKoDMeQT+l7AE0h/Qrcp2wexL+YPY3skya8SYJNXXMR+6kSLJzoJMtmEtdo
WzMrshhg9lZH737NN5sJUtHL+hvnrca0dd7wChoQ+6dLzTSf/BbNRX/QP7+W1ql2
gMz4aZmMLIJ+5YHgX9Uwq+39A7XrViprz49lHIoBzJDPTo+0Xj2zfK5lvSYO3xe2
YzjbuWBdKW9m721j2aRodqMfPBUVbjx2YeFObEfkSHVF/2QGtcIGAlEXyj1bzg64
ar8WKi1DiNwZeAZl3PWS9wglfnqJ1MDsM6fxFZTqfDhrvDyXOQnAGVd67TJo1h/r
YSoJG4bCAnIW3GD+gUUlAC5jIdvk6UCxAUV8GolR8zu8NA0+eU1EPwK0Nfh7uKAY
Cv7AWdTr9zw3NXFef4v2d2DEThjRJkCKZpHG0TI5aB/rD4WZl3Eor47+MWKpOeOP
pQclrGhdmA8+XKkx9G3XbyBaeYV/Kins4S6TeUqkTpPNXX2wKaLhm2PSiwFdsXjl
Clgg5Qtq6kqcHHRMO5J9cLhM0A4kKMlDnf5kxWD5B+LtuihKS0WpIDex3OHl2vZ6
eG5HKBWiddXNkOy7Rcn/8pAeoKBVl4QSCDqZrTslZXrOCi0UjnUhr6UvOGeg0pf3
W1G6XmF/nLluxxki8KLN2nAVneSH+G+jSHIiStv799agl3/m6vOkuVQJplirpoFL
RmHHENCHqng4XDu3hHRCyKlYSAeieiCAVm5GkD+JwVyEaJ6h6CZXxK7B52Tu7uX/
N6Iw6Hix9dolbuI+pECsMMzO12KC4sLw0e1C0ooOTcrRv9giEZrGleoU7qsD2H7O
sWANn0b4RsL1gCVAk2q9shRm/tp03f4+mCxwrBptE4w5L+KD1h2jKHRmCEoH4EeU
/D8IjjJDeRS4FOD4zvgrF6oscYdBBp5inkMaF4qUCOX810YC8B8mC4y7tPx10LHL
kkoEpIxt8YZ45DrA3u3355bhNQaqObj2MDNvvR+cE+i9zWyLcO+bbrdRmWoj63KE
lB0slNxsOimlzyCNphQrFA==
`protect END_PROTECTED
