`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8rMfxb3BN0H9TWRsOoenVUzVJepmsVMBPAsqkyMxkc4hMiZLgAZBGZr3MYdZYapC
jXDuE/ZnNZqYjHbwT2sNMBVrpk1jm7+arsuSSAxNwY7R3pxG8jjEgSAQaCcCLXUP
g2ah46yTF3gwRMkfmbsJPL1/zd2bwHMqlrDxrJxLuNkRZ3zoPaOyg8TZqloP4TGr
RvHm9glblDY8B2uiNhIAcj8g+EaGlm76e3y1HVy2qJxDc16yRFnmTLIjAf7ncSZz
sfYDQ9193yagVSY2QKUY4twOsN+7iV5bYmBbPn46hrA=
`protect END_PROTECTED
