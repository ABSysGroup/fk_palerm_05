`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VIWhX3jr1t4OMqY7PxzxecmUKtjWljAMch4Ud547curyuaN0PrqS+HdfTEOvPbbq
cYaXer+NxhJLelWjNXXU/KqYkeyQBN3eVzsl3L2fpV0SmTV2MJqG5t9b7Y1Muw/u
KR/JGr9E/dUsMdJieMA0liA7NQb/c4lSTdQTiG5/qDXWwD0iH0xuG1D9WzgIM2+8
VYGTqmPQFQPZHZ7lwdGG1+M1tvOAXU0f2qW6BVLpQMVygn13BOjZwvANJ0aa98f7
VqpKGL2FUVnXRM3p96SqP5mv9GYO/YujEnNGCussEuRxL3NZ3L7nr2j4wKhmgT3a
EG/wvYkdH8D/5oX3oL1Xbrni9Ybd9u1UK6SSQKAIa6mB1clwtDoCgY3kmmh26IHS
BhlNb55NnA6VKqooxuwWslp8VEWNO5Vwkjo6T1P4bAXjY3VsSR2EH/tsdDovMwCa
jDebXQzLFtqPeGYQiz2IG6qqktlg87X5zu3RZfyyB09RGwa46qDr2rilxWkeU4Wh
p3Naf62Uwo8RkTSBlnA216RO83QFVXpy15leafRGRo1AZTeAt7Yel/gIWyOXP+9H
dswL+3GKPl3gUCE1dKp7XdtljDZTQRgiWisVFRhSjAo=
`protect END_PROTECTED
