`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aNWRz7+MLBMH/dqcCPsatakxONWgK67mz7FFJwFPcqlWNAGHPMrIo++rFKOz3E5g
oHKWZT1C4e3KTOO1tFgiN3H/VcuL31yOjkF5IdJ4dAbEsueDjBKIkeP2vnIy2qgy
B8L86uaMEb9mge2ZJxcR8SyTfRmQX4rBt/5kZRH8a1C4mQd7df0YFyQF74rzkwSh
xyk3onPZ48jZy8BTW7T/d3ah+XfsQrLmU/vekFU0kg4TPMrYn/PZ0RUdz8OT7c8p
7OZSmwY9THwvHYVL+dOLEGaX/tJbG21xArYNswkv/5xy2vhASmJrURlPJnlG4R4q
HlTJLptkUz5t2JHTrpvT7BDiVpvQ6Jg9YMxj2XyfGJ8P9mh+nwW9bfH1x1zuf/aZ
vCS/5ORrCPhyc4TqsusJZ9T6RsHcCNIVJfhxbOxLnUivEPG3F/htUYvEeRNRig6w
4cD4GEL5eFCYNb6N2BbNiiSB/h8X1en3IcTYhWuwil2Xa1QrnRQNlS/2RUSSxaAS
sxKVyD0KvP1h2wmG9l2HNgV6fkUovy40PmYjCnvVnTWdR1sQYVgLXrWpQJfZ65O2
`protect END_PROTECTED
