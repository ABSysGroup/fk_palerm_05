`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i8Q0nemB9c2Lt45kNqjtkx1nEB9pKn/kXmnv0s04Q8f4YwgjWwR8MAtc+isUTd7t
NG1y3hUuenjBpLM+1pgoU2uZ6g8vATRvB7djjhwP7zjLHOIWO0Z+A1761vhlJn73
zR9AN8jCynHwFZO3FLR3jwvhH6G4Z3+Ws5bPa35tQjiMvyWoenbmKXnDo7K/77Yl
tJVrj4pCREM6XT/7X5NG8O5mupGR9Beqpe/R1wXd9ouc7usGNm88evGOBOrp0pGM
q411WNpmCEfdFBv+Eztpp568FrPovDsAgK3SFSRruZTw8Qjpe72lbe1FePZuV4zw
EeW95R2Rh19BVa6b6J4lCe8T5+BCa4swcJpgPTV13EOKfi2ZTJoIYYZ4ZhnfHNvj
lAZKjlvYoHWtJs7n5a0igEsi29EYZUfKPKPK9XKiLkXaedd6JQw/MrC9oOcbKUbm
YRppHSWA6vHoeeDeBQFq0z+5vAcWkD8H9xOHJBmQXn02H7HEm+exwasfoJ6tIdN7
4p0JUqFCjb95bWCvX8pJ0KYX6zomTYIZuLMnUeXBiPdEVQvk4Ve+epWG36ngHfZy
iQXvRi5E+n2R8ruAjapxqVC2jHC2vs3MPiGaz40km0eIhW7nbfwxE9LAaYNHfUzo
yn3XunpdRGqZHrkmbrjaq8jc0yXARv0upMtZLpzbaIkD8iwgrsT2jJv+2VUf+Ju0
iSrFexWi+ZewyXH5otS28cRmZcZNTuFx2XOQVjHQKeM6RRcEZqMrX00LK4bzVbgR
KqJV6TIk/xC/GZDH+SgKAMQEOSWMedXNojd1iW0uvI4C1W4/Gj7G7nNjgb5jDL2g
Id3drgJ5OURy3DleJbJuzl6QdauCkrsuXh5Bwz3Vkje6n+CejT2WmI7IZ3ySnYog
GWKSYeInkH8uKFGKhEw34EvWBYVunvowZc1YQS1kF+7cGaN03taow+E3VEQAwyeK
+keh1JQG4nv9LCDCi62QIuPuCJ9y0cN0xBChTQvSeUkeZc242+5HVvPzX4ZmoSX3
KpaEEJzS0o35YXHQhKazfP0U6BLM7DdGfldXVkG6l+OCYZRBLQy+tRwMJFZnsiqy
cfYD5+S/Un1Z7GX+D80ySDsJ6TmZRQU7UNg80ujhWCbICxnYIOSW6ow/zUEkbch9
mJVJCxuS5pycDVMRLYg9NmMEEKXOZhmNHsQwOkxh+Rawe3roOck2AetU3IExyKNn
t2AHlh8MS62+uoTl8FkM5XEzp1xK4iZpTOwW74AVrlr+VYYTtOBgTSPpA3blVDoU
k3HpBPhyFTPNyHhFhOxTaYXbDQ4mEqiHX0wEyHTdFSJWSa4E8S545YS2q/fgPYZA
NmImX2TrQG4nD1g/ZdVOSfv1naEin74xQKfUy7aw4bek2MgWWo9Qt3dDbk1QsTu+
HyjqFriL8s20VAHuClmfvHy+payMZ8v3DjTUdTlpj+Rm1WZ1QYkkrCgQh9jrBEE9
VsYQzNr8LvJOYSma3el7/CqdlOn0RnbFLGaWmR8n3KvvwnYGT5+u5DcfE3DgSuM+
exqbAz6Toi1O9WRKcyb2KL8kQGw4deMQxeD9AkDvXSWopjpNWFhEd4/mfzLeYadQ
VHBS/HAxoLTbbDww+w2ecUoDsCmsEYkb5JYJg7Ibc7nAyZxn70g3NSrJiM/X8Ul4
q8kcjGWHahYi6PRs456otcFrI0/LQV332ZlmiX4v0aMldfs1aetfLQxqDjhKeasI
jMXjKWdRagL5ZyZzMSOWfTFoBaAQCyGTX4k4N6mEjr3hRkmUcmRbotR63yqoskHi
RYVPSMeVbYCKh1Hk2T5B8t4oQJWtHVan1r9ydb3V60i2S7/SZrqpT/jlGsiRhPjl
2u0LkMhY7Sz3pv8zWTDKdMESNooz9qsl9OWETp5Bz5gkfemhkFMnUf/XOlOZR6OY
zKkAMldM1EG3bN2Y4LoRyphInYsv3wPU1kICyvcR7DgO92YRqObWs7Aj7VYxqwgP
Jaf6VtlePbUCI0WXkO3bSEhIrJiUD3y5Vyl+UPeI17E1uelYiLMkv/NBi108dfl7
ta8WBjkThqxGmEHXIgJp3oMh4jcaV3agMSgSJkDuYTrC64iXirsvp9aRh6e11MvZ
bZG911CQPG70fYT/1029bsk9YMDwOnzl3B1QRJd3PiW0s2qKzHlpBuENGP4UvTRh
rUw+HGxInqZnEqgVhtpZJVHapjF2DupcDVwaZP6qX8me4QpONYjq3opLd5EPDPjm
M2pu9UQLrmiMClhYKvlyEdT53qbD7pA4hXep63k/Iicd/vE/nJS3FeD8fR6V8cBn
efryCAIC6PLewNoRxH5cI1VPMnXqH9J6sO+hIeQ42n/FU5B+al+JNMxDHI0ybrEL
`protect END_PROTECTED
