`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tsWC7B3WZC7OpV1+61nhcB/RhUL4qQCuq8WqdU70Q2JqErSuyE0N3iJz+RbpLLrD
+v21iyLC8bT+5AznmHoy9/D0KFyp2ZICu7+E0Lp5w8MURP13tJKGdjgds9tbg/yW
RfVw7QZl6Z746SRNPN3l17DZUFhBCjiG2jsyZIwO68D90t7iTMGxXOKSG0P5VrKG
mqCH9dbFP03SpdCvkJ/6SinWxLGN0UaI+e6ts8GIK6TZe8Ti6PnT+B0YhHk/SAjr
C5Mqbc/dNcfmcC8i7ZZHnAqvHsir/4Z4WdXyBFFFjqcBhhtPM4q3bnrOfku4IL5T
2+fH3KuIsSa0fydBZQAIYt5JQF6znoatkh3RWFpKPcRovnB8pS00Tuz5E305LjIE
Ck1IHOyl96ugHS7YLQriMbjI8qOs7uMNQQOnkJChajrvAGFl/oOtYmbJYH1NbTe1
BnkeEcPTYwbcukvRDoSQgdF9BxIokooKv6MQRUNp5QdJfchUMtA4SmuDiWpckxIZ
SiyTd0WRxevCU7wMJHvCJozIvfM0lSrIi9taRr5U/WDCoAfKLG7rjVIq89sW91I1
ex3HV3156GRakk5NGbOaUGFjwL/vkNSGQSTQ8i9LxQg0PDfk2nJnqNGt+nFxvuFZ
VYEYo5zbwy089rk9HxAoEA==
`protect END_PROTECTED
