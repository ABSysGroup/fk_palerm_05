`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7UKU6cqHgeJEJMVWiHgMP+NczbdCi7JEfAYRWj2MNQD8xbXC5+O3Zyxpk7guKFoq
jy5xAc5KXB+cpPIsYx0h2ZTT3FEPMbZUUaGzu389ClQRqiaE0ek29bOAc4bFayFo
HLjptRnhHWiDX+eopVi2dZAEuulJjam7G0mLsjnefJvYqUAybzDsKacIGvWKpFJt
jbFX67/h87lzLtsteARLHf2cZ0XEWWDyWlVlW30G+bKdaoPzHwQBSTpIowFa5YPy
YEHTVfdE+xzC76RVq8e2UX9uniC4OaBDuRC1cgzfFtbfz5YK6Ixd0aSdce/vUKdZ
/1hlbdVzpLOxxhxsGNB5nYNYpUFR/pDkZX9jjs64nNOXM20qQM9bHxBCmDGUETLR
oonnSujnx9hMvXrTodS48jzBTkIZ7oTbwGNqsh6ZbC3Vc+Hfm6YwMXinej1UivCB
r7J2A0IIdpM9rgb8JHr1f7fTSFLzPeOR7M7ynSv0SuutaCDUDuEIEYe31hSojmc/
MZA4ZzArlTj3a6pX+HILrg==
`protect END_PROTECTED
