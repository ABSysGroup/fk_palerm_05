`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9uINhkFQPok6M00YQa8xVaa3miuha298Dt6fx+dh3h+93X/KgWTVOpAWIreSJ0H4
yHHtTx4/P575L6mficVvPOph3+OiK/WUh01+5Ggsp86s4FIMQihDnXzPgTO1OXlV
ilvHBsj23BIlLLarks2Iw8VUAaBsTN7svuOkY5jTw6M9T76RV3YqBJo5ZUvcrBFz
UMnTJUp8Zskn4CVfbdVRWTMTNjUk2nd89tJj7G09YK6sajgHVmjP/hsiI1/EWT5b
7/onL7De41PBfg3Nylj30+s+ENeFuLejdQ1GI6BnCYfMzDnlOY1mwnYPw6U6ouv7
e+ftD9/nG+49NaolqkJdDsrSxsZvzu1b3QXVXvhn3zsroYF29SLX1owR5NckgxbC
1eiH2u+MzEKPhJEOvJp4aPPynk2azuSAQIEsNb+Ls2UZnYMv121Gj1O1YsUEL1Kn
rAmDti9wtaqaR6PGsTtWC5fNEk6vybqOgsx1EcSX4FoU/gyVqE/mXFyXvcgHuHHk
2Q2gJaZWPw8X6qs5obAIeFTi2vyuSB94pdt2Jgecew3Kafg+GVlA7QQDx/wQWOS6
JEpkrXkWvNR0THijspNVoaMKtR8dj4Sn69KeSkZ9hACxjc3qYjedjvT2g3fMuMmc
KVo1NzydO9UPpJWPEnEKFa30jEkUvJKudx3e4uK8TfXEsjfVxJnqTQB+4HpBkEKI
4rWRO4sDFT3btDPywrb2F+RTcNdoSGoIaX+g1JruqRUWN8xCWb0Ei+5lXE5AzmtW
UTOEepbko4OD0eZzJS6NM7VyJhFh0xPr7KnWsi+ArsqTpH2XiSFQYHGEPUPfUgd5
JWXq+mskMNGvb2YjwoleXJq6NzUQdWUJYlyJWdv2TBRkQRdN7R1xhzT8YOkkiaqf
t/fiMeRvDyeUzurOiCqDY2ScYbjxDuQQdShTCZ2AnYAKQcUuNa/469cFnxf/HxtW
ED+z/a+xB4Tu0xpnVvFwY+c0VBP+99JBbV6uJs2AyQxMJN35Z0MZ09MENdci/gvE
rzoQPaqGnaiW82oQZFWQ622A+bz/QQz/tZ9QR58styfWHEN178ZWYdxh4Qhdxfx1
aJb4jQsThXUHMkCzK+hDHg==
`protect END_PROTECTED
