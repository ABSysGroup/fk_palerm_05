`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YpVlntz2+i80xCOwPYo76QKZJEDoO3Yo3tWwNGuAlVLRzKkWxqmMyKemG6w/05lx
CRTvwa+7u8bMhXWsk9FjGewLy09mx4GxEprBy0aENTF5hMoejEEBmP8UzuXUHQZs
GVXYqs/O3WDHqM+xL2cZm6797WVkP56FNn7vHZHYbjHdE2B4Ui8ui40ARVL2FTPS
7xg3OhdWbrUE05tdm+vSoFtenkUPxj16oG3w4eP/A4ghimKyss4F+xc4tSvY27GO
F46IdIVcauVdN0ZSO2FgZJqk2r9UqbiDmE3YmB3zZND8+h8W6SOn2L1a0sE7xTtl
Wc6K14/oLD07WUDaov6q++P00zASRP7IjhR/a1+6cdB51DPNiM18yumymQuMRWJJ
xkB773YJ45Fa92enGU1Teh3CTr97qj1QdD1oMxZL1c9sK6s58DR9TMd5JdGkk854
MPDyneJ6Vxw3mFSF8ALqcfZ5VjFTJRHaqO5uQyaL4dixjPzz1bPCDa94p1znPOkO
aKf60AtIL2k9c8cDndFCaNtOCipACEviiuRPCITE/pTdFQnZUTkWYaY2Q4e5y/g+
36sgqhPD/MpeaHC7jvQi2y8DRByVmXg48z+6tkyhQCjWw8lzhZt6TAQdGuEAgH7u
`protect END_PROTECTED
