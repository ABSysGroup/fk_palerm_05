`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w/dxMZQmcAIAVc41Sa0YAkBFj/ImP6fa9ppHkx7jCdLNPL8PiliBLullzC9xHc/z
3nwMxiHJKQukkwy+2P5z6+nKyhvCqWO8zWiFGjHPvuJyM9UAkbfsVvMH+EwGv6sY
bxlL7sbqzVQZolslXRh9E167HC1m/Z0hVkEhNs38+aRbI7Uf/ogp2dYkouxsDtAQ
KAvTI5uKl582v2J8+IVKgwnbxA/Fq+THUTEP4nwYhyUJNP7WDudzrOrRhk2RHbR/
AtYAW4VfDvGiWxSWEGPGdfNSd8S05waFSGOLUC5CN66HJdRtjLxf2L/0Rpu1lWC0
3ls62DnTat91CB0n0JlaLF6qnof0B7pslezqsVMToKqamMXM1pYeQ4UaPnJMJsfZ
+0ITAqGbysHMxgDv9z0jGnm+8dt+BfCMGnCCI72uhDxksMzsbr0Y3EoTGat6+oc5
8aa2q55nEJ3W6rC5OnFx/w+O73fVSK3nQcw6Da3X109V4nInhKwa35t4okJv71Y3
fdzgFHlaY/OsX2Y0d9SLeRRp6rn83xvyG+NUim9jQtIWQtt0UtkVCY3q4y70jVh7
tsFRX5EpJdCfBJObz6uBTemi1DJIulHrDFyaB9VCjz1CcN24mP63/AzAJzwgNxeP
9VEs66BUDp/Udob+8ExIwR3/YoThtUtOVOQoJltCggOkokd/RCcnxmdEDtWQgW3X
9zmaF4qkO32R83+fOXiMDwvw9Z7s8MC32dDmMO7Xn6AOOL96lE6iaTscXoYDEYph
JVXBMNhhSUdJeNAl1O0tRoQakeDlM9Kr3gOV+gG4XF9gNA+x0KJ/CMSZ/2cBx9th
/3mPUwcWimBayaFuTZea3XoxqeirCmtxTsU5cg8MmP6B6Z4A1TK9bett2ZQjqFEh
qSHrut7h6XuWzFwhEqMep13Yk3hr0VTA9uFVqTHYa+B6PoAmxJ1Bbn9293CxSfZF
SoRpVfc1cYeyq06z0SU8FbUAtMa+6I+VbxBHlm6xzV+EfgKivyMxG1oWxfEzz5F6
RODqOqP6PZzgU3R4N5zm+x6DIz4U6DGUwA7iY0Qu/zLhlCcmPqp0DfZasoKBsnsJ
A4k9prz0lOHGIDt6m4quXML3u1c8l90+Zr8mXDiSAhzoFTkxg5BJgr3ug1FL7/xL
nQNmgqk7js+LhCY41ojMNKoNBNc/pBuHbVZLWobO5AvEe50AVcePF/Mj3h2HFsqk
FxQkoimOssTmIPbbbovH+e9qhU/BkxjMkjkp1uWUogBSkvvkR52DVhaNH06hCW6E
OCl/SJDopRs7nF+59zMOgbsVnlqbOEV7Jbaqeo4WQH0IvzGBCpeS+JkexBn32AGI
SZlvHte2vSA0CbKUI+Ec40RuMUfKL1PrPXDE61MlE2SPs1XwDlWfQk3GGLi3KExA
u0QfVoYtawkKPnO/sEkbjyVXA6lPaH1O7gd5hFiHAhXb7qkCoPS/vD/2CIKyXuyp
tWbJ69e+xhQGNRnHYEcVaO+3rAsccShl5WHv757yiavLPQtqFe+V4P0hh0R0Hnc8
o+KJZ6cx6nSlrrfyiq0X1KoZPdrhQwd5e6jjpTYmkdH8mN/MqA/u9yqmOfBWsQjn
X60TH3rXXCSPGtrKwBnAS3Jbbp9CABsWjGXdnc6OVhfSFqPolCTLoEhZOEYz/ZSS
4M07hNkyG+xzwHWkq+oZPwIYdk7Kk9HXcyiK6fMHu63ci7LjKpEbB01WBLXMk34n
MG+aLK7vPU+IRFEhNxlLChmy9ubWL7/4qPa1tl1HUvIEJLpiRQOKJSGoWAyNd6xA
tiQd/0zetKLv7yjAH/WjCwVU65q2eS6w1y21bMBvX95x+M59Z/k1OGjrMorn+sHG
uDfZKyOmxOo42F2kMk7Ss4GCNU/NUtS8EkDb65w1X/r3etO0MhPzdeu2PuaGEnrD
TvrrZptG3ZZegbZs22K5iOn7OAFbLNLwQ/1TGjRGsImscIP8zVvzQAdAiZRW6LVx
S5GV4fZeWyhwIGIfVbFN3dyfmSSpSweMil48BA8/pEEvNPWbabFfvFaJHGZvQ0+G
1o/5D234Pzw7oom5lV7vLXEsDax/hFsmE7ub2tnlb0QbQY/22rBiA0dQZsf7DvBn
CM+pOo65wHkPwCwlcMkjx8Q3GX2niUaeB9c0R8oajmGOZuuPL7WjrpXb2xsm3p6D
LWxn3ncKa/eYzkxin046E/Wmp71BvE0WEULsZM7yf49bTl71HdFOhYZVlEGLQI+k
WYeGjMi6Qcg4stz7yHtLnqZHxwLMnm37YSASP5Ntf+aeiIk3v1oXikukXOjA8Zio
HNUq22fqlQvh2gEl7Fb4aHb4TkIjv+iD7s4z4H+S3fJCpQ/EThQr0AC/hEocr1Cb
+ctlfBweaOZsvJok4APm4FzAqqSIEnWt0xk1I8Zdtx/gumAtBam6L1awrlVAUcjD
81XiJtAz/XB2kFmOwglG8z/0Aw67L9K59oeulyJyKDjYriG6pvSyhUM3lMc8GuHv
o5S1XI3qLeP0hOY379CSbCQRtm/Xg27Ome6fCdXQx/XmCKlpxZ2rjnqsi/bSjQXH
WFHMGXg0oLGCOqisby/r+urgy3zR7tfeMrexnrmJcT+QtADbkpkAIqGpHafNmtaJ
V1v3JDjvilOh9QXwKAREgaKPmcqnb6ULCG3BY60j+cv/rfAuBpyq0SRukVeuToLl
BRqr0zqpF722B97PH42P8Z7z8kMfPpGay8V8bQ9i4rPZCjMShBPcIesMHeQzWIp/
lScIEtEnCYWNdFtUO7sycigA6DR2cDqmpPAG9neM3JdqocENBip9KEy/v2oaJx6G
KWy0L8mgEJg9a6/se+Uw26prP7+jnzE2l6whvcJoggbYYNNZ+vc89qrBOOPu/UqE
/+nq91M+jjoj+pKceD8nLs/vrB3px7vn4EVa/XOewndeOwhi/FbiuUSqsJHDjnhK
BHJCyMYnetL88WCw+8q2xwahVXpqMj1QxJ4TQYepHkvOAoZ37j03qnzICZpSZTzj
kV0Q8a9QxR2LBKyUZVyEyPX4McrbFqk0YBnDodnlf/S3I74KGj5alrrIYFNJO/qK
2MRVEosbhMpFoGpx5AKp5giZNcAB8t2VwXLaJ5H2Ax88QGJ/JMQGd9N9yptoQaxF
ID9z9slhyNoHj9SfZm8ymmx01LXslpsxUve0SLFreb0AkBZILtvSp7tCFFLRWNUf
nanypR2+65sGTyTb0dX0d8u+dOBkoe+XYwvdnbEGCm+5x/J8DTSVU+BqHt1yNrHN
nlQeFKCZZclY0ZF/UK/fJx8pzc6QK0RhKS5vhuQ0MOEAQtvqXratNwqrbQdOpxMe
mPnbh3n6jRBlCk8p4lPvoz5i9MujZ7gvrjH4y49ZjR4t/tthm3tMbJg/RKNCcUeJ
FFtgWtHV6Lx/M8/lALCCCos60/tbIVAduu/mEUGCFEuCG47MOJbxGO2VA9JjnOk5
+mjZGCuLGAqszs9t5Fkh743j4N/JsZwdGtzUvY+Ngtkafn7CtuVxC6cXR6gMOQeq
Jg498ilYwDaGdImwgbZyPQBvwE1ycN7tSPNeJK1hOB2AYC/frQ4iW2TiZ5gN1vUG
MCQOZ+djBEvWNZvV9QxNibnjAXmzdQL6MlHximSEQGD24CPuOteiY9sl0fKEzLQf
ujlmKvJ7UcajtD5rRLFqotUFQIQczurKyKocE7e1jkvwx+K3mZgRigiWkLRvBEW8
Do95XUTpVxuPoB6REnndVVkN9PfeyvpfyOXNWdW/gjMV0J0v1w31iS5QlExB4Z7a
vbnZdWFKeIrTEcKrQ64O1apGKi8eCKDseWvDoffHxWqagdy7MkOWoKril2R8hWNr
Rj8zIbWkarTploKnm7gQegRfmJl1jjC6NtxqORKTTcaih/W/RO26RQwENsYbYKeD
EWrBJn6+R9DdpYnpWBeBrn3yatcGlvsE3jzJJqLuzHO7BhBSajs5LPL2gQMGJT16
PeR30n+yRy3H94FsqQGX74Tgq2PskP3PR8/QwTAVCog/mrG89SlhFn6G/kbiIBsL
K/fm6AKjN8VYAwwwtWGEQqdzRur8R2daH2/jQtWTBMyrdZYcN7iG3TqAfmrEfybI
NA2Wc7XQG1SjGHfMPM/BkurNtVt0WdEmMTwNABCN1XMmQGrnCiQC99Hk9zCrYmPj
JbxZ5UATnlzOC2Q4QK3pm4NMI8/99TCr3ZQxjuqQn9E1ig5OWr1wOodWHHK/4Q+S
V7kt8UTznJfau3pwQpC6jf+69LUkNJB0zqE2TO4V77YPbezSvky/d694fYN56hp7
OFtFN49hqzbzTgnNaZrPSOymMN8gwCOJm4nSPrpszzUoymPMJtBe8kKzLs6l/JmR
0Sg/3tQDKZYFGDTLJTvDJ3fLRD1OAeRp68RuJCtLPt+rU1l2NbRkySsCITtrQYE7
`protect END_PROTECTED
