`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EL5jh/tO+X5PpJVlJYrGVCm0nIr9jstI1cbkxG2l1kJSjpWUOL11t73yxawLZyCL
5gGU/88ZjArJFbs/ywvGq9CpsmqF733Eoh0YV/EVSaHIzqRHx1JnpeIewoPd+ZzN
A8f6D42LpquDH3gW9CUi41cseDbj2wHBBiXwuHPFbJbtNjLhr4bE7A1QpIPijVvM
MewnG4EXm7sEBUmHpshXW60Ehv+/2PXjte8Bkc4lzE3qURxjhCPqz4d6pcwKCi9N
ld8xnXxx8y6CsopDQcM+zyPeH6aiGFaqeoREf9SEyfiZOuVinGrnsxqCVFEzwrY8
`protect END_PROTECTED
