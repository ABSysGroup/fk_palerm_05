`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T8ATUwSybdGW1qzWCK6PG6huyBo/XvG2nChsvUkvHt3It58GtlI/i+VILDvD6ZN8
as1nG3bHF84ZkFfGHAFtNMJ1JBZyFdzgO9AK/1cQ7krAYCwgRmD1pO6RNNdqEVQY
TGSFObFHc/XBFKWhCOPxjnuWF1RcgMLRzBrThjiH4NdOojbvsQxL5vsbqIEOZksu
N/jKE8d09F9kt1TjbGwb1vH5Wd4pWU7e9STmfanqj2Y08Ynx+kPIRG6fdnue1r1Z
u94Rt9QibIpm2tXAWnN4ZPVQtUcuSRn/izNDIiohXOf/aSnKlcL8g4JP2aNQhbjN
MxPU34Z5ylS81RrxSF/UF1dTVGqUhxvIvCrlLGYGITY571+OdSPKKHJIJgkoZ/4r
AtAKn0f1zn86TO8g6M0xS+YfC4vwahA4dfmYz1ffsYkLTvhVmMGYou00ZIlDby2S
MvsdQi+HhQ1erlh0ZOi6SCI4m/tJjwCJ43hjzx8Idn8DE6QVytZr9dm+kFQE60wL
yGp6+WJCJ1xbZNK6XGwjohbiJYSaNN5F4xW02g6tqULUUV0N8c/eCWDMLllKeV23
nqmqzf7sv5yiD36jdscceUNGNqSXIfhDP+G6bXzybVHZtMxS/VfQS9H5gaAIRkrZ
i9pMurtnohIEJnwiTo77QyxzgEBvSW8zglBVyMtzdMmnX06Dq+0IjDU8dUNSzTi+
NTI0ww//hX3VvjsvcdJKbQCvQdfBRdeJzLIyUUZYXG5YxsRLzcH428tujxCmDnHP
FzzoiKyLugrl1gnNnDJjgZb8W8JP/tjOe6pIMqsAbKQPchZ1rK4oMCyCSmIYx8et
vgbhvSu6+fBtibd8NrWnYhf172FRs9PJokzPFj75GeeuRpPytpHhJ5fXRt0DFCY/
Aw4G4srigfpYG1cximo9POfwVwbQUKporm3dhWvdnhAGzS9b6dTpTydYN3z0DsdH
U8jhNIOhMg5pwZAYlPLfXk4qSLxD3jXs0cPVRoIzMHioNgdWOEfqapKW2T0+w6jk
sLN1dW4GSkptXTXLRyCemKrgMXhZ33Hyj+qVqrt1vWDTozokwvMAQMgV9YbTEbb5
V2gN3o9GC76egpr3ZlGTEj8NhHL+hqN0lrF+4QIhIr+lgGobiIzLkzLWW8VmbTDw
5kz0h+hhVh+qlDgNAhpgD7mAluXSwmLV28bjr2xWwzuzyzrdOz7lcmFIBzeyK24f
r78yZDXQACbz/NF67QjhTx1CxeHGkMJYuNjU4XgPwE59TeEospHoL99A9Iyc/dUx
ND5x+uhT7A5DYsGXiGQlXytcu/WUZuo5pypkBjs5b4dmx+Xf4st+MteAggXKrnze
FWma/CLFqn0hWUELG3Cb3rXzWqTicqs/ycoaysoKYXwH98dCh2+aV5WL6OQy9NRm
ea+l9wayOvEqQQdbBZ/41Q9RirMCnIc5gtHKv2qmZDpBx8aR8u9I15AOFzw2IEMW
ut70eCSqR7u0I2IEvULsUuCwKLOC9vB15iljbzFFXsDsqEmlCZAdDte1JRN2wzOO
v55jHkse7dhAFKzQ5CwJbheu8meV4/TDLwk9ONC2yqguEifxvTVS9MGUqN6RwKE6
CfiU6I+gm2D7u5kIE04o+KCpiTInix7EgzILMLqcyx+K2wa+Kyy0B5NWImllcx91
lXIXiGqLiJTALj+tq2fS059zkCAXXjMpNwIyKSDvE+5+pLEv+LkLVyrsVZ1YpEJi
0VS+E0DBiQsE5zPbDy8BC7QjFFBAjqD/4RviBn9POBsmtVykwFpqXBbvHcOA2Ub9
CTKx20Mjf91NbG9m33+UmaXZ4iZeMx1/35GruGYQIOEMP3cm5gfDu9iTefpz6B9L
oNl6kLxQbh4CDKcLTGjbsWQIsVS/7OcTQ9hBw4rtq8hXt5GYx4ZwPeOCg0edMGYJ
xHFvY5KgiMcxQSB2+uBEBSUYNT9d4AsWDhwf0FE2MtQsVZqLM02ZljGgI6/vW2gW
S8kStiGK0wF5HyDyC8a0GosC5C40F5v4NtFHRDIhTdWnQsvBaXvbqyUubSSroS4M
EUubyDFPDFGViuSZNR7exneFQaUtgplSHgnftdsg+PfQhbfUq5owKyN14aTVzL+0
si064ttwn8or+8IV6vcng6qT4fndumyVQdaPIoRPcDezAdNre2+DBpwUYxyZ69d2
85hRZLnKd0G6nLe2SWwhFwRvv0NGRGSwh2TCnVpKeO0/1kWkRNPEcXWPAXMBXQvX
JXy2UYuXhR/+85Om1/ZmUuuX0ZYpyXVjFe4k6unKGV+YqEPXJILX//irJMjXgGbx
ggDQCOQ/D8rG6bJjosbqbOhClGtyKwH2X1LqT07xxuQVEfr8SQFOoYf8btfUde7W
IiQtfoKWKVxovIoYerNqcxWwiriFCPDzGQZWZf6Eiwaa3EjPs4rU08UZo8AAzLSX
KGie7nhCCOf44iT9PxgCeYzMAZ35x2szg82aPsY6LVPMPbrdOAGsBCAuwFq3zZdO
TWvbLbEcHR79EWaJuvpoX3d/NNHdS8M7gBaM+/LcGgk=
`protect END_PROTECTED
