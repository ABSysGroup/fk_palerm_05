`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IzwrKekYPl7meN7OgCfF8gf6HucbiuFKlkj7jo+BbDs4tKyVEP+m8BkIg7c60LTf
XF66bN6di+AOwxK5nubPs6hOls+KoptYcae3ujEN8JEfOtDQnsZImZn6/Hs9nbKj
DDT5x08PxoocpGaJHPbDkr+eY4X2JgMpWGkpZGr81GQ2TGZvoGkbfn9jeZNVk04b
cIELiecfYPN3ddjt5JR66+ok2PnafhhjuQNry4i0EGRKPTgP1s9F81P6KMfl7gqm
zPyebN0fRCC/f/F3yPEIdqYzhXy/6zQJjTDFpxSK2DOYGZMf68GBiPsHNhnsc85A
PDAqLEmG3WJm+Rk+rOJfJmhvt8oG5zM5mlrNPKQiaWvvWvbm+Zub9MrgJ6hM0WIy
cvfSJ0Wr8PPBI10wNVF3bX+GTF2nccIkg/4kd1A26fAN2dMadqqo2Ni+clx+nDB6
T4GdBey7knbaNgX9gMRXKAKMD+fnaV5NNkgr8IGRMfodNJSYJLKqMgvMolTNESuS
vI5vlDyMW9VHvPRPEP5SkFHMoANLqkIN+TD5Wg1Xi5VUksVnJYYbSEFXkiupL+DC
Uad7OlS4+TEaf2sus+UC3h75PfpRKzQWUtzFSaMjVtdWcR9LIkhxDE11bZApVyGb
uz5fa5RGx5zcXAZpFCYrkbrt92+3kgKvcin1CXPu+30wO8cTakkuvo71zdNpT+hE
pNSwmnoDpYeLCaItQ6J+UYewnksIeiBe/FtPrqjwijzKZMpho9s3bF8iSayGrA4N
rzWSuwaqoSxeEYlfD1xbE/46vDDxXlfC+d1AtPW91vbFAC+EHGlSB+z0hNd6himi
Wu5KH+9C3C/Eyut3b/Tq7VYuDpJijAfchcdkCtzRgudI2NCkExKh87/D/Dpz2iUh
3ZOFUcX9YFtlBdj4I1vQfZMtGHSWYt1XkKhdZpjnRCH+Q8pgR7NzKlMxiswVkF8n
yE+1Nn1HXoL9ovzs1cvnM4Bbc661SuZA+oSsmta6UefHefwq/MaHLBpYKJj7Wm5U
c9MY6p6k/7MiiP4EtQ8jDODa7QRBKyjTcO9z10dB11WOZyYQGLwup8Qbo8WbnECZ
4mY2YyDSD2jIIT7229k4O2U6HQCs7EdBt4GROo8mKrcmSEuRAq6v37iBYmvkitFL
+1R1YOvvv5kGIbl3VKOtZGAAAiLQqIm7cJL/lkn5A6qb5gcNDrMHcLxiV3O7khsb
7it37CW6nS7NwCrh7i7Q4TMVuk73Pawa+wOD07+rppSuim3kQMZjUACjuWzmnIRH
IQ6D1DWiVeahCtRoQP/pMdmT/tPd35Zx9IeMQo3QF6d4QbtKz1fewM967kC3D26l
HvUk/SAbLyOI5gcnVzFPCSGsVWDCueLJoerBMY71HMp428JkXw8QwHFtHl+zxN3C
kCNuxi4C3CmSX1RL3atq2GWOtuCNsdOqJSG3aOB7c1OrMeSb5CDV8S1d+Qm4/PSn
Uv5Z92ZiRZmSEFmqZNqE9cP/wGrm7QEx5aiWRkEdrcmTxFIzJ4QaNA5uj+Bc0Bcs
An6LPCl5x1d5qWG4WSiF2Bd6d/R+XSgW13M9Iy5k5BL/siR9VP2x9kIoT9rfuTrY
xdTSOFt6U+axqzw9Bq+cjiTqFntJEkfOnDFIJ0U+ec3V8GLTWvY14GrFsMrawfi4
mVAyveIiwPjk9SH+9mRSktpZ8Ncm/yMWKXwfTBlarjWhJqio/9p+OwGUrViLhaV2
me6H1H9U/Wq1JEwTRCACzfQhG+0tHnCoKjAVLMirXCueExWqGWJbmLmDNoGqzt8+
wv3hOLn1dtAWiSs8Ml0gKgr9XFyWDc0eSqxMcd3g3GvLGjpGW2Hdsn2C8W0eVzxF
JkXByHK5tvo0ffqMLgRfWHPY4Dn5Oz72Dn+f3TTebMuiv4frQAm1aeZqXLpYeqLY
DNoEiXMbgrOsa5LE9yB4gq/y4XtXJ4sViKANfDLu6onEirisqtgNt9GMsq3UdthU
sUK90ssSa+BI2rT46iKbs9SnGMa0SyUVp4v0Zusmr4PUoE/0OSFVdq6OlJyFlw4Y
SS6Yrz2mBypGJHhiBySRheOzNsCZ0LyZ+/2WSDcLM/r2EMq/WltpgIZHvLUuIpvD
r7wSoXyctXfCQQsybGWve3NHiNL9uq/3z0uVl4JF4B9mCZDozSwicyniCQ2YA3xb
s5fpYfKHy/3dwQsDL/Sadw4SnVEwv3ETOPx9D5twcyIFka+w0GcWHs0BDgl3Be9y
2VwrEwVXk+42YfgveEgC0Hom5XFBcGt5BE/dfxiD9TZJtyTLsQeDzc+XGELkX/XW
tyiQUCIdVn67xmHsrm3NYly6WD5noeb1Y6SiVkVd5U5E2bB9ytrNf/ZoQhEa/GpL
8ooHP3SaiDH49G8HbcwVCDd3Hn4yWIkM1glEb9NgmvYpqWAQwSErg+XKSA1fxu/w
3fBoAzV6xZWvypE3Po6B9D9ajdQDxtLVsJXoEs9+qoG1uABopjrEZp22UHK2EKtN
q83xLtudGdLmcFABnV3kMOBX9tclo0sPyMkr50rx3G3hJOCx+pIA0et8kvtpwuG5
u7iQM/yb6puaoo/kSSZB4NXdMQT9YSPxTyrNBSxOpD98DenL1JPa0BsulPES5mD/
M0paivf8AecwTaMF+iYWoFfES/0gySrIyGUDpGzdNURNVWWa82xNFLt1x216GwTq
QO/eoJptIz9dO92Tse/NNUuoGyrl0Bv39y71UGe5Nsz1ukrZzTIy1BykCmvMyKL7
h/OdiRCl5b9j8i2pSj/VevIpGKCwbXnPs0QBkPZJzeTq03qKJW7LyfLMdSKqHB8e
NuCG7YvQibGr9IGlNaX/dHpqfpYVNVZ/Wj/jc2Yo2Iwj59QlSZ0uOdemydKQ4BIG
jqg6zHxr2Gsc+XkT7MU6GX6KI6EWhGoOsklpExTKwkbJUgG2fmG5JWsNi2iKWlVV
tKsri9hLF4MwjOI/RiMaZ1IqELhXQf8mndmnAKsZmnBPfa8iLz8q3q7laOxsjGqB
CxTsnyNyNi31CB29iPDsEA==
`protect END_PROTECTED
