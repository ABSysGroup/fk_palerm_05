`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z5U/tFwBei679xpLKV/N1Jec3cPj9gaiH+zJF4Mn/xMqdB/UYbTedmnNesxbpbN/
SAily99WZylveBsMx7FXFc/iTb+c6e47EVaCBZ79uFvWuRNJpJcgryWlpUB55lFw
uchUqScDvQABcI1wAnlzu/I3QvFbDOqu8bOLbbra4lrEfy9IBnsTJ82BpKnJw+nW
ylWsnN0kON2m2ynh4EC2hEU15oSdhhaXwRG5mFZt7Yc59gAfGMDoM60tL85F6LdZ
Gcjtj92Zw7B54GlIddYotjYUcDG8mS0zZiwtfN3GLtk=
`protect END_PROTECTED
