`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q+WsR0OgxNUUutS3f8Tkp+LnbnYi+BMprSnaZlnDS3trUKmRaQ6K4FUHB/w6Di1h
08vq/bV2H300sUvc72zwcr2vnUwhgrzvPBDRMDqW5aNdITgqHvOYBevXo5m5zTJu
jFNDvksZwbrr0fu0qEJE6jE+S+XFk2xB2Gcf5A//mR1QZY3KSXWnAiTmtfUBOPFH
s0o3oFPV4CqXhKrCJxGx+j898h5Ro3xAS855NIfbVOMs47klwi0OqAVFanjDpWxj
YIWdvPP5xa0np452lMjbM4ek2jtdjl1IVzeVhiwJ+s7fzur63tt2Yn5F2DfrMMp+
GakIpyv3S+cGIMTF1tr36buQk+Vo15ExktsXwC4TrsSIquPDC51V5KAiB7IIh5Y9
v76AOm5RVXrTYHzzl8qk3L7fpa0oR4oWlqmzSYkAGhh2IdnOMBblAPdW+iDT6BQR
TeAoAk4tzkzIkGlPy0aaD+wjj/Wviahx+ZCf0llZv3gGt0G8GKzLwo+hONiUwX1k
1D/8gZYJMdgtFVWFQ81sFVWqMCqDxWExNYNSCp3lE9a172PwXFfyJ4oWC/4UesHV
5P2iJ6zBQ8LN0fEZvpM1q9wiAUtbwmZgdITRmnJo95KwylfVEpWjXxQU0P61mt3S
4NjVPmSP8sgjtlGSvJ656M+F0o9/l3qKlsM6pEjzlpi7soKdWdoxHhhjXSUgoyYr
nnv5FUHXyYuKOUYNbHdC1/pCbCrRpppdSJ8SdOC+j2ev1sGRIp+ZkVPK7DzvTlmT
pe6TBvOhvQErkEe4aVk07tkO5PDCALw+vPAo0NXByNq9CTAseFJr0d49HAlJ9awc
lOhPFsGp0IwbiZYWP6Qlfg==
`protect END_PROTECTED
