`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
quvWjLTC+CytphYNFleVamYp8+HYTHvqfWBQqx7TVFamcUOfF7qAxrcjX7Addwvs
KThDhQDTirvZKDfgTc6ZVhHey430re3g/6pVMZapOHzZo0MFd9uiOJVGhEBqaoND
RhkQae8397+jaYrhu2D9pAxGtx2+FiK0WKE2qWgFG4DZjwhNOfVjXywcPUOCi6hR
z8FcMP/Ev3wNFLYySCSQewpQagFIR2NWYt0Qfca8Tv+x3MrOHvpowWBmBNEfO4DN
w2YKt7Pn/Hra97jHJA7+3vAQqDdR5XbkR7o7BGHa/9MvA0eGTZp3bRShjF1XPb0b
6Ctw1xBk3gCH1/EvAHlr4UgEhE7qyMBCmLyXvpSY9Eu8W0Id56Q6JpcPPVFvAbSF
WS9LzKWt9NJ5gUXHVeHiNFwd2jKMBReM4GKlyKHSc8rE2cuq08aV55n4m5ST0HG+
nDYgh9GVUdM6Ym+vuYs0/6Vr2+CnDoa71/Ya0z18R5CmbUtqS/ADEonkU/2SmNWQ
XebaeXolEo58CsuJSSVA7WcHZTZ10H9GjfI55tCekyrhi7iRyAMO3MGoJaRYE/xo
jl065MH5QaFHmDJRLviO3YpQc3Y9ftClSvX4/jMXBX9nD3aBq85pkvXTJn0RXRlP
/DLB6sYkNiotR85Cw2/0EBIyzDFhA5pg/XsFgExj3D0=
`protect END_PROTECTED
