`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eq6PnKsClMeycdcUMTqiyaI3L4SPPN61OlY6O8x1omqgpseeoiEKDB1AW5gNosfw
5A9zUzyTPKR1xTj98ZWPLTIR5JXijQx1XsuSLvBcoG2qMOu1ItkR9tCmBxTb7OVV
6CdC1y+6aHdSfKjVVxsSE7HZxQ+aoFUQxEqt8QLABPJmMF8P5y7OfIWHGJ+5Hgzd
K5jnXHzq/o1qcAf2yHoemogztNrqOEskw/LuR2EoSITqA6KoHzWH8uN1lMk1GD0H
wVstzi1/N96tvXYGRNvFFA==
`protect END_PROTECTED
