`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nde9sX1EOUawO9B2k+efkv6azt9CDeFwFfXPhyE9YPq6fupekTxlk/bDaWTFYKRb
hiHNhx3+P3lJgS/cBDx4MWgb6FgVl0BxABz+ypt6oGMEBynmLLij4+PdK55ZNBHN
VuFUZgTA/29yPoIaIAqc0yhtT0fGOToDkoCKhYN6bH3yEUxXTH8PsR/OBJ+Upksj
V4JqIHLOXAqRIXGGEqfn5Z/uB4Umv+MNAxqBWiLN8+qCSHnSMxROsm/aQnJRM9B9
Aqg/h62cC3eDUbwqt3UP/eTrLnb5ilLwArF2mcuMXIieIAqCobQBu9d6OuLRfRue
yzpNWZQn02GomLDivuLGbw0Nb1FfA/aiHq9cIgmMUJk4T20Vnzbry05s0yv1dZS+
FlcMBKYITrFm84lICqm7KIpvlw0q9if510xCHeh0m5xS9VSl78FOy4bAHmtNfWJO
sksbvaTF9lTk8gP8nMtFDg==
`protect END_PROTECTED
