`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NrjSNT3GNYtErQnj4gzTuQz738X684TXhjFrjMruTRFloELp7CFgeWihb+nV1dK/
OfuFaayTjQTcNdqvE1luXAdIGYkmbrNyzPdD5FPFVuP+Y5tD3D5yH1KpU7V8TGkU
0zd5b63PYEjCuk9mF/NfJ3QxciP2vS9P6GqWVdDOMXC4ueNIdZaQhU0mn+bJAXzy
oZNSbLjR6rG0ilu1LIPC0nivZmVgjujN81SuQUDbPbfvAM5q7ZyYTwBf+8awIkif
5ww0CSF2UKFfSUdIG/ed2Woev+xXq37GDhlTLg107ea+hQbedMSYp6FNwjGrCnBQ
PlV5Qv30QXZvnLYt3s8d1cRtl6TIrXphM4YGhfv5cpMJOmOAbtbUy0cm5Gdd6K9J
3fA30zEBWNi1X190tLx6KKs1cg3DeXQuHmnIQFRiJQm2IkIQO0VgMScWgN6ricwE
sP9Zxl0H+7oglwAqw4OZM72cxQjTWOMgm2d3o/V8pZVfETOTt4iPQrGkuSUwMBWH
L2bFv6PBRxv4uC7sX1Bx8ZHSBjwaFkhAJfzAltyVEilBfHi6Wc8VMDqoIyJ+KMof
HhLp+KwTfEjTiB1f6AfmXheKXrnSIW+r1/vzI27UOB4cYqechh4SdfBHHodnbihW
TtEFeq6xHgPBTgQD3RTRnQ==
`protect END_PROTECTED
