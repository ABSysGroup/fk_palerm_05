`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/bqrsnRLZU2t1bqb9RB2iBEQtTI7QHO3DZ8ghwyg8sH3CbTTQXkT4Ft7oquji8zB
bXs+Zb37T555zvTdksx100DdH/T0vYsQwL6sQWpOp7S0f1DhkKAI/Nog17adDb7m
IYM5nB/wh9EFBqRQ+5BuCr9FI5i17llcApvac3v4QY7WZ0O9a69uRSUFqY0V78wh
UrBT/XFhn2OaD8d668zIBzElJslO6dmP7Aq/ZCSsFqDb5CueyL3lT4Xc7SBRbR24
G+Z83wFOFvLJpOywVG0L/Q62hHEicvwBdz0RAVXDkL3bqzkFdH8XiyzJ6D729854
gMY2I8TfkEf8voEGJvu8lLdDvjqneeCLd2y6eJwcbwtY3nEzLv4rpidhivsrIfY+
B6DUw1eDAoWyK2R0zrfIaKDCSzg5irDy5eS6FHJw+/l0Es0hQBobGBI/pf5HkmMC
0Bjpv42alwRC9jLLloSJGKLbGIvTvPmPmj+Ro78n52ET7sL/vcuR0XxYywxs03Ok
od6heQ+qLe95elomL1l1Q5+hKKLckimNGfJCEHjyijfNH5cZoUYnC/6fUBD1Z9Ds
ReRFUb86dDH1PSM1+1wbB/24LjyZAmBu/on67ZEKc2ZbkmfuMk/iNFcNyrs1MqLv
GXZSBDFEVge5qQoGjSopX3mcHufYWey7VcHZq4J2QfTAJfG5tbeWcnlGKaLJLAtL
SLBxL19yx8B1kLET85rqfYuVnjRTSwaWEsh69yvjwsMo3r67XAA8NRvypf6H+Il+
Wl+2G9Vi4UwHdtCmGezKA+iMaIeP6Y6aT0AISSM3jCmwuQWwVOOBM+Fq5TgkZghf
CyCTvlhSf5QhXo5pb7dush68NhtXnl7h9E8fg9n5QLOV984DUuP6qVBfvWdCyWEG
tR+ZGn6EXrghO2QSyo6TbpNZ54S7WZRgH9hZ+QhS6Zk5MhYRSdOI9ZmVwD771vWQ
jHyH4w0vewikWzq0eiz8NHCQlUzDulCikauuYM+savT253Fjz1xYSN4hEkIC1D9C
KNZ9PhgAmAWbVsntU4gpNcck+MtD4WBKHATtdDAHe2RLPO5WezlNwVRF9IpABABt
KqQBJN84Er2XFqFVYfZBtYLwyRfsf/vw5g+RY8woOEI+hiELd/rtTWgwUgyDKY3o
NctaBWbek4w1e5o2ofJ7ZG2K293AMvM2/O+guM++Kn8UZMB8rHTWWDtB5OdInj33
u07IgUiO4YZZd60xJlX3RghvOiQIdfkx7BzV5YDWrhcbl0dpmntBn/HOebtI0EbB
LGI8EnRrJJxGF+HoAh1LA9SAA35W8+EoLH2OF0SH0hzaSbUErDiQWhsGUC0qVCp9
2sRdvsHrQ4/LNTaSAiqRT+JVaxTUbmIJRVdwUPjwYvsP0d/WwW2d0obpxxHpdxIM
2K48adQvrml2flMfsx+ItDgA/EW/6yDh7zXh/etAP1PQRWPTtQh4yxz/zwQGeozO
QbFx7bbuE/01cAE9+s/S/ukqJaFrv00nqT1g4Pveqd4xeEC2Q/gITSvYfba1ZoWF
eTremkclOobOCh5Zfa7F2/WL7JIHv1a79R4iZ+vEuge7OQkhFVtn+2xPaAtOzeA1
Y7zR+j0IB38KkDi6j9xpn0NkMhx33d6c7tugnzH/RHEXeCt2QdnrFzL3VI6O4ppU
P56HNwGbYPaScJGCed1mCkunbGz7629lus5c8GujoPG/62b/CXEspIcsdMn8tFpe
T3AudqQpzipyWQjDwfnuws5P+hvEGx2h6kTirUhw6G0PCjg+1nOdnWPgm/blR41l
mar9xpvs5pdf8Q1EptbMfN5GULuHMD+AHgVjMR7sdCSOtbx/lqO5lVDBdeZsku8Z
3vgjUqoyw5Lx0qurDegMGwOO21UwxMuuutzv06B0mdC2OirscZqwre1uXbkHibq2
DnKuOTg2r7anCIVcG6DjvP6wbs+4dCPiMyTwFQ/5rN7pP2LXWJ4yF53ALDy2VdPi
05UYEAyd9eNSJdEERAaXi3eNKemNtGko7+ps/BsOXMQecLsxFTSi4ioWSKrQyIpc
LmQB78iknPetvsVYgUbAQpYfvBTA1lLIkd9nAqIH3bqK9Qz37LpAqyxkXl6iQFBv
TXiIRvg0SDa0hXW30hScKfSCG+FWevBj0Yv/nhbn+uzgs7NIme+uMrc6uhAOtZK0
hYEoeHqVqu2HbQvSpCsgdCVs3URB7jh9vPPnsv1QUq8/meIZCq8op/TPN4l7fZRT
vBqohxXeWw2hbQLMQWDXg/J7Ss4gQ5WA4aCblDvLbhDm3dp6bGVukZTFvhg+JmAT
pA5gDE1nksj+d9717nGoAn9XilpO/aPPUIyL2o1w7te6Gk4Y/H/0+nFxyooWuEts
wwMoD9yK0fTLvLZWgFvWyuqDsskjQ+BQgVO4T+exKY3bXYAODQFXF/7KuZFjH8o9
0wUHHA5rCE1RJfuq4hLuXEIl46lO+6sVGqbFKmlA8XLBNK6J8/wGwWm+KL5Wil+g
QHC7PlUphiAqAT+cK/i9T5LTJsM3VyaUk7NXRQYcki/9ldlmeswWkwL7aXV7CkdC
zA6TkSEK5toYMAX1IIgDf+MEVLe87HOQBed95CMazNU=
`protect END_PROTECTED
