`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IpToOKGIPHlvmG+PKss6Y95okjJZLvmwhaXfu14rpwsxhnN/jfrOrhQuZNzaBGSq
/Kd7nHm4On+iY0Lv9/UkO6fLC1k95VFY1XV5NoaDoDI8f09XBhPNtYjioi8xiup+
wE8qHm0BFL5FVH2TSf1x1+BYRtqJgBWlT4Jtks9XUHGzbJxmXjE5j4rDzSW3YAg4
h3OFB9VJbhFpyK9Eypz97oIMICt8OCjMQeZ0mekIpD9MGeEmB3+IVxhNcQFDlS6R
C5chWe0lyfp2/MT8IuhU5FZVP6UeY1QKLjboy5JI90oM3IUu6zr9HcnI/Mce6PnV
Wsg86Zg0Y24nZ/gGxanwg1fbjVmOuxoe2qmehlZk6BrUwB4pAd/bGhF8uwRGI3NF
JJYPksbOphbvYrHsAs2sCxNaL4K1/umap/axsk7nlOof/JT4+SM+VEgLW3gEmhfu
EVG1o/XRswuZUWnbYgbWAU4VCNs1G4Oyb3wQnoIhxnM9c+XALCaMhnr2vQxa/F9H
96QoJh6Ar8TBCoT9tchzbkm8QJRyp9+4DmL4nxjyh9nfXfutN33O8Nh448kUzV/1
pV73SyIjTYhedntjzPfDSN3QZZ74R5MDVhU7mJ7LCSGFgQ6gtAbX//+wyPlr+IaA
ZNLfTnk5I9uknVGd3BYuKusco9Klub+GbWC7hpHa4KfwTCU6Q6tHxBSf/YBRkqjs
55a3hX3M8w5AEDr3Zmf0oboRicH8yXknxn3RFwa0BLMtlxG/tJ3Jxs4UFeBmrSPH
FawL4OBQJVfkIqag4ZY7eXusyBhKvR/++ytURuIuvn/EnnPHs1CmG57ekI2ojXTe
D5gutnF6AqMZab50RtXK/UQJ6M75dmm+t5RwqNFdwTCiZR0Q4h8Ut2/lk8miDFV6
T1J4cIhW7sGfwaJpAi+bsw8tGGBdkDQD2P9BizD5iWqBPB6vliUf4SJoeQ7oEGAS
GM6v8YvMdbq5tEkmekkevvNJ0GCyvzy2xEJ6pyTJ0OaDgqc/0ScX4JVM6Rq3kDzh
ClWaAnLRUJn4Ltnc1/G72cBC6yE3Q7JL81XPYjgJRmTabqmpWWjoIWrguaJowyK/
opHpi4SLMH2k/G3Nib26bFpebOHVmai+WDd2qjJ2Bnzj4aUH+v5UAQDop7FyuL0O
IETPLRlRLjimE2YMUOmJ5FFkzjGkr+crYmFGo/gUnLYZOghJf+TNQ3K6RMXFmkh4
bpwhSM6BzDVpwu53qM0FObKABsafclur9lxawUk9ThPnO+MVNYy5xB3F64dOgxYE
wr+U/CbeHao2W/ShomFUbh57o3SCgIa8IApEuPVxhYNz8zlOpbXD14mjvxmlX16X
0kdx7t7flbKzV38DChmWoSS/pK52EKeZ5W3KslFIXIjf8c6RaCIIXt8qvDug7Ucb
nYqt+GaIy6+T/mexhJd0LwzEvduvuapz7lcZtn7lik/NitmcA0Ki+dqKO34F/le+
YpS+IZC47Zuz/ulYIFcLmrP0plB+c34GVxfg/g+LqZbDOJ0GcVUY7Iu3xA9rz2wY
O5MamNPy9IsfeC4ylqdgiW5j71pmyOXR8Up/l3Sgh8O+4k0gLLlUA1HjlQAVb7ZF
Th07CKozFNgoPUtBvL9xG0jruUwpGKnEpcNLS/OG5lbCcQ3avjiVqs1tUo3iA7Jr
B43T5VPah81ULIUZg1whkxN8DZic59MU6xXSlpQOIW7OU9xkpwAPXCSEQgVpjS1l
sqQO2l6+0GP6UElXmu2nGQIZ9UrxEcABYV3wqXPhaVSktpE45AG3zfQLvkmGMuK1
PIv4f7n4PeOmFEyUskJVeMrQsMcFxP6oLJV/wSwCDNOWLZrEIWrZsD64DVZmWeJJ
y/8riyVEbYAi0qFR0T6SgcYIBbR7Hl15GKDrm9v/tsSDzb6RIEjcijx1xq7j/9eS
yqLsB3kBSQL3dl/oOXXTchyIsbYMueZcgfG6DjXJficgYb9OgrdmfU7c13QvtJw/
spvcYgh0mgAxIir7Z3aa/GnB1hhQQV5sB3keovlqeOuwAYWMl2ytIlNuhKtTn6Iz
kvLxkuMU99KzBLTdd31XKH3h2Q6kmNBCPugWTQ1XJtGe8RBL7OsywqO9XoBlHN29
gxDQbdktuUUtHYI2E98E+HSpFWjA4F+yca3PTXy1sv5K/1bJHnU2QtxWSlUaQK1O
DlmfdATFnYKcq+mED2kUpJezEbzR8Mi/VquwmWsGWQqTiUK2dQPOx1RL3/DRyHWO
Sbq/eY8oPUxRe8rjANWhS0damJZ4F6yqum4m4+p2+dn1Zr1ONMosP0Y1e3q9LAu3
`protect END_PROTECTED
