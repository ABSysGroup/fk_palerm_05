`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uuIwwOjqXbH8Qvb01J3kXN8cvQg/l3FuV6+2cWa11nLFkrdjsf0Vt3PJu6E+v/xH
qRzjf3dciPfm1nispS+9whO2PnH02+hQ9emBrOoj8y5DUqBCJWzzLEqoKbt+JEGe
DQ6ANIAguXtoflOKhoBSLBWUf2S34zZ9vE8mJfJQ/gPB0L28eSXQEo5mJO/7oDjM
chKez9Opf8q6HB5c1BsKAlfeYCs4fNjrWy440n/cOzbjaTg7tllTe881vmn9H3ML
aiX2cnDTNKDtk/pBrtbQP9+ND8obcf6RuyDT48bPOI8MIYOlsjmbFdLhokV97y6/
taP51UASuJ/6Tkw4E8cKR2nPLkKPfYGZyQdtDeupkD05HIqyb7LYorNkXXL9LMSJ
KmRod8fL71A+u2vvN6m+wg9Jn3UjkIaBP+rnc+SC3fZJI8IeXjhxqsyxI6g0ICU3
dxeWBGEDjvmjgjuPNjyEzl+wXXz3czzOX9z847diGv7aPKGmFpAfxlWfXzD/83DQ
8DOP1Eim+IAPuLHLJMDNubJ6xnwm4syAgUqXmEOwBsIX/gh57DUw6PGQJSBw7uCj
M3+whmYeWe9UmoIgnsf5eY5mz0CkLG2KFRKKo1r502BDpMHNK7dBc/ZKOzFQqq89
OCnEQpZf/kJCDKG2Jujabw==
`protect END_PROTECTED
