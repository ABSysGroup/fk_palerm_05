`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u0gnOEYT525hwiv2kJom8txFrnNQB/XPu+eCqG2KD+RjcPtZJhIeL/7jnIHH4VXa
4gQEcucnqHxjfYpHoDmhz8vBnPxOpPPIRF6MVf3MnHXY85c8AvAwEer+6MGGF70h
h6BCFN/vzpIuxh/iFSCYG5fBaZWv8jJyRRlsXa+0zxyOWc8YF8qK2Z+LULxCcO1e
JIJeRmiVoa1kwH6b/RzZmxgbLtRR6R3jmgHchYvQ19eb07abdFOMdTn9OIh6dE+g
xg3wVyI/0IFUjCVBvyZT1u7CA6IVmZZyBcDgvgeeMhwiGY3WTylrRw1LLqHr52Ij
Q+72It0iuX9au4EfpQqnoX4hSt8Bvx1pxzzr1fgUkKHRJdiShy8NPR76P0QhbCWp
ihha218xp90k+2SSM97d7U/SCav/7YQa9TKvHCxzsXeWXoT25K4ysxKjUxdtVgoq
0FriYCuxXiP861V587zBN3ktfqho82bEpW9t6J443l2yLUNZB3rvIgzwb7WLLuo6
pvEnYOPJE82b+nIkhIYed2uzuqtdloMl6UKm3nlsm/1i4uw/LpYkpw1CvEFfOv92
46o3SboJ+X+tc0r4KNZJQwUB4AorwN7Pf1XpNK1zaCZncYYsLwEEOM5qPzdGZav+
B7uuagrwcFklhyD7T/+bg488altqGXIoMiYQpcXsQY+4CRBe6xKLogf3ZCcaxqjt
+1j6UI1q+Gmo7eJkTWfs3r7gGhrRaQKamz63M9avWHMAaVsYVOeHR7dFs9x4/Cwj
MRy2mumXS7vXpPwyrAKVxVd9R6EosCWj1JlV2zyY3lQvp51RRx/fgnS+WEt/dMR0
noHreXH8rnZ8pn67Ulg+BvJXIFMZByUT1d0xeBhIRHRDWoj0+o9NQ1COqnqw1s4W
qfb9pfsq6sqxkUQVulhtbvF8E0e+CA+urgBtJVq29iJe0jnOq92Zd7+NOTiekwr8
OeHKfmKHN8Mpx6IYcqgDhltg63bAUsr4lB7tZYRkrYgLrO1QyIb6BksnnAKKMTV7
LL7k09PYkYCWLRxp2GOfB0KA3G0qDSHd2PWCCNrqza9feYwt/OfPP+6D6h5Ps6a1
zm0GoXBKmJQUXIpfH3xgqr2jBFrS1KFMjBxyrMu5pebjEtsMS0IA/4vFhUcuPD7x
s6WN5mqXGiuzpHlkBqiPvGcY0WBzwXAU+S3IUBOOXydYE/3pnmsE3MXoZPZiOmTi
OvlaMn+7SGv80+Hl66gUhQ==
`protect END_PROTECTED
