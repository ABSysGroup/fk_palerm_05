`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
liZamKOik41ECeovIq1AiEtWRtb7bwKwWraliupEhzofH0rzffz+RfMqaLTQ8kQk
nbuMcDW0gyb0f1jVXIHHLVyi2XYioY3j4sDS+UoLR9OTQndiB/5kfd7tx9/Wk0uQ
ovejqkjF3FitFSMJymhuPePfLvc24rueUIX7scNeKvq7eB+PYyl5l8RycQcDSAZY
H4x2sxChB5FPih36ML1iilNCDsYvxFszwQ9GctnLh+l3n2TcBxEihZp28HqhBISa
MWBGBykvFEr1R+IUSC4VFA16bYZhNFYheNY+0aDEfBDO9AO854Una6rRfmKyUDRk
akifxDRvW7Eko8AQQ7jIElCrtISjmPF1Kz4CE8xEjm8WSf55smEhlcsV5fwobEha
boXPh1PY2MhjlpBVWVjqsv5asZdVIPrrAmkcySq64kWzp8+717R2bpJ9YpYihq0v
FLybCvrDgXlaxtj3lNbgnkVBfepWdXZZJqanqzit4b4D9zPGvMGcSIZMFplvNKJr
rdQpj3YYtDkk+wP7BzL/t3NAJpIMMy6nAXdPONKtZTqf4B8bHaX7q/yeVNQNOYE4
r7gUQ/5q3A1UYS5OCDI8yKoVwiKttAqPbPzmos7Ogwq9UlknyfW4BUnAgrBCMtBN
GD/y5+ThR/FOIMhBByO41GlevLOpzXlzpl7RFtya4KG1MM8ykPCzNp+bMiqJ4xAK
e5Bd5KOaiAtAhSEdoscakNREwNi2jE8I4R3IBMXbMKZn4mGBmXK7SlYM0DSs4cbg
t7qxsMsRQQc3hZGabl8J9A0DSxIHPsa4zrJ4PISAFfon+0j4anGSD9gNP2iTT1io
OJsJ89gwcWFXrFBBLPiDhR9mhNsAziqiEV/TjeTHKtH5uFNj0LtcjRoEYwFKaq8v
6Z0zGjFHAhLNu+3dNPQd7ABZLO+v3OBohXIpBqWtWSFZ4uTZwxZqxs6/cupJIqN7
v8C8xX62CQOQVI/lfWrUKgTFI83gXPL6YEjotUoKYTGrg2tlnodky5RiOPPZB91A
SCeHMvlFxk/JLAb95lBV8gnm3xvl8ZlsRaPBANMvlewcsMlqftVqmUaHmsFNDGaF
UO1XbxhboZf5XekUrORcDoox8IlckZg2qTTfo3x8+ackk/bKTkGaLCyENtup0Hpb
irtphTKb7pgwHe0/1zY6k1yoPAXfWj0ttLUrcp0lsAfNFmq6zGRokRYGoiM7AkDs
K6lyXABHUlRwqWsetC8azvgp2M8ENkXOWW5Q9OyVkjxCKUIDKnhPRGZxRQg9J52O
smZaVEqGuCBKWftANMzrMi+duwmI1ogtOKhoanfnnROff8DPivzIaC5zqjIqq2fo
BlwQwx4DMMNVAt3zHfHSUMURAyLWwSzYorZWL60+SD+sjBPc0xbgeW5cGJDNQYlo
XSSTtpMyYIXLyI4wE/UN4s8jMp5sb2lVWKZb0vAZSasFEERvsykduqFQJgnChLek
PLPgDuAGRn+UiqeDxLhvpWAM/1bWYAzGSVXeQ2daqLI+EhO2caAye8E+DSds767v
0qlPRzL71LX4gh4TTw54Ov/s8O2lPBPGnEnugESqwmC3klYNLkp6hKxb7KbljV3h
KoFK/URwVP6AWvcwg0jM+EeHOcQQGgpERnEuNnfrouT6ktxr0lqDZfjDIbfs8TNJ
rEJ//HmUoQSaPt9ytNLfBKtIpJslMoSf7Ieu09zbDAo0dLDuaWWmGLJ/VCgk+GkE
HwHBbIjLZjSz3xDh41LPNaxnJWtpTNcVCq/gRPrawQ7no2yxTedckwAHiOJvR31l
lzLpDOSTV30NU/sNEXqnGIVd0UbyxOxOOttXUoUQlrSHBCKS7CqgBEOJidr3BtOA
1Vw+rXwNqsx33dk0S5J/i4pzc3WMSDykC+JsK0VI1zbh597aacGpSczYELhuC8Wl
ooN7FQ7CwF+xvsPCeBmlvA==
`protect END_PROTECTED
