`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fpGQGY+YVlm5yFuc7Bg8FgfBk8GeRN1OnSBWzEXl6tGK5amluxEqdk6S/Ap+rFQr
izE/eakPycJwlY+sCqQlmrDl76K9cTVHIuWo+dSBvHL43vy2OqB+stHz9ax9VVwW
lvfK9jGM99A1Ymqy0LkbvYPZqLhasYX+rzRJQXR1T5Uo8hOR9UA6qxccydK/5oNL
JIx+NgO2vd347u02GETnABG0cbT4SB4EM/ud/ESYBZsofUko/OieowJKKoqWXznw
Vj6QfPcY3k26AT9OjaPbyA==
`protect END_PROTECTED
