`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
viuKtX462HgRET4WvAZTe/VheJZSXPSO0CySw4VDTNPedxvRsIPejUJSOla+5Sbv
mZ/DgP9PGZtdrDT6jc/aPZUd4UY5pC+WiLwWAKDJS8sxNjLIepIJm6QiztDM+lhU
SSNy18z0qHR0tdcCsrfHMitczfVG3J9idhgvwBO+ijCqe8cJgLWkshaNiMrh12Dl
MKySGx09b99lmY0wfjuZMcfyAkD3Tc0RXB5azTOG9uKTB3+jqkIj5wN45PbAOAnG
TyPAXF13GeZQfAoWpMa9VoUqf1gJD9zeCuTvoBvYxejNnx2oCX92zfUDqgc62jDr
jY+d6t2aUgugnI/g3DxwtALxW1ZIITwU5+7s5273LSE=
`protect END_PROTECTED
