`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9fcu+l3LfpQ/6Srhbsy9A5TDgN7AcTWuzGG8kYV972vU9WJVW9qZcphtjinO8eD
zyU9XWys0qs+cIz8n4P0ffsn/u33/DAV1k2xmfhWwwBi3vfxbn3qBXD699p+Cgrp
Wl0TMgcrU7A1m6uy9+mFrMxFL0M6iQg8FsYJ1D2MaTW/ncdLIdU2otJoT8JnJ3Ws
Tksa0+HD6fzi2M6Icv3mPggc5lKR1OeFcklDoqPK8qhGrP8g4erOu46ZepaV9cE/
qh4KdNaEbzjksnKDrmgZ5qbI/8Xz0cfYwC0mrb111o1r0BiGI/L2HedYkKWUYlHc
WjZl2yLHZCOFjNt3LBvo+A==
`protect END_PROTECTED
