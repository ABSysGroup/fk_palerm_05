`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l0NDvByGXqb0sF9DX+WrzA7vo1DP3Ex6IVW3Q4T3ntMHKuupEsZq6wab1gruAAVb
xp0bFWZyBQDmH8b1hsuytRRhWq6zJbmD0f2m+RJQ5G8wLg7Px85NZM28omCNdqyo
5BU8AnwLSHPsLY+XfqGs/T9A1L6nD7KrqP666wctYkaQsqD3/JYiaot6zt2LIKVS
dglalYY2ot8Al8Hbh0D2dbT47SoGHoStMiNfz67Hvqj361wMwsKKYFpEPJR6GcKp
bfEgir1i5so5CwHyQb4qhFSS0M4fLOVNL0YnH5Rgx4w=
`protect END_PROTECTED
