`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2dfGU0sBDqJ3U6uEVRRMG5UodqYIsQtOz9FxtcfnUO2v2QLqEKvq9vWzZKKho6dS
iVUX+RuwH7gxaoNPpBfv04flORqO31eRkPd52FdH7welEYti8LBpxeXn0Horf4xr
WLEs22kirnuNqF3MDZ+ywaCArys00oD6w8W2ECqmbx3LQHiS2/uS8S+s1qXWyUcr
KSQAUCNu25MpC2Ht8nQUL1bDNfoxG353kw/ByurxciuVogepFEydrX5+Nb5j6DlQ
iO3y4apkW5Xd27+Aj9WC+R0gdskPO4oywSYtthUINjzZVxCBTHIWMukS1h0Um56y
hl754NOa+mPAK35WTyd0t++r2h9AEASlcd2L4FO7COdb0FNGTASHmQFO3LhJhSDZ
ubj6tRZJH8MWJbMwzedrDpRAxjU2A2Ty58EehRBImclnM9y+8oWjEx+TcHMK8CnQ
HdW0o2MEMoAULICXZC16W24CYlmrPKVeaHqiloQQgfoC7XdonDFNd5P1ftfNVDvl
c89cB/cSU7J0CO865Rxag85mI+Smb5aD+qeAwtUXc3DrGcxHZwbgxooNTUpUu4lQ
8ch8EAzNbhyPpdV64OmZvOe2I7PPYD9Xjz38LZXelXtMIAR0eESKgfyR8dU83sNM
WuKty6SGHpX4XrX/NPDoJr9o4nMZ5KdqKsON/ImYW8NahZoX7SVDJ6/XtzzXST6k
/56ZYJpKT5d8UBWhxnO8XJATrCh9eO8+uhhQFPkCXnM=
`protect END_PROTECTED
