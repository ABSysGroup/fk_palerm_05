`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+SmR7a1+9ezBRXg06/FvVHHkeFfaVxlJfh9Ygz9tw8rO1ddu+4N9LRMSt5+nwr+H
HexBk12bLVAYYSSNNdA7K3ZQBQCNyPZqUOR6kP/jgTFTut/VcheV4t6SWjULDZ9Z
wEwvonGFQwCWfodHvRUTynaOJzZmfIwgq2Ch5GffNewbjm+gcY8bzQfZ5vaH884X
5lt1P6N5i0qhRLjh2vp+47HKAYgBUg/j/D9Px9W7keNVF+RY5ZgQ0l/faVHnJS/M
xt/z91NYjvzuRyV5RqpcENKXy5slwksB8MU20E7DJ/mtjPXrMKqBRK9xehb1R1F3
8k45v6oOHBtiCl+X/IB+7GYpo8kpIvwRG/wEGy3xdAJRZH4EXKZ55n1olWSlLMO7
ngjnWjzxEeXOlsI4IO5GH/iHMMYXf5dSSyC4Fe3B0ybc1PRYg5gyozbDmiBzaVVz
YFv1SoxjCtEURDN2knWWKV0BWcLlX2Tma8x6F+sqdjbEyqVe2E5POspRv8s9ZT2C
iQ7EtXSBTZZm3VWXmcLM7OMqJX/0VZw91OcHG/N8VXhDBqnkpyOgHHzSaV4OMR6M
ncFaNtowppzcFDLIMFgsSoTUGuq8sc7pvY+vr5QCjxZ9I94+wgmlsKGhIk2Yk3dx
uWyd4Tq5lklIVnRMfsyRbqtIfVPOaL61IoW3jOlDu11nHz6HvsPNPT0kHNPI1xJD
pKLCztzkRLniZyH7/gJ5Qw==
`protect END_PROTECTED
