`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DNyRmxn5vZXOKB1WXVUSsUDJ6lD4NMyi4DnRk+sr3CPZML5oD9LxfeIxbt6B/r4K
TMZOTZKrfw8SM6NaIvY3UJilnGP2fVBrTy5lKLa+eVccMKYLUY2g5mdLDpad7AVb
NFuVIS6C6iwMWUGV8hSIhGfZih9cXeKCMXPBEC/sfmPvjTMKoHyxzl7uXn4oFPIw
UYiOyZhdjYd6g48Bk+9gW3BjF99c2fnCiQdDgNz57/pksJYBTPQmCCVjt/mR5uwp
xeTCP6s0JlzN2AASG+pxQA==
`protect END_PROTECTED
