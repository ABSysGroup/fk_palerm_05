`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xBUk30sEfkagmIkFUIYFcVa85bBz5ILNSzbi1cGZoqpUrRqe+QRmQoZBrUPJtj4r
971/Tez++6d9FqlcPbbNKHWD3q0FfmpQxde6DKNWsKtnXwBWBO86wyJfWFc3b3us
/g0r718cKGi2FEnyluw2K/GqU+mR8/rvAlsrss5weLzbLFfvcoU9eE2ofDsJPtGu
NC+T9/YMGjBfz7LY1cgZQ7/m9stWg1aRJpUBb/1amRGWhGcIDDeHEGcvmgX6CE+1
JlPmv6oucz1ObTMyxLiG2hKln3ijjM/9EdVDbB0hLGyU4iuZ29vTFnFFxlcymxbw
lEJ6B3NPap+xHyevmOXbE4TAn3bwCQsRMrf+2RK33c+9zZ3Vqy5Uh7bLybgyh8M0
HS135NyljUV9IzVJW1k0Q4rSPxX8qm0NkI5+cDizKs97jkV797tIIHCmDHnaI5XW
q/BcW5uvhKRn7vIcSuEkoO0e+ChE5guUq+12hADt1/Amn2CZYGu9KxrqOUg0d/5n
PZVAKo1KirASvp/KJdvFuPo6tTNVdX9aOVg8HXcfbym0vdFNcG+fpZOAxLP417Mq
WeTEWI/Ug7yNm4dnUSxMkXsAWbDb/ZWvTBhU1jfm5gSxbIPmTl4P9LvaYnOshDsk
Bj7eGiANZgriky9ntx3f9ZjwzkY2hN4kfqfoJATakx6oYx8zhyP3Bftf8+cOeEbR
AogBr3Ohae5wlLJWLjIkN3ym9raTYbYd3f5S6Nm5GdTTdL7dXsm08Y9RO3a/hgZL
O7EbXp4tCDytOowXDZw23/bNwBbMyYSs6lP1QmF8g8yhSCD+FPII8F02CiwU9VVM
2yy/yKAOcK1MT5deWXP1nOdQhvrNNFo1HMu5LtfhXPHuGxfXWmr50C9nMBIXa+br
HnFJzJUfMYOmpuZWZfj79xEr73vMw7opQZcHQbUxdki3f9LVChCiLmlje3H6dGey
`protect END_PROTECTED
