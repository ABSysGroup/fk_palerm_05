`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UhPr6TBt+gKxa/O4UYCNXdhYEt/5fqGMzmRNIj9PYbIX23voWRDc69apTNj+rKjU
ORwcg4Or/E+p4puWL/QUhNvsDADaXHq0TASqywmogn4QOsDfbV6tkFkdOk239dor
ij1s5n5g+XjCTlCfX5Mi+N2QQ0uzZdwBLFwCLaiQ/9KmMlsPuhr7WdlfxnJGVSfQ
kj8ipWyps/PPjwMYzAB7bd6X24y7g3pBaN1qJddOKXFlV+hcanZE7RYhms+Ah2v3
V4C4Lh3A2w7k3w8ET85GJu5i8OFC48fhcLtMybMe8Hwjr0OaoNpOxk0IWV5euoLm
0A6wRqOQrWbjgzWaz2B36MYBb5bn3LBhbErgpw7MKcUU9hMFj45NtwTBVuImzc7n
lmAPjiA+ai8HKRUMupdmHRqx1FDecsj9AKb1g10kQ2QqV2q/yX4dwX6E5+IxZMHG
uCEr53FZVa7CUZ745oWqKAQpQEKGDSt5syjOoeC5BDNMDD88Ze6noHSydNQ50ESu
RJWHCOf1vg6jgCKgK7LHhog/m5iHAYS0InMkNRWbnTcAHa13VNkXQr/nQiesJU6j
uXmJNJ8jv3KHPagDAgwIZ6ks9ULaO3xWBIBPMUsBQOU0I5yOuJSl1BYxdmnnEiXK
4noeRkylBi8R2rogT/22qiX9O72yPfnUEF70vxAdoKPFbUc8gA9dVL26yjpv1CZz
xQTmMt5OpNfnLjEu8xZgdCaFWLtdfEWsaKrpDo0aRKH5mpCIUb2yNZSzqFCUFhV+
wCShyG+/mynWne4QrZRZHeQRSfLhm/FOJ654nC3BSWjZmWTsudF/HEYQoht6dg50
OV7EDhT7hZt9iP8GCdfkPlXDvlwJhLJitree1FPOeEYdW6WAOjdZO49dlRIWthqn
DfHYHo7Lw5Ikyaekgmx8VBFahrEdUbpJ3lsdHvSLUcq8KJDizmikLqGYr29PAh7Y
K8D2uUTFTYVtFTw68800yFI7nXNBnyS9MuT8lqowO2lsZPaFaZiywgZTm5lOpuHr
pmdK7sQtOiXfdrsHdwo5aq2qBq9uZLnRJ+1QHvkvr9quE5SAGv3PGBH1+YEXiqnM
BgmiJS5anrnjv0kCYo5occcsaZBpoiH4eMx+xkmgi4aackmHDayVQlRculjN74yF
LUUdgWwwkA9wCOmnNG479UTyFiJ1p/pvyxMXwFPt8gdJHsDB6IDmZLpSXLF9M2oA
CZ4/ApwJjPL/T7RbojwiclvcUFtXXQUFGCJQLxcErianSvIyzyxMu5/kn5M6pj0K
2tt2gSgpwWzg+UsogU4O/rkVFGaBHMlniIPGlAhCLqAXxsjtHnl95hH+kYdUc5UI
Y3GJ4a3d7Gli0jrqSuoyGhgQrypglKAukAGB3hkBUHYPyXDJd8IV7Mnkgi0KNfgo
V+EWeyh/LA0C4NOr1tJOm9rDH0vl6rH/lkUgMiurzOpWyS4YdMoqsha+tBtbtp9/
v6huSaK3oC+2zbDftzHFqegrF6pNYhuH8zCMSrJKni6/QYBB2nCPN+nU4jE4e0yO
xUwqrU4XVL7XWPKqggtGt7BF1z/HV9pGIPu1Tvb5rEnYjYnkVAqqJkuQHyQH/GJC
iQ0RQ9sW+Y2seIc0XvejXTsjp/DPlH2Vvi0U/o3/HSE3HFIKRcX1JwVwhPd836xl
FNjSVshlzMudCrTUVeUnDkMl/MMqFWKU0HPbGabFUZ7hgjFk6jxosKKYDvbc0JMT
V8y/K8BawMjR+IBe2qfsrG4tZAQ9fNhZBOsw5hkExgJNSIIcWo+LToxWZkR/AKtL
Hsn2hHXH1jrAyEyqWaQBd9VurGNvRuV/WQ6rV8V/810yMDDf93zOwa80EedokNXM
uOGiUkjZA2ZLypDYUVT7MS/b6vtjLCl2rGpDx0BQ6puFLF+EzuaDEQ0VGra2JhsS
x1zU5qNFHLMIPmv/CTSu0r1YP29GpCe2CgOllAs9DE+NE2Fqy93owsXUx/SOsQXl
+FX4eaS9hNIOPK4GIBbYSyABccFzQO8l70b+5tGDfgbuQ/fSGHg9S8XSHvu0gUc+
N7AWZob5X+5e4dtwy/XZYAN49bGbFN34mCvMEzXBdsnviYR8vblrcgwkU93XYDwN
AGvnwxcamDi8joa0RTMrGijxsxu1c77gvn5E6H5GBfXpa1KH0Xg9sW1La1qtFGez
rMEiCO5ELn0AUw67e46EAuhCMkgnZnvwRaoyZgA0jQGY2T9n9XaovWpJxR03TJHF
iQbNmsifPNtzvu660diTEtnkkm6esDd2K8SIS/Ia09suZlRxY+rtiKg6DoC+ALx3
7B7H7s3rCFMG8Glybnyy25gsraJQjZEynrcj3d0ZINm+hPhyx/Vb9uYnZIT4g2HS
AsB0FYW7gQOOlU7Cqs6DndHps05gVAN8oEQyIh/sCSAI1V9ahgfWEHgkTyLpDQXl
u+3WN1N1RQTPy9iQDBlpVrpEgyI2vNKJDHrOwvc9ZTVDlVIwGpJ9wt8zaSR86B7l
9HZAD5OP5fZAvuUx7LxxMP6B4IurH7O86wENSWv+xD8Vy360cn/JV5mInfQAKg/M
BWEA30VghsIhtrFg1PHdCmi9wabTBpO3r15M7DK5NxSo2dHnYqkjSmXB1inuCTSr
JQZE+zeDzA5R5/aauIsrAqCRoerfNjxNgPFVDJaQo7duZFhWDqZog9BL4GwP1rPO
kwOg/y+pDcryOyD04gg5cAkTMV0n9+hbWRqsltx9VB8ozSco+Ko65f3XalOTaPZ+
H2Sbxv5IyjhRw8mrLzTqZnyaVIyD1bBAFZo/AaNdxjJKWIptjY249X37AU+HnI3R
DIoqCexE+c9xGvxgNXo/zS2+sivKHCV5c64Eu2tDtEZHgGLRnw9ouXbOMWUlCTT5
JekEqjKfiIzNd0iWlPcn6rnhSL0sfZmtkcBwbWP2Vda3D7Eues0z8IqV+cnGyaag
tHALKAZX7KaOyw5g34+U1xJyE5bcbUC7h8wQg1hSTjrngIRY1gE4zXJEr1Z9bpp0
FT2yz4S+3Utu3d42wBc8OCO1ffmHBn5OrUdHln3oeZ9j3Axgh7EO1athcAOMYMTr
roBQXMPO/v0vb+vNESUoCCEbKqxh/xAu/eBfJxnkbP2XIh5pm/4Chdki63RVZt+w
5Pi7XjZp7aEMHZ+siyzltXomOfiZLkVPMlAUsxcz37igyDWGSjgnvzgA4GLdgbKB
29zjWfCktKic16KdH2S2pZW+EOc3gXHmBLgYCUMWaEZyy/hDfYCLUIoIPyCQHXmx
gO9fZSl8V8FV7G/ESIzwAQP0NoD0h3kjERRlRjsz8laMMwgWjle96Mtr6VRgH0J2
AdDqrnJnXXTyHbkt1TsP0r4mz96uuONpQqufbumOoi/ZZbmYZro1wNiapPWNjHNA
SEHA03OXy8i3fl1iPByMzVIjJK4D0SxBFQSsQ5GqwKUxsyftnUkOKJCCZ5VGzuRt
KWUiAcOi9WUMv/ENW8GMC3VMP/luVVmg0z7GCWxCMN88wJddilyPmdG5qD+0PPnd
Shm3BwSED4qpzAtgEcui0YsiFX/jamOSeYN8CF+3VLi7vhVLVx+3PBoEhVV1Kg0S
Xp0HSSe8y3cunzwOSXSZETBQIxsoKhIiyb5Gk1ICVujrePnqfTOJLJ6io4IYTYbn
QErenx0VG311UVHZlv74h+ktsT100yI+OxzBSTlslSJzdja5jFvdV8a4KjvLgZ0n
sC0ke3ICHc4S62EmtgmekfjRs1lbC/Xqw0KxkHHZc3QnE62W8CchnxeU5gxwyqkY
wIUA9SmMgW+B9GKWF7FAwsR+THSMYo8y3dolNWV4dn0mT15txktgyRJWoYWOBeoP
UGopWj05NXVJzU6yTfQdIP1Q2hImEZeUDudOEtDzUiZ3l/7UvOzDoftXE9EOk3HB
sGXCOUFCHM6aVBpTvpECUGnAGKoOU7yZVn9pnyaRgD8yftpG85H1k16FDtCztvKe
+lUgTM2TUC6giK37x0jA7DyBwjxNf+bon9pYTNiyhDMar/5LuiI8ThiQe7fYv9ui
oxP1lZw3YgIaVT6rZvoyqWaueUGi1NBokKHouMUbi+U6ed8myYEwENBBMx+ydULp
kXiUwGswrx2ZUA73wU6bTjIyb2IzL2Xrc0Ye+xVgJeG+yyCGqKtcoHEMhmhVk8p5
DbsCos3jhFunHzvH3nn86No61ul7gNTIDBDeXWTypWbp5IGwOD/AoUyYRDIo1Cso
Hvjw/18ov+/mqf1l4XxLwEwr4BUj8km4es8NddmsWckC3EmwOb7RlVP/2MLRqiWV
JbMA/uKtEsSsnT1x2reECeG3gYBh5iGVAwBAs1+ozCkM76WIxwyGYcTHyR+lqBFE
tuykozPUtCD9fK98Ye+VmqJQe2jIHM4Y7Ig5kEss1QlXy3u5K9UTnpswBN8ivzxi
zBziNIX2IYwnGd+7wSV7nkUBfq6l/MrdacRzdX2pyi+6SgjjiCHnQdOsZTEIh1en
lVJupfyVmQNBDfR34kqFYcGIhhnX1dF1BRw8BRwfjJFGkPpvsq1EW0V+SCAsB8E9
FfBx7rmQBM3xFBV6Qa75g124JYaLs54aQEs9XXXtInWpG4gGU/OGFYvXU41Si2B/
BU4sGZXKkyVptRp6u/eF1978F+kj+IBRSTn7k0ZJhA8hFsYgUyaaR+XQynxnaMFj
IwAWq4gZO5UUCvMAiYEfYMB4/GesscLmBEi7kyvaO559cKIc+dfZW6LTaYBsYST2
8AU76KnVl2l9hlPEBpdar3//he/bVClLvOWJj4zbN8+RLaZa2JGEZpndZE2aLWtf
yoRhYXm4nRdmpL6eUTB+5Rl47hK3iYZwACV6ehe+gDILAQLypdujx2Imn6hESEFO
t4d7k7s0ucc+8O6uz7bRAGO2n02bIYKzegOGdJ1S70U29DHw+SFredg5tzoZjQqh
/zflWhMkosng6G0kxbPlEoLUEvoblkcmJD2DCJGmQ2AsXIpj+UsU76YED5Wn5vBP
Q269xXjG29WkXtJa8Pzy/QivdqJbUxPAmUtrVTpccpwM2swUktzSKrK4cO7igtzH
O3s13+IemJjoz0h0J9aXDqZZSJoTNCGy22k4uFSxnx/oYzXQpYDuBVnEcgQqg9JB
QMPXaxWYXJQVwz92Bqh6kQi8ien8c6p3LWAjY770ih11RkqGWmLF1K9jdrNj5tQd
iNBStlITwWoHj75qPlVDNXdaIsrXbMWqnaIpg8olclU88+CPf7W41SOOQFEHepN3
2hDAZFCupGh2IYOPxxeimggCf/TzuPkrRzj3cZMqCMB2fW70atKXMuJOOEt5SBe+
xk/V36BjgCB2lmYFnHnKO2wnJkFAzTwwt8RWL9fEpPnXTeQUYFqGjgTDbA0I0B+K
d/d4avaEtENyo7YB6EXrzKeD1jkQaT+N2PieHaYHNJaP/9nLAuPso0QnkbXoQKIm
p28ZyAuvWFKHXzunJ4b4+jqPw9qwpFnPcJSYLNy3iIxRUTlmED5EdrHc8bVB3aiz
RPShH4wmzh/+1zy7mf4MUPawoqiuaX4XCCWjX4u/UiD5a5sv6R1cS0Cg8xntamKd
+zKi1r0EQYR8B2hka8xFhnJ2sqvlKhZ7ha0r0CQOYbPrxOsowEk61QNe3zlUuvJX
TR8guL+ZIbhgo4nH3eNSX3jK1Ywxz2Wrw2nnA+sWHdYp+ZWw0US5nqoP+WM1sgtD
BU1sld281RID8W8wkkCPncrK6UqhwmQ8hLlsP52ZjLwdzzjvnG1dF3P5X+hC8Lci
+Ws54YG5iR9VioGW2OsSXi+ls0Gulfib3sYnuCIbh+qxTIPGBUcF9p7XGXG6Zxlo
jiys5QDvjKLzRl9a1ahJ5A/LapajhAo3JuEmZQKTyj4l7HNX1hYaKUc9N8zbzOId
LjPxk/8WhPUb0u+CZMh0xLyZ+WfbOmw4hBAy6JqeF0wCkcUuLmuj2dEh3BUUsp48
1hJVP2sBJwiCwxGHYr5oi2dk3pBj7nH4BaKGeAMnzKmMXWr6ZNzhy6yQgIfDqFrH
kLARIQEHhFm4CRulCW6cpJjiMtdx7+ETESOEdJ1uY+7KJ1K8uq2lDFqBZg3417RX
yZuoTJ2uNASjapYO58n6DVPMdzdTyfN0lCuEEXvk1kqPEh9aHkPbhm+4Q2Ylof/l
WR/oXvHgbMdj/CqT22jNa+NUPSLaiYMJWHh4t976dJLU7kMuvFLO0y9b19CkhULo
L/JJpxV4v6GDC1/syA4HUJWNtUKl2Aq1xhwoMy+VWZyAowwtsoBxjtUcfY5h5bEu
Z0h55agYJ6r/D1guAV3yFMSkH5fMMKzBFr63KG0Wi/+7la2aYQEQV9hGKkda8HcN
LsqAigC1OufsAvTdfG/dPyu8HUbOA+tW1Mr3zZrlD6RD4JRLsivNN2ZjR3PvUI8B
wf4HZW7NlcnS8CkXfCWolM5zZjo97fy9K4kyBZkkmv9ioZb8E8ouCq/fSAnBLuLm
NaDlTf3QR/ClPMhgAw+v9NwSkW4qwAy0f2iK/nlFLcVrViuSxciqW0nRNAh1nuj3
x4yHgtAiTk5rOAeNPxi0b7YCpS6029ZwZVp5MVRUqPfFoSzhu4nrZSDKNOppyavO
A3NG5uBcav7E5MkbZ3kqx4fAAkra9WNu981nI1rVpkg2jBFjNKBy6A0g5TIl53H2
cDBheC+11VGDy2xrpkJd4yJc2lfpNDbbEFkXRaFPWDHEUSp8M3aZv4EOZAUSeXVQ
ZA2oSXc+1EMBqA+4tjStm14oAYjXkTADFPkYSWyWAkc/Dd1dPwpMD3YwXbbHp4qR
pE4imnrZh/RAQLg7A75m+N6Xclkm8I3CM5lQ2kclMWZV2OVcu4bcICZNVlZ8rThN
k0PdylT4ysS3sY0cY7LDCWTvonXY4tJQnpDH6jHHaP8tUneL/0Nr2xDFgnV7CKNn
ZYgcm31gYRNMtC0JwTLBPgwhJ2cho6HsP5XM/+4EU/5WTJlDLCsYra/TSHmRdN3V
0S4nXgvk9fC4CG3TzbezRkYvez/qTp5ixIIgblzA2I0Yy+cDUFMB5ytgbMHRyiPg
opQcNmJkigC/TjMA+1nSO0GIS7Qp4H1VLkxyEPtWksRG0S6oJGSX9by+xkfDatcf
mio332/gkLzvfcA/TE+D2e0r0ZkAonhal8l67/mgwPkmLPeXn1rbE7pGn2k1Y6/A
Mg0JCwkySzOtD245nD7M8Nc7B3IsYEOeSdcRZTl0fQASa6ipWncXGF81cwLdUBoI
yOr8TPGKV5RZX/2MdTdxYUH+tX4ATMCvBVjZJkKJompjGP0df2j/hta7aWX8tJs4
wV+tEQ4+PMdEf0AsW81u2sy5IlAXeizWosB6B/FUuL507p/AJ0rH//vwgn4YA7po
wLENWDwijhKEPYdcW3tdYE2YB/gHKGUjDdcxOiBGhV6rxgpRCmwsx0yd75MNWOeA
lS2BHOlMK5N5eCKiY1Thu3PuCMejwyhmmN1wi625dKLT6SRGcDpykuBiw24cAAxj
P+vFJ2Q+Ag+5wj1uBd/X3mraivZjUjV5sD9WZ0mxE1xWFFIZ9Eqbuh224wVbi+al
Wtzk3Y/OEPlVQrIepF4uk9XfmT3H0RLiiidQ5cIfEd+FRFprLDRQH/8fCjGQni7U
Am6gAUJ/TymWcuEgSJLUjMF15JT1NITtxiAlVaqSzKUH+b/Lpze9adGW5twaNxOY
iH55W0LW7I1R4tqLosQzLvgqNbgMK0ktfvRI8BCRPeF2uNjB7j0nAATfcuQSXXz0
oIP5vr5TnCpFJksnA+AF8WffBMY3ZRNYbZ4GNx2xCUay3NlZHP3pAFy6XaW516u2
a8MbmNEfZJawCDLuUWiZQdcAeDKwKZYnH/FCn9hdN2zS9J/k4DpJDzFcX7a3w6Li
R2QN3QJbjKLDIsrwj7cvYMW+/QTDJbSt6TS7Bfl3Y+cmUMldhR1+sjIbnAuuVeNy
yceBuVX+cqie7dI1cxHGtMyqrvDXfQAd7lfVmxVlvz8BUsnyv7+uelRAIpZNtmZn
0FUSHpEM+BBuLmDnA+CmwUA1FgKN8Q3rNSe5i6zud7gCnIGe1/uFyz3kK9QtVse2
g8dcK7U2AukfA7/fEjMvlu4MQ06QIzgFWlUZH0AcggL7IHiP65KytZ18hpNmHT89
jgd1D9LrVbXDaV8n25w6t6EfrcQ5usNgnk9xyGNuQPEyqmzoe7edJ8WrcbNb89Yl
b1/+Bm0f0/eUDG4fsVgZPwM+EjzFjWqGeD7jhffHsPgpWrEd+/AD0e7vDaQZfE2B
+ZZHJ7kFFhX7SRVso2j4Cz8CXNzXcaNoICe0bfX9j1XQnGT9Xm6JB6/1phGkZjuj
RrVaUcsgyP6PD8KfIZBAQarQlGW9GScQVRGWj7akpIJ6tI4Wn+EZ4bVL2GnkNRGv
vgwJLuFMmxg647So35jGbvH3EqL3ajjvPMlpLJlAL50gErkHLdvKysHnE8d3PZwG
phBTqBUTbpxyDyuoY1/X5bow2PQTH8Gu4PDWPASO6vUudrlV9ZtVeoqLUxLbC15/
pZrW1pm/SsE3WYenmNvnGnsE8qGi/0Fc35rrU7JqgGs2MrQMLHOJJWVrI2AN8R8K
0/XkRcSQuufJ/Cm+jgwEfblVbVP2S0SQ9XP6vz4gEG+YARiRVzM3xPpl7hVr+/N1
c6E2NfP2kHJFeJ4hPB6CDk0zI7br+gGCiKsJbXXyl/bIR9EUgmSk1MtuOLum0uDw
rzv7CydI6tcIE0CH0BsMuO8IMcQMX8CfSW07jJFkgjNzMN1cZh53GmiyXBwxl1DZ
bW4A/vGJO6HfKD5XOj1vwr+Vd+XkfonpIH9VfG9Q8xJ3c4+rR2xuvGNB1fNxw2Af
bqcvOva3Je7P7THB79BgDKNQ+le6sLgB68cNX9W+sIWz30CZX/2xpboSFlX5/cVV
G9i11Ex6YwC0oiPxOveyVwdh4B7MWrtkrm16Ug33Q3FZpxUwwdlDKpSqG2e2Znsa
ZWm87LVF1nWPwdH9fyAV1DEs4Pl102CLUjM3rWkwdFTKj3zgd44Ms6imzg9/2AlV
Jw7tLHvEIB0KHpnH/KX2cSri0qiNoKJXhalZLfEpnII6SXcxfjufXyppC93wOUl4
YlHApw5MicEcZ9Xb4NFzVafnLWOwH2bMkD41tA1XR81uhGOr1+bc6CKk+SGCUBcz
kFgbrOYJzo5esI6Opu5Tz/r2Gh0XH51ws5U3jKEnPqEZs+gWnOPtXYE74AYiNjhU
G8MkqC/dLyKb8MG/WMXkFTqZJWjYpeGeXEVTOiMrgiuDUDegsqVP+6j1ZwoU5W2c
cItRWma3plKfU06Rhi+rCPTt4mYcUjBLCqIdX/i1y5xmj2M34HSlnqFuTcOWLTqm
Az8QrCaY9P+wCcmv8ztBjP6UAP/vPXGNiUlVS8aSLAlUVPXtdk5G5RNyOai7p4l8
MPRPxS0+etVsBB4DTQWmNLMy9WiCv4q9WSVND/C87Cc0H10B+EGvg0u6riyOS/h7
s0PACVFSDUr7hkQ2OxXEkJsUmxWTLg0NMVxhmQNTp5OxRDlVwTlNwQYelW4GZ4VU
FDDKtTnBXwtJGuvU5a6tfp8YsBnymW/cc7K8TGRYWvOdMd/ICktUSZBc1AcLiwRt
oQ5U1zMPx0ndKao16O5LUqGZILH+wKrIQ71AYm+7cYQJuCZ6RTXdRlP7jumZC1OE
ZtzEcfaNvoHqDO9IVacZHA8xRRIpsk/eQUnvJVuztVayeVr2qsg4kRXZawiX610u
aaiBFu/HXleZ+a24oLxmhDeyT3oq2oEJJ8qsm+9ofTDhIpsTokVOWW8XVosL67Pc
vwJH0XaDmspcunzDPcv5U2xB7pt2Twd7QY+fbm94S/qaScvg7W8Cs5Jc45oqR0ep
UBaylAD5gbGgXhJXdcg7HA11TpIAMeIEtv9Mv0ClvdmNKAYc9vU41bBp+x61g0Xs
5Uoob8RU9gWdJecK/k8KzGQLaVCN9E8RXeqAKWQ5ttwqRSBtjnuhUaxE0WpktLzR
yHxCv9HghAQxOYDrqAz0G3Dbm27K9BL43kT7hjYy6FjqbWPcZixESvV7l9E1lSHN
QCPhArufsst7HCOcrZXb4zihJnDUg/ex6U0y5kVuVj4Bk7D+CqIlodnbJ0LFEFHQ
WrjkJEVHThbpEIxJdlMlVmgNtIn7IvkOLJB94M/JotjGbcdp8nv0w298psVwrTl6
z8eZQt3nH4ygiaURozeibw9XjbK1wmaawf7k4vX6ACQiBDzdbATVzBbKsV8TO6JH
m3pd0r/ieveY67K4Ky6v8JuJmhn31FDfMGMp+uy2NBw4sK1Mu4qMIBJri560eQHR
XnnjqtzBeSCfdDhWRFMpM1GXT3MrPidZtjCEkQnebw4tPiMCIrwS4AJRlXD+r6Ya
Gp3ZvDZskKKMfQ64NR6Xln9Juf+at2G1VkADsnrWwoGRyo4639VdDSWPmgOOW6cb
m3DTWuPIvoT577OqloqtNCZlzYTuVqQ43DKAgz4hcXA6j5qVfDuxJ/MIaOXRwaST
DANhpJNvfKLDUhnKoJ5VoT65817RnKgoVx59yXUDiBzqD0hGXxsyIkDU68ucb1zU
qPfPn7Q0q8ze44QxtJxRPaHri8DhHWApwAGo2RH5ynK18ATeLMXwSa9jHOau/Zht
hzPUijlPQ5hYAUr+n8jUJNxXK3n54VKE47yaGNnGL7HK+Wz9GB58393rRYQYIbrL
VyQIbo/RDFylCog5VVZGax75jRnZSQBCCJWWfvJzPUOSLrf1ntseVgvtNNlfNXUz
S/B8bmYvdwiFsygETrC6gciBzkcBMIRnSD6e0rDnyyFNTLZMIuf1iK9955IVbncX
WB+zrFeE4CgEJRKofeTX2OV5g/pa4bHAWb9d2MoqXt2bgcT0Ee/0YXyZZQgx9XtI
t0MGc/FkQTtdiBU7AF6Tbf+eZKJskJjhNKIBrvJx7KfOCzXxnwUDHxSwW/s2Vzja
nVtafzn2YqqMzn8Vy3nCzztOy8Eef8h2x9DiDRasGXrv1mYmKr5BdLH+19GpVR4b
B11n2NBT3mTa/oICgDyuG0O/YOytuFb/0FZ11O0Sq6TRIJ+V4QkWXCRfBdwLDGlK
ZawwGq0xEFI92W7IOjZKNowCcUL15d3KF96yxqFVEpCnZVnbAj4Ms77ybF+JcNd8
G3NB56eTBG5+fS9qrDXcZ3+HD4i9eW31v0x5xBLuB9z2SUQB/SazCydi1HTEr2oT
LUX0vseqJ3adgx0vyoQicdGOUDqqZLRXfnQ56fMtD4NwGnQkh6kbW47Pm5zEJTrY
zDC2EAPEqv433o/BgFvXIb3s6vVq2/uZTQcZwV0LAMbP5uYvWn+lpCKmTfarnHFf
FxYiNd/pTqBe/UwMB5WqfUN+g0tlSKATo/5g8AyVDRvhLeT4S60AboLx6wvz5o/r
cgK13b/7AisFPefuomRs4Xxb3JUAvKxvwwm9NxrR7/IznQMeMkKk3Fghg5YSlysm
agnrxXI/uKlNfN/To+krbrKdFSL97USYsy1TYU6IfQmdiXBBdrBLVw49JmL1ux59
ZRUbfV5SIUgz5rwiJPqEzyod8POFIM7impJtLN0dquJbsPuutcni1ByKdunhqZL4
/Er8gec/3GLIHctHqbqmHx7KWBviaaQnIATiHwgGSUHa6gv+ojbbiK6IL7AXaEDg
xnwgfmesQOL5QlHmPo1YXzz6lRdQe1koGePwA9//bFOjxkioVuUH41hPRKf/SWfk
AaBhpKNz0YLJthRTqvX+czkVPnsyqYPl0zG3GIzE+xISe+y3LEeYqRz7txzDwW/B
98Twy2UOR4zI0m1mGQSAnkd29AWnFu6Yid0000gd1qSqxLZhQWgkbkjMaweFPIFv
SU7YF7qe8kI4VzzPLWzA/eD64cVt5u9bGo5p28ej2kOfK2/MS0IDgWhsozrcJR/g
LvgaN+1CnLMEl45saCukl3prMl8QkNL5PAPTKps4SG/dsDRWKyaZTSCL/zi5JnDD
J3yfyHeyOu+MfMpRTJ/n4p5FfIu1wlLtgfjL0l5yFbpKLR+OW/lQe7kVRpl5fRjb
aWpfAnMfzhpDmCn92BcU+DO7Awn6HdSap8Mf3wZ5FhTG156eK1VNlq4pXdQyTPXR
Cu7V/zpnbub/D4DX8mSTVSxWvQm0d8TSgeJppJnEI5GDjS+OHAcira5a268ovFYt
trBoCEFAlMzHblOZY/y1XNkhLzN1zBNMwlgIJTqGGTBaZE+yr65rQVSKuZ76p+9K
M9H5qTZKGp4JOGSI52j4Vik5RnoFNb0N83Q0kfLg06qMu13LrnB3OR0uoUJIsIw0
svUrwglpASHTt6LG4bUwOzAyVrI9d8IdGBnUSbJ/nFg7hbTG0ifC+p9DzGZHMUna
EVA8c6ks5wT3uzDVflie99J7mfM0vD/QLXGgeUCN7QyM31Tuh/eMGWgURt7xfAmS
t2uNrIUMbZp95Zd6PbJZ4HxMfuSkgSCQFXmdSeOJmcsQ7cl3IguqN85I9kfQQWTT
keWV9WHECrfBKNmz1Ny52ZjtQaP0DFNoUkfrtub+YBglEeDCadY3tUDsKjjH6bFL
AZ63tXjAdHfoNLlfhVUML0Xma5ZwRQTfsNxt91ZmL/d4Ou0mVLYEnPDdBrWFQTEJ
4/6CC3h8PojQZU2RmJHc6H25c89YDLhb4+KEpPOlqSIUtpCvnit2DDSQUg+V22d8
kdTZxuLNKOiuGYavQVT0DiT1IE5uPkS8FoiJ0q6uLDrevrnO/jJi83a2lG9AoRWo
P6SfaImw4EVsDFIZUTwCaoRM2M0zIMZ5Z3ZEpQaJc0siSltzYziC+S5tRJF/fhCH
FM+B9B1h55WFpcXcGv2rWSGeDs4IogiITYgof/Krftt32FumQuQ3118duil1TI8o
/BwnNNP+ECrb1S1HMySjlCSKkWy6d9pB6RSKMHMebNtxmQiM6IoihIBCW6KFcSXv
FxD7AtoSw3WVZsrdUTwbCDB3eLu4JJk8jpM/iWI9LhrnbNfYtrV1HHQVo+SCMtgk
P4UEtK3MKdKoe5QRCrmJ3OWJykttTKkGThY1NzPACkOSftxOklviJl99hMGYKOk9
aK0jh2ddBzKYw4e4HgdWruRwgwt1DE43CjnMHXK5pg/H+GtMG9dYECZFtWW2xrNG
8KAz44yC4aMRRlTdN0YZKMNllihKkmNXQ1rpCsc7hEODMaoffDtN41lIhHNyYsMw
3zMz0OJR21VJuFiqrwKo0N7f4L6G+5WYKQunmuHwsxCvwUYDjKtqupeQzPbP1OXo
/UVf305b0+SAW5IOLD4X3v1wmDbk6UxF8F7anwIzf4F7kMCqU8Mdki1bJBesUNKz
U5iXtCOh/qXj0y6koF7Z9p5G8s9lVWV/lgUgdvLw75UHdMgbumdQam+fwtW0kkBi
t7fJLSN6Y6sBIgQoQ1m2GYwxvhv+xLl7otGrBafJhx/RWVpchZPpsdTvIzBtZoJX
6SCxHxdGhsxcKhWOa19kS4PW0bvDgDZoYPNsSULEFbJ2TT/EFnWVg+v0L5BGifmh
2ztWo3Efz7TcgsZ3DLPGzzdOY5mo2Nn/GbtpB27uCYwSfHGB4frOP9185gO/veGv
823mLhCCb6i46dC6MUQv5UyUWKvwtfAlcJKd6oovn5SP9SAwUnlOqVB6B1wfBh4/
BpaGp5WGnno0/8UJw/kHaFc8fEDI4qBJWDDhoTkUEY8xhxr4gq8Tkjtr6r/LCECy
Wh/Cow7wEkYoYBVDE0vAEt9aSCXWP9s8CZr6fp7Ky7eYlwtuaQjcwf0183/MvSuF
DKmTZpx82FMUfXD9vtxhsXWNzBU/e/3jsJ2UCrF4vFzbHEXZ7a5kiio2YAVivXMd
h24haJRatv0rmQ2Gmd+RwYytKU03thqz9h0aVWfp/DuC18wwGVJEQ91HvUsi4ra8
3zWk+DVDCXflolwFUym0+FSe4cQR3S0TV+nukFM3kTZa6xOHmx6qxcVwpDG1upjJ
XGHNeMgSiWmw0nUMRNqQZ7BDP3hKNhUP54Z6XdrhvbSvXiVAQou+sKZKnIAZ46j7
7YDfi0z9JDeW4rcTsh0V7BFPZsum3ZMYNbnNzVlwwbUAICIP+YhPFa6d7I6c/ruo
zJ3ba8V6usPjLn0C2lxJ1owWV6HrrjnjA15bsVidE7G/Y7RR+gl9wtsLtjImHzDQ
MlQqRgoeluuKH1OQdvzjKjuEQptSrJNQrEuX28JpGnwfHg9vX0ucoJjGPAS0+5Iy
5HWvVvkgbzZvjPZ4NMSwHXwT9NvubnDym0QFJ6SUdf512EHgEsrrHiV20h5e/P17
esuDPMTGyR0Ci5giHi62C2KaZi0yU85fIq9EPt8AyHZAydMFekWsOlRwCA5uOdac
K1lAcuMCX6pLYObVDPn78GgLoOSr6sgoD7UfR9VZdXThqJzn/t9aek8Tz5ppOxf4
2FxhuBIn1/AdQGpB6xWT3mtdn56mvI84nKruRo+kvu2FRjzMu0vPMHgLrBayU+nq
CqgF0B9nvg76NTiSPtr8IMWhn4DFeLpZIshSfnkOE4m8EQdyoe9PiL54+e+HtGsI
r7tszRaW3uLLHuIQI3jpl87VmuixFoacX+hUPOa54KX7lXrPNsvYdtIsjZAAA497
dLbzrq8THCzj78hVoptOYtCNjrT7pR6iWJ2JFEWcXJ/Ul0zDH5GtcytG82Uv8AUk
cv6zxsFQccu/Rg6qk5sX5mXjvIWxJLlTjDwiq6y5+Z+TVtw/LthF1FeY2CQvB2m8
7P0AHZkyE30BOSH258h+9PenXX//lEVo7xI57bAsnfoKUCCGLpry4hGrjm04+dXP
xVhj6dduAlNpAifAjXmBQuEN7gidPFxrQPV6Kk0hGw0MbrWYaZNLjSh+8wPClqhQ
F690Wu4Y8uTMBnfoRTVchxOC4XmtzlUfSkx3JcUrtV8jhs1Z39eSODGZytAf+12P
kizI0kECyeaxwGEA61V6PITcK87p33K8DX6KZ8nZNUf8WXcYwyMI/dTsa6JLW5ul
VmhQeBsEJXKYBrG85PI5wK/g+GxwS+uMsihzsq5/gw2aEu8DlUB2+dFeMeyHXBco
JSsm4IpWQ8+2ME8IhqAOliLLqFi0jSzlYJNYHE4jYQ+6oDNBgpmzAB6v1uOJF5TJ
wic4RP56LhLQk0vjGX9he5MJ5Qr+5flSSN6jEWLz8NuH6iaGtzbQs5XIZpWOLync
Cc1JWqmlYODy8+Cu7bjLWzHZw/8hBFGq7ZbXsSQM7P2glOQ/GIYM45kxc8Va/rTW
jfDDfvr9DnBRIKUzb1psL69apl/q4ENOu1R6OLQ9zCRkDLe0JVPCk8mnfQKCtFFc
XL1GYk8n30OrfsEtplRQiP2ksXLvbr/pD8FkuGecZ8eMtg2T9AcVELznT579aHFz
4wFEd0kCpkyHTnr6UbbKxwvIwv0QPX4VFFB3vzAFYL4lfJuzMAm8GVXA/OQJTo8N
/ibmqAmEWQbQDn2DCl7aUUcjkp5lhm/5gAnqejVvTioAXmLB23Xhclo4yMny0Gkd
sqpxQDc8GlX0pYN4mu9i8QH675wO7BY8oB3CH9rjpn6kutIOMvxwgPMHFvzVbug/
W6r70rS1N5zjNFQrf2Vzyx8w2xhzC7P7VE6KXI5S6yO5JH+v+G5eA/2vSaD86Hb6
IgpC6I7scu1Juo4a7cCeqTExQtevvLcYFu6acfMvk7UEnf1QbIV1TG9XG3H6QoKm
9ZbnrOIVshLQjq6SLFxKVIFoaTfknwqYG9MAt75y2tp01PCikVM/c8XshhZ3+dfi
V5XrCK4pGivmUcri0IZgVx6BepG+SrwmWg4sLE1h74BODimCOsqt4F4HTeOnGy3x
E29VTGALvkHLUpImoq0RekJPu1g9BF7cYATgDzFwmk8tl6u99H07cn+EiPNhVAde
23DezwamLS5oJpLhcTtvvbYw9MchjUSvAUzfLA9dc8HrQRdelLRJA3/TXvzVZcBW
/DcagCbmsOUHmu7QuPDWRP4Tn1E1xsvu/btuiQb1lacrjRSDaHHU6eiBJujSneBs
6myzzTLuMIq4D0vMsWsg1ENE2vqYwykvvQ2qOACP0AY2z55uW4BYK8XyUO335nsA
I31Mh9EgLdObf0/KACUKAPcx7e5QWnJ1yoDQK7yemnxrqcm9RFNbW6ZxMT3oNTI+
BZHtb7GPhTGTMlBFt5GEJOfDQLaebfCQnHG622GD1ulLrLuSg9IqYa5rI/jteP6v
KJADUAzXY9ZDOP91xQQS9EGmRy2uN2WBSRknVg+Pb3MJZ63fjj6zIt8C0RrU4i5j
hb3BhOJRI0cEErz65j8/UKGTEIKcbhZrmY0ltapybxkLDmGXr9jTGwQYlCsHvVnv
+lYIPeCbv9PaCxvQOQsFx3lxx4F5YxQsio3cVsl0OMsyqPXCHL77P7UKW2NoRe45
GYpXSwKJudC0s3L4PXmLLCoERhdeSxkv/s2VXVw19482gbxHMZRtf8FuGNIEaNOq
EYL9vomVJHvwQxbRIg+T5fqY6JaAytkPaX4AWfNj0PAO/d6cwSLPNYXalZ3xUYSq
3CHUZ4UPU+JPfCIkMIhT5CxfNvFy3rXyHtZruvjhL9mz0DzfI7iNzT5uWFcf5M1O
EPKW/EAG2yJiR0QkfIZKi2fsVjtyY9txnzaoKPoPSj03Oo9Z4/ohXjoLTjgk3ni3
/zBXbU626MSJfQcjWsUO+xAOlOs0nq2+W6+QPLLnpxMoWv/Y+qZ04oMxM/QkYbRM
OOsprniknVz9Rux+URwAynh3EKuztNEvuyH9hQHk5pNCQzd4BzbHpGd6Olaur1p8
DNNgRGGwA0hmYrbfNuWStcmlibV/b++kJld25cV3bSvZKJScRNJnxUtP8RF2TMRq
ey+F5irMKT1ImXAiGXhKA+imi9ipm+TS1sB+2XxWfuaZONdGhCotDQHIHNiL6wA+
1Hf/nLBESbkEefCFX7E+FjTwzOQ1GggUoHoqQJksi2tz3z6VEhAvvsKIUHchOwKH
/HndQBMufnVPzy73xwskky9hbxeK6TmakJVnX9mHvpzyr/IqPQZseJ1S0AQDNjgz
jGe4cS1oLJGEgSnqiZNu4vD1+ikDvh8K+afaW3iOSrx1aApgVm+qOEbzvrFdO/HP
wy+6otO2mCVwXaB1Vf6DRjLwzBIrxQGQIdH80eqF6dk3uKN1tE8edbqcMmQ8L4Qi
NYE3WdX3W005f+zXXp5d7+oXfdK1vM4R+gaRkJ5yZkCdBDjzb7u8Wx6zZzkk/Coo
qdqyYF24mYGlLpDFQnpsHXUZrudzbnWsHaM99swBLtsz5PRZIr8iozdxjpcVMm8c
2UyOFgCBsWigbfQ4yHOxXpFKemcM6xHCZuhWBj0waQi1VK1lJpVfj1O5Rd3kpQMQ
ISJ3Mz3Lp5lsmORvFw76/CXcraOxoJRI+hwI6oHqw5VE4kqPOkMmPIVa426Oa3CA
71eO+GCupL2pqt9lGr1vOam3vszVJPmNzreLGyVWXXvli0cHiL+QJSACNP+veTxS
fHdNcDw7S+ObRJKRsfPedBNB2kgHo3LPBOlzniUNECqjyuMOPwkK31+qJXWudTdC
OJMe10iktkoE+dgsSGislkGp2iqzr/pMn69oYAUMiuPkcuqdUkdHN6Uwumy473XK
TG6ksodiqIXi5yxTOEU6i9YxuFfGV9W+faP3fR6ywAqnO/pHPey053bYM/sSel1k
t6MRGCLMqKBkIxPkk4nupEAsbqehHgkKuRkgfrZtIfL8pl3ztajLxjy+kZYUUrIF
iDxb8I/J/ZnIzD7rI06We/UFpEBPBYGrxyaHjVZY57xyyIOMXzQiZXG+jg0Hv0l7
b0zfSBfw//jLMCkr6nCnDtdI9gwjQmbczNrT/6oXlDM9oNXUvPbsyG0Ys7CFHiwI
2OoCa0xB17+RS9n+sT8xffNi6EHsOgdmdfSPUeVg+LjAbxwLlt5cLbo47Bk4YhIj
/HYbQRvaFnSwIlwc9FBOgKH3Xm3KC+j0h4Mz+lGovrbUHhKgJvYZv9GzJ8JbaZFd
+9RxCtEiX/H8oL6WSgNqIBXt/m2zG1qw5K5fCkcmY2Mxjc0lq/7HvpcIUOS5c8jc
58ZdNwzR4Xn3RxMAUImvsMD6vlYjYG/bZkxK4jShRN6xPtr4PeVUnT+EJOe5OJ9o
ZLsOTNmO0OvU3THkl2L2gt//h9Uk2MCS14fdGLUvhZniD1JSzK32jtOmLYqQtROE
YQ3gpoSNfKXrL4PRK0HzOzikIw4hNBFEqQsReGhQxfh3pBBkOaq4IeF5sDl2FkBm
GU71ssB1geLxaECWb8O7vmhVaGBeVMdeU71mtT3WCy3oaCSvDgxZdqTlqUg/HilD
MtwV2KgeSqyKq6p7gDvZBWm4nLkEfIvk8M3ubLQo+ZlRUWeOGhXxteGp5rRLWboe
VaPcCkKIT065IEC2ch3GnPCdK8qRSjGfS8cHlXo1EZZGFp5JEm3/Zvu5dcPDFlSU
f2LlEIIrlJr+WJnhEPobTCWtFyGVYGp73aT+1/r04xWVP1zC9kLYRvFW4GWqHA+Q
mVx21eANr/9dPmFEFXwI77eL0s5koh0v8EIEA/G3J7wUhCSW7c0Qagzy/7sb/CBo
VLuaUwmHPEmy7qgXxh1Sbve9+U/b9yXf9eIhqqNQrkK6VkWYTgn7QJ8FKgmf6to3
lzK4iZRPorsKwzYwrJQXOOBo2xFJ6o/dQZ/XZZdTAH/C0itMgX8dRiE2u6rFavuW
hYie24n+5DvOXSb5KGF6ZzY2BvZHkgLtorCBvCOf7GAzX13q83n+5FgYmpatPRF5
iLxfC8wszau1NoUmQhXt2aX2PTaZhQx5yhzMVYStxzAch/m3kTxjCMANtLUbQesz
7WcyxupSQDdAAfXGKlxEZenYocHHAh96KmmWi+dVzvDidugdoWGVBubKbaKIeMGq
7j+vrCp7FCe0tMRjVzkqWHmDY0nXo8YBfPqGdgkXQ4izTqM67K+sMTML3ZxGmrTz
hP4A7YyXbyk77eBrYxgCIQ0S18BIyIb/qxFg5eQG9CTroQutspBePpeUbgCGHv8j
RCYY56c8ZpJxAje1/gVUg4ePPyh8Es7DhaE+Vmy5WF1MhooNhrzgZxJ3YLFlSW/D
cnBAT0tfVB/vIJz3YyqRa3EJ48nbGeEezCJU9ItDN4jClDb9R99+mpo7wVW4B4Ci
SSc9VHSLjeXXICpUnFOaC8Tb5or/ACGI7kmL0GcvGIpZPQD0Pe0f0V96a9gwjG7w
YCL7PVC7OyvetwaZ0LhXHghABW96urpK5L/1b6iE1zl4dL3WDwp0ZsyzwquuIT97
UyiZxzpKwxS8BZ9Wc07Yqnn19SoIHl5CGgxOc+OZND2CVUoeluo0fL0bE3Q3mqUm
8wxqgDUzTzAs4w4Zjfn2mfmokBFtk7oEn4gx9ilGKxWHH4brXlETCRishAgsdYJZ
wkRwwBhhou5Pa3PP6B/1CkK5E/98ljBuxeAH0st6/w0zLYlHUi6WDTgLWVPawwxj
R8KJdQKVE5BCK3pRsKoG3Kn3sdOmvrz8kqEza+w2QEooLzFQK3ojXazGIXeE9a2P
NAUtVzUh7I4DOKmW3jmrWO3R5RkN1z58ajfSxTA/NuBY6DIXF+SUlOo7G1y0fJGI
oZ1sdvRfFaGj+6ZiBdrdsT51myHr1XvDxnyjevaGenfIuAnek3fAXGxWuJBDSv+y
mEoPQNwna7XlS84ZtGnkjeiGQ4UG+N+1aC9o0uYGxWlVus/xIJHWEz1slVSMFnpU
QO36axSW1EgYi3tvPhm94cjxOOcVSxTCBTbPQPWwtLGDc7EpsIUXJZ60rZfWSe1x
yEiHnlFEO2OLYRjnp65jFKF8g1FwbY6ALu60anxvpkbbl9n34mH1qBfrU0VeA/ZZ
HlGfkFRV4+aV3X2TwU5o8dkkACV86RVQFXeFH5/6i3FvgKXPSKs4UiWFM5YZq5Pw
A2kSh20yw0FC9Srb4CuZTDZDE8PSBjwBtPAdEX24aHRTAZ2os1x2isLtipquj3Wb
a8SwrbNB0yzAH8/IXMnsixcM1cpUqkkMzYpasFdpJsarqGN9EkTz2rK3KRsrQqm7
8dAbKD3M+ZYcWo37+5Nvr2lnzfLHbapiUvftRNV7X/2q9BVmdNrCG8JgRj89pyhB
Lo82MjGvg4oanPuvBr5nNobqg5U+3oGkvUAhLVLxkaxZ9oPbq3odUtw+3BGwRtVc
4Ah2dcEsv9eQ37k2bNbkiJmlkBxxTtAI8kiHt5uqFnqQFyNyUqZ/vP3WWUwlaxKi
1dBf7tDAFpnjBLXP7sXSFf5eRzWzt2TleUEVTjvq6mU1mZ0urLU/y3DzxqmcY4YI
q6WgGBAnIIkrivK9SlqrQvp6U84wDJE/1KK7fYusBdjSu1AUgjNdpvNQXC3VxPxI
qAPjqf3lBrlcWmxqaAhk3YeIVNYKXSz7XMjivTZALSfOqb8mWpkCunTF0qNa52pS
/iSKEk+U8DQeTy3eNKQns+1foJVbD6A6QBzXAK6arizDUy3lbILF5LZ8Gu3zIBvK
G2C1TqjaDvzTpYa0J1u9V14wOqTrBr+Dfrkxi4Jp1MyFzioFRBL2PAH+PQvO5Qhi
zq7bwjyau6Ea2AvuSTohkCcbWfrOGHt/rdq2ttSlTSfGSDe/NnZnvB883L/yFWgM
7tBG6U8qCCsdOPpf82F5cvSkvV7Js4oqh2HqNi5WdSR2iQ+l9kNCdPMiZQ/pCTJJ
WC1HFAI6VZncOth+9PLy5MDB7tlPm0zbLYptjn9TObi8cgkXi2sq7wpuRTV8PHh6
wgcgiD0RMngr+X+N1cgoWhYIe2Xxa1HZOe1amLgfnJgco1ZnvnY+CveT9dFeNpUD
Hn816Z5S2z4xvTUPtW+2ppKhFGdwnK5eC30+yoHTZYZRKe6HvJakfmNwdQj45mJB
6GlfrZ7l43+U2exJozyhFrXdQjz168pSa3xV+4635rB0lwUBcy86S6cqQ7vie2oH
P1CnoWM2j90x+rHkNL8+JQMU0hV8FB1ZebQtBBrGmCzzWfHICNJiGqqQzmZ0YDKb
Nc5fco+W4ztSxJHB3d1bnIQWOkKig6xaspIMgslriAAGnHEzbT1+MbpT/g6O3ecf
Xp4+VG10ZgRLw2T8tIg+C7zAls2JzCZk3Z2f2ut/F6aNIA72ms1ssnu9nIfimhHL
BlmzXF/ySxdJEJ/OO1maqKhGdOjDs6n4UDYepk+ImJ0jjlvU04lMy81a/zfKwwcd
T2pwgvhUiiyXo3kIyk8HwKu6NZZl3+tcqcJ7pVqhIP5VlQG4WCnXTrg5Dc3G0prh
l/pVk0gh0cJWoY1t9lmgTOoy1H/WIi/mQeloAbLmYDKkPPTEBtT7vU5hu2Lz6To9
uyrdsbZ1oqLx3j8CsINA6wOVwX/3t+5ZYF5/nmq+6ReJuExaSxZG4QCipIvOGSjT
+CYuWNdfNsdCh4uB+0I7/JMnSD7/x9HKA+7PoBljiL80IdFH9WmqPNUyUBIUSUKe
h6f0MqF/KRZ6gfsaf14yDFVfP6MoGjJKVhgKV8fLa7c/pa4NhQGcGJ9e1jCKFPyl
q+hymdNSFJ+m2wLrH78PP6CI0VTGm96gO+taHBDtJoD8gss/oBXax/xfKFXKMw6l
+HLHxN3jym1MuQw7dg6m7k9pDtGOIjKDmVGFJo1MhravozrFmSysM1h8PsyPPwDb
8dbKsTGYNNsqs/WPW69qzRxWB2AgyGy0TceKp+CFERrzEb6haULvde6vu3T1kc3C
9+cSN4A54qvQlyoS5cbLYB8Wqvuq85Cipuf6yZ60eTbDkyO1LCgiTcPbRm45V361
IbSycS90V6dZH2CCS6v4aJfno5qZBrzMxP83Tu4xodqR8JtHBKQRmfjaptiIj5Qb
oaPY33y6dNb3BdnLPNjByBiARniFcZGp/m7PFKceJx+M0ewmL2xXmHnFftzPERVx
0zssnJzV34Lg1LSR01RuhfQU2f9ndj2HC5+UtBLwGotDY1QthAMt2tTLgDBVyEdq
T1QRVI8UewhhuR+60kAXI5xiO51Ehi2VZJKWO4bymkbntxHTkG6P4RJF03fqqv8E
CF0gwFk7wleROnzOZkqzCop+STA5yhK6isxA80S55ge673KUQs0545218My0V4jR
5WajPhzYuGFJkKspUzArqQzR0Vthhrn79MzKZlnAfjkvl8IspHnUgJlmJIZMzdlD
DrqwqTx76zpFpKsmzP4QLU6qZMxP+RCZW+ftbos/lbCikdQTYOHazwTxgg/9g1Ja
FbVjQ79ZnGAVGsWfWbbCflin54u1VKswjWwrN8ic2LmK4JU8JIFIDKBVFd7TnDfV
e3n/TWKyQRrqUF6z56UGGbG9tn1f0LxFhINB+Lu+7PGPI0kWd245cCj4xFqPlqDb
t/9b5xCirmuA/5AOrDcQK2u08HJERWi/UIPqxIBnWaA9soUI3Apq5RoD4vnJ1hX5
qZNUPrLaOTZ3wM9U+5gwqqKbvzL9MWDEVWucrxPi/IfdvyErGIqwkMOqj5S0FxLs
xLGXPay/NyQBgWtkVibBRImRJMY8TWBbyaFQ8da5nW+xs4uhYbI3gSSJiyz1d44v
aagMyx6qnBSS3K0/X0IWMF/hCuqs0y8KxYeQCBmTwJvMuATpSpYCSBMqOHKEnsnZ
Elsx1X595R5hKLIYeucSOnioqbU524PbOtueJX/Ij3L/jaVFoA6T0yIKqlKibPnC
DZTTaHxc0MDrShz8SlnILhCdFZldYdKiKTgij905j6qyUZlnFqMmcZKgclDoSDv1
rQwV4cafxjYauKtSuCbhr00ymXbFITM0CyFzbi/pCgBqF+J6POA1KcOgf8cm0U+n
v9ZPwNFsrSTHpocCqY0fQgfNC6bcnV6SdbAySVrseaINzO401WjGvMy/6w6umSRU
8wF1oXIxtGOQ3wCjNjU4u2O57ulukN2IzHu1Mpnm60p73PROJNM07xIN6Ad285yL
hJtHMMdLiPuu0zwd+3E7fd9Z/v6cAGJCPV/odfi70bAg+14rUFbR60IXmiD7OEIk
EqQ9iADM+d/qbM1TM9pr3BON16UhvpG8K8FU6hV8eR74NsD4d232TX9buolyL6GP
oiIefEQOoW9AgKRq74C1ix0ui+FXMl5OswfB5fIDpxOsYd0xWJRQf4h+9Sv+XZ+3
tAHrVCaAYltpU8bfaig7VSv3QTF2jczxZkBLVc+yn70/0JDFIglEZ5JsQ8bhT4dr
GjgJTheN8WyjsIyAtKs4F30tbaOXuUQjIP71zOSdn7mn9engwdGs38jK+HfCSKWq
Oi521dRf54BgTPw4uH2d5yA7cU3qvStCbdlICCoLSoWy7IvoGQWaFWF4MVXGxF4a
0qRssfcTNGspiXQWenvkenMtieLgK89+tRGWHawXSGxImpqpXwmNsG1Kuxmr7JVR
iXvOzWhQpGDjVjEriI/WRcH09tTGHIWvec/E7IKYcZSa3vtMVSVI8JfEJBug4Mpz
MmCnd/IsOlv97sw2JedI+svJNdil+OkNSLB4009516bLwS6dEJO3265FEVHE4Y+D
LXyV+Wd8YJ9GdJN46GbAG/POQq5H9GifUry9yVlfnlK4yPZoSMsu0DEYyDo2176r
iBpbQmR0P+rkkzD3mAz3FG8GFw0S8/trKjp5riDivlm3fBotQOhBxZA9ab+w1mTd
OKRGr83Hv34pgAcSq4NMd6nB5f2xapW/lu7JJS7TnPWWbJNEuIFoZAAeHwCb7lek
G43hhGBowjy2bAYJCEMf5x1TZq7fHAn8uSDAI8dCs5V01HIMbt3Wap3RqRhy+kPn
nIVrjjtatva6Gac4L19LZVJUK+UO+Tm5RLChCpYvKZvzGEB1/YuijhzzQkW0o7Nm
feWCm1zYaNPryH/BPNu2MJBKD0O30Ox7sUW9Cpl8QkdvwjqQ2M5IL2yAmAz6vVd0
m/JuS1oFz1m8Mja635F0VXUSoxLQwBuEBfzB8RI64HkW9oQauUH5QQROPYQJuBNl
GbsfeB0l1DSHMMkgy0PILck4rDPt3TQBktaUVV27bbM1Z1v1/y6oqnK+gRpoQZhl
fOzn8BqKkcAHeh6gHxJm/4DVyJw9KhhkFLCEJiyUFk2Nsp8B0cxp/4SjQmZuOTsI
uky0ap91g5a4FwmCIEaOJCbJCLKe48qvoSLVuG5xfuRt369UwdmUhxMgaC5pTs/P
EKgulsirFfv805avi6X5Px+U4RiwHcUi3gfI9wmuZxuVjj0T/z/NbRBd7/077gN7
loNTI0dbQ6xCf5rqWq3RtO7IHMAc0kQ6VXRtqcMldGoNa7sANEpCE7oRFnZuxxFC
xucJ8E9s6I7ar65F1s1XLrPLoPsDlZ0KqPfIy3xyt0p6E4EdCwZOi+mLRiMGtdjD
Bilzp6uUgS5eJVpKpfnD1VKD/ppVp3XQMt94+CX1neD03Oq+KAF/qgfhK+CYo7Rl
tRGLR2lpTZQphEISeb4cMO/Uj0fiWYIRS2irBsBrXeNbdwbJd9P25bYPFb8OoLDw
Rqa7cgyCOYD/IDbcHPmKriP5FU2ywsIIY5uHeEv7AZ1tohwKnMzd32OYKxsOPdhG
dfLzknIJTZ3tYR3cmAC1NAEnkXJKjrRhPGKHFjGftVTqm1FVCn06+CUhYN7QpAqk
U7SYL1NoGy0g1TQ9lCjeYUpDSaTmjK1mKJ7mzD4BMCpSSkmisp4zZc5XE/R2PzSP
evMtnaxDEYy05lDfAPUsf2o2t+NyVIs/WXxdze3DALE7zVtVr4ipLi8lqEU0k6lU
t8rqqpdP5E0+Zh9SkPYInbc4J6Dqy5Xt6sB+6qk+r2SRp5bWzxoG03jQLj/MPySh
jT9mVuL4uhbB/ddYj/olRRXXIQR9SwvNX1XnvqNCQ4SS2r7jglsa5uKctOQgX+uv
TugnPjsr5VWHwcElnIakqWXcrquuS1rfUZBGLH4Jlg6H6zHDsHTToCsaiqMsNaDx
GxbTnH2d5TH3pmWbEj78MfEz/beEot25paweJvfjfOV4YzUq8+DK9y+IWqDFr2Rs
h1ZEkA7Vbr0kzd41Nn/y4wf65+gcyHp5dIXPlcStqDuBWJhvSjAu1fHkpWz1uYhT
uJOUq7w/2u6nPivEE3tGfDbCcDfN/OuM3f7aDuaV98u6eBRNdXvUXXFVrjdG0N/S
QFHLDSL97GqmdFUFv7koV9NEVki5twIGJfWaEx59EC5rYm+njEK3Q1QV0YK7ht2b
m7xyBxQscndaREVDOcQwknbpN7KpCQTPnDgZnLN7TCmqpbGtsLy82LVaCTUwe5pu
pkCDOia/5Lcxb199Y3hWyIRIGwMbJCoZ1B6eLIBxFh562D9mAHkufRiBH0wjOhCt
HaNoG/vKtqGdRn2aLy+db6Z4O2m9+hFuAy0LGwum7muV/jDoth2ybkV5XXu+RTep
Xdyto9e5Jgz2+6Ztzc+xRuCL0jXVd8lC6u5+YCR4jGonhq12wnvgr7cTSe1BZQNb
gtnTcGjlcHarKKZINODnWd4F6VuJHpyKBcxkEZsOyJ3SZcQU1+gdVu0ilyVFWBpo
HItSfCiGI5zxfhSeGt0aPDHD3IjcPygdiJcNOlh2WRhoIBrcJkctjqM/RbhMKM7f
W0tIpRVbwz/vw0GAQxZ85tzAO5pYOMuUjold3I7zqhiwqvZpQ2CIQ8rUVQi+k75e
ge++yENJalKuWYdrj9EttQfihV0P2jupWhT6bGa9sGC9O6EMVw0pfafK7fPEBLSQ
SQ7OiI5ObFeej3h22l9fxPq2DsYnRSDGY3set3AV6CrJLRkGKwDQXvT7+QukbVSW
l7gpq6aSi0qK10+83/i/CP8T/vHrYdbenP2+BsyPajJge44OwSXcVP/T1EI6vIyy
h9g0cVEsYREX3QecGrqse9v8D2k96TyLIIYuZjiluQR6wlkEQaA/Wnwm+gjtejD6
xrZHIa5XfrcVBnAUbVU3Jp8MQp6bwLAYhMEZh0+yw1xafsw7Ag4rS+gQTYtj1rmC
9f80RP+HDmMq/S8JzHNyYJsoQPIl9x+2zsARwAwhMXtEDC7sf7RjUvikoTLIu720
5YoRPoapfrCgiN27tjcy0fSHaiPcn5xUjo5Egh3wUA8Uaj9Zqzhsb2NgYTMCN8wO
T1w52Ox/G4iq504clFVO88+9aGNqW18IS2xIBHniiCFuFTBfX+tP24wofyx+MeJS
JQ2TZbEf2ZgEfZmFv/s7DAJ7XETg8k0T91e+hBY9BP1mum4v0AtCedYznlzWp8XQ
TcaKFOuqIp31qF2ONDOaAWVx3ZyFohQphG+PhNGnYBBvncr7VMHHNvYGQ6L/pijS
VMH1ETv2lXD8M22icTF4G5jclnv/ZW/8U4i9/zxDGWdAfGyNWXbHT52FR0U54Lmv
tkqn1R98YNT9ZrYoeq268I9dE1EDF8LZfmTrWPQcw4x5f/uTyA8XjImhTw3DZ+fH
gZcD8rlVcp6lG9aHwZOzXDeO8eZE0KoxTqeN+SCOP9xvvFzXRqLj3BdethHAloKH
tU0GCX2FTup+NfRwsS3gJIqAMJF1VsUPA6XlU+5CpqTh6YgdMvfkwGvXURg9NAvE
oYEX0bsNPODK8BjGl3TLc139YvdzQwz4K91mo3DgXTsv18at8yi71HiuJJQl1Pqp
evv/fXm56QMgGsTrvy74G3MP4TKtonKKu+R7vTE6d5qltC0tnGuuOm1Ca8pzsMCk
66qHPMYCwxhPL1Vc/t6iLinouV+6EsJYbdCRSez0ax6AyU48+Ybq5FWCw5FNPkPA
7zICa3dSuyXISUA+NzB8R/y6lUA94RkTXT20oYbKhHk72GwBok8JOxuB+VVk94iq
eobSwqJxpRoRA9GK54e+eckpjTrlcPz8+XfTCwjtaZTfrnC4lE5alh8hVqI+rtXv
iea3dd6iha38tJ/9gbM0Oqz3h+XCyhmbGsbeM4Mv+l+tSq7vMhPsWUw4aJXVF/0j
BGgc7doA9BYFywW/bKPvGLg/I/6gWjwl1URGJZBSamfDEItZfLnEfawWGIVPGyV/
FyoLLtz+B3qAJWRyFj3s2H0hBPy/HWNiCqlrs0HXiAbwG9+HCCCZw2DHSp5lAxzz
r02THITSCXv2019eGYwrmBpu7ZaWhiBsbJAHS2+PzI0d3XvAHTs9pJYYlgz+E1Ml
UOJ3Z+cECEKYFKzRIKJuBstU9I9rQ3pIcgkK9Gse1Wld4XAF3zrT5uptI8G7w0Uz
ki96lq4lxJ3WY7IaUbOtM8n4Vk6cE1kuoepkhswsOZemjJCcBkcyaLVNJvY+XiR3
1Ii8uug7eL8cpHUbz6rB6P/SLX+mEeD1/cuaKYvUlTEcSrT98dEYYurW0WxPQFug
oaf9PHKE5zFTI5wjdpsN0W5Qq1JR0Jn7iHpChZ7wV87/ctDP7wjJMUkgERzyJsAN
uoBt1w+UNA/eu2VKWSQ07vs18tBZoYQBbhJRFrq+NSA6sy9kjKjD9o14zDRChKUh
IRebCGVdG6G8IQoXjNsplwa1USHO8ZiUm4ffxBDFRTdLozrhcsBgpwcYspiraws1
411zAEd55raoaW5nHER7Bkj6EeJXH0F0nhEW3KIL+i630+F8KnxCNxmTgY6zbMFF
uDRyOxXG+XWNPM2TEctQYKFw4wYa87ykYMhXJHrqsEk7D9bWq1CmLg5mNjNTnuUO
GrMgfooKO/8rHymaOHMrrHRkfz9Mwj/0Y9DJU/vdCnqei6ynmBMhDdukld2+/nwI
te9qgdIdyLfmX2qhAHLiUw4u/vyXk9LkIlrLxC49U6326XRj6lHoQ1dmYGZz1PtX
7fvEZ6/QHXZZI1WFYMcTZKQqTJvrFN5+jWsayMEn9fS8PKAMpDtrAe7sagqwu8Cj
d9fsvyYR0NrFXkPvhz+j480Wt4SjF1SSWe9dMveXmHkpzGj6/AyryeXLFFCJ4wBc
e3rUvOVZHDJeB2BXUMQs/vVcogJHH73Hc3jcDcoPCoBmP5tZh4GK4KcUwjkum2KY
0XUaSVClLUfXpxo4thswNIepg6NlruiDMyTGY6SeCrzm4PQhv2bF/eR8+TF5z+H1
Xt6LlgYvzRGLm1yzSas3qJ1ZjaYU7S9JRjgIuLFUiKya8ytx1kV49shNR26EEk2H
pqzZ5satNKikXs9UZ0RuTwS0irOEzluZrQ79HEwCps7qN99qHktW/ToJDd1XAUVI
GoktCY3TL1zhWqHuWSm+BwHqQNQO0d02y7kI+f2kwjpNHknYdgpSouOoVWUfcNDQ
PDQBoBJSrc9xdd0WvRns31IIYD0GDugYaYXc7Igu+KhTWLt4iO1Q3NIn4JRJ+KK2
EcPQqyEbhalJlAbhJd0k8RFCxT9X/kTWFFYbxkYtCwKU6cTRGN+9VpZQXHQtb/FE
LAZ3UVvgHOS1ArYkbU6Bfym/1kjoDdtYYt7SkEo9rz+etdcGEVfyZEpPwcQEEO5K
NJZmIIGTDo+HE4TfGfO/O3h4Y9bwgRQZtZpS2/36Zj+WSNJ/ehJyie91XwpRph2w
hrYiT4CyPap41FjeItUdCOz+WtaQlzg7z7U82q2Tz1dd6gzXXGuVlJSe6C3Qz7Vf
nqH4K2d2HHKBB0vYoJKHH3A0sYXEStr6fDPr4rRRVFVyOTTUGVkD4Gu4U/jtv9Gp
h1XF+/L/r1c9Wtu6qNlssfBCzfCH2X04ltPxH2s7ZPqRxofYBzfCAanCpo7GML+5
R4EQn1Xf7QC+TkeP2HWQCGC9w9z6+QW7naeFKZDcJFGco1Y8hhSFFEokdWms1J8E
AQm23YDYJOHUstFzDHR5mnuAKjExusDrK11YIPdI1Tr4rPL0GS3WtFn43C4sYDQW
756YbhVmKo7fpOzKq3K4S3S7jOKMUTiNtzSfYc5vCMLFlcAl6upn47rWISom8aIs
9hSqPBtpYnLCphsSttUfYnWUGd0UjU6qylhz6pPDeDVkZC8+2SueH7fLU3VNi+r1
Q8hIarRdRE+o7rlPC0G6xAaG+uGlBqm2/LCr9jNqBwkZ+lD534hPF/uKT065G2+Q
quc5QFbrTDl49HWiUQDRYUKbsftjkOXnlGzWJrCZudQtE/y5iTjRNlPaZXpus5Oy
FtGmAm+BvhnYmYJY0gi1RCzQZ8NI4UevqgEGKjWrzmekbSy8dX/FVFyddNiV7Gnd
83l3QpF4HtxtiAmaSMPjJzn0m8LwI/KR421A355gZ86uZ6OcU8PG63dLxbJhZPx2
fOWjZf/AWc24gh28dauJF1zdQrnbzXl1u3Cn/+njLpgc25VkAdLUA18BS6LLw96z
0UykG4I1cUwOMbsbmcm5jxUCVThBLYlxMw6nzTB3gIWP212grBz6SP8tNHlnGxG4
hDlR8q+eNWTvBISz9MNyWhGKEOy+ogPOk6L/Rl8Tzf08RnOBNwVkN3IicaDiLZyd
PYof70y+z1O8PNYIKWfh9t1aoSxdvh2M0q4uzeaf5Rfjqpy4ODtFa0LsWNwLqmHa
02vIGY5z5PG+HXs90Aspdi6tXnp8lvK/iv+BmD9lR+564j/NnlksETz8GW0b5JLp
tWnYG0ppCw2X96UjtjCx9Kh9kt7TytkcyxT9GVD86YAGgUwyBVljEBneAuIGzBfA
afKAs1XspajniKeLyMfcbkC42JX11BjbbjOB6PWV8ymqmzdTryH7n4evABEjGs92
uAB1o/wZVEUjkmnlkdckXZLNbKeOKRE5T4eozuTZA/YDE+Aej0Kcf+C/Mqc7GjeA
oICHbFSPmbG80PR8TswG7/n8tF+MrMfDHPtHtO1iOdRxcExo2EjizD7SJJoJLMFO
YMAaWMMWP/dllhX0biUPYBplcx7RZgS11jti/qQ4jNdx3FsfhJJPLzy7LH5D1gjv
MsNz7PVVn1wBChE5+DrdSnKxEKSxgJJvaCjCQBIjzIPhNRbJLnE34oLAVTQogJKJ
pqDCHrFEbFlhuCH1ImJMBLYrm6vgqBqTUMMO2T94N5kIzpvYcip8Y2BWYxfqoe2N
w/OwFEeK1ueMWJ1ihBDIoqOfnwTTWjtGR3jfS9cJRzNVHA6MK8M7eA9sCuWqemry
Xq/OnLNcLsQSXfoRxjQzbu8NLdgTMTR29q0jakH/UwvzPNQSn2UTY08B6aLjwYrG
66SYO+OHH4PhbtCCb54F3/4hMWtc317DQnTOuF75m2wvwy763kMm+2sNd7LwgtmS
By7/OYEY0trfXSm8msoFeiXMeIGRvrSyNiuopE0geIkYclbuNoMRd9MLWp9QohFn
A30hX4bcSVLy1AgICEvVPw6f4Amw4UzHL7qIIue64wEoMP2mNHFkcYwsjCISMP4J
w8e2JzuH52X46mFDLcyOis5RLQucGxYRKwVEKz8v1k5bKDuCbP/oNCRHgPaJPZSO
rf87zTd4+Lovklq8qLclroRz0gyYLaZbJdQ4v+e3wZdGQGNUY/Isyk9xftpnXZiU
NqmhyFkLTUiOK5AY6HPoeO/TvmA92pKhT7yjOP9/0MNj4A+bXo25TrhFSfNFOauz
wwEBSUNlpoSExC3dTY+9Zb29TlHLN7M3qWuuEfHE6GQGDv5LxRIuJkz+Is19+ot2
nPLxTAPOI3JGy1eiPGk+pPI5rgZKMpybjah4g3V4MJ/FRhnVVdY8j91FTs5jWVjs
tQjStYioiUbfhgO2FIrWBDgvKA3bzuhqD3ltwjz9fHOheOY8V6WJ0T+Sqks00dW7
Rv+phht3Z1AHO8K8yhWEC1JedP2wRoeM/3bBb1qnhsLGux5O9T7S46iv4N4AVlRq
+Sda9dEPiVx5yL7egST0hu+gY/XEL0wxqWviggO6B66jMBLyvg/4K6hhp0P8QfQT
soMs72bAUp7vTQkqFrFlwTEqDJk/uNi4kojUVlCeHewOpl3Q/LE8FDtxvvchlRS7
AbcFkmJl4Yv/2Ahu6lyRaGtPtqmEs0CZNLNDRgqiRXjHXFXrgKrpX7KqR8377Eea
mWcwv6cYqY7yyJ1SRGaPHvULcrlU66kJwkPonfp/4pS3Es9sAhFZ7Q6kKqx/9wkU
e8G6bJt2cYwjBsNfo1byI678WvxjxroeIg3BkUBQETmGGKyRs5tR65TGF1knkpNw
u0UEvl5123104eWKmklBGeBibordbgX+KEgM27E1uhpFUpgJTVPssjg4WdyANWQt
K4TxEYXnSVTTgFYWwATDQSeFY5FxPacnSQoK15IJshl8QCZ6B2XO7/IO6xXqMh2E
H/F7cQBOn5i1EfiC+isp3XfGVBvWN+2TqvZFvFvuVSIfjiFaXwaKMD283OXKDJhN
OX05IG7d5TvR/8H/Jklvnxa435pFPelKTOmKHAZBv1TUKl79IrOjGkwYXmwFS9Y2
vL0JuIqbPo+eJ7xFNDr57zi73MMgvRPNJ+0VKaz80ek2u3YhEMet4HD4qYCEYDnl
F8NrRGI9O6jgTkR7Dbzcn75+bDQHT7H9IqXY5HOpWcxElc5NO+UrfYnEvVdGPHXb
kL2+iE+1gNsMitFctL7QRZpCRx5MvyibriZvZoXdwDqgbad99pJhFj7u+30aMhEF
CSbP0IQrVSXPYsohSjsPiJ2yFSBC52AvK7qnr+lYx+cu3DlxtSj57+4i+6FA8roy
a80ghnYn8FybNygW6+yyuZjZ/ahUlP8E+1EgjxE3ANu64b8rO+R/P1Uzwy/fo3ow
E5p8fMifaPVkBnsadbavz2E1+G4IPMCkCDqJvLK7V14TG+iTPPmMK6oCpfIZKaxn
Z5LA+koZbkSxNXx6fAb0Txf3cjwdipoNxqpT10ob12KNhDvhpeYrVGznUbRZ6gaf
7J442fDYIsPTfzxjHcoW8QjmLX+5lJ5YlZ7H/k2fOHLdcz0yfbFpa3Kqvwl9rnsq
zCS9yjeXoxx3+6tmscKbUHCB9w4geUG/slp/YoXMh3pdeOWcSdPolbmem7sueFl1
D1/br8MzJos63r+PvWq4T1Hv6NWRohCVMs/wOmvpL/HU4pSq+eJcNh5se4539MbK
76ysmV9+U/to15PJbkQ2tMYSVokNCBrYTXFGfQtHkqgnGYk4viWrucRJMB9l4Mgy
eqEji/EPceHsIsZ8/4HexZ7jPkS7Pv+cFIfKtdvb3gVr1fiks0Xua9WhOHcLWLOb
Ll7m8MkZxiR/sE5cPyte8CT9P4I9beErkZS343gabt1tgo6Demlo/G9mDF1Gq8Ti
18RaXazX8uipPz6VRW/rdgCxs1dkW7NsPaP4eOlKhSQHutqwG4C+ATFIJ1i1XBXU
3YcKiJDvBJJWSv2W+bxVqaCFWeRu78ViG7f2Ejzy98cfpF6it+oGe4zVytPU4N+o
rzd4XiCYM3is4zN5X1iUVOyNjivZqssoWXQAo5xkeySnaOBvF3AVoEGtfPIrya1E
9jZr7ks0XJKW05QPDR+y0mGdCeK5jNYHWeCwq9vzy2e3HsPnzdFh8DVi+DmU4Ami
b/ceFA4xPgmj5M2DoEYZ9PYwQ8sSRRtByrQr8ab/pYkTahpsg/3Hn8FgL9Dlo3BL
soCm3F7jJ/NoG8rwc+8wHgQ8C7qS4UIFwHZgTk0Xp406LQ0+nbMrkwDB12T+jT7z
zbj0Km+g7m8fcxqgJgJXR0PVbFV8rs6RXNBjmV3sIDhEGTzUezb0XFTlKB4txM5E
tzf+QClqWgwtFQzkJNBTu03MhaBjuT6OFDQFZ0ewjVvTZv0CUYVjxD68M0BJEk2w
yoXkDS48ujua9DyDiNEJ/e/PPIsYFdBWfc17RGNSw8lEoXjYn3MVBOsE2Gk4ZIcv
d9V4J0xQMJfe+pq9OirUKdeoRuOKNzD/7a/1ir2Hi6Ce87gtwUjNU4L8lcp/e/+D
ayFiyTnV3yJi96W/hCSSCp9Nl/NioO9qhxvx64xJkM1743ac0z33QCFJnHt7l1Bu
XBTyapGEwBOccBGtsdB2VGqmyPNfvZQ86Dz9ZqDCpVHJh29hjlg1RPAHnKd2Z9cE
b68VEP1atd8frKM/HMfvHUsfP1eTiyr0Sut1fmXdltfbxcjEv3ftRk49WD+KsIin
8uvLVA6qyEllaCgSaBWPr91AHTC9Rn0YZQ6p9OLV/9VwCtul3JwQmwegEFlQdMng
LKraBHAwGZOqJ15od4qWoLA3co8G+lNscpkCg1p/9VtyNWQ0euge4JhtKDI9GwbX
/g2ui5C6NsqBZs45BefQ3ROaol8On/wATZqx4R4oO/D14zGKVACPEWEVCfKZ9OFD
1TG3VBsS/ckSMG6rdiuuJ4V81KdMGNt7Lgj6Rq2tGTvfLoFEJldW+d4PcVvxKq5b
sLU5JJSHpa2QNh/RKpuLJKF2qQAqSoY+D+/Rm9yweU+77a0YpTYQfHB79wb55I7S
EcrAx5MR9y/YwBI4MywP/UFyUO82cEm7V0GSf1Cnc3q9wVLYAD8tA3izExIUVZDu
7aotvOPbDhmBuRAj2aONQzv6y1x56PR5hjomoMJUL9C4K7xkDPRgrrKd1C14jWAi
T+26/SV2RKZEG96JEh2RRFfD09Qbb74M4syLFnhb6X2cNj/9u1SqpOhmbkW2shql
T99/TPNgbSjUMPOh7JjVFz8c7ggjeb3Rv08j8pWKoS5GlsGb8w6OIKrQQB7VDEqd
hu8Bs+xo4utMwUEMBB6IRxZydCDcHVKBuiDQhZtrTRe3f4qXXls4kUX4Bs6L3atH
0WM+O19RxwJscLpAmWxS6qjjI961jIqcuedmz0mZGQvbdfYYdbg5M1768gtMRF0J
68IAQEm0TCE/aWHjlc15vXQsbbE8mkW5IB2U3oDMATPuxL3jVLUFqE9g51HB4Ny6
qqsi0ueMmyF5nPbjkCNhwNklY7edJVKOiD6EZKBQYljIAL5yVCNjMSAb8kVo/qcY
MMRIBADenQHyN3luh5qhx/6J1GDcanXEnvKosrJCxZjmmQMfqt5PoLYu+gwEmmDp
gy28BmP/6aKc+f4RGSjGO9a9a53Fq5cNhaXBeEaHROEOh/vEuw5D2xJC1YlQCFal
MxWYvKxRJLnaLd2115lnK3vc5HygHCBzCkOapryOV9jepJZ5zKxM2NEWdBTrPVWe
Fl+YAAP/5ffYzfQxf9dSkquDHQu2R+oOF7voUQFAJLOOIwV7RYESirPjL1rdRUq4
GmxA0YYgWFThD4uCAHhhFcOO0fUEpgKEsFaSecsKNCWqY+MFqvXXAj5/mmfj7T3c
e97KpNvzVF/KsOlExKpWPOegm+e0heYU7/LA7bhoX6hWjBEPgePt1QVz/1EGRvIT
3r2UO+uU+or5kcMRb6Pfu9mFIef0pmqcD5mLiytRlR2HwdkKtNz4tBwlZ2A8Nbz5
MvAa7Zml95qm03A9k5Gts5WKrInlI7zNhDNqTUxnosQhM0KIe84QslEBcBuKtWuF
WSEVYxulBHQMxBBS9VjcPIemLP3i8NzoMnYOyLgbRFyPeZWzdz5Ao2JPvF5MUQ1r
/WcOU1WnW25UDBrmtJEfTVksQd99BHPfhlVYXJwUm8Em2Op+IbNgKW6bEubtdKp5
hC3P3QK2iZAL8MaRePd3GtFrucqDM9PCTyduXqsOs7uuspO24xl6UOLYmX2YpcQ2
/r7Wpj71PnVDVC9wZec5Lsei8bdJhpVo2Eb47s6xJvpqdqg12gkmHvxBXBrzvwBh
SjS+RHKg3yikSQCUBccWBCEc1FuECyf1GdkmovJury2YH+qPjZthJuEpA4ocaxBX
BtROqEepBwia8Yfhdo0mv+sh2enBxVvae1Wp1Kp+7nYm7sRcMv2TuoFJz8+DwsWd
P/fK56cC+JQGPdZxCXiqeqLZ6QsCYn8yjJZugQXi086p4mvkecrsbpXIlP+XS+Sl
GfEftdAVcTS8VnkPGohfQsLj7+m7WC1HODpNSJrefp7MNWDZD1ZmFBjfKWpK4Wlo
Vv/kt+2cfkFfoNSV566iEvaq2MAemwiT2BYWSbKoj1wOWuus89KVeiBo402oIITB
vzxYvGJ8iOnLnCYoMXNEIHQ8WpaN9R11IB+Xy5iLWFPQfViXp10J5I59UeZ1qF0/
MEvL9Cq+Wo65ssylt00aVRF2dklNrHdX2XnnLryBd1whZLJz4iUzXWHamocsF5tW
j5s4InfOzLChRiqbarSx2/j0CqYW2qvdlPUZrQSVZRnrpC4o0sd+70kj/87IVJVw
9oLXL2Jz4st8KjfahH2xjCs3duh2slX76NFsce3CEN4JlBseXIgm/qaeUitxssRX
iCHSHfqNDF9oGu/AmFrUnytfLp6VP4qcUCSngsRwT6d3IZPNdRaNqcJcVNCCF+P4
KjFfMVm4MEfFkNs+ZnV+eBk6ywb/LdrOKrbOZRpi+hon44b+ztdpvdzKcxUqps9A
8MVYGxPAOf0Hw72GTZN5akF96HuO0fF+/nmViYVCnrcWL6mEEIQyAt92IJjbGmDX
yoTg0C/Ieopi5Wltkhc3ougpXPzw1O9EPLJlOcFu1poDgC7JmyQLNmuJmEBhY1VZ
tYL7CJTnhmpBciHEe5pQWZERM4bENXqHn0K8bgamLA1dk1OmV149TtzCNKerMzXQ
4zf+otWqbmEbo5iKUcfcSaMIKgwibafIVxt5BgBvIEZ8+qx/zu4A14PoroiWW5pL
1O9oLoxubpShCuV2xHU0pw4wtuIyvOeGOzbYruCn7+qFAPM9qypUtlXQEa8oMBab
DHDzckFINx48zPFAdZ517ngpfaVi8EtaObRZMmpxZKFZ+68GdN1rgGTe4vJfix+N
gGmDUC+W+ShI3zFbKc/ZJSLdCltHADpyBDUuX9Gl6IEqTLWh2x3N7ZGVUgJwLaEZ
mkmkfIu9fxe1OTSWuASzQAxAYhTu/sqSh8SaJD9bxnWfxywoX+dw6qF9tNyU4jvZ
l6EijRY1nLF8t/uf8i0IzNabukQ4DcNzaWyaeO6SNRmAzzVBzICNk1A6uOVrffDa
jNgdfi6G+78Li0+TfHK0ZFg9+JSh8WIn3BtOOv+9fQQzT2HScCTNjs8mTcLfy52p
QNtdactYFiewehlTOWp1fYc4RQ/a0WQWKzfbss5TVkHYjXKyohajy5Im+67Dk6wR
HSnx4hYgCrC12RBMk8xz0uGMMQDIWjzXsZ40VV0AkVlbKbM/ys6bmLFfC8miwNoS
5Bv75na9JsoUVHYEe2oqOY9lw6rdP04auP8FjVxo9Li+ifMt9ktzGOkf0YvHnvlc
vcIXgyvP041YUBruZfvi9J27G7EAbka/oAdggvfsrc/MS4EeSIJla5TuEs5m8jfJ
9ep1I4ictQ5l0CJvsrpJm3qtHsK2JmKfk50awSL3LgeOhj5DpA/iQ9RH5En9ScN8
rMmZJcMUpKzPk1b4evad047WPHIfcssQLmaffBbzRkSMmpQeg8ZvSIAz8q3Y9s9o
XV+kAIrDC4HixwcAWPNqnU7UyWRwCb1w1vEPy5oqVw6nOqUcihoAkKnahc7LxMK9
us/uWE8iN3ZxOoWu4aFwNlKQ2Pmc3d1zp490z0nhAftwleQYfzY4cviCMSpX/n5S
oecDL0VDVPmw5MWHVWNZm6jba5hMEx/8rsBE5u6O2ZSuh9/iLXhkYra4aTphfHMR
TEO3g4nCnH8ljmSXOP0RRUZ8Y2pJxCsQRDjzBl0VkPfr+hMm1bzRJlqDOUICdOgT
QYGXsQWnjSn3+qIP2CRXFNK9qoXiJMo8vcJzCOcnd8M19hm/3ndGoAl2tuRX+aN+
+iBzVF+TGvqTi3rGRhAOkCi/to3p95jrD3gyStODuKR6iv/GeVP6XnfYTwccDxlm
aG+RNDNGxfqJCuNdBTAII3wItSngrCHMIENcye1dwpTHDTYUvENGd7FVXhR/DX8Y
av7PwplxjmiS5XCvOT40+w4dBWa29yH9HFHmnrx/4JNJ3Q7uqykVbta7v3Yt/AGO
XFy2TnauAOxAHBo1hhU79e+o++RXeh45u1WHWtyR4ebcsKMINtoByqC8NYO3mEv8
DX1UlSY/4HMfAAQNpnnpMadms1QRYmgLDVxZwmbhCenYJdm6zOSXhqH7B6ap+tEG
MCPPOJ99tvKyhsFFOODDqK9SFzhXUzoXZUeuflZfoycSebwD1/yJz5L0OlK/h2Y/
D0JRUi2tgAi/jGpy6mNO+xApRmHJ0Nv+ZCLbS0aHiblHjnKA+JggtTFojZbV4l8Q
fXLrhTO/JDUTXR0knzWAlDR3iISSil90BdfYO+vHCfZNO4XP4dxy/NK/+PtDxwKI
sM3oITtkyUgu7VpQ+HLSB6WsY7gcg7V1VITLe7UwylHhoG6rWmYctaraPOycDe3U
aR3boYOqeFLDwictGBuiN2ZnNkUrN8D3aeUM9vpGpRlvIBeCU+io8LaeV4oqSErr
+mkMANxtVm2jbdM+M0HwF0LpeqtiLLNfKY7W5Whu/FyoCetrgCMt1a+Ecva5JrqV
5UbUGL3rCsNfZDhjciG0UBSo2PAEpjQuPOvn64VmgBi4QzURCt3AxZNmC4IyC2BQ
cHEO/QB8tXBLJy6v5+FM+km8CBYtgBxwtpFuCx3SzpDJtgcFGMdeyTfPMi9D7jtX
CvqjU8I4JS5n4SMxUx5KKZgZzmXcjbU08OQt66hHXZKvW6fMX5oDEVyjFJnhFfGO
aIUwr7jDlT2cG7uLyjBEEClA35HH8DQ+b1OIkj9hA6F2vqfrjaO3dY+dQcoPz/RV
taSvDjFWy9j1sxQYHSFEexjivAqnvKbQU2PaxhT5SvXdUL3beN/nIvWqd6UVeqF1
+ul0iIo6PzXpopYZ17Tbd2ZEWfHvd3LAM5BTi/rw1mfLQ6MzUs1dWVerbih8Yo85
znD3jnZduwH7mCMBSPNc+SFrNBqAhSAEEqqw4ffpC4oYrpxlhmXn/Lw+3uxJpZYq
XDOLJz1zPw7lvVdtw9MM5QS7qN3QW0FSnBiOq/hr9H9sxD3sKJGOt17O7IZtdPXp
XvWao2jfsqhXSQfZIs6yI07oK1b+1MdfzAldRW43/OkrpkocGbwyb7exjLCGa9Ho
FZMaX7p5m/MFBnFfvwbHbRllMLH1HDBb/yUWixwCcpRW6IKyir7kLsPXC6v9V2HA
8brqTc/XBredispIgYdtOsgNsDUyz9ejd/soRipeC1ULQBtUQ7pCd/13L875OkrK
U4uc5LGO2Js9xujk/EkUAh8VfG6VSfZe/bQxnf6bwFmizBSJ0njCEMnP2BjOn1oQ
I3W3qCEAxCPMHStvmCHQuMxsj4PFKgzLByYDMfnseFfC5YwJQh8HnLpvVIWfQK+j
ldIqvhUiWUVLu4KO88bapX/fKBFbMYtOYEDDgvlLdtGm4YKu8JUPzlTohwNkLUSz
/ZLqYleH6jjxZFxt5huIOzcB+5vQ1AHBrSGnwyEBkOSdQn4aQj18Y6/h7R6CqKiC
GEEtwSucOXQwtjL0Ep1v20/+yIUizVqI/6O+uRxrqMCExBJ6xaQcSRJ58yOogb3Q
adMB+2MXNpz007xSqHd9TRNlfiJ1FJDvp40ZuufJXVwffemOI5BsNb/mDnBwJoVK
sY5xuaiQDRX38UG70VtXDrsReDmdS39b3jUy1OpLJwBSpY+2acNlGKAeMqYDIkOr
PL4SNCvV5PZgu+qYBAPUsJ8JjYYH+fcH96KzIAFjGBogaHVLb6QEIxkMOhR7EBFV
o54Jpuo+VfMfIFBfa7LoX2flX+8lxxWhSIgrRtl/aJ8KUTPQGYU0oSeq+90C5ID3
8pzv1hyrwvSSqoQ71dDhtakM5zoxTciqrBbLOgVfJtegex/sftnKU9h4HsEguzTp
ge3wEEdJUVfM9GfRXWLi5+wcVdAg0pgEWi76Hm8uZgMqoe3v861OEuEOUsk8hdlk
ZZEzJgOmh1clYd86Av+K241f+AdWHzsFtlYxOZvXlKkqHoDRYOqj+KWHg7XRrMrk
wrcJa4+xKxMXXH93vzCmiLtMtqv8DpCYhd5wxJrMGkka5avmZIe+Nfx3qnWr5Cwj
nQcA53k9fe9e+1ex7j0Um/Lf95meCzrtW07xVG4utaVQ/Yaue9pIVvZG+i1X+37r
ROfNpmFZY8CzP5C75H7TOVOAY9XTam0hgsFwmdDC2BR+k+J/NBuTi9gIhPflS5NR
W6dS9iFc9qd6e4kqiroKAYIV8jQHONMt/3XfUOYjgdrlc6ah3CZF4t+DNeI9shvu
MrMxjL8zRyiO3pnXwHzriFlp6tSwBbMeDAhng8gec1AJOSvtxYQy5NBgtbjPIloO
ktlsI3k7qIvJ/nFYoTOubiTEUEZ786AR1YeEo7jtNQRGmExIDeRuSJaSTExBGYSQ
1FFhwa1jomJBTLxZ87pWf/kDlYwVpv1Roq94YFpjGuQY/1BfGcl5zTy+9nGwKniO
6aycpOPaaBMD1yb2aBx3djkaHgYLw6mhU+i0sYcjO8/SdR53EtfbDZSXvdILmmdR
pZyi69xhFAq+2mpQGd4trA/DGIbtRgH+4G5agZLMUW0ioP7uOcSY7JpbRtFML1Wp
82OP7YIF1D7wMFZBZ2tvqzYAOz0W10+cZ/Da5JAsRSqQzQB2vrQ1Wcmbs+Uq/V18
eooBj3MR7DrvtHW+A++5rFfZWtWGVc9b/ILLvkapnTfgLgLSjcl91a5fS4uQ9S3v
FfaXp7wx795tjEJrzCqt067qVSpaT4jUUWDmO0jFnJ8cmCoGa7qmBBxJjoxvyuEo
ETOlFm6fzXk1Yl8obrcpY8aVF8J6cnScR38pCNVETpwJbGkzxg24uarkqPCz/iIZ
VjdXFsKC4c++pV4ZWABQYqd3KKQNTrBBvYo17phh1B76FKCN26fpTLtZbjsEmEDW
ynsh0CNt6CS1txGGvde1gXq9gnmFeUpckyLzOgcHijA6TMTQh1lD4VZk+jaCJW0F
YTjESI/tIFYqR87onb2qgPN2eBG2uQi8D/fxml/revmI6j1l03oPZUjb4r9Oo1pe
uFsxSdOK8HN2zdbxiEjrJKR7xMki6f828s2XrqQM4Lc1PPVoAzZpajBb59Fg4Res
lXRL5WxiMGGyDzfXutdWufNM+LS4dDoakDNdLLfNhnFc+Q7yAkbVPGxunZbhodEU
7li6HerQCDjHjqK7sHNtDjwUyOBhRn4AfoGIMHuHfYGsiqj+ARo4FyJ98kzVQa1s
KN5kQev0RLQ3TmGENR4taASxX/JniXfrowP2rgCNd3cdqqb3Kwre1T6ox0hK/uLR
dw8TXq9ttBPdNmiUns4i9CC2PTSTlR4YOLaqqeooyf2HtI+2Z+ptwzAyJKveNJTs
gLt0Mxqm9WDyhZIagE9iEtczS/jvoCu6jGhCVP7ANJRIEvoxrdo9I9rQ1yE7dTZ9
sN542D2R3Yw7iPSWqTtchEX5ZcKXsaIm+flYysWu6Z/TcuGq6zhtGoAGi4rijglh
zTvuyg5YYFnBvxaMhQVzdt4rLIbhtgxZZ4blmeRRanRkSzokNkmvZ2hN59hQ6Lx8
55p9GmlKob14G3xgkt+q3AHQ6uv80oaDZ4jGZsex8GpSo62RiGCkL6N+WmShFQIa
cQKLhhXnLSsC6i80HBWRHcuqXPcCU1TOV2+Je/TkDO4RqfMMSMjXfz0qZgEyOlGq
+A0xTNaYbAxantayVoCZnECMIgtMdZAzp8nTxggF2CuJKVzRPvW8n5/VFgvhJRlV
EzgEc0xoM7LyG2nnLoNbOYGEWuEikt1AzKPFJE8kzkPjHPphuafv8J678Sj/nuC1
eypx5u8h2tm5dzUxOB59hOQA547tl/TrvaVlfTy/8cIhBTO6HOqzLT0BHVQvFUR8
g6ociom2QQVt3uuid8IpR9iklUHowDgomefnExtARB5Mj0PKI5+i5NI5jVReYuez
CAs467feam8i0mzKh4mYv5CVQcYjPvDTMITrTjDIhQrKpHW8RfLRn113kwTjs0Qb
pVTxUYyY0c4iiRlyY6HqFlHKYVYHxdShyVovwamZnxkCQqWTqTrtoJ43hgCOkR1Y
3Lvc2+Ot/G1ia4ARXPLtggPpVFL6IVTWjEWb/JferGeEuzSUMBba3TgbC9TZrVxs
o8l6D95VHXck6V9qM1udi6umDaiqa3GdCKQ5bWA+kpg0AoKKV40FV+tXwAFpQZ3z
zALHMZxMkc1+K8rGUAJaz2pPKJQo8O5YuittCZJXNK9jsvdE71HpJhVSOJVFjsPX
19VgbTp01Y07JC/yPgLC5HBAQEV29xxDfE7YaFRN87Wm4JZ1gYHYriDwm3Fep4W/
vQmHr+HpvlhCs43S/4Jamd4tdIgtzBbtWXUVgLNDatDxX3D/4NrZ7FwciqKqhmeR
wHSxi5FRL7tIr+5Y1qtexWRaYUXlryvH5Dke83EFuI2Dk2dgqmL/gmozO839MJeC
bZMOnCXkbW73AfQ8OvxPl6lcsrVXuctue+w1e6SQhqD7NFn38orCzHX/DfKuSVDL
AILchduN87hW5q1Ja4XRfSQBInNVLLBkv6D4E3xg35WKIrMq11xaHGP3eFuJen48
Jm3d09k7Mf3fVaYhVATwAWqIO2Geg5fCoGZx0+YC4gPEtJJeFRKo0tjwooNhXD5h
qWgMs2du1vzfyfQy/VYMqurDWTr7AqQyhih6IjPgcadv+ATpH8ym6hqMbbHaQ2Ei
zDfrRU511BYp0a078/LIxaDCyNtgjyLP71V6X+Fva3w1dyjLr6txbGKeAuqb+I0d
0pcCVCqd5gGOu5affNq6w76KRMkLuLLcaCwwkPTOAnpF8CYCQBfPaRZ1SNVqpuc1
2TXRm2EErEVv53NDEgQQTMNLpni9H+m+e3ujcS7Uj+Nzokebrwa691qu8PVV34ae
G3nqFspMR58kq3x6dUeAlCqO78j4BSHNgsMahFdY9nOpCiEEP5E8IaTu598oSPse
kbc2GSqApXJw530NzP/P0njXs4+qtAnKAW0CEOZ0QjDC4SPu9sYm760HRcxTE1x3
7evABP6pMUz0nyoxF1nahzQpkiaEY1vgmoXdYXy5lyYcOJ1E2n25Bo+CWipbc0+G
vdPegdUgHxfw3/9oDmX0shGw9WlX89QW1PC/bCwDbysICly+e9Q92qPsafJv4bwV
xlCKnkVGy2cXprikRpzoVoKwaQfFt4vhT6oizz2tX+fpwxym9u3MsOC1zBWZB1QD
0JVWd6gyX2+QnW7xibkyrZhY3Tk6ZbhVdRLHkvH/LuzCxqfwrBqIgJxfcOsf0XKi
lf/gLb8EP/sRzacLM8I1ahIShdtfh0Tvwg3RDV3ht0mc/d3ZIJJR4srv+9PdttOs
rPnE6+/HxceennndJEwqPwIuSUksxz56bv4PZw0wYX5Y+TsQRIJzBNz80lagSPQQ
Klx9sfMIdSJu1ns6ml93f6z1o6+bM+guNevC1aZv7NGbFdgZ7wqYwimI5Dw+sIPt
G09mBEOlns9S4/mMyuYE1jOVEJvNcGOTTH3YXGrakeR1gW0WRNAKwcpln77WPY9F
he3Qe5kisIjUAsgCGhRy1iWkfLgU7S+pfuNdRgcaFdKFCPDBj7YbnSUYupYmu9O2
jW1B4uwxPX7+5TzaEX7dmnEHvyvqtmxeFNfChyiQKG9k+WQGm70vJWEkkyPzng00
T7Ai3eSS9ylsxlam9nNX+o/hSc5yt3KB11I3RbU0xR1ZnpSbMdyfXArfyEZpJqz1
KDV9eAlhPbNV1HELW98CnQX0ecrwgLStZ+jHd8eolFGxikxJexvQ0dD7pTM7EZ4O
W/WVj435yqw8PhUcVoUNbl3sTLVW/Dd94zYuRmbgtr4Wuqm6aJ90pN02P50M9xS7
01XtxarqZep34wzCVtR/qLS1/bShIhCqR6EZqgNSZHvRhyiY2EQPIHvZlD3aZedg
2PD/KTr2+2ZpuBy6Iz7BBX9hmHG6Aq6jkIBe0dFsns18Wq7j60zSZA1eiOkZEstK
DVmdG8UbTFePrvvX7FeJgp6xzI7AfoYAIg1svKLdRy1kfhDozOB0TyeGB5HVGo/B
1DkK9vwkXbK+VyCBnCo8kvVmG+scSFeHzQP8n+Z/RxhQhGQgG4j/yY21DUD1HnXY
Oj6aVCMI4CpXxCm5748YGVwCJQsg08vhZMdruDloIp1LQCNOyZjcQjvjWAuaoTKW
9JOo8m0MgpmrcVn7FAtZWNe8i9oEin+xmQj299flTNS3sgUbG0CZ3ybC/rZ4Uk+E
dTFvmmctB9n5Q8UM+6fRthJHurJtCE5x+VHpwevPr8NiaNmubO0GSk8v+w/OhO9a
T83AglzP9lyXZ0ri9k683bZSc4plrerjXbE69qKrdtjT3dxekPGHOFrpc2klh8Jq
lAId0e+RVChDZSqNvW3Dw0NXHHuAV0Mctm2QSxQ8VBTb8IYqlEHQybJM+gmsNiuA
djhWjdyOmKA1oPRTaw8haA42Lq5zAoH/PKe+uEZJMcJHohqqTHnPIALzxyK6Zq8V
Av2617ZJ9RW3p68LvIazeQJLFJiEmkAxZ5JPdT0dq+LslavlA2UjilkaWTVk6WkF
zIo0wXtpu8wPF1DPKwT/ZT7WMJmC56iN6k+VmhEtLH7VDyveRMmrBQR8MxT0EvsT
4X53VMzyJ0BA+ogctf3D69l/Z9FfoNU6Rutn4tYKnrhH2SlBQxfgVTvbozJMIgDW
VCYI88ZVf0CzPMLsHQbu8Vb+KVINsH1eTmfchmGJfuAcJTbmdeR/P9ptiLTa+yUC
4ajzv0abB9T0GzeHYYOpKk9xqahOGal5tGy7gzBJLRB2CjBJpile3Ieb+PI/i0a6
IUh3whAKev++Bq7DpdzrUJirWTeTyBksnbvlOMEY1BRZO9n9wYv26d6e6xrjTmuT
0ZVBap1a4GenZ9cwm5iLGhqu6wrMS5ZpSZ+hopOFh9qdqnvb8K2weXZwjZs7s4AT
Ty8riAa+LHRgDgbUc6AGj2coiZ09oDNBzrOSGvZ1sjzFZLO6J7Lvu98aYWoOhhWr
KWQtpDZNsQips89pFQXGdp1F7/ptIW3JSIDbUAda6UjxGu1bRNR0DcsAyPAIuiz0
u2oCSjnDNngDX0crFr+s1JirB/EydZi3gJmKOn7BKXnRc9ffwYX4GowleURIb1RO
yZAOZeqJwWpFb36Ye7x8GOxtG6OvR1RmJn7/VYD8B2l384uo58apbbFYqjC6iiDE
aLeOKXjnQlCcH7Dn+mr+MxuCEF9GHWVwud5yKRbloNltMTIDVxbWgBodWLVRhor/
/U3Xc/DHmUBXS+9fP7l5POmuCUVk0RMOKa6IiP3hPw3P+12gnBb3YgeQCUFGUbMy
ahYDbGsddhtx4CdeO3yxCWxlxummFnMgF1k3ZNfs44m2t9cmnVRWYhwfVFbacJQy
l13i+H3zhCOwr3rvBk7XzKPobWkA+9o92UPbvfqKYeGLecaDtkbQ6b0zjlMXBdrp
71V8qNYSq+AfvILTD1WdgPcYtq5BxnDI3pBStxIKF1qZ+xnhSUBcyGGQ9qR6MkUr
cGu3FwplI2+HG2oop9i+IQzgUJdOFd+ehVqg7hIJITDElfDJInSGslGhg1j8pngE
tpuo8bcfU9fVNn1BQQd3nKYaszbnjCV1g7hM9tGT1MlIJ2n7rHPcPkpn10P6Qe9t
uHJBl4UuAy4zsYKI7f0qw5CRfn++WsXGbA/MYqUOYl1oDJM6OuZ3holF5+dT0fC+
Bu9CMrQJl0vZZ2oTNGlFSEOGgJqdiNgdg+49pNeE7si2AW7nZpmvgNHLtSjhXM3e
AGmm2UrGJ9Q/920R4I5Novwbl2sTqNy6ubJ3/hmZMCFJdSxv1PHDBIPjGAAV5aAS
LgfxgyuxYIXRHXEzbAup8be1N3KUGM0rE/oKvMKWJc87ngYKxHo4P5r2CD40Sfiw
dZ/hg/hATm0ni41IfGhxUqZL/kmS11iG82j5MUuKQhcPw2/8bh8wCqFbGg/bmjnJ
YzgyBopF825rrrNydVb7ia4Q0AOoH5/SXxReFy1+HWw4Q+R+20L5NyS4v+NSwUXH
qKqYt7kAGhYepL4fCoahP3DSJN9hvz04t0lX643Hz0K6U3cI8iljaZrjLLmOx+i8
zknYhZz3MnMSs/+ZuVR+k/oKGhIKClFb2PEGbWJjyVU5yxMrP9HuH4XpLTfdrIKa
hObYdVOcIZ5r8GrsUVPJbjuJKU0lPSilKnGCJbNNE/ENt8WRcSHXHaxUo4v1rwpI
+R8u8fOlUsBVdcPKHxaBc2XA5GMrIjeTlGiPHJDhAGoGMe4nDrPkm7MOWfA55PyL
tKkgsRC6uiSicyjkBK4uFLGH1d0/IoZPTtAxYbET99zzGYOu94SHyKNjIFPMJ2k8
+VyVErlKHUUheDF+5G9gp3zwSBsEFBdw6ALQ8wOowOQfnJonWHNF03gcaz4QBjIj
pr7j8u3/bbeQi8UXFwY4HyKMVog5iGQoadtCgtrQxVtIP/527C7qEFrokCzV+3Lq
lsQz9PRiuYET5Dsx/lyZRJO5h3Mwac0I5teteIVXtb2wJC+XFgeYNu/Rd36PLPmG
sYaU3W0psw1IZKKn1eEub47noVQ6YzcplEYDKA2aENlNAWLJXq1OkF/5mgUsZWW8
0MQXPmWYlCY2GxLaaAQcx0t5cYiy9vV7HxO9mmnHnE7IpobQGTouo0pUZbLsMmjv
KdsSqpPglFx1AA5w1pCCat/fKjU5DkOJulKz4x+PooCawh20tGWPGjec/i3eJCae
Z2UG4R2ksIQLCgfJspsayoC6YwrSjFsbp6n9PwTnU0sRSOzbwBAVd3kShXrIWxd7
UrQdBCmeul3h2/OfFKSfVlkQE902aGLQdGbfJpDSAUVxVrSJh0MN+WEEqO4Vjac7
0nwEipY8r0tWDsh7Izx/uxct2VjO0rJQoeGXAbXmmG3Dtlwgy/QxB5EaoPFTpbMx
FUQl72s5i8BHvJeAm13oN2Px1iF9mkut6TTQemxeOWK/u11tZlqZnxPSaUWgyYjp
wg1Z2liUOa5DtJk9ds8qGeXdHxYa1Ld8PWHJ1bkkbmqGamKOvZGldD7CjBzq4B3k
05scRtbWvOjBusZFYojhtwXVVY1rF8qJ2wb0zX3oZmzNDqZH0JFTW+jaayP55Ewo
6to5bG6KxQEGFVVG0MHC6SQbe9Dt92oes02zzRl/Far/vswBmOxGd0Y+JLg7F+x5
fETkoh6d2KZ6ao/axypfGC8hMLRJT64LgZOsGHZ/Oj2wAm/T558VfdSssfHMlU6J
tIUvwdTUA0UjqkYOuBatbFYK+M6Vzzdpxn18CBRQ6Dsm4kZqit8sRZjrfmwN0O5S
vi5PSkHZi3E74M8GrE/9Gk7aPuD72r4LdA3l8Vv21314czhpSfaj1KEAGp2m+KcA
tgWzF+YuYnBh3xVtgPNdXIVBqcgRY9a1aFBtWHhHa8jUVfrkCvpf4Grm7KMlwLsc
j+WbvjZT5llQvBnXGc+BlOZ3WfEmR6fN1W4PJ0E+5O/oqwDJ+UwhNheT8WTfx4I1
Imslry87RQCs/9Oulpe79AuXvHHeBJM17DBRlFBrjT/LH1qvXbV93AZErJm2MYZy
29gKWBEX6dJfWhCjh505wAzzwzQQyfKKm5oD4lsdAro6K9vcsQqoaZvPPpg4OrV2
9Y0Hwcu/UetpDoYobl6NqZvxlt/ngK2QpZnLcK+iEizCAGPWSc+71PxgeZu5eSkD
QtYWqebJwhmsLicUY7DOPTr28citWz4G064fq4lAY7CFQ0naR19fbbfKKpf299dX
385AEqWERGupZ5g7VXa0SzCrRYhWyw2FAaE4comIBduF6adIKreNe+qa/fu95y1W
EL/1+Ft5xa3MZPcarPt+ZVfUOF+rb+GHY/+T/IRSIqIV56221bnVv2BUHIIrihaA
yxm0+FLZGhaCq5+cH9bHHK7bLSDdqox7jglTgimgqkfRxpRIRAnEMdQG+rii4fGC
nigdNU8sySx108EbcOW0ebNtRU8eLrPRyRyWySa2krJKdaAGI25s5PlzrlRRNXik
s4DjgOcxIwdhoRRL0qXJQZ25uHX+9jsb6n4TJLlQjhbndpT9ePqMLZc+dm4ZGw+G
5LjF9HEqsm237zzG6Tuywu+reQ/iMFvanidp5Bni+AecCaDQZMrBe3kchSNRfGZr
RlPFft+7qk1XoPBJoFZuEfFxuBstAkJQQq6m0uiGOCjyB4LEBrtJtbK9R/gU3KCS
E5kvdNa0Gwk/Yf00oohMcu1FqaZRdB+SWEOjrAQodP9/G7BBLwzCnBFnp/QuaaBe
SfMt4sx4uQZL3DWVxHQpzA20kg2RdJZ1iPyPxlQhXy2si58ZQ7wod2l4wj1ub/fK
s78qajnfBIJw2VAcAWd0NLhH1YQbon6vDaLZnPmgyDloK7ym8OGXm77MNbvHAmpY
BsWtcqcpU0xvyhunt3kYAa2+ktDthFvwNxmlHWz1siK4RxNpjZGUg+u0QGbciBMG
w6m+gRSwiEGkzfMvxCr78ZztbQ1mU5h2TAv1NtVqGifj01Z6aft1jomdHh4B56IF
NX4N55IQF1PRiF77G2z2OL8RKz4Q8CTvdRe5A9kLK3NrvdfJBAtbvGxFahO+m2gZ
fFrls+8KSZn0YdcqJ1u8RJbn5uMeoA4PDk3sEjl/gKfI78dAPtjLfYtMSJp+PtW7
WmNjEuJgLFCRFQQYmQFEdCxoC08gGySFI2wmIxaDcJD0vMnF3pSPf8FrPNNekQKF
NJ5GroUsPthjceKc+96TOQNXrGQPC6uFMOuyIhTN36Rs1IIhDCK9rHLX1o2n954X
3lUNO1KZGauOvf5ltxnaHBl41w8X5ZToifhSS/GMO4n1oejkDCt2DBdqWyvzAHLz
3WBcAWUY699GfYbpqBsbQprg6ILl39qtvZemCRgm4N3VxmCmUBbNBftK/BQmJqil
El0AX4MvPZ+Ynd/G8e9kT3hcO/DviRuxTWgCZ5vLggZkgPWZkdxyoCguuh4evWWq
pHniwOdzQ+3xNYLSOJfkiM3TYwwT6sR2IkwugT5+3sM/I9SRmukQrPGuAyGAACLz
7bPcJ0ukYcRMDa8q+cOcREolDEoOTP2jlqEoxAnNz8Lho1wFGPLv52G8qynVmRqs
7ar+imaqVVBAvD+V+2M0r77toLFd3MfTObnYYV8TkgI63THNXPcqxCeVBaDcWLNx
nmAIrR7NnNYutX80aytPPwixH9YmvjZ95oFJ26SPuGvuxohDDfiFGlLc+XUhBegY
LHY0NQNl9/uE1y8PHuKwG1C17ih6zrVgcjBOziPTeb3nPXS3/qHvPt3Z+SS5bn4p
K8VNVgPTlpakFO0AxxuM6MnxFCd8SPXNLFdHgcCDeRdaTOzQTCYY11MW4lbFwW9B
RVB2j1Ccn6C42VngIJNN5YI+kHPNa97oBXVlF4wUOtzrktCAhr234yqt6Mk/PhMY
C5DWCTG/kmC5EqmUB+sH9TokbBheK+R1DXZp4q33SnMxCVw+H1nWLVtCsX2v5aT+
8BRtKayeXZVc2q5iPZm4HgI4nozjB8APVlwQVDJjhlZnzzKNHuLfOSYibs8zpXDe
8HOxT/ifRxDf7Gje3zCp7rjzp/2ENx3HiInV/FN83cTcCfHDdZBdgHJVvSCsk97A
Rkl/+HbOuATMpjnW1+7qr96pEcQdkLo/oacdO5SP0CAn0dCGIaXNx0dqD12Zrr55
7vWQDTJ4ob4pH/CYH9V6zC5h/Y1XOvw2d6zUdKDGbAQ6XiRW25tr5/+XGDS4j5Cb
5CAKSxfo+O8X+XNmczlgiNQoX8pq7epaL1YYHD6laGfbUxs77gATgVpIZK7Q0VRA
GXKgoBtGEtrD/Dq57Uwx6OnImXY83oxgVnurmpIZnOaZC+EHmjDAdy/G5Hq+y8xW
7Z8mnarfMEdh42+2cjpc+xqj2rol0aaWQokn4Cg+I51hdpPg8AuYI3AhDJDFIcL8
CdRPKE94PwhaHqjGZLSPNfENKPOyzcpWjmWQ/ouhyWDkFq2617VxOy+oTUmcz3JD
S+c8YuwvR35rKUxum9saFNlZybr5IJSzqGqIbFlfOBh6cmWyCi28B9ZngW+n9Mfn
obL3mF9eKcbCqUeiRuTizZCWinE2MEo9pyItY2dTM7Ha19e8snRT0zBJFGLw1NZ7
DkQR0nfuRYlAP7IoV1iFMx5DOdeSuXiDT0vc/l2nYLXLarUcJkdIRizY+IMk+l1Z
`protect END_PROTECTED
