`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
81j0IM6g/Sgpblm27TOoyKQxndByw5Q0RwMwXxXqCqryiYDScfz4qLl46LeZtJsU
AyF3LkQYd6I+LK38biVBLvXLDDBiEqKXCkw68nU+iUEwgMs74+mjAVEs4w4/Ad1z
/I5+vugb3k0KFfYI3KO1v7q7/rZl1ypEkIWDHyt1+KJdD0VUgyrgApxd42MSH/LQ
kIAlqVpLDFZWv1I/vmEcZKb82/KspV1P+Pv8xjmUrZphSg9N30n5+6b5/QTwDmlR
THs/o9e7hQpJ8KRQAp7JP6bR6m5HMa2m1jKEvCl9sEwOzGn4b+hmytKx4dl/rz2Q
WGr6ZYXsoiSw4Crq0FDM2tt9QuUqFRSoh76/Nhg0Mvt6hAkcPfzM7a5ObylCPPP2
nDaQACHwpY23vgbjUep9SjeWS/AzdNxKa7xVLr1SgY76TR6wEFRE2usPhxQFW9O9
AVYGJlnoTvVBdw54DaU1QQ/+HY5K0LDwE/faSE49Lde3bL55YS0VsApjFk+O1cqU
d9nyu7r2lnzOgUz+E5X7SjjkIC+X6uaessYadoyw2erxsVG8ylR9rnKmUAoqx3Ot
iF210QgQxQwBQSWqDoBdVev8XYiSaJfTGeY0MZ95jOsSPDUu6G6zx/V+z119EV9Z
YuhairoY+aeIqOL9DYbCEo64254PrV2CwAVwliWCD+cj21RktwWTjC1s/7s0OzdE
7xeRkrAUTw6OnKy7fiPA61OsEEgK6OV6uvZzR6JEUeZOByJuEOZvIrs6tHrVpjIU
3kNlgkO5csppiMKgoPe1GeOBbfwXwro0aZUdBM101b2zG+eKotSbCbOcv3kqQTOt
/x+tFAKTY2If3w/grAgz+p9SQd54M0ChaAN0zOwFodk=
`protect END_PROTECTED
