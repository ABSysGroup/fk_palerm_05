`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kUFgwHlw3fmS9vs7AB2rrMJpVM0rsI1EPCl7ng5MTkYFA7fbs1mjBmAHcRYgJmo4
dZcnIBvRiUSnRPC1amNZfudiNDlcTiIVYlx5wV9WkPyUu1EEmBrSHalEs5ZvvViO
exARfxYKeKkutZz/gXraW/C0oDSK3LxLtq63nTsXL+GJFD8rPLCuF9ZBxleWFE0g
fmdzpVi3w59vlM9WKMV9hTzvcUPN5+XsCQRE4IpXsx4kGQ/7Ce8yya7y+JIWr6I5
Wt9KQHpWR3CwovM8U0P7MX05end092mRKj/LVextoGGRhBpFMars19XV7YvK+f3n
C81pR8FiTFCfV5SD5Btv/7uPu6cpiSMei9EL24Geuv3ibvn5kudvfp9WeY1tyLRS
XPLr7DHrbuuGfbWospYUBtO6gEXtb/8PXWkMqYNCZG3jg6+5DOTh2UDQf+9IMpR4
xhAJ3h72L1bk+7iO/gd7UXSgpu3UuD1oU4M0a5ZBX3r2ADdtoKXKZheG/qii9SPQ
gfnB1X6J4UEIQcy+EGQmRl4gD8p4vUXlS8Symw4Peaiy+rnVa6XCWKQr5GINEVjc
ieL4QR+uINIRmXONs4WpB0nVJbEPokFZPt/i+K0IFBEVWhr6RsQDIaRNMEqUOMM8
P1vH01r/xD5Q6F0HZ6AtYbObAQvu+Q9yz15AVfxn9vT2GomC6fmPzp2ymL0zcGnV
HNWz5w8HCb+zEOoQisscbrnwkzkAfGrRDUZM3mCVEg9wZUNV7sn7m1eVXDpU233b
InHF6aMjud5itcGRVTR+MM9DrENZPHgCcZtjSeMUrbCc1Ou/D2DwwFll1oj92RK1
9rZYROy+vAK7v1ia5EFVe9+yuhANNqPqccHHyv9/z8e3CuV8i19ESeQxwzZwoXRQ
1Ku4ljU47oP44csgClJ9u6vJQ+X/wi49GCjY/ElJDQXN7CbnS5wM9RYpC5N6kXMH
Cak7bxrxtLbS7LGKKt1Zqn+9zI51yzrRiRC1CUuyqiCDXD9TSoPSnIWcJ7uaXg9d
izmAXzU0ahhL46gBtWbBClayqDnGD+NQEKAwO3+be81FXSz1mrUcTdpGagQiqaBN
AxYh8Z5JiFmSLHd6yakPS9k/WmdnDlCfDV5zKoi7xNg/ZdRoHVcQeuZvMjfHqdUC
AjN2ujElSuow3DGcfknOi2S9CvQQTuhVXDXW79Pb8hQEH72NMRIPgZBlb3ol/aeg
+LTmmmcTZLo2XxF583j2tiTuSuVUh7IdJwJ6peWs/1kk1iYgXgw12w1EYNXGwfTA
1jRD8L1GHMiC5fxBKz3ofAGGBEpc8/Q2/kgqB75okgapA8BMdHyJ/ONlgr3frhfl
bUnHXcrVBozBuCGKBxyGSAgoa4gdhCcks2ASd9er1fadLrMoLEsvXGWJxr8cUUdb
3at1kHyCdAFHXTQgPJGXBFl20VTI4NMnq+ACjEl6AL+/vmZ5Uw0Ke9Gb4MzsEuzs
bfQUSLw+VNYFDEQslrWt5WTEjcTlBESYawTKqOmqP5p1cwC0+FFLc3Romo/sxWtl
5IL45lAvZS5Gpp0vEeOQA56wdadIQZ/if9sNMXjpwuPReDMTDndHmd1TP3p2yxDb
6dIZmd1gn+WYExIQasS6+qBu2mAAZIGQ3GDCgP/XXHC8B+qytdfKcmnk/5lpPiAA
KfJlw8BXdcp1eidviQpUdYDDneJoPVekJPq8lNqlfEsx4zhUW40xbwC0bFGt3+Gh
Sci+OM9KR0tkQCucS2kJNmXKf18+2BisKfh1VGjzv5U2A9sNK9bPdGej1fu4h5i1
xvEg1+MAKldocYqZ8O2lm/PnrmUZPiS4zq23rLfRCvxYGxBPc93+B/ssP+nPTFI9
PNPlFvegJDcN8s5+aPfFbfASOA6OgvOUBYUMYiwCMfI=
`protect END_PROTECTED
