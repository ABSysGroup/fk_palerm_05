`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WapSJ6PvJEUuyGkWO7ZZpNxQXFbEOoBaBEhr+KEPnBT81Yx3lwB39/IIX+dEiLmJ
w7npwam8TyKYWQBgbXs8RYvGFmimTfrp17xtMSc6/ajxUAXU/f+fVdZ1sJlitZA1
reem5V/zPE8wwK2hWwUUvAWo0IHksX1jgbeO090l0tODPwTl4UZjCvkeNSxvFjA3
1+cDwuIDXx27r9Vbpxj2yMlX5Ic+Ryw7cMfrOqIUmv8TnNIH6/GTf0lhEMtYiYcu
xryafNhws4ZMgFtwnIFV3HZoKHML+ngUH1eo2F0FDtIm+V8RAya+YMDh9hi2OT+C
pftySXoxIpMz/RJgOPPOGQ==
`protect END_PROTECTED
