`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ACjsHKR69Um3eUiKAHw29s/hvXCkOav4bU1azI0CIUb/ugibWRldO2Mrqt0knf6m
W19vUoDixsZ/VmA+5ZS/S1kkWSc7Nx5OGPqDsMmHK+aUuK/m2iebXgtoPrJCTEfR
Ae6UdOGGPXdzt4jPJOP0PGBtLQNNeCNSs9SW1LPj595hokVh4q2+4A7etNOux3bk
89dMYeJVI+CUwPI7VM70gA0Y48UJedZIaSTqyVc6toTXVp4fZzDWUKQ7kq7IX27S
NXEvM/i8H4ASUxqonB33O/a+aE+aIyLs1WkIJQJu8SeYa4Rx4IUhysQ52fcOyBgc
2KQ8Ly/GYUB6qjgZqy0G6T72I2x6iov20XX+SN7bvaGP45UtLaNODVhQnZ2FgEcC
V1fVmAeoZAPmscOz1LmIc62wks6IzJtKEJNRsm586BVZFYIMTPMXnxqF8CFlMwVp
bIaLWvoHk2E893EUkRKfccxL28Bl958pQCRL8rvZsF4=
`protect END_PROTECTED
