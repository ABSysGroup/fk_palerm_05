`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8j1ah9AO+4+PAUCSB3tAuMQrxrY3HLxYIbx8NxqFRpa60Pt3BLHc0BWJ3vgJvccW
m85C1jwH/krOsthDoNvfKgKBkb9C2eBz8Q/YJVByvbNNcxxpt4nooInJaymeZ/ff
GyVDZtLMybzkVYiGWpa2xmy1OE/H8OhcH04oiiEKXCRBXWP0PZCn1yeKT4VGxA31
RUC69P3+AhAYeDdKNWEadpH5FNj+dhWsLteF104bn4NB50iBkbqcxM/Tr7YrhFBE
9Xho1kpEO+SyevD9WhhSE5q0IMcVZkUlnIqyCN3ZUOzurUcm9wR4ryeYLywfki99
gDUoCfgs+wxjTALrMIqkxcnvWuvh3ro+fRMi47646J/IunIN74TF0ntvReeM8kvV
k6uw77m7pQSBiXiYWqjtunM2sXpiTJ69Q2M8CLZr/SUqsmhUHj8T1jTL5BL3GOE6
GILpXA1Fn+TA3oZcVndTS0UegfziRfEN1g3tpW6yosqw7fECg3orRfJqN1lUVjdR
h+N4O3bugLBnn7PmCEErV3eLyMiJj4YiuWedvvXnbzjb/ryRLiBkqqFChDkd81kU
5r2BGjWyy/hC40oBQSN08TqoNFVGbPN0VouaIezQVbw=
`protect END_PROTECTED
