`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4mvw7B5+e2rekhLQ3jMHVfg7LbznFIGvdrPScLQLHBgXw2K8NV2EIj3tiaWXeAUv
tghK+P1YWVqMgfhrIAhYNQokvwhOtUOVP2V9YbAn33a9Tx/F4OWMbCoVO4KSDs7m
G+tgFl04+i1q7CeWEeW7nVm9VSlXGuHywB5yQ131n3syi9KVwiPhEmsxRsf/amEW
Ao9ZGlGK5oTKRlF2BdMEGfDWq7F3lvY3HUL2HKklU0eV6yjLDCR4J1HArvJXxhI3
NlctVkORJ4f1LMYgqSLR7xJCoPNpi1xbzIfnZTN8/ZWqeVxiPjl0Fj1bWP68DD0E
SwOBND3Ns+QIfHHbJ6K2QGHYkJPN1sAGDVwysxDUYc6bMfdZDM2l7ubo/wDxyBL7
mi9uYGbh5H8nJ9ODnAJG59ZmdpxYvr4OJyuNsOQNMUJlziyklG8BAWxF8fkgobWP
GaTuPG8b9zhVuJtFEj9D/vMZ+iNm/si8LqLkn7oEzQiilxND27YA8fqU2lMRi5z2
Sm/2WdewwWLMGcAJQxdUrfTxzSWadlGHKMqfg0S+7I6Z3ycKPS+B27g7FjVp3h9U
rDwpm9kXw+mOrsGDBZXv7cFhG1WZCmu0JmItBlNHWZFA3OOzP8C1nzQV48bcQcrr
NWd61OoozHwiJketOyipxjQvXt0xZZpn9jPGQO6v+p9xcJG7Jh1G4qC6OMFjXzaJ
uBKRXQf9etgFSm5tTmMcXo+cUEjqgyn7av+UTX0+L5jGHpNSjjvzGDKLUfxjlG7y
pR2jXfJM8bzUEmzBKE5JBw==
`protect END_PROTECTED
