`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FKRVkUPyj3HcH0qzq3S8/5s7vU8JZN2RWUILV4EWCmypsSeryiqPczeS6aj23YBi
3SIp8deheARGD8HRjhMv9q9yxUKV1je9OZ/cVSyiSW1jejzOYLbjLV18pXpZacAv
N8BggaGPH907JmU/6Y/eHWsFusNOQydyXYOrR4941ceOv2rDap62MwwqE1Cjx1eb
q4iouiWqHG/31RmW0GBZ3dSzxwcph3zgq2kgcQuu5KN2qAyySW/5e2joYEPYCX1P
OlePTpwdiysqojeAewyonK5jnweB88O5KhXsBbr+dotp8UmQxjD3Sx6ZnT30IZtr
EyyNcOPbUTpqnT0YBq1mkMhGcGzHg1I4H3YB9qYb2XPwMPkKTGwcPe9l18VLxPn/
Me1hHWfuWiW7EPrq6pAabaunxIEPxmXvVuKX9LwdxABIJQkO4svThSQOpWCGstOO
By3VnKQQc5gJ38HhUwHab1Yu/NA2e1S5EZrgB/ZsQ2V8xLfQrUBrC/sPkgc9uYLV
`protect END_PROTECTED
