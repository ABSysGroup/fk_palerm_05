`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
50mHKuAIbntC2lUD697delKmrhZeRWzvOxy9WCVNrZNt/pcMC6oWG4lPlCJT80y1
CG0DPumxT2Q4S0mZKtqMAEozycrwGHdsk6HFROw4b5970S/AwUXMbI+jbmZp+vw0
zqFPFKE/Li/VRTkSSdD1ElY1TC7GgDeGMf5lmZS9lq2KTftOancuEckMLck3ifNY
djxU6ekyCW8Uu5UV1Qws0Uo9UnCmuc5hgllhYLLDlmX3xfr7EBO4PwYaRz6ysL4d
O/VdVlANDq3Tv539XgpP0C5a6xfu+VduvaVb4iajY88CQDE2GrfTacTJtDDByIO5
ulQZ6ryzHloOu5xG/ImBi5wbs4qz6r2o6hOEvKjHu463+0I9KTco2cOVgRKLEMhi
9oNdUkLKwq9oFLF2zXFT67lN0rSx4DBZWl70CnXdeZ6+AkBO/PFpaSVf/69ZQEFu
ofm/19VjRiJ9rBx49ohoqHt4qcCtGJB9Bv1Iq7CZsYiTG50DZPZhlV2e5Ey7F+xR
RRwszH6zEnbYmXMIlVY3sg==
`protect END_PROTECTED
