`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cZ5G1GFXONy3/yHYTsFPUkJKBBwnpkQItsXW/CqUjvbHAE2ztUltAfl9GfYHfpgK
HTTEFh53vf0i5fxyCwWXDOoFGICKvMS4FdpzjorUi2VMax0GaiKKJFntCHw49Grh
gU+BIVPdxgYW3BblbvowRPXLGGFATQ0HudZg9pOtfuQk3aU5h8VycvEpvjXRgvvX
51JVTXPOE/FAERXc5rpDJm9ope01aGhYV9GAHO5evog/MRaV9mnVRluBhtTLJQcz
Aw9eoGsQVtpmWAipXaMNnwRxDKqeDnx/nUvPG3drhbTykgGZEOSQ/nVMUzeIZzWb
nZvPssfXoscMqdfJFEfPbcviC98UpXZvLi0JEjKtREYumI32MHuxF5wUQFjGag3R
vmJXfWJUp50AxBlJmH0XdWM9yjxaQb5R1Q++4sNw6HIfsn7KTNl5DVurK7lTUg3L
H5fNnCXne39gfm4ZcrmZJi1O6/FCtT5wmOAJD5SjZdp9CPOuqO9ImUJiQRjaR/PN
Sx5JuaKVJpj4XWeimtxSIHFi0JJ87BRPN2XAHJFZz3NGeMnLvDE/XhQSnqu4SHQN
0HrDy0gJUT1oJ2wq4OdZ2PdXnLgbgjMT6CfZ9jDxS3R00PdAogVk8FuhAn2seNKi
r0Fi30qZOKf6QzrShICF5fgzjPhQdkqVqQfbE27+XifyMy5sakItQbo+C2QG/PAn
uYLWLk0j8afhSymGa6z8sepz81oCC7Sw7lZdKc82v63W/EJ9GL1qqYjhH91Px1ZQ
+DdV4Idt61pVNoI939PMKsJlq+9oEVi+O88Wk3LXOrAM9SRL0EWzD+cBYc1NunDw
f1MyXgSjLrlr7xmHQzvzO1j9uyIXMRidg01LOIKkR4yBvZmadZAiVN4V0IG9BQzY
oWqklyJG1X7donYsQWqACvnAET7axgaAHT5WgeKYUx4oZTIuisU+VdUPc2VLAgIW
q+aRhM3MnJQvtUjWCQ7B21vsgVdmYJ8zPq42LFf2+P8nGu2RdUST+9CbJ2F7iomu
+zSlFfC9/7t0Lzw7UV3rVPO0J3x4K6UqhCtwVl0/KdWk1ugnsTmmH1qL+rirWzrH
V0hWI5TcIOCSWFklO4QDlMMPK9YWOsVOqo33Q8bol0rNPsTEd28ruc1gCjgL60Vu
wlaceiw23bQc2hHHk/35geOWzkkZ4aVaIRx4Mov8JPUCZlAs93kXBipMJSqqo39G
0G8TJY3QvCB7HPZ49E583cQTnxVDo8D5Tjt3kJAnZAJRmGM1flw2PGcREZrliTF2
+XCGGMwqiWa0kC2/7/ww/dNarX7RA6/qST2IF9jnUCfhWV1ng0s/kvKbP13MWEn8
7e5OZF9E6gpT8iH3GSVL0iDbXE2IVGLlqsqxfco8l9APktwjkKEZ8zeChptrIvyr
japZUR/y18uVWGfSy8nUAiec1b1hz5KqXEF8gp72ENldYE3HXjGHPKpoTtueS497
isRjTECPx4r4t9eg2IroZhsuShuWTvP3KK/sm3Ek0HaAvHcKp9jsQot6xFuW2vlS
WO1NdrPl+SQNyCwseCKo19QKa8tIi8XRADyn08zr7fQYN1PZ89MAkeLUkszDqfO+
SCHZ8ju//d07LdtHvnXeRPhz8PnwBjNLwdTXoI/SGNNNDs16F/gsCaW2VKoRE5sw
aLNfMyQN55r6eEtYqda7cAhSoxqakWHs/ksNG5F6CAPKexnPd9l2FxCpXeiOwarT
4bOeHdqa7C+czyhS6k0ONNWYkviCwij6KL2NoG9hGW/ai0D1Yz5LjDhe8laQMS69
fbhU6ICgXVn3Wpr3d0OAmhFTiHy9P9wcNW3dfWMixdR1MXAR/o+Ts0DBz56CqgsW
BfsSIpthxvfRrr85PLDN8n3XJIrTkYvVzoIKHTA6HnjUa0StUMPEVWUbXsA9zzWI
gbhxaakfZkGc9CjMwZU2E3eAFQ0xCJeaM3rVSK4G5JE/gg0sL3aID7mIIOk4su18
wVUypv3E4/Jw3HWHSnefSk6H3zSaUtrNvrKCzksOExojZRFlEtEpwU5rqTvoJNIH
1TFmAa6s6xBAl8MJEl0lumEpBAXOH0bBjcKRwn/OlhsrquXBqLDmX1DNYwQETyBi
qNnkuclrbE0eCwv/8oXdDv95uhG70D/9P2y51CNNkTE1FJB2wC5OAOHkAXGDMIub
QDjFwW6ZoWY//Q1mVU6OoqqFN/pd22dWCPf2t0tI7GYJXMmKbPczCBHrGJloiJ8R
d9dzoPtk6rWpVth5sLD9Xe/515ihVFoUj9BT2lCPL0E1MkbBvwOmfoJ4ZpvwqhFc
SFR1oVJj/YgFaLAB/bXaCBCRSMTWViO5Li17Sxr/SMb3sjJDQeKyG6cCMAqwtbXD
KfWkKsiTjrGEXwSoAIGVkzcQaE4oudqPCQpXuMDXXSrkL515zTRQ1SeeAyDYlhec
mmhtBMsCu9QfN5FvrIbQeFr8MxInBSNyAoViauLQgOJpjDgwcC4N3/kVVDX5aKAs
DSEAN1qTqMWdDB0P5XMDUSpI8q8dzxZ778L/NLq91vjiw1a33MunHOivRimesKFM
BxvqrA7u2TvOJqd3u46F+aVct01OQv3gGtV9wn2at8LIYoSJQUdo98tBUHPTGi0t
6UqPWkJajBkG7pwcwjaq7Oh8s9YZJCQB71oX4eKOS7Y6MxQVLIvEgrV4bVHwJn4j
CgxmqzEjwYOpycqj3BFroZD72/pLRZVVTPIAf34//IahHP/cDeiCDovjAGBfLdla
yJo7h38iUlmIETitnDzc2QAMpynZtq21Nx+atzm/XSl0PqZNOmKDQkn0ljQ1/UcO
yiEiDzUP1/62Qedwq2Wz4gp3stZ8yU0LsK6InlsZwPGiLiBu7Cs5HyCkIB/SH4hu
4xvW3FEaYn4rLE2mxkvca37eSm3iUtvlHc4Q1IK3uDd8R+5P6ic/pcPMOsxtMplX
8EKnTiOKDw6gyon7sZE/pIPXkN9Z2fYr1tYh3UqtWZT6kOJKwl/tA4kIC3PsBD/P
fOFkRXFQiUes4GUHarBGBE2qEZ3Ra37x5BwZk68p4ZVgwifSyz43YGdwIl5G6/Yy
/iwUho0nkT8FmxAyr36hljKc37NEmrvVgVKp8Arw5Cvm+6lBv0B5FbNb2HdNWoeU
KvXgOi+gp/epdEPIyE6qMce9rySR3jUNKcnG6Mc3PWGC4/i6LK2TNxY5k7RxGtZY
ZO1tU5rr0wSv9cxgUPFs0kahGguKJiQf69THP6Pjymhi2Q6b+vqsklbQUXB9Xt71
U/loHRlbqik/d+7ODs3Q2zKGAj5btzWzuQRhTgNg1wFs1pYoTpRu8pZ6gBbKzuGH
jPxXwelV3uKeIh+cxNJnSJTIC829AYGru72BQBY7bJCqVE2YtDSklRbRcYiAXzWy
KuIp7zJrFP8A+pePblB/w8P0XdTA4sC6UkA55TcirmJ6akR7eVXTgg4WrNsARg/z
63dKzLB6/Z9M5aZFQTdmIp1VAfTm18oI7nEX4ux5g/dwf3lZP7Cf7HKl71NlHjiz
NDeR8cl5ZlFHI16sWd7/EeFGndAjh1BSYnCtdDsJIjEh4L+xWQ9+Bxbu3jDGE4A8
aWubn7HFUCJhENPBB6hN2ZIvjz8LsW6dqthcYOelRTH1N5PUw0a0O5sOOScpm3Yg
`protect END_PROTECTED
