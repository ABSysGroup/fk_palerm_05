`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4FBTNC4E/BRYwvgVBVxERAC5EJKGqiAcy4J+I2/GZeFGalmxInbvfuOYnbG5QZTP
PMwY1bTp09i0noiuZqCLBKy3UfGaaHsou0JtMyz8vG8fSCjFQU+eF4DF0NEVltxW
hcjqgC38BXFQ+e0z8S2Os8Quf5tEQ3LbEF+rSQPlnrcZm/iL0YZBnt8KwO3HVdnk
mVbjhW5y2lE16cnqAlMQM5SPhVq37LuwPsZF8KhU8ghSPtss2vWq54xWFcrZ9MQe
I8tOYfx8Mwiw/ZKvgz98LcySaWqO+7WMqtAyhnO2ZPcghIV/BnpBF86Qsj31tQgW
dF/t4k4rUSTvz72AmeHNTO432vE6jhL+5wnh3N9x596CmNLi6nO8wMZsHZvm+V3w
YF/ueZCY+vnja2C10+hyaFkAHZPnOXu0rhlEpie/dlfLmCMIgUSXIDqnDj73pF0X
sAgcl8EUUBJtplb7trYKuZIYOynCqbRivM0lHBo6JiqXmSd5UfNQrLTzTotXtRJL
j3djlcZ9w0HZxzulRN/7OY5U1l52Q6mcixSwmMA38ShoT72yFt2C/iBytQosLoEC
kK8KmB09ay0CFI973DcTXu4c0Fb1hkKoVLMGLQBzjdKfDISksGljBjBXR+jCMLFZ
BzxY25HXQ2UEWu7OO23mrdc6RocBGOrGPzRyPq3/tHQkK4yBDkrIngs09ZFKEnjy
fQ8YJnIgdFsO4vvR5F9fCCSFKr5UFQx/fYc4RcqCnPLocHlThW+wEvlbnD42LG5V
7rIlH5m7O5pCBi1oF+Z0BdOIzpFzTmnwceIkiWB8H7mjVqkJyp/RBsaD77+IY2no
oZYWg3SUK1VHIDsBxTD+TnllkG2clDPrUvkIjwT+rtXrQj9EMcHctW+kg1gKqtfm
dxtXiXEk27SsKJkdqKalyXIJgum7Qcald7AckZG8PyJtQvhJXb4pirB8ZWv02ibv
`protect END_PROTECTED
