`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rOnpyUHD3MqBv2Rl1uxu4UciDTVU+LwWStRq+BA3upjjlnQRpKe5aCkaxd2qFVDD
YSNV3jvuv8AQ6Gbby2Ih93SEKv6lAB06r0WUwUIvs2XijOn9SX+OsAEj159e1vNF
VNsDYvc3tPT2ZoPQs1Ctto3OWDarl2TxUFuZC8W3TUUGXtw0rs417AjAwAZ0GEbz
FwXV8Z4m21SEZUeA9Qd1MkdpxPK2mzTXOzSCH77v8+ASpxsVi13Tx9ViDQtQFoMC
WmIg42ryJOgCCkTOI0Q9Eg==
`protect END_PROTECTED
