`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/7gXRSz3LPwdzm3bkcM6pkJujp6OP7UwCDAtApN+3YfOYArfv+/PlppYTPYf0/b5
9O5t0/hsEy1mECifVGR7yhDF7xpzFBRZhMXmy7mF660woDUgYyajq+rFE0/9rxus
FScOJviHJc8T+62JVKTqyCmIgFUENCt1Byzip7MfFQi9QhY7/1bREdU0HZ89p76I
3VFLcIdrv/pKsUb24n5J88cS7AMFdza4h7A4EjjTtmAQZAHWapCqheLKLsCN0kvL
76JFQ+3nJdQZbeNyuXXzLDEUi097CHzUnc0Vfa9igfiWkuexjBd7LGr9WN6UwKQC
wVNxW+1yPnwS5xuJt5a56kJ/WiQgdr/ITswLIVZKvHgKUON8LWMPp3eVrRLSaste
PHtXZYx0WrlBkuhbvaEKXRi6rBUH2Ffj4zwbNg7Be8SnA10nczMvtIV54eGBrBeA
`protect END_PROTECTED
