`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nJDJ8kXaiCKiiM/TXqiyDNtvrfJ8z92mhIsTna83TT5PVJEK/SC+u1NJADWQ1iGl
z2mr4GzJiazTbDYX7FOgXtU7FCXo8W2hVqT1WkVOUy1nH5JLFW4uwx4HM0YrYcp0
0Zd0csrDz/FcngUbqlmwFqHmPsTTYrcfY9k8uqbZrz1vbeOUlXQOzKK53Q31ImgQ
Q0t4R8oXmlUPkQFJ5oIZWrEE/veb1zm54HqxkDa8rAleWl+dDjcFTAmxRTWMYYkc
orecgXTrslE73UrHp7DaxgR2CvzGpqMHHk7GhlSSD+w42Uki4vensRA9T0UWr4/2
jH55UBV2h/GPAl8gregJ8oOhOAP6mi5aay8sQFdD6LrX46FbAFvfO/HpEfyV3nkx
NYPRKT20ufIAHCUomSNXhdfU7qYmV03LUrOmBwFx7utqxmB8sqEBQJ/yLvFVVFew
Z5iaU8wtFhkWWrD4cF915QdZNvLsWOQu6/D8nDl2KdCNdtf5yZwN8Nn40lyium4M
`protect END_PROTECTED
