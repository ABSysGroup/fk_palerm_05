`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kADYXZ2QYq1UAHRLZ2PwhjQBbodzWfV+RxDO0qWI3PyKg6eQJ7kokKDZc5CshSAe
6FMeRfjF4WPxzGXTcP/OnJHLJMJabUIbmZaEmBCbBPtVTK0Ne2IAzdYvUaZvg0JE
whspYUjGoiJRHjGN/CrUlApQQS33a8unbKW9Q46QNgcu3QuIr6SEaZqp040tE2yM
aJtj45Em53UvHJX0rDmQ8zZqyahzUWWxIEWBICtu2fj1ul1J5XWnqXpsF9V5fZC6
zCWzbMT3m+0evOkSCX2OAwjrlcrvCN8DJc4ElOuybKNn11u0V+K4hoResUlvFBtk
JLfYCTN4QwC5m6blskd6JVaOu6N/HcV2fBTeT3IZ5Y9FAXxG2jWjwIaHKCY/x4Q6
5dhQLCL/aAWZVtZok0rK8zSyHPmTuRcpz+ScnEiISA7U+XIsBiywnLZgoKpn0YLk
tP5dBwK8HqF8Di1dbf8M859gErUj8RuSSZ1ep0JYZ4eJZdp7zqwuDywhi4ZIz9UA
yeOG5Xd4jmPkHnwMPvOI7b9WrNnOA0j2tSfSi7oVrW4Zuxbc//Pw0RQrOqxAq4vs
W+KYKuqQQcXdUV3Yg0mqFqc6zjsxNldv5nXu/iGzs9w=
`protect END_PROTECTED
