`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mql9Pg7GDVRsc5pGSDUZ2tre5Hyrh3q/FoqTcDhhqoDuoRhn5LY6WAhtHpnng9Wi
75tIeY65lKHVnUeIFuyr6NOFGbiDKGNUf9XRANbPK9+cenm2Z76f72+2TF2JCCda
GM3IFEL88E+RNMeaVxtROqTyY/ycq8diMebLBWMtgvzz0ElCgOIpbiyq661TqLT9
Rd4sQaN+IBUEy2ECRwkw44iRVl0FTKorslmA+xBUx00eqJ/z4hqAJgVJeeDaAxvK
3bFvaOiDFKpC77TN+a0MjspgYQZnO0xxXl7hC+Igqjj5Brr62iVdyEhnU0ochlA1
Da352aX13CqH7ys5NVOiKDrwTU9dGA9WXizFjSCR+ktwcX4xzPT1jhwsHRuHb+R9
rTnyoodpiCWI+D+VlDt8Pw==
`protect END_PROTECTED
