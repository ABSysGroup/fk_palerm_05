`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VpVxfebmK/RtW02wajm+oxOAaE5H8CFx8kIIWHw9Fy/3PmdP9qsAKFUE6PDi1VHA
EQ1rgHtczMR60EJvRiLBNnmlWzzxAPl4q4n9KBLMc7OTa3sDP1S92gyAH90RlwVC
z4IEVHI6/9hzy97Yuo5SJeLRo+hrjree/iMHzO/5PqksemthUaOuDEAFQwF8vqMm
oEFwmICWSnZV0Rqjiw+yEU3bBISQNpgkyr5bMY0gWyz4VdLTnJkyTopR5AvB55+5
2VkRmBN/sizunDaszmnukeFkDkaSoqrNv3zP5v+F5g0rfKg40oqnpQu9KtDwAtRK
4EO/6fjcKwhnRmwgHwVbpWLR8/lVRC7PUIq8nce9tKDZ1o5pFuDxEiwogwtk91Gl
W9SR1Uzioy/E66j2CMPSLdYDG5aKz4/ULxrSyeyhwFcaY355WWF54xQRzISkhMPw
jY5IMNYirQiFsCKkyzhaW/BLBOwgRViWxOP+fl20TAXo8qa6JW7mvRDnQIlxRSuT
JAWPOs8xQIJxuIWm57E5qd8dGG1LU91ubQSSVCPajYFxfwpeIIuviCi7LmUu1EBB
ms7ZwNysSPUyhZ+l9HPkMoTRfKgZ2JBLG2jkeiMXu3H3i5oj4Mix5UAPSejfHPTb
bfPAXSR6xdQimTx1VOYPZfMXz+Q2BRk9Enx3VJFZZmyACf1rukMwI25fRZiRRXJ4
UTfO7aw7ZE/vJUnmWgUybNnpK34yio71habcwgd/gRM53OhX31MfSalNfaIZceE+
e37JThy2q3+fBGroK80G8Q==
`protect END_PROTECTED
