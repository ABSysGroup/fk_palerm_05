`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FhGV7Ff8+1h33wGcFbVxpcNhmapsCYlThufr4DVehmkdR+VHyUj3Mt6saNoBVsPE
EZ1FOdppQUE/bDiiR66Yfn7h4EhbVrGhzuHFecmUyhblmif3z+HtGXW20cGIAJrt
IEftcHASjS0XB+ohRiMrsOmN4LznzVnxPIId/DYc2JGxJKmjbQGEWKlORytqJ7V2
E6fmUGBALTFRadbmnM4lz9BCDxt/lCnay1yxnRTvf1cRDYFxXwF5kHLR6fDvmpWo
zucKTyn8mpaH0Dw3oBvbNO66fvdT+sPiqSdOYtNNP5Q=
`protect END_PROTECTED
