`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PPnnJ73eBYC8Wl/gtT4rcwy1D8iz0pIZ6ocHQWFFAjjjFTpwIp0TAhyZehmrr5rO
hnavIR4z+IPv7jFyiaiwBDO9bNSTm2WWumGYIZnmjqt0OhWcY7EK87mrzbfgcK9N
E0B5H6Q/H8vP4btuWsF95RwlY7SlKuMKthfSe+bos3MNS1C+8N0a0TGEbc9tw+OZ
15z18LRTTBuzSsveI2WhWUXRe2WJ7M0q9aAm4V6guDGuRWoeY2liIk4ljbmET1SQ
aKYqLa4loUinyb5Y8Uvf6txwHjVZ5ed/0C8TkbRSYhuFo1kVlOmyZr5V1h6ImIbU
Z5WgKEYB3HIV4TLdfHcY/js78XczOffxqygNy11V7KCN6rkrzXIdMSIdAmMb4Enw
FZpQ7A+5P4e30bjl+c8Gke1r65XRcPkrqibdAx8Ly3etUmKtNcsZ+mgGl1nMnDC1
j6CVOtBS0lal5DWAt4G0roNnwxFttza5OUZRgWwPTPnsrjQoAmWSrPzupmeJ/HIt
iDI03Vzn9bA7ldeg4RvfYnuX8NNl77jSE5jj+O0886O03u4ZrBuUi26FB0crtMHm
xytSaCLgsBXZHagnFw5wpfw1cwnwxk1F+Mjrqq6J6epQNw9xcDkyyhXl6Ac6hYJh
1l+xqY2bKKJHw2HkrmkFYvdMh1pFJp+MtA8dA+PWy4+dPINxm0IKfqaMLbWjUmPX
dwoEixKKenNsgBrTylMvSpvfhG1PL/ODYiDjc/2Ooxcu7q6LcEMqkSx8Y1cRo6qO
iPDxIVe91XWHlwNAIS5nQJqRHtz7xk1JKyY3gW+sHSvrDMZTKzBHpt69orQ2lZVl
OaNyDdNJMpK4nbCac8fbDvVBrljuD+s8qXT3KtWMlE8MIUrqzj/3QuYAERxPkuJI
Z3X6wN0aAgr57niVCPc6LWskBomRyTnAFFvgBOdjkhQXzQMqs5iVOWh7UUW9HcoK
g8JsAepcoo0K+umCPQUezr3Rk+RqabZkIHSvixFhxh7STfwvQwv8Kibx5FM5zqgm
ZVDtPN9ugoQeRx+QA+hLp1OmT19C1dXgjIRlFBxqXSLdyqV/Ys1bAlQYxqDoCuP6
s8zR5aFXtszyjTRCcoFOVqz+Rx+J6FlNnmiRlfyC88AEQUM1qnYxcZxbEWT73r8w
`protect END_PROTECTED
