`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FIsvCigP/Fx7fqU4isnrYd4jRFSDazerDewZb8Pid9rTza9ZxFl2OyRpRX3FNJmq
iQO8fz2HSkZzO7Xg2tQfaZ2oAJFxKvBBlbgVvsKjV/CoCyitkPpEyIyxsUajRt8B
8SEdS2Smv5Aqv1q2em2upVHv7FbMi/8pUkmwsOTc6VVFTvPFWHZkzjG7gcppNTID
Ft908EvkYF734XxdE8y9CYtiR2bQjtsR+FBdM8oG9yr5kOOrOuwZEjOj6duBWrF7
mFmVMR789ky754qLCsV+4sOqYrXdnKkfJhyE14ymOwAViLA4cVM6xw5nWEjStSho
R8qEL/us2hmxZj0K2jrDXRBh2wyNNp2NkI+b/cNQQRT47GxqAuEGkhgk3y/fb4BG
lkFlluJ7EYQVxnt5Gl6HwsiMYJeDamnJsYZajiSKdFOjzrLN5gk0GhGkH63A6YlH
pkgW/C2D+hAhZfeEGviSkvIHbrYntXxxwlOzNCYE0MynT5tJwl8P8htqM3f13y/m
NOjxzFOzTpLnKi6aNDJhc0oEHDRuGjDL8w9//Lb1tCfHwH5mqEi0S+w4tHLFw+sA
K5SEXO1f78VehZB9rUjsUlybR7TpgtoWwbzYedK0wx2+TWbNg5yaIdTXFAjAW9f0
2Dl1jHqsGma73vVRCEgBkghJFRkzZePuvDYJmDX6to48UMWS356YKKJCj4fjEYdm
bhPRBGhEoG0dmk5Vj2KOjjRP333ZJiHswDrZy3PTBw8R/JRjK/4ygvIeqGzewWnh
IkNK1qdUXQMFfSP6vx6rHMSxd7LCbpu+LMdJ09i5TBo=
`protect END_PROTECTED
