`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q0ZiMN3sr+T6a38QO+dt78qFUiLeP7MbiHpFNOAwGfIuLluu1FI/hUL9bRumuKzV
yp3WIGrx6HijmHUd6dGa757y9/e7+kSRaMMEhiTio5wYDzX6ZEYIt7i+9H4Vei17
5R3ltxm43dDzv7GvT+GqTqTuRv+TVpF8Tp2huQJmGt2/NMG+57HM2yN5eJpc/R8H
CqehaFJI2HVDSBwDQz3o9DsKejEYbQpJ7ihQpyJcIccemUp9rVyuLk8O4DBKOo8D
/rI09uHE9oWvJ8YRKUGxBuHe3imqZsmuqNoIE9kMgKdCcS1OxGlWdsw3A3JNlrvU
EHRh++dvi+xvSFUzVQo0yVNPgZ7fEGTuZa7wWANo+sqUHMEy34gYTI2ybI01NV/I
9Ssk1migylxvd0vd6+wzsg==
`protect END_PROTECTED
