`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SR1mZ+Uo0jXaxYERak+EoT/MvntFXt81G8u8JRwDPQjiW4rr2TogDu5QfGetdU+5
5S53FVtePcpbQJO64VuQPPRZgZIWsdmE5CD1R6/34yCTBXmN0G+A30/3FIsSIFq2
FP8ehRVIZJjOjMWIErzF2fSzAFOcLdcocA8djJsmZt4LcfyiXLsO38vX736Ss91C
0RZ3bjM8NE0uTy87lDIaFLAvS3C8CwATutO/wAfdhRknAiQ4h30zk/9o3UTYRAfT
i+R/QwsYx3HW4xBqZ9v1/313Pj0VUaGo+SiYdg6AWuKCUNLEtkKtSMlG0f4E2lPo
OTv5It9tLdVzldKCLkXNn12QRCXbduQLGHT2tRmdmh1E+ZpKLGi+DdaAfEEfC1kr
oUxJhqy2ImJdPUt8/43xgYMqE0OYP/ctoxchuN471/3iW0aGIdjFSRszN+8GvsB8
AIvgO9xXxCm+JpcWHkSaRSSdkZOk0mb/Pk27cZUwXIPmya5ejne8kKUE9eibGJJh
MV+eIPrWPJR8gvRjdkghMY5k97Zaqz79+xkKpEQEyH8zT1ItBTrfRa7CABoV/MmM
StU9QMOuiyKelP8DB4hCIzdh6bPuzPBRE0SHpy2Ebf469vc409lZteVhskF6nmQC
ajrJ8WCHs1eFsLh2KxI7dd8cZmRoef1fjeGaGTzKDwyLvS2UhV/Z5Et9//PqVq3q
FYQnsuObRSTWBwcA0JMfGL7c0XNimiVAfBNzR17W5TlemiNRiKoO9OeVBGpozqYh
4GkAcBOgI6zg7BBG8BkcMw==
`protect END_PROTECTED
