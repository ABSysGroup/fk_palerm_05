`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zwvefDUqHIzA22ZYbx6xoMHOCdKmjqRHDAll0iRXr8b1IlxrTJp+ooQ9kMlnhw1h
4HC2yfBAfHoqKgb97MatAAq5K3GpWcux/OipSUJFIcM5X6wOhj5qzeiZKagstxbx
0k3maWxRDyHemSgJsLuJh8mYV8PgL7WpvTPK6OD5X7AvH2BvmYHbmT6RTjQOSYBr
fqgZaU2c6nMY2w8hS2VC42xGbqW+97f7IujUUbuwCg8IUOW1bCTHTDIYRVlqiMv8
rJgoatDT2pIlG9xkTdV70YNNXT9xtqEMtWgVtHuMF1mG75y7xJxCPofioeW2/JTg
kLq+Gt2lZe7kywR96uEZZMWlVb/VLvmEmgX0sTP2HE7B0d7DUiG5RfoDK6y7DT23
wz18jxu36pzs76E0xhD4SFSKrJvNSBzkyVdsINLgOp2+ncWod09LtsNZvk+2xhjT
unh+/PIrWn1hqf5zfv0DnJevvtp67NXLeXul0RCf8V4KmSfLv2dnUFuxU2iyynr/
a22APCEEUo7fGGOKQxd5H+7+umGugljt9KdMCfnG6yxXjUPipKaNQISL+ygPxOWr
20WDcv2/JFJBSslbPNtM9UZqA2VkLiDQXO+CqbKMKUfW9Ot5OD1mVrE2ZgaNtegm
BMXOhoxPiem6t5JkeiKcv+lcJOpsHeMneg7MybO21N+liUq8KS3K52nrAvH+c+xv
/RvDZQkQ2bwyD0sCFWtIPBg38EtyFHC+4mVH2XBw5PWFQI2brv8A2OWOCA8dVZ9B
1LUes7V7PieEt3YDyePM0sToe76SDmbq5/oHx6dIapN2RAidz1ZyRTRJLW/1szV3
i+4PyD54uRRvgewXt+dIWVnRRHdDtL+o8ABwatKhpDIa3P0NiJAZezqipV5xg+xl
3M2ahzKvToVHy26zOpf550B+eMYoncasgzNghogxV/Nbf2yS6ZmbXLsHSIloOJyD
cYh1ROVdw6FTlMCdnXOmyVIXIjqJpMw96jlDJmsh+C0GgEXS0uc9acW3PuFevhD2
MxWRv18mwuc0dElAwuER7wTnRlZX3a4OuAFBYM58c7Cndx4d38PDWBJkIT7Bm5Zl
Cvh64Jw2esraLx0JZVm6wlUBuOn0KtzdAIFkg2M5M+O8T6DFFBT2arhzbUn/VWAf
pULoGVil/d5DJOjqPxY2bt8eWLt1Dj/b/2O3zc8X+9cr7GsQynS7KHx03tt5DUro
LGRg/YqpBOxM+53jsflXoCUKiOpNvZs2uH6w+EzqDl8StDnFp7BM9BAaaMozAFtq
4ElSia2C4tdWNqXVAI5fQXPfMIwfLW0Xx/d1xnsXaly3muyvFfgIpl1zh91sKXqa
9xvjXf4aV0gAfZEz36smnvRVWTD1y3F+uiaaiDkoyYd3Eo5JB48vz59uhBoUKDkb
CHGyTRFts571p6vjAUc/EiKcKOIMXJJuC6yxspycCo+rAtNmMjlqhr1WbsbCD87E
B1dsJ/28kUDo90pFSN24Au1AWJtkpPf858nCteUKNykWiCbQvSh2ZVkZheksrLM3
yFBG7MBd+z4ZUHQvg3qNsMWZt1n+68c23wKO+eytZG7ZtZQ92FTpQN4bYi+K3Z+H
NNcYVllqx6kuLFvekEgWRtRDOvK+eRQBLPtKHRUkxEpW1SPR4QAPxzFEn5OMSlSA
0qDUHhvSJh5Rqa6Vc1ymFPoScyOu4OoncQUh+g78V5HAS2GhqYcchwcx29ZkjwIh
`protect END_PROTECTED
