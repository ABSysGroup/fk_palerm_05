`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tBxLDQMVljHXVl+Hywd6utMG394ak1j4nRkZMIfezJdTO7ufMu2kgpTQTRMRQKBJ
RivLxHfw1Qr+rWl519iM5rqeEoItXTjdhNGIV7H2+bb/sOaqaqtzauEhGLv9cL7i
hNyr/+IqH7ys1bZssKpNmvzn2tqPPez+QGsk3OJVhfhWQmOCh1YsvSwLO8Hj32mZ
yoPwXH1kWZc2mcDbvsy+/rtypMi4h4mK9yKHdOfbqljMjm/5UdnYFEvwXwEH/Js1
5iJT3n20u7qO4Qq1QcC8qhbiK4bU1G6PVRJEy98z77h9Hs8ieZqrV9zhHRAdBCH0
euy/gbuOzpbeYfEymUOzi0GHPwqjjAeFIByW0WkmMJvEh52CBofbI8HfstzNs9f2
V6Nj9BBEadYc4aj5xL6+ylERnmx5t8+dhFYtWLI7SzVXsUl4k2CP+J4yFnPsaiBw
PNxcPHBNQma/JQbkxImEIvbTNOeTg14Hob1RKCTCkDrd6stvRAZ2uSIFdjuZRNBe
WGT5PernzWV4/yw4BXrtB63X//XQmWSnfb9p6+F82Z1Oo94eTT+0dmX0TfD7MHsv
JwuJ4NKeLv2kd38kMLRbCvk0v1gMScUPEPM3gpjTNd6sNo7F4tgrt8JyqjYBEr9S
x/urvd28neNlYHJ3ZaajcDR2SXRD2OA06dyJUbS06agwZS1E+Yz9XF2N1+TPWxtw
O6GLthVF7vu7G8VzVcU1xz8AzY3TW2YSZ5wxHw6NWIFuX2XdSaTVBIIebQPS/VkC
6d/uNzFGSIXKL4Adz8o5lA==
`protect END_PROTECTED
