`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LRX+FXoQPFX1uVJcojZCHFz6XyGwgb+E7RCaluHEla7PEPzjUyU9Gzupoc1770Hf
yCXCgYq6uOK3aCNA+7ouOjLFVfg81Z/bPft3cqBokiTusFpMCHKBLbRz7JDuon3K
CP7VkyV9wx8CpOfnZxBKFMmAjlAj78WOiGrn5z82Rob7Ir68xxkC+e/rbMbY3sla
KEW6V1ZIhtU3z1Ma+hVEi5HgnmJVDmG3T1wE5HgyjsZCmxu/MUh2ve22bUOFNwRi
yX5K4LmtdpAd/w8xAubFuQ==
`protect END_PROTECTED
