`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LrhLdpsr+mfjRjLMhnSN6ClyuP+Wb60Iuc1w72BYeNw7x4vynuyv1HopPQavnNgp
G7ucyw5SsGAq9v+NSFyL+I26eaHsky6HJ5osuQtEhzz/FzMV1YGCNRdR9YlTg2VK
8RrQEvkyWpY60TBDDcvJ1LnNa+F9KM4XOyRJKuvwIkjl9O49YGL99AzihZa5q/m0
EKjexdktV7U20GfzqAmoNR35JuU5svn4YVreRfVIsBkxvzCpgHzX11qOSK8SInHT
87cEh53J0eCWbnNdF5Tlr+rnQqy0LrwMyHouuux+u2NmnkkRCZDlO6xTSpDGH8ZF
4NLRUXNnmORR3jvjUwX4kOn6JEhGHCl6tcc2/RBDf/LYRMkopXeqeEpaFSFmJ3KV
Yc47nKaXtJDVtumyOSEoe68IHFSya0gp6/UlF+DtJYQmTW7GLvH13nBGHy4koAea
HoBjBqv3AU0m10C5/gvC7gvNLwcQM7R720MsGklOqVhxyKjjzXJSWdinFqyHOsIG
mJEJu7MPdfucirW4KYQwD3Tx/WuR2N2H6JF4X+ketp2qCJbxsDVAJuODNXZshjQz
bzAdxoXQOK8KtVQsF/thuLVuO91igVA0xqKgNWLg1RpyOWp0ORe72WSRbPFoI36e
NgaADW6xG10Oxf+dm17DPh+HyvJRLxU9BT9XjfeV84n9E+/tcE0l6FpRHJi8/VRN
HXGlpXy4pUtMvLigpEjb9xLNGRpz8zkm66uW2ZnQaQbZIHJ1fhGEuhAsuoXr8dMT
qjGVBX2GT/za+rUA3wOMIESvA+I3HIqKU3Q9C00dCP63N457aELzVLnbtOF0WR81
OnP2di3pV1vNgUBDiGhZeEQLcNqQoPEGz07ZY2vqEKIyQIoqD3ZL1lL8iV/Zpc++
EVZozYqjJ+3gRr0B77EZuZnPnebAzgeq7AT2492BJXIgj4klCnmwwV97277QqO20
bAZAlxcy0M/xseNwrO/FzSw/41F62TAUoymxFT94crWoCJ8lVMqLTaXnfj3gVOF0
/Uw8Fptglgjg00bs0NMFpNlPlsYvPP9Ji9NA1aQe2VTqYPRsZAUOxUs7vMWs4hRC
0IhrEXVrUPG9Z/9BItGa8QKvGo1dn7464zJbCkRHqhNGcia6trRxqhmXY3iWdWai
K6G7ZT0Z1PS51lMlEYDQOayr0XerwlQ1N0iL0NkJa+ALy7hrTdIZg6zOHY/sBRE2
sxfz/1X0dfZ4No+t8N9B5BUFoyPlHaqMmWzrBDMn9VrXvduRdQsghQu499KXvjlx
qx5SFc4rbWNgvUS10xmU0h79l0BEyVNg/fRdovpq0yHrmvSa59SxOYMV00V+w8p3
JsC2rOfXm0YAiVWnbY+8IvEbSMaMB7iRyXgRzESVayooUdnFpazjXCAToINKusLS
HdO2WzcqZFDetLIVXZHrxJ3HPRbQna60yxP1n+Ykg2mg1K7rbFE2MSnL2Fo1+TYj
a6JSMg4ekoVCtiY6APqcc3Xxx7aFZ7bla7Wt3nh73YDk9Hv7fDASQaklpI0T0vAh
x+sZ5RwQkXyoJD941yVZ4VxKGPLfduD6KAho3VVECpbUo176VvEDonvR4aXUQh6f
YFNMeFuuMFTZNmRHbw4UsQ==
`protect END_PROTECTED
