`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8C8XC8uUiZr7ZpsdBJZn+tVJMJA5SQtvvqOKXt1eFM4wU57R+ootqTKtmwYojFhv
wFCvQ2dGocavCXwjOWDGR0B8c5ee2gWTwct/ZKQuEEpID+CaSGFTiHPpShAk+xE9
NznWpdp7f4W5fuQqeKNv7CtA79epoIhY8+xPtNJAFKLoznz1SVESsVqvo36I3vaZ
h6NjV1fVNOADKhRN8NJtgZBV3iSgbAv+GuJ0u9XHFx++/JcqK4x/OX5VqhosjiT9
Q1LyxFj/qjC7nw7KAW50nxZN9pdAI8tig3jGMOD9KKB197AFhhzoJGl8UEF6ESXT
5IvqKhY3S0X0LBPR6vRhOz/RreRzNpe/xwaSuaHR7H93jdbruWcmwnvMOCi+XGDd
/pXXF4wlh8k1jcAJa6G+GleRg7K6urAdl722cZks8Y42E3rQ6A1jIk5ZWCUavt/L
z4+nA2KLKdS2BTv95slR9eQeu1kupLht1UsZb5lG0bMmBa7i3HklscVKDb1bpaB7
LefDzSmEhtYM9MuRzsWkWwIwC+6X826HiH0J9JdXEpV/o8/PxZ+G3HJxkjtIHDU2
OrcGjbX7740rj+Wo22AQtadG+pGdbZSg1q8Z6baPc8sFp2rW585a7r6GBOEhiB3J
HNKn+6CBweS+y/inBqUMRiQ0vwYbXgG56NuUF43qIi6njFHwSvNip/fjyRrLZfo1
kdE8CFUvT80TJqJTv4fMpm5PzgS8zb1BS124Qy/8qcjV6fMfvDQDulWNUE/772Jx
RNGaxwp2oHcEYg7ozTnSplpxqtSdFGbONwwSn14aa8V/AvQu4gftmQa9ud08Zw2f
vwlXw7alK4l4Zr5G/F1a5fWckH3JppCJUXCcyqvrEEBJl9vnfOWCcBKUXpW5Af02
nv9ibyEtsjY6T0lCEzvzHwnkDvMAdzSea0BpNKLwD0rGA4PPDJvajp07vY2Aew+V
FR8fa4CtAolJH+buGWQ5QaJZw8J9PjvcKMWeEM9Q1B7EfVTTdnLgrfZecdh9bl6S
JBewKPZAqEa+x3lYX4YHqmr4kVS3zcq32kqmlJGsgjb6nIgfs4OYjahMTbRP4EON
5t3+hsJTXE7OfdBqcThleYlscbEhp3bL9nzqnJWZfVhi1rVkAHU/6slwO7lFU2Db
b3TGKj/c30xAzv7rcqBt8/lGk2qYl6G1PaE70fdlGWb+Ll4FnD9xqQjyB1gRsLRZ
F+xZzRPVedlECcAJ/fKFMGMV0Lg5dDPtYLn6M/JUnykEA+mgP0mW9ILXCuRGfw4a
e0p13fadOEZy7gFfIv6daq3HTl2Jh4wwf4aOi9TBOsjIDfMrVWvkt9FLK+n/ZaQf
vpjA3bBMVBiCfismYbeE1fSIJG1KEdpF+4o7CmEuOqPhNGRMEk7WxwUMG2a1j2rT
bggi0K/8kb/1NyXEbiqhi455ck/i1DdQnOXGl+FXXDEUrXAVRPUDEiBg4Qve5Gpu
DVweyUL5UXCRWM1K5HK0gJR3zko09tnty9ZFTLDhfl2D10imDXTpR9ZBNZzsdp8A
wOKtxuzevuVDsUaIEhd5b7kKhdwR5T36WWmjZIWEZ7j06vEIwZug8017psHYWgy/
vaBieMH4RTgOConDsieLFyrTC0GvOXMVd5m+YpdalH9dPHacAsd6P2zCkWSHtnyA
kk2o30Os0zolcbIEWEErt3kY7DkNIdTv729PXp3D0NsVcAtP5756i1xnXALtvEt4
R76JI2EqxaP4C/5PAu0CWGzfUGB3oqC1SHPyxeb7QqHNgkrrMjsPFB7h0dS63ktS
zjTTVg+Yg9LQk2RJC9z+iunCZ8zEHxZhl0NeM1mVHuIs7n5wzcULZ5Dl0uXAeCs0
M2+df91+fkPxrsWu1CwJX45Fria4nVkhQKtwkD+8bOTW9zNtQ6VCIwkzhbPYriGZ
YVXThFKRSOe3kFFu7qCGDCuDhoaXKGuA3mvxHLM+uJwBZPNVbJ6s5DvYzyDanGgh
Kyc49kTPiCeu/3NMsJ/l92r2/9plFl+aviF5F1FZ7YLY71r0Q754KwyzH7zhI/Ip
s2TbGQEHz2JAlShqUEoHIHtoOJUzgzVf81J0t89cnmTddlpzxgcV86pkOYVol5GG
v6VnayhED7z12b5gNJKtHRDcRK2Z30huHRUMkGi+lxO7jytg4011f6DfB17Sjysy
4XCCIqAeuKKwI3jn3a00DuNZ99Mc+uKORJJUKs9P+R8BTKPpJQenGWzGX+vaH09G
bqkDvM87Ubn29ccnueP1eIkyo17+YdSxjF1lxyr6TkcDpO0YxMBJUYscnKaQWsYZ
Jv6BLnq9D49xUt9fMymXLs0JzDwTk/RiYSJhSiXmOeML3XrT/BatUAHqT1OCvEm3
ZtDqWlxnmVnbm45gwTjaQgRpCUzth4YQ7CtFJ6FMCCzAa0yicaRE+S0lJXj23/HM
LFH7xyPgJHU351H7nWLRpzCAjJDWj3ronxm4hWhTWxcoicLpaKuGr6X0Y/0Jxt/3
JuROhN+mjBcr1WPFiK237x24YGNn7+5HTBACjy3fQDKoJLuA3k87mwi7zV1zO7Uq
NSskoMpzKFFbDYWlq0nljOho2GT1Ovl5P8Q7ZSUu4JemRHoSgO5pBrKAo63LbrMv
Xn47zTulv/G0Pdf2uuN/5zyBc7bhpdMFVDS9xjGmwSH2Ji4grlfjtDhB1EMxdgVW
970F0So4N4G8KT7hDxdzOlCbg2YhYBGgmOsAQmJmgzW8MtSbxFsEg1M8WvA86wWg
MaDrWA80QblL5gAwuCYb8++Gbrq1n97ZjeG1fxdiiOfpV1Jic3zWEJOqYrfekdgE
p8YsXsPdDrjaOVsA9X0MFEiuV/IQw+L886HKAPMQviUkDjTYwTc0K46qUSL/Sp6s
D0O5rfcL47ONvlNPm+ZlzdFekMF98b/Mq0qVECVfaFMFxrKVFj34ggbnbmZEcp9W
Uj8cLyyZtxN0JfFn2UACtsXwsUa/RB5Ccv0u4GxrgPRDYUykHuKCesdELlrZgeHz
uki0squITAA9Z9Ysmo5mfz1753w3XyF70Wka2Kw7njiqetuCynn/DtEomQN7QFiG
X3UHrpKF0gZgDZLHCVuXPDu8fK+fpLaNcCFGJey9c3P/PJuwB7rNG3b9Vqu085LZ
lA/dt4Hm6jJKb3qV9Oi4zYUpCilApfuzEsIGOcokn0zfCskhDV3QNxmE/o+9lT9F
uf0ZA09lH9QEWsLwRkHFRjti8GAXP0+Y7AnDDAuhePYfkPDTTQHQCQ4TbWOgD5Kr
RGeBGeCqWT3IYmbSj1XU4Xve1W0kQkSitkes1+Gf2aw2fTHZVNbEzB58EkntCrH8
FUdHeQqPVsUu3xCLwnqycLVH65rV2cSqz72skbjLzcJnMPmkRvMtn96wqA7tfPOO
/6a8zMyEJTXKd2JCoI5wg00w6gJziY4DCwD88IDoyz3uBEEBzkGctvEWVhe0OnaS
MoDHNEVx1v0TQHdMLvGo1zIkOquBK3QhvTSGbnBaYnZKByyhMxb4j48eVul8wLLe
npeWl1aruqoXta5PqLxhmkGlhzHoq4TSS9bftWQraD2feC/fKE9KZbXlM7r3hu3e
/DBnRiQS9jcK0CxTXayHMdFktAuBEH7LHBv+nLmL4TdQNCtD9hGjS59p8tDaliRD
g+sHFHvJTfn1PPEMxPX9G9SD6Syu0JLZDEh12jenW76jCPPhmjG2hSKpACMBRwNi
wl0OXl4pBU4hsMjGAYLDOY+wcfVXJU69ZAzwPVs6Oy4W32VJ5aiLxpfo5bLjZsYS
z0mixj8NQ7kjVJ9haZzcpXnvPk+7XXqW/QOfwmQ802pUj43pRjCizriUF0AB0dpV
A39rvpZc5UANZFm/Uq1OXCFjzZ1gNF+KR/sKodgAuU3v8hdgySUOB/Rp9XAqIC76
KJSX4KpLCw4n1E4fDoVeVPmTLuelK5CMF4iatGG0IExlEzlNNHXhW9fmcL/JR4P5
xWOKEm1nsNf8wy0iKdviJ9j4MQEyTiVetQHxXC0uf7IO1Rajy2YuJtK6wjHrq/bh
ds85QwpBD9veSA2Fjf0UDdN00vFVtsvdg8uYSqcTJKKgxe2z/c1mDHMnQ0NnEHWs
ngMGvF98MaN7r+jDk1N9nAVDuvSQmglTFPoriUkEzySOPcC+DS9rz25aWcpl8dZz
o1eUauAkRdc01aPfDy3HHNa5jgdpcImU2uvgC29rxX4/SM/pdErWVetRa8yYGZCX
gFXUGEHVp2Af/X2RCjELqFLEBSqIgbnVDF4DRnQEQ9/XIMdW7SHLrXzdHgyNL3ic
a4WdF+uhehTC2W70B+/53PmhwLbm5GdQRXHDQ3wfShaPDLFhE81c1howiDGt3ssS
fIlmsrUfD7wnR927xYc/WMRZMd0RyXMgFZL8i7XSh7iRbcXGa3pZKVdy3y2vM2JO
p0RCawVCjIzGIUuclK+wzcmgWofAO5W+XoznhmMKHB7Rbsf2+fjSZMKFCWy1cxbw
D5PIx5MxBmAeE6mVtUOe4ODwRn8on5Z24LHQiQTl6F/XvPcEvs0HTwe6EYiFopbc
cUbcsRxQJvuUFkglQkhocbLmfSL0TDINJzheIqcZWK0AdzrEptA0J7sq2FeR3QBm
0sx2xjQFA0LoNYoQIHnngwXvbbca/MKobOcm2pEF75Kg2Uo6YIQFidMvrBxXC5mG
93bjM0iqYF0ET3D8fu3bhHCD7SUk7wpVPcH3N0f8nxtjt9RW8XU3SQXKFulgVG1g
dWq6Z/IFQJgqewg9GtA6znsiCjz+zAV9pxGAd246Wvr7jIoSGb/SeBx28wfiZF4H
w1zkOiRI2QYexobGecoUdshFHem/gN/0tObIGrmMzmNliGOSC/XLaKFFt0f0msUZ
ts8i1I4LY0oT6P6mxBTbDmeUONLkhf1+1wm/r4RGXPxwbw6+/8ye7e0fJV7QsdiQ
XPLQx3NT0d69IAWJ405b4OnOXC1/ocas3MaSkw37rn3emS5gBYmYL481oTqfQahH
FuZWnqmFvJYanqxXFJ1yIVWjfWx1aroirYVzqWedl+HGJqVqQ7PazdsywfFF6ypV
S7XD3+q+xRZnpY0wClCStfZLIjbdLKhsnhORoG2/atMaSL/KDSQJ922ekr/ovzWM
JULWKfwiIixFfjy4wAB+xKwxMj7H5T15rMAWgcHFpvVE1IxLpY3DVIb2gyS8JHPC
Yt+ydWqCB9VapG11ZcaUAhqsfCBaRwRjoQdpPsWBn6zk1vhsXZMj6MpNO0z9s8DW
OuqEEifKRkR7SgIo1orxXScZAPmqCINnW61tEeYgIK0TQCpj+xvvOMNvszTo58Ca
wxyJwfTn3GhmJE9Zq58NduDzPIlzx8eVlZFcy9tS9TCbAk5HVBgOLcD0YYD499En
r9cyxW74wQG7uA/BO8WxyoNYRsJUUyFrlCGwdpQwjhYNbV+BDv2kb5GLn/3/x7MD
yzYS627YT94RLazl3lx7CV+7K6ImYfUt2X+cvhn0piqnaobRT0JqVNoSCsCZA7ZN
W/HBFgY/Vs+ddxBdBf37C/DTFWfVcpT+zeks51fHx3hpGLJp4cAz3Zoim/o18s46
OEioIY+L7HdQZorYPGkQW/OK+JyUgbjs7Wfkifdpvm7tIfs1rt+b8FHeXD+JxlNF
LcoHQpyyc3vPkxd6W9A374Zos5XjChIBrOx8pB83GjWNxPmso+5JiMyKKgMKfeao
cC3izA7LwvMhmXCOzj5iT4WJ+vXweqpJu1WH1HAJvCW6shqpZcepnqVvmS92DFhJ
xWWnG/JbFqCxQMJHexyl7GtTIeRTsI2yS+K1thxkhR8dDgObedkHiDjRMvRKjSby
eLVe0ja+IDDraZEFfHNU0WVOBtrpMzDCorfwWPRCSKGN01nu7IDrozZb3zSYxNc6
LfGLKzDGvoy/Nn5Bcoia4W0AvN1tTbZImowUS5C4mg4Xy+VvYtsIJ7V/zecC2NKh
EOpl0H49sYKzZuCZ40rCoXJYjKFWC9P0VNwx0YvhW5bF1K6XsKn8orbqgA8VoUA5
OJFXgFosVhjx9UJcZ22VGb504Gz/pSqaCf6Xc8nV99IRCK2xUzWPutonK4U10Or+
3VCyjecTmO5lRQOivMohe2IZO4mcMHOK3RjGvLq0uQmz9qUVSEZa9Bt0A1ckmU9d
rUS2iEAIuB6hbGRH5QDFTKDFjt7hJGqeil8AMZNa5NSvn5cOQGQoM7bsYRW/tFD/
TnunQ2e+jfku4WjQTfYmarF+S+Zkjk0Uj9aO3iwz8EkCXQCb5FcDMctefyUSt9Ag
j+gaGH8+3s1RnOFm8XzbSGMgvN3TOgFgKqka6+uwaAwnDbOOebU31FHiR2yHUnD3
2ezOErzRwXMUHWpieZ9acGvx4BxsWvSZprPJej0TPEjFKG92e2FWL4HFwPbYXl1v
h91dQ+SWtXe6O4orBPWdHjDnDxRSkYscIYt48VovGwLY/cZOfRaza2wE+U2C1N+s
Pr8R+XwUeXNlPEA3qZrpNvOUtAiLEvfW0fi7J1a58deE9Hl/TZVUFOe+luJAxHGu
El1TrvDCE2j3MaR2XUAzRyb5GSJ3GvvfQ8+V2HYJuYozqOJknMhTjpsWrlmtE0h4
SqkHpdT8FSywKRLUEa6LG8DtJt4jmba1tmJfP4TJ+lrJFZp/ZfcAvlhhO0/0swKs
uokXkSyzhVEUO46lUWoemq6prRJF5rX9I1GV7gKmtKYkIqOlPzmceJwN0v+GA7DW
JorCUzVtUrc8eSVaQZz8O0l98f4hDLFac+K/DW0Gr+Ah5Kr3uytC+rWf52nmbqgw
Ps4jhtF0QX2MaG3/CEwDh8yh+swCklpIv13Z32PIIumL1pa1rsq2rbXqNQ7U8XNb
kJtiKFWhh78QcGeSjqLRSp0DF6mNA4TEE8DTgFtfM/devKJmh52xZQCbW0tL+yRB
tFLR7MgjXZk1vsf1qQEfwKVB+wcUamt8Tqx1YoGc2E7Uyu1fGIpC931Ar3x9fkoc
rXqLjdpg1XXl1GAAOePXbcJOzRwU0nWOCulKjXjX/pl46kneqzYjnxcGzC7JCqD3
O4x2BrQFY9rpU4ZoNtV+EuE0cGkH1fjYJxQxHtfZ4g/Roban+Y28IUXtYA8M+3hu
Z7+AhW7yS2U1+RvX/mUs8tccH75dEpDadolbECe5lv/JitG1ENVLmFK6SYHTgufn
mEwvE54YKX7rcKAKUFVGQzVYWPK4wm46PbP+ph6I6xA7gDG6Qe51Bo+5QSKrywYQ
EmscVp1GgGrFsiVQ4J+nlhKhfpinN2dT5YLALvEVDbby03BOSgtyp529zn2fP9gZ
OxIe8BktDqRunW9iN5o111b+eHXyga166W05tRwIn+rzgV3WHuYvCIUqqg+DLF2D
t3WrUgL1NONaA8F3fQkhO56dn/dOCH8SL2q4XU0y/yjvK9IiXKLTRQMP4jEc4rAB
BC15td9liFG2hpLB57YZ9D8Agh5338Ep4VLDBCcx5VFXA3Ox9MnDVO/aBDQ9rCea
8gV1mXQlhAciCGy17RxPJ6Qlj6EcqJ7mTqE8pH2AkVNS5bNtxT86REsV6xI5Dzcc
o89qm1cUFWSnATbJTxWmzBOXaEKYPmAp8ZB4O98Tncoa7LXajyOriOE6En5MDvAu
v++1NXJMp+YwovY7rsfqgEOpsHzsteXy8oeuuWTQ1G9TvqE+7wbgDVB9ChUVeQCh
iaiowT/7ntjqhwulmXvob4CJ2Fri4cUz7bbWXHN/9G1kRBkmu23T4o+jMubkZ8KL
o9z2qvqIEPiJ+IB2gtwCH8y85zCd1zqxp4b184m9qc3NphoYJTIFYC4qFbSM2GCo
lF9w6WT86hTNL7yvD93/utq+q8VjiTZU3CEawGdIh/VcpdNP2/ZnMvqekGDG2oRL
FSlZXsOqbd1Yy3AssH90mc9WXbKOrL9VogUV0Tu6GvzJa5vHslYRkCIUJWbnvoVj
5W1TCqjfB07GZOLMOqd/ysTtyT+52BmdS7LN06+Dyqfe+JvulDILo/RUJ5NJAZfT
To10XoZ7LWP4KlNX2Sbw5sGGOQ3lWEye0y9kNOcGv1Vkk9abjwGLn5hCg3zTVNVj
cezubLozvlwKKyXlj60kvKZ6lAiCjaXjKaeMBo1qAcmlakbAPJ0rLq8WhZwMmku5
H/0t9NfhK/y8sZ9ef6cZDqcfH01aCp2ODiw/37yYTZJP4KHZZEgt+1nmHw4QgSpT
BCWUhIMQFOB0ggjk/Y5FqBJ+cSq16QSOvzDVea18CCH+gSDsbaPeTtpIzS+z3cav
+JE+wERgQSLRGnMvQRDJSqrfjA9R9Ife1mWF234lmpwaaYkUGE90SUFmnbHsQ0Tc
1ThKnHcND4a9vdtZXzEYTchsNyz3qiEksolmxIbBNj/z5VcID+sajJepyaH2LNx2
5a/9A0EHjzw00AAWYl7hR6YUfLhy3kiYMfrX1gC7uOoosDrsJ9NoBgFR+TVjUrmk
SnZW8ULNO7n7+r5GOOpAIZwnNDcfUo/GxdAdYtSI4FA0/jK8snhcVRHUmmaBv2pP
A9BG5xdqT05bJmM1Pb4AY6FPj5suYqhyyPNcSU8V8G7Z1RkMthuA26F0n5Vxb0L/
dpG5szIeKi6+ytEwc+ytTIYEaHjaCx4edu0ObfewfIJ1+XwXTsTuZAN9W8r1+gqY
sh5zB50KLnscCRx9WbToM8CDgBFlTxaq9BgOG31Z8C1HKZM+sD2pciiTyi1BKE9I
KJs7GJabhycNP9f6tMfqNyPlBtUverZfYwe4tn0T5onlHl/4O7d4w6aOcZVRm5h0
zQrDD6e83dyJTRQFImAyJTg8QkIWjUcqn5TeYMh8zk225d212hH1RDKNpB3PPuMu
TDgpqj7st32L9/dKkDZZLWP3OWZ7su0zid8llwq3aCiaaLJ7Pux8wee61h0k2acA
cjbs7JAzPCpjlQM7671TnpLCJH1SAN9yURM2DgCoKD5lbRbr/qCYCj5BWyKnOOS+
3IdUwXu4g9qea2YyKpaLmzhdIoAAgSd+d68yocFFM0ihtxv2mHH2aM2pjZ4pWTmX
RFK+bJwrrnuAl1MUFDJL08Z2RFs6FAJc5rf8yjthiv2snahVEXcO37NKJ85YlQ3R
Q70comzvOK9u2PGfB2euU8xy6lxN1xomOdMPn6WGogje0T4JaVFV0/i/RuYK8o1a
DCSwnHQvNaZ+z/EWu2uN+KdTiJl2mBmK9gyFqgDOZWjg5B27qhJvUcy8sz/0ELh0
QsTid+hBRnQxW0a7pDT1pw2toienV7Yllo70s/G7uFm/3EV1VY8ADZHYwO2iSYtu
WUJLW60RfHWL+ZVjwWLe4xJb7EnyHqnrNI63d5O09UOs4GYq2bEsPaXk8ra/e/KM
C+uF1AcJHzqRLxu+EUz/rQp6XbD+eSqs897A5hStPn4yoRukrHZi1q2SpUXKgq56
s4QzwXkKR3VGwGqBCSwCUEutNlEcBFbi2K1v+7PHZQciUSODbh/B5bFPSoU2NROm
WBlkCmuVd7XVmaqalWZb/ILIMRy9dtuq8DS7R7/XJvK4s0sIXEaMB7z8iJn8F+/V
kGuX8Ek//JlMWOIiK2DKAt219Hp0NTYXizy66uA0TJg1Z0LVCsgw9BlSuBtfacZ1
rV8B06oRXD18YQZ8HQ8bBUQ4rL//Dy4a2jqA1bJa4k3Ii/dBzpTVTeXppuzSlqRS
2IMA6tlL0w1KjaBVIO4J//UUOcZobckScQx+hy0KD8Fzd6wQ4VDMgsQycrc5xIBY
Sdd63jJx/JJYV533DOrrE7binAB0er/D7ZWjPvpNGzNIqc1q+MIn2gtRdkJsQ4VN
SyLQOxLnUcGvvkP/sII26elMxN/1Yi31XC2r4YRF60l9qaDoTg6xiStjAG3l+9y1
sXJr6+s6c8qK9BNwvBZZbIwg7wvviywdZMOosbbxy+nNFCnlRNVOs1pBPcb+TK9h
Vz6BSArrwHO9Dnnp6PERUy8Ev42F8P4D+WPlP8sREW8YFRlOxhQhUpa12YLu0SPR
GkbC6vc13aQvQtZ4EQgqxOpStpSvrCHfqIsYbNi/YJr+pJir6dqThzuhWVY9+V7P
rvImM5AXmjuQCmqVtBwWI3SU4rMRyuv+2weperp1Bg1msgdWFBdKqj48VcWxC2UV
/iWS4Fwwop2j4HTnXl1yeHz27mkPxVDZtbYDewR6dA9Z9e1HgeLql98GQRrpELxp
NY+OvZSuzosubBDVDuB6E/dCD0iwwMIAfUs1wK5kWK1JvJDmYlxcyP5pkFFnKH1t
XYY+optdRnG+k++2RJeCR4vZ/yRxP4Lkq9GPt2OtDjbYkM+55GO6Ykg7V4jzha4S
wZ1yjUwyalmuNzkkxNyg7MFTSRi25DFsEmKLHwvw8lZt9V0Z6PONRM6fISEYV8wP
ifarp3hNbAaunoZDHTMgvlsZcZ8LTh0wyVQRPHQb2zBCzTFfyvSOKhlRyoYB4tRj
gv97Ax1xfJoRK9vLgzW7m4VHsUDmuGp4J4SvWkXyC0wZlBAeZksnjz5Pkxhzwc8l
CfcL2UUH1BiwLXnhYroaUYRCqkCNORyRAeRkBDRlKYP/wko+7S5VRx9olrv2VmNI
IxmKEgwGf1DBFzVANuPYFyu9iGlvR6NBZSpZ0Nea7TOK2YpAF0zzKOGdbq+Dr23G
hXCj41U3IRsHAzXDarzxNmS0Y4qhxD6SPnAkiW5txwoMCmmSd+dlnrHgz694oqta
v/T4D7m2qu2cXEMZ9Tw+Y+ZozpO8PkSUne+qVf5YWBtll2YJx1N6dDAgPtBE2Hr5
XHzy0/UFBmI9eOiXRH884f/D6TVYYXq57PWaKOXPxkoU5/qfJnZtjo8VrAIYQK6Z
31aLm4c0vE/kg6SDtandgq8zDFAopuPmgiA36CcsklFktdwu+vv37XO/kE++sKeb
8RkiMrNa/SZVuayNvMGydCQyvpNHXQrD/k9QFqc3T8OsoWlMJSxnYiN0zmckrPd5
CUnua1+WeHCGoA67dNTq4aLUUZ8+9mpVdrRT45KQT8ggLYOo+qRvm8oyk5EpnPlT
wGXwFj0/PxhkO6kFuyFatPdqxiQ/QM9lS9lJFp2LhHATxYlJQR2jIhVV6q/6nu8Z
BMH0dPOXX9nst93rgn2e4PxVsHVqmtvJiP9ZW4oGjLWNq3MT9j3/22JjWfvu2Ilb
VNCxMZgKp/rhAUrZLZw/UJ+6SISK1FxRY95yffbGD6KDFsJXDQQ7AIxkNJ9EJTA6
rD+46ff72xQ/sYWNrHAOM/ufY6GWThNjiUQlEfhe8xV1VCx1wQHQzY8H1bqYKHkQ
Re/KPz5xNRiSsHAcOgvk9rPlPhQK4uLjXeal6Zn3AAxADCX4JnTf/INRX5YxAoe7
8wmvZuiz7XVn/15lu1hbQe6hkDLCR/qTzkinaSb70uLTkwh9gSewgLsxdy20/AgW
UqxHy9gAbb33bvFkYpqoi2Yj/5axfLtysJonn408UCGP13thU1QzHGiZT1C3adEc
squZ3JIE8nVWt0BEonTjxD0inSSr7pl8PpEoIj62SYpLOY6p3rDKdN2RKnG1D9HJ
C8mVGvyzS6XLPsWzOszzbco8gdFuSRcPZ+lronYvG6du5usSLN5rNBTJdy8un3dU
Gl33zDzl8jFm8Pxt1LRrSMLyYRqzA4EQgI4LCXvrNb/JZVZAQ0C8jvplIBi7ZGbg
9VWWrYnurQKP2x1vEnsLhkFY9qVxyJfMGWfY9paRR5t2Yv7WL86NhoI4FPFwoGPc
weFJOtgC6LO8rpU4Io/I4IyZKUZkKYUmetND0khPD2IWVZ2JNItvrKbZsAJe4TXa
ALhdkjBgIH+MmKUpidPgfkseOZ2C0pgjJxe5HY1wrwZQtBJ+sOCcH5buS/tZ8xyI
C8as81GFco63VhnnDcHmXcCr+3GBAdgyrt2NY8smOTxt57/7e673T90FrfHDG2F4
mUURmasozaRJvrsb1wpYedM5CFygsiQw1YDl7fqHM65DF9qLBYISp3kfqUestl5A
bK/Wphn1HrFrXRROUD4Qx2URTvfaMaoAfIlJ3bWLNVkCc6nhYDXPBDZNDz1naVw+
mWcQmSUq3R9mWEc2haZKerRcghEmbdfzEqRivCAYjOZAIFvhZfVpY3mKP61mWT3y
A7XhQM44fGNGfUmIKIHynYP1WimEI+9f/x3ZppNJEsThqx1x7j4Tql/kectE0wy0
SPzTDSpIhqujn6YbFucGkvy+DCv140Zs4hUpPdjxCi2IxO0W9dD/wavLDqsUXk/d
9H+Qsnr4c7uSHakum1YXugkRJly+wxkvFOgw7RABVsJkKVLsl8+NfueFfZzgOS+f
N8reOwT11VWwlI2iVtn0pUff+3wnuv14rIM9fga6C4rybfQptZJE9vQUVZT1e+OF
Y3zHcnZ0xnd2JooLJTmniHCmJcaI5StNazBkqnDxTyAgJObVSpW1/B5Ohe0RkULe
afcPtjGvFd4TyiwVUbwz/WGeBAeV0Oo7tY+Bbb7MgbFwEda0fwlXJxg90oQDO0PH
9PYzLsW8co3ADFtCPi9SKHELyYD1X6Xtn5Tg4JLo+Ht0a9F+Ddnuqk9OPmMa0OJS
5VOW0bhA2jwf+dII2S+dsxM8ngw39O0AEQLFzQ1yqh+CGyuFqT3r1aIiv3eif9ZM
U8s9dPU+eS5glPNqMv/ULxhVzDQuq0kWk5t22yCrUBEBJUiEIJSYdSlKb44wWZ91
5mPrOdTffEEWE9o7B/mel1bCgIXoppH4m+N09ip8iZ5TAiDGLJ+M8kwjhuqPN2tF
FaGCJjxHRa9k/yJcqwU2UxX5UO+vQXVWzBY1AGW2aIfHEOYnXXOOEd+Wz7e9nnob
lT82tT3iMJLNQ59prtc2XgDufgKTSzD7mx77fv+1cpTICJ4F0fg7748evI8qrqRc
K8yoi0DFZUVXcs/cmxdr8TcJ8El6OLSGJDbGFpMoAUIpagmBct8yF0EfnMERIqAb
eKB5yyJmph5Bt/igOimgH+sP5is12IkVDIO2yPLpFpk2wqQwLYe9N3MdP+qjzsPX
hrdyY4dBYM2PA+/hHOVgF2pz+s0ddtS6z+eSmt98K1fBKlcWYWgGMq/BpU13SJsU
Zhiz3d5cRJSLe6dJ2UhH/nQdPwG784F76vwJJ/Qz+aMVfMmci4cyisDOsm9JBjpM
dFL+aNTiW9hgM/feUKtgKzwADZ0iOjsxV4KkGRyj0aFiKBQGJ6fFcJSeTSPt0VtO
95GHpd4fg24Z6KAEmOYXI/Oq+Yk/F+mS/+UaVBnx1h6crmbivAsykyCkvbN9MRFL
epa4FvDvrinJZRmuS3a4DYYS4OY49nqbT7jIE4LO/2W1umdED9QxgaahIKzS2Vz6
2RQu8a/4pgGDodKbckcxN7Zd4AbFA2nPh5dcZ08i8PXs5Zp5rYLyv91bn1QHxMFz
mi1TIDcNhanBAL6hglYiF6gJyEOtkj6br1bujQSUn9ibPLtLF+bx8o2XlxMu8YDo
zEdwsNp9XbOYiRt6McQJ9f7yaDsMMWLNFAjMWOp9MCVVUD/T9OyMqAsoKGXT8gGr
ZzEHsyic2NMbYeNFq81DsmQBVnepDv1/EFrDxEEtFhU4R4EG75mxi59dmo/iO1+c
EonvILE45dO6JuUvb1oHjj0m4zCQGxcNfgaao5NA5iVOkUiTstSGj0fD1Ev0DCOO
WBssr5fh5Tm6A9JrzKZ6YaMMZXLDxWs+V3iOykUqjngl4b16dAsAIQdBfkP0bqO8
0v/Ru5t/2hXWtqDkIlPn5rJqqMjMAEZsu6YQychCWyvoVssLW9dFNG/IrPjBnbs5
tNPjHVA1ldv50BrB2e8Ll26w5EuO9lGR2aI7oHRp22gKc9vNX5FM1sbNKzWhtsPy
+2GEKZ08JwThayQGFv4/oWAGsUJFPj4GJu8Qr6cKX3Z3zgjKpWG3ranerrXzD7tZ
JV98inSt2WfGt8dRm+QDl/+QndrGpH6obguJGZzqTCa26+Ivm82ZrV87Kf7ASZ5L
yyv6i+WHKmidxVSXjgz39nAyS6UlSrbf/jJnT20csRIMuQJRn6McjJL1doE7PVdW
gQCr9GgqAemsBOXq7ecWkIA61JM4IISBnvJhD0NZL6TYrSXdGNHXgeECS10JfdlH
4ONrNX9EwSoBiqIxvp+4XiZhCMxzD70u4hStxADH5CGmgwvn9QoBYU6Fm5sfJjxU
fuF/V0TSCBGEU/VTTcorSv2YJ6vv7K3MriB5TogCvI2k+D7G59pySV5HGv9wWNRH
7cQEWgMpY7s4BwxFERmDOHyACusRo77sFM8L7UkS9YrFDF5tuIVUwPLfLoeu3Bfm
h/mIAQTDLK8uMdIjEq/bJ6yZrhfGNW/W4GjJ3iudfnEnhd44xmObdL1kap8HtE59
MoEUIEkLu6aGvWzTPtO/GMcerO3rWeqvR6s5xCsB2jZTdF2uzRhJvB6Vci1c0iNT
Rhj/N4cwVcjaau77hAbwc/Skz2/vSKwx9r3D4oe2TWVdh42cAlxrIe77l6r0BdiX
QTOLDTv4EjHB15ZGUaozq+nN1YQXFscbgvnm2IDbYEXMpCU0phdhiYDvOi9SPKzs
mAUxBpet/L92tgbLQmHheem4Ggk+TLi++717e4SucollGVY8u8Q98o3CSD/SGjlp
5YWCcfVGRo+DGxjF9nGE3E9nooNMfDnaMpzARPTGXA9J0wezbFVAnmAHHufUgZ7w
SQHKpuc6QdEj0nTEwAGa4srji5ddB7CfvJWNBEIkrQviFRh2boWbnvfTUI9ODuRS
yY8Uvu7a8Itx94B11NAw13ZnOnCY6QkIA2KPN+Cv0mp1oyuVBGqerO60C9K78cAf
Ndpo98WhbXFGAMDtD+S7fjgddxPKKaTiaQMSDo0n6/cm2RHw7mxwT4iVoRoRETjo
Y+fLFg66VK8AD2o2XqrgbHvu/uBtEqSsbkt/BoXLbQ0w1yMYCiT6aLi5ylpfXs65
8GZuG1ZknAxcFcOs4wE/pM94Vj7mPWZCM45d3c3bAS0rP3YWifNWYeSBSgpT/s1Z
nBVsbREpsEUmAJQPDYD77eFdZ1mQqUHVCKWD+N3fAKpaKrgn0EU5VvJ2wdTzSuH6
799BM/jRoFD3AAv08ijVv7gYLgaTUb2ulTAKSIIHUOySZuW1otrp3QMyFSimtRbq
w+It/ZfabY9coH7gg/CsmC6NJHWBj137b1skA4S4AjZmh7+LdPMrAW1LduTqUNcJ
KuCMn88Hz2jYaM263ZzBpR4qk46fVE1UAzx2lsxoItzqawNXHx8NnPLQDY5MQiXc
sI6Iz4A2rqSsHwDePYeN+u/+SrVI1ZaImEyGEGqf+yb3tyHc84kwADPEHI40L36R
iGG6f+yc7HXDnQC1M5UK68K2eG/IVxDietWX8NAMCpOiV2p3kdhpyZXG84d2P8jJ
d9sc95XLq7Ib/2t1zgcAplAAmEVoTeuC6ki3M81oqSgc6lIXTUTOHIXIv7oOA3KQ
2gu1rvJtZo7RoFCaGBpvwu6yuFl+rX3VJQsJmXBsoF76geKGYSzrnyNTsb19utR2
9ViXxsL39jDKOknDRLFNxm97pHWL7Zx4umOfrfSl5Tzw7VsOOLZLDIEGQZYnawmQ
Q6nJEhJVk56paex2LTatXPvx5Gpv4EvtCm70MDd4xJIchugKxlyYkLRyb9G22BTX
W6kaEW/xlosbK5y8uCMfpIcTMSU44QoEtnloG0UddtKuYzlSDenMNKWkZ4Z3M41f
5fAR1Zi7rojnHhm20Zy9sVvaSQ7Y8d8C2w16buePRT8VWToq0OfTVne4RySTvG0P
mxCHlcmWs7RXfa+neqMyrYPwnLpx97y15TYi3qtQgUB9NxqgZdOgUBl8PZhhIZD+
jIwC+0RtczyIMjGAvnMmg/D+m0I7h5NQD1Ci59o6EOhM/ib1GSJLdS4RJIuAlNTM
VByIrbQDOvNo8GMxbD6xBopL9CI30tT70ILm92p0m47Ows2ijxFSbLVc6uc77D+L
rRdB/H+XBrqS53ccz5ip/ofelbzYwIohQBIW37/j16h/wQgOvUQb5gId8WuFSpSS
Juwlk2x1IlOUMUzP007bcbBng/yfxgWy9aWKCWdg8I4zqXtmrHqPRgmF2lZv1zUF
noIzCNXtchxsqR1F85JohouEXvJ+I+1Mcs3RMafU469xlAMkkdA/zUkIfy4HohLS
3AOlqzKv3Ock7JjiqjDnwP3qb5mjE64vN1x15DNcMDagxhn/OfkEZtZHRNx/uk3o
rQ37iERO3bhPEVhDc0GqWL/EIVzrLa23fq9eUS1zHIMNl/W5U8gM8k/amRhOoqrf
6HERrvK5/2sLOJhFZ9HliizdzJOMB/dlMhpS5d//xvCdgkl0ZeSyGtEiZ5cyKi0h
7oz0eoZTd0smHZ4rPgzVxan4NhaWja2EOUmZYEfu/w3DOtRO6cqA6ZEna9zui+mk
JiWwtlUB9sc5Kw7e14ysRZ5MdUGilyXF6w8xrt0QXtxJNmc7cwNXrIb0WBLuav0J
YzNlzZo6yEs1e66Tn3NWH89hodpkbk0QZU+xvBb3YPdgxCiCextD2XwBui/2XLe9
paINY4Yv2JFO8Cw831N8wOnmG3Pm6GcoUVIQTMGSN2CCfvykKqy1yehfBIutXHlF
V0DcL8KHUWxjiAm3DNKNgjrVF30DYJzZOD7QH8XROOIZISk/0Wm3E4NhqnUpgm8g
xl4pHVbn1SU3pyoV04FkEHA86oyydt2+bfeBFkdw+mzbOIzR4NP+lKTRlCwa5hFU
i24U9ZHP0vQ2K0e0bkNMuc4BR7G3mDpRg6A387gjjXcsg1Su5/HFnVWXBVm6zX5X
AYo5LmTpqtxb3Tq/B2tqEngNPxcbxiqUiSsKD3IYauDCUZrF4iyU1c5X7PZf/fUa
97qOajR2zRKFBC1EZ7kwQfaJDqJPhSwOv1oLBscoDsIuhdxPoVSSLBgfWx51b4s5
+dxgc3LZ08cHKvB19eXo9h+e2y+QvirBlImMbrMU7ax6TJlPg7LVISrgoDuLK/2z
4mophvTlt+iEm1kdovM9Oxa+R8RySUi0XhLQHZTDoAgbx8QluNwie9NNKKxnkZxt
RO45FIYt6eRZ6gN5Uqi+6vJ75gQ2F+beVCXqKbx+crOHOHHYhSPtlxykIx5TQwAu
MiAQThWJDNS5b36AOkAiDlOawNx2r24DvA9onvuB0XaBgpQ7VF6603UjSpMPJu1H
Nf9Ur/TnM6JYOwzkP0SIvQFr8tnCFI7K6q3yHX5JnqUZfvkzZWZUJTdkqidaRYXF
RiCFZsByRXkDZe1zu71b68fJ8mzZTP63/uebYdbRiznqKri+f8k9OoT63ES0jyBH
l/BwKvSuv0lHcNq+uoQYQ/ffeWrtKuUwDTfI8cKFSVlrnNYSSYZXm8cuY4DRgqq+
+HsTSeI3IGMn+ltfMTYGVxAh+yG21u2d+hzNRVMCnWzbTZp6vkT2TSR5JCAzu2UX
IrY2Dc9hKKQeRJtKgL1o/0xGAb1g2Ep4l5sWLWvzzZjD49CzTI6kYTBb3UFRZo2N
WCfOmdg0j80h8z4bXSVoG8YJSo8fj74aezQ8rSnPkBIW68O+3JkEpP7WFsbN0y6q
AAvMgfB+DTT4xKHlGZnsXJUEisEicRzMiNWbwYCcAvZ2dFC4v7M/jLWgDV3TZUXU
PFLUN6/Vrk21WqAKKD1tYFCxwYz+vrOwTxdFkUV30I6QNvKwW4UqFqWrNFK6F+jp
lbCy/29qcliSfBuWw71dJE2MyDGA3Ipio9w+Tjyysyw/4Q/vfck1u/KraKMXla02
YJisR2DWzt9kuuaE3evDDsQNNbD+LZBRflqWV+3PhDCi+EoZ2ii8xXGnU9omVH3q
6bSUQTLTKJKO7kbFmL6xaPiWsoj0iVcWL/Uc18Sx23T18ZZN0YBrhuTJW5VCXeNe
p2B6aBi8bTJFhoLu8vPHFjJdOWz4S9XBoq7nd+T+r9KGFdhLYGre7shjr3wY4ua5
vVnFdc87ZfDSAFErJxz6YaY+ns9heDK7UiNp9Y6a4t6emlX41EjtLWtLqiQAVv0t
OaOVevNx9dfZlS0QVPKLrscWaan+MiOlFf4hkE7ad7iZo2cu/7o+JKrUJAppFJPa
dQjjxExlL7J2H7aP6Xnt1ariYyZ5YTqkpKToF1BlQ3gcNJbBCgLwaVIm1EeLvH0B
yC4flPP1TGBiaG6CE9Ixuare6qGTPTAlYmNSk3f3aS8ywL10/bZHK4o+jQ+FG3jg
txWO1d9zbPk+YfAAINWH7I5CzMVJKF6/6Nvql2s7dFd/MlqiRUnO7J4qZ0nD7hRC
Rg/RA6AJEh2arhS0HnWBHj4diByRs1QgJy9fDwRSwHVxNjr19gzKDRdW3bMKCyGO
qWUF2EkYMj3519mba5gPg0BRF5CSS3/plzUA/Ss7hqqMeB4cdbee8bgZ1QgTRpcg
jEODRLJ/8H7ABnnvA9yV8e2sqOFA9+iQg3kSNS0yOrbAHGGoYdrdxOvQDrr6JmLH
jjAdtGSpYNzMAnVfYmo1wIBNdkicSuRfqfKhQrph3xgD2OagtR28TOTEQbYPcjno
V8GEXsxWvCU4E0S7WVPvFnCR3pZy+UY9AcYgoBjtD0QbIUnS6oZHCyanJ+IWhWyL
kzfjk1g0sjO28PIkjvfQycJqfdFj4xVeAWPX5FJ2mU/1z0mZJdZB1Go2M+1czVpe
S4tz1YMRUwB8Ifb4A1wYFGcKSuoW3QuLteTp24pm+DIozanguUQTzyorJXbQJopI
RSJmJa7bRnZAb8P4Z+XkVlIN+phzrTqDrHHn29EyPg6dV9893uHYEPgKcsJWodbs
b1+aLBEbWqp1wJKP+X2kKyb2erGuAyzvMXp6pzwb5m0ZFirzkyGwkeXkhfFAU1UP
uM6WPwqb0hSvbXoMzZORj+CxpLnlWEm/FTijTj6j+PUso4hOGLwLn8XmT/3k6NEV
WcX6pcggm3RRtqZkMl8mhTWhG84EutAWj5MaxHe7f2093XcttdBOY7ohE4ZPJ7H6
44r4Ei/0X2VIpREnUk2SRPB1JoKgqMdeOH9+b6B+q1mm2UrnOl0qK7+GNBgkr1zJ
b8A3Y2ya+anLsqGq59Fovef1STl2zJYygqgWBlmnayBFAiWwxtwMcBfmyPrttYHB
8LYHvNFPIe0Pw6mDPQEciDXRch8c04o1gdH86UjvVjVzu3PSfxrHEkw6cllkEqJX
62qp0qDeOEpohaRIfQ/p/kRAQW5gvRwdnclZErhK05MYndbQi0+O5vEwgqP6RzE8
k9yKfj1AHYrnPfDgGNugqz92QQJLefd3T71wo4TP+KHb2JnuWFY9Agt8r54sOoyb
V46hoJc6Vm56GNlrQ/b4jlcHJtNfAmsBDg4iZJM7HpEAxHrVr5QX1I9KY0AtuSTy
BlzlFT+ZOIvqjW22lwIyVTEDkWG3/armaZjR1EKbDXP6IZW3FsI6t9hS5FRw4dsG
9eLNoQ9dKB8B1BsNLGaJsjmYUH3ONzSEo6l8l6RCicIBUBkYQcThOoYjyBMfXLB3
Kpf21B2ddoSTrhl9zLBHp435MUkP6qTO+Nipe0wjsnzPgcu480ppCOtjc0B/tjVk
tZ6iqekZA4eCn5ykuGRtQvKMWc4RxaiSf18XnE5FLK0nQKDx+l12mbuoTDaqcnF8
9gOoAJyayHfLZKbE02EBxl8ltgN2hUfsfh/7jYk8ybNAndZGQmcCNfQqQ/JuWVxA
lmG2HsFX4BynJIVAQSVP5i2H2FGjdhCPWZWyb2yuYI8uQ1ial68NE+oHmikizqe7
xyvSbIvAGlW/HjFKD0IdobwyR7RA19K85kYKMBQtiOQ1Qf+t6b7Jsua2Ct5CJ8d3
9XOQoDXO85h3Gv4301QElT/VuXIT+e70waTuMg3N57rc40YnnaBhmcbhKjSwNbKF
IhxUGU7hqiu3yJ0t+MElDKUPLGsY3ylk/meiaR1OlJOa102Fi4IcRVd4QsVEk/lI
uM+XRkXJOdZq8HtdmkUECkj5ZxCgKaK1mdzSKUWcQ84S5aHv9fdlmIwd5YGdY0zi
raRUgpD9a70Ygjt6kwFXdcL+POj0Lx3DtgsJWNVhcqh4B/JV5BcG/oHiJkxbSPuW
XX5bz0phUv2YDn6I4Yc6dyB3Bwnqkw7FAS5HILyEWX4JIxko2Lxca4ubZzBoUyBQ
CUrdwmoSFqpsqSkUAfrYvKoZsoNcznBEUmM3nzJ+wj2rzjS9SMn/MxMzqbSnX1ZI
NDF0V6gYGAirP2YeoLJ5qmegT3Use5dPSY11DfRXoGkaKjXNElRZUCjAakiD7/2v
sIrynSfuj+CYXt5bzR9YZqysUru7BwDyOFsmz4VFbsmKf8ePhU6sZPPOBe24sYXn
9w1b2zRYnm0sHJ4lmQmwRNi7volz4c6+nPAgXy7m2qgYdrW1YdY7+4KbkpF0AO84
OQh1310of51bm78Mwhs+g5yk8FfNmSrPbMVQixbv7ZTCjYIStSdQEGK/WhtTkQrQ
IgYtjiWV0WA1mv4YFnfQ1av4dNwscoO6TPcErDsQS+wgrfOp6ZuE3GFF/lRmiPu/
aJSDf7mLQ9miu4BJBqnRZmH/XpNezYXuoou9kmUv4N3mAsE++3ooraO7c3aC4hJn
tm/axwds2KDkcgxMMyTnsC7sV+2KOdGHlNkBCtQY8IVsamIerE+JZqGaHri+ekPk
q3GQiAC6ChEfbB3vfgOvMgObErbYeRjuAWTFktjooyXBv4fH2B7RkAIBNgWe+sSR
srx+LOdPAnGQjWG8za0yvJH6i7YgKBHg0peRDbFWiGRm5UGkBsK17PDc7KAxBuZ1
dnIlkkl/1XdnYyXDckxIguHL1+EhIGyJyTrhDa7cdpzzTzZMjchWTa9nCbkoiGZm
uWnUIk+Bznqs612Vot+VJV+bVTWPNQY6j+Ir6iri5v7fhLB46r4kOUo2OnOOHzPD
8hFi5Urv3UpORCta4LheIOm+ndCGPL+maAmVsZCM/5zZ1O4aSVZ5AXxV7A9lDHL3
lx8rD6Yr+AVeJolcu8sAB+x35N1kZEXny68QGp3w9Cryw3J9amX1S0C8nY7gABMK
d6+CpqqKbN2/9Z+SPHK/Jy7tQfwb+Jz4pv2yLFlRkifBdd2nhZNSg8iGbp3A5cMB
3mt1H5uSmVUtqwxEoYcTQOyOst9X2pfhpRJVAQ5cFwxWTasMTDde5jVnQtCzN0sL
NF43Z3MKk2FUuGQzv3Z/xnskEEcU16by5t3LhBHftB6sAlKMrAressZ4T7nLF7ca
L57G9umFpTHpseu89YdNR00JViDAfXhVBPXok1i1iWx2R6YBRi8q7FaQwGJHlUTc
0C2a6lA1ass3j58eOLysMLorhX6iCA6kzoZx/+hOmQrdk2TucM8Bixa19/KE8tXg
0QfeciXxCK9Z5OKAq+Q8D+GfDYrn+mC4g3RMYpMDBlh1YEtNxzRk8sZcuIE9eMEA
Y8BdLQFbdwkrLZxcNEz/7cfYQ/whHsskR+T3Z1/aN4LkbkXv+4sfRYkDiAVpM2EN
+KUHGewlkz657sQwOx8uNHJggKWkd8xWps4C3WKA8z558kKyk6Be93qxhv2MsZ1k
8gClj4uGuwEp7mme3I4uDpdIBxxk3iSb2BVEM26K2H32MxFG/xZ6JkgU5QdXU3cD
PCo8uaKrEKuE8BT9IBuoCvNS3omuZPW7f/v9RqHFYrgUHIDQqTabjvGxsPGQ/BBE
iWA2jOkf3dW10poWZqJbeKabQyp3jDar8HAd/ZQ1HPbStLa6NLiDCTI+2tKs022E
a8NIoasvYolmNzRyZ8Yb3Fb/WAhqd3P6d6byfuVY0Y78ebO23MWGzja7Q5F9hKN0
1Y5oPbw3RZ8i2D4aF8G71D6dH+bM99lWt1zrQpRGiohUkNsCCFcYUSfSqU1lSv1P
9tYrYwuTBkb4YSPwdZBJbd/CvqslkNEcHK+ONv5HcjwxGutAP1WFEoxX1okqTGlP
bsEt0ilerYH2rg1z3Bxt3uVtk3gDFbxG8YoYAlQSavsR4K3JaVXIBeChRddNKGVI
Da0/FFnmuJXs5IiHzMW+p8BJpZ7cU120bLkIMu37LRXssOCSyOI7OgeTJkXPcLWN
ttIqBQDhMsmPps7PUtQ/3pjGvwNXGSWmWeYujG/p+pkB2/+RYYBCM3j91ArxBmlB
Hu/R6+vZjecZN+z4uZL9dhoVghZ94gxwHrddcC/VxvQNUXxgJ3qwJS88Xx3Z7TwH
85hAK1J51VSz/QJnJsN79pAAltls8bXQ0A7Duj13hTszPfikOfSxnPGxa+1dS4OO
TGgXVZ9z4Oru3INEXrhq5b78MidafndE69ttMgm7XWj5Odmo+jszJwuclU5M/knw
wIkRG9oFGNrPC9OGBO0g3l6nBjGRdDQASFUj8VoYy1g7AbwD89dtKrNLOHiNwIoo
Un4DOpYm4G1Lk/zGuIpXuGjBRCEdsc30W6LBCcIjL9AMc7jr1mmz/2mLUgWTWONo
BhHYavdLvKgeZ8268pFwmPynHjmEfCr3E3APF65koMmlcuKTH5WkVRmge0EBjoIE
HEePD7+nMw9BftJ0UGzZ2jYGeO14dU06inRqSTNefoVQAEvF59zrhdgyOzL1gELJ
K49jL1G4Xyrv4hJSoUic4RGkIzvnSQMsk4KSx6fbKrsmA0yQGijt84f57zach1kk
1CKvSqT8vSBdm5mszdoKia9kayZtRRhsIG7trwZS7Hxby4xQ8pacV8IJIifc4xrZ
BjfKwPGeptVi3h0LFsa1jBe+G39xDXtvqSAeGgTb+IItvOOLM1aiUprwO5QuOgep
cx5HIQSsAo797LqQtWEfJi8TLes1Q54Ti+KQPLzuJBVpb+/btn+xrMLNTOS8a7B0
8mgS5gcUr3B/rSpvaSMC4EZ8cTFf63TMosX0i44FUC1vxYpR7eHxl/OwOc+ZxIjT
hVchhSl7qoBjhebJ53/R6lIk9dyFKn2jGVfvtoc1aWkQti0GAlIqD95vxd9ADyZc
PlLHlrrdUyMlMWTb1txY02DK7VWDZHZB/d83gK6oXGWPNtKl5d/yAy9yX69twVNa
nIwozy4AMaLmD4PhloU8GVtAoonceANeaueHIiTdorwiHyLcv/aODUrJh1ec0AnB
O/02LmYADabc+dj9kCS98nVb/Zg6GxE0Z5pijDMdQ0+V2RET5edxOFm47JiPMvLd
naqowi7vkl/BaPzVFjZ8FOdkxm0IqzOgIOzn1dvCNhnR+sh4Uv40EV3H9dSgf66l
7R+UqTl0AWrEUZeyXad9Z486xHcB8jMJtiHLOxHeLZQ8sw8Xr91eMR5/JckEuVYW
yQPwWQsWjv0EcGHrwoyy5eV2Lby2YSQ4/d2OzcgWcBsbT6Cyvd3LW+BQjIPiacM+
lt03fNCzWffG/1oP9+PrjddAvqoMZnip94hziRIubn8RgPOBKtq0a8x/A1TV/el2
G2tfr7n+VsljBBY3kp6113UdATT3dan15+pBp+eojbjPs8AQtIXJl3b028+FNRqb
RZunwe4xrSvOn4LV8Pqe4myA2qxYvR/1SiiIQ0nh6M2IAJ/FDYyoWrqNseFuggB+
datYzCTvAOm4frOOl8TjESFlFj26g30oMQTV/yU9XoNR6ch4J9ejvOcclC0KTpXo
xWTqUP6fM8JVH4Gg+f32CEaOzTSQPFn9GBCd8vMPdrSqekKVGw+F2bxVU1Weq1eQ
HqyKoUSexb/6y/224tIXocruS0w1XUwdauToPfixOGXlqbpbrl4SHNXFFZcDfEfv
091SWcPafA3DpJtuQbNAhW+t8s68PjUmK4dWjMKzakAzt+yoaQOXbnQMMHxbmD7X
lr0pT18wt7f4ILPjs4FMUO/9Rd5pMtOHmcyNRjkNiKDMp0QRJgWbNQc3W6wHo+B6
oZM36O4mVfxJa8NhZAPJuef5qlkUO9oleRy5vZJN9mORPJ9ojSeDmpKHUE6aPXzi
UCNFtFnp7VvNN2OHasjuekStIfukb0KH87h+P+Xcql7/QBwhiKzVJJCOZgb3cdSe
Re3Pu40MbNUQcJf+mm3OOdaMJLi9OLnnyd7ZoebBvf3B4nQvZtDf0/Sqaspnc4Xd
TVtffcUw3jPLNq9cFQ3pCkz1zeTth2jrESh3kB+FokpPxi4h43r7lbGg9TZ9H8Dt
BeDbr1nYSBwnlhnRjdD+oaEmu9LOp0jiR3VwSphjk950KgDiU5hu1drLTFgboJvu
W1lJZCWvSd3v9EuvK7Z7ICvbOXNC8hM1IRTi8YqM8MUHwac71uC08PvCS3yNdkoY
qAQ91HjHjqyaRyjJ8rG2MbdXbhcdJi1X2MiayWR6udUzXEkJyZ8ABQwCRJKbuOla
tJ4YEnnXacBmrVv84c5kG/mpxcsSZAgIheOap4VrW4CI7mfdztTldGH2W68HE1rl
YxtIk9XEWq6Fbut0OyyoTfcrLTQYj6T7+LST5Z7Tpd7gjnFt3CBCET4vU+JIuz09
MNZ2VUV85x/uGMYZ9DtA7eDkDCvwrEphrxJku6UAypUmt/NMj7WX4tGyPN+tVmsx
mMo0+OPk/X+LCS0izV/Nq5DKhooDHlm9Eq4a8tyZPROfr5tou7Co64InHSkaBIcv
c3tBtrx0KiAaLK0n/qVJmyQxvNpXAaACCJFBM4nf3rjX01e7LPuhBHHJtFULCh/e
2NW5rMCc00xp5kagR3Riv+dvmjfLXVrLZmaxl5ND7P3GAf3xcOcPeqK7XWY4c5is
bXDw+glLEhWoUCt/97XMz47qHUkqT6H5k6GbYkLs0QuRrrFmtix1ZaqiEA2I90jR
59R+xVwIzuk8711wUz2PiCQZZuSEEoWHNpRGsr9cfFTMi3Dy7h27wjzkaLJNa7iq
VSZhybhroYCBSgksnJj0WMZ8TiRU8ojGy21zqOEFZg6IS5HD9Hne5MVj+TYmU9ui
6Vv0GTQ6/cEDLKphKZDI3akn9CVT5+F8+PfR3gwwaju8PTCbb2fKmVMV0V0R+Kn7
lUNZgEvp6l6+n7RqhElNg5h0LzNzQ/JKH+Vln/nmUsAFZYO9gG8gltOR4WrGv92R
due7Zg/b9DDNMr0JKMKvwgemiyIKKOm/66Zs8PKrMYW7xnAlZcUpzDG0RG97ZiSz
c39XB4cqhztza7HMJbcRG9mmvfakdOnHT768+VW9nTslX5LeAHofWGNN+N4fJScA
JqIsyqr449vCCZ1eavisDhihDfcMG9EN6m0J7ytCkoZBdkVBa5hW5cvKcgOQEjCo
y98x7Ua7N+/63lXfaUcPBiYGNvRY7rzZt/eu4c2nkFDHe28BZtnCKrQ+y+3DAk7y
Ob9ZpclpUaebZxw3jG9cRXcdTEVYQEgaHJeckOHlZc4EZrEpDQ3GylVp7CoHR2vl
J1JK4uUfsdgjs/ePNlAfBIPrKf18FFX8yJGpbLS/5iO0N/qQIUuaOxdRKnIFB6KU
HntXaP2uiu2lSu1k3z3p79JOZqNo1zC2MriRFO3eNlH8ubjGrJt4Ixlv4MhCJRqN
Uy5Tmhe0J/TpmlE5PfzZUiW3aOUAuy4J0aMnhKeBbFr0q9sIm0cg+gYQSRJUbY4g
GgqZUe0+r9pWhkuiJFNIlDlfIvYrR7eXaTk9GGTJ6lGOAocJOScXzSvc2zklWXul
md0hihLsHF354kIo3Kx/pnM6/t1MbsoXg6IAtM4Oa1Vgl5Dp9igZonfCaB2AcG+s
UAziwz1SM1evOOFopd0mES3ISFaR2ZRdAdEyRLLzA2DymUAbryjYgD3YW6zugxFd
M8OAbLrGWVeX5jB3QBcz0oFU5hm4IsGLQCcjUG//2cae/XFsaDdm1+MRYAuTyo83
8N/3RaIOrtRUGxBPKGNa6BwRJr+MH5UCQC+8Inl2pPcJmTDFnJ91Uf6ulInTZ65I
W6i6rVwVg/GzVyCSngJU3Gnie/XRMIF48sWM3g5IDumK1UVyZd1bWcYYT1RmMocG
TLsXx1qA/9vsYh8OX7nxeVhTnMkS9UM2GEBaKhT9T4Y19pmLChrxDw7sccrJTn3q
WcAvVK+QkgMso1a9ig17kxgT2CbI/+YNg65PogcwgHHyPG7FTmWP5nqeuT2RTpOG
kfsF6Vye903XR20W5LsoZ96FL5UdxanOaTMR0q1N9WRbQg88n0+sse7yVN5HXL0S
4CYQ6yOxPGXKoS4KkCom8wil5uCCEIDeSp2H+8O9mXamyv4HnmYIUkJ1mC7eTfwU
WDQPLvNV9qpuSdNgu4noNnYLcRIFnkePKw9D9So7Niiq/iQWTqK+4kDqTD3ebLm9
WWmomZJ2n/gBfAK7WOhvCM83/qjHEOo2YDYsJdd2tf/Np/LRw2dNfK8TY2XYAOyE
j1c5jCqhy/4cac48vADkELy8c0cRprKu/I3yTTfXBzNs1ygenxyBiRwqrOLS/MRB
hQ40sl5W9zNl9FECKDKF51CawipTG0DVMOv7eJdTzsu8yVDW2VM3Wrj6u8eY2y6J
gjES27g3+kkSJSCEQr8sE8iXL4r+LXl6OGyT3agn15EIJ6ZEUZNcvp0yrSA4Kmlp
kl7EsESx5cm233z93L2Jf7REyVtOEO5k7qgcU6JBv47B2gl86siebgbRTYuQI80y
FliNEyZpQmxtuwElgJpenz6DD4VgjEmtwOYFjA4QMHyntDSyb8ewL/vvKmBkDsA/
0wvpYhzv1hAChlNIJ8LGbWLaPU34rd0Hs58chJort+oaWXU1v9dWHkM3b+LwOsbx
1asc76dbAbu2Wzlh8ZV09lAruQW9JmZgRPWxFIqKTwwZM4tg1R+PsJjFW2jA+g/v
kDpo7IQYjpyl7EhRAMhbeIF7BcrXqq3tqMiTqR5C77OoSLaG/3g2qxmF7+az5CYq
FLP2bPFgZsLZR5TNyj9yYkOMKNMigfU7Eju0TnKfCHPD29Vt3qqfUVzJd+2hWNFM
RKxCpzuG49MtwCy6bbRfh3w8ztwY1MLJ1BwGTbUujfHBWX3Op96uj8VmG4Wu8+3P
KzZVLUDrKPeom8MjYQY8UC4SOXObUDrSKANXghbk2BHrCGI1BMpZNwYEThvHF/+R
rl2nWhIaOjgkF/VC295oSaYAbX/RxPsHPLkGNvLqQj298ID1hcYOqerYcCcJRXLz
2nv89ZFWPGZAeZf2gYWXQy/kvRbieZxgzZGyG5wqNLk52iXFu4kD7QDnyiCtAkNN
x64RjUM0/Ptpnuf1tuIo/w5++Ofwoi6N8fsV2v2bsQSgEx0kkXNhLJBz4rH6owmD
C0ehn/WLx5r54VlkR3QVpMDCqc//5iQftnEYLqnriow36Xnd39erF+ugyswUgv4y
qhqAbPYxmc+bU00fA5+uSN0+zo8mUzoLuO8EyxtnusipFZUhDnqjFvfGvDQE/kIw
JhjUE+Alathy3kBADYwOE3FTwfNdgT6JuJ1iQQfJsVaFaDXTjogJ9EAoGeimaa34
1mH3PNqkMF0PipJ8WbY+A/KXHSu0QedcpSho81wnDHp1Fr8y7KlF0nCxEQR67kFp
7gaPlEpU6lrD8mj/5yxz/YepnijS1r50YF5GNgMy+w+IBnnxKYgMcQM0QHqj0JJD
tvgpElifN7S5m1qufmEDSFYBZNL9Lt8qdu2+WwzhR7DHkjSPvZvZIpSFOIriADcN
0bsIuv/KUuHDnwT5Eu1nvad+guwes1XMvn9SLJUYPmHQ0T6v89cyk/RCqOEoD91m
yZcobIw9G0KB8eVfgpk5NtqNshPKkIkkCblBjcYLPlfuhmXHdTqL7kFTrOs12c9k
qbBfxCZE9ie6ZPzv6qsm85hqfyP5dw17ymQ1sHVu7xnTXQxYslbByICsNx5V8IVc
WeoP5ZgHr5r+81dyd5cRGGBMYy8yZvJrpuybj4+WFonLNnDv2bdPL7+VlQGBI/3a
4QHbK6fdLEcquKIvKm8QxjC16rsETGVELlZhly96ldxGkXO3nVhaW7UCI7FP4dhc
iyQjqY4IBYPevutFRcIGo1/ws74PvLtup+Lox1C5+YehvwyMd3SgishrQSgSs3wL
GPrca4Uzb/24SkMJR32QsCKwKzkIhtwwf/AKAKK2RgZCrfIWrlyj7cZPIbAzy1WG
P8FL+77KwY5T61/+BIfOufPSFZhjEfoaWkcNx37u/N7INkzLd1buKnDdKuC0ljlf
3SHf2P+ovusnCedLOKdxWymwUuposLjG/24HxdbCwSdZTZeDwmHfhzVxheLVE/Wy
c+B2/9ONHh+ZEjPeA61ySdG/buR118HJWUdsfceriZzfpD9oC01TThjj99w3sM8+
f/m6nQWw1EStmufCnvy0y+ivwhloMNvwzJWQ2NrfaLsCg3TjUQtx70AbpO6FW2gz
YIHWgaS4dXq2NhWONYqtTzCiGz5FPSSx/l7f7yDswCHScHI4onUHFANq37DuHfj7
1vBPRRVrSC7b5a3eJ7OOYrE84NLZOy5e/SYNY08HS7Sb0gY8rMhTgklhIEjlhkZH
ig2raxG4za0hQ9pNZMXGECVM953dlA4F1amW6V90a3mbVbYkslUtnV8gvjAiui1y
YFsGoK6UkFPPjY71ruignu4Lb0FtZbNekTGhB1JxRQLXkRS9qp+JeXDwIhQtHbxy
Okj6MAkP3g+xhIe8A3THg/GsPJ8lH0gx1bKMHnjE8ZUszaF+UAYGt0zvmh3Bxyg8
9nzTZIvUvGI0S2mvpPsrmPk8TDgi6BQWdTt/rI/lYfX+gr3KZTw1rUfhma8+EkCg
Tf2MLm8+6Y25yGrkPVgRZbc0LMs+P3r7oH2e27WIY1FB+lQ6AJjf6TJt5jnAqUI4
jcGG+1uJUoEz8HNyrChOfg2DLnc5jhoDUCsn+RnKLxQ0LNCeuaS2B+MCk9/ZiqhE
mr8775PfTzeaYIrUHH2QpXOa2e8oAgODXLw+TGuMojBUoEfIcjm3jf1DemWuGLBJ
YQn/sc3p2Iv4oN+mJ3wQyJNxUXGKkL8M95ugu7gtOXOY3vyTrAU8XeIRv2+h47SI
xwbrSnAkYbe8I2lvyFOiTpktEaKBkaYYWINa6soXvzsu70GEjvIZdEXvAjssEK+J
uHOmQbn3YPZVPk+CsbK6p06R4TndmvYmRuC4uSxQkXuuu25XmYxpK42rwMMP6GRl
yALPsLXb5q8h1j/zUM091yXZTB/XcAsWNPpYTvjox+tukh6yE+541LCfaEDF5Q8g
PT84j5hFD++VYDJ8tKAF+GF6pLg3AfRRNzsSSMffezinABRh1prNTQKUW4cwYevK
9ac3B17TSCS/uARdtBWVex73wpzLEOPpeU2hZQHp+sIBFp3/LbYJLuulliVgZDXY
0d3NF+nxoW6VMkWeNfYL4WQ6TybVT4H/oetB00buZwKOgY/i4eni8UyE3pGLnYWg
z1MeqkYel4gp4iG+MfEOCPbSq3nEtL2LxSdKEhdDlOx+AfwmqApFf4mb1icLoRo5
ac/b23PfrFNN5PLmZyN1/BodLMhycpinibvzaypkCtO54ZurPhXHwrOGzYvnVwUn
+K88a18+0s9oF3btfijxOOUHtRe1WBQd+2Yarg2/haHaZ5EVh6IdS5nktwGVBBvQ
W4uouY22WvQrPsrBbekQo5ZLs2A1JcYr9fsFgAu1GrUzvLVcmnQxtJBZImRyLJzX
xkHhpOl5CjnKOkocvEnmlLxG2ChHyzpSoIPFv0k3Qct6O76+lODxpcsz9BJF3ADP
nPmJjNv4PIAYql0YIUuKAsl7V7xQcNymWyUtVvytEvON10HCQiVbQrSfmOggLRRc
ChmxlSwifT5BQx2XgfpSGrhwOgr8nITCALD+Fd7Gx9RRegt530DVpNsQR2dOHd7q
UwW5pt6qpooUpyRFrg7leG4mLK7nbxGcehqwlAA3TyBS0rQXJIvaed/PZNQKAo6f
bdUpvS2VdxJN3XFZQI3QjYYCsfl2HaSMEZ3fgNWVrutSx9Im+ph58p/Ha3TTRIjH
Kca99xnlNfhrSarrKTpBlB1GlDDEmO6u85gtLIoBHeTb2i1LsEBajYU4u4RXf1ct
lNz381KZX/yACdKgK2VUKNJTt5YackVOixBOaf5UPkp5cCxCLYJQZzfflOkEWi0E
GLnz9dIwZDD18OVsQRU9lxo7AL4x9zHtEvIb3EjxkjniPfHbxfz29TQ+rrrQOlxY
IH33yTeiB4sByiYHthZ+njv8VcOafc0LAqls9Gs42rfV8+7YY3ikpN1zs8jvntdb
c30U/PEDZJerVJ+6p7ajmx5yIOKBABF6QL2bT7sZtE8EGnNywiBvEOHMlc5fJz7S
EzkqMos5J41G1foJKX8vUnacgCd18F+RlV0NF1Io+/kugUu9j7G/tptGi9ItvQfO
xmpFdZB5wzr8Sc4UigY4ihXjhkVsNfZORnQanK3KCVWMf18kAYqTKNn/uhpJYCYJ
0RkpIKcJX21K054GBp+i9bYP3yNH2aqk97CBaHBRNtWP83nXTZRglIvecRkzwzkn
pGpaVVnA/XPbuOg9j73yYYnnwSR4xC0b+cGYuqXIufYu/Wh1uaFM/BFH1tOosokW
nWQmo5apvfaOl+vJe09km58Ijo9y42Ya9X98QP4X6xG2hs/SWAkHeQZ69zl4r7ka
+jrXPUcreO7k+cWy47tW69smu+vAweElKIxhtybhB4Wsgx62j0ctErXFB+igs8zS
M1WacnQxtOULiqjH7rI9jBZhkZfOW7dzQFuchp0PvM4j+ekblYysASecWkhaL/60
gNwmw8cTquA/vkzkg+WnGKKuxU6Wgqd1SpNokiL7Rz07AwBCLyZMgf2Y+2o8wB6q
jCwklReeXMicjORxODrIxhyHJG7a5+NABRQpaZWQssficsfN1GeRbBGOSIOMp7v+
/RkvxhiT9HInaPac4zYp9sHbZCVAU7mgJ1ab2UKPC78m8G3QLYfGIyax/WvDCrJF
uzjxXqIZqVTB6ltNqSI1HL4s7odqjRsXYJofs+F5XeyJynd/ApSahBdxbJftGpzR
WVEM0EV6jeExd8XcNhR/fD8R7+Q5PLYR5cnlK+6z0bvbWqkv1aYM81q5fFHkQmUD
7q46tzaO4uHktRlwWoaRB8DryCdMxrOSDlup+Um5po8SHrKmpGfYVeeSDzonguh9
+K3rmV6wkbqikgg7zfCNXF2TI6oIfd8h9JI5nPwXdM7KDSZbXWYXRZD+E0TN4dXc
29mmjkOYez1mTh/6IagBw4IRqN5QaeGdIuxhR+ycPAlNWLA3CSaRsbpHSNztKOAI
9+mvps/zahn0kb3y69QBlOTFdroQ/33lPCZtK+B+1w8IGqn1SHTmqXEUICXRhK9C
/htiYwbTyfJI3NkYYrVy4Eaws/vpBzZq6ledkR4X/7Qh5vJbWj2GergBMgEvZ+sn
LveHyZY1qW4678YmuQt8kwy1Bkq84tttjO+tziFKnwwGIicWfAqvtIahiVfZWwlB
xl84dwyeHX4Zkru4b3HM6Rlja3GMGd2qtOd6smxN8nLjEA5RGO+SV8PRHPXOP9Yx
Q4H0JGFiWCuayo4Q463OJlcUKyUAAXG4kPqmfY7A/Heofft1mt/2YV2e9SDVJMAa
hiakCDFeoCO2z3TtI/R3RwU7wmsULSfIM/CHABOQfUyApn81gvUSSDigJJ7eeU/h
EWiRaR1fPgYzOXuj8/0pGvchloCzoj7LHpbBcrHp/DWe1KD5ZvjJHdVeoMSirv+q
DrjIP8zpdvrt2GUSCVE2ojcuh8Zm5uYtA5TmkIon7HDiOytxb8+cdB4eBWi567uN
zyqqjBrBSg43x5gKnhBP2yIay5za5jJ2IbwsTnQpA93w1ln8yjpe5joznmEOE37o
kEae2zqUfMV0w+YaiYiRhMDdqyTOSq3JgX7D6b3XqBEgK5eaylN8VESVFpwX1h87
N1ykx2b4TMWqOenIFBut55GmgCHFSYePiN6u5TBNjHMCxQu0gJAVu5uPqPsH2Gvf
W/yy21yP4IVqp/zTDbAShz1SEIbGurdgCclRGp0Bn0NEPOlneZV83zcvlCKg+Can
LyIkG5YCqSNdbf3RF73lfrO+5V91oC6YvayWtu6zbA2u0QXsRqvAmw2tFyKulY+K
NXEjh8Vge+I2mvikHOEFa/VKEoKf8LPBUoWmtKmVgAj/5jdU662E8UzumNlZNorm
PcbCaA9LwvlbmYNf2J25/BJ8VA37q68Brp5WAuJOJQxSrpq/6F3o9ZiOSf7kQpFS
UgFH3vTUea8oY2Qm+HoKijziuJk5VGKJo3swLzwXS9OMUgwnHt297vGsBEGso7GY
4uzLL8qm+69ucmVLJWQLb8Xc4QXCZF42qW8repWnIgUJJzPZJCC/+FrMc65wxOU6
rez7LBTldS71VGIaEvax7pJ851iCzEtiSlOs64j5W90r2V21jX1pfrnACwr0S/wF
Zp35r4Hq9SmvwvZArymx5kyc92aVcKlK0DLA1KxWzVA4ese5tJ9giAYXjjhI5SoN
M76YBLdCWW2UJn4cLfWmtDqSlLFT9XXYQJBgdVCOvHLbBvNLWk5T3J9ThF+V6ABj
sWqBBVZbZaC9J0KQGUsoQGDcSHItWDDINXPunvvACTtCoGcT99mqArCcifef3rct
aizZxyxYhEfE2CDKDFdFH8cz34KCU9zAJtT/paC6QCJX6rPc4Mt7bsl9VdgIAsuS
kKpiYOteFqCkNh84FLpJdmJTpVkby9eLkG0NzMx90tSUpcoGZv3E+pXxXGgfsKh6
giyZ6UzdWob0kDnA7e83UwGyeEwc5r0ul2hRaz8xZVzRWZqVIYzvWWswMhhgTPEp
l8/1QaM6YOKZtf4/q1Vong8O6Sjyo0u9dlyawwTvEwFbhnTAcOv4LhJT9ybdYqqg
MveuvPoo9s6YW7A3IdmtdOx8DPP9Do2kN6ypIk3OW6+oz8+21vCVMS5YdinXtyMv
PpWXhJbgyGxUMWR++onXsc49vMckK2ojhgAFb/VEw/V4Zr+3kR587w6DqytiIVuv
me0N8bipCJ1VSTI1ltCt4z/DXpCEZDf76b4bMorXz2FT0NzJyHdmUQXu4/N0fEvl
ZMuv/XRmZLHbMCfUFI75Qpf3o8V0kAc13K7ApUnUaDYi5WlMLo1qdeUolH6aMuw9
ujoyb0CpvZHSQs/HJ5ybP1FDOMdAwci1FgYbS0xD51SM+H6RRspqznic5zyhFSGT
26bk5rHkAEmE2z3LUM9yF2pqqzVNl+ych6UabbQEw5p9Pbr6yugjbHsMiVeBTgbL
+WbQbecCKyF56yr1xFaV8AKnyRPvEwkdze9W7Og369t4Y9AUv2sbALkEN6gQMmua
TP2VsyfuxsW8eUd+nyAIwCloDUbzdJSfz7P6lx/xsWWU+lE1s6FXBel9HFd4RLXT
Xoz8/FKiqniWLZsLt+N44D/y2H/FIVV56bjD+4HVeLgLtuA/IEr4Fbgp7e0ovIV1
c7KgmzNKRiR6XQ2W7KpOmHm/DNlLCYeY+OHxOJs8Kipy4UW837Q5ymRwIhjQmdja
BZ94+HkaVuPrVPfgbR0E502ypN6wQl5xn+DLbL4xDHmC33icpPN/WSplYkqy/cV0
Ch2u5cB0FAhu5Fgm6G+AvZbNUhg/qXLQvN2f06kSd0fkpiZR2xG3ZTRCy1EN/Ja0
V2MZdZHfSUgNXKWAwkp2qvxATQTDawGqB7pLxgoUB7bExSvUh+8B0z4Yj0ys0GtO
lYXH0kuDmL9s6DubqYjE3KhedaKFc7SKAL1mzijiMD/ewqD5dDQe1zbf2HXY/LtM
NjPlgGXd9Liets/G4G7fGvfc775j6w8me8LbJc5udpVHrQ6V7Vf95zHtUtdt4zvS
VdCtDYZD7hA2srKfKutZpDOL6w3nXQlbNk0ut7XlLK3QUGPyEzZmGDjQOkmn2r2o
Qq6tJgQWHKIgk9AiX0VK12KYueNv03/cpNu4L0enJeIjT+idI2YSPvCIzpnRRGez
VbZUqA4Xxgt1wXBIx7Qi3wjo5oKCgXoDzxtfEufz2Dh+xy9mPKVVG6k+6HIECEFH
mMuaUjV5QOT7fHIJsl3WmEp+ZXwEq1dPpKaVbRnSqW+KJ5u9/dQerJTJLj+0s43m
9A4m+YLQwHPwYC/++FEvrWlfq0VmG+KUTrUWroB96vCg84rl1lrZvIIvxKS8DDUQ
sRDAz2xPPo1psYLPhdcBQhXUkxwhWJNSfYY+YtQ0CPDBFNqfSFEI4BlYSSQZBqtD
yVxECRH0kMZlCDkwvFzuwQhAo5l+wc91J7aCcMRy5KbR7ahwCkSOadgvbH4Pkorh
3x9SDlMeIFpvrcEUm4/1Wf92p97pyszOxCExnuE+2DE9DnZeLds7KByozizdreuG
nFpVH2Djl6rBtz8LzYhL5kSFx6zBzIQbtm8oesA64KCfL0UOaueUoiqSMCoLvCIF
0sp5DJM2Fl+6zzDEe9v6xrkHf8W4mVOsQQNuC+MamA5BqQeECqQrh5eh1JX8nNVG
zliGcHC+VJlirjK7wcI7kRjIWwC+Vb8KgQwBInllDW2/+TS2Xj/BllXx4I+DgI7S
yH115nqKB4hE0Udx2PDq8CcvzWaZvp4JcNUifjyTadGWZIw3MgMKjY/rmUw2zI7k
rnceqh1XuotgjSmW03veflF6E20iFqYNXwjgwwV7ygcmIzD4pUbU/3S0ptDqqexQ
FB73w/XShAMDlmDdiDsXy4B3mbu1XK8rLHuXKS5mgCIQ+761/G2DvdeqY5BfqXQj
ERVzNiM6u4UYFt22cXVNJ4DR4uF7HIfstF0RHb3HeY0gx4CWas4OpwqmfAlqLWtq
9/Mp5f/GMKBiYcS95WcoYZtswVFjOtb/6WEM86uedAQRrfJuJ3IhBkX+ErD7NNHt
QMpc/30rP6sZfccvLBv8E/yHnlZsgb/xhVEnUBZTeEZC4HAc7Sr1bTMSnRG6G7X+
JIK0UjR45dRUkDLet1lzfaHH5AC3fDJ1lUH/uxuPG+omBwNWRZLUSZX++wInz8By
xMnrpWTOpCHOkQOOeAJqjgHphjB7EJbGX+V0qXEvUsQ88Yt5NDqyhrx89o99Gi04
tRvCm6Yk8r9JzdAQDjbyT1N3vckmiYG2qWKn4hO5iMXmGujgXAHTGXmVGqn0SPWz
rwEYQIK0c7wQVLh9ooqj4UeYnNI7ONcWq7EgEvuaxGBzsDWwIJ2K6YArVHGcLnrp
/rsaHZm7CplIQpEmupsbKW+A08JALyJNnkLEmdutvHPGhG379BVX62ZdHx5ISM1Q
MypfemGcNyN0gXFqtUq9d9pQn5rCxQWWXTlprd4JbHynMXJVormj6ef8KtBJHlKF
fJW0YF4+b6U9Y4BDGssVoT6jMruHUyx0M5ccSvFyQygdtHYbReUW3vrSuqMNMwie
cPZEJO+XeopzrIKpI39C83pxwLsAi2Z5Bn3Fna2exkQRRY/D4g73Kuate8qDdVrt
j1rZEVYh5OYoSvdPmAQPPizolCy1XF1fFDDI/017cgxZRgyt7hrCus7fRDRTKLxG
G+yOXJQYVndnuAFJJ/TSEkEMKIuSjzRhMyKC8rB9hPup0bAq/FWQ3HnRmrLX2UB6
XfhBz494mgxgndiN24/HTX4lXqY00hsyGRR0XSmiVkJDKNSSeP1E88w99ER2CaMH
8ycUI2Qbt9zLg5hKumDDwGmK1arUoK17Nm+ha5t06Cr0RoBD5bsyeBmzf1p3Ap/B
NC6OVLD1zNC+Eu6wrfELkkxYTmOW7h59bk8cWuPzrM1g9dMh+/OK61juafE7Ja/w
jqIdf0bZkaM4q7thBCTOGrpjnYmr35bElv9e2oWF+SKK00wqN4So5uVst9y49ikM
YmFoToLXqNqKxBfbK8Xtl6gt+0Neqsz7AtWlXO0ijQOc2yckxIDAoDxwF8o6ZAnu
DJPJW9E/LrSXMndMVC3TqRjp0MbJl4dR8EebrMRa7WRk0CaSmtmjCeaJe6FH1oBH
TCV0HrI4XmXPUiLTsDwLvSQOEWmTcn0XcnYcRNvZeL/QWSwWLmwxFvYurQQ5IOLo
zR3Og3eNri69hoyc3goB2QyYgkpbfEMyGfqJoajRRcw2dv/i9dE6AIUt2Zw4cOeN
uovOnRq+lsc0U9hzMgEWNPbtYLMJqh2DWuaBgs3rVu85v40fAUugBbgBDkNPD2sr
JEr7D0SyJsSBaRsWDGPGfE0sKI7gNAaat+MxNN/tKHAncFpDUZkKn8SIiXcV9Qef
MLJ0DIRO0STIz6FqbIo2fW54SzjCjuNJ98mK2F7h0BkLYNgLnCGZ+m4rG1fhejm8
KOTfOvPYGEKDGIrHDKI09DBQ0Q7LFmw5+XyBw/UDMrXAUAC8MaXZxttLy/5ce0Gw
wpgmVdj72pmSLLqfpaQqTeSiBI33I4gVaby7gTyVNI6/J08tjFDfmhARuOGzBTIy
M/hUi64uMDJhJauFbvxIep3Brvz2lCa3RFhV7Ai8OpIjggsWju5DfOz8BFznhK1W
iR5AsOV1iobWfTLkvL05SXsGJqDVgJ1kqEJZ/qG/PgdYflQjtq6QkbUFAbcVjuiv
amo5OcwoUVG6yPVJBMZZWelQb7GQOtlcqTroARVfgZrviQr7aQTVnHXY8XJe4eAi
8V4togzFsjoOYIurctTQnMKTr7hddlD/l5tocQ2+BedbBGnO32YIJUcGw0/FMQKI
Ulk/yHp8vlDCMiDdNHurNN/5wni2RzuH35NQe7IV12W4LRFbxjRKAdQg3qnpl/jR
RgckAjZqSaFohbkzK4CoC5NjFzk9uAJEojgtNjEy2cawI6/tDmZj805umLTxm61Z
vNBN4ALO5eQl7yrMcA0xYoGMlPeUvrAutwJuVbVjRukNScUf3ajzoQ6XMra8OXYO
y2f87WakEwldtHDvCBJO0p3UPfKnWxgbncyA6iaQM1xa1glQjQ8GyAf7urpv8dTI
R/+k43uFOI6SB+RI1C9SUWnIV8fDC8uKeXvZte6eHvNqvekIVOh0KK0CJjLLw42l
TaOGoikiKGT2W6MzQpPMPIp6l3cP3y2ko+v+kwZZOlNgBaixUmeAIY40Scqtjnq8
AzpvKLcAcJunmGDhh42jrVIxje6yv7eAKHfuDRCkBtlAEq0UOMjQcvL/KKR80/iQ
OgylBaZkyVPswTqc/G54+AwJI1CVM+aFzZ3wn+T2azOu6b2e3zFx3b6k+dJb2Rvg
ypYpudTmoACDJ+pdlQVhoRkKWM5qEleRKBRAnIKqTmdhhffi+OYoDZuAlaRv6900
ebjlChOGHGKk2IF4ukupl6jYfFyXabovM2I/LFxvsEjkxF2thFvNxbj8XWLgyB9X
bLyjB9/Nxie+rulLlb2th0obzrlhXHf0vJi0Q4G33oSbmjWHevf6+JcxUvmsIePN
urS0TzgfMkmnXSbBXIVoMHFH8/48J6DARSC3NKZd8RH/AENQGeji/Y4gyxnVfHdx
I2FZ/4a6xubgjRCJAdvIbhltGyExzGi+bhhCMMmsjePGbHuEd+HbJup0eChShQsm
gRS7GC6grC8KnyzhJQe7UiVP2ZLmQvo561KdtiVDNi3wXTekB9sMI+drzSW836LO
KqCgHsr5hCdTYICzJ9csOv3LTH/0+ybL/qCpDXu8dqEn8MZFC3N313uOcxv1verY
jfInytoL1n//8Af7lBOGIAvE7PQGEglBuTauko5yTDnwyQ3+dDJHsSvByLVPHA+3
yC9HOmcTSgZ3BevLjBEi+o2clSEGrgiSr6+Y2V42/FaQQeBT+gFHPmwfuB79TDJN
8xGULSjghbF0Hkyd3kj7naQ2jW+0Sq9RMUY6woNeJpnxuQHEg1e+qX2FCDZzyUH5
925Ik1Kn3dk8+zQV+xN5RBDt7oC7iuRM0UFqRuNXKWrDLCa+yCH5W3U94lqVinq6
DqUWhPPLpAt7nm7UhFTkCCFf4fDLyDWVmI9C9e45oaR4mIeKOLo8uwaUDXfed/n5
4EBJeAsaMZYQ5G61X6TxXELdn3hgHSxaisdGOyViXyAcpmjPlZZa40ZJRJKbL/gr
PIRZh90oVzZP9Rojxt+p1FppXC37hlGgJlqhxGtrUi19BTA2ARSfVZ/o0oNPeAfh
kkhdW1YPFZJ0qiXNEWoaKYcWBWOpx4LqpP3VYAwkE7koQ1OUlL/cTxjEF2IIj0MD
UgDJ0hsYq6Ah527OE76SVIVEZUlrtnZrvDK3a1dH0+mbsqAbsf6ydNwzXcQ+h25H
CpgnUe8k5VmivcpJm3DySYWb6q/t3kTNkLvFOxJdORjw/AXsjr/w0HrIDeZD0LU8
dY3fUJHC2uaUMEzCYPs+1bd4si5Bbdw+OneTYnG5npg3KUnDNmamSjRsyl8vwKW4
1yb0mgE6vhaViivIUjrV9Fiovd+cBHDrfz17jxLBRkFkTqUbgLsKkh4zURfdbawx
5mkLDcmM4z3OZYKltZG+3qr9HFjptSxTQS7O4bvvInht9JXrSFJK9HGUp2DohsJ6
43Xh//I/18m+8XVKWumhUwarOr76ReyWADHlPYEVzkL0D5RqrQVzNBdD+bX3KyiM
Cs26tttLpWhVAQphxXekK+YxvEI+l8+qSG7i3HF16QRZ/HJynPBhGAIdxWcBc2eU
IKUS/UM0DKDLaT9p7jgxEGQFabZ9KBqqL7LFbhDWOuNKLtnCcu4TD/ibT/LOrPUV
0s2c0ZDfRylu4uHjIAx1TLnuU2CTVEIuRUvG4AB+1vJyr0gLJ0sTAhTK7ONRvvBe
UB5oLw9ij04t0MX3C2iQorCCRp+9NQYcv8On1qZ8DlyN5fHpuD+5Yw6i7/zkr3CH
HsFREEDoxzMTJ8fhLUYt6HGOQs6zvwRYbZPqyQ4ausMJ7hhyfcZkPnj4qXyKcZqz
1Eoo3oFHO7MZTKFJL4fHaxitDpBeIpTCz4VB6k7gNrj2zcG2UGbuXkHmCjRJWgCV
S3GmFBdzrM9yI3tDgrA2GNMMxeg7gZ2utyhKDfKIsOWqQJkiQ05Fs5wuAunep5iX
g112Z4ZzmjwE+xjcEQACfFjJZwS0PZLyFuENGeqRwlV6bUBX9RhVLu1JtHI99pFP
PHnGy1vIDabPxfcCaiKuCoyN4Nv4IA1dcD5JuJTC2Pdp2hXBklux8eGwM/MOPNa8
jVETbo9RQXjwENXdR3/7GrvFyGdV2/V7GhrNY5JKEi8bBoSS6J4bx1xh1y6M2wGq
Mczx8XHBCiNS/yfpvpKh8YGqyxhOkfiDvFfgz1MjdY0B4HdLrScHNVOo9NbwTtPX
2GLr/BA1FQaWk8e9LzKP7ITU9Xvj/heksxGu+Rw8EvOtRxQ7UG74NxYByElUWxie
2YGAmrN66+kNfrh5TIQ7r2zLUnV9LUMX5/QMwsX2mVGtsO+SBppYOL6vUy+UaLR7
8d1wqUYJsnM/yWZgrlMUQh5UOUiZ+72bx3eE5B7DG7Wd7d9mpM1gN34GZSzhV19r
0LNWNb4zWBFUWI4G0Fljv6KO9Y31S0Nb0NHeripZQ0Mj7ihTJ/m5ht9tG5qieBi7
sIMZMbDmx0qRnbQ7+64GSvcKpkr0N5mRAHfUpJ0AttK8LyS8Yk630K6GxrkOZxZT
X2JBgmtF/Ene7LwpZP9D5kFuDi9wOKjHTtVMew27jaBJx1lszqqEfapG0ZQacv01
z4hRM6o54c9JgVl6r9SiVi8DOxmjjc1EpvPedsX3nYVS+geygbyvahgVsdj/sVJG
rzIVh3SzwwK6tPdbBXXlo9M/zQD/d3AihEFhRJf1MxDW6ElqaUi4kqr+A6ZiF0iO
PAEpde7PSSS7rHlRszNgtY9pjzCYEYy55/jqauWs5CMIVDDyhViPNCwhYM/TWkxl
RQJoty47dMcmXH6MbELaizOpcoDkU6bg1ajykuSImtdNOIvUuCT+L+PLUME75PPw
wRKY0D+pQi+VLI/Sv96LKSrqP9ibJzC9EHLz4GhLjLyD37fD/w9szielwGIpeFXg
BQBq4ycAuIupSxGkhmk09gaJ46FJsIiw12Wlz4WspTj9FI0JW7vLNe3bNi8v9jZq
NUmc7hl+gTyx2MFJ5PnByWdwUW/KetqEcYDklkHZbWn4vw1ebr8ZRi+JAdjlUM8b
MDLggzX3vUd3IlKvUxA8AsRt4Fjsn6Vb2gW+R+og/JoJBsJggtT0hbPcmNuvDJta
/4UbnIYCA7o8sQU+qrkmPg2VAuM5vsXHvqFLthUsj2BTh83VB3nlvnbLIJktickQ
DfyhbDsV1yRdzsrFKSwJAtUGD4Zgit8UipH5gcKWWh95a5/mSuGWo6MM+79t3QFa
evt4FSikFF8pJ7jNhzn62iZV0GZLQ2sOiUf5WZOv5/vchfIKnHk0cGSP1Ku+lfAb
sLHyXDVn7sEXiASPxyP7OvOHBDP6uWi5spu0CbLM20avrt79kUpFQLev6lWkk5UC
B4xLlDYl5Gk2L4QHMQvRX/c6DS20YchXArPKyj2mq8pj+1UvJ4DgZd3nTf9YV77b
fa6gAolNKva2gjN/zBC7vc8NehDbRPd284vmZgckIMlh5sB9RbrIBiochlgK4X6q
7naYey8kXhH9D0Lvg0D5H62PFD/U+JFYHYw9Cda9wzqm0sXZPP/HM1xWsUs1wv5W
YN7KlFvOIZglUjfRtDLNuDltrcr+zFgJGE4fuhkS2FgXISh8B7pL2brSDs+UXbIk
cHS6FL4kwMG5IJfiLuX/5boo5y9JHuLVANmVLcfKGbKW23o6e7148yjjZLOq6fFE
nklwcZDUXRpFC4mpbfy6r6RMXcY1b3RVM8JUhXfOjeWtasIz+w9KXNPgDMcsxW8T
n//R0t0oKKVXh5NyOvB+49x4Shi4M0JM0WA4x8SnX9lPia2zPFbfczqOH7StmRHy
kmseszNORHrD4Z9WnQ7M/yhSi/PqXh+8jdvhvTU5Vv+N+ZL99F7M6+NWcwAfd6MX
ZQuI+zJPP+HERL21PhVgapvHNLSSWEhrWH7725fPjGrAjYRC6BqnYaqy4BfHIJUT
IeCnWzPHKv7NYf5Ko9x+cT0rZWQCBiUNt3RPVWyTU/Q+NxMKfHl9rOAnI7oQdiqd
rp1opjD0wjCiDZFWXoV9JkK6lqLHoBgrfEC6i97v/LPBKKtv3mkNRaHajBfqIUDd
IiGnK7KZEDaZlhc3ji5L79B2nUN6mVlPPMXsIzKnkQ+bZt/qwGn/HOWdR3aGFkLT
KTwGBtcMWaHBQbGLYZP3vdZQQzbdLCbTa9Ao4DuuTiyhJ7h5TxfFupcvN73fDF8/
CPN6lFIRgHkVxzTYZ53nz6AXTCdDgrQyHmhsNTy4yqLL/cuCe3PP+TYUyln9zFXJ
cfS2fDQLRkdP12OHMyi2yZ9AaSUVZrK3HuTTLMDTZojBTdMgmo7ISb1iaU1uVRM0
+HM/Q40hB5AlNFl8MyNC7NMVGPOrUDrfhYGtb7wM1TahZYuUOYOqIQvTWcqNVDPS
STpNqBxUEbgstjdK/9qMlTaQgWPbEYYUdvbEoEZrBPzRVcDRazdOHOBIPgkxiK9U
78B3Eb0b/N8KJwwjeXF8NEfZ0I1QeHC3YGqtjRAfainXq+OLUA8Ht/mRgcYkoY49
tBVKcb+29s7LXvvWB5i0ewGAJzX7sly1RcMdAZWb2qf+H/IdlOcMHERO3735XwcM
RluxVpTZGEuow7bgkDxD1tYLGQrc+qSuGVuFy/HKSj/hd7+oPzz9OM+kKe6gq9Vv
ChiOgPHT7unoO1SHS0E4gAzmTXqM1kPix3D9dScZcOkIucQ7UQ48fWBspFsk5yZf
b66CnYu/K04g0auP3QdWg0T+rZJxp0ol5GL/Ft6lRt2nV2PuI5Y6FjYfCP9KD6Pl
gnb2v8DOM7zYiT22uVikixe7ItpLiQplANnXn9B//rcbm0t5R1K4MFkGLEefPl8j
EFdfdIgUNhmn8OW3qVifHKaIImKURhJSqcUVLDe95qBWndxA/GtBDz3DzpEDCVDA
tFsIhdtYDnJXrYu0lHasuKy7HMH7uQQpJt9/7L7DuShazCEuVLSKvqECUuu1KIp+
C6FlKOB1LB3duoIXzFWlCOyQGVHgbMyhZszOwWds4kQTnDRfh8OFOBEHEEpym1io
ocfm44oTLZoVHm+yjfcJiZBXQP4FWiCQwue9oKG5atgIO5/UYIrADwchg3/hCmKi
44s3cRMtVpQCtznIPfPZIq+MglolftPXR4barhn2tldxMtGSMpl/voia/AeNsjBI
6z/1w+I/YHGGCA7rWEYEkKutUwkTXymuLPbpZ89AeX3eVG2LagYmAhsf4CuJW7Wj
D9LWfGgpDDs5eXoMEUyGs24YZrYHRudb2VU72e00GcU7UBrzR4z1dxdGipI8ZPUd
8nPb4zwKiHih6cN7aSZpc4ElhkXtI4yb2RpXNvFXydBFdQ4OrPIOVcULxISTlGH4
4qvW/wisseGZnVxCsZz9amHhBPeLPAdLuGloLyApEJbX1asokCispjCoGu/+BcAe
hPl77s5/CnELj02wqoe2kR5GZvKuf7HRdWzFDSVp40xhbryab7N7I4WFYjE47XPs
j83vjHCVpv9eMqE8NO7U3mZ+2HJWzXosihpNtuXl/IbBApf7gEXuvoUwsm8s215Y
uYrqK6dXYj7lsvy6HhqXpyHNp9hwtQeqS0Cuxnd1IzGkooyfjo+HVR5s2BsW4Ne5
bYmbuBAy4LeJC+cy6EqfnEf3KERj16j0xR2XmZiqTlyDBEBTjWFoDynpmX3pEdgk
oBuPvy+xJCqtPkTH1cH1kM/1RKd7RQ2wzzdCXjjxOtHxltd3mDp3xY3Md4Cz//r9
9naIA2g+aGps0QTDAb/uuFwy3lWSLWGG6oMP1IOfOJuefrAdZBaKm0ooDPFnK0Wt
ReUzIZbN1JmZuK2qGxgtBSDHU/HtiUd8uEQS0WZalXgIT3pXctvo8srYgTNtSWa9
M/h9qFlWJy23MycNZNHu7UIpQY0h5hOqb70MMex45YNQVsTtGdh5/nuMYPBcMEOu
w10C69Jy4xL8uv9LsnedNbftE5DhUgWuQf0ITUnDxF04Cv9kcNSC1sie2pl/tBzA
Nm3qSNw9XE5BFC5+EZEkbh/FY+vGaG9DfeiVsIP5Fb62rpEMd1i1c9c2EJ7xDuki
TC7s56I4MSgSpJ5IkKz9ZqoltSnTwoMv16qZ/2aDA+0E3qToCkIfc+ZpwfFs3SXY
C903qA6y/1PtuM697aSTUqFB7cQR8aSzSP/S9DJZ6oTNl8Qs+wtmqVS+5/O8TAJk
CHvQVi2un7frznt6r6xRJPXsrjRJMuWD6XP63Ux3QoRqJDyOMoVUdp22y8X3nmQ0
Vqc0sKs84dtSr539lByZEi4/3hpXWRLHAderfSyLD/N+gHKmJYzAKzM+d4MgSXfn
Z3lpOZ6oPbWTh/OkliMiGMXxqw8rEJO5exxIECGUiI6MLuAujowj/H5tQPM2bDAm
6Ar0VvmrUZJCELj5S4tExg9AgglZJMh99xzqzlFRF1UWRjTVLWDimU8zevL1Jlpk
0hD1yCY37F4fCSDAmsgWcaiGxMVFiLdFM3XgA3JfzObKHY1LJOa3cZHGyfbgC1D0
h8pq0t++Cgv2/SQNgvddxGsxGD47XWfc77tZm5Xqx0ocFWBKRMPxoGktTDez14o8
Bs2It8MAPv0Y6vxImY1tdIUDKUC/Fq22PzNXGvq3OB9tDbhL9U8qSIUWZtLWtuOh
oSu2y0WqEq8+pYG/pzrhUpP4JelGSpeut+1cW9cs3Gzd3R26h7F0CDdAVQv8YjVQ
DHdrj5pKjqVYTQnVQhG9UjiARnQUhe8pUIteUEnPGrH3YY9MhqhcVohdPBk1n2Va
63qTzTWwKI2+zx1p5kPn4tAFob/yiW6wiEqcYY+1c7okJ7zIJ67duHyyBfnjZSby
1XNiAcGWuM37tA7T2krLii+IgjhHB7dgirRU5oR/uaos0JVFEsa7tTedrmCRCTgl
pbXNkmUrTulRPhDjpNfzSle8eEN2sgVYsGF0Xd7SVJEOL/UeU8rkbGjMbesO9jPo
B5KCsaOH1oBF69Bjy3a/KZOE4mLKPfovgTrjdVyic/47LlteydoBCBwmuBByc8VJ
f46eg17dtEQXFmU4HDRGfSndRsnFCV1QUw/CNdgiKuzMHNqr3+sfV01vbOArUcqq
AbbqX+qp9V3WKTkFcnFaKjjmpYJ1Qf3Ti5QhFd3Jc9IUQLZP6jvAmhrFbQUqMAqA
TeKgYohqfpMoR9LPGD5ZTSJKPOZBA6qlZ8IXNH3i+I2UNQ6WL17SujodbvVPaT5D
B88fiNax+NNaOabgeugJj1+sVcIngqQpL9UVm3PW65Qn54zfePTOM3SQyKonK7b3
4F1Ryu3b2ziKNp9Pc65wXAfsze17o1dM0COGpcDfHU21r+ni+KOVORctp+n9WQvD
/J1uPzDkqXNayQ+yMUdjebhWZwxbK69zHHbbJykZjcfBeBayYhEFZSaukhZC5vOq
bVcNY9GkePxrEQJjyW+1CY1H/U6VymujS+RAxKJkyf/MQiwnvB8bIcLIi37lvsKh
Rn+PCZ7Nvab7a5lMijbJVjkYPOkRQxuYSeezVVYp0OM6NTr5GXTLL10aPvZrspre
GExbs816r3CfRXFUZF5XHcJ11rY6Ho+9SCpxF8bLv0c1kPKxaHj54KuC49doNa/t
vcIABbJa1Z3LE1c5WFPuzhiTRZJ6Xtbtkx20hoFO9ietcTUd6lGnxotXfuOlylSj
LuSEOGg4Xev8id8kozf6gfHV16jiXQpzB1z6q5hozw9HSQbYxCXIZ+K509rKHyYf
P0S9NSAhN26c9gLBKWAfFETDEIJtb5mHoxD+TfkRiTznvyaSxwRK0A+ZoqKon0oJ
Gb4FKATHWA+036txyOh5YzonTuMNAji7n1LKjtPXym5LuzZ1a1b01AhXdnkAILlX
wGvmPBLDsRqqirtQuq2ClZt0q7QuIBU8mrQ2/IFgu08G3KZxE0PAroDGCNOZ+Bdr
j/LjNDGbtqceImbTjxp8sVvATSKZ3l2j/mbSiei04t1ng4VXI+SSBcTKmPJmZAGQ
Q4pz3hnYRdze6kEb45moGAwGhgjdEFRtjxZB6FpZe9ENmNE+lGWxLpC5wQWUYfx1
NixI9H6oH+UN6AtU1WUkjojyafzWDUY6tPGGy0D9v56RUN5bw5k9mNyPJnYimyC+
xbEH17eKmCJlzrDUpu25xhpTdta7bmwMEEXLK5VCxL2G17yXweVuydIUkCjVFKCR
SHPZmeHZCMMf02Ae6dzGkcxkHOpjI5dFgKhmewibZHFTxd9g+QILBcgHLbf1CCjO
0VBK77L9PzXgvya9oz/NIE7qVrUcsSc5uvldqHV0YLhsYBdU8guwOr6KPOx403ZD
T7DS+H3WiKTrjz2tmT0eoAYeHyrmzlTnDXwztiv+otk57mFayKeHMN32nAqSVEHG
R53vhpUfa9VWnyBA2332FFJ8zcPaIGPUsNF1obhajTbGjWLYzhDd4O4ABMXueaMf
RbZfqhN/K0097Yjv+pZ1hXPIeA9ekMMi5hxT0657XSIGwRX79Nr8VUoyBp5Otjc9
i8qCdrjsnIeooy+oydRfQvbls++PgkZ6ipRU0z9EW55a4WGYKq8lg1kh0tpZDYSB
gFI9ArgL4hOji/JmAUD2u3qJGekIvFwpSAwI0ormpswUYJTNWS4MUkd8dK/CwH/q
hiBz4vtgCH46sQYIFMMBfYQOfuD1dieNoBIBoms+UzQnF1BX8yfhOpScJ2BNjTjP
egC/yWnt6Q+Jv2HBcS+Km/PghbF72vVYEvy0lXNPnfLcM6Vjr9IOmmEFMPXju67V
48E6JmpOLvJMyMksnKBy1ZlwuaA/bc3fiJF4o/qDQPR4lyFNdWLLtPZ1M0Y/FYw8
XxT1DqWtj5FI45ycykIb1OBVojztBG9IqWDi33rZRghvq+9MW+u5b6snBnICqdSl
B5z/XWbuntHNBkE0sLNCdQ9xKGh9uVIPPUxMOwrHtbYUyawunWAqIhErUCTvZKSq
lwG1RIdNOF+mpF4X6k84uweBNCR6M7rqCf6QrD1Ew1WjpotYrQYUABQg2gkkTKOc
E1mvfP0KfzmNdFbJJ2VtnNX8HNZFqw1S9iJuxkpuUG8JvEuSg6lk236GjvLDqLHY
MwJYWzSe6IauIBfzVCP8jevMxpRWp8BTpq7rvRHW/4gKeSDQ4hHFDsM8qoh4dmZ9
ACGS/2PS4I738Nmd20fG7RZFkBwEFf8jm3arF0RM5U3sQq8AjlRVB2y2UI7H08/T
oi72tzM4E93gIfsnxPKdcWsRpkyo6tIHm5GgykEQC6duVhqhTEIgJRLPh7rsIysb
dnF/HESHLyvN5sKbhnlhCWoOCA/q/fHNftera9JV3CRGH8zPz7GmC0jsKURZy0DX
N7+TwooHFZCvfCoeRchCRkAdEBYISBvv5noloMtNW9kHsHWR7vmxOyauvClS/5P/
cUjY9UM0CZArxV8woYD1DtJhZqQX6ONCRQXbEquOZZjx9QDKDi3bhsAyUV9T22dO
fZpHYVSB5lgL4gWxvGMm66fXgf/PUcRVdDmRLrr9e08YFvRx1RHGjtosZP2GG5go
wnIoYTOWt06LbEf3hVDE5fzYfjLYk04YxE6h2QF560TziaHdRXA4MS5Qs5snta+b
SBuZXywtTPNvBqCFFvG5R7QM5qqG7FEubfoVVtUGGJXM19jd3k9xKA3WELcXVMBS
6lG3vJIV1E8QL3OGfgqtOViphaa8NaoPuih88ZtoDHdAjaywJ20/jshdlhekXVxR
k9eE9iYefoJpoXqQWCpfHsqdj23XzDuIUJMZnRXQHfWV/lEz7HRlnfAwcOntHFHV
BVK5zdgpfeJxKyk9GKP3ceogEBmgH055N7sB6qO4Xi7J/0IiRj6w/5tP9flKArZ+
nH+/UoE3aHMTcAS+p2QNFdqnWCkOcmHh9WlQLzcgksBEu0kuyRrv+ti8O2ODAicn
2GB/bPRh8D5Nk+YlsgOlGsIZCWUznt9I3F027ms0SH0r1zptdNCx0fC2AEoPzlZq
NAXO4e05fgy1TIzosPGkDx/WPpADDiS65VOxjDScBnwBZQXLckoWTAnPeRMgOAXn
G7XspJ+LQ9iqbFlO3RJO6037sjzLIkvnYKqqjx7qcXOSJBv3jGfqGDS72JsMDLxG
o0LBBu8MKGDOImzae0jo9VMHddoIuTlklx0qEawTJ0oWobICdCU1rAj5GM7O4FOF
8jEkjQwJFng8otcpWwE9CboRMhA2rlom7ehGSvUVpO5FZE80eWOKuKTAsqwrthbc
JnYQ84eT9+xQwcj83kGRC+SEXHrvXa+BiwvvyB4gnAg0yQCDoxtOVzd7zJsq2Duw
gyUstIQlfstc+8vQA5AAoHWizlHoHvvyc2iLdbl7ZAmK63amnY5g+VWaOi3INpNa
6SJTFrX+tb+KlAUlvPS9JFG5+opb9Svlr1dviuA5yUWNIeFxLAPr/+RA73sw2eIL
BDEL5l9+iemWbtrWuA7fLopyrMZZ1+pJKn4zuObo53nrWs3nuZioqzyiLo+UkO7T
ZVsFU6KsiMmK0uvYvBGY4xl/n8umOygCxIfn22vmUDANs4uss4Pw2IMAq9YIXnxV
eoEUtC1d6j5WzriEcIZYLscS9yUz+GhH/dIKD1mpGDluWhixtDVhYrZ8sBiTCnV9
RsEjIl4Y0XFVSxwS6vcHsT3sER2wF24N666mjDEQ2o9HQlixZfulMncJq5J5xjr9
l6fy/dZP0OSEFeUkQXfx4gQ31wuB00qtituRxAOr3Z6vjKPYOJOU8X4BGlKOdEVG
x+FWpixVt/QyzjXk2KfI8XCob/Dv9Iu7FTdNtvkW6ume3C7Bqc7AMB6043GvZTRv
5yHHUJIRUsHtZmGHwVsR5LQHxHL7weDVQpz1Q94OrYlJ7OCleAYpVpXYO3lCZFNl
r709K5jsJYMafEhOz6qf/rwlUNu5ukRMpvljisELGsp8qIe/OiSrre9SQmyS97hs
axoN3VULIiCPMXKx31Y67b/Sz3p1XcnK9Zhu00E3v92Kb/17L256qFK+M+lie+KF
7i8TsjzdL+zF+OoIQmIwSt0r8USqXGPd74YAXQp8ANY0mUt/zwXUoJcx9VIx6o8q
MyIvKR7M5FnQp0QC2CTiHoieJWQwKzH1Wehql/9J9uekvuvt30/pipvgdqvIS3+8
JqFc2yWKyOOuzPBrpvG7dMZwiVSa73TiCvkWzQr7V5yHfyH/AG6UhJ1n5fKjHarU
pk6DtJ+uGLIzIsAgzUWIo9l7iO3eNjcIBrXE+QMwdjfe7kdkDsa/ni9R2+sDMSSJ
mYvQsmEBMyoB/JCT6jmv6oTE674i557FUJCWJeephFcbXL/cNlSTtM4n+Rf4Tjpr
EVd4H+I6prg5mso9+WUqyw4Ny0xIdyyQRDErJiMh7yKU3nKGQhyIUYZbZKVPsvsE
XTpGR605srmTa+Kep19z4vRnaRUc/JTwObk1LWcr8Kuzd14CzdDdE8rXcx9xxjzZ
spmgVorHnxmWcs+bZcXKJNb/cbnUVdG+CRACZHSWiNd8rpnZ8mMakB87Fi7q6HLP
5vXvnKheEftL8UrLVvYOofoLYz3Y+z6Adw24HIr909CfnSB+PSqq8cxlp7ZjwKzg
2hTVM9nmjGZcPE3lslFgFjjtw4V/bPzXV2C9mgjnjcdhUCYHCv6MBZCOqMmY33yp
xMACz5LtsOnQx/Ti6vYy82FvWN410iJr0+5WJKB+K9V5l3LUxJdR2HBD7fWmobIv
2PU4X8ZPa520NkRUZu3DYHaianJoV2sV8f0Lng20LhB54rozfj20suQPmnoEDt/2
X7xfxO1DvN4P/Vb6MXqyQ8zcCYEB9ag1qk8JgzSvoqbvItZMkcAay01oOSJyn14L
VoBxVE8PurDTdDEg9ptr9ezqpnt1ZLansGpvYmYjkc3lfZqy9xCvtrysM87p9Amw
U83pzaxCyPYKDY/jKj7C90gWb6lrPBFbV8ggglNZvirKtay36h3oV5nao9h3S3tF
q6cBV/fAeFQc14v7xU39G4LkXteRRfA9MFwvNlddGT4h0B46iOonrvF4LBvCTTeW
/6OmQktHJDb67iRJVG0V06ihwyIqGkR/mOkM/XYQ5tb4WXWk7odGXY23GiWZreCv
9GLtWyJsnQf20BwBxYwemhkQaX3FPOdns3EQdxhdmnM7AvI1o1U6ioRx75lNbIyW
zmF0L22h7H8WhWfO3KLluVLDSDHBkj7NTuN4HLkFmlIXgyzVH8l6xBHTLeKvSy00
PR3rkUwmFvEgZVHEy9thbNZC/sZPxrYzN+dRIhw1r+k4KWD/asaDgzNPANCIqgNf
fRKOpCFXjYxwntZE1fOKEReDM0I5qRn506lfU3HhsxfUpYodChFjKHAziBSDoiwF
M6NePJVgI0ufAJH+gQMKrFGcCC+XFpKepvPluUL82g2JiOv13IXWxW+PiRD+3Wqs
FlkiwqG6WTN+/DvRk7m069IRz/tt2BIW07cPOWKhg7zOeCSvkTtq0WDt53+KIKCt
1pBJFfF7T36/DEBjMJ8PaWH6I4Y2MXPnaw1XEYq7491Mg9NpVmkakjj72IzkX28V
yx9bVGo69o4RQZFmbP5/pA4cshBByieHyMe3zXmpLqb1D97XFzk7z/6rcokT34CT
9W7HAdArTibAeBdyF8SDa0Txdj3Qq2RYz17/lFccqW9VLNFReb4E8DwAhnM4Nizs
fQdvlhTJPJpN45idlCuM4vxue0fOnMB09a/J4fz6Mi1ajsJ8MtqnjibrGNy+gWMX
41EfZCqA0bxkJqO2z/dnq6nsNQ2n2LJI1EB0nWEymi3CMooCRSYzX8ChB7EvsNsM
kSH2ZZtKwEMb55Ouc7p+cBuJnAksxGCig8SKsnI+e6/dB38ISgFZrO3sgzsvkGLl
hfT/xZIFUnJ16bpCpPL1p9oEwwzhRL6SCdTVeWqbWQG4Jpps2gB+XEQGERfIkBMr
F6aSI9Uk0EDjlGGXGfSQnVw/7arQEP/CHZhLiCSXijRySjPhGIapKs2Ad/5VAVsj
6qE/rHaHxbmmHprrzFBHVnlaDHaM97/bigDN93kNGqlRw+SArClgHJ/ZzIkiEx3N
4iKVwIUCJ+a13QsJpppEXmVP8DUqRHEHF6uxShmsXQmM/hLRrK8zcowxMQFnRewD
9bdFIZ09fcBbLDiphN0DdvZrm0X8cTEK3Lm1DQqVwoy9HJO/GB1OF+7Xz6UXz8Ie
I4euRQao11J3SuxAeSytwDnvxnoksFDHOVjU3DQRw8ZxIXRTkdWE7JrRCyo1OmZA
+MLrXkCpfL4P2RTLFth5/Qor3qUAjFr93YxpxwtmmCGL4rKipVMld58LnRiBEmkK
Us7OYaNkaPJfF3kQwpQyr9oPox5+qxVUnTieNy4OGH+QvkGkd4MWMJT86Pi7WdnG
cF7q2QuMnrXEqy0bxUCKoP6QCwfaczb36k3DFIfijbGw1bfxWiQvOp9uJIjV0RKG
9iys0liWdSFWeMn5nbhf9GSpdGIVzvO1iT34IeQZnHFtFTE1jXyIzmKvSPPux9UI
KDZr258rRg6ZXGSvi8Au0LC7T9xoBAQJPOO749LqkA2OUmo+hQP6v68oSFrpRwY1
ICCGCqN//Y0pEvth+0S3eLgomkMDfz4F9a9dpsassz3O7prI5kTj2xD9X22tVFk0
CIN01VBDVHqo1xDfdgdam9nlJr8mIkKCsrmRXvqJTjereIc8t3U5LRswDRsaTL2b
D9LBGNNZ5Z/dymbcflqwJpvQqiZG3KleF9Tc/EcYeDCPGepoqKlHvksQjccNGNNY
5lpgn872F8BX/PKR1FUp1t+N2ccEou6Bdq18EmqX92/mAnuWAlADYHltXj7lGEjJ
doEv5qKsX7Qx5CvUPmXZ9+N4Tvmjn//MfdgnTBNdejvTES5+SpMRxvSS2dCUNmBy
1awPF2IUcT7mAl0nvRP12dNNyyT2JlrW7MX1WoxbqqRo8W25mZ1onKeqiu0jZmZo
owxPzeW1cbtuywSKTYdoEo9l89mDgVSG6+WiQu3b2aoI9BVabP4gWRboLzkWOh0k
lKL8rdIWkQpT6+3Dk8diMnNOroQEyqCv50PwhGhCh5BHqrHGuoMAPOaWWxE0kt8h
JWOLYrYAPIgYNMq405kIqS9I/Il6vPRVy4kOAcjmL1P/KISE84JZQfXp5GkxoeCo
dy+05UwzKGzroGzspfT941z1ewtyClUEdPDUTNgwyb6Lxr1Rh5EwsxlyK/vNYZ2S
dGBPnbJ24R0DERPvQCkXVHu/p47TSHWNMgmOHZ41aO58FMmlnuY300DOLnkj+pzL
0OU7/gybJGDQ5j7GFEJDYCvPH57s1khvsNN2eLVne0SiueBHT18axJVTPWXHwdyG
Orwk58fY/h7Fw9gTHtoYNwCqGTD22Df6F3HKq0tnY8RYRWPcS3yIx49Y61mT0RvS
kyvfMlS4HHtK0HPZrXVGqaqJ7avBT1WaAidWFXXXo/x1cgU2lpjKZzxT/YRySuna
H16csreqNlyqXVl7ufgthWR4IGOy2goLuuqzaUxoAf1RolUaGKsQ/X2lmRt5Tzqw
A9WZL4Tm/o+iwIOilebya6cP516C/zmoG58wyNxdWny74qdiJUjJDiQVMHqbACQ5
RCqGigl7N/9jpwlOV32nxMCwra1WPq0NYpM+YQp8zIAon5eDSBk7ta+UzydaMrH+
+ILlpZjHj9fti6dpbenWcEd0txN/6E7CoKX823xCfZkv0iFY2BHtvjvnvUs0sh8g
Qr7duuCQKGXPnBUB0o7rbN4Ha/HJH93018Oqb2rdlzEbYRIzvsdOENL1/0ZULnlw
hZrJ5drtKvvCXrHcwz7mVGJBVL7LkPJc6eY87D1K8Hlo9VlGsFH5k16fPL/xRpUd
Nmia2H62SjlLl0YOy+IDaEYRnVtqTfnkDXmfCaNVYPsH29t8tNrSpOkwzeO+Y2BJ
BdwNF219AOPJks2Z4CkQbWJ7ZUsONMngziHOJBecq+yquWg0rCoGx6Vt864ciNpa
IegQwQnL5NfjfdfolXmZut+1LP382gmpMX0mlECcktis7i+30WUQDGC2xgO2y+Fb
/0PlJU4b6owRm+GDG3mFNiTqeMZCTmkZ8u9J6mvAxL/lK5bStK+tn9e1U40+rpU4
+0WfnlyBnPRhxleKrcrh+4+9dI3KSN/tdVzRzMhPECBr1fNYjJ37N2BFcZOabNGG
6w2F2V/CRCMhcBoL1kfq+UKBrVCFDwcfINOo89nKF0qtqF02GNSPUlol7qhJo/oa
b7M5n3dHU5tLW5TBqJBnVo3jR9BxgxpdXDhNl8cIOMFhhMCr3/smhU6p/XIMT9nu
CJ0ytcqkk7Hc4uTlYNtv8b3VmepQ/CdB0exFGJ6BMuvCYHpgYkN18v07T85RC6Xz
EnWpGluUH5uUsCB3fT/BgmzeSGRf4gS2flSXmuScvo5eco2mTtfYh1H4OxbGt1vh
aJazDjpNmdWKcsZ85wfJP++uDlqFTRtV+FR8cuyVDSpA7zd/dcpV8bPqVdgG74kX
a1HwyBge+Ob/fIllMlc9gnowtt6L+xVAWYm/UHN48QKDEpLr1F0crkP1LYD2CV65
YUe62o+6oUJE5LzUmaM65AsQz7LYxbIB1N7xNZAkz/BGKpWcOYXWsYDeopdjdj07
BXqFy4ZmNr5LSOw/ZUSW+5ao3lElVoxWbPwFz8TkwF62wAoTrZ4RTSIkGdtdXFF0
sXu77ulPYfrx89UdMy7cY50Zzbk9O7m6AF1ppib8WIUp1W2hGkBewnjYx8kkKK18
ef6SGCOCUwZ9Z12MItlMFfDU9MkIzVJyBKLLxEQGMRrwL3w81o3fuNmWEbc6uP7q
LsdAzFWg4MIy7d8THI8Qujd5ILFRvtEiFkHZLJFVMvvXz43mfPTfKedCiseKfZNg
u5t+h7x3dct3OMnzWMfnLWMaIVrzIdQO4laDBLhixbi1yfN3xvZCnCeWNU5Sblzi
i0A2OFJcLUFfk0VA0ZLJRSlBIO/6PZzjK1KrCZbUECBLvB0VS/1RH4ovE9YlPrpL
HXVeVMrcBB6GojxJ1HDSH6WhfcQ4fNYQzEsnWM7vv8o3wkkHN9Mnh825upKh783K
+n1UtaoPN8LvV3ZcjcYFzcAgnBBGrbd7Jy3VN6lJTPlA0pBtHHw2bi/81WuIdc+8
JquzttDCkeBUcitAT8wHLYuAbHcBofJvmsROJUG69kFqs1sJHdEbcEcXH6D5xZjj
nY9DIS82OTGCV8XukxEQ0WH+CaapzoPEf2n2uKWLTKwxHQitsiI0cgV6ugLoCUwc
DI0acjd0u0tlp9T8ZqDVgSCZNQ5kF/4JV1w9qsAh66ZIfI3OaUH2eXn/V19dGMTq
fd8RQq1QD4ehPa2juoKJTMrpyTRbQpkYBRXtQwOBFgpcmgnN/4S13TaXTiy9YVTD
vWuzoBDgAPk3QjHAENkrXp5+MbsYlE22uhlO1qey6UJ6afV6YcIKc5dRxJh0TW8S
HxmsfhT6lQo+H9RLsQcW0YbmcsMgovMfAQGv9ubsvY/t6e2yV37vLvQgykWSnqPm
JE96sA3uYjVhfo6JBV5+sovAKgp67th6j3VGU4Q0KQuDF12uZI+KH36Q7kRw3tVF
hTWtrn0Gtx8BmUAtJorEOmKOH97vm+/8otnaP8sQJr9MSHM+7QvCJXtkJrNMHMCl
0eQsZfXhmUe1NqVKAEdjw51cNlSjn44e+ldfIPEibtgIcyXnZNWtKqqBsZSXUaOw
+gWwZUu6lyBy70xvyOhBnzPDUBuj/MaI2XNnOXNKnNWENNl/vAV1wnEoW8xYRu39
gzy5cP7nVGOOuroS23svRWZoO1de8A/iSQIlnDiT1nEVO1gb5wDZ+jUOpAqBX1Pw
emreNjc+b9UJDz1i8//7x/4fkbE4hKEnZOetwsJcho62DFPZ4dkimTRgBhqtVgbA
ruaBkkdI68vW4zflu1N7vYkvTTYetQ3SKaazIfygmISZfqlM8TxVRHhANvXM0B4I
/SDa9ZPIjM38u9HzSqAjvkTyj3+sqO5LNmwOzRytL1ox3xvQbdLO+htdERzutIHL
OMRXEzOdpCWgmuDP+Jz5UeKPZ84zCAOIlHWxuEaMNMfMs6ox7P421gVBdCAIIerh
IMsDBFVz0v2qOcr3tV+ywYwaru8z+i30xPDbboY1MoL6LadCMMiQue3Pff4Ru5yU
QyEhOOMCEctSl4DfYjPByZd9zYvy//wbhWP8+N8F6MyUh/f2tTaae1OrDA26CNu9
vZ49LeupuV2q3dCdojfnPKf35RQatPpXM7eDXUpzyz8xoJLLJzCY8BG5C+q8dBBe
r/8Jwhdea3zeZ7R2hVF04U7CxUXGEno3C6aWFXjJpxF24jYiWfdSIwjfNwtgc8rC
CSKwaOpQL37WLFz2/d04r3LPyiuvBj/npGjoOI+1vRo8fmpNGXtNs/Oug/Yh1kcn
UcAPuQluN8vZubPIxr8eQUYK/6vsLeKM7clHKgFaYsQMFd+gQqAGI/QitMALM6tL
pVhcNfr8O0E9svcJYRPaK10pTMuv5aClk/ELLkw+7o5wWfGs1feKVXe83LA5pg91
/6TWY8kgeLcAP8kp6GyyQFTv5cspfQc0ZKrj6pEvvfdi//lHnTa9ug827E0Y0BFF
tj85S2go2ci2YqMSmoElWWeWtVJSVBbRbk/+ksca6P/cSnspcNEET5zyK5+a1Y+i
9Kpg2z7Jh+cvwbHYIL9eS3k94p2VH91LWL/RREcFqaMZDNZHyE+xaOLNf1LIydjV
i5foGcMh2jDhWoc0TV5gR7XlQ7+woKCZh35jx9NRNnivRdon+1uePDRBnMHOqWL9
hNg21bBiGSPRW7Y1tO9f2CAw5tp2P3CUBTic5QuKaEwg7uaCB9Mg+D7Z034Mnvl7
cUBeEx6yfv4rxAL83vIL7quqfKKDGeo2/blIygMU45Jpwt3+0ZzNHw9HdesU5w0u
nlR+JYMAyONZqlTckDsfHg3GQThASpYLw3TitRkYhMgixfIT7IzNh7oFYAVyTG9H
ddzVC8KfJVQAsFK2fk2OzMp9UyOyFZ9KYwaPaTaRuuXMohjHVrptKUTC7LNYDOuW
mV5ZNQJY4Pv+4NeLOCh+bzV/mgRIrUEvk2/9KN5fcV2IQ00sQztAk176iR0oF4J7
6pHpZ/DTgU6eZ71d1GmTePKYhIfgB53tPyu7PO0D+p+QdE4Nwetz16DcHltL5MaZ
JLuCtsSxrLgfthslN0j8kYy/L9A4DtQpIhGdl5+ZCAzxtFqCNdWoJf+T55gHwJgC
F6eF68QcKzqhiKOvRKWnYPOasW7hHE610LPNZ7qKUKwhEjInH92YuMiIJOkhkUms
TYWE3dLfHmMYhb186mgh1/hdff7301JmQAW9mwwr1G4Q2riXHaRuWcJNvzO3VOfJ
XyPSe7WhqA6L0//htV7Ih7eAZ2CPtKqVEtEDxD/mIk3GycI387Pv5Nzizn9dBCT6
t3l2Eb99tzVHZTuh5ujRZIcbNIYE/Er/nfRckw1qawmcDhdOP9ZFzlyWg4xjg5kv
kJyqTWV5R+wLiogbnOrtNU5ruFQNobx+qpYJ2SP1E9RIk5QWrxEJ8DwAbhXxXhQE
SGS8V2fuuldhy2DKSRyMTeUJ8VJrCsliZZVu6mbHId0lIkxZbpI003iCOO55Hz4X
gsp0bFL9CFWOrP4c0YA3dX1NHBPFkMmLt2/JwGuus3ucd0DQc2lBcpUv5syJmVgQ
HOoT/cVrzx9p6dGbn2d4PtlPe+9uoiQ5aShuPpjaVJj0Ouq4lTKPvudYc6ECKHnp
EOJw03VVtASjFlCmsdGobfDBVP7Tn+THFV8ihYK9G0NqircTF+j3YVwas8wke63O
2CJiwWAz5ZNBMb6akT78wPP2XS92umw/SyrywbKJ2++9z5dlsfK0XmfdkHiXzO/5
Q8tJno9O77S+Dyqcji73pX/26LTlpW77DtRwlRz+UwSwl+QZYwWmh2yweE2DXIz4
xTM10gjxEjdLsj2L6Dm1f9I84qCWphGVy0pts0P2vOHF1jpumEKNHvqVKwBKoyZl
1L1IRi16p0lHaeMPDGh6hJaHbKyqCkRZfFwCwWAhfx5x09tK3MojRKKo6272Z4pG
y8CrTZW6f8/nFAAriGIwY42GOPYCbN/lFPOcDdURX8fmfSrnj55UeLGRwOCuTskM
Da5uiM1il/ntZDeDo3rUT7XPrchP5ZDyO41P1KvhhyjLQqEYo/N2u+BnDXz0Rv/v
LcYGhTp/qt7lkO+Axfn2u7cgsFPPsBCdzndpNBHFJBq4xzxNpRgTnlchG0ZSmmhE
yNlh43tEDmV9LA+LyBSiDQunqLkZL8UeCxmEKHsWF339W5OLRHYCLFrDDRPiLC8+
MqT6+uLebnjrVHZUBdCdrsW85QLNg+YAivG2m7iQE4AAG+/7GPZLXPu+WMfqxl68
uXXrwCyNmzheW2RrmYu+s+ANCJlVgaI8mCbDE/yBEgurE+5PuNzETExVgqk1wZqy
8q2P7KwA3RjNmPbLOzgq8RvMKbjE3y5F7+3sj01maa8w2Bqusup/S2yleSWuAXQa
eFhMGsAJznt8QJk0+OTs5tPhfBEHCWylKeqzJ7gPoi62vzdr2x4BbkSnhDT5A0sj
L9vd8yXzEqnN31xUjxNWuC2PHAD5X1ISXNbilGPmsTpwL2Kr/cUUg+4nMXbxfYDr
onAqBQOcyJINZLfeI9nwy9i0o5Q9WPcDltL7W8rouwnNHUtDGaBfdyZhSXsTpdcL
1JS4ulDMdLwfaBXdhtg428Qv6jS6JQHrB6i+XV/Kz2Xed8EMrhcN+mpACfelMetl
Laip5zrQ5nk2XJKSlYdGGU5njlrgEPbH6im0/RyRy/mJbVBnO0kyWbhybxHeH9Mv
VnSZYUReV5qGHF+vhDGmESfd/UOnT40mBqNs35zYhCHjYSIh9IxZlLS63LThxT3c
B6tIpCnVeE8W2gcdDLzWM/6NXiI7YdWFd907Fx4Lvp9h6+YNq4f9kPeAmB1iD3QA
Snq5PEjaTY8h4eb/rVwDEhr6V20s5ppMxu5N69/iQBV2+efjKYchfPB76j+z8whL
Ln2lsHq2b17Q+tId6LTmxqY3XNCadJf+8LfIXsEmSoXrX0GdYun6vzxQ/7HHMy8E
4GC7yM3MKVh2Wmx+HsWD6P0YXtCg4s3FtFiyC+hlZEtLQEmXQgvtEsNjRjj3Poy7
rSFIeYtWcMcxApaoBvKx0vHigRUPqy08DcCC6DaSjfddyFBy9qPVbN8SXyqnIV6y
mIHR5FSZov/kpH9A5yVhYSe5ktDza+2dP2NooTQ8Wtz17u6PpJom7MSHkrgNxOol
498XcAG5P1BH/fS2CQBFuAUzuHaTDSCEN2c73yliB8qCa1b11/+ZCYGaeMesyVN1
EMGneHGcWfiku9zXITNB83MkgCItyGEA4lacrKGgKuPvYKkHOxRzZIkZ76Cniwv7
3bHlt+4Bw+xv1kxvONq8ailsmk0gRPcVdHoJSByQLZDHdeELiNFrm5oy+TDOEl4W
VZWL9mNm4nfYj0icIjRRLPeMYdKn/fYFgOU2saujE+sG1cNfChCgUoHwY3efukG8
bj3SR2mDmky7aanHVwstlQNM2G2VlAkx4N23zPa1yr+gd+9x0tIpyw5PG7lhsBo/
CEA3IuiRZiSWPSjhhbKrIwcxiY7FyhB9iFf6mTwcVsq7t6jfZ2TOLOxjEAQeNQe7
qEN8IF+kk2DnvFV4u67EHg0z8oF4n8hzyXFnZ3R5O5JkHEBByrlUF4xNhMPnaL68
IUFvCd6kC0+0Z/pshsgf4JlEIuOVDwJNJLOtniNq55A7kmmZhiobwcZCZk0eVLcA
LyfUfvQib7hL/BcGRMGAQgyMperjwJpJqgTUSBG79jcFMbkFUoDLqPRYxKwmldpu
woiEYCB4Iy/kgEVmkUQIntZWlUNNXnteR3UcVIhaMncmPlQxnKWsJPlvVBLfGbjO
h0OXPqSuvsaqYsO1CLQY9B64AlqX4Zwz9dC0aMDNsLJsKVuKRwg0UNcBwFvNu3SX
rLP20FWy5XWuOqKDFp68d83Naw+CJWy9f/qd+Jp3XNAYHBJDXf9YC1xvm8nhcHcs
BrXJADAM/hvtAcvx2lV+GxgSIueBkbQXGX5q1GK7VS2Ja8A5AnQ/ahlS0urFYrGj
0FvD8vPIJ5PXw7limqufvRWAl/wYpXFeMZ+WLZkhb2uj04cpR4wVc1EXkfBSwAge
qF0DnXOzjyUsGfDNM9/EPNNZ5C2sGSy+ySEl/SLs3CXa2NAQek+RnLeayP1i0Scq
FvLbN6W1lgA4IiTRYzCs/MX78a74EzWHApUX0XRrcZfm1isyderYqrutTCWH9dms
uBgPueNaNgt9+ZQkowiNRxCZzPyg6GnBv4YF90IA2xLWGrysvYXDHjySRh6ZytSm
XJ+fkMgAEjYYHno/G50FgXbyu4XkVAV0yGEYwgkktp+f0BRSKS1igCiLi9Rj7Mku
UpY3AhQl/gr6OsSOAfP8P5wKzDx9IfbF6YCq6v7j9HUu/21qoI5NHt5JKBydeuKP
7R/aE1JVSf2e2iC0GwPN6KZVsg813yBFENUi9v2JznZYybAmrALcPRaRV86bvzxV
nDjIEvMWbPq1v2QfD1DHew2ZUfnW5ftTTN3UJtR5hOWOq9tRUJnODnjzvX4vHHCy
TQKq2JxkT5J+PMh0rgbAHvbMAvAd2wlLvDVEInnIEaTteVtukdhrW0TsQeufwcf7
qxx0OQrBs7hqyajG6MHqUtpLWMtb3O3AFpZUIvIp5uQ9PrbL9j6W4ldZNPvI/lZx
E4VBfOlJXWLjWaWgwtZ1K6DQCSzk3/GMnv+S7Shhx+Bs5xlkkXvTWzzunepSqLV4
WCAEi9IOf3Uha1/3X/ZK017mBIYGO49irY0WxzUQdRgG0DuYl3Sz6R1V0/kaCN7m
XyWj3hWpUWaRhyugLCpmatmynR01yBOWdYHlrdJIYMsxyteNfkPD3zdp0SZmst8i
2z3Re+peSlek7vCcRdtgMoWu7U2j0mXfcX7wBKN6oiTTSlAVtTAGHUndZ0We2VAh
2ZP57iYfRC4aURBgTEFb1Rakqwoy9nypnAp9J+/2HP8K9IW2MqzKdhvGXK5FlHVx
WY48D5EdKNiV6jfnWw47NqX1aItPUJYaqWAvXKs/Lc5oW4qbeNkgt8cauAVz9WC1
TpvxJI9gIKzNxcbiQLl3hrJi48MAl3PJugspbftbmpB5RQj17DC+zck7BsxbQI/A
8JmzeqcqWN1lmiSJez/3VfgrbertAiVZZkcpj1HfVuqOFOXt3YwbhN4VC4o6kg6+
a6uBMc0qRcjGA0vDRuIc8oGTm9t5bMSxjkQHekiYJaXzq0gsqufnYpc07RzfEawQ
5+HYFDox/EJ7WWIOttE4foJeORN0TnKaT3ezwyeyIfaLVLmtqqEtLMxeJ9SbiGZC
QZPfVejPf/Vb+LNtO9eZCtjQDX4v2FiJnCwrK+StLZgaWot66e1tGh2JCfOVWfu7
5JLA00id8/jg8nHRyB8Wf77C69+MryOBOVzR/bNpGeZvH5q+0bsaENVUddJsw5oG
DRyKUFa7Mb+5aBOXP5xt4tuF19k8dLrOOl9zAZyTsxIJIpjlVdf19obsYWdOwawI
FV1tMgR19/JH1jjJHQK0UnQj8iI2PvFAbJcdOLbwPXCQYguk/s9IJ7lFz5dO6t0E
vhSxCpXNI/qY6wmBe1l9uKV34+abD/KXVjCDLenLkvk/86/aL4fxqvZnq198EmI5
oIuhLQ+VfDi9nG/ckWTNptilAKiwVakHyCki4qOsA/Dj62nyi533uZTalBFyhi26
IqUChmk3qWW5vCz7eFro3UvasfwR9yhHyyYZd3PrDtSO6IRY8C9DKEImg30GnqGg
Lok/VimFRxd9EQgxAjgqi8tMuxxTsLmJ6nwj23Se+uhEZBXHIPRTSukWHnuZQtBG
Oe4m7GnVoIn6+/dLkP2Rrzqj3tybH9LH/tYAoKuOS2txLGMwLojJiE4L6ytqyWW8
n4KTfpW6EVIzvTiS/aBT688XygEN0tPwESErLwLOcryKKjBK6/B0u/FC/47Vrx0Y
NvA9k8UvS8CYe6VTWAP9ywsYZ6OLoALqQ/np0MuGvp0+iJAIL6gSSgQJEp6rxbY3
leQhqjcZqa6JqzlmL5UJ+ioY4pfH1m7rHSkFHyEcbtoSr5uowCJEBoTTuJD1HvpI
riIqVT+DwTA4kySZy8/+crNjZDKLVWjZLY7Snox0dLpYutvjVkrMdSA+B3cddLPB
smI7JpCEMo2pXdSltCMRjIa+1Tg7AySfZ75dLQhCswfZDHDVskuKVru+orfsmc7c
iz0XvJm+uvz8WVZF6VoXt16R5SdnF+cROZvf6dBvtmVIeP8/tERFAq4Oy8aCvs5W
5T/f5rMw6MayrsT495XD5j6Unc7wUmO846OGbeEci7r3AVzBqlKBFgRujMm+sdvM
zk3RnSHhH7RDP5VPmAEpLhrII+HKVGUgnfj+JC3gjJHGR48MaSeiltSUlicrqFvN
MhFH5Nch3BYl9DP/pmmDDCf+X2zTEOZBLZLTDk9tfnA/h+mtG+9ZuU8bCOsHjiJg
gPPq7BmUIv7cnEfDVQUXO6Bxgg9V1QpNntKVF7qQRRBw0wbVuI0HHkdupzqrk7II
wR6wqyxloA3IcWUPUeUQ/P73UfnWQ1wNZprDFSgOrymK/37VEzVubSw8MppThsWp
uFZku8RBx+ru74l+CGHwcGUYhq20l9A+2JrNCvnmqDE75JPUp8ZLNeAVD23eclif
5QZ9xgY8GzUKkxd8C4LSR68dmNZBRlmBhcGmI4M69W07W9XhNYnA+4vLFbOt5cb4
uFXfN3gnu4w8FWjJepi1skJ4ShQRyJLO7KQmd/IcQ04mQUfxjUNfTTVGD0YM0E9c
brfI1kwFaWHLQXUnpcoZ7xWF2HDP1LmT/xPCdg+6b05niEZlFeoOhDanPSmxYBOh
dpIvH0VP+QQTbNIogux2B7sPaOKC50uutryQ1sTft3Jc0MWpfiwSk50R2ZskGcX8
+43ZqGIB5PTu5vRBhEulV2acHsChKYoCkKARXjQi1MbE/zg482+bIoLkq6cQ4Qg/
3pFePh8FrNm4XIsml7r+LmbCyRrGw6EuK3Hr4DrovlCimoEP7Iv7SxjYjTQ3nkWb
ljVuwM115pYB3oWWVp/Ygyji5p+EB6Ke+CstCwLSpg08/+tSomSo9WJtVxsUp6Gi
FB6ZqR7k2TAKM3tH/xEtEzlS3t6ij+ZzU1J+/49EBdixyca0X8CXT4/DHPa3H9Ss
TjvziMioNQmb/f0B/fiD5kDfUJk/rBIqISrdtrsMFTy+GksTgkxTYUXY5fEPC/3Y
Wo4CA9z/XRYUcumVUjQGVhXyyOuSULvwClMJEuB/Xq/rEO3bkEBj6a2PXH/7XY7l
/+bm+bIYMfnPtzxfPSW/NUjini8NhnqK8nMu43AvBGZQBsSC++7YiZID1RTnWQwg
HkBq9Qxl3oeOGI6c0AkeWxPURSLNVCvzFwLbvgcgODPvPxpi8goUSUDG0LmW+QXe
Xb5OS+aGaBWU336aAH8/nw/iz30J/GOxV5IKTIYrhm60sMeyZ0IpyK947zv4cbu4
wDSRMK29UeZjcJrYDpIzUBugDvS/51zCA0NIfPFjYfkdh6kte37L1EDYzXB/MYLR
xXBlm8hC6Z6Mw7kBUJ6BtuJiOMY46qiKABUEl6S59uDk9e6YC/GQIfGIT8ZSEddj
N3AaaUzuLJVzE70dNVgLJM+n76Dc6WKSPrl6v7mo6knGIPRTSirgbCRgFiAbvzc5
vRaMnXYG2pyNGgDcvhuzSiy43cXSVPTZA0JvJvXOt8b2BMeY/xzgapSHJA98QUWY
3KDTgvmCeYlN+lDu4CGCeABSmxgrTKB6ns5ZUmEFB0TP94OCTZU2tHR2M8+lHQBs
0hHM3tpSxkfPi/h+hppBgElWt35dXeFG3xMOA2z0j6RLWTbIrxd2mpW+gqW7sWlG
5Ee+ul7VYVYoXqtdkmJ5ylN4Eus1XldUIVJbCvurTEg6JTbT+ex05Zc1V45BELO0
yOXf2ZNsz6dYPKYscU9fqq4JJgm+aUh6gf9pCIqnS2I4sftuVb5SD6/cwl4Umn5Q
32+Q2vjN5cvq4SOeoxtdn/VxBky7i6PfL8o/dkVI7r3qOW6l8RcFZmcwP6h2ejNB
4yq12gHspaG3At1uTp7ShYB9e/OVZ2DqPtdAwDFvwDTLTpMY2ZUkx2nWoasmvN84
yobPWJu9dc49+nv8VHqvd9Eww6aZ+sJl48c0WyOdtyHb1pv28SkGo2EAjheanAjC
EQN3VdPgCCGW40J5kwq/xjL/wAbtK/VD+O7RE50BKlCdw1Rx+3RDh7M+Wm0lYB0C
xUh9iIz70HqYiL1PhPzNGPC5DR5qkDSlZt6g/gMGXbqA1WNlxuxtkCbhjCR8B03U
m9dSdaseohX4mBPdNuk6fNGDroGi7MlsiINwv0ge5BTwdYjIyRgD5BkF2Lp9V8I+
i5C9oy/B1rMtY1uS7SnGzqP/gINDSHMesqV0Gj1IFcP08C5piftFzOpnzlSjhGWj
xDBtWPORbseHkyoi+PQAzxGnicli6SUS3k6erxE1BbravliSG4LsQMx4M7A8i8yo
mvZCWzEjIMOBTp9nhZtqkkU+ynYTssHB6zwcyLACiJQ+9jOrcBSpQo15iiazfoyI
RmhGKr/HuYJJnRY+jjpfWyMhWE8CIClHVxh/zfc4WkDKldF1SbTK4ZuMRTvheoKz
AN8lQVKQFimubPdCfFSMV1Z+89cAnUp1QEzc+whFG6MEOoK3XG6ebRM9TkrjBoMA
iRb3R5gYtkH8UPhEdsoA/V9NQvKagAzt3W9EZKfnzj9fECRsWzjQjJH4smBUYl7z
EkoHTq+EPOw/ozB1zAGeg1Z8YvPO1tLsaMvOs8rbBJ40GgSe6xvqNKXls35BYgtz
wwx87P7c+KVwm4zFakbZB0EaT6pTimuyogZ3FKHw9kl09GZkrRUzrI/OeF++wEf+
SXRJiNklMewUtWcd7YfOvwXuj8HzyLMqPyIW/bFzuxrNrfk5GhuTKSMZVRGSAVy8
zPRJ8PqnirU+1Xi/9wv2wfGIyAcYrNCOjYCSCT6oGZLllEnxQYoPjgGFp+TnI5r3
Nq7HLg22/G/YiAt18INtrZ74GoB8FghJW0uztCvhgf+fmEerlmzVtwmGcMvT5TpK
PCaacPIvVh0BSEoKB/hd7owLLLVR/WwqIuuMTAM9c27SHZfEMQ50wVwLEiK4tRdL
1UpxWVCHPy1ZeJzvuSAfH8J1hqjnmBdK4hij7Iir/PBH3HczbCteMsr1rnM29wrE
jCfOaqX4yU2AjyCyx72WU4ewckFZoRQyiF0nIZxNGmJdfzF9Ufh5ubdmmOMWf4BJ
A5tdBCWYNVylDIhpoh6lzWgK82LewwTpNkbHg1hNN2qvqX2DxTgLrgM3Sur7VO3c
+m/0DpLQOT6aHhQEmSeQ7uwCPKPdBkQeeWkQTeIcMiBGSqw1QVk0fniJ0HARdAl2
MS7ueQI00EGeIWyzXvzZBJRTZCYvftjnYWGEoJ9wYDcrRZ8u+HJRmZ1NCpU92kBm
Cpy/X2D1cZE87en0LEw9QfhAwgc806AD9S6t5hmB0sXfRRPXzYY4iybDMNSZi8/Y
nMPO0W3nZWqTNirKVnToDxsSFMOGUwEMAJCL0yCoBvET+QcB0kOaTPA7cbQcRqnD
U6V6PmUi6CFy0JjSkVQ2B2V9ZwV5ZG4gcELvTcjp1G6rtcbCmjelxPqJu+UplWZk
pr3gr3fX8SnNnHO3GFjlIzoEbw223YIz7H7C/oHegegcZWrgGsEHMySvAXao4JCo
RtelPfpvOhmCdyhE/qItnWKdtO0kUy1zJ2ggAxrRXKBhjpT2KnCgbsJo/HwVcPfB
bQlGoCPrfbMWhU4j3WUsWua+4G68HtJZBBPOhyIeC+jVwxYoBjqKjetHfiLhswzv
4xAD2enGvqm0smcZ4AmbLURuW8k/piWtqlswj/DxRlT2Lui7aeIhZw3ZoIaZD4G6
KK7xE9F8vI9tKluG/f4ZpP+Y06dy1DeWiXHkUjl5Ol13RSJUbVEj4sfh78EmbJO8
cBNMScPlSk22G7clKP2JD6OkmmXJFzb/YgeEzdRMRJ09Fszx+oEuomFeZMcDwE4U
MgA51+jRTXFTuI3UkePpe0EdkWtuLzex6rfdM7O+qASg13xjBpRsGpPF3Gv+NOfp
Gdsm7eP7q7OUQsAAkJLRrS3198ZX2lc+eFuY4kC5F+i0RzdsQ3kim+Jl3Rncipdh
wn3tsPrr+2U61h/b/ruA6REgr2rjrBewOxC1mFuuZQlON+8Ot4kXBuK0wfszLvRr
F2rjBKFvcxbW75gbOa7yrTEYO96COWGkVvFWlwGTu48Z00TZVSga1mpCOWS1m4gt
Aii5SiKV0t8vGdEvjYhIxKOfEHSJdeqSHQIzoP23V5qlbtcwmfwRLDQiuxgfWK0I
1tQmtAPpyoBCeZJUeFt4hp/N9Dt2B5e8MPSwPKNebDJLwmzz4pwjeY9QWmVboesG
4kEDYhlbpUJFsWyKPMXvtotWKQ88umOXqiFwFPNZCECGsO7OEk3anKgq8CqYbAhh
NmSkgUQXk8Anu7+cGp42mQGyLrZ9wZce91llOZNtGDVgy8E9CDUSFfLrZJ9+HrZ9
spHeG3Fr+lrXc/NOYOY2ecWc9aiWGmnCqsFr0AN8Nded5g75MT9knWZdRnnJyzHx
QfYlvxB8KfelRHxg9Y/ADm54H8CUAMB5MNoPrk4nAnodVb+C08I2s2XOYI2RPLMr
NT5/ZhETLvHQBS8xDd0IfcQfT6NrcA33umq0UHLr8d/1j622Rk9NdIRcZI4rTx/h
3KNYrd/vxEKn5D5WIjMJ+ztE8J/NeX6A8sFxpyX/MTsc0oJJijGeB7LZ9GUBdeqV
1elYtbDKMbZAUHCFXMrfHbBtuRafML5ONP1G0YKPbt7N8Spdz6HVYcvHlNTrUhGd
YWopMvtv4uNCIZWfqO9xIP3ILP7Lz6fO+opWX2DXIdktUYn+bT8L4fhmXJdFDt/S
4NnmZ3ZomdZUhlpputHf4ZhdZs/Tuygpu4WE3/pVwur2xUSPMWmvvnkDaIv7oAd9
GUpQBQgVGnBaShvaffHMUPGhwMvxvaA4WZ9++dgH/TKMWDzEdMZaaQrvtaRDSSHA
dfWBMtQWoX2f7n3ReJDmz+g3GhLvCt3Qon3+9p3/Fp6NiIH1lupyDcEcic8pdp2Z
YbLObDpYM4hXVzKsRAyWx5r/vzGm14Iwywn4zqmCXjy9su60xnJrT4x9kNQokKa6
DhlTbKx+7kR8Q9GRG4I3B/+UFhAhBn6fkgaU5Z+zDzRPca9S0qk3XJ7JNn1bl74r
O6lJajEcwYJ/dka+KvDYMmAPKg0+kBhNhcpYNuJFqHYMtcmmmjPfXuWg86oj7oeE
GmL2wDjb2dflAvprFPxLFKjra5BFg2b6RhFMmeDw0WU4MnNZBiD7DEvS/M43G1mC
+4Omybu0mKI0+qkERveOucawbaXD6C8KyVEV/H8Gzcxz+AmLJ3mYQp1qfF/T5kEA
vP+63KtKT74kd+URSfITfs3ja3GfqnzlIArd7u/BmYy+DNd8EtWZ70Qqx1g5ABtc
NQHiCVHImW9AGAOAuX9C2cBjsyvzErYYUfNLDOeQ3jXCel+JXz0f5smrQOdaYvhk
9ZUX6oBYA/D59lxgjwte6/MGbpagdTNsmo4tiiXxBR/8ml4qWD2hUVV7j4l4EYt1
Dz/pnUBhNVyzUBFo8QZ7o6SMUYidvfQsuDKbDH/VS6KfBuXmqxcbvSsLsw5vGJbL
mV0bT75vyj/n8uRs5QwurC41ow2IOv2FnzCK8CrtkCHkQStSCDiIOtZVUlMg0pxF
bE+fM78MZjNrpUkB7zhR8VpGi6LLxFLU6B8SdAQF7P/TW1vaoPwPCSpG2yssm3uB
DnmnhSud4FQKllfQxGeXnuBaHIt0/GqZAYo2IQS3c8D4qlisQSuSpVqeIZXjvtH7
cHucmI9gN/fVqzXVM4qhl15ED5Uj9KSrxzDqcgUFKwu4VqC42LCsHqXrA/QXVwPp
JZZqPsaJ3c4WR3t73IihqhuR4owXhO4acOGp6OcuKaY1BBCBsEUnTicdvn1lqIQ4
jRAN1OUOSPNqergGNTTYPagTYcIT60krtdohevWAJqOBeb9hhlY7MCTbsnc0aN4Z
ceogsFxjNsjNnRScFAeKmoAoyFLOG7yyYc4D8u7q04PmuM6EOpGygwWbtiyfRG6p
bpUch0DvobuwpKGgWpSurzbUcxk33214ZjPG6z8JFLcyQq/S6z/AM6Xg882fuWwO
koWCKfXpqk4ncT0Dw8bGI+HBcapVLK7rRhM4//89YuY+LKt1rx9Mgq3Xg69q7BkG
sehMO4vO0wsAUfoufVzsGKyzwmFiM2RsfURAIfjNs3B+Z7wv7w6Qvm+qQQqCvKka
IB6RmT6JA17VMg3UTkd2RuOr0i/EAheARaJ/aXOUuTi/n99iUt5kzthAr52co4qe
VQTn1yQy7ksQlM1bTCbQL+2/1xGSz5PNhZ7h860PrSAqBjb4+xGnpYyK7ruwRZZZ
+DESBe1dY7U4DHvfWsXwMLa7vkAxR0QeJNFBOJ5bYiggD+/tWal5de4pNvL+BFaO
SF4ziMl368Uvh4fIpozjFyVMX0uK6Q6hCfKVYNEXGRPJr/FXEXU0PmrO5xYRYNxh
En8Z4MGq5ZwFHKDXFon+Nb/mZHxoE43ZZE7BZLT5JnocAx9XR7TBhoyomqWxKKl/
ethXwLM5JfJIuzK8dd94gSDr1dJ6wxUC7x7JWh53wtbICCDI2HG+T5g+4qF0QLtV
eez5BW0SZdC6ABLpiqjmuMm2ZX1tJ1VUIDOZX2+W6RkJiNp7f0bhPHE4mKu2tMDF
NikplW5fA0kGHBrPR4nO9J83N2Ah8MXH+9t2QG/IK/L4mukAy3A7C4BMl0DEWzaH
AHDpIm44oSFRaBMuBBjDXT7xK80gkfOVML4b2TEHrSbscS8Ma6wJADzjH8xHQ8De
cZH6c2LEDUqsL1EPjTDWdLzPWai/jst/l9+EGSvh7XmRgC8MYWQlGsJ8O963KoSq
mQnwOPd6EdBx78bZ7CupqV95wzNLlcL1VJmhak2zdgMfscI66JJjglSwt2wigW6g
Q4JhfBEQgzIpxs4eXNWMC6GJu6p1SKTXqPC+0KHO6f35kwkvBLYJXLVEEH4grQSA
8E05iHJRVL26/u5Qgl0arLpqBVQe7Euj5fLgyE80uQEZv1XtX2HZsptpoQ/8brIc
cUIO+Foo41lNXLDPDsZnHrN6yY+9rgxrCtPFEnyJFYZ8iISPU3Bbt4caxqyT5nEj
X0lzMQ/LjBO7JKrA/wVsB7083+zR6XNi6W5S4b2CI75T6bu6iF9gFouVVLRdnX8q
Cg2aIGyl2INj8+3o4YsUGlAN1rOOMQmQZng0bXItQNxUqeYQn2LgaNUCIImLGIfR
n2v1BkrgDdGysvYnuphtlgNoqPeN+tcX0xUKq5F/v4RrE7+Gd+90h8y5lwVWFxUz
ZWE7jPqBKzkzyGPYNu4ASoP6SMZMsjf9oG34pGqD/irxYyqppISw4BScoUCZ2a80
MxMSSDUUXWLtOxdIkIiZ6v3ZFKwkOqp2V6iryXJ4ztLHl3Ki6e5G88l74NaB1Az7
z66CAPwVGt2ydUZKk2svmt7njJOq0LicpOFQD6aw70754uWeDgs+xnj/nU2sY59X
atHRh+VgO83crypqvM1ms8Lf5qqOa59XDoHzz+kaLsc458vto7zo1RTXMW+lvBl4
141Vbps8RNubqWavuCIZabz4tUmHKAl8y5XgO0l5qZFgydb+M4UC+xZAUXTdIfcS
hmp6Tajia7v1/AWeWthH3cHnBbIO8tygs+osaLMZB5SLkCJWncs16vwEtrIS0dTo
/Qs5Z3CNm+PdDolqw1LADcte0j+zJUPiLHSgSnY7u59L8mwEVE3H+z+NZExzOF8h
gDsNvzPtrDjT+X4amfv+xYhK+w8JV0gFM4bO7kYKe5vTuFEeWDz7IpSBh2K7BFeZ
vsIWrGdbSn90SlhmNYoyekGxqBhOFC7MW61JDaflGSe2wL63PRyhYIVnW4loTdYc
JqDOaCtNT2y7Axks4qYc9nSdVGMnmUiWubdY1Zwa5UyUqxKU3/gIPankgC2EnTs9
yYkh3GNMQOPg+78w1IkpED/tK7hEAqf7Dbkt2hjxudh+tMyz9lwwi25dTqysz8iG
ZrqiQxB39EvlXXOjzrnrXJbg4Xs5AIIzHTAOTDvSHo2KUZHHAlThgRFx9w4tZNoL
1g9yAkShghYTkis3KlHytmD8bmAw67/Pc79JGPzZt6Cq3Vext3afIeEhY/nzGtRB
9Po3fN56/EO0m54SrUdfK9N5b5gddUWqINzo4TNhDWSdOWeO5DIgDE11HUYAYwqr
cjiU5djFmdXT4wTtfY9+hk+69JlTjhu/3IUSup80pgfKDGof4474ijvimcjRyzVM
izlSmxgUmckEJLZ/NfWV0HceZmsCjpJ4jnFJVx1GhVw4ZDsz+40bQw5ruy8uHHbM
MBdsWr8THT0EvIqyZODOIBbzNBUr659gQsT/rpKRYhhNvi13U34Y/K/DbltRkPkm
9iWLdwYw+Pawqt3FZzv8BH6bNZGQpOun07QymjQKx3oQ9ACgsyLfu5Sl1Nlc/ydM
R9hZto9uiJWGmsQCwYOT+ZvMuvkl95G4KdFj/ooYQ6GNXA6GyItFZu0yOkE4sg4g
2hrGZ47z8lCCp2Wk+PjjK7wLMPy0OLrPygnc5xZrncSfyUbSwQcOBVQ4+hs72FYO
Oht1gN6Q/p+W02J8+nCWSf5DCwlCUelhO3Prr8zCwkeLNPxcfk67hIw6kt9qg7oQ
JT1aJIiijhWi26j4gdyDdPJgLwQNqrT7MNp6UQoUSqneFYQ4JAVsxZRRTKCWLo3i
vHm8WII/1sSYg9fbDNOy2mKBCI8Nzn2RFNzAgfu+BYZtyGk+t+ezb51+8xTjDmrq
XNzbPOg1iMBaAa3zYYpPE/7UZxFHFxpEKoTXncph0kDAGFChn2R4ycezenZXv79n
sVSSF31xwrAvQLJnlK+M1qjJ6FiwzUIMOFeULzYncJWrra7Zwabz6rWwzbYIUgza
UK113N/uCnWbnstHl9s0F1/I5ORtkwJGVg9JhAlgqkJ1ErvuB1i7z7zgdfWM+Htv
iDvAmG1AdCZei6I4VGRGFJys5RMQD6P5UtJII0Rnknzk5UQSmDZrqDTyV1QwbkLp
Bnml/g0w35yDuMsjWwyLY4EyXMC1ZDOi7/CuRdCAHRqEUz37ZZ6qTR8wFhx4yvn7
sokWBJh9rLt4kiKSbwGwaDbgaoKJRMDq4BKNzi7AN2acp/LKNjco25mOXxE9tMrU
bmm9DGSGWicpKV3LUN6rYum8fPDeXFJSQ8yckm5MpcSaQWExA45RdlWQQ3wVNbIx
EGCs9G4mrSfvmMwtch9R1yf3WZo10qqduS+/SqYxsyVaR75rkt4r4DLp1nPZfd2m
5UcvXmPa0PJMBVFBcB4vZ8rqe7v3qqz4mMAKBVUXOr2zgiEcn6COZBgxP6Mmh/ij
4w12QaDi0Z4bj662I9pXoIVGK+7WJdeukzZzSAXgbRF/RcICK7q0F3eqp0lQHjQO
CtL24HaF2be25Bfb9ilM50Xul5AJf6egrfEm8Gfn18SExwriZij2XFUn00lAgDhl
Xov8iBmcwD+lUGwLQZTfesnV80WG8GIdhfOVKbLj6mKnLu2TZVqGrrBZYzO59VqO
0JsFWIGp3lkP3kJjL1PN/4PewELc54yJgLIqSsamOsUL4z07/LWb62RtCzLnL+bw
EbgSUrNtGH1liZoKW4bUScQJQVBSOYOLNL6m4NRU8hN/EHtILZdJGsVZoDE7CI7+
FxQdKkDQ4yX9kkqJxvkeFs0n3b6xWqeg6n8TW0k9KmQoFY+gHw3DuygHSaxxNGJd
pfYjU4Xy8WOXJb9kqPjVQZe4Nle2E7PRG6XYGHnwy13MjOizoMU4mwENo1lviKNC
omn7qRG3POC4aezg6+AyJTi8njOlJrupnXto4TO/pJ2Ty8jh+P4JurJAS9iL/tZO
2xVAvNIP7Cf+/Z3Tx1hA0mUZ/Vv8SkFYoyTNngTv53wNbg2p3ngMkGHKrDXjfL8P
idLX/km2LHcWTvv3qO/95HbAWboDb7lI1MpGR2gBEXIFE0dK9l9oUxsW2XroG79T
t7y9MaX4DQC4/A4qCx75RMmY+lIlF9OeVZ6z1Sh/bcqaFolqyarqQGqjQEvmOFlV
NuSthgqiE4t0BUQZnkPs7sAqk1WGddqfYx1LjOhHEC7/8m9j2rtjws1uwz5vwKbS
DdBr3rQHOpVnnY2JoTiY2QWVgtuisRNlvsJpK9Z10I1i/zuZ4clTMA/7fGKnyvFK
d6HBCVnYGCpUUMMTX/NLT2eNEi7/n884gOg0uaBddyg1kduULp6RBvX1WC3U3qfV
Hm4D9r2Sp9APjyYxXRxpKSK2tR0SlcPCfw4fdJrct07W6HJC2lnOULxV5VxMmlxh
NTVQ91cB310O6ywjtm14ciGC+xL+m0YsipZiiGIL4KLabupQ5mEZHuzXPx0CVjBZ
LRVuEaqJDWyvNkvOeoXC+v7b2wJg/lDIcEddfeaKLXQj1nIT5dWSGqU+pHmRrXAm
ZP7lyywNIDFq8OBEClRW1vqN/GWcMCiYAl2gd8xEvtn7mBUgmmr37px8AjMWUM9l
VKoMXaa6OFJZdRCl7CgvG1653b/ryAm0vyabrMZe77ThRB+YAMU1vX8E/zKexlff
uptgLa7iiRuUFLFRlNDap9IitVg9m6Z38h16AAZ5B3S3xH9MQgxjVhFmnyhUvNjM
9uxwpbatTU1znbEuX0Sv3V97SmTZfioPu1NxpFXO9DjYhCXA9Y460GKdsp7sVRXE
M3aXWSM/fYkDkXfZgZoM0yIOpdmfV6Ar0RNtc6K302YH7vuK98fi/QHjDsG02M/V
Ggb+lB/ZEryhWZcPHYpz2HZd7yU5o7tfWtPXvVTKc0DYGGp0E/azklCTxufx92H1
ZMRw+33XlHa24XVu/wMmSnRqe0ruYTIHVCIz/MXBWwtsD4Id8xy5Kn+HJNMj66dz
msqsEt6L48jOGla+uq/2G20e3ZDZvXJDZa4CRIumtcnBcStZ2S9xaQnLRu3pCw2M
pUeSnwI5F/qXuBqCC+u7Hh5O2sPPsan2p3QTsGtNx4iAJMXx8ZexfWjblZhJid6D
RsPaOolpNQbNCaFYgP0MY0YlnQ4lWolyyXXir0K3I7KDShiofzvICNQcMAqo2Dy/
bnEkS181/9M8v8Am/iQdClgv1LISC2svU4PcN8XwH6nupgSHQVH13EI4ymb4jSPX
Jf2RvnKLyjQ290NZBUUkaWODySer0813rngsCG3pfXp9SxmQ0aWQpOhlYQX9w6dN
V/gtQjEfIaETwK2xTDxYJuKSe1nTjDeTYP1y5usEW8N9WXsKq8/2jmtG0GBZGFtI
jNdUyL0uPW7n07zxXkEW3XTqZHYsB5x9S5u+1liDThoQsE4TD4Ue3tlwjEnB0kMN
BeQ9lfZqeBsEqCPkGjO9vIgHZla9HJTboCTt3hmYMowNk0cr1Gl1kaUL0bSgXBYu
5+Gpm4HhSIWr4Ay0PH3V52Ti+7lKWWzZwtXXaPTkMBsU3n/DZUs6g8vwxO4UH2EH
rqkv6eVhYYdZV6ViexwSkp5EDfOxGw850d1Yv2f4BxgDbgmwAyxOTByS9JFVG2uL
ar8V+FJQ2hBh0VOVl/SjnzJjLIhfAyxgufSuxwbNuLsleNIXN8yFbnRr8KuCCQIS
5jaVCnxdhqEUE/KnRY0bYzHGIkE6Zo7oorXYseBsudNm0NcjNVvPyhU6czX6xSjP
rgkstWJm9Y925u0PqbGs4s2ExPjUmtpzZwojWPflN1Beer9UQMwDRejaq1iynefX
nlrdvnTcS21i/0+5JsJuUNYtxpPt9yNCkiEfyy7vKpSK8nTvEKX4tUDzWX31S6Au
be80WBwlCmYp0cpwpofL3DFTC2kH05utAFWHh0PT0hSVTmOa0iH1/ucmpNB3L2Wp
z2lYmvNiMrbO9OiID0SuChb9Lne6OY1XvnhuiduUFB26J4oe5vZ6SJgGMpXGg4Kj
uDn5yC2LFx5Li6rqtpL2l3/4V73sRAp0lN4+atT7BXCZ75IgWtPHcd1CSc/bhDwG
rOmKDE0mUdzqibYPvY/6EaceSNV6B7+SsVQDq84I4OgjJMPlqmhA6lwiBLI2u1/N
gHlzGzLdVzsVtJgUHzWGIZIUeN08LtFdJ4YgeqUtLzsTolQkCr/tHbgEcR0CG+YH
tKha47wqKuelgFjiJ6bINB+/a56/8kNssL4zngjwJjiCMfZNYylJMfAP5rNpS54J
E+qsEbgCJjbux12zBdvWPMxVm5LRDcVFaL7BtMg43u63abFi8r1oJTSFIzO1WHmc
535MMcJQ7MPx2r/1EZOewIuzYnNFMJpFb5oiFtUGh/CIPXt0gkI5/qdlq1f6X0SJ
azq8KIKPz61689gYwW2oWDHj42B3RHrtwq1DtO9fuL7Mq+bGcJx//zsZEmLYK14x
g1CUusBKew/c5Ke1MDuRNi0jjILYTZQVeEqHITtqPbDi0ojGTP/rshPkHiWaPzA9
TR+Xth9W1LAaRRxYBF7KYOqGuJyfI9H7a4H8Fg0cuTPriS/BbWc5cHrPBDaT92EY
2cMLVkGK8+dD4IJjwxeVXThMS1z2b3FuA3FJi8tj7WMnBfH2g8nNwNXQIjnFXIgX
M+yj2+vzg+QZGoDvLwthEWFxo+baIIXROiP24gNY6/5bhtP0zLlNuHpD1X6ShHCs
f5iWvgIcaxts/h22hdGmYAU4MuesUdMKO2YwKsB77sq4AZJcNzmCflu+qVk+MEeW
oo2zB/wYHu0pVpmlOqlBIfchM9Lp7dxVIuh4zs+m9p900OIQ5qSiFgSjokULBeIn
qPDI+xEcGopKOjXAznyDbtmuSZIB0ztLq5q3kLIfqn2uffijLPkC4CKijFeyXckT
t/efQa9FJRL76XNpDmOjvxrO9Xl3ab9V4oDDJwhUzsbhKSAowxRVUqvpQ9ICX44W
yIalO/NtuZ8E/PJhyYgMUy2zpOG/cjjZftp0668AhakJ96sDQB3h8DYek7joVkYz
xI0iJlq1TlmWMnjkIWvAE2WjBvjYAtTH66JKi6aW1VmFuWnWa6zWt8wJ/AnRtQYW
iy68irrqtHQWOtOYSw6zJ8GEktQxfFVDmz99eQsZ5S558tvGesxHWxIdfBJM1Xr1
lrbWyprJavfHudIDXRq3D2W6Fa0Y+TOAk/GA+A2/RlXV8eN+99woOUqBVs+DJ6Ae
I2fe/nNtt+QKMzGY3eIEmcNZp/giuyCMaCA+Iw9BqA/pA9zTL6+qAkhNFaga/Fz3
v5zsM4IJDC/KdzLt15Di8rwW1vZ2qKbT1fNrXVckURRyktoGQPTkAQkpS/J/ib/p
uyhZZaUi+xbBAgLdQuZuTIsL9sWBgFqHNX1BGOR7IchyAUb+kKgBUt/xm4Sjjulw
+zs+fjsMWuNA8v42gStEtI6uOuNogb3L5fjVt+DYPQI4mfrn8HHBPJ85wlDWGxpd
eGkvAHcgMJVgKbp8/j6nMXG4Nr9lt/tb4DS9ZzYD7Rwnm7kzuhiQrhLZCDHN4lTd
AMwoLtoYxu646+A8NuXdDSqumz/12yWHmLveHsmcfgtBcGhbrNcAUzvBPhC4Menu
oIIrzXCNmfr4LqWXDEso+RcFkfCQTUeJgtDuKUWeuK7i5UEiz3Cb1mvaq8te4Pal
KuzP14OMRtFk84Dd3IRHbMFInIOReC8DIaaOE9jIZMVf+gvdGPjm6s0M3TVQSADU
D8234qo8v/MAgBGTixqD5v1kgSjUztf2+QA+IPxplcGclH7CPY4OMFYh7RJY3IEn
TCOuh+jsvuTZg8o0+XKzf7WBrI1DAddULehToMvamQH2noMWS5PrnIdvovOoyBYO
zCFmYfcm+SoR+JMo/7J0sQcxzjtpJ19xbmwxJw1/46zWD9IX0PR36toDe8C5sqRD
5yl+3SD9dPs7a3hiduJq+c74kybf27ogka1UbsjKsamWxxWAKwtgDCGKDX/qoXLH
2umVKtbCC8vppkNVcpK9lhTejKwEyb75roLAfBVReVCKrMiDJSntl+jIAdh/ZJNs
d93iLVkmj+T88MZYZ3ov+YNzpds2h7Uwuizrn6B/DPAvJ2fIHkOSotV1rNs4m2Jp
6j4Xu4JYtOmVj+08HcE4d90xwt/z6NVI4BkYjA+v1ir6MWXWjPOBswy9TphNWtUj
3tf2l38ujMxJZr0itrWDFLZH+Z9UPz8UoMutVctjXXWxxbHiw1jYwXtOiua3DKbq
4w/Egig6I1WZtZ9S9b6R2/PvGD59TRIVBn6oZuB1HCG0ingJbYOax7UNvchkkezu
5e6HXY+kRV2uk8ZMV4JSOeAdllMH0qptfTXfkZ+59N1INLtLe+mzupD9tuYgYrDY
5U/SEBiFX63Kphv1rH+63uMGQ03C+tTK7MEjihzgrJ5vwQhXych08tcad73YW6iE
+jmRf2MPxUH96Igog4tNSOPTYnkjRKCPRIgnx6n0qxogQgIwjkzcBUO/dlpOV8V4
GAa7dMrFRaZP7eH4DCznbZoJg28A4n9SQ2/+3O9glGWohLQoPrdrEijF+nDvQfE1
vopdNUOGu9PNLxYij4XmpErZLts0iUWRMISH5nL6K+I8Frv1y25y5DBh0zdTlwCw
7LpK7dfTWQGrH8qrXo8ZD5282d/SuQunat1ObEjtdNgBujU5bocbqUALUGTzkhJ9
zbTz4mVVL8ABRM/KDXDlSmPMmYOrX3xdnRBKTy2OoZdZhmcTDA0Q+T2NqPfi4fm8
8d/bD156vtmdIBOUQNk77od3Y0FKzNCefX9Vwa9kN5LxyJ4jwKoAcNhkeSmpf4kp
zI3y0VjErCspz+I+MA4vNdFM8mnL82FSPh4sB57NxJAY5GQhkopM2TCLXHDZmzid
2wUL1g3SoLwNXtM0FS5fjZTf4T4iut0eZx/HZY2oCigzY1dUyR14ejIch+xqXT5w
/Pb75ZBs1jqqnT45mWEyMmw/psE/bamqzGqlgyKC4tw7Mh4Y7s26GPM3bWOMGXlC
yqJz6dAa24LjdyOVVsyQidiNIB7BC1WB8402qVTRWZR0ykE/ZVFTdTJugnx/bYMR
Gt371xlcCGI+VHxm23mNOZYx495xzoffdWJ8NIxlSzkGZ8Ax0yp2OTnRa8fNTajy
/iaVPs7+4kQadXpV8bAfuEaNm99ZbhFU5udB5Qjj5uWIvOYGieCzkJBpMzEc59Xo
gNvEGgVN3b1swKjpFmZO+DPooid9ik7r24ZWlWpPmWdNALQGqWia2PNno85kMlX8
MBArVuby7Qw+RT8br6yF4uzeZJZ8dVVfGs1bXSdm2+AtXnYdRWP8SZXdU5fkWwYy
4hMOa7a/KyEhmcEXh5dsdJnapV+C619CX4tvMXfC4vJMaPuBDRAyz28av5k+cjoe
9d8Wsewd4CtzXdJC5OJO85gYmqbtUaGfKjTH5LJHHg937r2p0UyVD+00IowDAR1H
c69PEUCxivhi1DCeictcYsLz54o8hs6nUwxghl8G1oxyWWzp4Ie9hDigU0LqCcdm
wakX9qqh0aBmEM7pXdCNzPyiNgrBUznZNVZ72cdkmJpXl14ZLHV3Wblr7iPENRI/
qJXUy/RwX6vnbIb/6V1YIoY6/U0sKonZ81wpR/l49sbCz7nww6V0Qn+RgbI86RfA
gywrJwxa069tLxFMJ9aJLCl1PNyfvchHDoInmVnD2JXO7gEuMZqNheuMd17Tt85/
eMI3Y4s0uRhBrzIuB6Vz0+nyAXGC5vARCg8vxvWZnl7uiWg+WIUZUGPkVAbts9ip
4ALk5hh430jVYNaAssxL/DFjS5t/vJKfpRKiuLoSzBskOq/OhyoDVrRtNBUtNuOa
c8dqL8TJTB/ZlYud6QOujkpYoiWxyAEjGPE5RpxrGLVpN481eBYzrnON1U2+rR5K
x4FmeUOeyPVs//jNzgDsaXKjmkMLIdstiozillXAos9bB4bTo73iProrO+0plZOR
CV39HymAyA78o8w3E2gEpDlHKNDHMFja2sesEfyOl1/WpznDSsnjowmynwsXl0f8
zFsb3o6KeFqtrVSNKGZes0Bx8CIKXSL3jpfGliZh+44ivOQEgKRLcCLXPgw1sQPL
BfTepNhZaS49DTIT6cyARp5j+VGICLEs9D3JAqBcLIBSb9/VoEp6S9eKJ5Nn0WM7
ElaFdf/RqEEHZRvQQQvMD5jldAQ5X2zmWzb0j8E0MQQiFEAQ1APQrflyhloh6B6g
NXVM2oOW7Oishm/1WYpot73Wmuz9HBlG9dePJ0hWdSAcR2QxPcaD0dpzpc9dSY6D
zFhGkSs9SWrD8OCPod8EW62eh6NHbZyNgtnEaQKMKF+GMVmJCpuWHKAApf34vXuc
iIfoPV6FwN5mG4CeSduGnYhgzsay0YcynH4pq7F8qTr2kCZsl9TmbSyRoRkBmriS
rPR6qn/mXTJorCIFB7SvK+X0Q9ELH9KZehY+4YndTYWW4lPoOXNkMj0kMzKPbKHG
9i009Yhx1ayJzbjcRfSvwWpPmIvkbd3ApM+xJw44V04etMxDOl/b0Mmn8E+1akEi
LnaP44+9WDA6scsVGPL3T4DJ7WQ9emnmJgoogyX1grMTC8ZbywUuAtsMILOTXHdW
aDGNVY5GTdqDapPTYNF/yAXlgdqW5UPR8XCQqlzk7B1dKNqE5SQH6YwXamqOseLo
s2x/DfH+9YWiAy7PZTaXIfYO/cp/6GsZ0/e6YPRFSJo8bEClb16L2VOQ/RTbk/UJ
FgO/TGXLGeRwSm2iT27HMMOWE2vdNJ2boMDlKNMkL1yBgUCARYUgf7QxXEjxEunv
37mKIMAf6kA6hVNmRgB/OlWFzJV+2eFYujN+WjSm2XRKnLbPHKe2Csd8653VpGM3
EB7JwoFAlAYPfJVrefJNYFTHBBl7sLLcwOX+u5xo87NeWlbIr+r8l/0RLSuyBDnb
XNJkGMVwH1aahZwad0pEpuHZCB/raZ0H4nQelNT68lUW0OtdMbMBJRGC2kCN/3VS
116TN/uPOp+hMvjpLOiJkWE/hfe7pD6lUftJdLqZtuJ/5mvdx590AFfbpd9YB2fs
nPa1QWMZvRY3c9uk5IjQmddxHCE9vV6HCJqni9qOC9nn81MJ+T5noMlvIGjeEPCe
/ywoDg+phcZqF8qRfrLLLzNYh9n7YuLZvpDPe2BglEcRIowDtPjcP0Wu6SboM0kw
MZTUBJzaCnomdb0WjecDwWWbHADkY/grvToCNHtaP70104iV8ugSDDSmT1X2cIbv
tDwDTYSAS8xJnNWqKtZ8tsYXc7S8q8x2gNxvHGuEgdLD6P4+YGNAGe+QM44DL+sN
ZUG4C3fsvXJ41kTtdep2j9ObDxYDPb/YzNHlJzugXPGStajIe9gJHpJAtoO7GSwl
79MuNxIr6rx3i0vGRlCJJoXx/cZwULUz6TAXU2JS4ZGfbEQ0tc4UU/w38T/cO3Wq
AVL+DcyP2swBNZqq16bjr4hNx82cgmaLSzemcWrgiwaufQTx6LTJ7Pyeq1MX1gDo
//DzzO0nc+kMUd9Z/0VkbnwI1eJ/KK+o7Q87UKn5yODW4dx1khIhCs4FesDYo2ks
kvaDYUKMfjUyCrpiH+JqmKlkqOVGIotibyu6/wwlJJcUegzBo5GtdJNxU3RXr8Sl
L8GsdkRSYTOHRpofZ9n/6yX/qaZgD+84Tpi/DzfTpi85ongIYeFhBOE1x8JdECsf
rnZGhKDhrtBfjKj7f5d9dXygbgyGBteRyYefRrjaFwxDjjmR4wfI8JYtsGrWQRxZ
+fcLzLIBqJ/cJEhQSVJ7OEnT5gi06d/Jdpvco1KOYB2hucD4fvmipM9aLAZ5JwMf
KiASPKEl+VRu6jFht20pWGr+xeAE85Yqxp7xRhvkSRxJU6eo6R8UWNxYxIV7ht1s
jKvZYQEJSyjPzvjZmQsoUjw+nho5p2q0obOo99Iq/w0DM8QXzTwMMqH5ZwHC1q+8
jFdmJ9ZkEDH5Y2OMGJyvtyoaDYXXDjdo5FfJcGUqCnySZbu3Qjn4stWm+PZ27qqK
cSK6VDbjPEM/OBPmUKvAoQNttysZt54hE0wcXV2XiJh3cVdAsOFVWdIoITaUGdrf
qNzZFjsPhsz8a4pfpSfKg53FkK+kNQy+ExU2J7msRfV+mv7R0NyeZtz9xiqO61lJ
V3l0ZKe5BdfGCqaZzf9dTdb5OACcII2ryNKXm7c06ynsFve7b4a8X99+iO0SlZQz
gE5+WnftfHAJ/OtmFYJCFm+WRu1C3VY/HjQIUMUagEgxPGA6FtJtIAMpuBMPtOKn
QDTGgVQfeZ/6gxmGke9WV8NVdiQQzlssb34gUU9NVVtE9lZV9OKyHltTfOwUa6tJ
Zn6aLAboTPmEOOB7PAfd4ISmhWMgQutZEsjJr66RygfRBNXa97JP9mQ2OxHvERVM
n193rbrvUze1LtkI/kG7h90xJvRP5f3lkUQgCLXfir8gb+rv5qsOu0NNGpHqSQYl
YN3FT8LJ4VWVYEVGpxzi4RBxw4XnAKXLtL/M4cdGJSColwLDqNQuXR05A1tPXoDh
Lb8SPKS400GDy0b9j1Zd/eNy9iqWkkKbvnaApanXU12H96Y5vevh/acedl91aWk5
zFDz3ZKGhNUYMMJc2Kbq+OfVVrv1/ZZLtB28uTSsLiQlf6JhLsHMJZq8+LWVciyW
Qqz0Ku05FJVk3NvbLvg23cDl6UWynLLun/UJmGW9fVIBVeFHM+j0JE5h453H5roS
PXs79C2fqDc5gskrD1z6mkFzHsVz14O6BjaBt0pgf9IpzQ3GF2coHOBL4IichSwn
J5EyX9t90TMiDRfGwfgg1zQRuPC3bLabl8cjXa77ZjaQj1Xmq7FCN5SU6yZkRcrN
+PdPzm0sJvHCqGcG5SmVLXKfTKTeiFTzBozutWNL/b5ddutRq2ynpvjzubYIwOf6
eRq9DsOqjPFjowZ/KMEQk4qg/kDFwZ4uJfvWq2Ug985AE84zFHWLqoPcFxz965Sx
qqCBBPrXxIiHvZLrBN3OH8vQ3zUo4tx568OXDm36tLsxvErYmTyyw+T0TdmtQ7ep
Aqb0souHnYYM+4OaLTp5vuRtonVJCXCKOijId46q+WFtJR8DFbll08la5JmkYbcj
0LS9VD5bYbW+NXUrnMPFy3QgUGHjRXEvB2uaDT+sVxwTt/Pv2eRNtiC+C0GD7jml
8jKOgAJierPRCSVmFHXvDi/IiH7lKzcJla6xlBuKMUSoLBEdHHXAjvKLLljFJY66
KO4LYWwaKXBLzVNffov8dvETzPYKXLiYVi0neM4K6QjW6uJ4n63Eoza5TBrEesYn
JgJm4RDTY1w0OLwX8dsrSqtC/2RaRD8T/vUaCL27cs7NilFL6zleLoZU5jX5Po75
ZdmWRUpb74gNWS06tnKQgvI/EPxscJ2/BRhLx23yWI7Ts26PO9atbpWXfnfxrCyU
NvHYk00o5ZfRD5XZFpK+dTjiwnOPIsvbi2nckrKGL/MDDfBQLh6su6RQqnY/6gId
4LRmRdsKZrkfnMmJPW3BljLIHVSemNuOkpDhUifvHiNKyB5LZH0UOKsrE8Zf15iM
Ch6PKCSapAwPLc1oU1rm0JP5d2KymUW43VDHtB6YgfYUxIhh0So8xSoItL316z1f
JxPaGlWYYVvDSRKSuNT/Uq/15YC4lc2eTim3Sj2GhFbw7AxFhL2Os3CNy79pAbgb
/VHEKlR3UxVUakZMAvaiSEej9gAvrUMJ9bbCDhASeZ3xDZSrjbGa1s59QKn5nXRH
z4oq3Q1yaJM6HShfZdAReDNpcO1EIzkVBBTRlWINR+hST8SigoYGy4+DfUZLmqSW
qKGNkSbDTzv+27bdYuIIt7aBkpL7dL+TRA+5PSLUDAoqV3dKF6LBZGIc1jNM6YrA
sjGDDuh9m88tOeCSVWKDpD6wcmgWPdFYZYDFBIxBh+A321XjYoFM83y+De354n2Y
ezymH6KaiYZPABk7VnClReSZqr8K2xXXQZ3VYvRGLsG+aC0P9RYHsqmZ/IeDZ+wG
XIC6xTwCY/zmyTKdY+s0XR1Ka1LZUuU4oKDWxG1502aTTT+ym4Erhow/rJd1JrfH
2nxNVFSGE5H6JESaA0Gq4SDkv3/+s/pngSCC9k7OMRbyQyw30VkMx7mMD9f30CAD
2h4jFVYkWMU8lw1t2OzhJJPm7PQ6PUPek+QSamlQq8lzfS0SUXExPygnpPiGo9tb
mHrfpbGTtCJuOtdKkVrXEodYTtFqcKzJhZL0kB7zEY93duOeum+yHFnieVOmsocI
e0LyMbPJ+w9UACkvTn/7GT0mtuYyQ5he7BVuYs1MykgwRzroiy0M0BpARDYUmy7J
16sV1UhrlC/rWVwlnN87+B+/7HJqIgmqeMN6pTTpBgBouifDY9V2qAO+Hs+MCq7r
U8aR3kxB1c2KmlyN5qZjVM2URvAjo78LrPTDa53wD5SZH83N8575Z3aRNSH6mTbp
BVj404Jt18pdaGEP8XwF5Vc7pflVGsnPWnIwg8TOw4fJyJr8SLbYE1O3XFxVgy4R
jgBLPpgsCU2Nx56ZrGyxKGJSrWZ8sVJLn4xu/RFYqKlShuFt75z1pkkrtAnX16wU
mOX+lHsEnOmt2+dtv61FMegDwnpg9fhRVyBtZ+KBNUBt0MTXPVqXZFwOIWh2z50y
E6wd6WJ0CMj4pdOUsozQT6Zu5vB+LE6zisxveDV0p7Bw+WW6EXuosG3HmzJ/YSgE
7ax1HTQhfiW1z2eYQY3RK/c/kXBkyvOyfPUsva1yk3D7AdrNcf3VdQH1zq7TktL4
4xzH1L74Wzbk5x4U4Tb4+/PKXG/j4aIlUVh44RyolirFzVO5RRd5CHBc+tb2TWfe
7Pw3sBAD6X35guDh6q6zs/XMON5kC/NwGnK+IfzNfHNFs2REXOTRpi4EpRU1RFAI
vXB2lyDyV+13/zctdPeZoLWAZUDKQpIAbXGTmrWBpJ5+jfxSTrL96MNznJhf4R75
Upv36y4aYXU208LdjMiPjFZusaKXeY/Lk7sgmAmV9rFwGRxnVeXg/P6XW82Lf/Jy
mgtXBjhCm0A+l171k8BHF3jT5uxf5zzyxcAoeSZGOxtXb093yqnwtHN8ttk+PNWu
j5v3piThRkq38nSm7HrDfjXZx2Iv53XOkDv0E8Irp6HsQTq0b2E3wmk6oMczayDU
kbco6FXF4v3hTlNtJ4FIm/xemR507Ib7CIJYt2fsti50b+xvRHOavqp/WF/7UzCX
XYK98HEjVCj6tb02IMpVEYKPQYfhDQGaqbVxi4Ya+UoW/Hk8GycsZLaDw92aKk5l
NmqGyd/PbaL46YueDMhIC8sJBrI6gxm/swwA2z1u3XPDVCVpWeV4gPnx0Qnyqpug
SA8Yu/AHeV/F6uxYTY7O7bbuNYTHrb31v7NlADxHcUcw9jLlAQZNN8raHVGcIhaD
UTtyMtNbxHtR+h4SxrnJpFoz+7wb6vK2VYOemcS5ypxWNnwL1sIsvsrPd0Hnis/v
lgtfA6X5F/+v2Vd4MfPHGWowgmZcvEDtxz1IwSRkETYnlLfilbESgwrR6b49VTv9
4vcomKOS7y1WkNdjWg1UjCTzQcbGXna9raT/Tcbe6nB44GlNovXCgt9rPkouWXhD
b+9SGtrt91tUA2ENbQRiAq473pplpKFLq5LlaxHAB7UPH1pTsXBaNkq3ypOZmPpx
YpUuJEBOAtV9l232Q/nBPOLIvs67XZ6aqS6jCHx5TAh4zzu2TdLDWfhDElAO/Fsd
X+9DjTTV/IbiJEq6YmdNsTOjdKTV/yrgmmSieDKFHuKdhc1ESm/0/kFCTYA/wudL
IjxzvD28Ur53v4f6tTLzUaX39flWkcIClgvQtjTgUmY92D1zP05V6qfmB98g8TnQ
u8K6bGXU5kSNy1cv2DXUr9j0gm7AwfWVf+PU9DAR6NsQRd9ExlcT2LjJ1Q9hqV69
oNhZLj1dinIC1IRyCsPr8+p0uC/QAANXPqU2IaaBybHuQtlN24yGW76UpmNC49t4
qC1io27VQ9zfFXJkC0ffj4SARMvgROH+ijMaqsLoxD1xQ+MNP94fB3IeG1Rtn6cs
o7UI0V8xTUqN8TAe0gSlERrE7AQg/pwLJ0HeMwy1UBVrqLwDhCur35AFl9aQLBeA
FKBV5penc3FBCoSHqi0R7xpyWbCsqF8Bq3hW9BCjX2u4l6SPQp2snU7V3tmJmS9m
CCubbXCN+8xWJkP/vWKrtiWf7YBbbUPiUhBIbHr3lDMBptc55wDLr5t8YEmFnBx5
LOplp508p7PSCDHpadhoojmkqQ3DgoGXKROysOfyKgHn0lSzidzDkZxNL1nC9SzZ
Atuz0isq3QtArFQyxG/wlVLeBio/j8nkxhIAWlmKC8bSiiRyf1oZc3qxYLwICYqd
+AbT98l2KzzUbyiI8YEoj6Tmwgtacs64qMj0ZHPvIUmB6eMTqIaY/GIPzE+uj9IA
OyBNLnTlTRM6JomjkQn+1Ske/0iPVJL9hF7jNIZn4nz+Ljl2eK1Zky5RTeoAPBu1
OZpahhZlSUAOIT9qqapuOObEQ6q2yxf8W9U6Zxpjwy7cPQTfCO/3O4SG9c+zzy7e
GxiugjxL3NWjGkCN/M+MjC8gGoz2TWKmnrpTkC/43P6mX5L6bcnf0eaXw9i0oKga
KL4HohXDS4UfDu9eNOiHt/HJxoqLaO71p5lbPa8VSy52+WP4Onz0j6cZfgZUwbm7
tOViAUND1TtKYG+DUiqtBzZiDVVrJR+AckCXtd7AUuxevojMH41xQtwdYgifU11u
8KvTUw0y/4i4N4GYzhn7FLgXgtgkWYKn7bMu2GUJ8JNsfGtm70OmWPjLRCmRqpOT
87XM8fCqWHD6PqAi7Y/HP5fyUDrW82UBj8nskfvepWUW6FsL2/CkGzDA2Om4YMk3
XwjqQPc33p+eTp0SsqDv1DIkUTGA16aUMikiDT06435qrFLEY4C+I8YCRhmlA4h1
Gea4lzZqxmdQMvOnlsSLGoa0aSubytkvj2/WlFBsQyWhKF8crxjoma7M01y7Q4j/
jR+6t1aYJhq71GrgqzS4RAH+4PNrBMI51K1+v6N0olSG/NQXkRvDyt5dMxZx5Ws5
vloFSB0MQVfpeB9fqz/wX+Qo4DW9s1IMKcJorERXMWBZFNScBbiO0/UO7lVZJDwd
UYBLK10As8AOf2lggq1fjnryUqLObBU4sQIHEnpodpd0m8KwfFgAtpykKuq00DkJ
UEgkdKlrkgNJINW3GTjW8eD2kf0G5qRXXACaQz/kgwDlJkeRYpPnQJHDYHk+QoUb
ytm2k9sqXA3QNiSFXxgWUSnEM9xWfHXV9LbhNYOHPcDT9A3JLpvlOd8KGU56GjRT
Eb15jg1MeZxIqNBXlGEABsuOLKTmnRvr/QvirWBe9kzDWlEQuFOb2qREY7+lMxGc
YWMpSvdJGIZ0Dj0XSIxBz3Ci4pwkoYjAfxKnMf9/hp+wxC7wSOxbggpAohyOZp3J
RZtLvpsU8uBR0nmdi0eGwmrFaS3Lgc/fofsTO3D3nQ5hPSylbx8Ik6iuv4XkQyMe
cgIMS4UDZ76HQpNhNH/2fom8t59g1Lv7b1Lns98FPXURzsPDbCoWYMuU2D/EsA9K
Vvv7p8yHB3newINHB3vbwtD5XmLEmVXAlg2/UBzPfxYcfYdPYdZMvfVBcljPKDp2
zF46Q6U/8xHoRQAgNXiGtvZYfzHX2CguYS8uN7lOcKLzBZpLxKXgnVbJ5vgTf8zp
uv2DWnWj4kbpJwzy8oG9LrGktvq9cZ0D7IirBC9KSiU34Djfr3dL+EYhtQzkW/AZ
aTpfEj0J+hvcDlmRnJJ2VBGT+Ub3GCRuIod8jJAw1d4YWWXkuK/pemb0ImgHmfpx
KH8hbQrNRX3kP6NXNWk+TyVNudKWEV8Ck4h40CZ95yox78n//N3sF7+OPjzQX9m4
8HSC8onigcjw0FAnpk+zPrtRfknGlQatmUy8jsvnyapHOn0pA3mn2zpERIet3Kq/
4YszoByJvgmNv1DeWyrKmI2UKdb2bFmIiAFve+RAEYY5CY8NouZ3f/DQbtoFJS4H
kTTvnykqYOz+3qOrL4MZGQtyXGy7AbhXCbTpM/GvfcSJrCbmxgGfnukGFh9uBz3r
bR21mIYQGZyRR1Tf8mFA29eQa4/xOLfIuLJOoFaAvnYWWwAfmg7Ca+kkjjgrP0LN
YnUYvSTrnjDseGXILd6HBiS9gVjXpwLkRVXpEpvzoRMstuRihJqsgi8MVp08lqlO
/tpfcw6VduNRV9ZLbIxoYIj2me01yrzhV5XRQwobpScBDZrsTXJbBL8OgCypf3te
eknye/ycCVgt4xHTPpf5R6KNJwGERWzxmAPyNkG2WoGYMwtfN8OtrKyCH0TWeNGS
JLRAlPxFjE18cmuc5ZVGRvMloLEn+7Ng9mqbgbxxz3YrRYK6pZQWb6hDjobrRTv1
9TkqTo8hJvM0laDKsr3+hjXnsKktwhD27WtFeBbEZLR4S7LPGaipRjsmnaHKiAib
do8+mQRYZ1lLS7f4dxO5dxW/63SZcMybOCoezzwjwsypsWBBYB4jX4rGzZjc3MT2
YCDx21xFf/Dnt1M1Fd0m0IrCZLiyTHtGgZDmOVCU9kFtqy6fFGOdWbKqofBcYexh
Jz0H+OWtArFlR5NyA3OFkgbsUaqWg7h70TWzWBDpT2b4uy/X3mfQaVfmjzF7vKxQ
9L7qOgtkHKF5YCh64V4uGF4uF3VjE0I2W+gl+NdYuDn1SLuWcZTf3g/6lFnOSx5h
UZ7oUpsfrpD5rB7xiKK7Ci/wqA8WTJwlzs7CY9GbKSwrdEXAsnA2r+xCRdtFphr9
aAHTrKzNT6OEPGGTZ0HSQjkqX8XZm8I/6VG/ftVg62Z0rH3uVpoQCnmTzqk+Bztv
LmV2IvgHyjvtWoujlfgo6VufSRTObYpjM5h9cQX42zw8HK7QiuClNgGPINEhjZIs
sWqFV963hg86Y86HAGoYo2x58ido6oMX2zI59beVPrBJXtwn6ZLSUT3CnCZuZ+c6
p+d2xF301+S+W8Bm0fY/KX6+uK7cSTVjYYGX0rQbsJIdMKEJtOO8eqZghw0RetPw
qyJkkxsvLgsWAUPEnvqV39lRFR8jZIt38WilSSyaFljNm/EOb9gLZGca+JY5Asf5
DFxI4x9cBvyiGbW63JSgHDWLRF4yOu1YVZoN92AJlEehH7T8njyuP/VzYqR5VdMQ
JrcNH2tAxy/+F40DVWakKvDsunn7BkWxwJYHl+0bq5FiFZPcw4P5gKsneoI6ob05
9JjldffR14Peetw7AbHKHtShHTPzwvc0lyzgDVgAB7aiAd3giKNwRieMlHjk/Bgr
Py72hAyinX9zkQXW0oNepXT4NpCoel+fIsNCFo3oWwP3erUj7OdY4orBlRZYX9on
hOy/YLCM2JeCVNa7uh6t5ZW2UDeOGBEmZsaAD6i1HJbX4vreGlIE/yOJgypFhJ+a
Ck0ZqdVJq8KOnU8Ruv+qkoIw593z2NF2V3dScRd/iwIF0Z9SjOjRwrEW4Svq4BsZ
OYmeHZAj8zHdD1Ylfyk3BIIQrJdlFtsxVLjQFJbjbbpQGH6jXB8mJIWLc/pyJPk6
T+Ge+TN9fRpsKZx1qbl507zDHibEmUrWRvAvneH2WHqU/1Mb8waYzoO06dE6q4dP
XV7IubwMFeUGEsw4IgafbnsuJGrnq+zuZIyWSliCMRNgAX5pykyaiRWcTyTczKCb
R+7NTX3ODYuodeODXBX+Skhjf8+zma/NXNRfiR6qW+Al2f26dc/TRFuYqg5LkrPm
CRDHL9oBHnYu8NJSs18IHsxWCzDoZM2auWDJMPGo7m+GMAaTfieEDcm92sHgV0OR
Hg/bjzqReQgaCQUt/qyz60JSV199gF5ydNocceCxgqndqbS0H3v6YlXeCWnaN7nE
IKEVwjfCXXZoQRli0o+siPgKPZt0tj1u3/ZdXguYeGmzmmIiXiL54wxOpMmaJ0ld
x3YvszQ+ZlYhNVtUQYAxTwr5PlMN8OL5GT6e922d+vKt1MOR/nEwyd1Dg3GpnqzQ
+KskEBIaW+MjinPFgZ/LlKJR4wZO2QNKhpHlcFDVhQ1I8cBpHpZ6iXws8XQvbhez
lqZQaF2/koQOQmUQVUYswoO9gTJiA+Qdb+2+FrXPZdq3584uNn3pshzE624XVGfC
kj7cHGyi9dxbytf/NbgiuZsTMq5gqVMId6awlyWi/EPe0oN3f7YlOVmthmKHVEeQ
PC+S71WqI/xTJeS1GAiAOMP1CBcGct36V3oL4cNltZ7VDigQddDX9H2ApqdDG4Dk
ieq19LHZlFNpaux5rYqyI2fxeEWfbAAUmGb+BEC2x4Qnhn4S0v/iSuPqoCctQWIY
BS3VsHnRmSentqiT3zFkJ26JiD9aThLZoah0rW2Nx3QoYMVdRnBSnRNfW5b4Vh9T
lzlCcIE5kWPIGOValwoP43R7S5N1vY5+WkywlRCd/B63OQNrx+nsMVSExQOhEkGn
ExWeHy/ISUTg43otw4TuHip83FgyMw85n+0hKzF3xzVSe0wa8U9rJ+0ObmP3jecT
eoe7HeOGM3zZm7ZxE+pc0X5g/ogDi3RcZNLxkyvxxegQYZox+ACaQ1XpGlOwTD6r
X7nkYtZf+ShnYH6wb6KFUPcFkznWt2tpXe9zd2glaWcEmoWLIX1x79dO8x1KB08h
di2qS/AaPtvnz4H4aBHk8oibqvsKKM0Rc1EYCxP8ry6tI+YeRRYmOh3R27TQQ7p+
x6uGL1yFcKaRX7DuUuenmg9Lk1ivQLQQdy5EQFKMXEddX3aGpDvI/dl3+Bvukt6v
JfWPuWMVIKJhRHTveUv2GNtV2w9/tlqmvgeJc9/YuMYhCO0do8xec/y+6pHa2+3G
+jmbr+IxNiJdsJjKsDSxd5O6mp2inFOXfxR3TJXNOlYfvSYiwhz9THnpMjfyXLoL
yoJWaezr729X0LVngiFx/iU0mJyncqxO+1c27XqpSaGnr3HJv/juslO3Wh4+6saj
vPgCS9bYSM8NjQNf4hzfYB9VBlkGtZ3WedXO30jb0XIPFl1j6dREAU+I713ZAXdY
pH408YfD16fRf9fnKQnpRSGJcpeTnKReSZN7fyx1ZFSgjTx9i622z0viXxpxEXLK
dfIlGxEDbmABPLHf+4QQ4C2iZiAaX6UTIu0XkTB82JLIwzi1Ji56GKpjaw6E33nh
vx/zWlQTWMWjTMGjcZsdc21QNJ2s7R6I3VODxHI/4RDbKS71p3BtRZIZ1gX00i+I
txAb+OAtKmLEO5kXad1hDInNeQASMsEB/zxSz6XGzXOXkzdKB6W7l2eTYuKiw1pn
GarNu3gXTu1T+lwVPPP6+4NVi3l/9l4/ocXMj0xm5/kSh6W7r5dDbblvouVadB4u
ShEeDsrVGaD/fiy1H2bAy+4mRa0JO6a1HoqPHWkYYV5VhcOvKCr5+LImM7IBN+2j
TgBMH1NNGlA7LA8UGXAp2NoHyYcoS9+npUsmD4Zj2/1wli1H92RDk/A6Aed6KtwH
V8E4hwyU7oSj6J678STdu5Pg1zoVEt/3vOcR1fXE1FwRVzt+Tq8gcJFQhDB1RKYK
/KC4K64hAIG7bIjLKWUvX6j0U5AMCAA+jDllHK7bUF7quANVsuQq1UEBNKAe06bL
36/96rWdziycooCIMHYyXB5dWSFC6az9dU9pLqB/GYudsgnMdX/HtRpv2GBQBCc1
eEwvX6PQMRPimIriBoiPE3xZwIfVDHsnGxXcEE/SuJXecUxlmWBNMMiAHJx9N6AI
NaJOHwQGnfr8GRH2pG4csg/BDdnpE8NmJ/rgswdueSIpYQBXE9bX04EaHgPxZcR3
CINYuP4oNj98ZkNhgp11vUKBcnflbJRphTBvCVi6PbRGcf96SiMME38itSPXzuR/
FHMZ5hFKkpgAYz81+Uga+zmHtDYvB6mgDnGiYlZe9BYtzGhEHy9N1EhFSB1s5j5e
lNW5UwJg2FAJsm+r373Xf2gU8TKnV85VdQ6e+76RtgF4fFN+uCfF3/W0EWcAqaiH
5zA0xw27kImyxIxeEt3+qoA6f73v4Bi2I9JyBr6B8OXCcbT6c81+X2/EJUjzuSNF
7Uieh9kkHyfZm+ET7SCsbQXXwucuhlHA1dlC1E/bfuAic/pQa1/aOI4l+CxOZukW
MKb1+geOxerP4aNDB2I/cSKVy/otwYb9GOqcMtyhmLP39bd4rwNxXMLhju6onnHd
nvQwhNcH9c8zI1gR8h1ntuZm8wOIPaO3FTH2baUYwcVqC6oKJAxnN1v4ggwzl77F
IOgjjG2mOeFHgh0dFY076ftIYddXG5ZQY4CtGNfhAGNrriGKpbayFXno3t302GeR
M7Fnen/g0WKa2ruGL6VNaWtZdpRF0QUnJza2gtihSSIqh9mqF1dMczDM2Jiywc2o
QLMCTaFL7ZeGjFaDpCAnWYadRmfNfpGCVYeq5/UyF5/vDk3QmFxn9JVauyAQqF/1
8lHOeCHkcmJM8TRdVnz5Rmr7tQymGzz1x1Qw8iQ0OU6KUl0n3m8zEWqwEP++PhMS
n31wPywrpr1zvonqeZehuuxp8+eyWC08GIqNv6Evp2XoP9Xf6E9ybcqFd3asyEuV
KZ7n8fA3YR7Ex4SzVdm0pMGq3tpliwTDWmAV3hn5v0d2CUzgF5Ltz4RsvvAnhQvi
bPb9/OCTCCcUpMkRmu4/1zzwmq/zKcpRQvvUVvRPKENi5QZMNGmkQhG84JCv1sWs
BuIVoY6RG/y0k0w0jwxrgCozWG1S+ys07dB4frTZqArC60mE5TCZCO2/V4IzEqjN
jEr//Ycz7jf6AgyCgchshIYRYJpOWMutO/OaPenRDEX3hQYbSjEHIGGwTVKXRRVo
dhWmfkiLEkzOhovSHLQawoCNmEKaw2uRwQ9dSZ+qtxeAE/TxElY9VqcTa6ERwKcG
fWv/slXs9CqcVi1cjEwegkY1/d/otPI5IxQKjBGripnf9zX1pdHvPUs1Ba7K9LER
bbtMU3ZcKIYlX0+cGnlVyMev70nzi5B5ZemYzfLDGCqp3Af9Mr1EykIoGCOg7SBL
Lb4otZftEKe9+7h7CTZHErggtV845jzunFE+gLGv0ZrPHPXbrdEd563wPwBlW9lZ
yAnXg79qr5mPmFCS93DGQzmRkyyVF7VuaGgauSDpZWeXcrb9pK8qfe7YQYzoJUDi
V3DkG6vOuO3Pw14rDDFcqhon+ObkRyQ/dOo+gL+w185oqIuQZ6FDlZc250qlr1it
hjRR9aszpBc1qCFKQl3JosEM/Llrnfuand0cE1Tn5F/+mJoV/zcI7s9ID4v74GAx
0/okzF8TTPxTs93Uw8H02uhTzxUjbuBlzQM5F2miEruJsmxGz+lst4po8KgcZz0/
jRYNQ8wIPRecKm7xHyD61SA0NytgYeRi0Woq/9QGksxdWlNRZFaaoyjCqvB7sWCs
PrZ6zN+VjU0+67Abvon85VUdSDvjFIFcc601gLXwhSAXIUnIXzFLmVkNQmqPJt7m
qJR432nJZOc3+k4JXaiTj1Pv3AdRn6+M0+XkR+mlfJqVnMGnWDGVjZF8T7QdL86a
x1eJm+r29KDOGDwRKzKZ2X85d9Q2+fEw7PO90VfyZFER6ASZQowfrd/IlQkuuuVl
p6HcExiIs7I7RWqPDr8RDGwXOdh61hps0nksX3d6Idax+bos/N/ptPLUEUJAFU+C
d1UcbD2vDssu7elea+XSnEnkA75mJKN+oh2nvNIYh5OY84hFr285blcrxwds8j/k
vqEhymOJB6Cj0OxzMqfTuG3ImjrnPAy4sQnWfsmgXJlg7YA2oMpdtAQv9ix1WF6W
HmDJjsAprBqsZ5Py9Tbioy0OSW1Sv1K5t7KsdUylGM9eNUO/g6JTqFdD2xddsAEA
O3E2wLdfRrFeBjkzdFvA97DrWqIeCKckjfATw6dEPUcK9ZVJbj6XC75Y9u4aiRUi
rSHqUOEdc7jnwHfj3pXkpC4eeHvgByFFK81rlGihOdbViph5g0pjHUUEKFQV0z24
oujxwC+41ptUKe9/mwSJKtVBbmLEzt6lq+gzk7qxmseCWpEuf+eVMABgx/nHTHFg
KtjEA5ZaMQN0dEWiTAU72X73E/lqnY4x42RbFv49vp9pEEj+bF9hYQVqKuU/j2dH
sSEPcFLPdxKzftAIttUh8zQ2NX3QerD8Pekur4LetA9mfheSx1XskcGe4LqOqg4m
XAkSs4eOPBn0NQ4aOj9ax+xhwwT+sT91M7GpXd/+1RFq/kKMMe38xn5eNJCgTgz7
o9DoO9EuVq820Nve3N+o4FS08GNuKLpn84xCPDiumrb5MWHvtLiLnzNtqQG+Sf8+
hs7BNgaV4yBMz3OxObMM1uD0KogNl2MsWG6KL2cS/UvIacg1BJ8sNT8nsZCjU/FL
L0Zg+6GG2rdjeC1ULtCgEnmb+KJNIe4esemgCmDQY+BYO8OsDaYGTrS/BVNzFaJu
eRDTttXfJ54suAfohICQyeISdORPvdhdffj6sqVT6ufDTVouvg/guVLWnZ7FjElH
jzafHpFob0N4a4biaUYnmkyK38qTBLqe+InhBrHMbaPn58EaOYh68iy4uRmLZYJX
iSFs38zvaM/CqbKh1Cmc9SIAz78jciGu59+FPw4lxs7XsvabYvymG9vedewrsIFs
GdSrzZ/SSvbOGmG2oPrCYZGsldhQVz0A5Z8NOISn+QZIvcaC1F+hUE2lJ1IrB1Gw
Ibz8wiP0wX37WwYJ8hRkskSV5QH+RMZRulyoqo9LvzB1zmDKQn5Ki/uVIIoQ/4XS
Mz37rtIl0pOWU3gmUPo0TNR+YiLaPRLqKp0JaqcpUiKAZ1DwmQL/qxFxyqcdmrSb
38OPEMF32cZRBhauXLjq3de0B+weHoT9474vCvqJZ1bpaP3RHO/jst7cottF/f+M
La2NvEX5wkDOzsyu6WUbKvuClbfWQHbqH7wYtOoq9B8+3idtIv1lv07ZNkYZNpmm
Y9wdNLARgWjSA6xJnCJcKp9Zq8XM7uRuxJ+kj9BbUt2NmsLzmjiwVV1zIW0gM71B
nR7jB6zjOrcCtHshF0nct6GcACLflYwPcCZUb71ogZ1RuRNib6JsIyK0eE+aBfRE
xky86sJ6Flud8LOJdQ26wWsV6bTQsNXXPQWaGSJ5regEZNclzuek0cvTYRCK06Qv
ztTK4XX60bGsJ730J6p647+8oszOZI8C2MLgNSynIOwNRUnKxfk6h1n3+YDpW+dX
lUmhq5Xu8g1kVu8VncrhRri00w+fWUEYs5p/0m2f0Av8ET+A2FNB2GBHHU+y/AUo
UXfhctn4ajs1pPeZT/mrfP8FzKbxPWG5Nvfe6XLTtjslgB3/OBX6hEJdx7+mceRW
ZVH3sfqqDAcSJbsLoV1C4/YBzDe9yDj1PIgjEk+kapG3xrMASoaBDOgEE3sXYxAt
BE7MiKbbSEDBP9oRcZA5d8k6aFShkpsklktvHrH7p2wEDHPgapYrL18CHwPaESk9
ABT3gDJp/2dThHkJH5IMl0tpKi2i9UkSK01Q09hfIjncIo/MhRt8xOTWZoaaLAvI
Z9EAEQTgwcJmb+7Z0MGQNS7cCicQhoOfy8PsxLo2qRH3vBnWSrqOr4lLK2nSvkIl
WEj599yvHHDIQVtMxp//ggbkkHi6wRFo53r7f0YY2cH3yPP08gf7+kRgUr4hwW60
pNbtQ34Y4ysFG+m0e3Qzn/X1nXR4VhLPSceAtMbFPh1J15N7HK7Y12OqIvNiGF8l
eUxx8en3xDHTICmb0tpA0O1wUb2qhu5FXYE4Hq7hkz/nZVniOG8whpTuAsarK3E3
ZlUDf7QHiItXDvTgAWplKa3ZPbovY3AF5FMjJQT0YoiGitUjd3S0c5NFK6gkbsPH
kmcJwuPjUkxN3KJ3quUa1BqE/hu0ZmvonV9LSmvyuYQOZoErkbBDjKzT89KvURQR
XIbMQdo/T93BosNKXOWBrBmffaRfwYSrzFhHjAf2qagoZgkVmaSQ6ogGNbPl5SF/
NgwuCU7OEcP7GP3oTJ7OKCQo294lc0kdKNamIzf6iGutjvJBGfvI0ILBXf/RRe2x
G00igms8vWhtXkc6Dqd4HZh8+jz+BvET/4MMXzjnemlpxjROuprdVUlZFcMB/NY0
jlKyoxMZQLeYhT8s6dIzOPYWQmCSeIReUy2Z748lvTQDRpjWoewSkNu8YbPU+lOm
FDzMl2W1PFIIUK9SP36mz279wOOEcgCz2otDdYhlBv/ETCxIAbYqeHJQhyKt5acy
L9ad3xhTHbyXZd497I6JYCvyewU11YR4HsC9d2FC0Q0SNVB9Dg447Z4Je/cjbivc
45OX7METynH4AJdb8zHflnh13hVcH/onyMaiItanjh4rgA9CqE3qkp3ibxtRdqfj
BsZlIsiVaGIIv6vhj5IcbenhlE/lhQaSJxlvBzBMpzqceRUUCf21nMoknbleJc4Z
R8/sdBZSmuxa2qb90VBKHe8lyV2tTnb4W3W7ox1QWu9WTRUApeuvnXB7gnpIiDMC
k7eQG/QKnvbca93Lu/NDTspbhO9NBVK0GAWd3VB9/5PwCbkP4+f9eKtggoeYFn/u
ac3bME61+r/GaBkDAF2MeuKxK7JGBD/Nq6Ko/Md9KEDDkUQDzJ05UTUyopMpXfWZ
HFENPjXlbXLjIMrlxqHlnZVN6o+MNm+FIUE3gPBwn/UiR3z4Z4Xt3D3edQSmo0TX
EwAJmwLv98nNym85vHaqbd9N9UUC4ZYchIG1Uf7x4VAODMBFIZUTvB52Ck2m4zA/
R2e0zELNrpZssIHQpJtoWM7T/2MxS6v0IdymCA8yA1VyfRyI9QSnN09fm3V8/dgC
5/cfDxIHgA0DfJOf6PRBoOpx0nQdo+ovim6kz0+LkGomnDSQkgAOS3HVm3pJkTPl
ZfOpBtLmco4ZGH1YjtP+JhIcqSUz2Xg3Am4RwGqTZ9y2PWiV5d3zRW3yx6vAJ94s
VL7GeU2Iyi4BX/tSQld1MOsS6UdodOBVravWBiMa8fgxC3IGJQpRrIIRto+VNDXw
vKco7CAi6VVbCOQXFsYCTZcJqgpD93L7M+QqtC66x0ao6I1qsutau4K7Fhz06tlu
kUZrmbGT4vbpbDGAefa3GVsE9FZRZYpCbgaecd3fBRQDUIvb/8LIw/v3MB/IU2oZ
41bB8zDPVbxjtKZwT77/jSC/yPDkkqW7VtMp8p7RVZEZlNLo85j4K6S+GVDyKfMn
IwEZ6mcmsXyAKmHVdKOxFezRjBMcGWzbwix0xkBcCkaer06+ycEUZea3UoiOyvra
aVIffTBEghNzJIXRBJiK9hGzecxyrPbnCxvZSoisr26+eT23T8dXSY6+mHcQ+rip
S4/gJyIJ1IGLd//F3ENM7nXnQszE+KE6SA/k7l0nrXHlxJRIYdVgKWPOmbCAliRv
Cvw/6i6dL3dheU541I+DPDMXOk4ozG0Ntp1rAj1xh2X1YLSP1Ol14rveO0e/PVB4
GcNYlZXFO0bP5lcTAHa0OzZwmBXIvOCZFoHWGcIEXXwj4fuxIRXNeRiJq7EbJsEE
TIXE1kPpidYxdr4mu5jyMhlALpoTxGj0LylsZU7WwG8+frAZ4Pm371kzQeEzHRNi
5CD6J2SfHXWSF/Xd3WLogrA/JDdKgv/1mVAwA0g/bycCZ+RxEqByJ3uo402yitdr
1jDZQ4vqvAdBc6VTEHEDdWH4Lh22qKrTtwTC9Zk8ev59baqgANRdMuLiYjp0HSx9
eLFlDuoPgSo7yobNPGk4JjwnEYe5TytavmHEviRKm1MXIhW1w/1udrWlX0ndK6ju
7w4i8KDrLirC9nZ/G1kpvnU3gBQ4sGgp7+SaP3Bp8NFTr0s1zFTjlBYvJR/NTLT+
x7wlSJ8e4wYjEVzaY0jaOPUebSRiQFTkQdQAQZXi81BMvJmrWw3jMzDxvV0Tcsk7
tvu5wBeP2z3VURXGtrnfIdqYzdpE4RHJ5xr60E23WLa5yL7y8SAWh2jvIYL7mFwp
d5LlRPadRUnsdkQW/fNg67x7vdwvlBCYhk9Q0wlzrMwlcCOlLH44Wfk2RK0mefwR
UQrGzg/ReLn5v76n19syvCLmicNzk3j/y984vrCvC+QFd9V6Zsq+T4ZWCATBFNA1
XjUE+mCxBK9Bz7+PyGUj3ROo8/jKQDLUwrmi1TfdDzIGJVuaI9X7iuzRSBqQMFFs
29Meo6pGBR0CyF4vHt9Ym9bYL8NuU/vZ2XnnGEikPDjYIv0bK4vpZQ8VS+MKh4Dp
dULFKKuAFsBbU32VQQYs8SfGfn0G2+JFHMa7EetpjGmvNsQ89IIz+K50OXHdrYUJ
ePOho2jy4pfgWRuREDYJfrvSEK99aMyny+oqBzAr5Fe9dMFH6zAExUHW2HSk95Av
n2B4Eu7enk+qF7Y8Tf9/h3lV5CgyyNAbPOGMITqOVi3XABvKuQhw0OBpNsbsja1S
0p3ITh1IYCf9rPAQvk2hJYReoRUqWvRG0O714Cxc4O6fFh0/f4+zHkyBM01kzAE3
YscReOsX5M/dSlcUSYh8yFf4NKLZB/HFfMebE1eesD25sYY9LAHnnzLxXadRkBsS
4T8xSZHhwkhzX/rC9xB7inFUWURNKQSO5+8lCSPCfU7s6J47/kkg8S+1JTTUTxEx
gm2Pkmk1RXJkZm5iKXNLNPr9fcM/p+eJOCq2hi55DP9O8vqcT2ZmD+m/8hzbB1/P
ahEmcwNvVTxwkIuY/v6x8K1MfqCWGCGVkFWXtvzbhlFwCBPJNFVptpKkk7KoyWrI
LpqOXpm0YT5S73tU0sr/W8P4TbGBwhm4C4L0s6mjeNyeKqeH4l4nclp2ClHSC14h
Wi5iBExXx36PLBRkrMtZpdDnxs12AUXOqA6QYBREFDIpjQ3yI/5Ij2gg3yjlPJtf
vCu1gy2OaRMdRfDNkbEf4ZP49Q5P1wfxmg1QpQhHQV8W8xLx/5Od6QqPivgd81EM
uXMxsL3AK5hwbQQnPI+xhpxtH9iFiqSB6p6LHhoOHHcAfFFY3I+77kej9SMDWcId
8hAmnpfT1GGsTGif6Os3ZrKdqPhY0gMMFl2HV/pP1VNTroZdUGpon3IPaVIanDgJ
iWYairJ9/YaRbBTvsZWRsb39JIHBm0ICSYZd+AfBN9JZxRahUeOIBv1YMMO0GXl7
sxuUCWEwkWgzypqiRu70UyiSXJ5C9d3xJyYa9mandzOApYkvv1xbNEamehUq2cfH
HgmvRBRrBT/rYacfhQ3Q8VSkwW5sdl+ME146YV+Pkkgjs6GOeLmNP86L6Cjvb1Uk
mbKEWQhK1q49BZmsJS3BIu40FS1g485BbXqcfJvehwY3CcZP54FNp+PU1QVtGimM
L820xCbrnLLQl6Op4kWyiU6AgpRwrHc2+zAAlq2ENviBC0VfEhMkODNS63sEJ5w6
ps/236KOXGTAdW12f2ptB6XQ0DU/N2ztJfcpVJn+Nwdw6EI8Px0YepK4RBStftdC
izUQ5MAP4bKwDX8W2vFMz5M8r8j3rt0n4jmlhisbXmBMgijPw7PAFQChIjqcJw3G
w1CX6ACpm9w0vZTOLtwOrXoDMfa6HrTfmvhHGtaYy/ZTLfkqKreomTT/lK1HhrQf
mEGjkyKR76xYa0wm50TBlUs8bMjlPebCd6wJcjo1whrKFAdN2YWE9alZOJuf3cRp
QACsx7pS523NXrWtK1iDmxx2zMrUnIDdxe94N9pdy8zWzr1+O4SVCcn+kru33GDc
WCkBxLTsTRNFVZ91hyEYzaMptk6WC8imJs3aJsm+H+zK+HfFBbxS+9oPH2vOcFX/
gcgikliosDvaiFI5zHH7dRvKQ1BcguB3LEG5KWfm8ZuEfbEGHWea1eRgDeDCmwbU
8LKkyMr3ofcVmWdCb4cctQEkqowiSNYkzn9WfXgkmG6vmX2MmKVjnF6N8vlJYU/y
nmVqiDjg8IAHI9FLr3alq3ZRPJ1+DwadNHs1gZUrrTAtMd/ZXaJFf9q3AKuyFUlL
lEklOHGV47nupWnuaUEpMO7P/8tzthz+GLmzrzEvGqsc5/JNQANsyHv4R5uomfWG
eUpMLETuCHw1Iq7tvxAtFVKhhhWYgDtn3J6GWO7EE/1lzX2lKuesleq8iOHK6IcM
TjPohr0TC42l+DK+WNnDlvnWPbQCnZrGJtyGXH+Ua8Co2ksf7EaZ7QKS0cMQMhUM
1G5fSqHZNiWJzVp0W4jkbL+WWBIlaK0U+MPWsaWDSPqLQ+KXamBkYz1P8mc+nhYq
U1MdI6jJxwxgdll1jURZXlsAy6rZ9T5F5WWF48Bvrz8bAP9hqlkJTSmb7vG/1mbQ
rM95sqtjdslWX1c3QlEGLnzxC7dVnFh5lU87U86b2ZzwPTu9ELZOeaDrhyNJPau6
EOwFT025IwNSiQfPFN4T4yx+PAq93p1uhuQYyUiKD8eJbyw7MEyb2QoXZp67oHu+
vHfjeh6hDcLX4DHBkg6vUKF8a1HYgix0Ds+xCGOBfJiYgeR1xPi8KyxI6k1ZsMZr
1eVlH3lSmKsrehE93TcFtkeGAazv+zxEa2v/1w4IxPPCMj/iVvM7/6ldsViLGov1
SG4B9N5oryttG/uHTyM2VWMnbVx1fFfz+f6VY3TJVk12Srtu60lrpCDrjT5i6mgo
fckxBCLOHcnkYp2JXWK1r1nUrEMEuVqPqZmMWS1+De06p7+L61ncnF3rP8xtMl9y
G/VS//QQGnN0QG4p4d6dKrV+ot6PLJGllePqMQEXVc7MU9j5mFaGYSR3yJP+ap+V
d477ULU4keZTVJ5aM58j5p0170nx4yimeGS5N5e4VERZzSvemd+KoEEnuvI2wF4B
S2lcTj3pUXnlwujP1hZk2Kwkju5sZz8CAo4sIC3iiHllml24RaFckr0mUv86X6NP
9M8alyvZK0lwRRO/mxxL+8Wsy+o3p9hFx/mVjRGjgv0o2E81Uhua2H6RyOrG5Nm8
lkqz4HbkVTzBMH08yxdDY1eN7eCd+XLx4h7qrDOQwC/Y95I6iTgUa/5Dm9oSfjc/
n3nm9cK9pu5xPJaMrJouhgOtGO2zbPRbHyFnPKYyIhLvbE7uMU/LbZ+U927Qzau9
E+iQ55nfVXWxQdKTJx1tJyg6asIVtX7raLWrDkfXeHg2wZr5+OG75L7AhSwe+u3B
Zl2zOPxCiGVewa+0ZuG1oxZ3afCf7FYKrYC+DS/Wbnhi6V5np2rgpW+SIcLuOaqr
ypDo1s0IdFP7hI8ftIK6A6jdmSDmnfZp4/iFOrfg8m3qlrVbb5MYHqHom1NkN9sA
IPH8w7dl/y0UMnsBlad5+JHANjcE+kUDJX/RXeJDshTxVuaP48OiQR/cHCg9NRgV
oohQ41oaCGOvjzn9Ls94vnVzal0wb2kAQHn1jz5WMztFRmJZNxUdIF4X+Xy+opWM
wzJG/mCjsqRGWZ3l+/w71EJtRMOscI/ibJYevNYng7lbbqXB7Y9c1hxgwTLk+vIA
XGBMKJkMIKDRhClEqpYII/kbJSy6YYj/qyr54OisZEdtqIVMHfxxbGM6CJNXLpJa
tVVbFnFN1LUGkKUPs+CU5YVjXbZFavOG+Sinl0iYKHaMk8w4I98F7Gxiy0XjA9s+
KnbAq2/HuCuekuZXjDTTaGnzF8qY+IOFVXU9MVZ98V9OYHpORa7HP0gR65TMeolM
DHbUbqhV6irK20po+DPpXKwDUtHXpEmlDehRxXCtpZQOWvu58HBy916+DvDNiuZI
c6+ohTInD1bCjJFlgsjKIweoacWFtu7qu2m2JoLvIXopHWN9UR+6ml27fZ/Go5Ps
MUilfXxjSUAFT8E+bAH5hyRW5OKPnDgxyNClr1mvuIg1OBPiac+GK+ZvGVO8tsQO
hGDFMhHcpNKK8Go3kMh4rQ==
`protect END_PROTECTED
