`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zjberxJTiAuIsPfMdjE8ZIEWBxuXjHyh5x4YhUAlQRIlM2Dp+1LFii4+BaQhixMJ
N6rBOGZ0mHkVEget18egXmyG54T0f+snNwXT54ev9zbWfTAGxIG/D0PLRFn06aQa
L6RfsBvOzGWAqMrtnk887IfCvlrYCZMiBgOtf2LqRHY4L7UlaFIwoKMt/NqgKF5D
L+HJxWp+OHnOdzQ0aEYVHH6tqVYg/u+yV0aNixtnAL5hZsVXXbEPV6Wg3s46xGL0
LFJkoE11gT+9UaQ+lmTdS20wUpliL6rLlrTQ5gMBTANzNl26X4JAwBnJqoR5GfY1
1O7IM5Kit3afJu/+0q/o40/AIiVp9Yk3sv6yGuEGhb6bLKQs2NDsnuQDugOhR4UN
HI8deJoOyHC0Dv9yL/L5H+IvNeRLK1YXPUeWhqe+OD2dBaM9HoGtJyMf0YW6XjWz
Ls188KVuelonK9hXEguMkLnvT8FayJ1aQvGMYhAtVYj81ucG16hxpV8oL8wmvzcD
u5Mrr8cnkdooWfu3JD7dxmNGDFRTgDJLECXcMQ8jpy9zYp+ka1rQ6YD1O7AoLlLg
tOA/EHAxOSaQTr1IN+osvUVr/GgM364AMoSo3QcEdkzzbRoaVwr3OBKbJkwUpe4J
+d3LxZkbFsjJjxz/2q3aFQ==
`protect END_PROTECTED
