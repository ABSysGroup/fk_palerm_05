`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gef/xBwdEaCFpYpCURG3MlBfPhZiRx1eYdP+dA8SBcEy0nuIlmSrFSX/vIKXPGZP
3BvbN/aY9FlWtUxOKxivB4ytEf//XGeOywcH0YcyolBgLD0p9sYmqodqtJ1Kj0yb
ymOw9FsDRLnFBfq9EBCRDmmQKkc4h1/isxyFjFVCGMrtHeU/ujjjzFl7JpHD30I+
2Dgtik8i0S83fTMXGEl3DJYTmPWIasYtisYnCBJRd3qgFCmdc13mZJ/fN1ATIrSO
zQAV0zOlENVPZ0k0YRIptw==
`protect END_PROTECTED
