`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cCE1bZMBDBo2p1z+v7ARvUrrB4D1nZ0ai3t8krCV72EnsxNceCQPJruXkKMYXZR6
+cKK9SMjpxZmdZ5SNtWvU3VNJxfq1cw0vGbjl0aWo5hStexdaoZAzV8kPCgrVyYH
5PF0gndrBPX9nygqD1M3EdNzOFBxxF6VkyRIidvEF8KMz5oHUO+oNX2WOzEvB+6Q
UK+Lmg96znswrhNKEgfk21TRdbBkwDpLyFCaiETPzu2bdW6Jv3K+JbmHHX+Za/kf
aVbCpl7xsy5dlaJUmyhiCpW4EysOxLcfN+oLF3LAlAc=
`protect END_PROTECTED
