`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6n3hD1BgZnlR5JDkbHbLc2ZRyO/w7jGg1G2G5309lNRUu+/G+EhP3BuzgH1+sia1
fkiQr1AScf9OAuh2Difx2IqWbE+Yu0liWwmcBIUA4OLizi82LSxwMJfV95vOJ1A9
+OEEosJoy+EafStSBS8oV4Ahpwjs8lNPvejlPjHQLpvoeL6l03xuOz0I2QaZSSqe
+1c9TJI5vzxWA+B8aHrZJMffzBwmIreqUltMbitGXRaOVlhlcvD1/ITpk7fTX8Vx
E4jQ/V74yzH8QGKTymvY2bDUjg5FQL4m886lBywO9dcOJVR9BRCV27sZt15updaU
wOAPfbSoABvcLiuI9adgVkiI3En0bxcMnqdx5lo+7XvrzNzO/kEzvEuavkTWVoKT
9VhkJiFVroXSNDKCnG9ubx+c5TbaCH+ss3qA8IbTQLc6fLN0aPJ8epdj2w6wVoAE
zrtFwJ8ZZsjY5DLm5hk8+SlJ430bUeiOtsC1IacyQiW7MrgrQzEjJmgx3sTD1hIP
vN5lw3B12UoMbzD8uGuxYdE3xU2z5mnR9X1/OOgHFgt1x81yeCGmO0zRZF2JV5ts
pu49yKtuNM/9Fskh3yEwygrlJdvqKox4eQH+2gSvL9CCNZh9T7q//FHm4WN8gLRS
j1Ed76hu9vVV1uil18VrOHZ65JOx6UXRJiqZzK584SWNCcyIYkI2X7t/2XqqFDTQ
16xCaEI8BHTslqFKq+yqorcwfJS0XF+AWOwEX/yFjRIhzFINiIckOfmwtZdR2c4l
EF7SyXtfrWsA2UQ8qCNr02qMS99ps/5mLRiimRJ74LxH5oAf+Sfcotkl7Upx+arQ
+boI8VaF8BXuK25p3V4Q97vBLeZUPlzvWWvANFoQ9pc8ChAd3tvWkJt8f0TRu1Fv
2ytWW2Aau+dPI8LwPstznwEB2KD35KcqvXBpYALWH+2nofjn84YGMY5YUfi/KqKz
pKWSX0pZJnjIm1ZT9cN/spQ6U75txDyTJM3nHfu6f5FPBov2fSmxI3rn/LET7Pda
5MMST3SDX+Xl9HXm09g7SMGO/4qfNhI8I2TGuPvcRNr1mOtfAb/bLVnmm0qR6cSf
6ZqbjkLMovkFOUa5D8WW378JfL0SvGlwPHyzMz4yXPm/zDP/xhBADJhu9G1bjkiM
WBwMQb6AsB7OJusZndWFQNw7TEquPC9/HR5l5Wi9qJuu9Tz+O9NqdMcF7JvI1RJ9
ldfjH+mJneYDknN4m0Dg6uA037uIDCUjPH5Yl6gQOR54m51mIQ0mwu3Z3U80CQmE
v1o67BrlK8qHG9jywEVfUcFRw35o5xzVFK0spDXO+Aq8J7+a/ejE6GKZ+ClgYsBk
161eAcQG9oR1YoxNVJqYtHoehR1sJ2yvdItFv3pJj8Rsro67j9sta8CPGuS74azi
lanFgRKD9umSdwWaSXbxCBMS6tt4tBLQ/8cSNX5S32S5aU20sKg+ZCuLFzGksXWf
HNQouLdB5sPFzQdmFhTem8QPypRzrI7ydqnvlI2qfwSwV17UvoAaa4EP6ggU+Jqh
nyDsGuOUNbJnNKkJKdZFi+9/2QgxLs2AH81fc4+jn342xaYrCUEhQ6/D6UV5uIlI
DZz0XoC1z6gljC5kmTjzVgUcUf/XPSd6ql6W1/pS6JpIMzLuYXk7rP3VWwT/Myzq
XAVbicTIq63zLixprec/mrM753zijmBNqDX9zZqerQXv5nWGIPJlzgpiApPS6Xxj
G6U0PU89da+7iBwE752/Nq9SS1VVxdIbJ8CHvjx3RigOUJ1fN3DpVQ60NggO+7MS
xh9zW+taydFsULfKSaroBi+TwLZyOLBny06via4YlDDaCvfEf92L/7QEjvvcbibn
Z3x6gLZFnNnpPQ5XYFipu1EIIYDz6erakh9VpurO2lsivzZN5gHK2PBpzMxfqJbC
+JY+TeRyIqQCdOcJDgRpwZoQPc7pt7W2xrzsXtpKomOOeSpFAhefgItl1XgzrtUx
uTGonCYyN8MLiVmQBPaYAaE6hNrtK8LHTLBoPn4i8m1D29TIeqjB43vMPiTWWQMF
NBwJa15whDos4Fo0tyAM5kXgRy21/1jtR7rRxdHwgPoEOvTovCkYC2l6bTYptHDP
1FW0WLMyCq+rRLPPbZySAvROJ70RuLHSNbdJ7WmHKEjeYf+tRWQFWhLLKNtqx+Qb
G9KRYpSgnw++vhUMFPHUkykMAdEev4MjdcqJnY2fZbRZO5bUoI+6zWbeZvlCkf8h
+fPbjM4J1NOnU103y5FMv+rP0PwElqY5XXYNJV4csp4fUZ92dIBOUF3Hm2pKrTK1
ZPSSGyWXhB7b3QJkuUhC38dqYCIPoZ8uMYi2KIB5l6actfp7sqO5XTxnFuO+ScQI
9FLlKMt+HGP752frOyaFibdK2QzX6+Jr8NBBqR/DMnH8At903x5F6MrQcEaE8YxT
86UWZa1FOOk2+kvaqvNLxjaNqIIHTThbXnywie4ehzaXCzztf8Qfv6YdJA4KxrSv
F0HqHH6hSaj4g33Wf+od7OjWS71F/v+WWBuZsEssyuIZp5D1hcLPFqTzxyzsRSLw
8MUInEDJbLeMmRP/sZKocb0k1DH8qqI4XaTa49qZpIC30q3sENXrvLLWW8duRcK1
6ljAo7S0EKFcAZ5R5h8r1/+TdGOP9k2SWm8RQDsmEnsrApYwtCFCyNiysLtTlR3u
tB2AzCoB4q7GSlsPP9gGacx/XPAZjXgdxkWQ7XH+JY34yUugKLfmv4+viNdz9GR+
6zl/oO93JZIm06xv/db1TXpxfdOxFM0ueKPrefH6bGE/OX1lYzotuvpn1p12Pn/3
IGae7cI3sKDZqKgxB/ECJlmN0jjC6utnIYLIlob5gwvcuatFNtglm6N4XsGWnJwo
xSqmbomHlqLnfSAtJqknV2pNw+ve2IWv7ipCN/rOeZBb8GuSx2QlPIGTcVF4bpsF
gqc85wIxVWiXFGh7qu+JQ4MukzpS1U97LjoIVyYyq/ekiFZd0YY4Ej4vUZ9Z5R20
j51S/VYLzwfbg+dYCeZNJOfOGjV5/plLtPkO+N/BozdXYyRMTYDVYDMmjvPIcKW/
CQdhbOGljA3Lv9wsRWQTcFkdI8GCrN8zFQar5Sy4YeKFcmdlDARkD8YCse/kX4wr
60+nDRFhefXqfilSycq2YFtWvH+F0gL+HW5TQvieLc/cZl1P+ATjlfAniyskpTAH
KNw+LFb1fwrEMj28L2MFHkRA5Qdn/zn69VCtxJRefzcqPmfqYmxWBK/Ysk5oHdpy
jT2WXz/sLBJJd4veEHOkaTVjXAwN7fq4U52FDndJGwXHjGGJk9Z0ceg2eJPiDew5
ZdKLn43T9VqRPQ+YRodL2VkQmoIAO0jJ7CkDZVS/pBON10ePdhNQ5Heij8cJsrhL
5E7kKA+hfS72DlXIRmnOIt8WOMSYS/q623BSqfTBqMuzbsL6AAGJ81/Nr44R6R+1
/kaC4qThuPJOToT79yafBDDxiLMyjYZBVACiUWxMGW+22w0rXNoelqBwS1FaroCD
HsHvEVtu+NOd0NAipbJTJIjpJgkup4PDvuLKAifoZ6GhpWFv5TCgcc7AGCm+Yf+Z
ucHtMT1ZXcQ1SCJbaL5koZm16bqK11VVCLDu9BhX2CDumhfSGFoOix3pnUfZ2jKs
rguHOZ85MhheF9idWazaMG/G9AR54VKWlBmGoebQoNDejZVhX6SAaRBUjxV7nKqS
yMbfatbPidroobThZ880TvqiqDGrc0EMZFLuNdROUSR4tII76emhTD8VM2YDnvOy
B6iMycKlsTXyafRC9TigOtQPLOL+3x+ck7AGtzwz09MXyCAITI7q5p/QxA+tfLaI
BmXgjKwEEw+qxEcABOj8L66wibpsrl5YnwMfN/gcLu3PkkWA65FDwAdkNveJ53cG
OpPGA/+w4kvDJH8swALpWRCuyx480qUlinGIsLM9J7FdPovDMvh2ZAo61jDkLZli
CrK6PQR0eXBL4Si5Xj7YIR9elDI3qz/sCeQPU3qN85RHQMcqNG/+5anRmCnxok0d
xmHHSzIbW73SAgri2uME+BZ+BSxbLvPug3yZ0D1c9P1gLuZXBsfbjb9B+lCH1O4k
TbYEhWiZOPloCr9EqtFbwXkBx3CFin5iS3py9hCDRSamDTNH1eQ2beGpHW+iNvMF
Onytty0vPF15KK2Jf7IFrb1I2wIhrCN9Mq7JCOkrO/eQC2ktzkLUQ7HHFPPzWEAe
C5bZ69ESndfTLn5sHRO6jrOM7/vlF9XO+m8BdlRmsS0kCV9C+zrau2grTW5v66LW
+xHJo0MargD16psMOU3Zyn1YuzP9dkksYW3LWCMIOsX3JTJ9Xs06QbadBGWBqXxj
1sfDu3GPSoilzezrPuGgKJRyu5CVBFkRknkGKMeMyVZ1D1Vcpc/edlquXqiqP93x
Cb6tEaxItiO5DkScQWyAwP88SEXyiU9kXXTZzV5EtBz8dGapyvgI7F5sEO0feofF
VFrSJ8z7fiSHqjQxWT+xZQtW12Vm9qesgszkR2X1GDlU++7zSgyuwo+hNKijmaGh
IiPoatXxuUAPfgbwhTrjEg9Z4wrX/b2h92sm1S5TQQaBenm/kerAg4py481CMUVY
1ubG0SLtkv7XKcjH5825VL23/GN2kCucvHULj2ozBQf96kv66jXq7juYzkRIVjr2
7P3opGr+7Zz0QGQSMwlHsr1UgzPKqhj1YtDMrWbEugDrD1AQP0XzEiQx6iMwNG1t
1q4gCMCY8Kjsq/+FSIAhwDDykgIP0tIwuBH77ZLTsRLvxyult0k+2grvBuaWbWrs
QfZ/4P7LniL6730A3Dr23G1urVBj2f+jh61kGjSN8JxsNE2UoF+NmheWhWa2oCSM
J6g0vdE1i2bZzzifPtwWijb3lm8tyzXQpmWM84wfTlJtGkzRUd64Oj6ZOEHYTsXl
+497Elhz0/2vPAnlwLv6eBrUTAp6O39lepX1+DXfm/KTbJIkxNwFsahM0lX3Vo67
uIGIjYc6hOV9EPY0tADDJhxOZGuyhJ5EPGbEz7uL8YBJZG7bTITvN3mPFs/Q0Is3
hwmj0QNEnCWf1z82o6JBhLDnSo1HFT6XT7iUrfjabYzgTKSul5zS/x05p2SzXQm6
ld810GHUZQceJBmx8mpp+xE74WeX3c7OSthBvFigUNuxIf9Q0ww1sEAB6GmKxTnX
6A/l0VW4oU2CeG2yiENFziPo0lIDzX5s7Rm2/8m3T8TvMxY28c2uCNsVlxiZFFr9
7m1LuHsDPQG9nisCvOWmtaJ4AK5DwoaTerFaACdiWlujVxpi92C5LvKo2ngUf0GZ
jaSzanOg7bBaR2bkUfbKXS2Rka8SaRLnCH+hjsJjSa59ukYXK/Tus0LL0MnnIa8o
vNWxNqHH4en54OebsjgsezIaFtc+C7exi96SmBSpKh8dXKnhIhmqI74J2lQyr2zg
+wqrtDXRitFblUvUPL+cVdd9ObkFzngr/+iNPa6sYNVZpOgXNAL9E3g5j60tFDFH
XjO55kp9kV3dEkwThzuTmkg7LU2zMBRJ6n2+EzRPfLIqXqKH24sGmci+zJJW+nT0
cGxDD9PjV6BX20WHpZUhEnLk2Xe7kOJhq+xeKxRb/ojRC9KC0zYDhnbybfAgDC96
8Fo8q9fQmYTyg2No2Xqav5oKvxKJ1JzOW5CsrDxmWixt+k4llAX92I08Vpxaikdi
xwWKdwC7O7L0I4whkzjXW5EW4Rd7s0p9bd3G7sH1wdyR4zu4Nhvd64TS3S5J4KZp
1DV0IMFphwF6buDX+yVAVq7ESRDAFtjNWULBo0uW6SImdsyqjsFwi63ae2DkPOOT
yKrgWx2yL8q94UQRx66dHytuamU7Wb3g1iqYi7g9GK0f37GjclAcglEV0L4WmQ6R
4BhYcCYYPAkGgeoPj8D5wrad1xt1FYJAi86MtLqnK0VXisfaMGilK7Feclrhjs0P
aHxQkKKpdLIGr0Yxxd+4pGzZwne44j1e4ltLJKjOMHju6m+6PlhtBEhZ55l/V4qI
ewsZA0/VwlJH8VLwhCpQeA13HMX3/vhUPI39jfbjxatTpXSn63jECTCW9zSg15QT
XMWd1x/pQdO3wCVpY68l/QjZx/PrBxaFi2dEFWdp4REeJIXBVbNfuFUnZ3SRnwBM
p7NhMRCFCfrBD+VfOTBTCB8Hp4nODsISoFCxzz1pN0z3xGjbPvgDzAL85oFYU02l
b9BPX3sLyGAdb1ldGYzbfaJNemgSilFC92SAO+vgcPpqwjGzOEFEV9F8W8JPH4Ce
4qIq1ZHx6Pb+GMGy5oBoQ3V4VHbty3ieVE1/x73qx9SBDKYhELM/Ea08pmlRDnLv
UjQDoai1mOdOOJWPCmJ1Q0VZRM9jjNXgAU50/pU/pWvWe2bMexZ7w4kvwfZyvTXO
7xAdgfmhjEQDBkyHd3lRpJbybXY0mfmP0HfX/r5MJPEh6mAxJl+sXaJhnAutZd0z
lQTiizbl5r5ovBWOFo0qUBgoFUjSe8Kd6luWbcquCmgPKXaYLTwi9uEjPb6P53b8
ucge/vVME83IqaeOea6SNs71VocDFS/LC99DuGY9lakKm9dpPpvtYdPEHXQNSntU
MKo5clloAj+eCO+s4FhkZafjjPf6Rm264WfVWQMQJOJ+tBpQKHTHsEZgWQ870z36
vnJ5sJqzKixHiwSKz5d0UWe6SHkoRQQ2Oh8vDHCr8JcPLTkAxc14EOUbogLCxE+R
cf/qdFIIcfVrTc9Bsr82reX7s6FbLsGaj+jmiG7YQkT1r/7nSTq6tE/He8W7Z2KI
MGUgYVok7visFw7G6vHE1mvBKipq8vqw+pTaA8mRg+PMaVdiOd7RzuBwjDNxwlb2
C/+/MBPV0lKvVvo210C/yHtasy0Uj7IKUEbbf3GBcXUqCu5iiclufUT5zBKiZuDA
obYIcICFXy5Gq4C/AGMKBJTca9YDW7GwZ4iXsGX25U3HT0S4U9gO1FAp8jctF9qA
H6vYU7B3DgFZWlTl3sLOKNlwmhHZWK7rZaib93h5T1najBpNQf5fX7tYbxnM86Ek
BmQaDa1cu/gkq82moS6fiF89rAwvFAdbrPkQYeHRquepMEouI8/a1C8YV3tdGP0A
18gqbDhRm8WHbh2tVTHHea//+DWpFld8XVofUsetnv2l72R54+ccaS6FjfZve6UU
q7ILODGMZ853dcd8/XzVIUkxN1e4EJ0mSM4dfcPYQPqzyY4gXRQGgENUV8elWkMD
IKegslcpjLGbRBQ+5+evHR907z9X9fQkOdS1BiPSZukbv0UU7D8RFB3J+cr8Fhl6
yE0CuGjuOpjPngTmzbcwdPqMR58ckw7UGWlWVRmUJ8DHGD342rqCLopXNf3wTiLN
nY8OKpv2+ZbNKr9JjGt07np2XCwwu1ck9ogOt72iI5NiVT3wkGS9T4kq/g6r3Wad
g8tcv9x1tLYCofnqmdTw0bIQmRXy5WcfKJWrIpo9aZq2tkSsTNj8fc9UpI/6/Lks
6pZuLtugCdvtmm7m9XbrZP0V/IZGXvev2f/eK4JM7S+lzCDphcPyTiHN1RKx3KSa
8hiFMhLpQraRXGcRAbnJi7dRR39jB+M27AmTo8OTyX4faRcfct6dybQ8Z6L3Nlkx
AqO2b1YItNryHsLOQWrQ0N2Rr48RD39STGg9pvjmV6VtW5OabUQSveHinmz7LlpQ
tKehTGAfvgJWxGyLrCQJCtlikpAz/fM55U3yHwMd3/0DGjIjowDp9/tJDj+wWQmQ
8+jDma7jP4wI4jNR89ZAVZXSDDwjVVN45rDSWmBdnHLT7NgVo/e5XEhRe/bm5j56
EMt711rvp0InD+D5sExZHZENvD4FCB8o66k18uv34GwzAClsAWb721+xIak4vl2q
pp6vaZc3d1IZ5SdEQ06fCZMF/nyBUhrSRRJo1lFKEgawek3oPQ9edJNCwgjfxYyT
Jb1hcxf5vlC4LJ1m3xJxxzZxvd2FSi97FpajTP7wg5fHDZxxI/IiSgKP/HSHaQmH
jp5Ttd9OAm/v7FjBfqG4VN381EW/uCc3+8kVcRN4vePcgpHe9NrUSeCGGs8j0bz2
TFr80sbwZOWCnSmbHlTaMyZq2eHzS1O9qYm9q590GAyqv7R4VxwgYWyRBChiomb8
8cw/C2LTVozfbTzEQjqac6Rli+JB0Uo8cTkLpUOBNhr/XUxlOvhJKMjela1T6xyF
g+Sr2CxUIE4l4heCBVeSHxRrNiXpQA56lrhI0NP37ha60L3mkv2OYZnG99/oSuac
WoeH9MFpFSWcIjrGkJGBP5AR2cA0AuOZTe1Rdhz1GsgDweOxkKxABNkrX1282ypP
c5Nn8BHht6pOD5HYyS9OcDgFj4ORYGxvMy+jehQEFt6RQhW7sq9fLGYs54Y8xj8t
nZ91sGVQgy1drykL4Fevr+U1HbIRwrM6G59S5929EtXAYM5cZjGMxd7ey/MXzMC8
dYhFNUEgMqMGJtBEQ4kxUi4NPEe9OFAVSsyYgcZkzrTOMNcDLHKaJIePB7+I8Mbu
TtBIhfxj6IKXhVgGcCMnc5mFgxWAirD//sXNRa6UPy5CzwCd3aCci31ABmLJ5LY+
Rd7B5NnwFCsgCVG5aOpl6UV4md3MBG9NoBA/qoDmhVPNiyw4JvDw205O7yZMXQ9E
hwzupPtPF1yl057zE2cklaGEfQbS2sobUyktwzR5c4/Uqzsw5pT31CqqaZU8iw9b
NEzUdZrGcTSjCvQDvDLGb8FK3MgY6kyl7w0N8jLagH8RfmXxf1v0DmsQ6bhSAOXM
UhRqsu2qglTavwf8Z0vlwfPHXZdsWtGmFdpRXv4WmCCHCc0DbEiU8kxeKinudkSr
9CYM2Vv4EvX8kycaqt9lmSXkHEJUZhOD0pOUFgNVMhjRovddAHemZ+6zdDwjJ1R8
+l97bBVhpW4pRHfSZHMKVEsrXWbTdhr3lucTcLC8XnypofZHmFK5/uSEIpIjWqf7
teMPSz/6cLXX5PCfvKkdzeIyHyyyz/ksahU1b5v2o6iWjVdUFkLvWXj9vXnqMzcu
80Ovxjul+02raBjW95ngqMf7chy/7QWHG4y/ynhWaXLzATfZ9C1wRYmc4rpHOpUz
IkYasVpqbfma2CJeyCI+8xZkig1MfLQQaqBqFxHICKW3ZMpNf86M3IUY9hpfRlzf
OxgcPUVuYfuOw2v8Yx06ubQssf3vGqbTj6/4JIiDrnJSoUl35P8dyblRkfDpFrSv
SknQXIwQOT9jObiXA60LJKaG7CMdbbfIm6J9mAMuhO3uBuzpQ4eFsRnlXzCn/mdh
ZfYwfI8CltY3b9XAr3ZUZrt1KnChQjz6TCJyF0WNa2EHyNf8Nu2l0yYji/vxI/Jw
g0E1cSJc8HE+W8ePd/Rx6a7e7e3iulJYSymwISDYGRK7fnVisTaVUILWEdxVUodZ
x2R1G/+cFYXNoWXHHAAHYAFXNIWJ+mFtfeY9hRtLw+06X2Kct5it1eSZ7b52nl+u
hezRhKsjdII48HyNn6avqrSgpt3lKA6FPEyHAUnhi5+c8xCpaj2O3sH8RVMh6mY2
0+XbdHG8B6i0Duj4E3yHClzUH7a99VyRlM+aJ40+kGtUoO1tyNFK257WOYq/GdcI
QKSxCOul0m2yr7J/tIe6aDikMx6UyzqifrMIqEdtMwlC14kkD3jHJoWT0wmgeOpK
YvBx5n2pChhhtdNj8u3GzV8y01tp5wVfUsS0aMsfs9hSGqROlXlx6nUVbpYUOCiX
CQ2puiwLVVtOT394B7xeVedKmHuVrw+CtgZO25VlgRxuyXht4cZX4+IKhkdAyISl
Qe6IlBFXjKJbh+EHmlPGDo1osDCeJOrRu2NnT4eAQw5ZobZH0CguTBZ/xQufVX6b
ECPvqWjvFtUJu6rZ74RlS8Dp6nFZA3rGkqhPOxyXnmQWInYmuwV5duKZFItEMONF
L2eoiHLFL71na/Vl9QZZYtDCONJ2tHOXSV4VEFREiYh9+yMaGzxtAXEcEWOK3X8K
34TqkjHX6iVRfwTNAnT7Qk9oeeItFN8IhWJxkDYJFbHm1O6ySfMguoxRJJCAuS4Z
1gM7MLUMmnaFSj+y2anrrLaNmRSQR3FD7d+97r9WzZWUbtit5ZoWmJScSGOh1y/G
p4nChj8QtQp+PsY8Z+zP7y9O90nk1NHkZbUEqymCVdRnr0taurMmfoEO7Phe2ztP
Ve/PZKOviCOZKRm32lYUhuoaVV38PIqIUMnmOMyAOIA9wXJNwlwamHDrhCJaa2jZ
9cJOAygZMmnTZJAc8VEvd6C4P5jDTzA17IVepz9kelSwTLT78NvJJNYyI8FwkLG7
f2+rP3vPB5BpwypNqWQTqOCUDRasP40G0B37uGaL31bGFUhB7q50uFTaJKpnnQqr
2kSnXKIo/AxVH6HpwA4fFlEJ53WT72g82fK8Y9EUSpGq4YV/vz8TKcts65NZVMOH
qn14HdtSHr17XvrekGqq+IBbx5HzsnCIi7Kd3p6noTK5vMmeMmk6Kes/u1OEnWpc
XFsJVE2zW2lf0y8nKo9fgWjKkEtrHSjdHkfBNFSGlB5QV0VmD9MA2exjddmG9lP7
PPg/xC9oSz8C3QY1TQwrgxfEgfyNKObM/OY+gv0j/bKejcovaRmzh+v5KZBDQusM
ZCsrP8lI4+bAX/hA49L02XeySbq/vjV66cwhLgC20BoXWM9bJeiXAo4SuPcUa5r9
BrTm/a53gwtrgJDHyyhVnIZoXaE1c9pp35/g+0SwThOpgYAkqu1phCsZ1XvdU4oO
R7fqogAfzxCGEryt53zjk9OzfRbzkeCQ2RTFACb2Tkop8vBZaY9KuCL5aRSjaZEc
yhwdbAa1q+q1s5f0XaTQx91J5ainpyhQVsqct2lKJcY3tK92W9HeT3eTIH4nnrFg
Tc2qQqJWDudAK+BfByxa+RcN8BPK4EdBKG4RDOlf++Ko5+Jaicnp6FgOauYdl/y9
t4abhlWP0LzZxqkKjoHW6IYQeJiigiuo3gTG5xU57tR/sbb/tmC2kUQeWxfSgU/9
Dt58S+A/AsVxeHSNVr47Tw0HRt5qUTfV4iPnJpw8P/7jQAyk1ekquXd3VIoIQklv
lgB2AOb29bq/P1r3Lb36WL0Qh0ZgcH6S5WITWfCvraz/bvEd79ysJ7B2INSiNVji
iL/55V6mF3e2k75IH8l032/MwzlkqofVFBL2BsJacrNOsyYkclwt6X2FKbfK4MVI
URp9a31VFRFkNLSf3LSWSMbEZ5DLgPQ/qjpmx3OWPdInBbdVpMhZlWB+thvr5JMa
ae+YYCQwrWvfZ9x/Abtk+lyz05h90nWc7db4mikkSu4SNwMPkDseyEea5Z8B5MLn
GFzmLqa/OzhGW9e2DVPWW0LdC47fs9kQC4lLB17SDRbRbHzelTwPwSzaeRP+TKE+
F+pqiPF7xZFu0vzngZMRnKL4Mdeze1YzLztdYvxVw+d+/xB9FCzDUeVoKtrcgzeK
XFMCP2mmqJ+cmXTytAFnp3SBTTUk2Zgctk7VpFXsFRKbau1G9EJanNmqDiNUlkMH
tt7DTS3Lf0Qj8DZ0PFiEzgHVHlmcYwu+GccXA4NP9Vbduol6lfL6vtjEns+D1U8l
HX3PKY0eyqc3JX89AlhTV4TqXPvUZ1AwPzKZavPgRBQBGAI2zMdUdhSnuDVKTVbQ
ulZleHN6OgaGS5EhokeoHQ4owjvVysXTwsP2UMh6WQCcby1kk868ZJMpgTpukX27
iSfTA+pWQAuCboyKMaelpNkS9DHcrv10RDNjDBYj/KH4KyeIVBkpNeMPMpqgkeOr
iRC3bgKq5DhH7grL5RYyK+OrNQh3VE9KoZ4Bkt/1INnz6vFxO7NBjQQ+XRceWdyg
UCz+p3GPXf4xFvfUNWnPj3AVRcyRY4/jzqVtS8MYOJJUcCud5DKuBKMOBI9g34qM
4jzFPMlqUY+uzVd30z6Ks+CTd7ADjXnQxjrLS1VJ4Aj+9mP0kY0eH0bbCxu1J8vc
i7TvpIvHiraFUQ1IuJe2DTcIc2/IHxGCzbxLsasrCCupqyvjKyHdM7xOLFRUYI7I
eBQU1Bj8qZeY/krJ8q4qrgcsXZ7HX7gKzSrfpSKXsM+TZ3JmI0BAe5FPngkd7OLJ
lFmLp/qh5g8guQtPOhlkMFWePY52vFkpvTHWoBQeqKdTU1lPGDHCjBvPO5erU7jF
OShzoiLDuA9ddr1Y3rzIrNPxgfXHzT5nY7G6VNponKeRpmpwGADDho+To4mwxlu+
w7DHnvnVsRbM0b4yHIkO2+tPf6A43Ric+oTg/KtRxpVROXwzNzwN43a0tn4sHZsZ
jGnO1ggY412Vy75LBs4CsDCKhFBI3jcvI047iEwUhBdEHUOKzO5Ky/u52W0iPA/a
w5+bFYsPq/P4nuWaqzlXqRmlhjidGcTafkI/HGpErgHwsbD4G/eUI4ZZZMgst8DB
w9ekXayVcuCdLQ3gxa+5u1SvY/spyqQ8YgpjykzWI7RB11owGqkpQosjx5uZAuk3
TD5FwAmqTHMGjafK/9H3KamwFKrTWNcL6nX5sF/7V4+/51D2qYtwlR2gC9QOhoPV
J30X0XObbisfni1ZxJDrp9YQdDy9eGfIHUZV5polZn32qfuIRdarS5G0LwQmLlHG
SUR2CXaxhs30ZCiiev+5zunA1ijCCXuB7GWO7wvnXE5bCfD02WHkbwr1EEhUKSQE
0HEye1acySD2K+T2IKTOVt8Z2Ryg6xhI9VucAtmbd8dEoMncKpc1eJKQdnxd0lyT
ZtOjQ5ltwjqSAzhbhTgM/Aof9+bmuc2ixvL1sTjwotdPGLPmY1Ml4GFuD/1h1WRF
mc+aithJWbBTvG/XA/8LN+USI9adPVzmCSRI77Gg11u66wYDYzx1iB2cEjomYDsk
dso9O/XKmX7ETbxndNb7MgXk54q46gY4IE5+EsJ5Rx5tiZ57G1SVmVWI0oLA3RBU
ad4DDeCCbZOR44M84MDvcNxEy806w8AirDBAY10d02g3nMNW0HCxL9PnXCxJCyjj
bxe+SdYNtKmNmGGZullFromqbrCnFB8NUeikFySuUGxbdeOT98nWe57pcoSwl8qL
BKoSArRZs4mQwdd+Ma8s02YXS51xGUfxbzj+y01K5cvC/oOHnQVoff9QvZqPHrax
BVjKplB4wfcaZXl85CPxLETC84vlvPRGl4PKXBFLsAl7xKoIIyGWm/4qxvkTSjhv
VVuwq7yXxijHkQg0TVkTfryRAlOcKTNecQLLIoQPsqc8yPBB09aiOnEUcjfU5N25
rFXU9MsBp6cMz6d/MtfVY9sa+O8r7UWOlELvyTmvyXJPlTbPZt9L/3/gpv6Aa4dd
wbQRjCvqMwR8QXET9nunPM4vFRu2WYMvevT6A1rbjOwmRjhtpAqgniG0vJEXq/i4
MKlO1iwp1Tp3pjQLA85cp8F90nW5POkUR8E25jEMdv7SY7vcz4yxufZsKr0upLSq
+gRXJVvjGKQv2iUc/GLErPmtDkF0j/NHy2xcl6az7tQ21o9WKFxmz0Lrvb/4wuPg
eAXw1viAB3xxUs+rCgv/ZswI6/YY8E73dHd5jshgIoU2/9tGQYssEjIobeMHoyp9
/GIuO70aW/VGuI2CnqkzK/JCpmXENXrO8H4MGfnlQqh/0NIH1c4s5zSIf1A+oyds
tyAzLU2SPgUYFMAxARREf4Hk1seKlH9yWXk/F46SlDRMqoyHrg82rycYPQ5ImmRC
1UtJXaVW36aEbtRwzG9ROa5L6l+3pulg9iKqYGEmvvpO7eCAJUCP7K3mrfdUWxzK
Ltp55iZHNoZYNmlHMdWoctQE0+yc0u9U4O1QjB3fG9VoMCGQacTn/Gm0v8h4fQH/
hsLMD9Cz8Q4CSrP0eQcZqCBPzpIO/JGxNn7dgmr4BX7Tow9SDrRkdqT5ScpDEo9E
90jW9Io84kM7MfmhUtyNL/mlEKzP+VcSUtLLTfBEqXVbzC0RDkxCCKfq0+TTDeet
32wMCS4AyPcIH9vm4IYED28r+Lq2HWkSYeoKtcu21XgH4ZISFy0Gt/dnz/DbzhJH
hMKWNX/eObjipnVRRU3jJxMN9rXHhQdPqp3m4gof5Iiy9SSiC2B1wpe4+t2t6NF9
8sRu95NnU7WUARHKd6rNBXbgyvAzGrPpLJwJhjMlZZurRqVdtYBlyFxQmUUPOXed
Zog7RyD9oHfBgV5SNtN5D3gWIuwoyjZ0Qsk21omTIQth23vkdHwPaHM1fX9Ty83w
BKBsvbOXIa8RObiJg1evQZuoRVwAMNyRdYURTHf2YRklcqrrVpqndBSA4+3X2/vt
oHtBYfSpFZbHwr6tGM5sqT6O0A7eb0dnrxH5ptnBcqzUNndbcpLAMPqfla3bMU7i
15DqQS5QEMlSc9brjFlfTVqt1hN30fy9pNPq/McT8gouGMc4mg00E5ee/cXAgux4
gPrlYXvOiNRhU1YFRFn18xIYUiBmJPmnb2EpWBGAcNc+Vtx7zUvVzfFMdEQM3i1H
e1S0zozVS/xvSpdEjZHh6/MeLCTlKNlRNKoMXm1GS3IganhbP2pGPgEGwGZhJ4gU
S5nht5JaQwdpatJn0PkQnKA/YmOY9yK7SFtsOJIGk+t4LbgpjToz7GF7eNUiEJp9
owBMv0OjU1Q9Z7iZzkvyMe777fSHAP6FY+1an6fezlGHKwYNeHhdgMtK954Vz9Oq
l+mPJi89G+B4UVW6I7lYcH1QK8Bt3QM34VknNznKB8z5Jf3AcapRdlaDdCZboeLj
2HlMfTljqDnlUtuGb8u/7aAZy3lW2b45JpUM+/sFzDInG2N3zcVFN3t5/cn4Ac2a
PR8gzN+nID264M9hN0HkhfeEytlLAKfFQGiwD+GxjjOe54pxxTR6wc6NBYoksGHg
wwIGafAniYk6BSwhhM2wgycTfGqDjE6oEODKj3FCIYoVU2U3HfQQiqkz4SYV4NsS
71o8j3sClLFsbAEt9dqNScUfNuzBJCeGmR0NFPIZevXQnpNaueVEbPa76ByPcfiu
Zs/balLIOlhLP936NcPKb/xUunR6cPIEfXUdZIVqUdPCBmKLzWoFpbbg+818hEqh
JG9toTXEqCrZp0n16UeNb4o3XyvGbELa8JpgkOj+QQGB9cQTZFOvhxhnX7lnrik+
qKI2ewmHTfAtS3H+9d0GZ4hFUCmQRdl1d3Q8BTvl+HfaR6uB+auiBix18DWv+6WY
wGJO73Y/DiTo45TdkbwvWrBva7hJewXxEkD0gVwKZXlw9BMuF2EkkQWAVbbejoOi
0KklMAI7E2K3OwvUPI+lhk7+TAaEpUjhgQixaH37V2gqCjybIKo7T8GZYAkj9s6C
VwpzojbGpia7q/gEi5C140IGj7D65ZlJp+Vo21jGEV/NlNqqKxuIqdERlhjo5CUF
6bLSOSG6bhIVgX9Wq3MnGzUr9lM8ssBYAigIHlj43BYyA0jPhLQj86MrtGCYt2fg
zMCWz4UVvVYinGY2kWykNStgLEe+PZb92NiGy6kW19yfMqVV0J9EjAKeZKAs1fOr
DYxWB+wm9b/6TPgL8rOgLLbf3kWtaFRQYEjGzQetPnF5Yqc5LidgAzi8Mu/87KLx
vE59S38cT8IbYBZP7SM9bVpFkLpONN4ktKU6mmobuEMByvRYb18gSTBlxuyektL1
rm5IV40JqytlYfNwWnN3/KZEvA137K65YQZvRI2gW7RzF0zjfCtpadHvBszHLWhG
SdLM0E8hYuKWL2ydZmagFVp1PlnYpGnJhWN979SlqH6J91ye96lzrAxfG2D8/g/W
MoZlJwsLyBUQ0fZTBZAt6R7/0yQyqEM2C/fNz1NsDZ6i4hOkY4pJr/Sr8dCLR9Ty
g5JrQSQjDpvyoI2ACmfh4H5Cfwfah8QbiY2PPwFCxGP1zz42thkgmctWGhk3Siwm
1RNOFFmVh5kRc82nlFapPs+tCQuM+ZveaxZ6QVhnSVgf0ZBWs6tOrRnK86G1xWSK
etEv6Trg0CIqJdTNy9IGAJn7vAzwgQWc/jm6NHbd357S1qFp4RS1wdywM4o8QWYO
RRnkCrFfuD+tLzIAgTnmLqcMcAKeJffdpLf9cMC+tOnJmlAP3db8kNH4GCgwRhlQ
lhufVWQv9JIVnQBmYq6inOTxght/nqY2jpjmmQruS6inqr//Vv9sqzgIaKHW02QO
g50iKP0vgO+YRm+eIvqt2OF57Oz8KvfJYZsZ1Zd4ytPoOAC+3pH57lE3NWU8Q5oi
fpFI96WQhokgHpPFI9xESYxaHcGlrAbqdgwRzV4bQ9WpP3ytR8iuFUYeG6Ata9m7
LHJ7tGPvC86CH7EKOHW6cJuOHVlofYNiCBBHM350nTTC0P7u3gFsuAA74d3+cx7P
vodJ0NGGK5Q8N4tOTrtVeALTRb4SYIcD1afxSJpEBgV8X7uhNymLu75vOtmHElZC
PTD/vMKfk7rUhwNJif440wf+IebauNv82AR1B2awe8rqRv3DvBeCME/LRKNr68oY
NF0F2M7VJGzCOhKQnTJFSQVJqJFk3kx+g38cdxPPKzbL4g9Iet2qIYL8Kl9n1sDj
BsMWEXGWQVBMdKJFKMHdRWB03sfKZzGbb8ZRIrojVQ7zmPlWuIxQcM46qXoomVEW
RJMjOT5K90aA/w0j4AO0hHZKuBz0Eo4+WBpAREu8GKS56DE2nHHxVb/KlSuaiuDt
veqgHs8HwdQWdDeBgphLlk2RDgkZR0vsTQAiWHiCIOcLzWKG53BrwqKveQLyp9K+
no4ydpAN8sv93wSXYaoQ2baoprZQRbGFhrSPYpYxwaRt5FI21BFHftRSmL0k+ZV4
6Cvn1c8Oif0bAP0PaW/l6FQqSAsTGbLYUQC0oy+84wbqQokSDz+NPnPUEBlb1Lsw
xxV8Ym9atMXKbtFT96S7sQb/nZ5gDcEZq+uXlexlJZ9MhFpxPdx3C9/nJH6bA8yJ
nrhaG/Odbpb2HPsGX2x9LQ==
`protect END_PROTECTED
