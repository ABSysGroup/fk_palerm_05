`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ETe7sAzN2QyYdWPXs5BnS9mRrsFWecQMBKm0LBL9POgs0BQarvK2iZ4opGbwelbF
BX5tY7kvNgPsoAN13E2vNNUffFlWgkNfZILYBc54+1ziHV0slZhSgAHkk2jXbJvE
Iu95bUWrElFJmNABdEoEVrJIP8pikNGPryRJE57cnrbHtyS8eojA60gUFW58HGfH
EbOZaEzWFfM0RxXVodS5vXwF7bF59wJFn+n9s0iJF37dVlIcs95T3Sk2lbrWwkmg
vfiZoDVNkkBN8UEPOH4BmLX6bi4joIdz71lfp6PGPKAC3jIeCE7upSVbvGep6kSy
ZrfQcjaRgNBknqJxHxJjJ0JrOeVypyxFnL9Rv3uGjxCfHwMpkYtT+ersxw0+/dyi
b4/IaMdxTw3N9yjxxtRIxftlAqOXaDvZiIHlxjVSQwEpsz8AqfwoNnLMwqf/qXb2
5kU4qHajsLtt1n6Ve6UJOPQ7glDLCojNgIPxAxi8AL1huFxbFQAEv6DtRGkYj0fD
qjI88w3UMxgPrBoAYcE7cqMM1gmnCW810ydOiNIR+NK1YPsperzPWiKwPs82JXKX
mdAEGB89paKdlqeuEnxyIQA2BYhD1dbeMUKMpFGt5XC+eFiGr6aE7B45Rioa7xoj
/rK1Cki/SWNMMj7Rnu9tVU54mJGs6elOXPMb80gbq85IIP+rTmybG/afqQ3R2UWE
o/sAcna5iFvJlv1VfXIQnhfd7R1MiPFV1BTLTDp5hOxdYA1emdgqG53lAqXWebVq
jkcYcwdri1cFAO1Clu6esryNYC2u8XZnoQAjPBQOOqlI+TLk7Z50ktR0rVHXqU8S
t6JV9EMH1cgIa9SrcQ1bxWt5mx0J81/QekqkmnbfBm/An1gxNK1LjVfVw+72Si0O
euoly7kCuAcsGeSU6N68P8bh5PCKtwCJ+yJh2ntxTx72kHvtxS80AhFcryZsKhN/
oXu6C91MsnjYRikD4I726ZKgs//oR/mDIb2GB6SuYA79TmMo8+3tBNrdftb9ckVJ
FB5OELAMfD5WInidZEPQhEDQsL1iUqqcmiBfSfuOq2CdJMTF3p33fVBaku1JHZco
oDRVz81NPkxypyxecJmbVDWwZxjSaBQZSKMMdWmQf9zEeDkXAUCvn1VPPt6Wx5FF
XF+u5IYJe0EsuiqX2Vr7t1hXJfl6h15EZDV+OuKz/OBRukzO5ESyW/M2vChoXOnV
YTvFqD+CWYu6c5tz+a75JVS/+EQHrHlY/mnKdMG75xxdap7oGEBjKzVfSsU0jOcw
+SuEbDTaXd9g2qT8c/5JLuU6IDZwfm7bSC1ZrEpixU6hunQgqDu2vrZGnK2+z6H+
5VgQ4Kh00sP8Mgv4jYZCzm0OEb6/xaJbdw2Cuzsd+Cq4hMcDS1faab2lZCy1PbrZ
ieNpjGdaSBOvYyp3e4RDVk3jjRzIvocBycfyzWm17+KwwcWTHLWPqSXx7DBAHfcA
doN0M/5VYfMUlNVNVNxH+jEVFZZEdoCx5Hn9947M3cSDQQkmWJCb59hpNhEFH6X+
F6Ed8+M1n3vp7CkkP++2y+t+LKGv9RE8YL1xVbZuBTdztcTcmfghxZ9f6Lj5MQhP
BZyWb18zOr3Kr9ULWwuafSYAo4boXCzRg3KQ3C6HgURKErRi/LSoBYKKw+YgPFFY
ivrGUKU9ZmzLi+Xi1L0Hi3adNzLp/q2cvX11TEKcyWj5oB4DzSTRPkV5oz4mFJut
e1Gu1/Xo1yrLJTLU6eA36h57C+dAZSV0Wzi3nveTONwwNivLGHC1WTm784J1P3ka
o3SSKSkLib8Ct7FAJBIv1PUfZpE6fgZCCcr8EhEz9ngNjJBswheXWJlF1Iqa0hyp
tkZaZMLucdKbh+eO7ooVyqFOpbtSovG5txbV14LFy4YK6uoOk/A+oOyfUnIIb9by
7e1pmUUpsmlB2WHLM5dcGV/riTVu+L2Rmk2BMisTzeFEa4Od5d7kie5qUjAK8aMl
BSCm/W6MVBCP9tO+XZzL/0UtPPKtTbDpA77f0C3tUp2nJDcgA6SG/pclXDPlcV6l
kBaUreIzD5sx/1WNYA41SMBM4cpL5hXhG+8Vhm5o/pVrw2+HI19jsxeiKNv1OG1s
fefc8q7XBBDEvbtNfdUERiKNh1yLVpiesnGn5xvqXdUtrLV/+Qc+MwNkIIXj/TTl
1p98wEjAfopzx5PyBUjnPj+HsBtD4UdHxWqoWBv4mQSUJOiVycY5VtRFA1Jqr9PW
KIFp3qluP8RVBsqT6tLSkRJzdI+jmdVkQXTdgHPigHUdYzdWGZJzvIVKpDZnjWl/
7WZr8RCWexzpEtf7BWNFGfudeut5f37jjjQVApAYoHR6FDKQpIFioHnBApA3Y6PC
uT0skPZWf09CFfn3KAF1tiOlnjny3Iix9mRjOEViZUsoDRkrdhzRR18g088s/nrq
z6AbYQusS6kP4AbmJvlSBYEmKjgVbM6qxJuQjPOMPBMLxyNLu2IoktP+nr8c9Pml
pboqPMOCNDQ/YfI4fLC/h+z11rOuVqwORf6FPp4ZZwtdxiKO79YSFOzyNMurAyfc
XjsihidxEDx4+EYktZ4tBiB0gmhGjRycIdu+ugGptOcNMTgJc8drrw1v40QCky8u
EV7fCJdl2rH4hrE5GLgJVAtkEweTxTcRHBJiwgPPUO/xv6E2ze3YVYij4kGJy3k0
vyIg4lOt8bcOIGlgjS3rU4U8rb8OAJBUIC/70oM6I7tOVdmUGCIt0CORJiONzanN
907SPdp+WwdxZjV8zF/t75rMbGJQH1kP3u3Z5ZFrJfAxifPY3ldL64+wuTR+IRov
a6YpY2CDr6Z2PfLyQY/fw7jW0QKdSLf1lPmdYTu1RDecT//PersPHyaP736RQEKw
OIYll/E3BcJrP0cIbv/Lchxv4pK2/cnH23jwKS36BPVos6x1ewghkccQQgGHLUqK
u8HB8/E2wU2R1mA5+Ocqm3InjLoKg8n5OtuhH+WhS4g/FTTx/DNhqNXvn0B26MJW
J7p+wnj5iMrUMaOp6o1o589e9W6fWdgkEu5+IrSbMlbltZ4p5F0MpRTu671rSe9C
RyVdCSd9U1psCWmiK6V0nb5nrjGiP6a4hbKzl3AgwycMUU7tLZIPh61kbb2tdxhC
ooJdQfyrd3PQwpg9+Y6w/94SQJJ3Oa5/5W1h2CWLRtDHoCNYWKMteUmZy0o706NZ
Iim7wWtEgfOmLGTRTFSbhXNn7kojACIVO6fD+qXKG7c=
`protect END_PROTECTED
