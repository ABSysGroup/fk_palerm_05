`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uAfoezhtvl5v3JV99VtWfuJO81Y23ZTCeH8ZIV0BMHrShsxJ+TMnw3nlmBc0WuMz
ElJuur6tyxqbV+wVnZS31V/zxA123Z9D7JS0vMsbf+Utk+6vHY1C1EDLona28EdN
Fn5ZxrKpjRctZsBnjnmnEBkE1u6e/xJM/RakErFkXTsRySxqsowEI6WK2wdOaaNS
H+DO8NE+A5qXbpXljT0qSZoEz0JxIazppssa50NxgxMVSobJXF03waMEYDeU0OCM
aNgstJg2XwzkG1W8qM2gVbavmZ+Cszc8QNF42mhPTpd65sBdiT/HSxTzXLjLmw4v
wKqiphtyf92mfDSQvOTvMU7ccFzinyy+38HP0Of1td8Sg1Wfhok7bJi5VA+kTmm7
GDPi67jxbbNdx/JY2BB4iUjTup5YqEcRV3W3wHJMcWrswn7TTWhiTM5F0T5lwkca
y/2/q/C3SrBwEkTWv4JTSpg7y1vzftwMmYr1rZd0vJDz27aTZ10dnLz2BqJFfAG6
02LWNADAqADWjA1049yjyO1TYMjwdqKmcm/acSeNNxEIVmHsKl3QxYdlm1D0jd66
hieCPqXEFZ6a2hWrkyyZjnGgxqbVJrtQbtgTECygynqjcYtiH+GNjY0VbZQm5wA8
VDcDhJPqSe04T9eZ/+bXxfoghFdttiAaNrw+9JSPk0Ea4FuZDWsdwLSDgE5ZBdQL
hYhPK6N7taTx+MqI+JsKEcY4aSnznIqPdIi8V/Gj46nUIbpgLM+H9V33OFndTdvJ
cgwYhi06rxNtoM06uukkR/tZj211mPMpP+LkcXL0mvWB4PyhHtY+84qcxvR+3rTs
JnCYlBidMiLoVh53i+ZBD9LdQAqBQEOm2JSiBDFZSXloVPYL1FAFnEq2BH0d3gzs
O5+ZNn3hpAiJhnOX3jVMk6+FAqiYjn/TR346fiNVmsnRgX4CyxBGfQ6qwwTStXRB
xl3V0kD2F6JvH6kpVsHPTyoWgeucHVpeD5WRoH2SsDqIbKYs2lfsVZHHZ1eswQcb
iarPlDKH7ZZgWl1/tD1fEvnXVUd+YObJCx+ki6O89Eg7LEiu50kslE5IR7tsOxxY
sZ/GR5R7Z4HiDXU5kdCxK87ybdHynQFacT2Tb8l3XAnEiIiywmWl1qglTAPnuVAP
JAL1mJxwfpeX6kbt8zgTDroWZs1W2ChWy6pN/beAEx0=
`protect END_PROTECTED
