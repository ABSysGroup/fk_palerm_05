`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WCvo5sgiSPTFfe29h1hZ4nPGqhOb8dlWCzHOmXQ5iDtcsaRk0uixN/Vgd9ZA1iLe
Uvl0skGbg1G/ewlKdGdo6R0szp7eq9zDwk9aU6FW45zoZ6+5Mz91elWcgDfTp9F+
DueGeNBtDL0UpxjVvXnx5+vn1IfMgy0Tnlx/p65Wbr0oc/MEGv8tQdD7CGFYDQbf
GEj5CvSCkodaTnhjfRpVsOnRFReHc+mPfCvxCFJi4NmuwgcIZfrvzJK5CKGqCnSy
xIkq76xptLsj4jQ5b4BNFJoFQGCyJ2i103w2PXlSRxfyyXQhuNJLj6jdiaMVmVlC
oQeyH21POBtrVNa5OkVi7l3F8KUcsTLNLmOBEP2oht/hma4jcqv8JE/phfnoCUrv
6sNCYdg3KKez9W4HmYb+/DyaWpqQsGkRv7z5+3yHJ3CM2y5XmQvX8xMbBGsl8vFJ
G6zJx7BPzznaq05P6zVV95J1WTB0adujb322AUSJxsnjO3GBF/cpdGPnOdwXGJA6
`protect END_PROTECTED
