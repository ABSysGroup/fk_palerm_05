`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AfbBkz844abvl43yVPf7cbAV0+j7SSfaZOc0t/WDZbVUVgWEvtX5QgTfvIOH+Udy
k56otQKAwVF/BRQpC/Rs38JHE0F9ccERoPRF64283i1kXh46EQ1A+1JUlE6vhdDN
1OZiXWAoqGh3FxnErsJRZzzRh2zHAJXwj+bYlBl7RFwOJLqRRlyKR1DPftUTnElI
mUyaxb59WN6ZUCRxDhuPF20mT4lXAL7HUaTvVQpa4JHSVxU5wR1ZU6cJNhbBsj4O
+gxAsHtFFRnSf/AZi7cV4lNj9amBSNW7JOGK8PUgd2xjduEe2+T0WY/bTeWY2iR+
KjMBXCN6itX+yBVWg55t50LWoVFCoqL3Ge+wVb+KsvU7fX5Mis3JNfu0UVR0DShf
s32QJMCX3oirIUmxxz1Y1E+CbnXnfTBA6NthgA8RE7CKcv1q5YjnlED4IxhOiQdD
ttJtGryy2kIMF9NIAhVx78nTt6ZJvwtCo4Gk3kHAhBHBm+2nIksDjBhKWKbUcyba
m0yOn+u9ku4wDWbW9ij3hjZAxWHm5NNF49eJRn4CyEFc8BCu+jEG+WyyUOogpGUc
Tv8sLBFMhWAaqQ/A5VAHUEvrJN2OmVgJOd06OrRVDLUfFaPwIgczywnwAQjHblsn
Ic4pQt5gNYjMCh7mi1JclEtsgO5ofJkGVvGT9BuiMvlh5vAc6a5i0e/seyAQAqN5
KVDa7sTf376xtMV4n6A/kQDD0xYhjYxRoB6f6gl4+ZOGI3GEPStn74CXWb1kqaMB
eiKxyrH9yB1OXsRg6GQxPLDKye5LIVm6J5E+I7zIF8zkqAbByv4o8cTRKXUwCVlb
A3oBSfnH4mGQEUaZdM8lDyGg2XvR1Tx12Erfv4JlipbnO/OjP6B3btK4HWgpjEaW
IOxF5wganaLWVLKFQMghLVuccvw+tgTngJsBZ0knOAmvx91gwIUJ6QmpPglux5hs
T0Y0icIFxFzCQNmQh40ShErJD38Ry1J2reRwV0OGtbvbX/sI++eVAtCV3h4Maux6
soZx0/kpj608+tSOC6Ow5BAr1JzHpCFUim6sUZHcPf6LzIE11sqQATmEDSRhNEzA
Rl3mKWaT9AXl2xt4QbaaKNR04utolUeqzzBFBISHzJvBCWr87rmh/yeuwGHhBTK1
huKBrzUQO4//rrKMPtEkBiTQMyf3KyFQkMjP8xyW9tDXL+/u2AlHvA05Ss8ajcr1
4unmg3S474nUcir6T6R94RVAuHwnXl3GZMZhDUJtpQtZUYs4Ko30NZ69zjkWQNfH
UX77FOLxY2JGnALqdX5VCie7jzABGGKKZh+elSs4H526j67zu0Ld5pkmS1Xv4O6p
JGVlX45cPdhs9m6ySPjKXOS4XDdWj8zrxb4LslnPGzA1kY72A7OQ1PvjRFyGedxp
Y3vskoFPipBq/5n4JDVO6NsuoeL9fn20LynUUa1eIc3Vcr33vSgCwiRIaCpJsT/2
aXvSsQUAsjLInQyFZ7RZ8Pl9i4wo6Lu19IxmcxqQQS2s8pk5CyIvonIdG/V6MtEW
GJb8OwgipwpkZUrCSGvZKU38VY6PdVmbubV4nhmuN2pK3tOyRtsBeCCAYYt+FTKD
cNJ83OVVd5Q2uwvgAUkaDH9bDOoS1Ivw64HHuCGQqYW2NK9UfKQjf9E4sxHIpbaX
dBb17Z4iLMbOfr/N9kJtoMq6PJa31RuDS45yJn30gLsD9l7Qp02V9IAd1LV/65UP
tdhRDziUzTeWJkYq/VPXmKOki6GJjli0MmlrYV5WWI+EPrrFoxuG2DCKE8djBnmI
MvmK9ygpOgaw8KEdJMqq3OZxrkEclz5mYv6u6+IkFJ39T4ofGeMjkOTEGglY+sx4
JkBRMAjAxqDNrPFi3D0XteT9+bpjKCamf9KXy827iJf2btiMPZpDx2g8GSJxPg2Q
NSJ/2VnYgonJ1cWeRKLy2M2or7zp+Uj7QVG4tySVmA8XfPkyDEIn2mRT9sCE0bYQ
1fj+sD43NUy1ecxkdR5OmsOPF5MW+8Lko9ziPXEZnlW67KKnwBjlIIyTo6G7boTu
D+hdn+ZK5w3zXP+Bc3SDRpi9Eu9Ho6CMFmRJ6bCrenqVIgOXZ8+2jpsG5PS1e2by
mGDuIY8emMmqeHZc0aNClWRBWRhfZJv0XAuKZBDnyPd1tqiltnutJBixWNZVglgB
TWO/5aVZGo6XdUHhBkKrQRJVe7xKW/97E5neRjhOOqpx+fwKJOJJ7jVz/8WdYa5r
LIlhL3KWRaEnJ0eDSXRxFqLW9bk8LWiB9FXM2DbGUFLzE/AbkqWxr3Zcb/MFDkF1
0ZUQ+KYT30eN6ITm+O8mNAtsU+hCDRtu0HtfJUfAHSG5CDJ5rLfctU6DifANBJdo
LSH2+S1+O7G7e9SR+iBu35aqJbLuk8Lgn9jBU9mBVlifB8yJyBWSWE04gfVpAdD3
bDVwiM/T5JUygWi6KQk4wAU4e5s9/N5JdtHm5Dn9vwAfnQcv+ei3buu7V2zXfzMi
bnK3A224bOQbfvEDyHP5tJh+rVgSqfLZHUV1ERgGv1yK9cdwxqRUWtV9uyU8pOrs
E/E6v1QzG+WtKnzQZi3urKzPF1T76jcAVn7ZRb6cjEmAEefqkbt8JSQMCM4H8Pz1
XUAXBhWLafAf9WPSJdFasA==
`protect END_PROTECTED
