`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hbHKjdMv6pey40+LWTZgS3TSqIvpI/Z+o0420PHmUVRuNBZcM42X0KFxxMpWMBn2
TQIyfBETQwk6HwIeabH/cQziDs8V3HrdxmjLxD9JoWpTKYhn35XQa2AyUovQzOzY
LpXX/sMmzMfbROyk19/jre4QXlcUaAFzUvNAcX4LHNeBEip7mf47Scn9GCt5O6m8
/1TtqkTFeViPeJw1wLTA/excaLmFutCORQj+zxBBULsve/kPTH7bZF/8A/Yjpnl1
xZnWxqJNKMqiJCXa8KjVH05uIqg+1yQI0aRN6UZnXvT81cHl4zxSHhHHiexvg313
OhxfMBBDj8ATFa95docp5FmuPZF5QIM/RPhTavQ2xEVg1LEDpfhdqzE53kYG7W9V
O7Cq7VXZ1ttcClmxmweQ3gFI0slt5skogxZKu29SYASCoBZuV3H2ctPHmF3Gz0dK
tbHcvXKpu+oJjZAEQ0j9C/wn0yPAhoQUpSJVkzi1LjY+2Isp6DuYodKzEQ4hkHDH
bVmMUCWnZvHMOEUPPVbDD4CF46hJOreFEZVdY/B+pAmSlfVnCqWuXuYMHek1zJ7S
grPvweizY8cOrNB6QZiEF/86GxlWyrfSfK8vWiw9GhuQBy6pVUW33hNHjWxZFm9m
3WKCAFFDv01kz8BanWb2mncXZ1sRVYYuve9clQMM6L3cusdckeqwO1Vj2xLrsi1Y
UgfjI0dtCeQVN/NiXJY58vnhOk/aqoInjGMku8oL1cQPGHuago7BlkqdD+m8RzW5
39q0bm8b/SJMicwbNBtQMxDPHFj6EGPTKDCWIcWsBu2DXcIY5wcFwGIJcz/4Oljn
8IzH5LRVoxXjjh8LAmYmbljR5G7U7qS6OJb/kBxCzrvU0kSRKtb7FglCzeiuneLJ
jXrg8X5hYtihH6fR+b5uc07A8fQeR5N45OIkCckaYY1ga8R3pqQBn0H33M0M1E7l
1NQAtvzgkK4RHCCh6IPNA8FVK1XVswXMDLOmHxkFcO8FnSGhdOc+EFks6A4ZJJmU
`protect END_PROTECTED
