`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zbg8VEWkwLxnK30LlbMMmE1YSAhUGEmpDGoiVddVKGIR/DJr0dpHV1EbSyw4hLS8
rC9LL1erE6IViiWALfvMuhQZ1y9IV5fTAyJXAWgADHk+5+j4D+MhzIswCfvdMyus
+7qEONFCwS82FXK98YSh+nl1PGNX8OUUyRIPnYnYRc9J2LsT1ks5hq0481gkMunT
Wuq7ycIdvihNgaUZWZg8i3g2UCanuyOPupFnabCQrpDQRTjOlwgVSI8e8qK5PT7T
lKevvRW7RKEEFbGS8tbrJhceyrbyINvds32TJYrcXWFU6cDwdigoQhaQp8BAuZ8L
T8DWYhutU28RTlX27oohZAFJR9inXBEFd7dexLiTH6akJPJ5Z8wX0OhoX6W5voUZ
9fOiauNMwHvGD/6I/3QXF9rkxbBn7wfvL/rY/3Zm8PuzulhPH0ex1U13fkNvwDUn
ov+m+5+zLKqgDdrNcn1aGF3BK9MoXHOvS0mk0d8RNH+/WEFNBs8cUIlyiP5CJpl8
R1iTVRMExMNHgps33ZWf8cCFPPCSMNk67mOSdlydw0uEs4Z5m9+24M+0AQAyOmr3
td+7VfATxp1em93AGsKIJPy9MkD9D5HlQRPB3fORjECGA2h3sCfddipfAgtihWiX
91S875YrfDiU40RUTlv86J3U+GGzD+EgonC4XSpdNSnMoqmIqGSygOQYYCoMqhn0
OEMfcOJY/VltqW0fGoDa81HJsZi79pHbFgd/922iF9JlFSGTPwpvKZ/LwSmgWh3F
9NJGgb5xjsYF7snMrV8ZiUNlm27ca1feMyKXLMpdYT8=
`protect END_PROTECTED
