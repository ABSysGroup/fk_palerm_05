`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Izw5G6lMSZG/gC38HvGdFxEbiRvHssqVfMOD+qF3m5jYPkovRF3V7INPu1yuYTWL
P2/BFqW3ToSfkOQDPkeBH1tbQOwdtAUITx3m4jlts+YP1HwbRZFD40gN3t2zkJ7Z
fzZZ1YLQDeg18dulKNH6qaIFs3ClBYSxsMvvy5wFkDQF28JWjbBQ7vq692+e7tbh
18Fof/2bNUJaClzl/6jrrPdrnEolTYj7hhRO+bGLE75U7JBEwJsNDmE3wNF9+Ots
Yx5WSmOl5ptp5Os5X9X0CAnogQfic/oo3mKxjffAcZrnjrYEozP/gMoZ0n9GFyMf
tN45OugmPoYccoZmillw0TGWAid+AzDWbno0kvhbykb7Ds6kPVwq1LIcGNnFf/SH
T0p5LgZdChHKeKmsO0NcgiJweCWMPOhcSxw8UzgbLi0EBywyQeN2YC0YVLoq6HYm
`protect END_PROTECTED
