`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cuqda6NkAdld8ZVAWW/HYNSBtt0ZF9kGe0LYpDtjeo4eWju+a1b4rdaLdBn9fTsC
kga24YenVLF2X/qZ4EckVUGTUwxAFtzrXXarlxQLMseTmF7jSTyC1Zkx35DgNx2Z
LF5MvQ+Bs9b2LhxJokVzpSciQ4yVtVF3gQ9NNX0On8fQl7nAgywyeWrNuZPNZLQI
Qxo/eG1fHRHLdqpLcofYvC/r22QueE9jx9dJIQO/w0r7XrxGJb2eEgeQusBaFmbo
H+sgbAypMLgrlfSbryiQ9OuUksY+im8WO8kLDtcqWREe0lWBgZcG54Yf4cMlU6Rx
lfFTyvniwFXFoas9pm9RCv6A89KBy3OZ9xnAqV/WtbJX/JvdhCwrzm7I/x20/p8y
yGfBHl3LGi9m8HzQf1gT9F9lGGKxQOJDTuiNSf8bxIPiro4qHE60AnMOPfQFxnhY
bqRxpdiLuKGCqf0aVDGEF6bPJDYQCDs6qwVdUi4jHd5G7L/17yBEYPu2q24wkkIo
UUGnADPJKMbQhP/PwxNen+f5LWkba1BIpnO+P7s6v+Y=
`protect END_PROTECTED
