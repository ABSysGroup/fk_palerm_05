`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X0gg9VNRPX+d255Uq3rw7GrriHiY6STzfp2q1nG6rc0Ps9OUKTyunX+y7cIBRe0X
jW5HNgph1txVT2sNPTUMIl1wG7GAHCnkGpvxwJWXQm1z57I/B6uhrMbdofG16Gyp
NmQL/mzcMHy/sMAoFEgB13sRzOdkpDTtrZBKq415jqaoAH7Fqpajmj9TU7Gkfgw7
1znAPKS+LDsXy4E/MnUzaLzh1UL3RJIoDGKD6F5x/nv0yWYUnVp4qXt4hsSP/GLd
T6JLNSRAOicXyAfy9inNnlcymfleCuS9Z2k1NEjCAziH83UcvRfpNSULotJ3QZU/
HrJUzTiN8q7qW817Ksz/wiwaWsMqWghrWzEAxGRmBW+hH9qwGPoOg92/zxtogfTY
1YfmcEBP/A3MWlm+QP22REfR7cjJUkqU7ng7bQcpawCvwnpV3kDKAv3X2A6JN6Kw
/FaiAXukth9TfFOd47yDZ0gvLtfDBrUjB+hQSYhPBQcfaK8/zh6gauVvj28CkrtZ
2Pdut9ka+OYIHqFO0f9QhYRzMRanwlegZnSklnN6hjQnVMPeI+wWupe+MYNQKj6F
23G4cQu4aZaHfte7hMcP1ZhvKRqLebXaXKwvACyFNOtQoUKC9gS471cxfwdb/GYM
1q8/SkDk9P1BsT/DcQ1xGlX/Lfr/2nVK+SkAbHLCfSwzaGLRF0qGHWWUphNOrOyU
rTBVRhdVGuGCHKD4vhwmdO0qXqwi2dLtHiDS09+4FjsNtRSeInVac8O91Gf2JuQt
2Rj41xrL5U8o5vLkt+l8lQcpK4UZ7IMGVTuFr9zglVKx1Ntm20ES7Yu+4ER55Mtp
uF2uDqNWggkM5LKhdWTWBCqh52fZMepp8FVJDHzPN39wcug59DicIq+ov/+8lJyS
aMjhlT1r/P4kwbxXR9iOm/t/w2hUyEfShTa6W54QN1vn8DY9Ah/XpR+pZ1SDlDdo
`protect END_PROTECTED
