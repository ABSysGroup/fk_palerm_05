`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V8+Hc8aX7wo9lsr/DWdg3JbxtItqWK/Yn/+J6jRFTHzHIFXO+z/idyda82YbA8rc
XWUUNuKwWPVefQskK5rgdr9tyAvw97RHiALCoLnxJls3jaS0vSZiV+B/U8PxpwG4
mA5nX5zZ45T03aThU9HjYcQXpStcAq/04YZh7rWXwMP1qj950H8OfobFsXmlkLU8
B/848tF4Eepf/UnWB498i/4CJo9UbJyKD5vhNkfQprCLHTjzqJbYowp3O8QvpFsY
Js1g2IULADgFELeMrk06dgkgstgVf/rFCovrSwKSGBYXeCMGbPGzhcWAJYiAuHCF
NITFArG28i84ikaD5ZEdRg==
`protect END_PROTECTED
