`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
34fL3eNl5JTFuCr9v0tAt3acWoGI9+nRhaTQtaupKbdvGJJtuaoctUk6pKiMb1Uv
Hi83ZjXb+EaLGC91zC4T0QXZbTXa7wmQtpU5qj235DakORUp5H4xfC80+M7s7+2r
WKkaBgERUe1f0YAB4lC9+xxXvo14WEIqATQL6aH7JHikUc684Q2zUygOrxhlHlyr
Ae0XU01y0Euz5hnYJbp5NlFrb0BCcX/enq8kNHFJryB10jS7yvpGeeX8scgcFVRN
SXvvVbLxMTVz5LwI933JMqKTgwFHUn/JsUF4bgSNqqIOWDvoDnrdF9OZjhXzqfa7
ZjScIKswb6J2Ck/vy+lE/0vE3cYfViUlHwrN9vXKnjSTI27aBVuZ64IMta4A+k0i
qDxwNYuBoEo0Ext+yF8qZ5BocYlV32Jc+jw9yiU7tQN9zCuU8/N4JEJAZnR+51Ru
jPyVIJcK8jzub4YxbbYvnYVsws0VOaolRk0oenwZgQOd2WQ9ArR3jSf95i68flG7
01CwAvGDiymirqOVdKGX5bwzpvpwL6dh2B4PkLoO1VsZmahwnuSNbRSWQpLHp+tu
Kfczs+kOljsWE7qUlxeuK9owANfTfIefP9AOap4r884=
`protect END_PROTECTED
