`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
id9rK78sGwM/AezijXxqEtE2Sq2CRTnVjb3dkHZ+Xv2x73cposPUz53042QjWXAP
qk00zqbKCF/HNqQQLzKdkX+jKXwO1umkCM0q5PQnSf08mOJhD2NXPeo+R+1GQoYB
UaDu4Z8p3QAw8MwZjvAIQ/6qkSCLeYkqlEcHDsG+xbOhK89Vd5GiWP9zQBqP4EhJ
ZhWqYh1K5SBMz3dbzSl/UaKKkil9YxxE7t6MiK0KMQwvC/WgEIAVQHnDfnJB9WeO
azvHafyoL/WHyDAs9/w1WQ==
`protect END_PROTECTED
