`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
neIYIN64RRvFp7DUmOH5DM7eJddHIuWupURwBE4JCVrA2FHtyO++ppGDmF8qeE5Y
c/TikajiBO6Eg2VMaG9cpPIhuho5zzfWLLNixm3cNBSt5hXuJE0WS8ueRZXztezr
4jf7Uvm6FEAfVuNQjZKfxHwhW+0bbP/jmh3xNETS02nycdLz+B2Z7iQwBvw6hUQD
8AQKyO8up5eN1VwpUsqIqhcPiOxLuTuLkFvABah86f9yRR1lMpxhgQe6yXshDHTP
5QAXvPyE9vO5le5qFTUfJ5XWYab67ecfIs4mrQmFGE2hZpLgEIGBp0+nGpbDHhAH
rXtf6V9oGgCftySC1FQ21K1Y9FzORUvLh9GEdNU0ZUIh5wa+XTw7apypUEfpmuhK
NddKpx/w55eqWcbjDcY4ErD3JdpDhvM4bAKHz5wMLw7frVH62UFSrjTJfVk2McAI
cND8Yo5g7GfABI0zH+xvu6XjJlF4gKje91H2CUvqmIgUk6v0ofuX3R+oLeH7jP0q
VvLCYuPprbIviPuXsU0xrVRTcsvnb3+Bo2yDbSAzD+V0ItPRyNjwg8sevCq9lzjk
kpJ8AQ03cXOTXGOKMkEfSdnoEzxBenIV+5OOxe4FcmWgpQcufpUyeNgtVARQqXUD
cjkU9cGEEOrbZZW8NGztAAZiHQnkXWb1TKtsAlBHFluIljwVFEEq5i/kfyUrwx0l
yrjlAFshA8U71I13eCgFtm4ZsLLrUlALva/GjrifBluXiKum7goU6ZcJ6hpFYItV
Wa4DMn3O9US9ZbO1TW19JUKz9N6jnrgvF/Tjrn5TUlyA+W0IqcIDoMaBqCW69Rnc
JNCvJhezUDu7IiV4JjoHHDANgqgm6jjgS2f7nkhm2UehriHMYa35Fzq57MK8VR9K
tHJu5lUMiSTfF/zwsb4XKdEMeZR9zbPeugMJet//ynpCA0c1iJ7crepOY366NSnq
BNtmcctLWZuh9epbTQLrvPFyobu6IbUuhSgDVycOnIZCvJfWSvV+0O5Xovb6sBhl
+RTqA5x4vRVQkLk3vVWWp/9Ay1lMsOZg5w7vTBgJCg+06d7l3zYl1x+u1qU8BR40
J46WM1fgyFjtxAzHRfltUI354nJrvJH8Az5SGOs3MKmtxMECEzzWYx52OYbIjbnL
`protect END_PROTECTED
