`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+mu7qLMzHXvVKY1llS/ic4MRtZCVK9VqCGBZMimJL16+lRjMGfGBRqScpcfYzz2W
7WWHgiQmPvS0eoSAy8o6TIdemDg8FAtDCDoJRCxWupdrWDqdABy39YMBChn+XCvd
IYaHcq4b67QjDLl5IF1iie0qbRZ3TuGinYXojuIUZBfpcHpBQOQ5Jb79W2vpoL0+
wr3a5jWvU93Sl03Jb5hKODE8fiVLVfYPatK38TxyYMoEE8YShFuK2ycDYZcr/dzW
Qbf3XpRdI9zbniWJi2f31E7p8nQL3eyszZfQ9OU4gQkGXJ05E9kHhj6MiiFCNB9m
ML4CGDCDB/Ayxc3tAFHSHU4P6q93vQ93cn23P2tOPzjn26cB/mvbzDEJkm313fM8
D77YUZnm7sxtQNLvBwCdeJJcWeDXzDdTbNeux+gbjajJT5akBXw9qImmOMEvVA2m
C6HIzVD4mpTDVmGwVnPKOs4wMVgh9cF01xy8WipKzqK4ATlFq3LhLNIEy8UYqIMj
yLOWm63vWBZNJp1JVoEHSGgiq2tceIP3FUiotG++F/E2nBQ+a7/gwZfwL3uqBVqq
4mdHGMLCNDpxDgmRC1SyS4zlatFOUilzM0xyZUQOv/RpLh6tKI+iUXOOSR52x6Qw
8OJYXsJDFYuOkmCpArZ1qRDa0DuwJkkvNWj3NEE3W4dM4ltZRN5Zjzo8lFaHJ1Kk
jDYZeU/ZxLhJhcR9kZ10S/sm+l3nhQLwz+QYqczYk7LFBeqgfGnumuGgd0mOmTqn
MPZ/CtIHYJfSuF5bDWv5DQ==
`protect END_PROTECTED
