`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1x8+Ygt/ayQ7qB6cFjIq/5qallomjhTyS12UMbP0FJP/+Jqr1nuHG6oTOtkvXrsG
JCvx5wmgRaR3tVK/quJIud5TSopW2MFYg85OZxEsckVlrYbZo3lTQfjkpjX1PY4L
oIITGwzqWsBWhZ7kWd/2Py96xbIidi2h2g0dAokefcs0LbuFk7E/MBUGy6wQTZUV
qKAeMfJS7YCASwPrDdKNFBMnxT7pQPDMDSD1m9IX7hRZZ7k9BbW8QGHLerfkaNrs
0tljsb+KEDspq+BVdO7S2bj+AssRPOICrWPeSEfgJ916zdrrwJbrw5WYWJh3JlCV
TRpMHzAJhrxkhx4fzby2G0ilbmMRBY1Sj5cl9xwtFOGh3o/0dLCUt8o/HQWfB9js
1fLC/hlA77D/eGrGYqnRgU0pslZVLZBSGfCr1VjfE0cDtQR/U/D5ylBBr4zPV9Fx
9rriA3MCS13Nn/dJmFnoZnZVdsLffJcuiDkqVyCiqirUu+5Y9WnfDcZrBIoI6FcV
5//STJ+BNEMKh9IH2bLhIPFQ1hg8uqlTwj4fcRERhK08pmDZvtuekR/Cu74D1Oez
3QHXJ5uHK8XNDt2pkdbTDcJAImmYuqQGsTUNWGe/n0UbKa2AnPf9L4raEhuAp/ws
Ac2CuUkc22BbVNSyyI3RIiLopHVesJSgz255xkh95ATy8bZJpILYBqZ1EzLLBdrX
xDqw3wuQNNrs5VPkKJvXKgPr99JmY8DeKDgtcwca6fFW++RFoU0Zxv4g7uapTtdL
9dROImgd3u7jI511SrfPLEurw/9NYRip6xDBm+KR5YIcPugh8pOWm+UKJWJFBpoK
Wl3c03/pwt1Qd7AjNOdX7dP8kHl4jyqxQDPXO6CTzStIg73O9d6ji5MqTkFHiyzL
KIJrgrfK6BwDiJGjQXrpsX8y1tLO2ZleaDCqzSZ/5c+WDD55BmhoyYJPNnAO4YEZ
h3v9TIf8NkMpZ1DVZCJegHKyOT9an6CkZfSZ+W9qqAWm7OsPHR2JoUwbN7dkst4y
MUjwOiA4jKMRON7sq1XRJ7fzVpxPNtZWGKp4V+ToCp42G8byprnJgB+h9LWx8NRS
J6ZHBqiVjmMokWwANPsRP8AHW0NUkfK1JGUE4icfHCJvlmzlEbMG4k2PoaSGsjHI
wP2MXbXGi6S5oYBJHMVGzXV9MbhNjtGLMgcN0WoHd9mpdZhJpFQrZSf9sRiGrwRB
lOftIXJs5/jgDGfXvi8r7W/jH+YzDCdw1yk3Z+ELTTxY5+7G5twGNuiSTC1FH2fr
Z2ksMiR2/IUAHSQeoURhl2FVEE5lY9ZniyCKdyfOaWk9boSe7Yj8V/oRA9Ux6O1z
dT3nsNRFX4UpPD9evAbThLJzUObzoeb1+wkIvwYqLTk3xcMpAoY5nwc+rz5pC/pu
GG3sIxrWajw+bTA9vqrTYChwDy3EXn2fRE7qtXhtHWGTuoozM6tsYohLklzcsWbQ
hIUVHCfmHiqJk2IYfjoxmTygGaZth29sLOWCxtIWxyJmzMnkVa4wyvwbXqYUVf17
4ULswKVspt4bSBjBj08h9GHiI4CFfWaHoBuKET7AzUtbxxK7QDDUJGVCiwxCsiG/
s1+HfDPT/1Z3wt3Um4wXS7AHRH/asu5aejGk6zC5iJVQJ3OjAqRN6lKFbiz5+Ex+
ZN2+CYXTHl1g2WR8T+vuwUSlAMLgrdN7aOSr2/TKrD0TtYOohIoSSB2enlSWKN7x
sl3eeocC9IXVwRe13bM0de7M5GPKahmoiFdq2Fi1S7arMpWyysu1YaqpWoyjqEI3
6jwJKMqA5Pkgv8wGRWrbr7Zgyjx/URq5JAzLhn6YvmvO49piigW+JfBT9/gtljHo
SPy7g0MyYBluk+tpPWFrqHe5tJSDeNBqv8+fi9NiDBppcUBTmoq3wzyZMuYvhedK
9RN9jDDuS8QGI5CbsEbGhPV5P8nxCsAFSFg4aE7cJWjWoahty0cXLWq8PjaaFjj5
hed2eH/P50aeBup6Tfi+xsD5ouiZnqIjk3kM03tdemlgEyVscWC5E0LJWoevSq0j
iCuVwT9hmBu2krmcEX2Yp/LiYrVEow3x8U3/6RHknGv4Jj6G4NST7EaUiFRFVPVL
A0uxAVYyhn+WpEImy4d3ePsDTvwpBQ5OOJX0eC9KxvzfNbYZsrSveMK5gepqBE9w
DvdpuMeWvC1NpBW4AkCNVhk9eT0Kz+1VjCNR/vVoblDoxUNGWF5vEn07lqulnWkp
yTnqErApI2BCZWwbGqUNaSYNvMQik3gNEfeY5I34YzToJn3zRJNeSpyFTGDdhuKZ
CVnFRCxpjgJUZHDErLX5igKPPZfrKonKszEl+5hQsX7PVTXYPZosDfk8gIzWXoqO
EDSJcuraA0Wumr+rTA/FcbGTkkXAMQAkIOkC42RxgULAAKm8QWqfycw5c0PDCJ40
YLIG5mg1JYG5cc4IZUefZunm00n5YdPe/75NRD9/USb2EJRIVPs2dgw7KGgpMkbp
vevzFDkNgFoNTQzhZ7XX1yLLn4oXaEEVZBolXXuksOPoBM8wtQlBccs/Id8QWOJb
ABjV80BKVaMD5etjUcB4ZQ==
`protect END_PROTECTED
