`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9QbKUAd1H9fJ4B7ErzSeTG6Y+yXxSUkUlR/yAD7518FFGkXrBl6LUHQ98flxiDH+
kRzjRzb3tF23S/HXk9hKkEvUCFV+lQ8lJef+b4ucUGJqra/Zsi29wbeAxZm6ABtN
atoD7O/ZMitmfVYDueGQpLfPNHiarAHQl7Nbv92PXlVoYp6ZzgtieXtvKWwezVfQ
Y+Rm8LuZSPdjAPiArhWBQpYrrfA1/7zEb1n4svKSWPfYBaOCrn8EHXjiMgSGeyun
v7lXTFoWegAM+nOER2ggmKVLRiIgf54AO/d2EBpbWuep1eIWAksQAT32tvvZgeXy
XGiVAGSqyUnyCSh+FyeGznjM/PQO6DPnbaYDHtMxdF3J2Z5KGuF1DbnYEM8+axyP
wjtV/D6IaAhPFfEQoYc+bv/5FejuydU0AelICMfaM++FfitXnrqqqyU5Rx130aLp
px4+h3wLLoiWqkJjxc3tE1L6Son7dJO5wmdt07ey/xrEoM569amsUZB65Zea1WxS
HFTYLITrA6ZQLsCLdMjXq3hvlYeVNky09qmN1QHSwB933agJ5BUlO9dDA+190Rms
t1t13/0FC/g5ZplJ8/yWmEyILJY1qsNQheyuYs0vQRJBGi7t8rCHXh+1Nknu7oXT
Jdgn3S7GHrrN6eYsl6xzbiOw8X+BB1ZNY8OGThvq2/NOWbVsTiYdaOJ0UFHQdEtg
8E8B5gwArMis2HPShOXS3og/B5wXF4zOMEaTBEDz2qGDBS4lFKD6axUvly32igy0
mnCv2WfA2/Tgk1ApwWphCb4MAU7/FYvovnp+k/dkNOr18zipDqd5ljfe8UD2FGoq
519MNf2S8x0pyjwwLOa1No0k03EfwRCwjf+IA+YMcUvc+BQEgwWdF5W7357kmDtU
N/oSpZ2wnAITeUzM6qWrNsLAY+6al5hG5hGyiDXZbiJkJNfn4mn+7freyZwo9i35
lAABCsW6o0t4EaL+p4VnbqbRL/95LogT4Me4PLIciQyJSq3EGiNp+tDB1M79LwX3
uaTBdKfgeGwWWUBklvJ3/XkMkxLK8NrDzCcaq12dP+DEFumxRG8zvq5HTLMSUllm
UYo6cOfJoGuNAGErOUOK2242bFFkWcRVMOjMk5+R6huc8uZQr5kocV0/ilbKVw/0
7eSWIHTvGRnOMfzHUUVsr0YBcxqwusUC0Ee8TTi0J0JTeCNCS2xPig11mFb72yrc
2BubNQOzCn4PKlIEnOjEHdHuHa3E25mBjFKWKoZAHjpO9e37vXpk3qNFpoeJeW9t
Rvh+R/b77PV9n4XQz/uWjVme20lBsWVyJzWmQNP7/2IczrqcWiXB6q+kMq/4uy0+
JxneM5U91K2CaRXv7VqtRKEnmmu6yE8Ry8faTlNQK6KDeDJYrXQRuF/gagymjYAf
+EJFs59HHPif8cVpI4qcHqLdyGaF8CrQtbE9+iQR/KJfmnOBet+bRxeyBH99snjJ
HjmcClK5W7UFnrX2jCuSbomXbe6FajHa89Gu0n7/OQzRMn/yvXhpRYeV2XiaoX43
RGjdigoOx+5wVJBzjAGH9ohy3+lapxjqVjqf71F7x0sKua0qDMTat2epxokFspPp
Cx7rehJYbWPB6cQX0labiuwIBAQtsV854u7DDeQOz9zkGAfGYGFq+kVycztv30gC
xinPrm1eCmKhFVJJ4QiVcQJpfToN0vVNDI+VSXmFFqopx8Jn0gJoWT0rRzL4Z2ex
5mVVcj/jETkwiC8crSG5VhDxnxI7JVgi+BIFUytVQ8ZZciV/eTs6q6hK/wD0Pn1V
KKoSSMdHMxowxvvcqRrpUb0Iozur7bTsKTDSl08/X41nW0c3QVxkw7b+k7Up49L+
NK0jlFTERVo02IASWR6qcfcIH7srD0XHzWIDQBLq8Zh/FZfelNks/MAr+HkzZE0J
9nCY/EnTlXQa3G19HYy8ggPDHQuwLDHK3fPXmaKoQlPAupg5dzW7QCJF7/xw3zBD
lUe0lQV4iDx+aJqqgdBR8VMdEF8UAqIYwjrm+BtCvhdkv5KuBWYt8lx8cr7DLb9I
XP/EaH3u5ML+nD92pyZzR0MaX5nv8hxiAltnBDRoSP4rne2nIu4exAHZ67Z3uMwH
spX7jXHyxrltNgEJxVgYtUdPjqnjae8hFjgVn1ceBmz6F+e+7KMVYCJxmyvZbVOb
NmNgYAy519npLWfpZrwOZAWtb+V+A3tuIKr8nHcBUqSjklye0bW/3p8sLzvRTNr4
0DrjLKJxWVqnVsAOtYpf3Fq76d+JOcR5yXuuB+K5U2sEUKwRnV8tUIB16+qxwwk9
JxuEHoQ2Jqfj/miKeZMXcXVC+OIXT6187DHVLWbS36/hd/0icbsuhIR40gBTnA4K
9/AAWZDsjcH4AQdnNNaIZ8JyrJOuwVGC+BURjMf+SjQ=
`protect END_PROTECTED
