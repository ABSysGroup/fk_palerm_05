`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xShKDtWxRaCGhgmltV5asT7dppoNT8KF4rcGnM8bUonPsNBxuQY4O/c5nv1iCyQF
kDIvnlknn1XxT4+p7QAiBjmWZGtTbBEjrGxSQreJLdtsX1EGV4gMRFaUAewIkUVg
RhwzljXw4YQWS3+C3lzZyh8200JF2YzGSfdn+SRNqaAkTHx2HOo4A1nd6EJ5TifK
jI3vR7wESJo6GkbYA44h7eBWe7knJ0WlYLauYzjFx4gLssrs7/6sli3bSA53LAh1
ygTL+SiLAL8B7YvMILWmcYYbYnBkmJb0TvKstbns+9mhi2veTF3d9B2TBS2w4AkT
og+Kv3HyQ+Nr4U7k1kKIwWxki4JBz3z1xk/S4Txo0PAe0kAsG89dA7Wq+jrHhYmP
xbf0f0AU4BAMN+ClBzxTxIhnu2LYAnjoaW2+Abh7Q3QanbLZpUvCM7y0oG3jic2G
0s/alH9wiXBhlJdEGjR1JCtggt7ItNNZ9OYs7qQ7mDI+34OqNr9Hx+dAga1iXv/w
7uTrU7puRZuKsnYlp7rok1cq9Cm6/Xpe4Ti3KUJg+B/HC+gi3pR77pBCRbl6BF1E
I0liHSdLAx7AZqYoPiMi9x735gcDlc74APV1yOiguWHc2C/zsK2C/iCT3xl0++Jq
/dbt/FJAc2c/16OamMCJ64CYGLdjIue1+CYIvTlYqXn7hj93lQlsj5C14/FKgSdt
+xaunbAIGMbfIHa4HEzlOFWYWgk0PB4L0Qwz+LsD0uxoxJfXhkhLCaXnkJjnhB+U
nBIk0Df4IkAJuvCWEs9GCGB1hf7sRsh6pkmNniy4A1Pe/X8VvBPJml3HcklBXf+0
tj3278PWpOyQkLz/crmiIcd8cqDLhosXpNhKNkEKquCdjNJigAsiTAm9SxUAo0JV
Q2KgExAID03kFLpIFqeoO+H0RGgIsf2vWyEzCe1boYY6l+wcOLrIm5SuE6l+tMsp
XIXh1Aofw5SLqApCqEIrgppizlni6ngpx81YejZDI/XNgB0Vd2iYbe7QVyobj5V9
imLWLJwO6yBP/UxFojrQIa8GgLEEth+zDPoam7JHaeCYYlc/6YKQpR2yfK8qVxNK
yvE4DnHa/1dOIjpjEs8Jq6jb9TAgHAdqr5qT4G0omSdL77oUS6r0tockn2+Oi0v8
XTNkmd/UjW59PCqKSQ0OnWvfAznkgmPCeXf3POr+tN1CygntRbPhR67QBNXutvUG
DLt3ILo50KibX1qWnWwk+QDmkE9rSojo+ufYC4BBNXEgDlvkTE8W0CLiwbBMivAI
uExAgJxoGd96gHjgGUBBY+8CpCnXSW+qHW+HGJP0g0DvwT+TxCC3TFaXB3gRQq5s
kRQPlcPZIqlDRMUHgQ8eY4X6GR7Qvom+sYITqcqYkN/taZ9OgboABd3+ZlVB6Cci
3sPT/C51OTk+BbCr8YNAFqiLAybdW9B6yS66OMaWlgRdiXHAikLBHXT8VK/kkGpb
QewFLdC0RMlmQhkKsCOv5i6SO1wRw/cjwFCVmNDktuzvSrn0csnB2JIu4ZWSYDN5
lCXpoEiHhWVQ6WvkyRSEtkJ4xt24yHiSLfMiSNzUm/HDlNZtvygMEQqKYM/zibfO
M0OmWB95A093NFOE7oBwuN76xBeSvE4Bf3p4J5zPZ1jGKmcoWKjTyzK1df0PdM6v
RHhYGvB6wQ4ccxAlPtHws8y7MaRpW+wxEz/g1P578S+G2kEqNaofEjx1uXW/Thtk
VaL+iIcp2X+WcA2kArrtTBDZuuZwgNspLIQ+pXFK6blqMpINkMEyVg0tpmJPWcRb
Fgv/NXo0SLG/SYaY0hMBoFYsmZj89ft7c5j9HgDThYQXeaMG3JIzXKcD6suFsyne
yC3gQbzmGOMpavdHzyJtgy8v/z+ck4e3sj7XiJE6t6cbCVBCru1gETeQm7ZjyZWQ
N+DU1a3Htao6eoIui+N/H2d4j+ITax2UWXzWvmlfpvswHQ3gz2sUJspt464zPbaV
0mJ2Re63byOngOjf/nCsRe0LPQz+qa9zqnHOo7Jh/iRBL7mNA9TLhyNvuIxvgXfi
zlfslNssIdeX69wGo+Aajbi0PE3BmSqtW6oLTyxEemcNptL50WBBgZbSwCSNw/D9
sh3lqMmEFPOKHYzxDN3LrCFQjaG/bD0Uqj481teYarOXMB0hx6ZRbUwPIhYQmNqC
cF8L665AYJPA6Eg0XP0LR2KGIWh3MUKn+WHEXIkKEaJbMMzKLGrg6CIbfFqisFrl
bgccMvZ54VS6L40gnbePVm3cXjbj9S37EWet2WXYULRrAg4dovWgWBiAtG+oulN5
irpZxzppR7P2KrH03bsAso6bc9kEfmwH8T5TgxEqjk+Y5NCG0EFmil/kNDLOJrFk
VwW0dA5c/x//Vn9pQekJZrs2TiG3t/mEeKjCRvY0bo6Bt367sRcElbDVIUviBbA/
aTgReQxKVO5YJbiDndu/YuCwVa+XekisVAw4vVPjNZur6fGhatqIxVrmZ9AHG6r9
lWHZVgxppPNcborNuoWRxQ==
`protect END_PROTECTED
