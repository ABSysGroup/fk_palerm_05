`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nh+JEqdZRGme8c2Yk4vovI3vFBdrxrk1pUc9Z99uvhGH8qlD2TbG63i9vix0Buvn
c8PtfSoe17x0pdMxbkrdGCnpDwQu/k7iszTmcoBQ9Yst9zTA2SHswaBEAGsf+Chb
0ioW+s9rR1MwahYOBLrX50AP/PfoQixrLFbX5Mxx33/9RVOUiVJYtj/FtOoajEfC
4mEq6I1zVuwzVrreSl1SAN8GqBTaeAQlHywcbLTSzLiV/z42jNVlaQTpU3l0OUlx
RLFE69ZWCoPUZDckEbeCyQ==
`protect END_PROTECTED
