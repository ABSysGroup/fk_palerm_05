`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NtPKDm4vK0G2i3jhv4NR6+fiklJ7nOSvhIkrOiDw5c5MyoIqoPJ+TX1MgLOjg2G8
gIrXRukn5hc11fw6ffAapVUb2wB7W2GX5vt5S76hhXDTNC4A8kg32NbKX4xhUgxk
XK3NoMyzYK2y5f2LSpsjWDwI4mRTTmRcug/jal6HfCd6aymKX1IY3uLH0aSpU1Eh
C+v5HfsXU+FTBzd2Gje22ejdkIo0g4nTH3CumD04vk6KsvAbb4Z/zBruYXaoOTl5
TX3Te6PnqQnfQ4rYm1vK3mqGlrKr7WIgVkXhojK4wVPaCcqYfKDxX1OVJgpnDPe/
dwqZfV0C8kKROs9yJ/RYYQVgRcgWbCDD/hAdGIoxQCY/XcdkGvOg4ee5f+TiSbLw
L9rSKlSMDt5lXrTt7f7RvaJ5Xg6Tt8tGvMDPOin5tIZLuQ0MorlUK6cvoMShylFj
l97JDrYpDvbTo7OM0TOwtGIPBqKBBomc/t4SG2dULDBx+pvw+2/xSluqm8ZINVsF
46AxdF++AUNjwGZLSQktyWiYB5/Bx14thkaLvYVsVNhbbc5RSzZveOBZtqYM5bp6
fPu65BkgE0QsEIpvZnOuAajYEE8AXMuV68fZiYOVfXwhnu8d5JJ272BPorPVc/7n
rnyGXJsUI1Eh2U4UG18AE+TMLBksXGj/2ULC0cZ3gpuXMjDOWc0N8cTzUJPMmZQa
Z0LQzZp+CXJgfAgaSHVgOxNvqaZsErqPjzYOByC5Ua3qKtuDwZw8fooaP72H7hEO
yQoY4FrTpOnVtYMvYmpRJKh/onM2v0hZvmuSzcD8HfibC/9Nva/AVHE67RbVbTU3
Jda/vJsm70Rd/1tkddM/QjSQH6aSHPjLwIJfS9J8UHziwjJ1RvafE4sBN23DW6TJ
WAkHqEbgHeBNBSmycoAS/4Oa0Uh9o363+s3c1NSqICt7QVyBsX7ovhFouOYNHvh7
3uDAQiNfVayMMLpnDdeyQXWJh/HHX4jh3fEkETMJb3PwUF+fGlOBcukPXwl08jBs
zwmeAIjKxtgvA8ZwryhCckrwLy0QWz50CVcuOvOEwb6gzRqL6ry/tYf4SGcIJqLF
kpKa+yLv4WlmXa/WZt4E1K6JsVop85yLhwtgEC2Bf+G2EXxsq9Q6yLEgH05BS6mD
boeto/nKIwlve4ve+7EtXMSS3k06uPy9IxIudv+WfoyYEeAabp+APPXWC8w/nEPZ
eDuL5ucmlC9b1VKwxlIfLIwSs1smxz6QZWED7r011/x//S+NY5pk7VN2Bj9wviQL
uufVu5JMTpL99/VipIGsKtcs5GoRjX8OwrKyMafe593HxdCdWpTkiQXCY6M6QeqX
JHTFlxnftJKeVITI7CHRktDsJF3X2FmZ10fZq+iZZYD5LS7BPyIuNT6QWJvFSyDB
uKiyrbiOAO2LlhLdzoC6XymhgxM43V6/63MN1Dm3x6TncjKDNNZtkn2xvoGhOW8d
VarhDV+FjfTIwmJXJ2/0EtUGsfNUz6C/p0cD5HjVyaNRPENzmeWR/T45SfZlmsLB
abId9KxA7FBBr57ZUQHyguqwEAiTjncpkQYv1I1QgQ8NV1pLVn/5mq/jfNIxS67E
9thYCtGrzMzcfOI/skFR/MPwRAm9khFxAqKUSeybI05NejudpMYzLO+8dxLA9ICx
3KC70Q53nVWmvDls2GQTQZSgzBf1Hu8UV5yaV9n/QFhXM2pDKLCH+5BIucgWml6r
RrBk4MFCjoZ1yz/HSCnIjAaBEwEqIAeP6JuYOQLKVnNRYaM4A4Z2y2+rFmAd7isU
JQEG7ssofkEO9ROU9v/XWrSEk2h+2WoSjjPQJx4xH9SvLfnlky6FXMXwW83YMWln
IY4pdUXpwzgqRFXqxPiY2cmXt6c21SIQK4evmUqYBHqOZJ91CN4fPp1dL4p3ZNaA
ZxjXAi4fdhV0zEgPYpXoGvDmiIioxdBFITNiECFiXKc8VWthybIlo+EAYz/6v/pZ
ZRuxwR2scTTvPNJx1+3UwTqDQv92BjXNFEu7oBR0l97LRglLidZUYN6WKqBMBDmo
KYEQYe0TVOlVHjzt1KzgjJZucvlZzLVSFedSo/N3dEFuShi3iGNzKvxXV0ARkLw/
2tsOxuyjmIgYewScqLpP/UMJeTCA1xhB+bQDDrWzg3MuYwsQke6RUEsb+0BT1wZQ
VRetkaG9VLum8e5fmGMvAStdJJCw3S4e6JKXPSt5FNaOP0xb6WVb/9VB3ahY48+C
Rs6v5MqN+DFwb3HW6zUeh1fJRjHRnyZ0RZPW9rUXbQiMGmpQbEbhyZ86nflfXqNG
dKJ6GaQZ8DDbtlIapBNcoeksyuHTHE9mkkxIQiayLynWRBJt8bw4H3LsZDLYCVhf
KvfbuAIy86iWIwJTGFZRw9LWjpHaQrA6/CU7KfL0acVEjx3r8QarPY8CPJeRMI38
bXqLLzrmQEfjCbsYNHnIZu5U2B5r5aMXexQ5f25wY/PIpks5EM5VWUTU7IckpE9Z
emepH7/sc1NzJ2k6UZ7ldsStfUC/zNt09c4n3AqrzPwfaHeGGDuvyh9KDx1EmtEC
fvQHTZcvznK5Pr63rtJduGloV104Cu3q8rEtTWromVX3LC0wg4iiPyC2n/PxMDFH
eCZtH2H4aEk17NDOyrjhhhWXcASi+9icMqT3fPzVOratFg2a5II58o9bLkI6cfGI
6BrbzEOdGQJxuV+wcBqV/YrNAVHlnsZWPDE1eZRMLJK9hrI58W5Zuo/ijPDUupjW
YlmcHXumQyYVN5RCYDcnEluDdPJGHRfEM2xl+Alo/AzcvGw2TP23z/2Yzgp7tqnW
Tr0oDstCKwvcP5zVygriSmPo+hEpJVpYsj3FLizyX7tDSPRh/0HGZCz9+7sbqvFv
zxOuOCMf3lGUUcbnYfXMG5yjLBELSWpsDcEWxZ6wj7SHQCvFctqEYiHZL2lV9u1g
EPgud7C2N8gsXNKy7LL57cZQpeWXMlndxuvlnrUgR5pe3pmxsRbUTh3yn+UXNPbZ
Rn+Hw82MMQ74EIp6jA5lWs0g0RjYLINpuFJO0ompdOcSd3ulJiDYYKzgn6/yFn+Z
FkEZ5UUSRGKfTEBZCUL1QGJashPG2EQVkn1SwUFsmfTL9FhT38u69C8v/MRQKM+n
u1rAhDZcoviBhoR7UkBykS0NYP7IiCIve5ozRcwQNzkCp6lxgF3whrW7OodxSFWQ
zXuazRjpKYd9S0/4/Gr+XOZhahzu1bo5BHR27WG31EeSsUZRlaHzTWKp0ylffvAt
xy2NdYOWlPPYnSh8TenqXCVVUFahud0/nV/bt+Vqg6yIftQ9QBZQz+Fs+Bc/D8Qy
94rB9OY7RMRT/oRggmmCFpDwZ5HcOGRlTZyoJCmsqd6kUVQWoe9JJqKvPGNk2wib
Dlo3dQJ3zueuVbqSChAP6bnOaSFS8IRiaIpU4rN4N6CT5oKPuHnw72ZdU/Rnji9c
lPbar8OhPpDYK5KRQEtGbw==
`protect END_PROTECTED
