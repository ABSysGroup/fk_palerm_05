`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GNKUdjeahKIJZvLP/YaGJXXCDke7iM9397ohYmGsUPuFiMsnoDtBVLARVA9JjlMy
qrHb7qa8EWLe88E+Z4J14b0/jM56OC7P8KQWtg8+yRsispMCJkcrmllCfuvQ7oTU
iRO/RWb7cNMkjJ/kT2TM/IM9D8ABCBaCViUjxv4W+fu/eRR8RukDsgoJlpyoBnbv
TVHLgh66rr5Ee+X7rwdw4TtdsakXlPJGp+DvP5rWwurgJyzuYYsNn7BPnWBJi2gz
24LVkh3TybN+bYf1HeoBify++tCxDnGIoH+u6tetrjf8a0VWviPOjySYx+e/WPiK
tGhz8bcQVR9ENZkM3d3bpzIMAQ1c0fzImXp8RdEfw7WlvdWTMTx6x4GM0nfArzyX
`protect END_PROTECTED
