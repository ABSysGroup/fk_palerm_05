`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jKQYhcsdz9Ee0JBgULEhrqVGz+pq6y9SLh0J5SVTOcVHTDjoJ30VNbxiJdsI8TyI
QnD1c0icUNefCcnDHwMF2lOeZ+Ptnjq7L0XKdD+QUS9YC6IAeEaYv8kR11lG/d5b
E59RW6FYBpk676TAEsBFDEZXtueKjWAHhURDZWRI8tsWpbS09MA+iVXGWS7SShvK
N/EjLMs3g87eeqV9kbXKLEC2w2BYLTQ7R84Od6NXj4cfu/3L30Upng640wDZwKrG
vaytbo4r+62Iil8r+XBt53pKuQlyk3BCC1DsVXW48aht69gYGRNA7I9ic0ckUS4/
3+tzSxGDNq35nes2QQnzW+0kU4PZPxfNL+BYLmoPqh+6qXLgP9ROT7tVl13104j2
MY2oe8XWvLl6p/eUb1jdv6QqHeMWbTFyEw9hC1yNeuSME9qkmapHSH7sk6fNMmxG
gL9ufGpaXcjLVyf5WFtNx3CeuhiJ2SnvQfNBJTIVlI5TkIuY0nLizqSu9D32PFgq
vtbWnL7vf2CKsaOcVXg4c7SgrV8Z7zGP5akSeC8CSXLKqHfUi1ok6MJWsH6Sik51
X6d8ZFgh0B/kv/ij+Wtzg7xw10Hj7y2kwVzWAvVQIaANFnYbeKgLbI51sdr5pC9U
AF+pG/Uj5tnAaA2ca5kvKQrDxAjZ4nRpaoqndOedu7P1N2arvOm4jW4tHABoVF2q
Kok3pR1xttKvJ30WCtTQL6Dh/E/Ib5E2PUDobWh8vE2V8BBy9S2CX7be1LrjBYrw
vfHdZQHFWUDvVYj5HimM+g==
`protect END_PROTECTED
