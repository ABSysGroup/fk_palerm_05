`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
brMWg6f42zNZAUwKE6wHe+UqS2G7L51DX1+DkRmSjbsaGe5iV3vnGLl2q9xJESS9
xS4BZBA9W+UnvbtDDJoWCD3BwqOVMatkDXOl9gQhe9otq5SazS5iaF4u+vPXwiME
1qMpiJOcau1YOpu7BYjQyVsSY7a//XZ3mBoywzGegfEKzZ9FXc+r0llaemuC1bmU
NsoqiZ2smoVklGeQ4Psju5ObZ/PXGBFDT++r57Tz4Sma+uMHUPRNBnoeG03J/OSk
n/jAM3ZHKt/O0KQvkPDnGxNivccu/Wl7YfvpAWM7yKBFHbKB2NxXouqeYqEMhvJR
CApJS74zIRqDmW9PkWmv68pHyxdaS1CbExf/11fmpJEP2I7hH+p3cXNaKHtWj/Jy
mzvABBNyAR1sO7d9xv9dRxt2QJOvv58jJJs0GphZZ8uYC2f9xnlMwTBy+O3cAyX1
Y3BJDGwNR1xYnpFqPcCKkF5GzW/6ULK3ATvwuH7DbGaWNt0lFru+cAs7VZ1/I1+7
8463dkTMjMm8GRbO6jhUeLzbGtoC27Scq/LnpobU2gFD0B6gUMCBM+BHq7Mozi/E
co3NRpPzhxGpoceHTbzGOqB6W2InJCVp/a59Fed1NfmWDG0pUx9pbC6XNTKrT2WQ
yTMT9tAyYV7dwUzd5qW84Gs4Pyug+Efg5d/fNJn3p5g=
`protect END_PROTECTED
