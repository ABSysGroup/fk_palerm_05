`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tXQ7d3BIyzlWv61pcOszhPcegL++3tH6/yVC02tV9WD+uzAyv9WjSn3sNxhEhTVg
8YaA9wbhtpwPM4CDaqwOB1glT+gy4AgKUcW4jLgp0FkDh1+WMcp1SDqS0pYELvl/
VdVI2M+AWudo+gRhvcf96GoWG7/WE8uqV9yBigYB/ZIFFswu53unTpDQP3/R75RD
RdGW0CyXYjYLXQtplKWjOfgIE7QsosiutLqkN+VqKLR5Z7y9Hdp65/fDGMzGiA3O
SaQsI83AueAJ9pyqBqusFQ71OOgdf6+nOGjEWSVj4HPCe3zQOQvheU9jGTXeKJ9M
4mw6BS8o/X/869r8XtQjVQ==
`protect END_PROTECTED
