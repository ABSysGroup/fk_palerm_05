`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
omq8R1A375YEZbiXZkwCORa/XU37co3CpCbJi2k/0zzECeboppRRp+Gg7nCrJnF0
dC6PogpfSBJD2lot916eBi0c6EnXW2hcMhJWwZEvTYYbJlKP5QQR/WHjdUB9C6im
du732SA/6v+oz4kas5JXV4FHGtizdohehe60No6hq5e31o+KW4Th1IlIMgpRyyn8
auDofPvsCeVDlVGr4ZEDv1HDYO5ueD4tHZ/QdGRQTooErldiY0Yx4rRLpDSZralD
JTP2xCr1et9cYaYi5xHGNdqXzNt/xSoGVBdifny9e8M6PQVZwVQwJxKQzrLnGL8X
FhDzNeFLbpRQJy6L8rZKBg+msv/L6cWV5Nm2szvjN+bLtYNn5xQy2r1a8pWD1DHU
n0TFZZRjZmh6Ow0JAIr4nuamKVEYr7AdL+b+QKigjBhyqdwUYey3eWHjtR+Jgb+9
gX616zxQfF9E81bD7L8BNMdUCSheCYVsgfJ9oUY1Qck1lUjcXGyZTZbZLOOJcUaa
7pijt/e4H/HWQCYcKX9W9N3PqbNycHQ/qnT3NRt8JBU=
`protect END_PROTECTED
