`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gZouRsFK/i10lkGjwft2PFl7rUGbfXIPuB+eV6cmCbEHxqi5C8u31eKAZMowX0e5
cDSlPsNE7yKL1Tc3+ddImv7mxY9Lsb5v50nDarN+gkYVPlSKmGVoZsEqr1OsOXih
fCHT0+2SVwr93FSMOMZXBvJghEi6MSzUHSFClQwSw4Weu/b30iywWcr26oeuLXY0
N8CQEGKr3nMLbHJnDM+Uace38fzMNVcEGaEfA8pMWPqY1CTNPe2V7VreB46JWk2t
J8W6e2mAlqBwYTHlOI/yr9/qiA/vbLgeCe/ZHFKrdNSKPAvOr/PGClKd7YPLJUZa
ZNruzjos/3Zo6BbVA/IczA==
`protect END_PROTECTED
