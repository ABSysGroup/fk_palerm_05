`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KRIH1e9j5YSrIHrgv3K40dbPTj9jxSZEWjPGg1xK252lVt1DyI8C7pM9W+WtiDHY
6L7L46q8wn2h71Z2wfhaiuXfh2BQE6rN2nZA2kI/ibm1L9gfuaQ4s1x/DPDwiOCs
xABGRV+kMmEZnmiEfpOVQVYEx7VOcdPTUdOpFm0pFMywUKBl4Ymf+mCeIUhrYIVI
W7mtPe9XkBx8SnAQ238ajnI4SDPmNubMWAr0DdNZAEsD8FTnPTOoT3XfwEH0K/f9
oQDrVfas+3nUtv6n0u8UrMPaJxprD+hhI+VuJ/lKJogCAHuq+3WLKIvcSL2iZx6t
73AxYZ3KbdMEs5uVX7xmwjvexaHaUCljiUEn0d19wQDtPAzPNwTc7U1C7NdRGtCP
5F3c/9akJhYHMANFOakSKsf7kjlO6UE8UpN47cwbTN6Zo/Ihf0qgutbuRWQM5FVd
J6euk6Xer/GY/2tH6tHN2PhtS9GxXjvSPp7ugXwa1weG3kKEp5DUwVBi6jBgZJHT
n/kcLgix6CblWG7OkRbBoWm2LGIMxr7vRTQ2IUA92525wB9iAhXtYJCURju1NKDc
f5g5o3wbvwDJfg0DvIpq7V+p89gqCHsK5Mvv5uEESSIp2qTIcoySsNxMI6TJrbcC
WPHEymYnzdogJ37lQXwzrPj4Vvqjen9omjQsPvWggCfHjerk+oao9EJZGc25ok8K
GJGO+jXNYjENLY9ICm64ft5ZiqTgMr+vS3CfDPBiARo09VsSRLvmAyMJ/6XmJ1nw
A+hGQHglGbt2N0IJbamuEELaArvJLeuBbGPfRU5F/3ZIb3iSHCkew5NO8jy7obuu
kRCS64eTDRtj9Y9R7++rHV5h82AePd1cyAHVatqnZ8MQVUOEJoIlp3rAce/n/qNl
EZyF6H87R6RlQqg5gsnFDRP0G76gqF0yQBvzpKyAObxV5AjPtQ7oCRxIEZiVJTWW
0MnL3YIG5ZdMdNKug2cRj+FNBhZETmKvC4ce9Hq01cfwrD/+C/ljiZEy5SHol7fd
K1F5yRV1QkADDOjk52AT12jWn7OJ+eR8QMq8NCKmDYdLS5h4vJ/LDrQwP0FYm+oM
sjCmqdmb9sKT2G8ja9ToHVO/wly+ylUDkAk4VcBH11nteir3kgmywAY2GqVWRIpT
vpFqxWYDKCweEHd2GohhNl39M0DPmIYtvHcI0mBijlcOuQW3wmjtyBL3kdrkncQo
uS0hoqIH4FlzbjzDllut+eefaGG8Cmuc7ZUXYcTB14Vd3xD0GlJo33JiYFtXgTwX
wAjqAg8QEuqEWMIwjczoJdzpDg4Oja0+aO97OrKFjHXKJVs/quFzbwkix0MjMiqr
1sXvEsNGUHHE0lQUOQZNBaCf7nGkHzzFjkBDjTHUsyHKrfZ8uB9xC7vtPiemeE5X
BrDYSkoNbawSBRNmugrfXr56xm3O+XCUnFWxuHdyjT10UzMOKa2ve+ekBNbyUXed
y56M2ZAXJz9phXpsvBJa1u33uYzjV887yIm3APXWCuMwJBLQwuvkpElqR/4sEcjH
uvac9bDjPrJ6Ln3YziJZHyT4qRLqb/Ilz8NMnU/cMWdlub6jRB4HqzZBz/aY7BsD
YSy7T3i4pITDvReF43Li7CsVtJ8iDof5xt/yBYTeM157R2CPJUtuUIinhTCNeMLT
TAxvEo/evxe3/PH2HV5ljytOGQ0kAJabhXxw2aiNHRE/CqgSBfrZrOqZCErq+GmX
sMR212P6P/LzAYWvniu48PoQcXPlPRbUqtvDZVZSJ26EZ6FjIaeuJHOzmwFSRf4Y
+WGplRjiCOlWDtJAhtaoYH3AON/1le7yGvRW8/FR9yDN9uAhdKWzyuPjPJkl9h+g
Cv964C9w16jCti1NpYvISSY8BubCzIV2TEA/AOorQO1byaus286BAEFnuNvx4vzd
kr3WoDicpH7eOBTtN/LJuNr0SctY5aiBT3fdz7NKPJFk2J3hipcMcbSp8pe2RcNj
8fqEYuJjgNj3nDi/fdqj7Fz9fbK6wZP/FxW5a1sV6tH9Go4FKWkyLRpM+MpJjJtm
zmJlz6v30SdCZzlQ+/R/zYV3t69YvsmvH5mNABRIeHtpw9RO/MbvGR6JzJq+obvx
oOO+Zt7XF1DXIe3ohDKY+M7SuOikXCN55bkqsohLTXG3HtadiL60jMOPSvUbt0s6
QUq8QKFgK2sH6r+tt0+6maRt2+3n60aFkhICCQg2D8nfq8qI/fRms7YZ/5tLfNie
KjG0sjVAgfBylir29lTRO5Dw3VnezfvMePyITj1WTRcOuQA54Dg1K+Y67fOLDgiM
zQ7nmC6w2q4upBcqUptFAFeBKlk3YbJISgMlwZw9UMCT7rkyMfuYB5aGRkw3xqpG
CULQ7P1WCwtidGXFq4c7LTMZb7pODqKnWHYRwhoKmOmymyy9T8nr+VeFVqm6PZXq
N+1HosAc68EExntiIsH9KKNo6ByqC2bRPAtOhSHEWuPVGsInZH4VV8gWzo2/2Jaw
oxx3WaSYOA/Remgs4M8KMg1N5K0IRyOeAI0znPbQsff2zHR31vUpE8wgFLiXgyO0
s5BWZqRMKiA31Uk9nBw9V55VjzOEllsqV3Dg3HHCfvhVE3JkW/zsu7IS/WvEpD99
7TsaKgSzPmZbviqxjDh09Yjv0QEudNcAgbg/auSuCniz5SsmsN9iQ7Cwie0fGn4D
kF1RObmajb0/gvj7sbGXBm65RKL4GgV5+mwJO7ITjBNZU/RWedAyH3Z8bUvnnsuJ
iUPHVOtp9VAS7bynJkUPOyXnL/yomdhODxemz7cVcn+pWT1+5mXuY5MO9GvGdSaZ
spAMZrBdIM6msTUb64uyWQWa93CeZXL5Gmbj4LHrgibokdS1uwsJiCu64yA7hOsQ
HAycI3dEAyCGehhzsycSXGAxdJB4koni40h6NQ4cfYAhLNBro8OXtZEIqfyeqEsA
wRDZnFlCU58al22TGcE2qJjV7B3yJtXX+Acrg3ih82+QVH3g2yONdvtAXwUzwgjZ
9WHzIra13t1aORQqSYCjRxhd5JYxp58CNvAqz0NEtAG+UnwDlpmgfSPWylCdVb4P
4DDzKbXwrFHkorXi5bDOjtNrdUd2VK6s1jbw6eP7n2Jli0zyu5JwqEMU+sIvY9wZ
Bj06tkRQnKBCORrS7nABpE17UKvCFYe8DHShqBJklCWYVzWuvUKzkDX0CXrXwMaY
kJHUOMFddJKYZFN607Fgjs+0Qr+/w7TK+pD+yNjSSLaMlbs6eBZlIIB3NfrQ1RNV
1Sj1yfD59fp91yIgO74+Yu3K/iQuEw91T10PZA3Ei+CsImgbH2AIR4bGUHM3SEkY
2F3ZpnsKebWK3sxS65O7e5gGdLoDxwfymZGG4VNCHtcyBsi84wOb79Z9bFsBWu15
21ztTqKz0yibhRGKOebG7yWkdhTELRa8HFOAMkQL8F5l3YyYDz1JgXUxkXPPs4Vu
AIEIGV1rQ2aTmm6ILTPDO+0/oe1TA1VbNY5sgEbzkzDzg9fGIf1Ld+jW0BTMRGZZ
IvfG0CXOQL7BqXsdJRj4BCuBnaK+EtcwopDin0zSK8Bt6WuJ6bNfenjAZqshWUv/
jrZsvSc7wrY9t3YIZ8GqDPwYLG5S6I1fNJHT9qzqEwh+r2FAgRllqvfXdhePsSTq
e3qNHNPixXy4mmB8dzRovctIoeUlUii4jX90bX8CED4Qe2sINPaZGDFlBJaGz1cI
IqO0P23VCZyzOlGQcQmgnDFuDXozTBMOYj8C2+Rab5kpr6LUMXW0/Df3zEr1Chxa
rQIILXNIzlgvv0V1mea909gbxWDbxYmstZqYSC+0M8IpA5eVVFJocpsaadzNOsm2
XNsK6GVEtgRMRknzoAw7k8fCwpEk6fsxlOb6SpvjTyPMJHpMjWub8hyBhecu/d7e
tIBAaPwqx8uBI2xXY1SMRkgTAEUgkVXnKKDwrcVE96aL2AOpg19RysmbmscdjNGD
tSGXSFNBEx7+znjB1pzDHvgB8vt8K18WuVUv4FkgFygWd1ZPV2sBYKwe3gY8Or36
MeDm26GUlj0jEZBoq7ewIpky4mNAl+gumaniVTajkuAaP9dquu7NLqsizdqyyLvl
mTr0Mw5BsUfYajo6JtKrJhyhLRT02MJ8/JnYbN0PG9T0rSjfbrKG3NjFcuk6l+ZM
i65P9v3G0TEupgrBF12m/QGWB/aeJe8j4/MtUgJ1wmwInBCmbNMZQQPou00cJVpA
dj0WWRWMVDcrjdK87xPtpJEPABTEorPyZqb8cc2jIsCcO2w5I+oQkXxUzVwSca6G
lLn5h/yH3ledv3TqLMSTgF8DBDUANTeSiwoRhdZBhMUYp9JNISKcFLZmsWW+lT8x
Cv/fOZtKm3Cw5r4DAbdiGgodNHFQyN44zHvity75wh6edEWhZVj1wiuDhWnx1JMg
LY+eM888TnVDMNAA7DQ41pygqehk2pegFUIPtZlrQvrnJ0XNd+w46+n20Yr/9PwC
Rzhf3NzsypvFmq0YvjJBaSufjDGBj4uBCfvtZghcaKCvHf1LLjFFijs89ephr8Ky
Bh3IQk/feUNfsnPavlAR6H8rgndYZJvduOOgW8//NcNwFHT80rZVZEKsRb90F0oT
gRhmWGxcfe2LRvHw15tcoAL92rxinAma5cZ/E+mWQAYcD5O7n/Vlk9mj/cfIhw2u
eFyC5epNKkoToJPilyHy+klnmf8Vadf2++OHaoaV1qxRmxaDT67nDvdIYsOoaesC
Arvwp84hMVclPO0oMIO+eykZlyrpFRqHQ1wgrUdt3q3U0nCE74jyjs4tDy1DWb4A
ei28mISlaJaOlHtIbK4wAh1eAeQPUWVb0HTEfgrdZ4fpcYfgKQwZcyh28Qoc5lvM
1VTOjuUIKtkHXP048D6ccM2qcoheMFss9vw2Y9+D9c0udruZRXEhfuWEA/8H8AAa
1CAGiINWPNodk9nJDu1zqZ8h1Qpa7nAHBbsV7ZNyje4xdGPuqn8bZqSIJNcR7D16
BHm9x87C+QZ/DuvpeaVXFNbSgX7UpUPO7etGEBUyVp+T+uORCXMPpMusIGytsw1Z
tAE2PcghZTonR26xZ8RITHoiMygJrgxUQVFJeI5auJWg5NrkXYFSKzkHv8IYZ2XP
fHvEVhYzqemsANlI5n4bpnRIKa9zzGxg1UqC4AXvNydeh1mJbm7ZikXxCc/msEfu
eN2lYTpTI5/NZnI+zK9QFdaSIVTeJHi10057/x543aQzf1dJ3Me+oMEwZbV2YQZm
QjMOI63WPPReeX46F2sf06Vr7kzpPy/uH9wtYNrhqLqDR1fSTzEqcuU9TJIjAnhQ
pbLGo1lncDUh/meMMU0f0WCKgO7zBHUierHBmDwIVnPcErFqp+8qqpFNJpFNVjMC
+EccRBiutkz+JD3aNNSfVG1DGuqbiivkG7ZdJD8pWpRnBWF9XztJV3WpMbb7+8om
PyF7G0ktxi9MwY84Lf0oYy+McRKpzwRssTROSA8X09jNmkocA09KsnD3GdTBOni7
rW8k1hHC2HgYGKemn9Te9IUkU4iJ8yu/C0/GQrP1U0Kqwbb2oQwVGB/T8PbF9Y87
vBB4CiXaZJ3m3yz6c9BZ2/zmswYnZ6Pl4ruHZjl9oy783oj7nN8Y53t+fviqVDh1
/lI5feCc4SSzN+8r6Rve+umGpWhi7PDOUUH6HJhG3T+xHguu933qdoPU9o+jzvJ2
GuxkfQnwyLOZidqsWskJ+pnoAzbHImnTiCH3ANJY2l1crMKmg5JGcA4BiZK/4vv0
3AVvGBpEIJTxultZbCKWuKJ+ehX1vCAaRVdETBNWoTDeIXuD7e4bMD2YlY4mckuJ
FKUy/Txqa/zUYmbpzHmbUJOIfXANe0VsR2p8Zif5Nn0V4Wuv+cYXcvj3rx3cNTCL
mqNqYpmcBcKfJ2jCC5Z/5p3NluHKeroAkR1r1RCegtG1aTdSNCSusE4wk+Ht6n1z
IRATGQW0usEfJsPq7Q6MxqvHahmx7/p8N3vrwTHtoEuaIqUkgx+lRRq7HO4hPAEF
h+YAUwH6iWTzNtqal62cp+DlcIHgTuxbEOkYhKUzZJ76dSKU6Mrl/OMTrlbTcoZ1
PJFlghX6SFVNLAhzVpeQoC6/4r7Gx5Io8wFnt2hnPMDMH1F5IGzk+CTbd8Hp8ARO
2RXr0vW1QhuiTB7IgmGQrznBkLZ4YqzdulDSgskwCBfUjpqU5lUcv3F6ODfZe7Hh
C5LPeQ0Hgx6FkPSldyuns4gt2FTpGrmw4pDyL9EMu5zcPDa6f4TiiGa2ath+dAnI
QFm1lcJnmn6h7yGfPXzF/yRZPr2+4OKRKlnw7/knqYyXFhnikR743JL286y/Nqg6
oyD4oSYPxyMwxhgEP1nB07s5zJ75yVxA1mS28OYPLsmrYLthaGhTlUYe9u7t47NL
KyC7FkyHUTWOmoTTtFm9+0eMTl6KEyBPvVkWAQlT/EimQAwu9MOm0cMC/ka4r2T3
VJ6qPkbD/nNiWqvfQ4WJOwnB3SkV+O49eb1QgdXQld6SWai0otTVs9zO34f8cqf1
gi/KRY23LlMHvVcL8TCxfiZ9d/tQGqX7jiqTO+sSSxNHyPeiye+NjPZPuNGPVs3g
jXnvaEF9eKMFHgg3iT6yhnAo0XUb9/hyArbbDjXSArjV0GzELUl33WCn2SVZRrTX
tZbYFKhZEV1etmTakKMSPpcxzEZNv6qBt4/P8mqq+vxirx2ab8kAxOEbl6nIrs+b
c6LmQ4K/6wz7Xg5aroFRYLdeLEp94k9TvO7hh5NHv+d2hI/WxSywMDxzyzJ4NFWH
yF0EZoZScuEVc3/4pDO8aCYqed1WTmiCKrZsNZhw+IFdxvPaYEPVgAmCOm+EpSbk
INRtqhgrW2BfaDRa+UCmwM+awlvLNqFeg3871Dsm7IFlKxNmagRpXvSRGJ8YLDrJ
ZAp9ZgReROlfcnFZJyl7erFM21a91QmSp0O5gylG6tMcP734dzRj2jOVsVFWO6h+
saVim/5YIRmksnuDuw8O52JJPugSWNx8O2VK8g51/cjjI1zM+1M16J+8BTiHzHe4
jp69sFfNQwpLLwoN9YEl1YRhYauvmOz2yFu++wHAw+e/aVp19HqzByvKgE63OVQ2
8tbznwv4WCBQ2KsJpviSpgIYrHazp0IaOCfeRt3mDDSrLXXANy0fPQnqzCQBKfPv
x6PJ+wUTPyxBsL+A4mUXvfEfoJ0AiaTqwBZdm8RdF7gfY/DErM0GcWzFbmMG+hua
jVfPcL4oQ5ukJYD4jlg00Zep90xtl0ZqTWIaOJr5Qx4WPmh2ILlwKsfxAxU+E0gb
E5+sjH01Fp/jyinHH6J4e8yXFjVhJLAAlqeTLxBysuWEe0SxYazdIe+U96H9r7iB
h9BvoU/fKbrvkqLsxNxILFFFl7R8sjamo/iJQgIzJVXv7qrC3HB3UiVe+BMgsim7
+A4X6FKhba9juBNYMrfDnNAEEF5tF9Olj4YnDfBPGI+VP2HZX6e/riZ8ru3QXstY
ah68YHuqYFLjUZdJMgQCShDfcsQHPBnKAhnppsXXTk79vEYLHgZSEvL4/CP2GpDe
vZl1uM8BKg+jsEJPaeHZmf5Cayi3Q0qlrd7v3ksJV20tSH3oODf39HIrBe0lHCMR
72P+Vn9ngNFNHH/IJWIMs+zhJJ7vUc6u1BxKu58FyCxFGZt38kD5ZKtElg0fWNmN
qITdAKqHQdzwOpMtuRIqnRzZHWg3A0nlqmfSswQALze0NVCEfLt4WyIRL2LwRpZz
KoL5hQhUgYPE7mKgyhd1KVgO70ahOu6zyamKELfrXTjwtiIFpIC7wEPIdHYvbT/T
g2O1gL/4ScNIDejYtrHzpG11sAsIvXH4cIXG5OzRzVN9wxZ0PZCkcgHy8mlfWtpL
GcKbJ/yF+SHQ+m04DkDOSoGUA/ZooCTxC1INJlHtSReEWsLXmZ0t2yDDxpbbOO0W
C2kLbKShPdhHhfzTk1JgHiVAqbKrMpm/T5vGP3aoFt6kiWNmXIxWY2j24Zgs+ZF3
Pazcn/ZoRJeLlvni6fXmnIwnGSF+z5cbb6gXoXMNQdzJM+rtnRVzSrVsu5AK3F0Z
bndruO/Q7MBsBJln+wa+3bpBAhUNQV/oytrGhod7X04eFg/yM878Cyoru+HpRi2A
qS2yrm3JPuw/oN9C8f45y/Mz+hVrDOpYbNphmOV1k8olaX6vtZoCdDrC0SBKoz2Z
WmguJxz9Z0K7+Zfcv8cAzw7KtLDHyOPNuhixTB3+LTBLkcWhczyeJSUgA1uwWxue
bLbwlS572NGw2jnyKpNEFUJTx51l7nJlQSp9Wx8jgdN04j9jn+kimTc78lhUFBAD
kKu8SoS3ecjX6cX32yFBr4KRhMJhvyr5GOOsh0ia/thfibh3Z0JO0WMYby9Jg51T
kk8G1ykyr1EvATTyu0632kAJzW9UFiMuzubuergRclN0g82Si21HWoaN2wYXCCje
6bhdkiMIGQa8GTPHoHdQY4DZcCRwzRO3B1TsIoIziTk4LVtJtDjhIexkX1k0sIEb
mSS1ZqCWPSbOGQZQW3cM7u8TcLWmb9g61ff1rQ3ALjOdQTlunIE+i6RNqmH+Xspc
mplT9YBP7ctAvqwLL0iCQnd8tKq2JC+RjdTumBkzw0es69rWBjbYzDGzQe6s4P9o
GK14GIgzT5eUZuOTHZFRxp3BJVQvbwL38mCmN11ziW4GiRR+p/aSmJ8DhK1uhNwR
GTzk6+0OjP3JQpTWiN26FnvjMjIIDvUaAk+Xz+kkEbD6livE11eTZ970kOrgGis7
gi+lhUcIryVvVrAgnH4ugTlK9ThDe4A6hjg0rP7zAWKxhMxc00/5l+zfHao3WtbO
kivmFirHGzQ2QFVYrSd0euY2N5ifVD+fMMfK61KibM+rw9yXRBQJpGY6QlaCx9LA
WDgGvhgFYjNaAX87ZZmQjpdJmr4yWeBqJx59fe69NXXF4wx8GxKTW0rDZsdKvaW/
LV0R+36/bqTvjEmZUtD+HUibPvSGeKtQtaZLhn8y2ntXBe2LDmPXqFGVslMrN+KS
Gvr4tQxLEvCn7bmQFyN5xPN2LV9DQygrvsRPcmvYV3ZW7Rm0Ypqui1GrBrF4IKUS
d7FETuC2jF2vbJJm9Fnv3mtHxZZ10Lphgo8oacG8rJTtHnKWeVjrTppOvX0zGWrk
RzS0XDJPBRdujgKW1htBy53g4X1vIpZoTeHQLWAmMsyDGP5PdtXhzFnYOOvMU9Bq
VenxUeLQBYPVZAcq/feR+2A0/wWU3wekIEJNiEgMYJzzvCxhuytsEX6O2esgRdgj
y7meTyOZrDR6BhMJbMCh83/5YqyIWnQSmO7rayhLCVh5UdX5JacfY/ZxWdqC3L2U
KYXn4l+Pk8+HfuvUqSD7+RXO9Q9CnkFRbyuCHE9PnsufAwbOnPO/Yxtjjz6fJfyN
YyOA3X3NgDC74MQlcB+BTDrgoZFlH+N7LeqqYdcF6UgiFpTy8MaWjTF2xJNtvneR
yhPlht/DOwf7xwZiAj/mtN1eRgwc0AJmudAknFLAuv7wtSiAmMTBXDctofugDplA
XR13QSjPyp4DHifjqwO4P8Ea1VJDBqGJzzZ7G7nsAmjo5j01NlDe5p2mImGCkWGI
dhgBaH5hMAicny6oETo3RnUoTC8EcAk4iQtd3mk5URnlqoiCqPNBf1ZQ1cUuWANE
6EASIeQY6/jEEUSpXr5RyCtcVmiOJvOsjSbL3j6ujj29qjVibDJJD9LaurG84tKY
D5B778FM0raTTTDFSDkWCO1xC3uXTe9G9ejZaDhGmBJaWuT0tIap+lJiXFp0UDsU
6ImZL7dHZVgokXifLSZGGugkcEEBDxORQHxPqaSkJdS5mevpLbJ5FWNmFeUqBhgR
UIimKluy/rq5PyDzhc9tGOaf6kvL+LVs6E0h0xUcK5ULvpQ8eXbmwsB7yeN8tylb
MhaCfjUXZD0gnz7Thb33n2kSD0CA6k059Vvx2vOYI6JamnN0qTfDMonrBoZm+ENL
oGHpNDGuZ3thqRQT9lr3QJ4jUgK5nhZKC9Dz/D4JKXk0jmlafzI0lfL/JdtlcJl0
LEHGKpKQezGCOlMKbQ9WMGeYj+rDnM0QqcHyYd3TyYyapGkaLjZW6bAwxWtWt/3s
3Tj/xmyCj34fmWyPliWWX9q8LNFTd08vTWIWUCYraJGkUqkOBhwz7wuRkCe+KdfL
1ut0LnQVAgTTT2y2ZRmCNi5fiDzAuO2SXNib62gtkT1D7Xk7OcaIUhFRqQWBWTzt
B9NxoTL3gn1yVZoOWt1cVJMkIR70Hxb7Pd7TYbJY5mGD8b7mGtphywo/NKac7qEu
i/vTZvzs4mqbpas1gT8eb+ZrRoOBHqCEDOXl5phQylD0/uWpWFWNLfoXmlWM1L5F
nlKhBpLQBWA/5k09Bum9TySD03pXkbo+WrX9892C86+gtfSXA7JamD8Ji6JW0oFJ
pUZ0D36AbW7ErT2FXiZ5QToz+BZOyU9sA2wXtDEHNXBKcvE+eKmhYjipYgBlQW30
YCoaIAaR16MKIx4A1NIihSJw16dxog3VVkhNXqAEClzPC+zK4FiCuaTmne4lCkHF
CdTExAEMRlLAwgc5kIkTCupCO0OWocybWeytyY75EXwnv9lZ9ZTXwFN9EsM6YAKP
lHvfpS9BUKWT1WZGAA0xwsvOJHjhQ01W2DQGZ+o97wGUoKgrJ+FYFbML1FDBPmII
eUJJEfcXemioc+dI7bheW0RpyqwVUQ5MwStiyuUoYvZbVGZLvqBVXKVJFjT4Paf9
qvH2BZmkkCUwUaowUwiwZdI8BqvRK18vPa/sj6hggxegqe0kEfVAVMn6qlbhVuR6
qKVaHBvl3XvFnB+xgKphsmdB/lkyyQ1DdCBgssLrdM9L2VFn6HekX5Sw3tn00DOU
DTYhoFiSSUy2TjxnnYgMkBy6il1dLScsJXD8MWDjzXl35+OfIRspTGce/dgg8mIH
osqFYs1UD4yEWVH3LtDe/7M+zq5gsTLyPIjdRjKxlP8EkEmtBnzw305X7ji/lcqG
SWMAH4pA47UoH/DyayOYCyWeiDmChs/MbFAWiJIfeStXAQSAvXm6viMxJtZ33thZ
x2fVt8S7pZ4t0UYieFLIjQQzySq+SstlDXR4SjA8djKZX+O4IYmb+p0xc0Z3+wqv
dph3wgmPFUbr4/sUHwd9069XUpI3jVksthNXcTQwtYlbkduCP36qWNI+TiD6WoE/
AuI2l29aqcer0v5MM93oTjOOYCVpLD3X+HP9E3ghpZTFKqv+U0BPFGD9lMt9Nd99
wFit8JrkmuW/RZfZtWT6mt0D2iYbSRA+lZzrk4INSTOvvllkFDYqFdmLu+pVFb5F
Ys7DtaoIasbE1GzbWfL3kbq7hrjuAWF7wgePOnu0jLqXh+HqFIaQ3ShQwghKbBkM
HOUeKPuwLc+PDYCvzqbBrOYsbJZ5NXbeGHc4qdkSbK4g1JdtDpv+nj3kL/i082ls
tlhXzh2HKOFxoAea7gpXpoav+voZe/REGzh/odUktAvdHVNY7/TCO3VJV/TC6yws
9ZmnWYE8ySzrcMqh75LuyUj6Z/HLHq3UIIcDIwpGrnVzHFDyWCi2zmgHr5d7sTbz
ZkHmeZBWTxhj88Wo2HsyUbnt+d+IjaVeJ0gXaTBAam/9v09akEjx7+OBKGuwKPcM
e6KwWC3Rqg92kNifdY7E81jM0KJtInRhHDGYYPz8AHSbXNEx7WSQRvVbt9aljbKG
fEOy1vClrjCAHbiCcuee8Dbiey4LTksD2smYqzk7efKZ2OmDAYUQQDQXWygRgy5w
TywpZ4OFOi34zCXXGNtLaydZWvexs9Jdt8HkLYlUnU0x3dV57sT9kca103NSxuon
LVXRIfxGXNSRSumbGsxaJofVu3Uhmu8+LzEGhUlyd279PBBBvTg0E8cxBXP1dW7d
wAv4OX7CN5zTtFotCWSuFLU3MtRZpSmQAzYU7m4tlfkGTBcw9qFprDivaIGL1nvC
T8ghSQFzUD8Mb2/U4bn2vMMQxZXkoO5SIk9crLxzuNAC3uT66Xnf9QyZo5yRSwYX
+H35ZooR7aC7ipdqjl/S+AR5Uc02xVV4WTatsIeBjN+MVdyP8rXpJdRtkt9gOPLi
4KP++W3LW2WarVXTRt4PbMK/l8pwgOJ6BFK3cmIOm/9weSfwU1wC5kta5tdtuso2
z28V9x5pm/8q6PIyXtYFbvePOhjhWeW8V+Sai/gmUmeTIpCqr2j8uawz3wQZo+JT
C79puA1Ju0JxGwyfppNEPE9zZqWiy4eKpxRnfW+RZT+1MK5Cag8MQTcxR4ztmQic
oLeKzmwpUVy21y44f1+k8MA4tR/+YHO6gtlTeN3Y1jo3D9Phz1qxRKMW/ll5llnr
HcjimOOBT0IXsE5LYR9O21dOtoiBdR7asTQzy2GfJn5HN3YWrFU3wYuHUuIoG4vj
OKCBljU95oeG+Gv0E68lu6UPDK/SnVcdkbJuqi+2o3qYDSe0k1Nf7fmHjQ5NygBE
cEPsWi2pYOdXA5giQdFAmUeB1MCRasYUbOP+8aYEoGyHOa06mVxl+Y2ldRLQipwI
zbKuMOAxF8Czl61WP+qJO2TApIkkskpgxJSy07c0PVCLZjwHLUeKg5UKR47dJb8T
IWlvn4eU1jP7HJZjbHgWongXsYrTJsAwd14Eq7IthYJndHdskPOQ9kH1Bl+/5gWR
DCpqKXrr0Ez7r9xI4PcVIjs/Jxig3SndXQjcgHNvdAmxiohhMUVoXjdAtZqxJh4c
/o0ngp3cD3Dc8WRbKGmIq1pJ0awqkrdLwAzzlTzZWJ3ftwsXr8GokXO+TIFGwa/w
Awfy/On0577vT+ZhvTh5w0xK9401t2JxrspdSlQnIvuUs5x8DxzuA4K/RtWs5p6d
0fYkgATL9BkR7paSmdp9o0gLTOkPmAgS+Xr3+CZNFVQMF0dHHOMBGXdU4TKrKRzZ
6wxZttq8dNVFWq8EAlvwkdcrJBedb4t+MTuS+PwrgXvDUrW/kcZsV0NnVwlyuUHN
Gs82OlRMj06ZY7gvPl6hpqMWpti0RaFKv0ywVmLlWrSdQpkQFGUySfX8hYgJJoCQ
LrxqTJSJYrl4whbk9B1u8RLSBFnVxhpfvsAqrE4xA3nZ6phqvUhU76xiM/9jvb0V
eX06NCBvAajP7hwUnMkf2g6pxV/FkVRR8mxdpUKGhTOCJlEm/2AdYdLuTjuBY2N8
S7xWWrsL+pp1aBp7EkFDTDH1vGXhcDz3o42B77t4CxoSN+PQTzKralyrVK5dLfeF
NHehgxmzGttjFG9lNqqoskC+oxwcBWR20el1OOEr+BfOiDOIuN0CZPyhm/TmrqnE
xZxr482t30B1JIgiKlwX48ZL0S2qxiMbszK2n3b2dwvKq8t7EjXG3RtnwGms38hv
T9yaDpFkzLaeNeB2wK7qgm0Ujm3Bz0DFlVEjzNouF95f+RhtD0ftrcRV+/UnC+vh
0XqQUeL/cFV8+fcBhOCJut07zxvIHYz5AT4EYlaIJaB+6dxGB95hV87hMZzodMl8
h6XRGWJxK8/SSz4WohTh6ETufD1ckM/qsjAWabP+oDgDLceRVsnrYjbgOFbeBGyM
j/Z/taBzStPfLi2O3/7ayORl3xLtZnmYCwkfmdQMPvqnJPndyMOrr2F42U0qOGHZ
v3UWubG37s1mRXuSEnRWINZFbLgB+jotSJh+7T2SLzYGXmryqGsTxopfTE9+k2Am
IEOx8dce4bT2fGOck55LjATdYWADoVOdRIfFZHpHduTXNxxDK0l74qNZpcWFhqyp
8GqHkZzPKQtnxug2a2SVkIMSaEG5hLPPbfaXlULAIhqmG31ilG6CZlxy0oO5nnPK
Tt9B5Wh9Om6xTRVkFASIe33ZEgu6JgwLpH0IQfwZcxaeYql5HIasJoCYj1e9FXLI
SB5+ycnM0j/XmOK0DD9uuMw8zHMzzZroB1X2PNAuPnfRS4eV1bSFKuNzad0yII0E
bIGVj4ZoX63m0/fIRANgF6lnvrmFMcuxpUaB2S+6Zdi8kWaCJ9L6GrQDzjLoHNMY
u2hYifVDKI0vZuhSwLRzPNilgADjEpJCnGubTgh9iZh7OroYM0VgiJBFkkZPnU2B
LjQ6Vi7oLv5iW0GqJcH44tu7oiNzZ9wqYN4/p2dOCXU+20FSHhLPyhRZSupWndu6
cFZRk1D5rKaGtLpmViZ38X9vxLj1mcbekqtiDGnp1yeoBCTBtSu9upRF0/hMlIFC
0ibHqsx5zhESqbO4JKMtEKO4Nbp4ViC4kFYeY2JIslAOk4JN7jHr0CsGbRVzvA6D
23xaCDFt9K6ZHX4G2UuKV8mVYtpW5RSQqV3gjWR7A6Rt17d929tT9nRKCICJjccX
E28rUwRj0/ERC5DDcp0hPG7QfdkAFWbmu8rFds2MzTg83YSoZXKqM9Iun9vtInxG
mwU9qkIK4AhDwjoEkrVCeNY/oNXBncmz3v3Q/TWWNmXac05Wp9Z2rb378dNzH+Sn
XyMFkxUa4xA+zvRF+6sD7CZPgHwA9Aso95BHYjI53UeqsGAeaP5TjhoeFan8wJmj
VaE1kgJ6kkga7I1v6HJpSvlTDbBSbQFMawjr/JslJZOGQVNb+ml7svj8JBHHHtaV
KepNke8QXyuKGDiafL1nP590XmYMpFKtQhNWhOCooDCFeYvllAgxWZEE+GFQzxPV
DqjkknVd4fenZQwFnZjBdlr99FseNbFaZ8MmpABRKDbahSHI1TnFxSXYh4Y9vzie
uEpIxdnqkqaIsfXDAecUCM96ieDITGQ70149ZWAKHovikuiuHVjWsaLCg7G9dK68
BgS/3Uekz3hngSUEqfTZ2BXQlG4+6sSdG+2lZXiJSROvvLpzVHiYU2E+9ROiqwXw
QAmcr64n6McufR2weGfM1tkM2znpegpAVDqve267sblpv9YHPuhmVRfzbOVeTZyp
XzVeJdCxmZSZIjaoD9W8P1tlQHFpnnLqFQ1i06kuJ9arxjOObZe8wv9J5v7VCArh
FFol06w/TfrKaGwBC7CKdQuftZWpZTuTj1Lgdwmm81t0gZ1GhGORgPj3RIofMkG1
m36qOBwnAHKXmkfi2TsVTU+TKF3000hjsgSvrVGE6dy/1pHQuyEKBwYZj9b/ywIM
Jo3/9B/I6wieFlZ9rrN2+lgTlxXVILvFKj8tkS4lpAo0AeCDzv4m5mefRh61Hplv
5TQUBTDfcAJcoydU+RIUCrAavbvxUfgnewEXGBpyjJ/+TSOGj+29Ns/Dr8Bu6IZR
RC6zzc55TLOW5q7neoDOAz7cP/dJh1CkN996T8UJRoAHpESPyATPp2I3Bh42b12c
kKWLIscdxt2atTRr88Dypk4CU2vl65ypuDZhIKp5dRuvL8TzJ4841ztvIqibbkaa
+2FfiMOBhj+WWSVbGbZafPGb2Up1DPDsDW5+HkgcOi9uivwjAbwLH5uuG3Rwn4pU
5/0UunQTPhqG+qo3eTZfpt3OM6q7EP9kj83gGQafywyPjWiF3q3JfcPXeov07Q9d
fDfmj9gz6dmg1yLvqQrGLA8A7umEud9kngL4SBl46DC/qVtFiY4CfwTrB7/Mx6iE
vO+Yt1zsOOWuziiuy1Qf6wEd4ItAV4KQGui+X28UnpDXd5hAPQ2PIuZDXARENw4R
Zt1gzGHwJbaQaQnBQp4VmC7pyWt8sSGSXvNmypHuMMcyThy66AiQXfS1TDFFcsy0
uo2fhAnhl6qdSGcm0+e3Y8/oZVjLKFKh3arSWP1m5H9CTi8/ig7eKmoxid0nNMX3
yBJAupG0idrOCW0DR8AY7bnH9SZa5y25FomAhpUt5o58P1bCKSPgztHPFIxRf4hu
HORQC24Apl0Or2xayuZ/FEN11uClYAM02WTp+VEVc9KInccBNPIoxD14osiNQTxI
bdwFD+wgRf9U8YReWKHivCooTI0d6b+Bpm5dhvQlIPlVT8ZPQxh7Tbiu/9kFCxAk
R+ISsdHs6GWnOiI6wAKHHUo1UCASdOgCXBlQO3aacYase9yvsKhUCWYql8oZNayQ
euT7yS9jQfEnWXnV/hSd0HtQZMFRjMaOdZaYK0PiG/4Sg6Q7eFgaU0nE7vxLrqcb
rYfs0YnUEzNkFR2gdwPsYzRge8KjbM5nggkXOvOREr7EtCGMVIFZfY+mxWodgEwL
jc84Sxgg7z9n/RsTw43gYyni2RVJjR+7GQH/AUZkFFJRdsURG1YYQRGrvwkFzqQF
u2z227YrAJiIOQqJnhUB6QbtYzdwuExTt877c080M49X4tioCNd1vybAIk48mcts
H5usxEiAQO32MtHq5fEKfvSQcuIwyqB+bAA3IOpDhoIDhdCrWiWIBAmzuPE7yGFN
iAFGSy355Xuf8ACCZJn3U8VfVJhLNnLFXYWDv5YlhvlJfPStNfcTLGwCTfaCQlvj
LoqKPOt69FbveMkZTQkrdwFTtLKhtWAYVe7z2/EOTBnn3uro3TUku4iVDaAQ5Dtm
XvsXRm+NxvWDC3WviPB1hDhRHYN/bqA/RGNQ+KeU0XsNMfYr9ZxXTRv64f4eh+N4
2xp6MDdmnPxvil9OAvM5XbpNUF+auEVb9FmHcgoLS7n2fcl1OHHlX3N8h1ha+rnP
rj2GHZK+eF2drvQidQIYrQrPw9Mt1mezD6lRwAy66wBtkIHh6iTaAun4D9KsHQHT
hOFi0czyeBZmsRfH17ib7eetYKIBGAmZ1aQyizuqAKZqXBkyfQHNawbj9OM2Irp3
9Fy9JtO0wC/Yd3BZ90FsLnnw9mz8gvfaUHvVt9CskSHMmGwVbM7OWgegrQMEsg79
3HoKL6Lv5ruhcUqPIXBc3LMjmcghxjPsmsB0HmtzUpBoqLUAFUwGtAwrYFbicWR+
pj9FO1BmQOwNN6OBnDzMDpRzJIlMr8xUD+OzjHJl7rgqvTtIdc0bcIsL5xhZM124
9ojbwApXnrYOQLlld09bJGTFaU9PkIy0/6in62hHqbylWwvSefalm1Lqf+roMn5o
3HZLgf4cTz8FkQgLc4mRrW099YXL3njAW6xAW7FAisZetb6EkWZY8sTbOl8ZgLR4
klu1+n/fvWhf39WqZIo/hSJNf0w+p4gBjD+DbQXegWgqkGsyn8xsrA+5PNeALssj
rFJZ1D5hr0PODf3NIwUYO+g/qETj40FYIUYiiWVle0PPyU6lHi4myJYVGu/49M+H
6OQ1lhU/KTcux0iTyrsRAeunVZmrqEhsXMCsLt8vhu+4TYTZ5E23Vpi5yB7Rn9/z
G2LJiz63iFD741NGo+atqPUG95GeHUTqaNhnVuP8idF+Dl17yhGPm/peG9iOqles
NwefwshcAf8pL65LAlg3xzdEBbTZ6cQNnbiumIh94Ba+xnWVaioN6xVlX32SzqnW
SeCtnCx/0Co4cag3N0ephnqpCWp7fxN9/tIijGpCaW26zyXkXSjEeBd7WyCPsnjZ
9dkNdtSShEdYodwqlIA9KhSH8/jAAYraqHOcXE27e+AHAzFZz9zfI0lpihUG0hjL
W5H/Up0mDX7Ge5lpnuhRMK49T1tNFlYPxbNslB3DLur3qzJcInG9NSGSIKpAUJ8Y
sdOJfYHGLK1AMpZjzsmOh9JbncvH4v9NFVVtvsVXd8Nz3aiSQe/DS4+CL7X9c3pg
UcgSSA6U9cOPXlmL/WBxuinRtitnFhVtUCLuwNDTDbVHxZ2OTEtTyYlU2fxdWSIb
fRCOnGGOm7RiJWm0nc68MSTIJbG8DnSprdPqaKXc9isbQpGiKo9V21NUlhUaeuXO
eqgLfg0rphwfanf8GnIx1LVoRnOUCfaK2f7J8nBdbF/jZ51lO1BhJIfspgQmkz1p
0g9f2bOFUBw2oPHSTERcyMUk7IXK1ZAoZi1oOmJD9w7Yw1yb27H/fSfzkmaFZWMl
zE2Muwr71Gn78lqzlwOeNUJ/oQWVcHM+5ioWau0WLARmBTu1j/sWvpNvfOJeX6BM
CkFYSFnUf8BFRa5wSjq1+tjH9Pa+PNq81UGMm4C3Wb59nN6Ykz+GhrVBvS/whrag
hfYEt8QklpqQnc1AeUswk2a5xa2NjM7jVOdNiA3AZthRzkaWEuh/Sgw/TTaV0Idl
5Yzyz+dfExv31jLN4IVs0QNMIOQBu8EzUvlFHoFN+rw2isNuekPWod27MkQiMTyk
Q/ya1dEyg/xyBLeNo2A+47DO8cTeUKmd2mzI8VtGCLI/nV8te72ExB5Cafy/cAJz
Ly4JPrHW4mWKnlyHRezlrUUJMMkMZP23+MDshO2qCnLdSHu/5ZmbjpAwULQVZN4x
XBSJQkNck40y1QszEpeO+HIofACohQCWzaNrjUs658OtJFtYIkwLDOa1YRtyhJ5r
pXnOl25BApdExgeNz5RdhpsE0coewR38hr7j2DmRzBwyuBErNzWnAO70rJe1y61b
TwFv6IvZjdBrbOy31oI3jsfeI/AS97QR+bUbU05x4+wBS8xrs1FH5CWNo1rEdyD6
FY1IlLjDufOPUMInC9vjEj2gpPrhE2Byfueq+XDdYUzixoCCo0N6/or/ZbxL7u0S
HnrvGj/dZFdSnV+nmHaq7zTiJszrlocIWfca9jP10RAOMjB2wNKsYGbg8ZVoAPor
cn6n+J1PHGYwYG8aVDxXXxjW7mOUFYf1uyxtu6zynTO5G5m5pmx4wMTVSWA/+49S
w2MvQqrIz0HQFOYdvLsVl6FbseL60L/oi/R0IDdQsMa1MNKtyauHtv9ZY/8s3++H
odoKT5o+3teRwsKoqNMTPlx/RjcHMV9DHPr37/M60TqSacT/5/ycCPbHS+3bt9Eh
xdPMZUQdd+4Lscy84IwTfxizXJ7a/ZehLksuzy4PC0iwxLD6lzXPm4nDUDNJvn/5
n+Y47IefQ7auP5ut1Q/xXs9ZICzqCG8V/Dt9VXAcixH0knYV3MpTqdeZ1g51eJ0w
xwTWGsOaiITWZV2GE1+Y1+rnVZnT2JhLy7Gx1tojfz6yxXwKmMzzVPJx9vQBlVVZ
RBAkV7Hs1aa4K49Wi4NkJ3wwwmPB58zvNFdAspGJgBzPRSKqFjEEdiMTvzB7HZQd
MiId9xXqdHBJWufqXCdxDqVaHgnlNni04UeGEerlOQ7mULcfObcKxk+LS1XqWOP1
ypQI7q41XyiN0wgQLhjakrN0uU/+tqNXU+vwzgfd/thCtawKwt6t0XIQ3FLmIhAk
dCI1vo7zMAeZqAA1l2jdAXm8VSlFgAwSK7A8aOy3Dpk+LkHNyHqQYngLO7Z3hQ8c
dZRsXQsTndJWEdzYVedkCgE8qy2HNvkit997dTk1cwuNKZNNKPRiLE7DqRcdffaI
U/P35FiNT8yDCCL/MbxWTt/RRBVu/IYoaaGQWVagUQAlCDYMjmBeA8TcdxJ/QuVU
KQL7/e3QuthN1g7JwEVKJ3yALnwuc1k7McGFNy548Y8jeEjrOzUw4yraY1rNTdus
9DrhdY1GyR6V+N/wyprHXKFZ7n4NoJvyic1pA01CONKQN3cz2d/gxSLxWvs0gux4
uHP6o7OBeSlaMUJGxq/q6nf5Cv9aUJr1It/cCPJmEiOUvSi6vLGItuygAT7X70Lm
GYJh6PprtJA9sQBtilgQG4phlU/eb/1HmvdBMFmgSC9c+tmtSx922KtvBiewZ5nH
XYPhXyIZn+oHQrWo+0Sr8MfANkZ727InM/Gxrfdcp4YwBugS7PolY4oXqAifSNqj
5HKJax5dbTDg/wVyCK/eLyGFOKGXB16g4WnmSmO5h78L9Fmap+3qCQcvA677Ngvj
iELnTkw//BVfONCgz60WubUf7ZpRZOJARBZ1N81LwPO4tW8ZQDxP51ZOlxeTZPQT
9r9zItptSGjttB0ZysuD3XP53nQEVUBOp7oHKGEH/W/sTc2jOSZS376z/WCyFMch
ZoD9nJnMjtKGn3zG1QfFFjnhpfjS3ifaTN6yeVG8HPjo0fUNcZE0PT4PkmCG5OUy
4ttAYrbBDrr33hGIOnfpgyiOgXsW9V1xKlWtHnzsp47laHFSsaczqH9VSniz+Rcq
9vEKSkrgt/AU4p1y22mU6k5UV6yL4Zo53KKiVKgkpTd82R/SR1bp1zb/nD/25/jA
E/CwsEKcuZ8o16+4/7nlHYMVQw/KhWrnpb5UgQUpuiDjI1w8FIM4QTxrUEa0Ut9S
LiKjOLU2N2Lyxgn2EDrbPyILLMEngZZ4PIzfSv76IMl5ndVEIp+6LqTmPJUqu6Nv
lUdA6un7wJT78Va85twsxBT7oTwqlL90JvRqFht3W2oLNl2oLwdC+nqPVL/PPRr4
6RNHtrseE99iqkIq5Lu3rGg3ROF7XQSnufT/fRABzYsaqExiXMjapwb4A7ch708G
D/3rCpLmUx8BtCeRcU7nUkvYqvklZuc6/IK5Dcf0aMoL1lmwaSYDzuUhrQdTcZ4n
Ri+GhSv7M6r/zbUohCRzJDxesBHyTFhksMaoP2+x7bqpqJpUUKPEdQ92U3LsoJSJ
aqmHYEqs/J6D4z69nbvgHaCNk/nFKP63Lo46+GEvMB8yxMpIYINTQqQyFLaJju7J
opzCBFXBFb4POtTgRe2z2OujLpjR/kuKclThO+kBpyK7PoIqLITHnVv6nS5qAStf
Ku/IizjxGZi73YhbDlHRl8DpnAbymk0UWY7wKvwuC3hzYnnqfjcZk6GqcGTdTvSr
PeSi/jedI+a5JHJ4jw0gCkhW08zWgb6pXKbK2xbbiSMsb1OHN7llqNtbHTLgn2pE
tVdihPJp6BKgaj5Y8rxhIqsDGml+usKgXSYXa/GyuFsVPiesOA0PNReDSV+CEK8D
EfixcH6JDH0MSKZkCqHmQfCoc86YWEBAMLyEooy6IKqTn4r94ODyZOfY4xbBfvVo
zcYH+ypFfDtpTWey4QieUieZXrvIaWaL5cL02vcZT0tsUpvtIa7ZQVznYUMZ+kme
qtCv7tIPdXLkDM2xgWIuFIZEJwrJ1NnwlshvqOjfIRoBWTyitxP3A5YrjkM8D8u5
BlqVvjY7v1/CE+KLcGdw6iZN+L6wkXQfuk+p82cvVqdFVHOZFiV2cOXMtbwXXf5z
pui0zDc1qPVOwS1TxU87A6Va2K76WnYT06kAONjSXlEaxvF1zhjYsOB4d3TlTKUW
lJ7X81kUucIbHlUQwKlkb5TQdFjXi4f79bXYUF3QDmQAmIaO7wvOY/6G/eiSrM5v
5j440hOIsYlYIQ9Nkev5AW5taQQfv3hHzk41lcFU/CbZt0cLve7YosR5LE73hU8K
OEUJKFUCwQkaEg5Wh79qVyxKCG5hfsVEO6QGkloUTpRKDveUp909dORcxVWN3I/W
hz20C1QYTGzCVZXWc/Aqwptf8z3M2TrN5Y9z7IdFBs2AjIAI9rlMRF9JcxR3mfK3
7yd4Y90Rt4Rirq6Vv0W0z4jLG93Jxa+tm2+ReGipVFjkDpUYCYzjH95FcJVjK+/j
3zkvgEYqKHVNIDz4KZF2tREkgydYWsKrjJWQ381fekMj1FAcVKGG1yGmQyXsA9KD
PauV7Pr+hgOCj+n2Gldri/bpjKT0aDlyUFfOTYPlwEf8dbJeD974sqrFRvlZIQMx
04rFiRIJSoDRfS/sycATdD2Sux3KJ8q1tnuDXaLc9lMLCyYCRTx99hFNzY1AhLi5
IQzX1V4MItz5wMwgaayJAdvPdpFfXkjqld+nnMYu6FAGxglAGCyXzuTY7xC3ET+i
rcFy2xQ17HCIIDy1dd39z4EMezqC5DvKK9PAjgXNwYX3IxV9IXXDreaUrVaOg9Gf
Lx55gRa+RFdIApF2JYpwKFq2+0NZYLSPL+JRefO3LYoMw902qjQcf5D/KxgwOGIp
IZz+j/hzCDEICHebmSU2q1E46/qjXB1NuvGtl0NjW5vUNuXWGPgRYgVbzJIiuvT7
O6bU2el71cyBb7W4FTwrrBQke4hM2egbZSNwkJ9L9YyrfpWFde39b9ScoX0D/61w
6yM5zvuQNFH+4zVOeRZMdpEy0pQiKYXqT+2anVzBhrTl6wbhB04TeSM98enKV6Md
MI08xDfuySt9raochI4g7YPTtXuLip2QIEbMXHpjOJGJftSZnSdvdm79a5yy5dZQ
wOdWmoBlsdVBixqZ0Sd0z4qdQsSC8IqpzUArfPgGhEqeHuXY+3FBaBxSTCwihq76
sBsVuyA2dc0sByx6EFyUT5k78OIbMoORC228aBSSeCYesjxhTaAMADXYws7gpbfR
GX/LN2w+MDkROV56omwhwGoxUVVba1G72Vd+LFBZXjmvBco/+R2narHjqg4818qR
sLMi8IjcLeVw4nXE/yrc842wTluC29rzRf39C9YWMkfopm1VXMNld7klA+LceQQz
Lq50Ut0xdYBlLiEHpMZ+gozPDoWnsBvZSLNP8pMp/x46ipEGyhFhHHdByOK4TVVe
1hK3f1e6k/OYuioy214Azlc73S651Lic1P0HDxi0ck68Zt3Kou4ONcr7c8wMIaMP
ggMUzsSDHiV3s+x9ICTP0bMoFgDxS9c2j+S7jl1Lb76wmhwA/an+HURIRDCGtmi0
uaHhgIXUICnTfJFqXMmPzGtte+7DU8O4hF0/Xk9kWOm737twyGNjFl+u39BbcXvZ
ohz4wFtCacIlesAefNZXbkS1PpyEBXUQ2jzBIWAMtk9wTCoY820ihzl/KOdNiQWS
Eq8pclMt/B1ntrKJ5b8DB6CVyazSmuTK4Moc47XGYMxFrgcSRXYx54LIWqI1wreR
23p2OkZ9sexEQRQWZrB2epRVeyY01d5aUKvXWKkAd2OZVVj7qYmjbfi85w4u/v6Q
Qro1ES7csYYyEu3l+9kmm2+ZMCXGjJzxtfble7Hnh/bkadm99LtTH1iTCoJrHanC
ervqE0JwGD4srWex//fLwjx7dvpI4k6gZovEjIPu7RlB9ZZx5+skYkqtnEMphI9E
8NIljSZMJmRXWrv1/YuKFZhvXDr56KTdGK94QXCaMWOp7JNp43hH8OZ1ZZUB56BE
vTXUTN/g8sF4nyTbkRnmadF2svqyohsfVS5G8Z3Ivd6qF93XHgb9LhAaylsAqaCd
K9Fb/dH7mxlHhl3Ytrh+gEnJCcFQxmizEZrSnNUytcMitb74144BjIiRVqVLbPnZ
osMKfy9p6DjoC5KQX6ENbIOjtcgQoKd5mZHTZtECU0LXj2Qf13jguIKO1Wp6L7q5
tsF9o22bxVaUZ0Kk5SvBZs9XDuIsPgB02U2FRmG5cWMrexztRaAxZlkM6mP1V+Ay
rZ7+4/nrtF00rpm/W4R3AC1Xb32SkpNGGxWhKemn5inXc2xMJb0Z5IAknIr5pzon
b9U0Vnnf5lXcrQdV92LtCoGD0QiDfS2IKls6bcNViWF21tvhJdc9G/GCD1kQJQfh
lMK8Uof3qAQtqvt7+xDynrJl2hkizh5GqIT/8dA7/74C+543QArTyqsCWKL7sHWV
06MbhhRtR3O81pRHrOQrrQ7mUa6QlOueeWIyKZ3TcwZjT5rSyyT5V8SwNzxuvoO4
SEeAss1TzIAoc+Na2tYVTQO7DevxdmzkxnqvUJ7Gn0hHsg2l7Q9cxie2NCgAKYis
Otk7fGrJokdcVKs/2iRe934P86ciJpxfR2B4gCqUTZzAwSz/WrA/QYgAbPhCdoXN
S+trB23RU5zRbiXeLG1Rnq3/QRNghsSbh2ny9PQTW1sRlZT8nU2LXwkj4Wvbfj44
KsglX3eZDbSmbYDmUxldS/EuTesFgrX4YRHCJ6jqIWxsOu+Gwkm91MZJhg9Tleu9
24ndTOOKW/g+NFQ64OMNfzKqxxI68GYvR3S41xktc0aj2x7oPD73qAG7hXqXnV/Y
VcSoldUK+79XkdCZi4Fr15uhVJwNJolSni+gb9MKKXOaSA6VLMCXrHArBlwZVGJD
TLOv3jMFCrixxB8gsA5dBrYUq2q3wBEkJBiSCIGvwvyhjzuSs+7fGnI8/nJQ5f02
j9f/8CgWJuACDcXjpgM2GqxOLve1isLovAQnnlrbko5/ZeUOFE2F8qGhn6r++d0F
ZPdFaDoDJwNGFa74MGDt4dPMEZAoWcBT9rD4wkU2mVEpQHmJSO0FcbeVcSz0J18Z
8sYSr1pclGcetJ4rtu5+AG9X2qXZN8Eu9FKgnqGcUBhfe9PZi1ztH/ruh+tNclbc
ryTiMginWmZsIqjXHQbugEtT3uA1NckCZ2Txjn9SzCtMBHYep2lt0fggUCVYBLMX
7IaKPTW3osBrmc3/lAeuxSMOT6i9gloK8K9wBv4SYnIZd0y/bpHM3XRb7CLCeqHM
o7zPx/Uj+1ErgPrFH1N+p4oL6u1yvQwkV0zJqEUY58LceOgWQ7IdjKdzpRyoXIuL
kZM/mwxTp2TyNOqxRG0yzFRYN1RTsnyx/EdAhNN504X3VGfX6IgyFSJJohZKekjP
EjoXprJdxJ39UG02+DKfjje/SdFwTYQ//auS4Fw20SumNouSoT10xm75PeNho6FR
3/9Fao6GAvPkqdxxoq3UCt9Z8GCD1cd6OhXeZZfxpbNYDNFxY5VBuQLSo3VvDned
P5g0pE26jUhDY5F9ELgcgBXiIpBDxzLNYBF/CFiycnW6InRtoOCTfK4PUUR9q1Zr
wx+HKk4YvsdUkyoOavyf2BDnOsggmwpjPVOVn21RZworBsysSE0kkxFjFsgujGGf
+vapMqxp4vMJ8pwH+RmgjTvJJtAYKEkT5VyIlN41cCpbbT5wR4uLRL3q3snzQ88h
xfryk9KZE2wZwaHaK2tOC+/0E7mV7m72Gx7C0hNjUz/3oy7jcWcZWwGR/uYW0ik3
EFLFwi6Ngh26nSnZ86hENYxO7FJnhUHZ+fykOenmCxujJh8gMOHj5o5jzq14A9lt
i3xkbNPM1ayuqe5npf/Iejy8YaVRHPs7DCjiDZU4rSM2FNNl7izVzB1np+n+hCwg
TgjUjp28w4I7CpZ26iUog9rOEu0rhvMTuLIMr6V6O0EZbOMC8QRl1M3hQcUjU7Ve
QYeJylOoMBeaoE2fcnFYco9oY/v5rUnSdCTfbCvlw1aGdOyPaWXbKmSQ17IXIaU0
JEIyvppY6UIDRPKB2UUctdxu5+9QChQbj7xhIV2ncsQZWluBTa2gKUbHRyHhzG5c
9a31fTNz4Cg0lDL7wZfpY2TJpmuRrjexUHDwDYCU4VvR2bZSfOkgmH3mvkfTKmJc
vSDvbBAll388dNrnDj2LMfwCfUH1fRtwJfwJqtl2h1HWf8hT/N2hEsjpUbo1Ov+e
ywOn4HNQJRb7mweYPftj6qcDYHUNeFHiQI03WkfVcVuCMphP5aYjEo/u2wE+vbmD
gkilYTan/pEkBtjGFIbRKcFbUe3RA0VJwxT6c+kIyWUR0ElN/7pArXbEtI461Sk7
odvIR9PcGM6FOA3n9X9fnbKKn/Xh/juGJNcZ5YwAKmfeXN9Qe0hEAG9Aq3EgQKq9
jlFMJ8r+uEzDx/qldun/xVIRUKM/HyHGbdTNkLDEfubCA7r25nnpgkj+lpsCv81s
cXDkD9dtDJ8WoRCzjrGUEdbCG66hdnvH9bc7FYHdUpV3mA4mM8CqtJ9J5ShsE7zj
v55s4OnA2OGJpirHbzT3hVY7DpzXEBNt9ZWIT3DMA4ZvGoF3x+ObCugtPmpIzAEj
t2kdZWyluq72ESYBhh//eIBQ3VU+odHbjvWoKnvwsI8VpqiX5GSGc8TvifmHE2lo
m4UhuCaV8lqhOE5ltHo/InvI94BFfLT7uuRu2kZmk8Knh/sOZFNd4LtEnw4C22YW
P0MQh8faXcux5Me3GDn3p6SdCQZq1d7MVN+CORBavSf5N0yWJYmYXC+ciydPD8/L
ZceIuE/42vHsS+QGqDsGOrNF3EYnBdwWgfqGST+McCqT1sGBG0FUsIJYc6XtndNH
ykGe2hCRvUFhsOabRac5Jw6/J3DDj9NfWxCozBpi+iiY77OhZ1kGUsEE5YWaPpSm
kTEvnNqG5KjV9AZZR39kQZJWs+KfqgN6ZeY3hyoarEF7saWfB2rJoRDSZH1MHsC8
rrYDy/sJhAHFy4vvjR4uP6Ly1x21Rh2IUJ7pIBSvwA7+gl6R36j7ND1f8GpfC8Z8
M/Tp84na09Y5NbWNfYKzmjTNB/lXq9x7SSfeMaipxeXO2ZJIGFbyU/R57ilPOlH4
LqUGTvmiT6ttlt1bBLshT2Vl/M3YCZApjZMxpWL+WYJLWTczFdd7oZtsfH9yGjPh
AWCshUbwARjXqAtaAkeO8Sc+dZTKMGweKFewHwxSA2jHzoJnRazcPRdAULWlYDEN
SjiaON0NOVY12gJxz8wbcDSf8QJEuJvsZ75gmltpLez4ke1dGp6KzfllKq4CmF/P
qEwFunFAnq98CQ20i8CM4gsXc9YpgL7ZCLg3OAthA6RlOZIybqv4nF4FVshFnUpj
pjBra5tqOii759EC+1nJB+ArFnXCZTgLKNzpOwPE1jDVMoXoNAy4Y9nctAq4VkIV
3yXNMJLkGdlejbsRDfPp1LwtBT9gUuCIo9VP4MhiSBIrPCuw4z+JJZZhPqDTqX3i
3gZ0Du6zYkRGQkWy5P5+eIKtxyXl6sSNKmMZ164/bKpJomMbNsGqpsg7oTVD4kfX
CQXBgcat3tPYpQhVCPN/Vi9RbE95pHJTlr5KgL2bUOD7dzKRBlasZBjq5ICrkycR
+onh8vuymwWVBzJOsCYk+NptqDaz3vL48OdtPxb5Yl+LHIdarf9oWrdmTVnugxRI
9j8xHKwzSHJ94ana9afVrhHr0LBIdnrEpkcGw1dw/8XNxmMydNHLu0ZT9zosovz0
ayLjBEc4qf4PUXUcfaKsizBX4qN7qNbU2jLqQoo0Y1Ye41fQX5p8QAL1tQOSJZYN
OkOO/zhlOeYelRcRj/VVg7nQnFUXzHIJnK7GPMPLlf6GHsvBZc4kc76JrM+Ey4nw
ejgZpa32Vd7yAsNPSpU/QXSs8UOYA/uNbpLvYnRaX0+uxD0x6Ifhs8meiuje20y4
ocR9kJPLsjYv/2I0sBRxGOa6VydOsS4opF4r4g058PS387b0fgo0yv0nYwYYK5yc
Q80dobeCPZ7AnuGxxkGLkqixEJrOren3of+qQ4gN1GAG86wo834H0ntpWs9FxazN
FlC1B38v9qXRUrukoUosH9Uhx+v7lPyJ+U7fBTwrcgZzMWtAsA3cEtbNK5KX6hab
EX2rGRLmrGcsumRXdmq/c89IYWSGHOKeZU/fM7H6/QGodslzQPGcIYtgaoPzsChz
gL6raVrHces3LKs2VhxwWFRomTlA8FZFFLAFIRu6Jz0ogFEV76qgJW9JtJOhCAIe
zrNtisAfYBiBqQc58rW8vf8H7NwRUbdx9rIThJGgBxL7lquvi/rrd3vGl9ff0xCE
mmGgX+8HX9Fe1MZWY0QwuY4tnWwmcEM/li/wNi7NqlaNkBoeug4b7xgAwPJKivbs
BAdBNWo0nJhe1hhTdq3jjd6KJAFRUoocYS0kBNbeOSZgthM/8Zo8hXSrnxrfBCYm
v9Ablneh6WvNoy1Ux8/kUMcn9dG3yWmsDjVwnhJWPX/SSwtGZzpYtTmWDfljAxno
vgsBfD2j5tfzrPlHzwTdBlOKW4vCWKf9TKAnAi/trHsXRkJ55+8vjV0j6JkCo6HP
rdiMZcmSLtK10u9UemCBgmlTkJERcLOIUWFT3XMiyfB+V02wqYUkYZvnnaQHuj2/
YI8SwjMYacGj2MUQOjUj0PDSCE+zA3ReWc1wSdT9u06b2mBaTDbi6jJg/CmaYst1
O/J5PA/b1J43twjDu4tVae17MJRR9m8FsAzwtb426azMx2Z+0rsK3kmck20XHGXf
8aaoD18dotmZq8kuhU++Z/MK2/npLCKBQ1lPqFYSU1IPXQbNFux4wxLZf07f2nzJ
LOfAhCNimx1A7tZYqz0rSEiia/0euGRNH3BPtNq9ssyR/WjWj63Yfiz+U/omVZoh
wTqNBQZn1C+B56eb7qk65YzzyKxrRFIiIVEY5hup2lPw1nT1g7bp/9JLkiV8pcG0
Sub965JC44fsJzfFaH5lPSYuhap1QFZ29G61YfshxViEcPRh12snx81nffDJLUS6
0cPX8F9zzrf+kjeNbVcu3HQNfXq3bGdbfx+AazFRGlLqlsaqGmLMS1yjyiEohA4j
QQ6rDah6bWM8ybRTHCyYn5he7biDIPCabKoIXccRnyJAXjJai88UMGDMFtpzbmdA
AjyjNBZU7s+cCDJFj3s3VCet3H2xam1ZosXokQOXwYqE1RhKQlxG+NJANbFOjodB
hRKAVxJSvwz3sZrGas87s4is4+ljXizrTRu4QmiUqqq3hd9KYhP2C+kpW07ycRtt
zz/robcTj9sq02ZrQkaAPwoq82bGsYPkjXWFqhBDj3W+V4iQ0QfVAEkF5IImJzNt
hhqGBg3sW7ysS10SBzrFMJTGejhgd8DOwD1OKtGX0I9pfizqK91rw/KjT/gW3cdc
ssdkvjvyUOs+3cYNRqPw+YfNxoWG7qywxVXL22s+OZSQNak27B3CSY1C8SJrNvsm
hfMj4VuDlWllCyEOAe6xlfTxMxWkS8d0m8MDhtr5R9RbpWKGC7jIbPl+XmlEo87t
c2qbnbROORiLNggrY2yK131AjrI5zFDwxaK5H/qaLGp4IxnvLWHhTo1kesNna0yR
IQTZ+e0/kCrGMyxNpHBFWu2cRo51m9B7du5ifUxELlWTa2ZWQEjWRIKbyjYiZJR2
X0O8a0cnJbJG7mLglngdwzdXQDC45n8wPzX6qqxHW/W5gUxdyQ5KWAVTyJn8i8R2
BX9suhs3fBoT3UYjmwoMWd98jXMROVF8MPdesO9O8Ol/5ZmwAbIGR+t7Vb8Lp757
bkd1XJEUduWqxUm0s0Iavs4tHUllOQpDI6DSspZnW8vMUaJ9n6nEjPQ+Ef9Rs5Be
zr1TcC9ZtOa/0q5CmGHaulzqshAC+X8hUzy1iD+vL8rPatuY19Zzz1PrAShQ7qMV
A3oZYRAUCRKkLNJujMlVSmuHpXS0bI5sM0qO+z51mKo3QSAlUDNxTt0lNF4hwPJq
affNKBAJ5Wtu/NnNficeZwW500LTZpNT8pDFwbL3dVml0HHsf8AYkAwI4YRasGgp
I9CO3SpeHnmZdUTxMUpLG7dXHacC4AQjHka8EUuSJbXzdYBGAugmOSGewIkMnUNN
V7o0gF0K6a6+mRfb3D9c/NG+4nQMF12FtQq3PzMM112ROOo64+MZQL6ZyBwZazgr
wturM5Aod69UPIohUSkluqFWYO7DRWlS/7SEpmjkUi+xhDLkptW/BRG5doLsyXS+
cW18FiedN35Rd1nyXB3ywyAQpkcPxj4JaiAWwg5dq8sT7JmrytVldxThMp/mFPfc
by044JzqB8sVXDi8x5R9nxM2k64WqxtgHvMWM4lbTALfT6IU8mb5d5BokXn6sc3A
N6irFk8KMK/D4MG5aDNo/eUivkYFHOxX3pmBtJifw8uHXfnRDDm67OBpmnZXS8iU
1JOA5BAOt0iDmHxAMUiM9k5ewRfOYg4isiaesnazbQ3mny3zE2t0vPGvnGkIPc2X
B/rtVWYZMfH04K88RKI3uge80954YlqYLvWgZyTpeToy0L5szXNUtFjZQkAAqcVg
hVziX9QPchuZ5CDTjEw04gLDY6Rk7KvaidGS76ZY0B4cYFNoeTQCQ57VVZVQ7sKZ
B5cLeKoRATP34o7j9A0qevqfK7Ntd6R2cgIZfuehjqUS+xzmOwZr6qIVCwrFpTfw
wtJG8DJvjrundF5eac6p5fOBWYtTmUafAkLEz4hHwwvxdP6jBq6FDUaQXmcJPnPY
wH3+0OiHKIRBCU2OI+GrUs32jcMXc1oFbC8D+soR3bKLnW40fACaOa2vN0jKHl5t
nEwu2y+ZbGQ1zob8aiEJQuefHsLQsKhHM1HGYeVzapIAFbp0+pIS5GUQcsG9eHSM
MZNvbD7cFkAH1PTPgFhtxFze5f7qK2n7J/n5y8aIq+4x+QrsAuiT2OZ775o1Vsku
X7a9TV/Px7V/Ku2Ho30OvkswzjrazFJ+Ii8qTOWgVQH/MHNo5FLr+yQMddFss/OI
bZ48UWu/gTKM13U3iDlTn4gY58C/izCzIfKxJGErWh70g1lcL+y2deXaxpI9st7M
lqxtnxJP01u1GR/IoaQagoZlbbTPm8HpahXnJnG4gEO+3zh5xNnZGg3fw+knNweb
2uzHeNHnu94WLoXZAHSNMD4sUD5TfDkcuPvTYpFmGmuPMJqFQ1q3yBLdwI3QX+zd
2t2YBPV3Ow/7WgjVA584X+laBOiIIB2pAljA1Moeot0BkUiTxLiGbaAj4Wey+aMh
jsevH3eQQ+8TKDRqEVg47iexiELNKJ3cDWygDW2CcEMKi/fY/g53FkbWxou0zjsj
gD/AOMXUFCKWI8BmO/F5/+12+6VJn68GoTYzF6A1tF3DQUQuXbWF83zhF+2tIV8h
LsLIpL8RuCWdApweOpUmsWVGlw99ZSk7SVVAT8J1wHyA1utzG0RCCUE99dfz0OeT
fmbZ5tI7bGW6+xMTamrwz7HiAnHk5fxtb+Zle4kGxDc/4NSlXfWb7CZr05YinMZ8
N8eOkAK7Mj+OeJ75Z7y+Ay6NCvhicsryUsgynHnFOJJPSL3rQeYQh28UeYbo96dU
R28d4DiCwG0pSGKxaaD8NGoqUI7FzpQG+rciMV/A3C3+hWxtHEuM1Jbi3zgaMVJi
R1i/VPTd/iLMd3QW/pbBZvmyzGuPi66qDSorsjgTR1aes7LQNU0ZWgHeFtwwB5HV
n7va8TVf95iWGeu3Jn4U5vHKNMMivwk3Wn2ROnSUl0AFeP9vsjLpD5Q//W0CAuiv
uRapUDsRZzkQHaHb94TIw2BVVyCoaYp0jdKxVs5HEwCKmtDRnF6f7ViVTdJ0TuuT
i4PpPEDhluMDJ5klRJqxzGBjHnrEpCK7HgGaDlaAy14a6dE+s9ahdpxijy9FLKVS
Y/Nh78sxTeJ2sOYYp3l6zFrR4MDn+QTn8TWm7r/v2s0aDQFbstzXGHJstmSUrsdw
PeRxY7gACzcC59xBvJJsiXzHZhvfqiHhsystoIb3qBVE/0yhdem809Q0bnZk1qIV
RzDIgd4hMqgbIdfB+nHCzi2V4I5+Jf7SjrAQnSW+PFQ26xwWtRCh/LpT1iLpsI4B
3bxemqUHN8mAevqv4VfbC2PX0z+VQaZgNVyqrbvSYQM70CsYE3g6VedR6v7REMND
MQmgP0uM9rfA3PTNxhOFzQ7mrsXuPK0dHZb9Fgl1M4f4XBW3VLpseq9Hc8ah1ufW
VyLDsBPF4maRRITqJI55FpNQ5Gkfa4t1+aQQb+kvA8jqZu8lFpPI9YA+zEjU0nR6
Q3+KIzy44F6XmmIxmNFvgxSfq5REpZUALJEc8nsReDIsKM2yLht1IIQGG/u2KHtM
1YYwAsMpEqJob0L3YR2dVKe18dK3j4YIoTom6iAevMOfGQevMfi7Iv0+RlRjAw7Y
MzRaz7XQVeIluS+xNuogg+oX0bcZEa91ibV34tMlt2Dp8pr/bqMSeTKifeioCd0X
dM28p8KdNEakG3mQCS0YGsuLQU1PBWYp701K1K3Ssf62/hkhP8tCJZFqrylZnDAC
EFYOj5/Rv8KwsZpfj+WL0pmqeNpKebdfgdjLsnvYZkqpZOUdUAPJP2rBxh28X+xs
PTNgOkYYVGDGVwbIdTZquT0R+xvWSgK5uMGBByehwbLfqQ+Y/HkIr38HZiozcstd
DENd8eMIjpSv1OkrnLGfr75YdD28y9nNI51nbwovn1lStCkOmt1uUdTeV3FSAJOt
huEhKsgu/2qAdCnXtIB96E2OR4i8xmaRYAKM1wiuFw1Ri4IAkSn70mqyUjBQuUCg
JhNArTV35A+oWQhSI8nC+ri99sVgFiYwXTDyF1jXmivF3DvQNt/9stGmB6Vn/hH+
SxSjcJO0XCAIYxNlFWRvSEvbV/8U9NOcqE//7BfE5r5BSjbeSsAMjTWrMNAcwIQ3
FLTJUTQcKXv2LyI/4VFl2nxkB/XwEkaktEM+X1vQ2Ys1RpdZEBfYXNhcTPL9doSa
btSzvAQhoybWUSCePES9wvRQSxYuaVf4+2dffa2Tl5FM4io6l+MJ7Zy1JUSi5TPw
yWYWfrD9OkqfTCLSWrD4Ra9AQAZTc+HAgBplOnWbGjF3Q/O9qDboaO+0PsnkMpvv
y2YpAPo0dDhdFAyeLrMtVAIjjWCIaiVkGD4QlM3cLNwhS7fbLvCFmIV0lig6abw3
Hakk88DUvGIEYveaxvAohztcaL72atanYA3nhcmsH3ZnNctY1I6RciLH5oxzRFQK
nBQbHFn9Y/c0BWB1ZUPhJnDxp6FM3NrTDmH687MTB2M/r6axSM3mtk6jhBDyS7KO
JlcgnZYXpW0jV4W+iJaZ0kmvgzFRH+onH7OhTrt/JqmY+zFcHb2lMCnVc6VI4Xau
CLAGvQqRIdoyxwamX++PZaH3SNAXPJhrFw9ZMmNF3ZguenkpraJsGR3B+8kMh2rd
TB2EaFYj9IYNwiBp8bKjct+f2k7rZDp3z34C8diIbgJeix3nQAlN+BMUT3O6zNik
Ptmxw3MKLNAwXgsoAFcPrzxjsHGh9dnkuKbduclwDLqHwWYtPIbPHvnIXKHcbcSS
ESxkrsWC8ecb9Y1iX8uLKW7lYWkuwZ/lMInymiJk95MM11GOfufhbnJnKZL49r2O
Et4f8Uy/vEjXKOrlH8B3uWwj0SZwMd5glY4N0d+z3p2CvTex+lqs1KAfgAKUYdvx
C1neF4bN3LOdEgWQOOSELPYSrhAr+pXpZimCtehVRqmZO3qFHYSIE+2129lJhXqM
VY2cZ2ZcqesowCuFrrh57LnJw8MeZBX6RZUzpvrLgsqZ+C3TsAbzvHlRpC8wCRu0
PM+zZM89qMOd5TqoR165lOXYYDMAE4H0qnRv4CgQvNq5yWr9DH4D+oUHtLa38cz1
nsnjDtzQBmqY260CYZXVNfWkdKgv/DpCM+ibj69kOdk22G6IOwttl7VywNEJj3TX
N0is/g9a15gTCN02LkcycaIKjsMV3dVfGVqAkbvXIXTCUGkyTSVSasVClTvIfgza
KzmtMG8iL7cVkCV4MpYzyLWdmd1HvPBeV2Xi9n3ag9OKDbp7uoIbVy2jP6T09Jpf
sG5/IQlSOgclPcV5q6yuJgGTMDa7hMWXlT9VD4B8Nr8sd85EeuV9Ixy/ag3En+8b
lfcxb/JKm5fro6dOqyAbHC0HLlxqmP+Gq05zFq9w30D2XJ0RmfHcfSf2Gli+qtrP
9CfCU7sJC5Y9NNeHJ8K43MfQ3dX8MtwU6Zj+xZ5GS54tcdQ8GBKtkjt0QJtiWjMd
rHBjRJffTEDq2g7wLF7Ogf+GWglFtJOdYl4evjs97+XmBNVBegDox0Kv/uxJa58K
/MSiuqZz1e0qbONQLx0Z71N9c3E715gde4eEtSPmqd3SLwesZHnZdK7BD6krmkUc
Fwuc+/dREYBa94VqDsm40b0VfkoSAUCHGJT1qwHNn/YmQJGy6Qn1/XV5PDiAXVz8
oZNcB/ZtlyaT/3AvntbBDc8EyAZmF0R9rwpyNgZmCu6QxwFYEdydDW78mFUVZPoT
xBxyBtBg5AScQaF6YMYGy0YKaaxX8gVqR6ramNs+bUzy1vcHBanYe2L2ZUUiKA31
wl9VFrsXTHjtyeWEhdzPXSAl8Ujrhe2nQFqFohBWtJxJzDZKsLMBEB+tZua6YrsG
lo0Fv9GAZTrKN13a1tEcaH/5QS5VaHVixpcxCl1OtBz4ZZfPoGnBGTY5Ewp6nSI+
uNtQqg7GTbDdK6lDPB2h445fvs3ME4yugMnuWwZA+qOr/dpRtKeexf6sHYOmnj4N
2uS56RsBTZnTvBjRLvCRecQ15AWU8wngYLiLcB+MZe43aXDsIdXkABVRdbudqiga
q6egHJ2YAua9SJCEKSdoA9aNQ9wq4c3PYvGS/XmfavzHm8BX2rcrOALCs/Aa5z/f
P4vL/EU6Z6UF0h1aj86r6TVQCnAsTx4SP1x1b9XNc/yZw/Jpfyx8W3A2x3M/cqtr
t5Nd3/cmJbQ+kd22rG3PEAuOuO1P7+HH4SezaqjalRynQVdQp9wGiRhEgJEDhrgA
NIzWFvjlBo/GOKczmaqW6DHREYWK5F/fNzQ5JZDjV4nVUV0K8yCk+6nhcbaEhUAz
y1EV8r3xnTU/DgnJXhsgEM61DYEw1j7umoBo9GqhgY22zAuriAfBkvb70LtekIbf
h0b4ISeFtfH9alOkHtGn/wmaa2WTPvIdEMf4zROnMcQtXHn0B/jSH6IUW+UyRV6Y
dvbW+6wJRgAsDkyEXhlKfdOUi7M4rlQnlc20fYQWXHxv+lOP+zNEi6tCIoEtjoRL
VFqfR7hQGuQJgQKSwf716TGvlj1AHHeBY0bh0CCn6KESFTeDE7d3dIL7BfzlvCPc
jQzg6IEMqwNe6i8aHklkdU2yx+Cue4TpjzYS33hxSVQrt5qEgqN7tVKd6EPcoyin
PiM922fOBgrF6PdPWNXMWVAV7umBvAQstgBHfXnAGkwZA6MODigO0YTbQxQyo1Ne
AsHrqel+XBdzQnAM8c6/lWXsMNF/qFAJ35xjzUipTor3PqCr8e0F5B1UH+HGYpn3
gmREO3BsyIy4fJ6aU9kmkpe1mYn4NfzxTVhBl3E+ynVjuVCTmVXN2H9t2dPj73en
6cAphU31ZM19pzAZrggq9Ymb1TusNvCRD1FXPHeIWQOoMWcUiCJH1HIRfz71W4wn
UihnOIQ/FLsvKOkuhqUJx7YH0Hj+6D/0T4uuaauuVyYisBpm3E2tT6u1kqwJuYsx
x7/DlbTbo4s1rkeJ+hfzqAU2JmEgPhbuAF1KQOOtnxMaoAdiMN5jH5mQu265U4Od
7K+Alj8ejkkrlb+nGubWcCM4S34EHMO84PrYooKDpkRoNiBkrDkB4yPUTwJpo8AP
+ysAHBXP7PDgaGspiojNjI38qjLhwBG5mBdva5YFlM9APgZh74nwC3oBnWx0QOcb
OsuypybjC+5P/WA7+J9MnKlH/luUaBagj29unfuJeDNRSnydQYVi2y8OOCsCN6qA
5dVdQGDHdJ0HdeU0+1Y5ukDLB2r3H0UaGv1pk+4GNGjfjWjxtOjnJ0F8b22FC5Bb
myLKONwzwa/OI+O5jHEJkZcX5mMfcgzIe7aSnWfPLueXTDenU5auEeN2/pXeJJyg
0L5ObeQk66erhXWVF0zxUR+l6lJ+FEHT9gU2Jkj5E0wfB9txkzUOPcXLWAQ9mY9T
wLpDl/Ikr0olCANZmbr0f0EHXo/Zx6KpLKAV+XUngyKWydTAOms7KZGQqROlhuQY
kYZ/2m4I6gYXEtDeg8+Rno2hgJdV8Gvpdy2oeKrWzvaYYOTsIaPj4fupMnq93KR1
/NTzp09qh9ldn9C6yHr9M3Gr3DbLBWT9pT7pbHIOWg/+NSz5e4S8nGhSZ0N8jYfz
kCpCQFEFYpsAawpMT+52y/zdLVTcKv0odWeSsU8iquoFlL4arY/TP6OjtBne3nFF
TiWSqEeOKxvT4BMHizNMnulXLfBNB6fcdVp2BjEXTSpZFdPAvTAHg4x3/Yi68VsA
C9lNev8jNsnfQSkGa299l8RTd3O6ry/pP0WxB4xWqI4UyOh1AZDumBCxXkkwDDHw
H0nUCcLwdggZkH1rzByAwTtEebHUz9bwJgtfSi92kSzjEXmGWxmwcejwd2Q6BTyF
swwrmwATApMJ0kS0JhHiWK5wn5BsuTKzJMNhmFwvs1GVHW6ukIuwk/MfvLyROR1i
VtURBoMRfE28zrg3xw+aNiRvqCWGSmmvCEuF8pBH2/ah1xDpCM401KPulXSXZn4d
rNX8J8BHC4C68SbzC7bKGfQI/f53OuYsBEDjDxKNBmuY8CeDglxd9jS3Yk9SdSMw
D0V3D3cqBPieNAFE7cMdePGvB+AeDaV/sCTbs2In1vvBR2fhxkUE8tLf+QbCTvPQ
JeFTJSVZEjXGE3UvbJCIxu1FHVKKCojAJNC0whAmXPSMaAxw+a1O1U9huOnq5WbG
917aMYEOtTdfcs0OoLsVw8y3GjYeYRIzz94pb5fnCuTKtxvYJ8Q/mvIQEsi+3/yR
8NkxWEyvBkInhdK6CJlRt+80u7LZHQ3aRmxWK8qpCbaPENYexPXLKzX4FZNHBlK2
68kPGzV0sVUKKvd8oiqyAVhcjqsQB6QM3XP0JioSF+Y6HsZaKz27+/FYM6k+09CE
u//j43e2CqnxJDY6bJAPz8vsaZ/G6rwttlNVSZKL2HlOkai6YU+7ab5pMyrdjSJi
677L+rNXtV/K4ibHisN4MehCf+F6kuVh0ytuRxbqgYq82ofQyedIqLWzbDsJ+3HI
Rk+KW78kBsX5cKg9qiRtoNFOMc7toSKUDGgnDWSa9sbqgFCk27Bwcd8EVsDnEjlZ
1BYhcHp2xfToWIjuMa6d9LYB8obGmYfqanhj+ATFQhjkgFIxPP39ZkOd8f9si65Y
FzqaUe97O2VOx39Wl0g1BSIA1CQNwcIoKiq0138591bqd2BsDsU5c9TBfQY8QdpZ
BTq+ufakHcjMI9PBTMtySd7Na1MPVuWWP/kPW5JvaX553JF+8p9sJssVnGZWrfr0
kSK8nqCPgycEGLsAMA1EnnOg28dsCPx/X+uN2fV+h5RLdHLG7w7fNbwK01y0h8Ni
hVKrw7UVjiSesKNBQvgELIvo/2Uy/C9FYDRR7/tOEmRJ1I5zjAfTJPeUKyPBI7tw
pw7vvXnn+TVd8X+QRVtqoQtDnjxJQAJsoLK7gWzrfTKTUD3u7mbQUrIHIp/NDHBr
7cRWw8AOOWh3xGifK/qkXXhzu9tzXnr0Y0+2YNlxAN9/wjoSbw6J5mnklkcOtLRv
yQIkztA2pIFidm1aNDtKZYMbpCHTDKOoOQlgkUpX/ssxmVI51rTrJYaiDWyt8v61
ONwzEs5luWFjaryXdVBT7QgTPHZO++CuC/kI8XUDGpD77lPCxmLlM7g98df08jV1
ot+HtN6f/89wMK06W6wW4/fUikL7cXzsxtlhxswyCewSJY1ZV0IJeyTN9onudnO5
soLeTv23mpje9GlpOgCeXCrjqvPK++OHWrEclygWlTdkMysJ92amYGj1kfXjzH3z
CwdH/3qfLf4VvutDT9f4Su5vQhOgN/WjXifnmjh7zo9xJC9uUAUX/0W0AAs8OdMV
cNAAmrxAdTcycW7bmMJ0yGpN5Huw86LIXhQf4v8cAq1XdkTYaLd83CaiPxnRBV0Y
aCcx/fweKJMeCIM5oqnNF8vCjA/AwaQ0eIbqUhdakcWxxGVG8H2u3eyVtKBFAECV
OVf/rgGSuD5A9LgILFGfAG7kGZCoMWJVa5e2Sp8iqH/P05jRlbhPk9ucD53eXl/5
tvFssi1TTZYzP3eeOWnwKm50vaakNJaxhwkfO5EqWRTXQr2IEolmxUEiVaEBKlxb
tZE3A12vFToEyJaB82DpQfaLqnwBukAXzp0Vpw5jCgH8/hlPTaB5/kW5JzeKF/iB
GREdV4wrd4iFJI43GSDY+Dgbkq++QrQNqFW046FVks+fyn2Xzepiqe3O6GsNjyLt
Fv0hb4tUvIE7ljLvfkMntvozkrQmp8N9WyJmjpx+kA0D3vtS4iy4qKHP74Z7PIXP
qXefccNug6939KhtJ6eKGcqHITsEViGncBktzywIPdk9Gpi75iIRUi1gmih9avFD
/p6NdZFBvH2OLbCzN6/1981qPnAbTCZJXNj/DrduC58p/f86YnvelUOehD3ItjEV
MrB0by5YFqvOFdctSCDCKIsjLdvsEZ3m3vOi5ZuRApPbS4MurtSlot8tGg6D4qH7
g/4bpwbEWAWgCMCAp56u6wbrLBFm/ztUZHfy1gdp3cl3goGUSIbAYCwgILtqrDgm
znvAEqKhCc5cMcdyKutQM9reG8YyRTmJd69W+/SGRuwFUWocO9vqfsmbPryyPxa1
1t/aB73ehoj2q01KMSnAyd+gf9pCX7mPacqGyPtSBPgW8jtXclbOXnFSrKA/LMBI
6OTrh0bR0OYWJsjo9xJ+g0wEsQEZ9TFaAdA0AgwEyYV5Ecbx4LLd6a/Bmgltb5Lj
8YcDzfAZSR6jr5ZzHqEoDJoW2Sav8EhgA8bXXO3Se1mhGAEfpxKVjKJ1fHLL4C0q
RixZFLWptq7U/6stbIqR34w1DpSGQHjqUB/EYO7G8h5KQEs3v6huZWSOeSHTjEmB
xmS9rS5vVGPee2hDK3l2tpMMJNadYIZOhugp7MYmmZgNkhU0wjA0AAi4eGIZ/cfD
R5tgH/nGxX6iIFlrCg0wjH6EzG/pk22ZtzpxK1CfrWAYbWS1z5DGqZUo0OrSz10C
I5wADCsNfJtdODIHL1T4XeNNtSheR9kwRAyFgFPSbq+wJ5YlmOpAWBhydfLJ+OnD
NZlj8Ca4vIDMSgvLY+Nx9Un75Y46IS6b8ktR6RSESoUJ0TjICKQ46H4yzM+z5Wuw
Qc7S9gdDOoATbIhNgaCCXvCij3KnAYHjSNmu8ln2FyHIfwXW3gAf6vtA+8PceD9W
Big1NSLVOjQ7e9KTJEGH8fC7diUWqsc2yWBoi1n9tJeWappUqOeBOFODlD0e+H3w
Il32bvXNBljpk6yBcDPPl9lYe7FeWHqSNHxxvFD+a2XwDNApo01XdajKLW0+47Qh
6uqaP6HscExyjGVubWgd3Z8VTlA3CGK4AyXaHhLRfbuc9mXP5BVft13SOz6CiRl/
ak6zHG4M4GIQW6gwuucyKwXcnRsmbpKHx0bevIXgbAEfQOPTfEPlZGSyIya2eaw/
nlSBQkGMzJFFYg8q7mWVplbPgrz+vR/qnZNgGsEOMCnAeib5SonNdrb8AgFRS8Tc
W0O15tVbQbMCTq9XYGdl1Zz2HzanItBQ5KSIiMYpB/pVMBodE+444nPxx24rl/RS
tEcO/411vq10ZxyrAu4X5vT8jj5BGbhgve8+ENVosqfs0c/4intiDr2DiRjhrIvk
VGvhPKDUr6o8ZttFBfSoCdcp77R/gu6pYDP1j+fmdoZn4aLDkF18J21P/kr7TdCg
xU+z7uxEGn8opKnIs56Y/IEqMcCU3a0lwh7PtBQrrhdfGUNjHcnWVa5Pqzgevl7D
fpm/hVtkP5fRFU9ROWorSZrgiInnCQNxKxBxpTrWXJY7IuEOP5OFslOoCgQV2ZFL
JHIXs0RLp8zGmlPNuxL2/RkGKCQBjvkDGNkzcc32yJLxgB1t5mZBinq9wznc74DR
6QX8HjKcm5ebbPU7So6dhjKSScpGbgzSic0uROhW7HPyZgXuxXMuEUS6EUbC4wCS
oJxAVDpIDgFvQNzfMcBpT26BTaNPOkm+5o6zq6XeWZRDcHesznOKqEZQ01XBTO04
xM+zMXu+KDCXKgVQ5ojwo9I1S8DeK+kdvoneeihyL3vnwI7B/Nf8JwaNUOdrr5nq
XC+kMms12+rnfxdAH9b4OO8sTwCfqb6n2/6EbdSECyN7epqWbVvxSoUEO2kqRvu2
ltt9Gv3lHzcCsUHOY10S2uQYtq4wXoY8b/YUkt+SrBC8egqKfsT9TgXxLEXscd/j
eB48U5TcLnP9ZaKqsOJNuYWEfRjYj0WE6/zwCIOLUZDfF6NEMjVLxmdr3lpIdrjI
zhskoz1cc0nNyemkm7hkstdfOF3kyQP2Dy82HNwLNcqyyOEAxMen94KBbl22xTUY
ZnYfp3H/hQ/HyHPkkekfqR8lodwVEnOApUZD6uqyIzhwGDPVtvzmr3I9fBdDokCb
DeXjf7IrTRUTngmTHyavYh59wGnLRSSzb643MbbvGPuJc8MSKANJypaKwMujAqWk
S/v7bM0tOnVJ+xJyDTPe2D8TRyNVUCmYLKUQVKd+C1m7umFZVIKU7cWuOiXBn8Hh
pP3CuBcoAwVmEUk5uNVhjU9DtyMlQgkMrIsxW8dRG/UVpB3ZXHAYzgGZwxRPYLRT
bTRSzfEaPZS030yGqFU1bygy/YDQeyLiiGY15yKAOvFuYlega5wfh6TvcAc9RU/F
4+n5fx9slfjaon/J7R2fTICo88ApYHKf6eaHyOmDUaA20JSMjRSjPLkbbyWKxlSQ
V+EpsTw2yAhuoSO3LS4tgMRLdIFa8Vthx1MU0+KLqDndL7V9xxWRzGaQbruR+R+V
i8XgCv5Mj02shQTgQlkUvDgmx0+86COAPu7f5Xk7hJc1jGR0/2hwEXe4+GFSBU75
WGl9XzOHLeKesxABT3p6NeASpV9rxQ3A4VINce3PP5wBQI7yvX0wFUKBjh+Wqn8b
L+YtjOGlTIoQAPM0lmQsiirIe/ZGVgXhN7aY2F17Rmw8x5LtySogmgP4EhsVGBXJ
i9Aq8o01pfTBKpy8kuGs5KktnCxKlzfXVszdwELC0dG4B8EHcbjg/xXq+vlAcxoo
SbKuOY8Agy2LDxxS8uMjtwsRDHKG+/jpDd49yv+dJbcssRhjIq0h2BSqA/TvsP+I
ibxegRIe/GQ3+EtkMHL4Op+XvJKsbUGi6c3U5VZ/IGI5XFe2QkK42o6VOldWomwA
/lChyINkGMTCV4WzSYt8ZhbpdnKs5JWxNgCWCkdQXMJ33CBIdVbGPg/Ryz1GM9VO
mJDVHqJLSL5b3nSa3um424wp+/elGIygRJ2kmeNd025lkgiE2ClTVSaUa47fmtJq
SE1tADNgxRaG3vYNCE+XrbM4Ixfrgp9tkHqUd9FSxEwSt8G/BtqhssgWreAusVKj
X9dJyD7CD/RDBr8/jffOCmFd00x1sjNiPbpag4/YzhPQ1JOkbN9/yT15G9nT7Al0
cxjyqGKOOYEYWi3z6/aukAKJd0O4uE7zWJZMHWRKW8TlGiLxOAFcIGsUf1zGhb3m
lyINtyCdiLcmE78xAFwcYY2i4awwD70AhqMaKac/tqUK2nLsA5EOpARWQFnaXBvk
aleTo10s6FJO6tp7YPgnql9Uefs10SWUrkgBUqdagP2mHJms6Ur4CoubcWCwyJjJ
621bfQtL7dRRj7htlaySkcWcZVXzCXAos8QFoXyVFx6ItszX3iqIp+WR+6pL8hBQ
61uiLQz0maRmjP4JBveOw2DfklmshdysAKaB/KjSWvvtc+8fN4jyLT6b/aVb9tAy
06yKY3ZhowIXdOLlijjeq6dujiR49A/YMeTxLYUWI8j+DOsZhxfsFqNkEMPG9fiK
NZ3mCj7op+0zao6rGWtQ4xQ841/tOCR9n6ijp6c7zB1EmH7s4M/Hjxn4Z7IyDxAr
dyz9bWl7DswGJuYcXLJESX1MOZbanveG0YNvvrnxUkHiXnZvIFhrWAClfcCkQsjA
+KftI8bcdAdJ2NMgMgrACgGHlVbrq0VL6J8x3tdCRVwCv9tSWhF9USJeHH3Qs6Nj
hdZa0s26CNxEdLQu95DfR6vkLJ2EQwUthC9RNnjiCXoxht2mXUajFADXLfGCtfWK
wyg46e8MaXSoXvTeQ4x5hRgm6iXVWYyXS1LQL+QCRROsNUM+eme5fAq84wK0mYy7
KJV1P1M83k4shypuy2XYs507Y6HBp8epqZY2rVaEGXcUTRes/GKtprs4N6Y0phsN
vPHUsn4bvakpDvqtV2iGy1t4E8QpgiSkvwy8NQdMlThegovRjd85L6YP9yqayDcB
Mo4fj5ZvqLgWY/OiqLrLG4nYYnbMlRkmcLh37jIZN8GDW+mjURAcl7ukNmN94DI4
WL3F7mhH07vAZwOkZztKQKbi95LKg++f7ew/fjVt+nTzlLwfyesWR4ZlYxcyCvtl
CHC91xW7p3U813DdEWRce0//9vuSYTOPVeSvE/DEQgiETPwE9+pXGp7FGwHcIejY
G4YqYWUdEkKWHSonx+wcd9QhbEk41u5eBVqzVGaxqD8EdMj7MQGgINz6eY4U+zGM
dCNlpOgSY41ylvShtMSF+1cWTAH9flxJzpRkqe1wma8Nytny3HYQsIW9ZD5e0PFR
WBgNNfZBdfrY78EEG4DZrNXjqfh/zrRmB0EHXkdGayI5ISHnAupug/jIpwf5uDK3
plmKuFyHtnM2/w9OWY7Kw+WKgmCFVl2v3USQu2NOsTkBcujeG4iNryFOT/LypaxB
9IHOzZ02/mLj57QdsRi8DETQgyJEzq34LrRuJWLfhU9kGsm6ViDUCAwtO2JRELDB
oiJHwdJ3+SUFBTby5AqOkJu7vtMHY7vVahtChnsH/cRG3yyNl8xdZktXXjxrUdaY
jzTeds9zqgjmZA3r6KG2wFCL5Mv83kcs1rV9U/FOHrDvB4yob0gDSmjO5MUafdSS
fZIEX7GScp/qPeRpPtGuLWpC5WF+xpeCC63sLAkuXER+1KeR5xX9iS8XQ8LCVbsw
qVSOCt3jVXyTagSk6ZVngTKGHB+dnSXrCQ3XdmZZuYxIeQd8vvfm3pzxOFr63bSk
dF3fI/Mi22gUd9W5nWyN+1oOVr90r0kHmtukWTHRa8Y+ZfWtwn7L+zXwatgGHEVW
kC8p7535x67F2ynk/gPvANX8QX06qImC2A2RcuDlsb2IFi3F+Y5ZNzqq/4tW6iZF
fJ4K49kLbaRjCJfc3xxkzcNCwgRKZJ6CWmeIl4h2MM0IVwQbYxmOJ5S6gmHYZGUj
mGtXrJiqqiHSlsVuap/9U3auye4eTZQUCDeGzmurf7VOvdEsGZi+Dew9hEEhtT76
2sjTyxUeRuLqD4mndaJyOtSmoy9ca8TGDV3bPBhQ9Nj7aT6KjNeGBzm99LNb75c7
TPyiUZbw+0CQ2WYyz20mSv/vLF/1xENMz2Vy6y0m3OZpqRnKX+BgjcXe8fo7gYu2
IRRgkMzROp8NAcCuFYaSEj2+BjqcSr9xKEWncCbgh/l84uvM7grnQ30NHQuWHMq6
v1DGhWransggAjKe7U3x4cZcyBgl2mpp1TwRDa8kXIxdVJ1Eit71LNt/xKXoTsJj
Y7yrFkdIh7bNIgIQpmOKmhIxpmdHIjdSNFI5VrEEkno74aUh2tNtfXt8Qr9AaGSF
CPqZ4dUixVTS7mUKHztZNla4LvK5LiGd1pQG4xlnQPxM2N166Dwt6dfIbDFHAs8h
e4+kS9krXymwtFQbyi8eLgzMazbt9MZvlLfEZj1ybACJiERATAHKwYpjLIHVQiLp
Lm6YWt5bJkWgaQhE9RmMIcUu1CoRnVyBPcVGAY6E9qo3P1JU93bBQz7KSDDXmBV3
tuDe37/9rpg6ODi/EOiPzM4DU8UBrNI73iLaAg25RihaqzoiN6IIG/IUwekOxDD0
7Zrk+bkaYqiUxgOWzfWaalfX/pGa+8aM4hJNemsOsq2oIXtkAh8IY+k2GME5PaPw
MuKoTSFHSTRNnjdqIHyFrGZ+rI8QN2br/4BsMtpnwUPsgsX5RV9vQE9TFe5wdJVe
j2o/iT3mMkIZJNTqZeGX6euhNvRs6BaNoO+pCDFtf/Wau40q0g+N2UkcPO6mBWuL
`protect END_PROTECTED
