`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ij+66iD0RTh9IrhAaBzcGDbR7nbJpBxePTJjvikTUhT9CQoJyZIN5isZJN19l8qz
Mw4zROhUlF4yOY74is3SF1TQym+1A2DgHCIfyR673WnYpSYpZbZ0SOHUzurmEBzL
KwtWy7Mo6kg8T94f5NQfHeVGbguWNzFt6RXQMvHN7xeAK/EKflOKxWX/2tqWcN8r
UMRcZu83kk/SDTfOb7fnJWzeXx5SLPJ49+evKKcaaHBexSeyTDgIo+rXuef7GTGZ
bid0i6QE2HcuaxIChYw3ISICUP2O5jmwl1XPXw51wqb5R7slErhb6xA3ebl7CFK2
Y2sdAFlC0IhwVmwwLGE4of+qJlxdr019upPWAlTiIQ3FdYXpFAI7D2SoBqXt0ge1
1Hdo/Kq/vlgj2iaUWbMkfjqAIxd4SjM/NcPo0xDmYzxnU5kIgAnzkVOllMfN8UF0
dYbACKzvzp6eF4V8742oZ9uiyz0IiSjviAMIDuzlRarJFfedW3bUwaWmWR+3A551
t9DxV7FhhTvlqKLOMHJ0YpKks9PlfHUuWiZUF+OW7hlQ302rehnz8QNqjU59JB9v
6s+Ktf0r5OtG4Lq9PxNW2ptJqLYVFsEj+IHq6R2DA6vCbQuLyW7bVE770UkLbeZr
RUfws4q1yE90SqUc0awVEfrBQAfIzxR7zUg/bMIvGJ1Qx/haAXjXNSqEDkDLi0PL
XfVJJxnIkOnXIx1U17+eBfTzEIaQjuRSabEi7Gpk7H0HJCmfOxf6wVeW3EHUA3wS
oEZk+XA+KugsjQ7y6O2IT7GavO0CDmna8JTp/F6AYDT0glG9QgVtNO6mFw0k5TWG
SlMWlrnfgiKQX2xCYdGeOVe0c5EbitbC1+Kt2Fm4A8kUwpqhms5ESkb0VO8kjSup
G/6bbL/KoSM21K1RSKk2GYGiz8Sa2E7adSzjchPQIT/AlMXWCHCPqnfNuZR0rDWw
4r9XEeTf/Sl5MxxZo8qH2KLBoy8XQC7H8sJxdN2/jXS2/XVyo0WKkSY/psA5zzVi
dWlGIYXuP0LQbOOmInVJYGpxYF24ZeLMPJiP/OJcGLMseKADMmGvobTBqi+oTU8C
i91ZyTf3RkBx8q1Uk6l5hhYfyubHsDBslINSdFo2a4wIiHTNAmI3nuv/8Dky6NVV
NHOw3HihUjPIpcWRoz7Jze5XWzznXXqCiW4OQKozezBmzOOPkJ3/ZSSuSnC1Ae5k
Vz3hlAP+DuPAP6+o9/9ChrdGHFxjyUr/pkgpipqy1OtFnvB0OIHTyXzbuWW9dzoP
cnCG4CtHnDFVLCprciCkOSSYMa41hYW8ULo1SGbf8fjXSwJfH/u7723tzgASsySi
riG2SuaXjoYMvPZJrgWgKyHkIjR/zVZY0qhKfemLOqBp133nmbJxAuAHpg6G+CZu
fWk06gQiuCUpT1/rLoSe/RpxtkvZ0g6edpogTeft2DAVdBXLzUXk9OPQuDDkCzLS
qzVj4aa5HB43BiEYnJTUv+Vcmz2z8YBI07CJRiq4d+L0r3lq/OwbuTZdNBNEGSIb
1OvBGGy93zdQPRBdo5/p8CnZkiWHx+G5m4Cm30MlzVVQxyTDfgfl7fpBEy0R32LR
Cfi85Sa/w2NlMvK+7rW1O7NDz+vP6dBJIRsjDibgw3V6u6HHLqpQkR00WKo2fW7e
dEW7vIgH5/nPcwgSPIXyKiofNJ2wfpn10a7yh0KDWL/BRDURdpYxlxNGrbM/cSUz
8KNMXwPeKkNTr3HNrQE1Ykgmy7OSA32x4G1IFQHHb/qJli2MCXncpUqMsHwxLwIy
5IWNT3pTVxCd6yzSTvSFhjNuhbWuAm/JYlDBQAwpeetBW4Fj4hWnWW/u8zmv74Y/
EyYgJ2KMVbUgTNHV1rf2hIblgCqfgHxfgWAqAhDIfMnUc6re1coOGegyvXzIcgWS
GTuagqDOPj8HFFJtUEVqp08Jn2+iA6sAPKAWgn5/Apim1BfjYUzKcSAftaSn7zrF
ApO2kJ6Eu/+tJHq/EJ+uRMkzqizd78ikT9DToLXZ23CYRpvJmmaf8xelWQzpSps8
/S5vpGxjGlksYS8saj6vg6pHxMTL7+zgYwSJYpT896MY6jmdY06krvpSuUrXe4HH
5lrgzXbSU7wt5o7pHdPjInNRonuNuIT2Gy3XGkQ36t8mmWf8H2Ql6HfxZdw8BEkV
M1tWCzOo0caACECCJStv+zuv7QILBWvusIsmLQ3rX0XoduMsAV4vDXC+4DSZd0FS
9QcPQQjX1J0Q8VuFaZ/rZnDDVL1ES4S+6hQccgBIKCP3x/SPFNTWiWnis2YRA3QK
CgbAFw43S5Kk0UnfhC+ipg+/7EvsjwpeBXrOJujo9cyW/5YBESdW2oTejf4YOjq2
o1+QgLNUVTItsijUH1+e1XKpyz1SHyrZ+lWxpn6ESV7C4pz3cg7dX2eXSeMBWyIz
SdlLRTVvjPKVVRK1QdL9eHyE8Abdt32YsKf+vkOzMH98nJoU03uNYkLINdoMXgyL
pf1HALN27NLKvEnxCbggdWm6gQhS2jkRpHDxAR+1+6WZZH/ZXACrvJrrUQYzcMOV
O5gSAFC6Oegk/EK1h2Z6OXmJQw+U4ZpYNLZcy12K8GIaLPdirjCb6bWyoXGF6Lt0
1KiX2yxKfWQojnlxOj1tT/pL+7BepseimHPJ+04Kp6VMoWNAOWK/MyCs0Nsfhw70
a0og5l8UnhuOv4W3keUmamY1Da2LSP7MiaLri581COxp4WE9BMwBeV4/awX5Kofl
2cZd1W/980bw+8msIxaAi+bXC776BVpzI3nbK+4nAqsKHEk31QEeL0bJiDlzc1Qg
LUPQUOhMPZNL+wjd2voq4BMxkKkzWqdY3/3OUZWsPnVTZJ/f/4NQtvsdRiKxhp5g
mIkT3xIf3KkwDGFck3YrwObmY+w+SpKF7odfxgkoMASARL7AnZQEAIRREhdgRCbL
NZZjjExN1CVHv4Nr9oCXOzXcK5AYENS4AeboxSzmDJpk0MSC0O5UtbKoq0Rv4f0H
pnDhmG/l6x/tptpuqD5/FEoGARNaZtlaza9Lb2aO9D+L+sRyRKZq//C8DZDxJXJx
+atFqrYF92sD8/FlKquFJFbk+K1d8qSQ6irWEWFL96tAb76JI7LKIykRfke7VOTK
BkBh2Hvk4FUhFWWygD0vxQjPxr56gTr0yJqVahRWvCEB2q60a15hd2oQxUvyhn03
ryRB3fheit6jJywrywRGB0xtcSelF54hYESrGU6+K0HKNxOolsmwGW2dIpoLVbN7
ooYGiDPMwOp7JjcIMNNkA4FimaTCxISxRFwG47jBmU+Q2eLSX3+UqCmjEFrfKVJH
6gkMFVUfb+16V4/k69ER9JaqqoWSHBlshaQRa1eyD0n6eeLWS/CqrFORwgOd18l+
y7BCSWoJuYgTHV4LprUZ3mxiLW++luKcpJIE3qbJtjpyUg022RReeD/yd9YQ9btq
6CEQisM1d8ezX1R+0soCmfdijeGZR4Vpxm8Kz9LjxFSxVNBdLTjNbp4KFlA4mtH+
V1vAMo/LSqzzbeX7H/YBqLfCqQPrU9HvfsLLZREUk3TKexiiu7iMTmJj4KuGLcwP
xntRNkIZ82j3D9QxmqEOB89HNf2C19FhuEQQWNA/MbMEgvB0i91hwS7PMhaoYBrC
1kWLfP8VuOgdplVvrtTiXQyanCynPaifEjgOkSEJMvShED/LaM++V9fEhUJ7p7J0
6F+2oDgtPB1VE+gv12EgibvzYZka6fX5hEWy3lWCFdpi+BL37LcWF22CGaQsvhow
CP3XOMUkV/tU23phU6XxOKpgZ5v2cpoOPJNq23xb0mnwXnG6tyji27KepQQdhF/k
FsN7OqKr15mcW8Ae/96iYmEzCS3ZTwHJb3ffzpW17uhiYE6T4G7QNXi75zn+jhpq
u7Go92qpK1UJvtNWSLg8X1BdgmvCf42V01t4jheDdT4UfOpMZbzi+frye8rzfmql
mKOWeRIehUhUiEY1dJubz8MPQGCPSoorZOH830NaXg3RHPeMt1UPb8d1BZ47Kq7u
S4b/S4/atwXtiFgRJR+oPfZNIkXgmBC+ZBGnklzJurGvQ99BxvQX4cnlxLJg5Xwm
kuYLEdWrnvJbE+QZU2O2lve4NoK5zNPeI9vm9B11tybkrcSMELl6RThxa3QIkPTc
iyV4FT61ClzvfqfMFLxxjog0+lx/lSuARfyt+GzcgI48xvIDxMsoGibYUe0cSmVo
4zaic51Jf5EzhwU+A1grfw==
`protect END_PROTECTED
