`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zUw8NnzxAyEPNgnT5Rg8if+yB6GNwrr2pxKiGgwo6aI5vFZYI+HabCt0nvhqFU3D
SsKM/yKoWGEa5wFX+YQN5BSzO9CdLH007Wvr9oznKIXssr0vgGBlqaM9WzFwHzZu
zHivQ+A7Ir1Gek9VSzyrWTjFWW61u5GspWFstijj5vSMZq36l2Any4tw9f74ji4l
0JFeMh+tYgPP/7hG/BvEW4DEEGRfTPnpbdfUGpP6Ivs/6RTISD2GrZ52h2KWwQpO
PVwyXVNbfRvu/pYVu7MjGyUHrmdW2n+SRhNGpozHRB/pHJJ68VanQeVOZmxezICG
ujFudwdL3Y8SnhDs94Ghl4stxYgxr1jthSGaiPhWDmuvzfxXMgn1Vr2prnBCcuPn
txVxGz4CSq2yeYoa5PG4BDf0ZatOytaB7cf/I4I/+/1wizwBTYKkZ/+G/9FGOKP3
t0V7rJkfU6QTGGqP2HszSmVmXheW/UjjYb/ynID974XTp3hdUHCRfs/VU5T0+SNP
nIFc/4OHVKhoCOUYsvSQH38NpXSWPHaXEJH9A1yi3mK3vDw8k+Cdg1u+gUfI/cxr
21g5v7oisYbDPyyyB0T3vImH3nbl1cKQQxwZ5EYhNUGAfg3g5BDB6FNTnDsbfgJC
qafGdqCGzfQ05IXN+xfCyxMKkBYoLjU2wwsfe2R/vDhJ8lKf4pMm7ObTieQZ6E4S
fPcKMHoNKj2XK88CUcfIPWKkBisfJVYwTupSs7meaEIpgldp8kW2R6lQWAa1ZZMD
2r1sHLCMgWkcEdqiw24FG5Tx7kEZQptvIW2ngM22Xf30OP5c9f406l8u3/+Pm7Ey
S1dziXx3FDVUIkJQU/K/EC1ZXZ8+PiXt3rtZyxfm9O7zTdKs13K/XoNlo/r4arKM
QEDblY2KCF7urudQ/Q/uA9JmaDt11NQwDxANJEx4UfxgqJjsDWOUDVnpNi8V0VMj
96alYZjln0hTSWSU01ZRDcaxiPyiJL/5Ww3cRPRgKRyv2nV5QfLwEqAKsAtOjjdh
mhv62DUwd4nswgD7ipG2RCVUrFtbz445LWjCCp/dLqYvW99W7be0jPBMY31cOFTW
5szrdiEa7KMFYWdRL675Pjy+URQGX4OusVCZSbHqRVykIEYt/CMp441vM2slTP2U
+zYyPEzNLQWChwMBwrSgApU823Y4X4CFfq8NvCbinCXyl0AdabP7o9zl8h7KBHnQ
y1KVBr8P8XtAOdReeEWtdwE78AOT1pWrUDJLHRodfbNIen0f1tWiBVC4guAfiqUL
oq+aPZNOX0plEvGfYUrQVusOmzf5jSynneNWpDAI4sFDDj0+ZN4Gt7xAOWnrBS7Q
mkVPlv9GhHhU7wot5s52AFadjz307TkZpcwGgMDnqEy7OU/JbgoRlmsrp2TFCppZ
BNBL0dTE6Sr1LkwECRL8OgJc+6R/SDaEAf7X0DqnbXg7kMAMXl6kivmyRYXxcPPa
WXsWPjpxZiZA1ZcjZywVBIAK67mHeTPgZDO5a3kAc3jfPvB6AiMrDRvjcPHofdNj
r75VqmqUPlq3e9Khn6RumtfG7FNSGUM1A4vwhxM3MvD2AuwsIerBSQFxdFwnfs+2
TW+cE5ZL1MUdG81bGS/BASA0p+EP/fw7xIKUQKSRcslYnBXcCpeOuLXTTV4sjOg4
fyXaLE3VotqBEDJ8eygHOyhFYTFu2bxozjnOo0ahja9lB9gV6xqKU/K+1qVsavpD
DhRnoSHHt2v04adgmgebULXP0ckLBBqn1COwrxNFd2I2Bd4OxyuIdshrqMwoYhlZ
fpGxMFp69KLSvY2TNbOFD7oLyEJeaMH9UbucLLhgFgzqz00fn2TOZ1LSNs9++koX
hHppug36UwA+UYX7qy42QY2fyaZpdv/11rxjMBRJHqMfedr21jOkQNn3fLe+k63m
q9U6JC9z1HLvzL0e6XqiQhfZDcF1k3+jy3goLjNOVUMdpcPmRxKQtBPc9PrA38N2
Xx8pPzQ/25NTL8aHeDhJ1ciXKb7HWHbfP2kn9gSplhMKYhRwl7AtELV2QFz4Y8HA
m4KuKoxAP0nYHzNwkl4RTjvi+kHRGQI7rHCzEthAx/4qnQniRt29/2JMhxqTA5sw
AhOnsr1k+wMiapw+BgXWOR1JGiD+5ZTDhwg6rPV/7DjRjGVAQmJz8gZ0mf0zA2qO
KVTWSES5ZmXKcjG//FcTt6dIZxg9Fb7myjvD1sU0+uvfwxJmapuOf7+vpzJCahNG
NRx7pS2ifgFr2VAdKGNECymCCNcOwwgJwL2gR9X9wzDsVpW6tJ0SvTJmrvQYCF/P
NuOby1gAH9eWJvtusJSjS62JRfeK/Sa5WF4ulaBvQJaLWczfRAXflI4mzvqAlqup
x1M5+2ZfdNm/hEve3l5eaal/yJdCcEZEcvPbckzG6tHHnUlnneCyfte7l9WGCLBY
My368JCP69i8aIiODeYjQ2GK2RtPR9K2iYdU3r77F52K4+kBW4CVeoqvK+6MfmR5
x1tXFjKBTd1GCTlLHZXNdkAvZTXkWUO1dQdfy2RaxqDeMZMBELPef/W9sGJ5QD1O
PfR3ThJSNABDgneXu31Zb6stDnbM16ZM5z/uAb/gOTKnyjZWtjOlwqd3epWb4QYy
2k5kFYR6mCNTo3a09b+/tTSr7wDrf6aVTS7AOYvHWtfNh4PtS3DlVv0+eh16NV/3
X75YJkFoG943HKO96v5FvYg6xpF39/TWpWam1Zgkt9qL6rXiWFLklToJPuCqr/lW
Wh1pSXMZm7TUxiMGXG2kTiNElxtk0db2BEFgPU/w3q3TAei4KQkt4AMTVIGDq4Er
au5+Xzd7OJEDuTmqLU731oMNA5DEEe0UKzFOfXCRuDzTkt2qUxqhJtytIwDPf4F/
AUVWNAHgzbv7+vv0JdYbMsHFm6BJm39IT4DQSk7yG8LQy0t6AKgc9HarKDZdY8bL
wyp67bGw5Z9y9BADUz8mOK/FJ1Tx6NN0t1VIvIvRDhp0YDg14sK522HU4OFZbERj
mjXi3vQuNMYJCWwlhOU5LDHv+g1Vhdbhr8paEnhZntRztPtXVEFQOwca3Hj4puS+
4IBZf0QvLnlcm59CQRPQc03RiO6VcqdPVAMXfadKh00HfjYh9VoCli82ZvMu7Y7S
p6OhliFdqRs0ORj6RHl33GqOxUd94WRHfwjlHm3yfpftEFwU2Jt8xcKWK8KrYTEn
XE3fVh/mHaAbMTorpchLQS625UooCvFUzhyaa4j1iSSa5hVvxUSpBa8vTo6gcsJz
9vD6m7A7tEw3v/Cp93H5ofnW3ttOOcJiqNsVbj+Xd0gRazZrimgoobMcDSS0sMcM
YXCqAkyuB1rbw7v87XQgf9oYEv929whkQOu8bJlz1KcKsqS9OLK9Q3QQ8SQE/mKW
xb+vXbxRgg08FPdxJpIWZEoIsr55+WuV0px+aH72B92HqFI2JtGKpOBs1Ctg2/z6
wXHex9XCE9QbKROto9XWWfzQH5xTjZCeKLtFYrm4DOcH0UYpqaeVCtkbfFMR6wuL
ivWUtwj+bSWcRKk6poqQUcwnit+G0MI2xkeXV9vfTWk4vhX4zljy//8qDU0I+CDI
S8JAeVZk2Qa6/YopzgmZnBI0gvgMrYiCUD9tuo8tNK+Oy1tMgymg+padVuObbk6T
371VuxZF83sFq6qSX4DWrVbnIid7g324EWpXnuoGxThzwaGrfiQV6f0caEty7+75
BZ4JSAt+zgOIehLzh02XLNDpd0W9lUgTiBUvcUCgv6vVKhqyhZEbGASCAqDa/i1v
JtRN6XzK1J9dMeUXYP+UBQj1uI+F4IpHy4A5s9jWI9rEsfyyzSd3mJQI3/xCy3NO
t4HGzBwq0csS9YrTPP+4RQvswU+Si3/Tmp7aswiza7iaQ0ZA2vVAEe5+zKkVTSj9
49nq7h9R5YVdiu9klLCuRC5RQ3XIOJycvJRpaP3rBFCwBrQeWhylx1EH7oYTG6yF
5t3R+5PR2trHY2fQoq1ayXlK90BvEWNu8eELn0YtOET307KpG8Riv9xPHWfwyE61
DLklohwoWBhYh1yUHsEWyXJ+NCd8o2ijxGGINPncalA2qVmdY426/PQl3ObiGahr
k0l6dgRLiMO7kmM+K0+F/CfyNG0iUNKQ057gIP2/yTkQjx+yW3w51VhQgJek9a51
2KtXVvcWlpstfAqyHgf234O67XxJJCh2Kpy1NTANJqJAYi0dNX8KfTC3EhCVSvk0
i1WpecM5kZFWEksy1+QIq6bXLACfmL3mkFsW/Oizv9rqv+ReiB95r4Crew9a4FKT
CiuO+bIwLyxkNr0l4mgfrgcfZgz9WHoZ/TL7DWX2QWPrXrVpSnqLfwIuQnL8puPE
i8F5rJiyan3+M1nYZMRb/65noqJClpT5k9jJbFg9cy/dfvFHbAZ2l/pU7DTPx01s
`protect END_PROTECTED
