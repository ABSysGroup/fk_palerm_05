`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qFj7x/e8YlUex7rx9uIzcIQghERoYg9XDoINSTHF950tIHM2WURLsEatUYyuh9FV
ECVOYHiX/nF/9lXUNYViJZpDYB/suqen4Q2jlK6HR8tR7YocjxwOavXVbwP48mhh
T7yum5OTWHU7yb9hmzn7mqhtOUf2eCVEYZICg8o7hAMrcdGs2kgU6L7PYfGeGRGs
V1EbnD/rksFzDY8K/IdQAXWwWo1MUXGVTLvZ5RcWdfR64AZ2F8LyeEQ4aYb/oJwf
KZSYhGGPX6h5iS0S/MOe7X+VoOQG+ePIeCvKeS+lovKD5idcCfYAsNaIdw6X8rs9
A4e1JNUskrTv3TFQ+TaixdjTDF3+76nUVZcElM1s7c8MpYKk89LAgfl2pW0BDNOE
uaA3d1lQajTc9vG1gbbD/eHT/FsMbT1dQlOURlXuEWpLPv542haP0adT0NgsvvJg
Eri4YmW1x/WijbFFVSrv2bpcKp5LAABEb8IKTMAHHBYLd/7Z7J8Sse/T0zpzy7u6
u45XfktQRiAWtrbw9Ey5La6FmXvTyV1Dah1bJFzLz9/zIKTCoa4csb1YsyKs4Yog
eL21mTaZl+m5xmlFI+S+VAEolz7Taz1oIYEoUdmKYVho84YsS0kvLtWrfRRNrnKl
8vQet7LeJPgVndao/pSyUEcret8EqDtnz8nVN5l6w2Qm6nYqKk/H4SSvnErlXKEk
YtG2Ps79gV0VdmtWInsnhV2t15GySk8wz8PTBoc2zEc89gZDrbXcsUUSJ3VGqwWI
pxT5b+5GaMJmdcOumQpcy39cD/GBpmL0Jj73r+kcMdRhGItbKkjdwh9fsE0t3RKk
XOfGaipRuhGm7DMjgGjzl685mJ5UTVOvImUIjKWGbqgE8EkY4XkzxHOujsKsdGT8
6HO9srDsjf3NSYLcYnrQB5O+joZx5mEW3G27rB5k5oZhqVVOla0fXoICfnF0dXck
`protect END_PROTECTED
