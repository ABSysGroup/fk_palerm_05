`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IISO4wr25NL4YNRiXRtz/bZ0kprD8fSY6HRlGPQHxR/I9fYqUwTtt4HIuvDt2aQj
QMdDcfBWXgtg5MpCS9RuIpP8Cggcxv0TpIetAxGdWLQNqRUrVBGlcpVKWqyhg7Vg
XKWaW0MIevrarXORL+5TFVuX81epPxYd5NoV5tqibIwlTq6X08H+8AZScdXRzF6e
AJ+gJmizQ56oISzxRGwi6eoA1TdFKjk+94bHEcdXCyLUD/jIPX9PB0alA0W7YTTX
hJT1h/LuKpxxwbw00JxSpy3x5oJRyIBwPbMSttHswQO+HHPaG4lhMVuFK2YD0PLc
bi40c9Ktbz/vScid2vg14ERDumD8EGgg0tEIm/fj13aZgIa3ILVApdJRvJP1jr0U
GTNgsTV07M9uPIjFCmwPE3UEvKeZHWX/AA6FuwLAzD4zrTXMGr//WdL0+QLZlkEf
0zG/cZhuyf3oHYX6jRvcYgw4M9ILc/2c/r3TwZPybjb9Edz134LCHXNUE+nEJfAU
pEmmf7+YlWUC+bdqpBnlxysAT6ij1MRq2kWyzblEWmCJZpTg2rMDRcsnj5gYrX06
1YFpuHbEqI0pqJnGFfgDL5aVSCTQReU69O3mcsqXbdEI+xvQERVJmbIVbxwN4Xbd
14/TCw7jB6NeiVllJlfXKwpVr28Y4Swue65vPE8V99XueG10x9sU2F1YwsNSIf9S
f9Rr7sikDxFpxy7FZfZlcbtN0XlEQijdVXkEpjbPD9VEJhItsEBg8dwISyf12qW6
8MvhXMhxWqPLemu1jbxiBqcqDVxtYoZj/yuRpBEpKdnHAJnDDh/8jf8dQz+ogb8e
bIiWBmxT1fYfZWqE95jWKJfGoL8k7Z/8bEvArGLaT2wIvFnkdBtRycYjUM+y8aR2
uX98T+CfNz4PPDsgDjm4p+YixvVNbGx4WMeU+t5nRMVK/iel4F8ueOunpEhH0RNr
spe+9SK+Zq0pqskxlXgPeI6cWflVPyn0HEGqwiw3W8w+qnOBCtV4dPYUzYfh5D6I
Kyj1ShDo1PDRSZVsg8bpHZovBBuzEP4hixjMxggetZCiEetzWpjtYvwC5BAHmNOa
uSs2u26KJAJ6Aa2HMdBRrI/Pkpv1a7yao7oGln9/zCsW6e05LJZthdUzgi5x4tC9
RdOQuctsuzBdl28NfszuBDx0cHmq6M7P/bVex/HDcVFso4cMaEE2zJUZVV57CFgY
mP4ubjgS8TQY8b2kpkp70emDlNtIFsaPtLP1TEogyNxvgWbZj0Dd4o2g0nfatQwR
MCSffK5dxMkzpUhWHGSuFQqLAxYbjpSYg+a6JEYif5YIM6U1sQKWUBdKZVCJ/RrG
q0Ezh9lQx1yJn84NApf08coONOAv+8TEjSu1lCGA8BOaJTK2y5rabcApkOIHgVJD
LP/Ldn6egncpi/fBXO6DT4S61fApmwpM5O2aiGNU+kjvXVcPGSN+Z8XiEvVBmmXh
3726Jv5p8rt1Zs2U5ROZINK074BM5MMAC9WmrDcE32C0OIaJsRtYvlSrVxnIhtGr
dC4R0xJJhJ7diwUtz+fV9l/DmlokWb3aTyGahVZw002bhHqpiWiN0duEnxO5Kp9C
RS+5WHWGG6CU0SgFEzzyqN68oeJOtg5Nmk0aTUEzgfk9o2hRIB3JPOL4QpUmupEv
jyj+4w5tOld0bZQpT13JC0Uv/qHv44VTODtxr4xckf1K8c+ZKfrwKcOmrIhv6UOf
lRRfngQhQB4Hev1DjW3b7U/5T2ayWPWuU+cwytoa4366HIezfLEJ+ACeOTMuKMx7
/No6PxxRBqbvWLisBPBng3R9AGsL8SZScB++Wm8HegUh5c8dEhVfr9dS48DAxj0Z
skOy+MCmudyh7oYwvg2t1oTxlAbJddZVFzuxdYMqFADwMbBqfdEzxa8E2VjD6Oto
8Avwb+FYLTHjOirjT7Y180EP9qMhCmxUJVfWCmljPVFnqrH4MmUWkEKr++/dby73
kGYmOduCpFp+8IMgSvVJ1AL9dl5AWVTE6aEU3XMl0oG+AE8QKf2RwAYiKd6WXYH4
5J5JsWIX89hkUuHUs/gz239q6wcvEjQbclz7EgBi74Zh2pMhE7b7fqqk0qiT3Bxl
wN5R4fig9LeqP8P52atZOkoGz6eCAi4cupn6lxLloAqb1BVvyRCHl1LOkN69zt8U
SM2mzViOjU444Ji1xJo2DnTx4H4X2qT6HntnKqkHpsKmQHDYfuf5B0JR6lk2VFE6
sDWMwUT0hgm2puB/XfAPJIif61w7oYpzpleXrzA8/WRrfXZc6fQIiRYQii638sNc
hLKrHOs3aNguvEAlafk6DUpcoMShkM6sx3KT1ZhMwe14hItHEwgF0YBRTkdUiwe2
B5+/L/0B12GCUIroxqRhEkLaKD71q+5CAi4fHMIsEYX+uMT7veWCioY8p8Bni31B
HFu/MwYNsd9wtzwja9GNDX5dKfmN7s1pFda/nsxnI+RcdDR6MB2XvsJkJIUcLu2u
VX3iLheJqI7RkD7DsRivwCrs+RyXLYc+EvxWCM9LG67I8SFF6IK3VuMB9EeX+jqT
O9JwnDWIYm+2dji8oWooRTwYCr3xLSJGnxWu9/G+9rAvQmgDYVPxN6xmuW66LYsY
J2JOilderRhb17pUMzovZXOe/jy9jWoKHlcwG+te7mr2roxTWU0fBbQ6WRhDL3JK
kgWEmfNzeH96JmM+Rj1ciiTH+nPEMtaKfLHZaIRtgZDyxzbqAA04lwmxnavDuM/Y
EbuFal774UwEQ1AAgyr+3H/mKKSiLbzj1qjOaanTrrvnRvw3oNcvP1vA5Osupk86
FymoQndHjjAVPEzicGTSc6HipBKw8ZFdJvPJ9f4NWD89mt40IHAKXmBKsYgB0YAi
AhkzTYTXiyiw+knY63M+f9YxNflW8qF7yUVSGYtshzH5K7IDBZCjVWb4viBPcCXc
TiRG4yWVOXuF5SIGKDfJhVhQlIs2rKS75gXX+acBkoHCMeSkGvW5DrguG8cb3Fj2
0Rf01qbfhTLABrxIhHbb7Kf9EUdhcJ73wXFtyPDyOsxotq6OcHDS+iMEFvgzmpgt
Gf40/+7qzgy3ymTLSBG11uUoViGI4oN9HmR8wL5ry/+FeShnCU6VlejWEq/ovuAr
Xz3azHRY46/gQYIDXoUeIBWHuzGOW+G7/ZKIVWcdxxM39fbCh+qyUTIzrcGK4CL8
ZqQfhB35JMjy+xJODKJb2Ptfhe16INNgdVRgjeO5led+Gn3EZncxitYpOvwZEc32
+DVquhZeg43RmtT3uqssRKoqi81g/L/a3KlwRp1xIsNMeCXMZqstBSE6g1w9eCta
8kXASfic5TgwRbSm9p1FnK2C3mgFQ/b9h7l6d7LpPWZraDtllMefMumC0uP1EyPa
dF/uxaJsTXoJr0Y8N2KwmTy7x0tq4ZIDWIYc4w3+WE3oLa6CajvuBLsuMFnMn7MB
VRAB0CI5C8tla7jteJ161kWtO6CQZUzbvfV7Gt2ApMUIdC3yChNvzWokdxI3lnh5
fye/dgv1VjkjnWkY/Pho0Snf9lUxXau7xRwGLdi50ZIlVdeX9zRl5lMB505MjdF0
20ugofubPuIrHQeZuhg4VSTZ67AuIRQUCm89j7XfsmG60bsfrDYh7fNLzEAPK6ev
9TwDCXy/u/xZIDQlOQFe/4yo/8TZ0Jj9Ps8LYoK3toA8pjGv7iJ+6ff4M/KBQ2OO
KzSNkyIn32gnjtWnDNx7zAZASJ552auVOqL0s4QhypcSsE+yiO8jKZ+klWLBLBSu
CCs7G+xVoPwXNDi1Ssx8e1lxFNsV/S30Cbq+gxfr+ES1VFYl0ZIeKib6C0+MNAQO
JVgB/GGC5cG3Q1riRRJI5Rjs9sERHkYCfCGVpMt5sleKJFNs4A477gU8UfNITlQs
MRcqc7zUAM8m/7Jr4trexWVYkskP8nLJ8HeJGQxowl+Q0B1+svVlEpaqbyUiVX5O
dL+dV491nObCLruFW4FO9pZKLf5B67l8mtRAGv7+Djt2nUmyGMbqwNjmnCxKyB70
CdhSy1i7CIxGRusEsRzBDHIXpOQ0l71DxjLJvNTI14PGOsDve8NYcOePDOHr0hMW
PhDLVsfCaqjyGEil+eA9X/d5l/g0wMI/MIjNHZiuoPNui6qOS5sRAS47HXbyrxtt
sejVM3+i+jTjuBxpwLJ6cZr9xfFXoiCH5J4bLf/OFbh785IlYnGpkmTUKkFDA9Bq
JeDRQCxFoxqCnT33duhxHNZlZ0WsF6TOP1zx0Fd0PIB6YMGvGnOhwwB7wNpAh5ps
mMw6p07OkdQsPwfbWn4Psp7a6rtO5FojeqBtZPisdMhVpgAby7Trb2QdTkN8+KcQ
Xt7OAWyJ10p7/xrbgLPJNuVVcz9bC4arQ+eQHl8BpzLeG53qJsFR799ScZfhhFt+
tUt6TnYycbq8J1gwn4ehP2C8EXnUKJWO9CV8rN0YrpUGYk4Lb1OFwZ+AuWhDxcNw
ysTE4bD1XqnGA+nBlC9Em8DeoA/9R2kk2gPbcfWLQBWf2szFBegZyhsDFzjCKLHn
l2FteYtNUQCLcf4ThmfXePRYOVzl+TSEnzwZQvYJ+Um2aooDggYczdeCbi8w8Zh/
/Mij5+zy+tGsocTJNvOhrM2+i1ztJybfWCB5pBVYuiC3Bc2/ENZxBCWfAXPDfd1j
4rEJ+FVMtMppw0JK0LWgWZZkAzeTg0rFzmgjxBiUaULfhOCFxNEpJi/8YhuruCgO
EmfNBp+gq7qjJqWnOZcvhqoKU/gjsaNlOqRA18ogFo+aXhVOyR59KA40/twI+nyi
NZXjA3H3y9Nv5cQiQ92osA0gCDDx1PGaxMB2O8JMVYqCj+1urM4fefsUtM1DZfFL
Nivs2BtdwOMEV9uM8v2uiE2hoFzvfErqFVMmNKY0SLKgh3gc00lY5G9KyvVuXJGy
ws3B6x7If6hyE19rCcpI0MQluSxmO0X/KDM2qFYGhNGMZwcpMcokkEEhMVLW6irO
OPPnPe3vcO4mrtBFbW6O3KD/zL/OtTJyB99jf6fOH6+/h6LtJJWBCxOmo4i1BGLG
e0C9hxkMq0s4OcsxURMgqHbN+0ZPrPKXu1mDeVSV7I7G26qy4yQpr9TYlLjx22nF
+zcXLL7gdAJhTVOvXTvNBrneGMslCyJqIFmL5YMQ67mEWuP114+1g0tx9DimBPnd
GIBpBCDpWZ30axaIE6sdvjI/5NuaquQpcs9z1xTL+XBFCe/6cvsbuTMKP/nsS1/R
iNxT3fuXnb4rFYOScGayxB1SNpRFJZa4dqzbAGOUncPDriw6lgOr1/13KHbP0gh6
ztJfPhksgvcdAxvVOEzoQrXp/qx/LxFUJlCM8iCFGj01kubthgN2O+xUohfwYADv
1V0olyp7ouZDGPOszsOzsapRi7h0NEblv8DY7FCy8oeVYHQhz6VDoPSzFrJj/tdE
P4YdPC/1CaIluHKkbaQkYq1iAZyGJ8cx4jBjKa8JO29keAxxL9qPoJVNxChNsCZw
lZkw7Gf8jymGVmX/nZl9LXr0cA5Wg7ygVnPAHUbZWTR6D3lrTQoDUa4LAKndUn8H
GOz9NVIeEfLrSld/JsVq7VNOmaCqYQmxYsYrgqIdc/r3K5vZfVHnel5kbJGH31LU
WmTyAkbCpJJ3qwsK7qea3YV+C0Pdez5f6fO46XHI7YwwmUMUzokNsZ0h9hfiw8nM
2NXvJJgCEGIknyzSy58tm9tmgLLhWcq4o8lmYLKpM4rzWrZU6o7RZqH0Xaz7ONyJ
OgekmmRkMzmQpSlPhjXNfP7pGJc1p+MbEnasTWQpwlqzRrTGLUWy7BtGMIgV5X/m
hWGt4KzMPc0lYO7ADK1/YSoF8Ec41sctIIt0fd6wVSvIENkI2+8yys/BfbCxiq/S
5NbQeMD8ZD1Le3KMKzRs1pExtCDCEl0lm19NQsD2n1cemLSj+yyaJ+YrR8h7AXdi
uNPP83Fxqn0urn5CkWQ7+LaAo87wlXUwqg2cNHEcbUsPREn9/Am6cuhqMliUpenp
9AuaZ78FmDphLq7MYohhURPmfY8TjUS7LiUgEFJkUrJf6FJcvbMdAVWMGno1fTiU
4mw6EN7AjhZ8k6ky1BvpBWVDBDbb1kMH2+im8NGo9TbfTT+oFSEpwWGMEqo9fzf7
Qcph16rZqYsJJd012ojls21bLLeypDoLoT29+1f0EQR0LHrIrxuhzjBnnjqPrCaU
FDRrAGPO174AXLwQQzCTcBcvecqMOunNyaOzxpJmS0w35JYkQ8uNS1YU7Lq17N5x
CFdbWoM7TQ6U7q66No16JiSCzzViVFNqwTnnFjPk+kksO6yxV/J6uG8XIr8BcroM
MUWkjuQ40/278LpTAK1WlaShALhjxZHPGoAtsiWERK9GmWoEhCh83HZ05xfpgGO6
753bc8rTlF/uf61cvdhZqAGMYdJa7WQESx1hO12sEhuf4J/JodPRWVddnsYObdMd
jiAqEFQlM11in+kPz4K6H/1m7OMV29h+oHCFMrFikUf8wZBTYP6AZJYb/EuEp98K
scEd0I9gMfgZEShv87B8oEkSj7ZtfVYqzxyyK8jdqmo2FR1KvYo2Yr2MrDCuIphj
Hc4EKGwyeBZC8BxmlXa13aRuy5sjv5eVantb/sZsXfTP34kKkumXseH65S5rInp2
vPN518ZiyXrR9e3iS4snJl0mjw+LrT5fEpSR5Ilj1e8c/lhgzKSsAEX/nx9DlK2w
aWPWqChkAqCbSDqZYCguZkbgcp2CkGEZtAdqyZX7IL4sKP6/B3kF+dO/sRGP18vX
dEYpUCp9m9u1FverBdr/ap4kiboSmtwB1hDbJ4bfGHL8z7+SIW8YFLzTXcLLHAeG
0xn6bUc73f70E8z+2Mq8NL/WKQ1c9ugN/3Qewkn7VYiRuhAegSiNctBV+HhaKrKd
MPxEjtZxdQWjA/GaXrbfPjbSBfH7Z9PSNN5IT3lyvrdijAuQjHRwtM3xRQt/HcBI
7455YXNifoZknu/tiXFXZpOHtd+lIwzue0XltFT7d6MLLgGMkPB2weBRa3sDIS5Q
mNAKUfecBNphR60mCfJiL9S4Q5bNIS7P7qYPi48HuAM4VP+h6nT8k9IoOKKA6EhH
wFUXFPXnOT0LC7pxMZqcYPFn1AqmxdO4qz9iiR82aeMi05VoY0tCmuLfJRt+OvV3
SATzCoZbtOkuCVYJjvRmjGb5ixRAoYzGllt1fXpsHAlptdR8ua4X+Jk5C+8yEryq
UyuZLI7beUwAJEiNak34X4ZF/Lf8AQD7NXrBzSDiXjKrucRdHlSVTiuub6aCQomD
FTGJwGBEnehKQbchQvoPH+DxY1PG6N2RQTc2CptQ+vleD9NTZGBnDWRxT86xywzg
`protect END_PROTECTED
