`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TbdOOQhwZa4VWyS1f5ah0Zyq6BLWqsa2UotsvDa9MnBvxnkp/sbWWlrCYCp/DYCl
srW5uu6ct1m6lbejy5qUVJMs74ikSQF/CSNOAuZ2V0ThC+AlIY+aj7JWbqW52CjB
0BgKkhrmNTSTielbc4WCJbAoHZktMpWpvuxseKOv14/c19DSL0aaUnSQz1qXI93m
qQjIFOZHAOb4VdDnQvCtRfNX5Zt1ziAGJfGZV14MAIBTqcAGUGzB4QBVan3gDXNk
JXvYqXlcLQh86rcRNoiPnW5zEXpm9V8czgVknEOK3ojLW+b8+O5OOEb8uvIraAFb
Qu5SDZpZ5qY4upAhxdQ8RKv1Uy3ls9Y7BhdIskWGaVERNL0wdmuGPfey8TiHNyHD
Sb4cBRG6jnOCXbuUXeGhmMrXW6uaA9Fb/SV18f+qnBOjEhvY2PTgUmNHM9xyq5hU
/J4EBZbiKW6cD1mpZjwmoEwT5N9oI7pUZy3rkKNDIuTtUQvXL7laiSyZ3y1wDUs3
fawkBFSujNAuNvtO1+h+oKY10+UnCgBUH6JGAhixPuPJoJzLuJ9MhVaW05EdwJMe
4CXxAH6nYG9iUs2HB4gQYqb3BLzf/CzEjHEanxjsftFFP1RHuj25ZQizaXjjAcV9
MeWw4Dlrgp6CLIZ+83frJBf2SXoJxsEZu0uwd4+ctKAHTS//kolWQr8BHXjGvwqc
UX1odkCty12zFREaroUwTcXI4M1L6SoBCi1f/gwY7vDYUZ2NzbRYJ+W0bEc4Pr8V
QvQLI1lTplhLGnjVNBdeRjYdogpzgMDoUr+bun+jWAedOoVBgd0i83lVVzZWndqg
+assoGJ/q5vyKCUd6Im8ffYYgr8vy+h6WJkIZUbKkLMEqRkNOZrbotZlEABGYMWq
1awCBtB7EykJElYKkgrOeZm4UCEKK7iqRLfPuUdGHsWyn1oiKF8982gkQFzSXjpG
IZlz6bD6k1oWFnhDFqc6PZYWn4RFftiGKV+XmL7yXDhlXXe9UNMLuCWZyKWBwUqn
D77UTejYc2EL3NQhd8qJye69mH6+AauHCNWpJ1KLXi9iaNUST6idt6DGFIcQLcBp
lDRI1PU4dbLw9K32z8dmc94sHP6mEyiow+ue7hzalzPxIkHGNBvipuG0uRZNGrQh
E1s/uqVrECGO81UVGc5jP0UH0NWHZ+7aVPcjkl5JkRZlGrr3/tizXOaKsVta7T//
vEgUCN/CMPHO8FobQexh57vjCYRSxjL113r/k+9ndo3JdxjIuhxEV/btqP5vPyWF
xYX9Fgm1r+kuQFHKH2FqmTee8emfRc2U6Y9mnLCZWXgRg2u2bkKDGQC6pHpkk+CD
HQvs9ESfe5y2p339x8zfg0FmjdAl+OZJMA2ejJZX15gkS2O4m8pAyEE80BhyU6HP
Kw0+vAlmujMviwW4i0LrCnTU/6F0oktXgqvTff8vQfRcwobW0XwYgNJnewNi5z1C
Q6HXxmXetkZKTA945ITbuv7a3zVtANDgAXwtdL5XSKC4FZPP7wzo1yMI1HpDMbt0
8M2c9njEUKuSAC/sQKtWCBEPRsi+eXUbD3XVK/iaftaSpmt5ozu+eTVesZhRrzcx
O+jF94QgdWJ1EoQyjpydyJCzf+gLCpM4rNMIrjDwAo+buspwZ1muPgVmStRx8vKt
hHgid3caGUHJKns0o/iHj59m+fLB3BLPAmlHs8aZpdlP+CkIvO34se8FrDfwY4Oq
klWnqagchoeIFjr7R86mcpLEF1oF3ItG7KsDnl8+isIYmTQ1zYNqF9M7c4km754B
FNuHkqbcCskTAg+5KqZQMki3CfdaiTMZ9nT441jgO/pf1dy0/RoebpEDXsIQiPDP
iJ3vv9ZRCkI6K+7yBiq+RAXo7N0n4/lpmzuFkHYbTWCcbwlIvVR1e3i4yVQusBZ6
dlRdjv5m9cha4s/ZRUatWaRxuskcYf6LDv/2fJpoXsaxEt9T7P86HlH5wBWsmOaX
Huwz1wsNDiL9SmhOsMaemlEUe2ND/0hvhNX06ZpgFYTQIm3aZp+xqm0OPVPH8Ks9
/nEzR135uKXiKClraNTEyPzhmuIu1ZfgY6gzQhnXS6N0XL/q7M9JvIFsmcWuoaUg
6c8fR8aauFROFibhrHaFg86c4HuNxERIph+zBRTk5AHBWNESItqbk8Qc+QRJ+wtH
kiaMEkwKopqDh6bbOFAvDavcLVlQjU4vUOZIUXQgMs3+wgPE4K4zZY/LxZXVqrWh
xo2CqFavt/Sq+KIpcjJH1HXVcapBzXxmHYvZRfUqgVHj4FCXqC4eIL+KQsVMvu/k
NHHC96PO4Yoqq7TA5uqYi3aGu1Ol+/m3XSxdJopT1oq8RmyTqA1XcjaR7NQ2umNK
lfqyLZ61R2OT9HkTx7YLmCBzh4ok5jGkvbMrQSMTQDIaB3PhZoinVgVG01SdGbcP
BSOyYv/guLIVxL6gKU6iGxE0OCCU07/T3432XOqjxcEr8igPPmBJMH1ig1OKiPhT
JdMS7dHDqVH+Kz/8496IFrWe+GytBSZ3MiUlEKgjVoBingGFbMJ7UIo3s8ordFxJ
LYcaPy03GaEbONxECc1+Ft+qRp5HnxWtLkL1yfS4ooINJ79n78t/WSG91EwCFsO3
Hg7o9gjqwl311fDD0Ov2gfBQJnCNtwio2k0jXvp2WR9voCvg8f9AKudUdESwZCJ+
1vaW/B9QAGMuOGnNfEVPGcP/JslzoM7VsJFkJvlPtS47/gosE9A/caxC/wzb4TPY
vhpFI68IYebkPsGBTDCpwwLm1bXQnOuvwrl9HY/o6NfbHjRBNGyFeRY4j1JNAt81
lgmNoUX8vCPc99//padXWKzjJwHhgyiGXjUKq+eHB9GHIu7UApGwrL0HebZ2kj92
bBWe2oTtX0zXStabqFc7f090av7inCtIhUa7MAxci+CIiuER2Q1cA3e3sIQOawCr
Hc9Eq5tbNK6nG/6eKEDfTWByV/eEUFsBGlaUNpNgM+a7JzcxJJ3NNjgon4+zNoFE
JU1w7Pw4TGmCeA6QNg0fjKlXFX/UklLoZjUrEfL00IwPi/OmH8bXwmDrt3YWxaMi
CWDfk+98m7mnjoUa2eyDtc9UliwxowdovV+OxAhbbwEyDoRG8oYUT3JFFZYsoAub
J+rvR85NYu0GiVWvD/5RI8XwTVtL3Ms+9dCebumLnkFTBY44Dcx7ZGyIYLj/zkcV
b+LhhWGs0t/n6A/XQotXQ6Oaw2xTqLiiPqxOrO6RUojsJctB3O0RBpUIjbRk+Gwq
5ug8dv0vQDH5yDX7kFnlSQr895eSHrAD8KcYV0ipmQBgYwdyRa3tjUg2fE1OFUJQ
SX0Uu1CU9x4nh8Mj2blxBE4rrzOKmu7eDtE27GbcNKxJD+ici8Dx2UYQyenQofDI
Su0Ll00tGw1SBlQwnjxNzEDoU77bZC8VeyHWjtOCwzmOnW/bp7zPXQf/z/UuimrJ
uUDMMG5vc2jw9cGOjhQzCjUMSuEscNcdh7cD8T3hUnmYuMIYaclfGBCEVqExI9UX
/cjHARHgn8F3c2ZzaC9Q4/QSMFmf2Ek1D5lszmcbVSPbcSdNCTVozhPFRyjg3yCR
oO1Q4KaqfTRYOECHZwl11sjmhGI9hKu55O3dSBKWpnXMyyRuiLziagRkVHp0NQ0q
s+euXVemwufhTEYkXRRJXkly8y84IoKbmibupVnMOyPr+uc0XJYWfAUUZVpE4AsM
P3lM7vMA5mXdwkbc1VACkcdROBwDHc+f6umMMOJtWGqr9fux3sPzNnh/la9+W0Ch
foqtKPHiwuuiT7vkcDI+F+sCvunY5+P4aPlhVpySiPM6xkLIawEW5HM+JM6mVaOO
KJTrfQyH4CYP35oA1HdaITSV0jiTnduGlymRrlGUNLbYQxtKR+KMgefKCS3Q9Pok
PcCGaahXTNqO4rP2QIYgaqm3DjItP7vKCi3n1zx/3sICB9WjgRuMEuZPPsfAeDRN
DaDMvPFiDsIxFPbU8pqFlUNuh39IxmscnjVwgGSyN7pFgncorivmhWDr4Z/kU1gk
fV/GWQGwuMwRVMr/emp5oN2ZfonNdiYeKFWk1s2Q/fEfG5m4zaxw0N8B+6QV0mCh
DXgJeZ7RKXxq5/YFi8KkFMmc99slvR6hCN99G+PMBYtjmnexQu++O0XKMnBJbfZ7
wWRCGWAmZOSkP7ENSTaFtHi9/acMNzhb698dy8aStB7PwrYqib0CuIClDtvBNtyL
qqrsREq6KvqMKpxAqEntxTyJn5nFeH1hauEiyzt3ek5jnFFpqwQlLjP26aHZhRRP
XE4bzF3ylewPVhsTZ6ONiJDdTuUX3Fo/1n4rBB9/pF2nvb87WNokjQiyMpUUdFnc
jZ5eueEs4DjdKjciytG128WatjzV1H2MIBJOYj70uD4I2PaA+6jv7nuCKuf7M4uQ
Fni8T5IibbwYI4D7CS0PrT1E3M2xuZhgar32krLS6I2fI/I82kOfD94oQkSTaLmo
q+RJVPGrSMbAl3FyNKrBETu37zxCmw9DounvXBCDDbT6l24848YF/FRbnfg1Qk2f
Q1MvzHb4dyPj78KkpKEzMPYjjOowcOMCQtIRja6VW3SYeEuZ/2SpGzduLVr8yeAl
/Z/EdclyZyp1PZ/JcdnXBxNbcSK2YmhN65xwGJb0swQpl/6O79daiIMumKZmcSUE
PNMYcLTO0+4kfJDvMwT+rsNh5InZ2m+PQBwEHxZvIV0lnlj0Q8nzi3agGZvc8aO8
oyD/hRSOeo/5Q+GGT13CxeGCq3HTcb9/JfHWuQVo/dVFYrN8CNkQMd8jJsggjk8h
ckxUYU14OdjLM8zbH5IiBu+AkheCblw5GyedkJPJ/am/1tYlV05rWWaZGIPcFbhD
uafZASHuN9ACXLhFx/9eWPlwmjCQYFmJsk7dXTd8osx68H6s8NIf6huraBles9Wx
C0Vz09a2lyaZ420PiKfaPg==
`protect END_PROTECTED
