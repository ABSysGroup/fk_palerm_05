`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kpFAdlZvvMHlHEZHAZ6HZ49FHQrcIfUdMG/Wpg+apAR+CLkQqAAVFEV/7bzUO5Zs
bI/Y39jpfYQSSmcFP13G4M9r6LFR5i/TXVX9VgX+bvRshrq2N+b4gpl5Ekj35ayD
KK+kp+EyTKTmVkabZr254LUOSADM7dlfMUBSlCrZkcMp+zb/Twz/C75rkM4jzBf0
/e4g6PoYs98q550WpVwYkxJ2pH/n9qlcXPBTpCTI0MrRaRv5JYwoEVPbqMGsJW2z
+QxcFoYAmmQwihhDSZRITQ9DU/hcJ9skSJq8mxnWWwxFjbirQDMbOvCfpgY5PV3R
98s8c0KraFRFm1kHjP1EaeO+njYTpmbVMLTJaer7TB/weot+CrmGrbMqwLx32ZFf
WVyHES00pIoNudA4X/2QveDiCRTGc5OdQ/+AQJqmgWA0DH8kQXrvH1qMpjnRAK1V
URX002LLmVsj3KjYganB2Se5Mm7DhiqSBbfUofvyDt7WVbJ7ZCENkSvNr6K9B6M+
vckyJgZFcaPgOCBpiWSzz/b1gw2i+hBcpXhyDZRE5cD+UXKJXBXhP7/fOD0qiSBa
3ZxWiOd8bj4BxKUeklhfNwsgvyqEXOhbPI3wuyvYn9GV62TPhnfyrMMSIxnArC/z
43nik1phTNbJBd2Sr1DFT2HiqtCCL35Hf1EugH94sRer+ATuxEr7wOBE7wLEGxUo
vDVCeJ8tU7B/ay9pauHxUWVausj7G0fOVMLkKPB0Nn/msP/dsTxn6V6SlMRn3HGq
pQ3lDU1f8g9Xxz8XRisuu7RgOWQIKXoaqaPY6IAAkoMEl8r/CGk2qa8Q5I7GAzqs
KbITqRwNsB3vwPaK5I2UUjnRq7srUwT6OVuJNbqTXlmr/2Ck4I/vIQVDIhXkwIxT
tRB3JnqHTGGQ6JSGzKIgGVj7cFR6wp460PgzQuterxmJNSU0/tNICVFkflO2F85i
dqpfYLPWt+HhtyONSxu8JjO4vf5sKyBzHlyX8XuL1jNMJLl1XXoIr3mpxK0d2hb3
Yp72dd2LoqH3NYOAAJiIm1tPaHRmMmKaA7Wj+Xev72Xb8ApdK8yLj3zAUYtABuZb
IrPf7wMuDvsmFkDNirEnaupAy8S6AQQVAr5Wj8NtDaRf6Rbg0hiTGpcZnyya1cTx
BixHqVc7m33DehOZgjWJGdCN58BV3co19dbckzned8vCWEkw2bGsli/eYWgnu7Pv
6OVAyOTSzhvQWlchU9D0ufGnmjtZEzRt//+ITq+azimM7Eclz0ne1pXeNOcJ0j2H
RwDXDuaBfiIyRM1xs9i1L9rp5UlIYpdBqLp+uAZHQBTWjL8ZLpOMvz5mBGTShiId
IB/f8vv0rhUMkcItb/aL5Y5yO9ANI8KGmgQytcS2Udm6k/O2i7p5arvKRn3HdjF1
AI4z7fCPqo8vnmcFz0qAjamq364gOa69kNsH/ioGbFwthJ7LZBddGJXnYgLc/NfT
3gepWjPWPqq8aSpZOx8lEqHig+WectnQ0zQ+ZGVzw8A+lS72SH9jJXHYEAlljl3u
xjmwDeUEgg0UqjEZl8u5j3PZxp8y+32N2rMIe+/z0qEQ05oJAxQm8WOFiFUtWLXL
sD8tIdokHA2JXklWf+0TZgxku75HiV0kJYkEgrOCGR46eE+tDy1qIWhQ5pXtJNOB
jYjkl0iyCqvV4OYKefF+3VkZAFx8ckT6Ji9tCWD7IDfazWCoUDHPr5WonjscGHaT
QbIdtmYfR9d52jD9W47j3h1n580IB5LFXEwcF8kj6giUSXm6toxiTOLOfp18V3Tn
DFMhyW5QcFn6oE65A373GVBDLzW17qcNb0gWuygSWNrsxbXh+3Bl7kVHP3ebzTAc
WIcM8v0jKy58NVkpJ8g3K9g6e3Yl5lzct78kawNEH0Y+AycJ53oyhJjPuzSLRT+h
14+F3YZKVRDXk2iWl6dUHlphOC+DfiRamzEP8NWJoRouvoVmja4UI17UPhgPx3hs
jcoqtwm5Tl+ls1j8k79se5/nr5xMgnnd6zbKTR4EV1V9wplnTAbzCKjNwBRRbovp
Spx1x0jHXtVuonViINBZiCqa4f3xaeN3JydvkhzSHIefpbFACeJ4ICwbUvouEoOD
Ar+at6+GybpE4ea3UqVwKQg2j93HFaerUqrFmhj0jZN7oFvRWqmfLtLk+qQq2m+w
UiHAY+pUzhIitAM8CXj7lf83HODGEx9cE8IVY8eR40Wc9nuuczvvKBVShfe/hsyR
2z55u4Imbka9s0/qXJ5nCJIPOHKVgGWnfdx4ABdu1BBO9scq1fpq8p9L3bcPypWO
3/MxFyyyp7OPrGV8xDzMstqBk3enPorH1QcqfDdvNuasbz7r2BZrUnehRjd5ETIh
mgtFqG6HLSYIxe0I8G4D6rSbX0T4yNuh5af1r+XwLU8b9g4i+KsrgjJqIt9to58g
DcQmgesmA5B7q+YsBNMF/U+79cv6FtczvWErVHTaArmZMu+PyW7U2agFXxu8FPcW
zFG5D+ZJxW99/gX4OLDLbESpEDthIaxZ66m0W9wMDeamR+eCBTWElfssvSybN+iE
MWdJkf2G0sBV4K9x1RE3C9bKu7T5alML0ppo2qF9aoCzxMpyO1wNU11v2oQt/vKa
Hq33BwtpUEG4Srva1UPGRW9GiKLfPyJw/4E0SJTZ4U/Iq4QnKsmVsYqt2hZveg5C
w4JOmBqgC48tOrVQCkiOCTMiuAfAFEBxG4bc16gU6TfRxB50pH8z/XFch5KCjhu9
AzSrZu8h+oWhG5vEiCD9nNe8kMMrMPeUXm9xdQGaiUZinIL48EBlyceC0RGw9OWi
6DLGzI4mGlijlFDkMb4/cFfX2/WmH4Req64Y968yl2M/ZfsMcjC24puJX72NdUUD
AJ7J2OVNR85gfAtZkep9ZqCW0eWozd7Lmw5tHCI8P7jlf8qfMT4T81N9F0HoHCxH
jvHvkc+oLa2cIxhGsGZlSb1K+2pdHjpbTRn9supBGi0=
`protect END_PROTECTED
