`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JLdlAcKxNSkpCjJ1DcTnYSQJSyKTpxnD1ZIrWc/VGKDOPIQfM6PdH7DssMLZQrkR
PO7uhZUXlVl4oLExMd5O7SLuLWBenANqYezYcZ3LJhWnRtmUysslpYvvHH7yqnCU
+pQ1Fk47Grp+Guzn4k4YcQeWqq5OdWjJYz4uRSUXQVxHW1vJTDagGx6WKeVO3XFs
/WVdqCjM4U9bpAV0vkO3eCzghBgi/uZcbnNN8DWbmK0M7sN+CjNy7xXGneggEHYG
K6iCFYPiV6Gedf7j0C1CuxA/eXJC3ctzyQTfzZSF6rex3k+gW1ao2rId3vQTEz1U
1jnDMUNGHEWMz7FztDCjFGFEqDoCRQqfNAt2ev0RNuf/I2f0kQJyB09GFaNgTvDG
/NAN3fvGeQmCDxv96yzN+VpHfLQVWLPC2r6TXW/Uy5Cw5KtcgB8H/X2cgym90lCi
wIS8Xi5rwGZM8gmuJn8PELtSq5BdUr3Neu8enEhtopKXh5ljmwNUnzne5Qm8eTqF
dpb6tdFlMPnpcEGeFn1fRuqV6Dag2KoieWvgp1sgbPERmuD6cpqpm3+lgCdeav1h
UtaZr6jRmF43j9KULtWSxvGdq8DJlhQzQYJ48I/D4sFkUsWO5IZEU/Wtj1o2J11M
9J1sZAkyRarA6ds0edbacac5Q6xLWjUaEZ2FEQnzx9oL5/Metk2fANo83WmymFbC
BID1K2qxPU0JsnXMtYV8dI4h7JfOD1roiIADGG6EX3i8Cp/szUdXUsVlTimj7vBH
05B6zEPU4AWTjYI+GwNRFise2BNt41WEwGZjtBAPcwHbkJfdVtKCxj5LjXYs/e9x
Uk/9ZBlu5Cv/QCPpByJ2udAfyVnEHyL09oVvaVuOT1R9gIDzrFhA2gTYi9n/27m0
cJm1Mdaaqn4KOleB1+X/EPa8USSHWPHKuEEBscwlNi+1Cpb6BBcyCiYFFtYEFUPw
sYR8NP+ftuByRUDXCbpNEmKJdqffyssOSjzkIi3wpY0jhHkMVvxYISyzg3Zmgjmj
fx1WENHVsvKLEKPmZaK9jTrdkUQ1WUac+dZT89ynh4ted6OsVPprsvUXAH1EnmXk
jmbWFPC3tMXkg5JDiTcK3Mf05LsIE/BTJwgw+ZSZib7qzWIRGCRrVhmJvR0MRxiy
ZCsI/2ahL2gXZL9hyebfLRKPMqjVXlUwZ62gSW6kkTNIt9l/zaOBPGZYauKt6DPv
xkAUKUe/FmF4vbN/h2E2hZq0bFQ90Jz75ASJfUueEVjARkM6vVjwvS/WL5XafZ3b
EYpHpRC4x+84pqNYY8B7m3yTuKyw9gaCmg/bCUq6Aud5sFzOAuJ3U+UlTRHWGnZL
y8/TtwjaJaDF1sRYKoejQyMEyJChZ/93Zid7jz+tdSQA0PZhoqQSszJINGbXIJxi
2ewFd4DoaYU6VPj5OlkQZn9LDdZb4UJyFZ6NZ7x33cjaLWxCSs71oD8dpi9T+W89
flqAwoYRPbOV2r9RVURDv2uOmqV4vE6cIMjCLl2kJtCWURVcqLWu9YQl3blEdSaB
vyo4FWWjT/fw4lKcdtKar71B559SDFm0JszCjHoswUgJhTHda+jioDT8WpIWqnvc
a2RUmJH46NmyPeUVfijLipX73dlEa0a+smZ9qmj9QY66vQzxBekYAuMZ1gwLFytF
fxKQVNYQ2zOkuTckJXsydrNAANoKtC3Yg3mhp6HGErFTjkZMQ06DYe+NqzG4LhkS
S5x/gW8nE4Dcwgd9c8gTYYWsuS+8PQNphEq3qgKzOQWpl/DNoeRWgG/HARkGN4hY
0cmk34NTbGtEuha8oAmc2zV1ZveLarj/UN1AhYArIdsUp9yYNRMvFPl3lCDs2Ryy
/9X4GzWBbRFv1tf2RdpMpYdW92YOGrowQ55O3Km6BNauGLRI8od1KUIyeic78Xoq
EodwXJ8B1jEH1BiEaBKiLcAydNlwGAKIcEkLGUohZ/rS1zB0NrNWzDNJ3XBBvJvv
6p0f+kbx3UkHrkWt2IkpLNLrOG/Y3RyTokRunFw17JvYEnDhADvoB6fdmWZ2AOtx
i7NPNZnm0g4A9yQZ9zz5ZDW/lFd8kuDTQQ53styQFH6XMOGIcBeFsLJMX5kWw0fi
clCJLT4oVPzbWoC7yWSjzidaTRyV84cRy2LrfofZGVaFtBqKdNOju2hUKej+Wa35
lKfIhRbw1ud1lVtZx6oqGm32tAHiFgq9f4s88xx/zrAfHBEnUsHilqOKGs1KTqvf
IDoraSpNfyxVZ6q4/+sfTOurhn3UhL217YRe84KeBaOcp6vN/txRg9iOkX6UTXv2
sCnn6x+0lSJJlLjEI84Z8BeaRGViQ1Yyh1wv8DQurYq9EBbu7aIc26kpP4lIbnHd
+ef2YjKl62JoqzzkEUoJMXQecThfkeghyeXFM+qXp9o4KzCaJQGQt/ZuNx3BdtKY
drPmOWf/PNEdisY+fFv7+uReCF3VDTv8utny/1ZzVWElLhHCov+Gozwx3ThYvYpW
I6prdJjHg8hw5C0VYhP3IkQgc1mTDrEGIIGFsMhwaZieXOItqiBXwnAl+xuWgg3o
YxM3WTS412hYpgoV+g4ORMO2BmwJByy0STAcqLcN6UfPQO7LRHNADOdRpa3F4gRU
hnroWYuLf88guJe+dUvarYgd4Wtgj7NY6HPbQ5QDZT14GiZnq7WwuL0Wwiu8etUD
5efQrO5SRf2KB5BgAHqSNAjAb0UQHKbyS22J689/HtCy9xKNBpVTcKr6Lt0jrahJ
+OXkfr+JvKcRxOr+OlwpRfp+b6tHaCdNrD+o72YYHvSSyj2jdyUpvAIAbCMn/nVv
tRBCyW/dEk7wi0GeIdd56A6y4veLY5PcMgwzYjNmimSkj4DHD+dsP8u5JE4cj4+N
xlEmyo/MmdfKxHOD2BCTyQd1yeDS1h5G86EMsI8ukBtCAVbdfnwzuTB75vM8I+Cl
0tvWh34tMFMmZA+Fs54s0gEsYafSJU7lEd+0s1MqQ/jtK+XORx5NNzjK5AyxF+gh
5fxTYJ8kSpL0LwGsceGmPnryRzqY3DrJ9Ca5cQBV/LlfBr4Qk7FlKfAu4wekY+W8
ym+0Uhvbf5gopAW74jZWpVUky9+OaWJIUsIYXR7oYGnzsEhodfkxHmW7BIxexlxe
EbvhxBul63QihoUjnNcmPAmS6tmGoEyKonSYu3fnAAtnx1tZf64MJk+hicmQpFQS
8dVoVJW5HtEFBHCBBWXVQudh6lnpHDFGDkFVWzqrL7zwBVMNYOvbB06+59uhD/Gy
HFRxcphjFvugaVNq0GLMjsOzw5/SJgBX1FVRmjf46LXzVcurIgJw6m9o/ESRXBFF
J7qcCxoZ82JQa+j+6t0Lt4okg3iV6NimcgXVXwyG0iHdmrhMwv/E7RdFq2NDf9kk
FCXOPS6mkE5ltlNkXQcn8oPlSK65fGTNL4KQx+xg7suQZaJY2+RuYXhWgVdr7jDw
rTSeaMSN6tRqeMczgsaNWti4V3s69sdyT4BJbhTe15qBH4MlJK+WSBg7MgU6ltkD
auKRJwbBv4lJavediQZY8wqyK34cF7s0sqV0Yb09gHxx2ApL4zfTqe9HhN7ZEOjP
B7fFOlcDllzckcBjg6MOVCByxyKbUjtId764BqRHWkpIPdlzsM3T3fLs5Ny82bPZ
XZLGdBC/b0qejYagxttiUUlxTHEuJh+QQ2Z37Y+5T1+9nOJ85givExmd/uO6LYRX
+HnRSFdNNElMrX8To/1sI2kM3ZrJ0QI0MQVM0ABgbexm2KLstMMtGGSX23at6u7x
jmWe3lUgdW4uU4greDLl6GYsoUSnbHx26AlFQ1o4bqLriILRkdE34Jhzvy5cAfx/
TcDuWQwtwpjEcJkwE2KjqjRZ18l+7F4Zf2SI9sMLgcouaNzWiJxQFJ6+NLZaBgP0
H8MCfeUfl6Jg7vrkRxMd3axYCgCiT36XViJQqoPWTDKO86xrEW9dMlsjDrmXB8nX
lkgRxYnvrW61tQAt1QlUC0tHJ4r8Vn7pu9JAvaWaNO5UT+NjgHWz2xCOFhbxzWmS
WCKLOF1UOxX5V6CpqBZQf0I2631ARv6CZSvw8zhwAluyjDZUqS9x3N7KH0yl06hw
NykrRfXF26oEuYzPMBA1K1bV2PNhSRArMG9qf6IMdj8pXnCC3hP7JTz8hmhhnHS4
h7Wb0TGmt9ta8a1Ie7E7NIHOehA4FYYGDhyc3AWeM8w0dEerwGwiNDpvrwEAzRWm
Dmxmt/VN0JRmh8mjWkodSATgATkaE/p3sWEglptNVNxHt33kNE8ct7hZAMmgxluY
NC0L45tMPj8JQVit65MiAKC4Qaa/bi3phpeAeVcMNI6oNHty39PgZ0NzbKsyG2By
ZKgmC89Hgg+KBh+n0rnSwZyavhBCwiblDfwwJzwvqwrroSpast928mnSHK9MZYCr
7ElLU4TMZo9FGPilMYngVb5gTZh4BlJeJio1c3O0fG55ovjSgl3Y5mpcx8BL2WVr
pHZupvwhavnsC51EuXRQkOPBkViHKKlI6YhJOrwLfGSeRcKXe8k0IFt3WUY8Iged
EAKzsM+j9n6Oci4cO7C4fodtFxaDkwrnGncJS+eeMwdLWSK+z2KFSoa/n3rr/MP5
2LNADK4AmnyRvsfpre+HpE6TMK3S/fWQg9Oojp/DHpnPQXsu+KKff2P1oj5qVx9c
Rx7Pve+G8UvGHvKJj/LPJupkCPpYC54tj6Th8wFDmOhchozKRjtwQ/rNivEGOKG7
GX87jb2r1Ya2hCs4PuqBt4ZnXgk6Mkv2XeoaNaDiiaurMIFwB9jmvI3S+rkzZcKO
W7EoiRtti0XRAvhVCAe0dZZm/vwxWpQPWvz+seZXRbrkc2ViGfFJeZcNBbYvTOyU
IFG1bcydw7K+cjApRRYF94YE0Mak/tJ/7jDtSVyfXyxYka0yHaAvoUFpXa7E4Djf
v9cR2doGjU3dpmenyA+DD+B0tvdChR6/WXSDDLzMYyP9Mkrb80t0aZm/LvUCVwMk
VP/oa6qyY8FemE6yVOnZiq34pWcIkg4eNWGZsRr4uSgcDvmpdvoVzbCMc/cuI20h
3PiTCBYZznLsqJ/950XTDMF4TJcnnP/Rxvvlfy8up7HvoPBzAInszNfNz9ANSLjk
jJquXwKz84fNioj9RbwJqUD4+TN1uReoqJzUarDSO49ywTO0ZZjoLzvSqMeYmUnY
uwKlQXzwxX4m/aOemeXcEFseaGPYPKqzLs9e2Jslespiajv6zhp2wJ4UbzXl95p4
Ai0nNTZRP8EPyxLYbMZgAJ6xK+2EaHyyR9dAnu0AJfXkei5amCS1DYbONyAKMKtb
6LHgA2NQCJ16zwZoXABrTUBZkbdfxgP5A3NGuo8QeHtRoqRDkA5P32vNyRj7tvnP
ntGDNa06/EFJv7ZkvYJ2MST4oA1CxkR3U+qt8tu64PhHJ8vvAEhaC/z66f0UIqTs
IKHAbGH7cc6yQI4uCd0xlBTvyofSm/e7PZJmvIo4z8MsqRMIlIKGAR0CP2sXqJKD
M/RR8N7O0Ad7mXYlhktDVufrsjhcDBLG0RqrfKDEkLBiocSPCZ0SLRpNMDu6ztj6
xNeI/4ot/0uHwC9dQecae2zYEn0fz34/eShHRLYNAK/f8nOXZwy0yvLfRyNSUr1g
3Y4WKF5aKfS6X4hvk8S4DQqoBsDLnMNwpIMDWjg1XMIEJ5eURv82CISzZn1JFE5l
ugpMN7dB7zlJmUl1BA/urwd4Hp52p39Ny6GOD89KQs3dxNm6u3t1jVxNgx8/62uR
utlEqI42SvpaXGHYhd5xmipDS2dBTCGoDlMD4LEDI4zpWZaAfFpdLkmjQL2e/nH7
XvyTlEFqJd55oHL+4OlMDZ5egi/fgmSRmfQkSRHjLs8gopM3NDFxOeMUnxSF/c0t
KEmDXVAHE0VSNGEFj+VyJylgQKcmWQKBJb4hyDEVLlV765qSECu9qv0s7H/yZER6
BgIlfO2f4DDEQ0XMaQKLIQyXOeJoXljGTTQVKkyKv8UeTuQYN//iX5ZIWcM1u072
ej8EepUdyLspZm8X7ppD/PtH+XzriM2sNbDP7BiwDTAi1KgN4wLl8wAsSp7H14cg
OI4VJ8mqUIDHLbLCNJDrV2OyhWaYctlNiGQL3IXzOf2zfMqcT9o//zZaQ3Hb2kEi
uDikoyMcdcVzjyrr15Opo0DAFKuiQbJmfziHRHY3mKqmfLKtDcJSsK24wInGJizp
rd+OAs5ReVzaQrz7WPwAA87vnJZZwf1YVqIlLzymJcRobB2wKopKGOjhS59JMe4F
7yD7FucLySnlH8OQ1i3WkFXN4/Jg60X1eGBhjjlLsWPBpJPE2beWwM2wYr35Kis5
73Egfmu0MuaXOUsI8B7B5BsGnQX5jjWZ/rsvwMgEKfQroVEVxG7fTwLPCfYHP2Qr
mVkWPVYbgToV0Tl6FJfJ2shB5CYQf33PJJfV2Gy40jJuEDOGdriz2BfJLhbMUmz6
G+ak28cNZZk8FBrFx8p8stYHcgds+taE+juypLvcnj7ceu3SYss4T/KCe8QavbF0
Ko7Ko+j8SALJO6WTK3XDHfiwa/9sqvPx9kCFkiESnMY4A3qs2SkdGslgN9SlUhBp
d6MkORshnav1HtZprHYVKKD/JGSGUspsjBR++x5+19D2MV0ALb1b90v12kvR2U4W
ooSMOG/ibZIozJGAXky5HMT2nHItL0JVMXe6291GJrA6oAwEHjT20UIXNv36FLSG
gox8kwPC9rfCLRtkYwksOdsPf4X5iT4gcspcQXs5FRmroCLBW7dnKk1m8AceUzps
9ayUcudtxk+xgNVLKj5gIw4wAeEyBdYLZzPQHHD8/rzHVN1E3jGJ/0LTEnzzeW6K
k1OHrzeVH45Dw/9vqLBY6kNoVu3nx7B8CoIVOXBtQsOii1COXLNoChil8EKQLITs
MKfUHswx9C7INY4Ql4nvHk4nMSJmZHze33KFv9rbeCLu5+K6RAVu1otDDr/8pJgb
/TA/Ejc7dDdD1RbBywzM0bHN4/Xe/KKK/9jU6eH0/cfn+Z3rMZ40MU+xo4gIk0Rw
ADMny4mx+VZoDDMkRAIMK9IlCEvOGZa3nF/4oxBIEXbmGHSwBnVPLOMgHugJlI1B
dV6BfDkzEr57Wa4oSvzrhbijiqT/Od2nm8qxGelosOs49+P0H94uXmedcDm8Zqnp
q27coy65bhPIUg5tnol4w6SaRijWt0zb4WSFP8EEjFeHSGxOe/DUOHQGV3HdVuot
4ctdRswz5Sn5oW5WQBH/eAlqlUxSTdwQhD+QfZI7a1bEH2kRzg+egyx9hq31f2/9
K+4P42fS/7GpPi8Exl/MVBC/iQcNQUj57s8Z5isUxz+4lWOF5NOBZJuitgx/6HK9
RHfBr1ulbAxiFC1aVp3dwSx4g5QrK1GylRpDCb0XiKkAsvkwvvqzu0Ftds9MZh61
zRRBCcy1iQYcSiLNVSP9x96kppK9lei2r0Q6x2TN4Bo5xd8QQ0qvoEPwta71kNVp
Pcr0hFmEcORYCInYxfQB8TQgUugVfs93+le/1n0d0FkD7IHXGaat7Q6CMrTkxMjR
hnR+BmvxGDOPQ89rOZXjHzh5Twn0WsEJatsngRXmNEG9k7LEt7yEIqy6al0y8CvP
wxxAyjyZxXVfbZYvXNfL9VKDswa7oVdSVCD8DAmE2XV38/Avbp33In2w4LE+mIVF
44dLYFI0foTdtes8ZWAWJtda/gxuWsmxGNuI6nbM7wMfmupc35b1CO8kUEzRJ1W/
9hf/wC4Xr+CwE6wea+VSrV9xdeABH8sOCQO/YC3ja9ALtd1lkxEUQP1yOwS84d1o
L4Xiu0PZqEgnjEPSnJCVvACclCDLqj2484b3/oCBb+HmmpmH8k8cAcYyKLA7K7RX
qR6m2zEaHPmB751/e8cqfXm3fhbUtr+WZrfOtHEI/HJDovN/KFm/NL8GXYJ+sSJG
nrRbNhuRVGyVhnAB1GN7joelizG7w3030TOCGZwwpNa0TJwkqngPmw693kJWqIhv
UD3Pqd3PpxQtm4l89O2ny4opdkYCYVO21ILsvPXgHRKSAX4u5fbUdgnU914J+iPE
iEymPQgqCqCgP4tl9VQhG7nKVkxJrGjxKoEjTRLYjP47WIcwr1atpHpqOoRdHLzq
zJz0zXl9NcWBgZxuXp+HV6fNnzBzkDaWDupZXFv9nGPAgrzuloC+goBjw4Xwlu1j
jxj0tFww2KqF1s0mM9p6V6Sb7vgbXW6HAyz4XcgzQHgYYlykak8oKSgkSWvsOv4r
9g2xg1e9ZSQ2a6nRNsL+KunhjlGX1KxVRsdY/leQqP5HROhh6m/Lug3G5vrvkFSW
XQRfq3SmVJ6/6ERB/yyJfZ8HMnxFz1n+cM0BeLjCWQvGo5h7pA26vEZuzo7qIGvF
mj1nzgurPrhkmttSeBPRT4RkOSw2hBYcPt/2KwvoOR9xQ7ArPNSU38a4Z8cBIf4O
qqmt/VIB/rIhOcrLB844ewn6YeSr2BJE23YeUepuqVNhmohu2XBF6LFMBZT0Bl0f
`protect END_PROTECTED
