`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LHMIsgboZuEdR1WW0yR/hAundwGS7qy0G6YiskxVfwWBOH4qwdmwvyzE6looMFq2
vXXxT6/BraVJEQ/dmPKGaPQbwNILTaUV3iOO38WgqPoDMMaX+QdvXlihYHD6LHeA
LI7Do76Lc1b2kRxonSD98IQ8dHNIrr6vQJbj14wkTt5t1c8IijEIfQdoh3akfvzK
IClmE5eRfSvl2WNtXdX6WGgCW2YS3u5cRksshqHnRUaZhUJLPMxNuIqyiHlT+yUY
1mrHRMAPeKqvOErjzN0BHVH62WeD3uzGq93iTI7Wc2nk0+jsBpiVLfl8HL+iYcXa
QNQizl6LNlmSgUqaEHFQVNFIfYBHhXFzxVGDgYqZtB7/vREPgTOg7Kcz6wOXIKha
0dZNu86wSrLgMi76WkiuAxgfstsoSvnUFfJfa08TCyT8A+7VgZSK9MzeVD2ECeT+
lECn8xxzoVW/4adPypYkmrDkOP8nX/gXh7Z5BhZxe3PbSf+9qInNUj44opwWTbKh
Zim+IveQYa3QD1FcZtzKSFgo+NwoK+XUHq73tdxzhj2R7db+tBb4269DCktx+rZ/
fljO6Y0C70uZOJXSdSHyJlIiaTIacWCzVC+j1EMIIUBOw6QWcicYnAQ5g8nrjMjR
hYA/jmlbXdBsn3TjPocAa42JRaNgThKMOyXwjQWhGIBaMUYA9BGwjBLBU9ATWpQF
ILsTWWebWayt/mb1vNH0rgaws4A6DFQo4yxBi3x3OcF8GJeV26HuzoY6QhRAhaPo
pSABk3Br1FsRy/KXIaV3Zg86QHn5AQfyLX1hXhntYBoal7TNzMxXwz7Wti+ZVD/c
dE3ySiCoGyiKvpm2y4DdjxHjOu68RpGHhJCHEydNLg/wqbrIKadc1EmlEv8cq02I
/TaY976SKxor6PC/M9UXWcCLichJKS4ZXU0BFTlLW5CoVU7jGmAUIBLV2YiQfO5e
TnpU9EtLJlMHufNJMAVMnhlNtmrcyErwyCLIXQxAsgVOfHk7B1y6CoGfRT//YP/c
zro7JJ1WWmkVaoNdNRfS8Hpm9+kFrHQfK0wOytBsUPhFCleYpcBRgC37LuxiSzrb
3bkzPb8RGB3h0eYpg9TSYdVWj+UyOkX60/pVYlfusZQ4IKQ0IGXJpUt4BgTTcSlk
pbF9/8cfrcj0PEUVtGKMOpJOAHJxnCT70tl/yVoGPwsrUEoXkmFt5PwJfXXQgpvU
4Q7R/2dRLhnuBfkmq/1zrWn8RxboHA7Zbi/sI9I4CDo0v4Rfu0AEZuHEGbwjMhrY
hhvHObnMdy3VJdHUTiNxdLEJTw1ibt6svDfej6qiCLoBOjvz1zY3bl2wHZYnebjH
9w+NJbkVcPkIY/2Xs3bmJ7d1riYEfmEVk+eNZRzX3DcOo8wdMbhZ0xLLmw5AYSQ1
g8MQZM0J7LBnlv6apd8hbvQVG/t48Sr5adV5noDHxsVZHwdH+3DMkcrHYdti1PLy
h1JJ+dtm7wuIxDAziS18IVMtAzw/7/1OrwnoFtsMNHFuuqWUV2hEsBuIZmNt5zQq
wmSf834C+alSQISDEzN+prhHshjX/wm93dB++tN1B4aGEaMWSgNDm7Cm5MeQvCLy
12Vrj4olijUGswHaEty0ngymRucHUe5smpTnxHjYuprKqygSLInA+U69POW4ME+O
efY/qD6syC9puirhbcxNDs2QBI1sbyXeMP+0l1JpywCcHOVGR/rCDNW2j9PYpsxR
Al/0gRh8bcQ+YPCcTugsnKXm5IWRWPeg7+IOQJyP0hu+YeU17hiFQatFvbvITf0u
eeYNXXPLNPNra1faT1bee7P6gXmK66o3fcdGmqMVG6wJGkd1tAk6em5uf9+YZUpx
IzUbA2XDu6Rb7xGacAjctow9Miwdfe+T9E1UkaX0IAOQAxPlvU3YaVHDCjqwym+F
E4BhhN0M6JGs20lRbn15sDFUxNlL+h+m3wh8m3h3KC8ivGYVeTNkA/34IrT8wDH3
PaV5B3Vh0hDjFZQpExUOtK4jS3NsMvENgYcaAMg06zYbUMsHiZBZJLoLdbBeTRIp
o0cquFlmxfxv+DP8kY7XxIHMOMUfCubukGfVvI4tGDaWM3T2bbaYcWM1whBMJREA
bKBiOh7VEtNeHcGaRzBUmdJNL0H8PULo3Gk7yBqkQLDttSxGAxI401e1BExFPsmS
DX+5aZWulQHcm7xDuFf3Rxm3VDJk9zgP/2/fbXgizPV90jinsEoM4b9wMwBWhDPq
NDtVcys1BFVq4XynMKXZp4vbGVk1LoylCAbcZkmWegSC7CxJvx7kD+Elr/wMx6cT
tzO0vcVMxfwVyzVdbHLaGdKx2SOorIGIKKa+aIaUXoT1SO8oUCWTxgZ9rtMXWBqS
5+btPdLJSCFjwA2WzkufLeYl1yAaQAHRt2HkekTvyPiJjrha8M4IRbI70+v1oYM7
b8X+fdWUcVGiOyWjxGjCIQO9hKvIB8kpbcv/jdxxpckrNxuTOGUwrtF5Fn5Zmk9h
U+CQW1Pojv0OVCPVYLYQ0VOSvSr4kW3SzfMiyNLD+0N4SZJYpM3qNv7WSijfXYR9
DnT2mqjxyJLc3jOTLn7G7ovRZrc2Sm/Mu613zYrJgAiIFxVRqmd5DysB9Rhcol+f
woMFFf9NRLnnZ6Dk1mkW4uZFqHOa8e0qGCB9dHS8PhViW9zhEl+rXGjDBlPSGssb
r/TRM4kHPI9hR8IzAtzpGVQzvWroe1skJzR0r0M0GahAm/vHYxZD/RN/mWtDgjUq
8PlcfH1LXRwJUu25fUtF301nllFXItz1mcjKV4H6mJbw0hi/XUhM4dmHzMXbEUT3
yIRl0JeZClqDT7lNQEAPkta11di+OsiSO9MYYMvgdM3ubYXJjDRaBN6GuX8vN5n2
0uDCVUPhc6afcWhjjlddgbOWFP3othERHcDlth9utU8t9doBjWUv7JzXdylC4qnE
H4dmyP3iKtmJwLzTHv54LfuwtDTl4z4kSX+ArU/6unsUOoA8K1wuJ62EKrVZHG4h
7SwNbMmmX+cyLmGFhOSTEsg2QTr+VnCLLe8DT0l2fhk2hz4do1m0of+Lix/VEMER
veFpxZ5VLI9bH+Q+gsAP9KKaa7htRPjOU6DJW7WZD+ll03HPQReLZ+6UIfOWsWDb
vCDhmgB045a2Mojme55FVNbZAXIHkTXBXvOKf6VeT/E=
`protect END_PROTECTED
