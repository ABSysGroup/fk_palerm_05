`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tmhJndlYNJS4uP6udyJ/06wvINCcHUmGzLyM314X+ti5k3aHLWI7sd4ZlYlkwrHl
2koZxuxqc8MRfTwr4mwdd2Rc4McVEzOaH5uH64shdTAI7AzKbhWLJ2ICMb7NhseY
U90cMQVtZNWgHuZb0m8ljKL/qosCMLJVrX/81nUTPQPQAEKgH41eXG2S5RFVB6n5
fniT8xBj3EQl0aI16OEL7X+cEfCPoSGibBGX9Bsgqv7mQInMB38j3yfhDdsklhZg
H5l/E8SQ5rlSHj2GTY7QCO0eTwu13UbEma6NFsJIOqCcN2EMb0kzwqGPFqO2RDRr
+dKjQOzcWg0XG3yf2dze1Ml65rCfJD48Gf1oBik4ZREfPk2cDrf+IwbBldkMe72G
`protect END_PROTECTED
