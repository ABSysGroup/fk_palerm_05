`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dvLh9flhGWSKyqjapDiBJyh9tQA7J7iVtU2lL5xn+tC6zS79Rl6NU9OZjue2B+Wk
dCwnVu/uqSV5YAM/AkRGTYT6CxJaHh/GXNnUJOAVqsBkaGwf4/ydcHvFLYre92+t
DJl22g9uSjFYUyv+JUbaYHRA9tRzCSyju/fIXX3LGJ0ywDtL0lCjV4uECHbaF6To
ymN7DhmTdNMqnBM31v29Pfd68VafFM8l8GRUAo/1M66XMaU4MIC8R8+0CCtsx6pO
KjcO3WyHYFF6VQHFfxkPz7CvXukiyZ+/0cbuaHa5gDvs1C0HOTllHom2JtDIpkj/
wtz5XkMa8XS5UQ0ZV5gnVmrE9eFS/kIGswWuaiwtINP5bZAYzr9QVHitxoRq4G++
If6tY3PfE/kxYQKcCrSJ1wZWng6vwASXI9t1lHsmGtk87SoEFmgIzB9bAt5l3cAv
VmEFgC2KURUSABzjYGcbj2rLZOiZtFVsnuCniVlgnWgI3Y89lLkGIpt1U81gY45X
`protect END_PROTECTED
