`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QM+aizqsvtmLxXgiGch3HaWv1kcgzoDEQZvdEs8anMHxoUa3+TOCKbQaFS1NI5Ff
0noM8fsy2IcsPvZNMgz0HOW5gw57i7lxHVwgUPqR+jDoaH/D+z0AEbD1zsKv/EMn
41lqYsfO++psN95P+l8k7KOQ0wg4rdhhRqM3qlAohnHIy/h1uW1s18XXsYS+77hM
NphJY9kjc6TN3BV35DSlPemTKzP/lL7rqVhLzOdhmCds31J00FY0VMD0kGJK30go
rBRrM8nhHJ0GRuXkw3/Adx6fMOl075NnEU944Ntt9mFq+fFZVNujbazdHEzhD79w
nyTBZfRp4OeuHanvis8FfLlVOjaok0ZNx65de6NQ3GZ75RPmGmJSFTjfxRkYXYON
Is244trLXEoYX+V7BpRIi1nHybeFOAUIoS25zr4Iy4nFKtzK/rGuw21WK0DFY955
DPijj3+VEmhzmhufAsYrB8OL50PEudwLWOECipi3iXhpsdXbwGs+iSeY42nB0qdd
6+k7VVREy/yf/Yah9jRNu8usJVEdX4TsVL5fgCq5u7XDwwIcWOacBo7q5asyZWwz
nQZAWnnjwxrPv03JbKBng3ZjkRi02sAgMBthbAcxSiTH3IkRGrIn9/GwOl4MZ0qD
0AMBtrcrzQ+VhIE6ThMwdJpt+bQVpZQ8nlz7c81MCNx05gj1ZmRRmuh5kMAXP1Rx
kFXRrAqxkkCE2y5fG0xI1wHaiEEKj0jvn4v9MmF1se0tPxSazqLFRPH5zG5Q8pK+
SDEWt9qOTcL6EsXhrUnMdePb5mgRQ5SrUHqjdpK4SYOYbGp66ueCNrwsyOxHaYeE
h8CldMFcm+tcobo+ASHAu8rLlXWznsl1h7ezK8OPB52+oV3RGzW7ttPd6EsfzGZM
IfodgSJbfuY3jn5J9dBUvE3qo5MbfzkOs/Q6Dsu4UZPD2U7gvbQc8ahM4EYm/piT
+/NjfBmuer9c1phc7Nh53tezfW4JzmpNz1rtZ0f+/A90SsXJuBB3f9Y+bORamgTZ
tgfQB1+ouRCUMwQUNkkgMZ6Lmm4u2CGNT8s4hYHOt0MMwNFFtMR3iFuISrtEhZnX
GYgXOY6vF+xx/18NeJ19sGkuRNo/YuiInC4VE5BSx3VVoATpajhc901cIQgIibnJ
BNL55o+joYefT+Uolbn/ry51IAObICbqdtMxRnwZ9M2OhaU+Q+/wnLt0Dcwt8Qcg
+lc+RbUYRFZnXplxzh34XyI7BNwq9f4UtDopp297mDqfU5eRtHc+ntK++7GZoA0t
psBMVNmCsTuAnIbCIrjiP/1278GG2ar4rHTrb8t6MFR+YZnPOtW0zF4x0JyC3E0J
`protect END_PROTECTED
