`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wMMETRfwPQN8BvYmq2pk4W9YciO/JuB5BlDQv6soPKME9ix+Cbca9kJ5tiQQmYWP
6pkYh/SubzK0334JSTTHYwIXYY+mfC2+/hmFQ80e37FlVfb11MOkrXOPHBreQddQ
ZemD7om/47uECtDdgcEswR4BCQ0dYgOW6GUh78w4Wn255p2B7aWtQTQ+l6DhhS0s
GbZ1HCNm/xN7AePw4OSFUsTigrhw5nbu2GRshR4/bNsT7wCvcF9EGBJyRiwdGize
zMNrJLJNqZ9cZEc3T1ZmJA==
`protect END_PROTECTED
