`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gnAmlDyorrvFXMRa2fnAj+uB/UNTTyfWG6GbYiFyonOMAQCGyURyClrbqzxsUgPo
l5L25zPIc+B5+3Cr8427Tj/8n5jviJ1VuynOdZCalStYp2NeGIPnvEDNZjYpx+Ut
OQn0XWg67LTwEVgBe5Rhk87a8yuu7q0jku5BZLLgLJ7N1tbqJGhxUo26zuALsiEs
GqHAtlWf79vj3vRxNslMkzLKBDbDbEtiGoCMLDKY4/ePS2eWN7dpSmutzOUbFjKs
P2moKRyC3h59xkPHrotDg+Lt6YFn4mtPZ3ALjb+qNIHZVvQJNf7R1mEddKLGvcfV
fH3b7+j5UPbOOvTA3qvUUYGuLY2n86OVQXgrKPDvTLrPUZVEbxFzrPbZ8N923kVy
V7V6IPamQCnUiimF4FcSiNVlXeMZx2LG7dU6+lz+lORhgBXIK7VFLPGjjau6fqxZ
vRPwfSgBvGHNefbzXXwOVVgKxBkXY9CeL7TMv2X5GK7zADefRbui+DWpER6UFhWl
ld5A4Ja3pcQy+ezmU/O1w3pvn4f0cmGFvxYcLqp+DuI7o1fxLbZbh8n1A76BkEWV
RlmyQrUAjgMXy0oe/zKH7kTHVT3xJzVC3jfcAR52nF6uNTQhY+52pksBnBwtgXqN
IAPJf1M2yitMPO59bDpRwixIHjvrrrccb1g2gPU49NI80HZ53uMNRGeV1V7MuwoT
ZWTB9SfNCU0WdvlftnrEmw==
`protect END_PROTECTED
