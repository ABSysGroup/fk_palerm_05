`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GRi1DbbABENPAPA3WaDBF2YWHoHc5bVUOaVwoR+MHk2+/mdfWSBoOVw+Aqvb3TJQ
1+s4CmboXKszvIzB5RjvNWXCG1SGcj5yyLHq3qCV+IfetqOfLNRLLJmrYJKZqOX9
J7cCoVe/gu/dN0yDtoH4mnf1ZxCk+EGLI7eiXNl1D78/prgzREZxavD5/6FCanbp
a0T4/4XgJogAlZda4DmDC/Y5slvIYAC/Wl2gQ5+A+AU2qNaC+Drgcf9sVCcdmfTD
iUPfThRWG0Zlo2TGC2ZoecGUipA6Wv8JQQFqBhRUcRaDrxmAdy5+EdbEPW1Yf1Z7
8lwveRrjll704KGp87NR5UbK3BWmQAF2tpdCCEKoMw/7i3dbyOLzPaaD7ylucToV
SLfq/9zum7TiB/Jxhdw4Gl3QaTuqpe9ctib8106vHCOu0riiMYssf55l0ZONYTqP
bkJAdNt6uQogsNeKgRyel29BdoieRAoFoAstisCS6P9U+IX3lfvLZKlg3CnfMk+K
jc1vXgj/qsPT0Mz7uz74vIye51vDrY2yyKk7rQOypXnFfhIufPK4RXDNRoQ9wPeR
8Cxfi3wLgCRtMomM6B47yJj8Bm3Rk0Jg9WlnNKjiN5eYCKp00FylzWp92A0ltXPr
iEe8TGxaDxm85KQA5hGaCbVhY+QLoVLJsJiHw9itYb4kRg+iWdjspXEQCSJ1bH7l
7uPw9O4IStNMbaLaGwsyZ+4FN9bKbHgK6KkaeZ7Q7bU2dgHaTyToxwSF6kS6pzDi
8y50mi7HHNziskF3d4xKiv29A+lloLiKMG7N38c7uuTL1b9pobCLgxAeCcviWxm2
wfH04uQ9y6G6khL0GPdciwsZpJnCZuL8TmEwRadZ587r6lIqpmcvcK9XlqTIthet
wArrZTy0GjnyJt4nhQiudruBC2fxCN7pgmxVs7Y93ztXhEtDxgvZ/c6L6GRThNs8
nLt49kzZ/njYgu1Jp5udyd/dL+LiqnTQTU5euiMBemE+x/tsOPEYO11K6NwUZXZd
QeBRGIheQtCipWpu4YRLPUfAaeSM9SJcH0B/GIf/1zD5Ic9mA1CgknM7H/+zOtPv
ZzxMviAPJBdKjKkExVQGwb4W4h90LPgXcHs9oFuIKGTyBZRIiT9pIXZ997iF+Tog
V3JnT9y2F3tpl7/bCGwy89oDLmKIjQt0hrncImeRM0AqL++yPAoRsyHvYXbuXApO
psNI/IRFx+8e09fCnsX9i9AuCSgbuOBngDt7KQStf+URI4stgFSlRhVPm1XIsh3C
EQ+L6EVo19Lkry4OrJHqRSXkGShRxQWnCnZ566KrPBclhbXESLZTLsTBDDjPFjVx
LPEmH3QQnxVxvqpUhodGbNXxLPVV5JcV/TJNRDrTHxblCBngJ27cZxkPqVp/XUQP
DQAS3umoOZq6S11Et5FazIC1/G9FKlpywlydThwyOFvJwdnvkC6jmc+Ap/DuBANs
juspzYar0SJFK66YS501or8sPPt6t86W9c2Lpx9JqDlTZhbSdU8ID9SpLZALxBSq
KPG2KZ6spz41K7Zh+kfUicqiPqjwXSeDA7mFhTKqjDMvrSf+iCatoQf/Cb6fCkBB
1rpIMw2eLrA+rB6l+extUI1HkfrBSdaH9hJTpoIMgdyphFt/Ikx1sI0aNxk4BtFP
jSLTdjqwRMNh4++JEpyhzfQOlg+IbgvbJbFuCsNK6+FvxcUGW5Gdvl1SkIuYouV7
vNKJhMhvdpYIATM23mpJP/edSazYTRJVGP6gSDm3dyq/g1wS03ReB0SCthyGi77/
hL1lPe9iUfdUEog75hzMEoI/6B3VsdL+yDtDJdOEwRzoFIh3hJmsvc0+wZaa7ETW
bT6od+TuXT0CB1iz9V8YIcfk59+hc0TCSQUzMBehR8vPL4sM5Lx2VSqEXdMQiyPO
9wfpMPNkoE7LCE+qzspaZFXygkUExNzk+BitD5YQDVS5zv6YqtukCQvEveilMGsA
+57CzPWDpa8C2FQCCj5beE5LgQv08wJit28cvL0a9xsQHp7M4XThq8Q8dlwMA+tw
zdsFR7MkQKHf1GfrCAGnF9wCbjWoGUKYapheGP3gxTz1ksOro/HnjAi9gTafi4T7
jHnwKEZwh0+codhX0TlnB/pXaSBWGoFHCaWJr2OatO6AlU9slo7mByqKtZDbnLKR
Cf9G0ph90SlfLHauBYu3XZEBwTELfzp2Uem6hDm0uX6nb6EPDBBPpNdUTZ/JPZCo
Ioud3rg1Hlo6YqKBmaHUBwZsNtvZ2j0K7O8AZjf4+S3NbET1molzW6f3gEF/E4bL
BwOIi/CPMAC9mkg+R+ThTRGS8/k6GSsuQTEoPk/JACQtaDcedBaPn9Ql7DWBqjl2
x9REQUCPzIE754kpkW66lCcCfpuWLa/0UvHrEq/EUPYgjSYmesi+HlzPm1wRoW5j
uriaV10fC0ledR0qBfWNnSdgk38Z6XtpFKDfm7Igp8dtanXVI0M9gMUaC/v82A9V
HsEr5AeEVSCXhWmmECvnuKe/QnoBRl1596qI4auVoOJZsqr/x47HAoQRdWN8qLgm
iEY9jU2ENqO/42gczEa8O2UAyhWbO91PvRgWla/8N+hyBedEPNHYLUR5EABOgziB
urSmnj25plmIn1xCOyx6umYods03jqDVSKaYT/9RNt1lXa6VBwEW4B7wWyVBPkM0
e3mNi5XN7j+iVuJmNG3NgERImaZCbyXN0hJQyxKG6PFZKRysuQFHTbgbcGf3UYAY
+B0LKU5XvqAyesISZf3DhlmDhtOzGwqUsuP4z4JEiP5Hj61AIrBB0xv4zFwb2naJ
nZKxTEm9hv5jddIuaeIdlezZbl6B1mxMxcvd+jRgOUutF1lAWDma9xdzPgchEZVO
0oV/2BkJ7vvWvS9v7lUmSBabLADRX/QPHzVvxge53gB/4j9yaUROpDo2ESEE00Ws
PDFhwKFlSW0yQmQXibT45pO6/a1qisHxVs/w++kGlrLKr0KkjAgbITSY/WBPSwRs
1T8050BVah1oZg4J5qFPu+UKjUKws3IVopFYZnzhhcsew0nRtH6hOjoNYJVOTHIJ
KNuhB+Vl12xaHACPoxto9BujVYEuwpjyAMn9R9olRkOZ1esTfa6qga/xnoDrYSb9
xxlakk0xQiuYb+yiad8SCZN7t1VOn7RnVSqN9o8wGz9tCeyOthMHg5MHDCbCIzJe
H1h7nDM6p3ft2G7YkqmSzbS3e22qpjPk97ePu11puADRVcTvrr1gSlK8lUnO3sZu
8X+MoTPTpM3ZHWr7Zg0AYKLtH0iuuUInNPsJakr3Kzeo2hTMPKaP2dzDzwybfgUj
/9LiZ0wUEFBfN80VwkYIuXvw3Gid/gl9rNbikIu+/hQ00AwhlWGXdU23kmma+b2Y
pncqH9yQO+vPcUg8m+e44RNYOqPO3b1JO5IEa2nkddNkzjNy2Grgz5sJjiym1Tfg
OcG6IJHNyrQPaJGYBJ543rXeF+0ex8zO0uG/HS+OHLtVU8y6HvWedygx8cKI9gQC
Dy+cys1pG8jWHN4cAVa1g297E7AedZdf3+XvsViIkj25yfTsCM/PaJvWDJLxxuRk
vs/19Tn1YKioPkEz5LXx6tg5KOAz2HPEXqyF6KNch+XwfswUpt69VRFtufl0dMpJ
eewj1+XI3KaANFMglt7Zq592uCsYBvxB6kOXt6wKpipqN2fJNrEeh6aqT/musPAE
/d8ztsvQLV9IEObW/d7fG9kA2Ai4Y00I7smm2Jnc2PTmPgI+PgvDy2xgKY8qf/MB
Wg7gV2gwSMtkHDp6zJgtzR/ZxQX9xI/lhvR6i3LXvqyr2yh3hZ/iuJh2VdwDID6X
ndRqtQyuoshSPpfdGuexLxXhdo0008eeCIX+0P98cMOCBTYfBUZ3mdUZBiIIvjR8
uUX85XFNwEq39YS+3BqGx10NEyymJ8JRGToRA4wK1TXFqLPJDymPP/sijt2YpJkl
qs0cfN0cjHyDOlwOmgDFDkr7qIHLyUSdHv2KNBPZPwWg+QtnfYSh+sQCO7FGgYPj
vIfTPvjuv2IJn+0Eh6Wf+xgoQ4rvPna1A15PdHX57Aoc6y+w6mFIsx9qB9+AUDTy
/EQlx+Zi76VWtiTasTmYerQWVyVug9/GOXeyE2i4Ilex/UAYSB1TrozOmIgUypWD
EYvvc3YPtR5J6Jl27UGryRe3eX57yZcH/Q+eeXRIac4U2PelYgbY96gA/B9FpQeN
BrHU2u5EnaNu2Rcv4WfKvIzAuuGOYq2CauDUn35Y/rSlmuHg0hbCdP2Du6JiAb2d
ibF4ov90za3gusvszohaKMAjDVzxceKMcO7BCZwV0oHLHXqh+Oh8tbmywgokxYXZ
mg0fYt4QMwivG/sWvsO+/kEJ6XUkeqhsiQ9yzjmcBxdWTzbqC59l7SxngCyCQGv+
J2MCn8JCJsMYcdy2qCnn8SNOAZRg1BeoWzOpa0OHpmjGeZua2kZQNVtHKt8IGUAM
cOy/Xrm6ckuaxgh7zMlr5hHqmtY9AbLvMd8bdlNQg4eCfgpdvuyiCBZLl5yJwmiu
/0mPky+4M8NCOQZ//4U+JFdA6nD6C/vq/XzG9Pgl3t7iiv2Fjt7RilbZBo137Q6x
5Oj5gtBwKoTD+l3GnIyQGdUwqq0+gaDZ4JwjBRIDFdGn2AjYzwut/Xuwsi+kRtM4
fw6RWNr+JLoeVPxR7RWtG/X0dBfvVvGjjlHWrqPRG2dF2lBwrvOyM+eoAiGGSVYr
b/GRcHbi8fm4jn1e6TSGlNa/MiqvQi57AB8bhN6aPN8ZrJbthQ105qVIonDRnXOy
VBiWdhfstFsPA64DtQP3l8MRLI6l0pd8ML474pjfJlBeKTgCDhCHWoYMeXaluijR
F14n++Gv23bEg8tNSGesAotHXh/F7OHgawf83/28CNYadwp8SLXP0ADxwOTzMnkn
ZOAUN4XII0x5yJESBvtQxRizrHBEcdiAZ+qthKJWdwxux6mINxQyK4CshHSmIlGM
2JQgb3iV565DYBW83d6IRZzpdAxRnfMf1Dwwp4W/z0Dagl7XCzVNC3ccd9jSS/G/
LT/a9iARpZdgPEs2jRKlrZ6dnDPx2U2aLyboW2lx1uQGQHgzyMrgb1v+JURAH5TN
PF1DEG05rCUKdmX6cqjPqSqN3S30BqTeVO7lRrwdncWz6e7+bg33tRqYIB5+L4n4
xcRuoMGXYK7a5ZtvoGXXpOXcYOMG0aPhrcGx0npzjVqrUnQ1shg7tjr5WSttlUDk
zqMoflMJkfXqty3oSYypY/27fFNdptw0iBphtqQJj0AFozrsqOGDlU1gRwl+jAAN
BDUHo4l/6bhb/o696SfwUR89PLlpMMGwv8s5059NqOv/ZS2g1nmSpxsod7yCnLvY
JN/bx0aH2JszEd6t58BTTl584ON+y4kzPqylV2jbLvVBqSQzK0Fe4CgoVya1iv+b
kSICEHV2PPaGWJIrHs1IrpYN1FwPwxXcsCsu9sT/aBFaP2hblf7KJwYRSoQvIojB
GmqsXKHXQGVtV6YK/F0kqFkbtKi3p/iVsdvuQKzT3ejYZYjFCC0WxBWmJ7XJG6Vn
VIKQeGq7+OcMcCq/DDOP00Z8HtaqWF7IzpnysPvBs9A+BiKW0icXhyRESyLBHsNN
3kFNEmtCynziXgnB6LIry/AMAtWp9oSTAXhSCOQAL3d895YqYtFEONzdpyo1nAEa
8TQPfAbpDMdlcNym+sXuTjeZ5su45I72dj3zhXdk60tMvv/QLzrsnFJxa2N8SMpZ
JdR/ZT5Tcw9vTAnEQB11ObGoSq+WmLtzFH/z55ErIDtpJBYih01oJDq6/AUxP9aA
xMYQF6p0iFuoS/2nvaGvulL9NE2woojZMNWvmBVJrt4nx0glGBiPWBBsI5u+BqXQ
bo0/i/pX7uZEttuz7QR59TUAcWbEXImXFPjiui4YqYWJv97kANbROJcEK0Dv1+1d
RvbHsd151nWK3jXr/8h5cCe7Mu59OaaIIUiD0pch65IVsCVJHyuITRAuLjLRkTTb
eYwmTXR+91AgCyIQayyoXdU9VeLoByu/64Ey9+rPgV6iBsVuZJ4HsBdmgERYxrm5
PurTGSBJaGIazHWOMnCEOFCjVpfyhDQweGmmwc+9k13MfejladrLuZ5JKt9hOYQ5
TdC87i9/ksBrQ/Mf0BHfoz3Gh5+2Xje8K1pf+tmawoYfEUBdKZKK44ag0aQr9bm0
5xPyOr/PN8p/OC1ttSDLPXCbH+nM7LjGCdMhJWOoTCQS2dF/UMLRUVrsTl6iRFg9
tK9sjPxlQbUFDHwMjeaaUbdxWzEcpis7GzkXuBDQh2laEo7WlrBmzcRgNywOg9/S
NRqL89uZbL5Hx9sas+gsBjTMUR+i58b9hdKNm5Ry000pjhB7h37SCvwcpbjUdtmd
AkXCCWPpt53iqs3umkO5CejCfO+SicbHksOSTUOgU+BDjXiRPA91aNHGnXpNADXh
ylNzKiQmL0lq6ATxyhVeQQsjafvUGTv63j0D5Z0vBzxelIeDGK4tVRFgITK15jTB
NnxxdjYNjjA7IxiuljO5P89GjEk5IBU1sFZYJZy2RoSNZEMdN1jkbuXxb5CdBWMu
xCJc2ID9/cAY+/ZLrOV7moDqkmhZ0JWRMP/1XvWYWRAMKEwrAOaj6OP0p0Ac/gr+
hylLLAT+LQQqk4FXQeGs/gA4q0xJfbmtqMbWKbYs6fMr4y+25ehv1EaH1685lBWR
57mypFndyU5Fusd0Rju5+ieJSueS7nJSnPPfg4bkrfp/VHXR4t+6hhdkLrOqEy+7
QLiZ/3C+6rG58FRB5K/TUszDouWJoc2AY3sGRjeJD4HbP5Og+jTBF69Zg6LQwBr+
+tlnnqeLQhPOvOYi6GmhtSm5B8lWgrFAfowqvoLK2y4D3wt8v4On/+ekfdx+6zeZ
8jXbyCDU2au7pY3tBj+o2Psk85aAg2CVvRF8Fj9NmKOzuuXaYE4i69038frynxcP
77rt33xF3oQaDXFRdkkxpAmxnAQzG1K90WD+0VnuMNNHzzEqOJ6dqjLCz6QVtzWm
InImmdS7Qwz2fyZmHIP6UAdU3XFh9LKc+fmb2NQpxieCXdofsHxAzz1b7q02OYSm
VG7qSx9N0JsA8Iq1PPztZgYbIcqr2oOd8Py7YpNP5q3RK/+iyEKe45Z8Qf10/LVp
17vf/fTNsUdNnDDyvtkpTfjjpO1jVxWAKKm1nTp/BwWce7sFXhqWKn2ebdIbueg0
nFvIJ4rqf5t+9+IlDqOdaz9tbsokazkUnPqYLis6q3zwrMywZ0LYk9q+tzlXAF1f
w7Z9lTWSGcg7izHDkIGLgfl+PkCp5PHKJWGc5lcYGYVQRLnfdDpkiHHfXAU7Rax8
+gyzglafCfws1sM2aoQQti9EaDMi2StnpWha8t06HCk9forWgsbw120DO0IHWFRW
JlTN6bK5znXXbzyIByCves+eSv3dcRf1pqL3OUbP/+jn58EYRKi5nflU8Fxn9+Dg
JDS+6qMXcIzU3l3rEg8JTCnAYSvmBOxNEmyzcXFewbAGM8x6opFByLxjdL/4JIaf
KtCy4/OeNbCxUQCFH9j0F1A0w7iT9KDzMIlRkHbG5+pF8fHY0bWJ1gsxnbOTSraW
WjVfviJP18QI9jpEn58NgZVRROaQ2jGBeLvHHBdZbDXxsvM8PhSDRVTohrLtakpt
j/eaKGfyY1gj6BWHlO56Tw105uIPSy0f7E+abbAc3eoGfqLuPmjnXqnUabHLgMeI
BqebGGAi2uU0jd+tFl3ED02XIXXFtnsewtGdbqJGAyNcSVQefKgQX23Y2h60oo7x
5E5cvkB+JIXDigK+/KJRTtKbWiALkNOkg75I1PmneRURv8geHpzF/mjjcbWzils6
ySvqLNj+AED3WIAwvoInm6tWttoAvdh9d6ZCfUSzpLVUtFupjjscskn3w8syoZUm
k6D5fMuPOq7Ugqfe/cEBilh+xkbVYRp6FNxU+/rn0G5tW270izZRqprEQ3/gbd8c
dRGw8NqHWzW7Y/ekF1EZBiofZUWBvNT3eFVPA32QJdcfzhBvZB1Pih9rTJ/I9JMw
1sdlW946WJdM8tZNNweVJB9TzufWVcwmsmX8Jkx95rAUVEvU4agKYbulpeFFHQI0
ChjJjZEap4rddUgkMpVHJDzQ3/DlJVMcrpJxxnQ1vDz1IfZ2/Rzo9WZqy3Pz9+en
WBxUcwDEr+VG81bRunkaR51KzutekPXzG8swM9RkFq4pwg4Dn6KLD2rG8D7+0RWt
Il01MjRax3Fhz+cmhAOnP6fQupT07LTxtgyOqvCxejKBYRK9oJG4OOrcdDCfOvJQ
z+RKAFWGmjMNHV6xVFH2FJtxus3MapD447/KupJUs5OQU4B1OzOOhf2TG33PkgP7
+sLM3sIrEv9f/YUtlOZFZ0EQZtQpwQDEaCVVHYj/54akWdICUfUHublLt2CqsNwm
ZhDAbCOqNesR0LXFoBdcc1s7fhgk4nn6YIPr2eNAzJgGTtulo7LI1vqeMD3Af8QW
Y4RUEWzJSCEKYGJCPF8o/Wo6Mvk8jpnAeqLAnox35riMuY/5BLyalQMrckOwGwRm
+gurIlSkBqBJsciOLfkg3Aw0hGt7f6xaAU88vcYq7FdKzAW96lb61rJSVXw1+PGp
bDpbwR+YcUw2PZwy9qGhRLeumiEd6I2mkWt15eRQX9czroEOQ8e/omGrfdgh9iIW
AdgKl//st1CRB0w7K5GFKSegNckLNP2hU1Y+SMeLKCwagDDjkcMN2XVyI5JcK8D5
uqBbKqwa5lY/70cvgKyCQClPiaOYhd2ZVXsiz5UX5H6LLgJx9ft/fgOXLsXPDhv7
D6K1+RGXOY3DfkeAiYI2pMKYKp7hhPYIlT7TviCW1P6pqA7zjUBFgOIwom6aCiXF
s1QpSOrvcACdx/6idLL1XzXpQ3Lg3UZdh4/XlqZniisdKtz/FQOPaRW6DfhG/jah
fyb6PZBGP4y48LpzcA6vTJl+ZOMruZQQLMnd9cogZjlNppoeW2khm7IJjC88+xi7
ME3gito5jAdQrySz1a0ujgN9aSPMlL4+oKMN/Vcz5n6moOUrieF8/81LJcfVTLDV
4ZCz1km+WIrxjH8znD019qqk5PNfiVyC/4rQkm2qnW45jD87ED6w5l7yi6b610bc
MClJ0c3X/j86UAZcsjriYbMHiqmt0z2I53sv2YHBu/dZp1QObh0UvzK/7+cJ9amN
UWFlYonZIdwewAAyocWBYWhDZDcikijwKwNoqdehAFAbCglI6nbJpL01beYnkSyF
+LI69t8xbUAnmEz2t885xOx31gGYO8cUt2UUTeidXccjDwy/GK0ufX4+/i5QbbJg
PhWm5wgQiPjfPQ+fEFdvcIg78Enu5olrjtWZ6JLdEMrpJG+tS/KENff1MixhP4WD
4QBRmhaCZS3GVwY3BoVQ6nvAhDRKoQIzkC/yINOaH49qI5u0OUFJu4Tm3GCV+5cG
1XNgzWN4nCRpmsrs7dtmuynvcbumM425Hf6UlfvS8gQgnvWIVLqc6MEQeIidNLRU
o2+DVC4MNOhdqIows3C1Vw5p0IOtABee+oMmzb0utz0ZBJTm0mZektyNIy4kaeni
Jvr9i8OUBVDBI+pdxQRXdMlcduJKh8rpfUjPBGuK6TcLgRKbVy/Gi+n+sUK1VMq0
hVd95BUKdxP8sxIAzRSAwV1pkWMhE00ONwMnKazN8YmT7shS4FK5S9HlgYeyvQne
iMGXhFH6etVclxYXWEJNBpzFQQIk3rOPv7S/7sNcWqzwA2AGzZklJ0yG3h8Zo2HX
VCsWE3Ah0ooMIUYocEAhCeMgeCByx/631eL8IDDhd7uRsmJXg+Wa9xq6aqHRpZtO
pOpS6MxxCCRmALnkOxfGRuQ9PUnv4zawH43n4yMuhw/tXIESsdo+LDlm+I0WFpeU
pGicmtAIbJYP7YmmiQgKwg==
`protect END_PROTECTED
