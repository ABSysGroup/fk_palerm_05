`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4gpAz8RID0ZrIO4MLQ407UUVknVb0lXQLik5w3tyJ59SZzrKODlYtW3enesYE2T7
eChSzVvEuPtB6nZxmY5La1Kh6ig3jq0imxnhNfLfZOqy/ChW64T+BczO+EjFymy6
rf+UBsb59Pr782e0Rpo6MUZgwDUordY1V0qi0/QI3ronLbukp+vrz/b5NpAOAKA2
6VlmpaXRISXzXpPsoFpq3IhlrA/gOpJxJQMlGbLhaMx1+Y2MHcKmM00f+9MFcw5f
4pQz/kOgO8vvdcRLilPIrHJne8mgQbDkPIupcysdwA0VYSowPe3YroeS5d3K9R7p
UpGI1QgEbQZuG6jzLMp7nZ0y/6obykig8lP0Drcx+DPNKNkeFlpixERwtX0q6jxw
FnFuDPC0fHBZBocArXtACV/4BHHjAIJ4Fl6M7LroqHx0VElMi67el44LmRoWtF/l
WOhw7LQqdefCKo2kIM0Vyvn/DalGY1dUGjo7QZot2tU=
`protect END_PROTECTED
