`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6NluiqztiYfRg5fMK/aIlTti4P2g12xMKbsBYBFav3Ij7f6E2u5OG5dvymrjDd9H
2+Cbz4mVFaHdJEsxLbAK/QerjAI9YxgHQKOqBNp5baG1RlfOpff/tujtXSfU4/q9
GwJBx8JbOYj1eCMB4nOtYc36vL71ETKS2UKNYpTzVegFjvnuVKLXJEc0q3wpbxtl
DSif8Al7iT4zCaG2FC6Itq8IcTwlzJHyYCcb8l6S4WFAjL9abNhNcqar5J9KxfN+
oyGllgURLS1ai0FxQjmuj5cC9gVXrDotms+C4ov6xwVJqlC8jx73ztJ1SXOIYgu3
nyBbdn3UrmnXb+a7YLR132PhylT+1XkolhpkS+Q8Ozpo61VSWqf/6ag4DfkgtCpm
`protect END_PROTECTED
