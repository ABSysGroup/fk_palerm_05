`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4CecloGz2tY/zpcuZX2q23z/MTxV3T6YpUEzVdbwixvmU4kMF6LD4qRfZm/D7t05
iEnfAHDKxEeeujN5Wa/bOPh8cMZ8gEIBGFLdiCwpwxRlJrZbewo3TrcTbc1vOSNg
vWQ//1fRtWovSdohRiDwWVDkDErtpgVIfjcpXUxfUfEbbtExovcDiabhKthFGfKp
y/PukEYcYlZaPgKQpNtFfb31wtZL+bt1Vq5dVX5Unl/IycYuiNCtaBQh+1DqrWe8
Xq7cyBcDiUcEHERtGT0uF1A8rt/Flh44u/PEmTtaamFIDJXyWFJj7+zYRyrrnYXd
DCyZopG0d//Aq3svxP8zI9eWBH3FZFP3Sq6EEtqVBjQVgNR+8K5wObYuLbv4I5co
TkfXVn0XjfpXNUnBJHdt/2m/yEEaXieexYQHjos5EVy4Dinji0DfQ3AQidbkpT77
Udc9/FNAZDhGFXsfxuogZgCjc1IImdwLb82hqXd24kfKLw2vlulKCbQYsB5AucIz
m19+vmWqfz5KJGEa3ZMEpvFnhFnL+AmNuMtI4D5PS3pCesZHGYr690sr/KuZ6gch
`protect END_PROTECTED
