`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wgv9aIhCybW9AjveU1/tnu35gNSpdFQqBoQUfQoc1mRaw1HtQyB600PLOYmxbiLk
XtnSGezO+kKGQzWO42NM8X8nccLYYmoPwnyhdfeHsrFKy0JYPRbEiFdvf5zBBMM0
ArgmUdz1VAldanCor1aivu9y7lf2uOzbqamOPc2JGI+DAy1rKH5P+1PenAIlL9o5
RMCB6Kyqw4Z4M5gN7UT7Bi+CLdg5Flu0cPN1Kl3YmrlKSk6LDmWROA1QYmmiFdYU
Ye6y3D28HpfSyThdSmbnO5kGRRB7x6Y+fq14QYEZGVJX2KJu3Vzg8HMFeHuxYkNV
9zesxpO1+H+ptPxpvaZKuyg3aicfkxEqbrEqE0LTkPUT0/baXUjczhGhzj52i8Jq
5TxTmFD8TzOFp3HG+1SdsPjG1gNsC8R5g9agQOVrMWl3TMBQwPsjyOJ3RlvlWSzw
En21QyORXaBbDzJJAfnGogOl6ozpcdjCZ1kl61zGN2eeNrcJYJq2fG5CNgvkT6yx
NbiNtRtz23VYkEjZwzm6jbFq0eF7pTLRernuhutABhqAz2S9eTpo2/lldHGW/lqD
ZAPwYAiLsfQzZDUsG53Zin1eedCwpW94p2QS2JXGpnATfUO/FXcbWgkwE0OzshX1
J9x3YWQ+W8nTBVgRoHtm0061tU5/P2UmrKs7K8G/4xtt9/SGYYZzTJbG0N8N0Nd1
iaN0yfdJ7yfuAg00tOYsjjxPHByemN5ip85Y00D16589zbkEbFVB9UhDQ05m9tW9
TYClxEvH2IMAdnxPBq7m9mtfMu+miiGcyBBPyezM3apmLh8LgEtHd9ffjece16/H
YLTmaaFr3oIZXtBd0TaN0PGdlDLHeMOQoxVxpwAxV/DYg62oxgAmc2zUJvaqhyLF
BuQwfJDkBR6Ut4/ygHW3AOvLgnyXsTGxnZhQzWwzHXutZ0/ShiI62d0nkBXI49Vd
rXgcCnaeTmz3rDdAlT1VSM2OK640RQXxZUM6Bb6CFtr9f2A9bRPmdXjEJJ6Z80j6
ZdH+eSiOFVl/WRUVNeZ7s5DbwE8OlwpVg7fAzPuW0Vyh27NVe3vWbqSqeiwFSs/J
W4nCJUg1jL1ie2sEVQ4oMj1VYG1ZY4d9MvRT5eaFpKR/Ml+WeQinFFVHUE+ivOiG
ffHKVZyCVWgqhnssttY3g/MfFhv//YThebhoygYAyhmx51epQ9CbpskLGQ7UWH+w
XExY6BNdxrkIKgywJ6hG8Jqy1Tc4EWQMZXCJP0RfrD9oGPq3tqOzFH2sx9FkpQcR
ZSwEvcctmQCGH0NRiDJEl7D59LoEgjcyMcemOXuFzuxpoPeomXSt1octMObukU0C
wrlDuIjNX77VPskU9lwhQFRjzR2gmJbCseyCeqo8djBZRgVPMihgaoGdVpAlE1TM
lO5DtUnumvRPd3CI3TNEkAUktf7XIULGVRc5F4I0i6SMYWxsiTytYm3iuj2H+bVD
gNc5Yc0Bf8Y87QgB4FsF+uUe4xNz+c/AOF483BetA025vQZwjrCOUSFrV4U472ER
z5DFbQsNbEAIVvrfnYSkR7HE0TaLPWiDlxKalbx/nkdV2Mwlx4Fj2CpsdeVQpqDm
3iOR6vkEb/rVQLTzod8mhmz7JZG3ImPqXl/aEI91wwrre8vzyjxxN/zT0zZ/2gj0
XkQIVQk5gsG3byf9wzx0NoQha26U8JydQMb8xxQav7N01j4X+tONJyV1CmjeLrxP
dAKFCtayAeiskJ58wlHMr74B5Zju94YXtv0IcCarznJjjxzak7S2B/anmsNvj/48
ySeEkbabpE12FLIp5DHnOKQG1tqxEl8vc6PZ6b66u3mbH1YYr5AiKxyZCSVEM8fx
d01t8zDlr2DDAlUzxw9EiSNEl6IoCjORBqk36FUbk8XcsDQMEUwfkQZonzzfNDyh
YKdizSzkDKQOWb6WQDIWMli3UGXLhGtweZXUyycDxwGH151/OO/oWC/H8dKk91s2
i4w3nG+yHnXU0smgsgk0XghHikfpozeFQ3g5W3iIa/NnvuJqAmfUINK0j6gnGT08
7xcXFlZNFc4YgzMEKqd7lbISnf3v1ZGedIupC+GwZ9m1+XXG4Vs4RkCLr8iO6Svc
fxzjMgMwEqpdn+dX45E3AqQqodwMBxnXvF3NBCYlw594Ho7mtzEAwi8+7d8QYrE9
InYOjhmblmTKL9YtA/UKPRPbNQtGF5bwErFV7xsNWpGayej2ynjwdK4TeMHCy6D7
TP4W51c+ZH/HC+hE98o4qwDqEjKByxL2YU93d/015Zc++CVnWZJG6kBokB22jQKG
4vymt2AsIVO/8bLISjZPoCKhuGT4rXVlCuZ+R8OcsorhkEHRToAC19XTKLVuhMOe
dCFMWvD0eGBE7oIr5LI8Y8u8AHgI67gaVo3MaZTV1jVFS4HXyLex/QQgB0mzs0gV
eyMJD5IZTqD+1o4mjdnThwXO4eOTsLzEfbe58rRDTQYly8yZPyGslblPjvzRl1+h
vrsghwNglZ2EHRAHU+PNKLgwEiuUygclnXYwqPUu/E5bVDIJomA+eaDHhhJJyLJa
AeQom6VXSGBoWeqDqhBsd9ao2AtDdIvZ1AZSG9q3IIxS9ZIaVH986rbsTJQ0upLH
PR81kL8KiKftNwEnTYt74BYGLzLHPjlX3hbsJOTRw3UiAu49n9WBfh4cw2AOY6Lr
ZP/gMx6uXGEnHg1juj1N9CvGPcV9x7D8FzYYNtwcRVIROW53QO/1yIqpunP0TeV0
EvM5kWYVBBBowF05KofnzLp0Yh+kbdcS6/xw8ZGsEJU/+Vmcnd8BlfTpoHQbl8Iu
6qORoN84e+GE4Rc8lx4jp1pE9qHyCs6Typ4sXIdXskKBKdJvX2Ve7jeEdpFulG4t
84FObQgqGoc48NxbcQfCV+KBWTSLwfkYdn4a6Nu01u2v/W3ZYcm7KhTScNOO1g97
5hPp8Nv5xHfWw3xXl0IgpocyBEvr6rYR3P5Gu7Ids/44oNSDM/4zVDStzngU1gZt
9DwSSOJq8ktpdmOoX4GTkAKvh9Be0iOgU4bNUY309QF3qswGzhsD7db5Vg9Y+t3L
/wtihMZWm1y7CdRf5FR448Lz6F30oObjZhrZ7zb+oX0pLB/LBqxJUL47AKNlcX0A
y5vor0PpJLkPNCbM1BJdh3t19/ACHpV8S+BhclSnZL4tlt6Z252nQgCEyd720p7G
/lJ+lvyPPFDX5Hbg2kcmYOtUR7YD7i3H+WbJoQx5T8Z6SUtklRDzzdglHXlC1ZCv
3oA6leV+QS1ku7nJXFi2wP0eha5oThVYrKDkiMz7acSpORLzF9SpRmvOHpiOGPV9
DhUGUqy37tsIJSqXHwvYJ2V6Kpyh/bzbIwnmSZNilTMZEokWzU17BfPZV5cxZAhj
7tSxFw3eJRzNOaBN0D5ZWwC4P4r/OB0NXESg0yu4tSxL5I+mA0WR9IMGgxPjCwwl
a7IQYOHneBXPfixs27WGqHHcM3hyijLGLJz/BGQviQNBJd08zLh0DWcooUrV5rVM
I7g8fayQo9asNTSg0iK7uE1zKijTbEv6SSndEUXajGuSDGIuMpYEwaGsdVCydvzr
4ZMPDsjaZE1qKm0N+NSmFqhT6yF+4O2AZEr2N0FfSz775jas7zJjAArqtMFRKsD4
oq13NNkncun9tzZCnpc2FclLrQaExuALWyHeXfVXVDfGZoeXhzAGYvZfTObUIDMM
KtVHsCtgLsiPvoR7ZMcNc34RI6r7+QErd/mtKZiAxQntGN8yDSqsPvo1CrNs25/q
62zM6ZnH0n1mCvC7aLVB2+juQ0E1xzBcmx14uDpSZ1XhNPuEPDZM8zNkVVf/KEyH
iZiPIoocY7XSRjbYZHQhrCD1he5iYYTbB1D3ZVRrUWHmA5eRJ0P2P4qUVB7X29Au
fEdOvTuArpn2N8ow6oZx38A1ogtFPbXpweoIcjdJyU5MAZrXWKxaqoqi2vEOpcs6
UVHaGnFbQyavQ+rv5Y5sDLGix4ierZuMiL6PwpV8U/5yiYBESLTq1LrgYf0tLyW5
HkehskxNcrCdZvdJi3teZIZyqOmje1hhHXvpxWyY8oQzkD4P0P3ZxQUwemOjWNY5
3o2w/oNvLoAsSrQau6uvj81p4qM8X0v/YwtwhdiNgqxNP1RuvNb9rtxr0nVdW4W0
Pjcwp0sNOi5dGZ4mTs3yzpi6+Mn1KJD/3SJTnx5iL2HKOIE7ZDNLiOneLsJB0dOE
lQLh4gCNaoYRznveKS+5eftyJA5e5CpzABpqACOdscUDbJhUtfnTVlUwCAn/aGpj
HtpVxMkgT5kM13cDrYdk02DY6bCrUbrB+X9t6u+Nm13U3BtjgA1MF8RQaaljY59+
h/DMgDu5n5nkJ41PBit/yE1D6CkJ0pG61VPtr4jxiqdbU1TVNersmUA+bz/uctTx
AfveVytUSko7YbP9Faawu6HJ/6pw07mE2bXuAkdha5ATDJqy0xfOETylDvIrz8dJ
cmGQDDc/DQ0rMm9okFFgryalazEGO0V3xUYKxeKc1QAQ280NjMGhnL7meA9cPAqS
ndvD5OP1LYLzGckhSUat/tI9DL6EC1nJPAmvya3ah/aYT3ORw6xeifwW4E3jV1QK
TpI1+rkwE2vw8s9dHl8DZk5AageFW1bAPF11ztq5gjX6+Cq0v7cetbsNwf4S1LKj
kEh0HQ+jZp6eApSVL8tDyJmzhqfhSmB3+a10Ct9mHLRE3Pgw/SFUVG3Mou2B6Hf7
UL8WyBsbmZps2F3f8+iJWA==
`protect END_PROTECTED
