`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QT4N9sTsCGsYQRI1+wOhg2f8I+ZdXOzpJoUQ7yBDFPk4iD8TH5ksBSaUS6fFxayz
FM5smmENAnhzT8dS90TgYXKysbr5K3Jf3a/JuiUrwpZudgJkdXh0iDepi9wvmM4U
Q3/pehLaswV26pEaYjfIUI7NcZuT9AIjjJMJPI3OKNBCst0eNcXRqIIDOFLTPegz
VXU01VH1kphLJ2e2MOUiB09x7glmRYQcIlAjWt8IfNw1A1dBNu8lvz/Et63/BHYx
e2maMZrqCSlBneV7+R3asYSpc2c/iFH1lbYJ6E+c8+6wgBCO+MlX9v8idFAE2nen
UU8LuMeVXIHlMW9P+zfDvH7lIPsann0S/xdy8d/Unt8KziJuctyV+0oGWvuJ8N/W
ITe6D8W2oj6BF07mEM1MJ0Sq1KCc925nKzsTrxeXrpyQloEfbSrpnW2J8G4vEbgw
0Z5+tWFCBwqeZYZ+TmSUKRtI5KTuDEqzH8Lc2DYMLkay0C0nRgCRrbP71d7SBJx1
bMss2uzfT3faXIJBRQBJlncqVETWBFsf5CrP5bzYfiiMNreZCvfCQxtCseSs7SWT
z1TVvhiT2ps56EsYYkOjO8/2gDg9Ls5/vTRdzl9j16IXLfwGiu9YwCN0wdhYC57G
csBZsyXfNMCEFSUYdyY3oEzRLdjVQ248yc/ggQWlzZh2HDAVpBZAhE6ejNtT7OxI
7wDVY4OWg2R/WxvOTMO1k1ZhewAY+5fkHh7tYDouBShay0w+u1wJOoBTrUDGDIS6
stfK7QkMdGc22vLGVrvrgtZyDpY7mFU4le1m/3v4lJaT2ZBAjdY977ySmX+fZ8xB
iGTerprvziosQ0LjoAauNn68Ox+jRB8NTgZ8YwRs6Cj3cTEjDykxpnjkCMi+OPAL
kmg20tG8lKrxFnKNgfYNw3zWLMlBv+NEM3uWoyOwHhtC8IcZPVXHhIDjVploNabx
PWCrv3Z0Aasbpd2E0dVdat62oUga/D8bxWO85xDlz9CsVcrwzjdKg5r8yf8JXSEm
uoEaQl018ru9/ow4ZpWN1z3Yu8+RWnvmCjvKFSnMazpcxouRrvchLH5KzX4psDi+
pQVgJ7I3kuxxUYyN4gqo63mG8eafM+k18h00LrMDsDNjdQhAGmLtPSuWkQF24W56
EZUF+I+HAEnRujFh2aj0W2GtM/JTiSEAp3UvsAGrX0r0lgZ+QPQ+ry+PN2m7NjFg
h0FKXg3QVqCjm5z9ACr/Z6C09rUkmszlp++WpdjqRsfTmBcaK2DK08xtTNEflHhz
ccEG924jBnayazO0fMHKGxfrrfLfWgx1P0MdCWcRMQ4fCG+I0ACg1INtntbQDbmf
UgTvgQJvnxiLPoen9JmZvtNk01fpY1Kh3HGU26xoBhKN5z/EnJZBbfnLVTtfW8Dq
BzDa3AE7NVo8TySmkRbM/f+o7vv8mFQ/Jwx3cK0dYuzJ/yZ8jAkjqo+2N5vJDv9q
IGM04+2FHI53xYmD5aI+3cbyN0VkyMLoAxmTtgQZ56eaxpWqV5xrXw9iLd7iVWfZ
pVDFBqrkkzkhHcnbjfZ5rnl5wjaODXp+1T61UVZmU16lapBERhQpaW1tPm/IH1ZH
GcWaTHZkj7f9xR4HEWfosos8CNEIIhwBXHouFRrtv9J71K784l3+aDj+Oav5ssnU
x5CahVACRgsLnYH/jsEfU/9XmGZAllDwgLokwDK17wA5E/+PRen7Vai0UH4qmatk
H/drtzaNTAF0Mrn/cskzr/ctTcqWoQyYYByqSBTUc0QmaYVfrlhWyyT7RWPCTbZl
j/rzqvOFJJ9Bf5C9VnEPwt9x4SdjcyI7Z4bPGVrAKUrVtKhHsfhcdiT8FSwrsauw
iwbGb0hhFeS3bYm11zedJQJD9OhGaRKc/1zk3EP7bTdDwwSPeQi+SaJERDmNEHIo
7lktYsDFsWi9oBMrqkqdZic/icmcXFRH0DZGkx4fqUEJv4VVPSROLWd3vN8Uuk08
wKLecyjLGhkgXIib0S9lhvuv9tc4t0BQDjwGE61SJ+YqXb8uodA585165Uw6h+0s
jZFyGe3r/SUZ7or4iKwMo5awvBbk4IhC/QmiODqzqqXNrW/uqiP1yS0p9GXmobSb
TPDu9ouRGRGFrGJrNd5POdK96lCFpsZQi/CJas0OdU0FBAEMx/KvGlAX3GvZV1da
bGKoyxpVGNqM+Gje/LszEgSwBVAO3Y/TqgIUPhOWhCJyOGwc8Od7KvZ7NCst0bdz
ZrO092Ym2cWTHUa+rFRUJCanvBK7mYfWUiP5q7nVOu1fy5wfy/2FpVll8oa7NTJh
ohXf4S2ITLQEmMi28A7GenbDQpTooiZ+eRVOqBUV4pYcpt0DnB9LyiGgWeQHM0gg
RjzSdOfHPRmfQmxOpxlNP6ZeGvgu5RTPvm1xmpKaMY5O1JJAd6D+kwFEdTLSsoAS
/diDxuXLmooWZ6TIVbtipVV3mqF7IhSLl7XEprcVf4mGZMPmlJoA+37yNFnQyn0o
rCr+GgGWL5775CSZw7c9Jze3nMNnXeXGRzh9Dz/KsQhx8cCukp8Qw1EozYGY31r8
Hz9nrvyiao0/FHcZ7ASQotHx7ymSbNs+MlIExEwAONlKUYnhO5AJs3lyGraAAjvk
I6/J4ZNAo+Hajyx7ATzrPofWtN4E26rtObG+e1oO4XzvZiVL/+2DEw3kNyWKdF3W
19oJShZ8FlahRb+37ZYeO/cqnbLGEIXe06BaAmNkt074sfrW4QTStPu0vx41kmoW
`protect END_PROTECTED
