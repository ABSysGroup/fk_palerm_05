`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GKlq4pizGn9JYGtDKNGnUbRFr4ydKsOMe7XTNmYoX1U3K+KzuL35IuYOYc9KAICc
rYZeEKLWFayYl04mSO+7Ld0NcK6K+8zoO4LQwHOgBD0faZOnNmECJ8gpQR2FlsIk
/7ik2t54dmY6tMP9k6y0Kq/RZZim0BLF2TJhq0BS+CWZmREJ3VfRRVVvN6ypc/9H
Q7uTt60va2t9pd3bP4jVygFYu3r9/LP9H/sn0VFAV4+qcGzo/NpJB0nIercm9RrY
NHGzqUg2KNnEO8v8HoLWe8AwaDiFXZQrF09z/nWKAqM5HmH8EIUBdFFw5eB126er
9oHDUdDZbP7PaJvpQLyDETxr/iwdrrhNOyT4lg7FRiZoktSSnHjAs/Mv1NEhZahU
9Jigv5cWOIs/ULYWppKUSJ4MKxgJRgzHOGvg0MDK95MmQ3Md88f+DhX1XO3Okqfz
wZX7MKqLtD6EZVYdFwSS4jbj37wZu9WRznNi3vNhDW44YL2SvW3mUEUsPIxxmFD+
L7puMIXTvSWPBP+XyaZTqki6nnwQXPz3vVHLPNoyKFjGbVdPSPjaTI1F1dk7rBsZ
bqdVL1iaklp2prfMLLe6F3W7H1Hl1Dmprd/sMrzkt1MIQH+GKwI0tESX0Ky5eG6V
YKou4NBoqoDoKhh/vNuICxrzNCyx7kikae2F/t8SnuK5KOw1g0gB7JqEcvWluo32
/PiL0+IEhTzetFfC7zZ7xHVpLfh82K8PRNaC+5hH/S0xjeKgMvULJ74bBaw8CpJ0
FcY5DSzcbwLcJLTDTm9fTeY+bfFpM8xc/KUJ8jZJz0BEnX7NJwwdyB7LFGgE73h1
9blMCoPixSqg6CWkaqV9NV628jkek1XfRC9cEb5QuUR0AK11ql6mAU87IOvIpEk1
J6NIit15602kDQgjlJeRKFMyyAgtj/h8moyqpah6LxSVZTCFRqymfz1yG5msibBR
aTcR1FV+AbYhmHy+0Ubs8f7X8DyToz+XBLRI8GSr2mtFJMZxJMRhl0z/0+7d0X//
pEfEFQw08ab9fISM+qeVnz9lQbdlfl+qAhQh3kklUD8=
`protect END_PROTECTED
