`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QaiyAjlcBL723Wc4K6AJmqbh3jBhkiuuWd9wIZGnTEEqBCxaLl8FIBYnf1RA332j
MiJQalM4jRI0UDCFHLybFXbsYsPTy7ifGNMnIu95B9FZzyP9jt7sslaOXKkfSsnE
wgemiGUk2JuQfZB2FUzqWbXATcxYrMo4Ay0qPepf6XHi5eAjd9U8MDemDIdIo7FE
x7pL1b7F4CjmHSWUz2pb0zs6VKTEuwdF//dsrH2S9gz7xraJZRFDup0YTUxYeTgl
cZ1ps4lIaR99ZPipdp8c9r5yf3GPqdxFfN93imYLE/9nRLjNv0Svdz813wc5LI/2
OIDMDuVHHFBUX2qvU0G9oelTjAHCEz0tIo5DJmd+g8JLNWvKw/PmaoTnhvn21/kp
jXwX3NTJ3NXM4q1fsv71+cvLykUBYgPS2O273orcd67iruVk8EP9DxMrWfVPlrf0
BQUbw+RLBqAwY5Bbbf+xxrzByaLzXK5dPx1qeb6x8Ijb2i/j5uiCBwkPslZQUtdx
dU2yaL4PpU0FSNvVDatysjlxTpog7W9eKm/gVg/MGMerrZfOw3QskVcIkENYO1T0
7GC4JFyoN7ZXSgNQ2x06CoLT4uNSI1AuT2GejURo3Cg6p/ASdWs7Zz6COyUADEDz
D3iAxdjvUSCDVZcVR7IvCzmcjMXtbK+7acCpNSiqf9noHmzqTgcr0HdXlC6qrhuk
qK5vOrjm7ct/Q1+wSBE7Gc2qLzkLDm6AoHAzpBOv+wNNpKfWWg1nq/hoEKqCX4O3
`protect END_PROTECTED
