`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qcwn88+W8+4Mh5oRTDITeiacF4T3WWapkgTOt4BlTqcNO0Gh03UV7VIcii7nKq7r
LWPTxw/6BUM1N7FapjmnCtdlWo0pOYLtPwUk33DTD7OVhhDq7zGpjRBHhJbcOHiD
sjgn3t+H3NnOVV1oc63HpCXBkEwGpZTzuSFJf0ST5W0Bk0C0yNmcE3Vpi1q6NFfo
1UVzZYgxNG1yuzwi8Hov0g36zD3TdGdL5fhJT1XPrIRVe5mNKfXKrudR3q3DkMCB
tUVPqY+4XMcPWwvfKEksl//81EgZhg8/+Y++ZSRxGU/eud34kY7levV+sxPtXCqW
zVb38Y5ZOMXtMPjKOXWe5+FwMLrAEYzYai1kNVdS+Ei+DhHzTJ8uLZJOM8m0FsAr
rAVl28Qg3i6nMRHWtji2GxSdjVfTZMecXe2gsWy6Kc6A3R8CKH3pdA5ahv12Uiff
xeqAWMCVxMY4FDYS2pAovJnU4CQromciSojPJk8JAKFDkDijDhtIg0FawmsPS8yl
8KXFrF+hytnL186RnKlkydKPP3oiclh6UeEYyKB5IcmhKXma9e/fy1Ecf5oxCtwT
1U2GgmHSf7g3Od4u+ITY5BmahQfOd8CzBGsk3gLlaSlCtVVrphp72RdjMALPCGTe
8ZN0PjeoNSerSvZh8OIL2j2RnBcD8QbJKSnf79aWQVHbjAVhq99KNVN7syO4f6h9
SURyqkldOlEZy98vqjgE2qpGFZd3DTha65RfxcL64GY2lD0QCPGOVyCDt2n2VLiB
ztN+I1s1U5Ahm1nosN1OCuMDoTiwR9byeZGUujnIhIf53K6ZMLgc1t1H5QyYrq/8
6HdUNgPJIzq+DGkBnq6ObSaad2ZFLm4sliIOvV1vRZnR/AoqdyML3gJabR95uJUR
uMt7BP3znx7vqS2kU+Dn1vVDTvfw2j/ClZgQK1gLUqjU/drY15hZuFISgHnaJhKi
CwUHdxkH6BJnc3VxKxvz9jcUrsvWJEJuBXXIX/TrMqOSK5NKZwpIvBBHPtsgR8ii
IJNOUTVPbPVJK+IG+GIgRnwgPElvoI8R5MqxGjaSo474oamotgbi012cuSnbV9YZ
apQ/RgMS9Gh+2P9OEGTYA7/AVGuLwj+LxZqggcQxPItATwgjPV+2i38GDiQUbemB
ydGSwPkpy1aqsmrEdVlZguGKE+HHBQWVRUI5IozbHsgINLDAHyJ+RgHY6xtF2mgi
HcLUwtGgGhSbA9WNXOZSJgQu/FfZcb3fmSD2qoqxseXfjLsKDnkBpNgvUSWNTRYe
/1FPWi+htTbJ1GVY/t05jb6LhzfEVUh4SRmv6cTie3JEH81/QiISE8N6cJS/czng
fVNzpdp43STYf8SQJvJOkVilWYljmUv1a0PDmL2YF9jMdZ5RcKmMqXjabT3hbtct
7z/o2r10RamZJaATBM312ytW4V6FI7F0QKbKHnUs76lC2O0c/F60ma/ZPEsRWLBN
59wRXN/K8EwUZ/7vHNMNNko30yRjCJq+bgaH74Z2rESJzzNj1ONI8C0Mn+ZPf5SS
CwAUFRZ6wfLm22JC38spS/mfTyE3Uqmb6rDTsZEHOu5gdeN1VZ1h+Ep8limO+ciG
3mWuPfOckeBbyjks93ONpefQs1WEcHJx+5Uabig6QaZbZqVXN3UHD9lD8/epL7r/
YlHdlUN4HdCk41IS+x9ZgISSk8EIM2a8+sbcF1BBphClosHtyaXykLWeqIinX+ni
KGhhE6cY9bLhRodBwe5znDdULX3ryTRI+ZQh1NwAD9+l4C+suYXwEAc/6VX5p3qY
R5Q7zB5Z8ijEarmE9TZLOYOttcn/Rg3fAi/q3J9IMdtJxtAfwwcfkKGhcN6DlRnI
FV15H8XqE6OJdZykquLADcGVp09JN9COYtaHjjja03GwJSgUSFtrZps16sSiMF+6
40vKZS0lR65e2k4wagvlXHaWOOpf1vaIaRPTcsLekKlcA0BH60x0SdnFwPojNj08
uq09AduyrqK4VNnBDzHFoDrdJjIL+rlfOetPrcI10GXOAH94zoUamZRdp1TtVvhm
MdEzjLS854VuQ1Xy0JjMIDA9n2GsXOUtGZVjXFN0hUZ+PAMV5Uj1baekL7jdPU5X
LwK6gJSQIf5LGx12tP9Z9uwyRxns4ij706+ol3GGbu1k+cv81lyRDmsuP0yP30+M
1LPlq9M643vX6UFNcISN4g2Y1Eeho++jO1ukJZtVhokjHzZCfOc2wNiRGZOktj5U
O4se2oZyAXoJMCPuyAuJ8IfENIpRtjyN5IBR+WrvkGddesMpr0BThpSDGUEkUuDS
HXmF2bnTIlLHrV7p9Dv6ohqdKrXAwN8ZhAxJJMt/MmuV42CzSNVpDX13DscAVgW8
aAGTIVl51yZIxXAqLoRBj3Zvexeal8tcuVN0AfuxAtAZkZ3Xy/+5TGH30B9zkIPZ
6djpsi22kgtMxs3OSSIym1U2WmxyFOVxNCnz90majRjFg9dFC6ha9TiRnUHKuhGG
hPp3uVfRGOBOiJ8m4g2ssd/Q2sZtvJNMUB+N0z7eNSnMBON0cBaxJrbnkZEL9Voa
NH1vsmyijU97yqTO26zJI9aPjMQ+J3v0ZYphXlCyp9aQpfDoZbzYPaylmttzJG3c
jawxbW66cdOT5Fi38geo4Dn6r4cj7M2P0NS7OJ7YWQ5HOngmkGSGmiJiYRxxSJAp
sh6W2uwJbj/vwWRmuJjA1qqlJ0PFDHC56WTFlr1CIXvT/V0cWDvNZ5Al8ky39Q/J
IfcG8naDSHw9D9g6SF7+/gJWOnfnQVeLOtENn8COHV9k3ktXNmmv7SkSyHck3Kg+
jZTw1skDRYS6xoxFc8j5f5xUAZpnxDAOVNibQ0ITOwZFlygd5pSES8nts3zQKiw9
bR+wEvi0fGbCvtnmlNOK0XTk43POUi1DgaYseM0Bq26cuyXxaBzXTlOCjT4orSyu
w+f5FSLjeZLvQdKZ39KKYq8xUeWg5ydCI0bMeevxwjy+iZ3nHdR0XWAUqv4jseKt
R+SWuJE/vWO5Avw40k8ya08Q3FF5iCvfaHelvflqXw9615s5gAg6pvLmOSdcnvhI
GerhsBb6mo0fOv6sCQz4qpcuF+QwExk7ZO6XLw934rasLyKAlK93xVuU4n4/CACw
gMJkyqQOFthG7b2pnuihbpfDKOH1unLpFo0czoJk7FVqHtW9K8NLnW3kN2ZqaB7B
Fz7lnmluOnGF/0qRLo92j2u7UF0XfiHpW9Fa7y8qh62XjMSzOHM3lzI606J3N3WD
P78U9Cb3IP6cbkdVPyxcGQ5ISDKk7dMXOSW2GYPcNaixtcCn/aeXas8sYhXopUpO
dMcO9okeMf+xxc94TgbD4CL2hNXLc8vSeY+dGvm4I1fHvQEIwByRBI7sPtSemz4A
ddREoXg+50OLoh+2DtmI51NvOgJToO61SrFFrIFe+fGWqAw5ccvTyUit77u+/UBO
L3KGdwaacnJL0x/rodvUyCaLF4dGdIDpxXU5c78o1iwGNqMv8W2u5R6h0qxV61f2
51upiXhbuitHEs47BBZDMAx6ci8q5DKYt13pjwhx+uBtyJEPjLmtVyNjHgqr8bsa
VBOrGn12YRx7b7yY6L50J6Eb3SUsPnuXlLtPLykml2HPMla0jmQdjYGnph0EwKDu
tSBaL6mpB4+Qe8KtZgHBgn21aOq6UqOaEjcUmbT+OF37/QOa3NV9WekX1PUJJ0Z5
PQj/U7qoDzip956TX/9sz6I+Av16BJUUv4xMbU3RWckt8wrMEBLKCrZ4nxqLZo+g
0hPGe2axvkGzxnShXkxu4A==
`protect END_PROTECTED
