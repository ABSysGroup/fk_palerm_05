`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OoMFKI2FPCq7JABf2ZqV462hbdlMwScJDWIGg2wTX/NWH5qM88HyXO+o2C6aQw/l
Jr+e6EweFo7/GEgnqEuKIoHLTSnK9k+NkFLga+X4HvkcKmvLWWyUiiudzyG+3JUk
JyCuEHprR7ds46PXRPOrbfS6g6tw9yAUuHmLrRHlaEJ96ReT5BzeY3DKMHOHJIh+
tGfnUvpZ3l+Mr1xR6KWLjtiJ6Dt2cKx58ArtGaZlc1ETz1mFs7+Yy6YUUQ2lKvsZ
4C5LvL7gyDaK5tk70jZgxGmRqyqGY+sp1gmAoOnr9XEFUAhyN4jdQRBOt+CFGQ6G
+yk4wXhkjeu4/XE488595W4fH6EmDk1o6ftT8oip7YZZmQCrVE1XYiA1zJ2uhfoa
fiRjfQBkQ8T2ujazg6pYQhYNR95dMxqQx3iKcdd3fpIdM3T1idq0d7Y1DtaMgdhb
qFzgqKcfP7JT/Egnjbl0U7YGOH3OISBMHZUcHbroTL4p3TVWJBJXX67Q15gIVVEB
wiYdkq0j63uZh7CJc8FMF1TEdoxMXNp+9rU7SYAR56Piv9GrirZljXz/nunZyWq5
WiBgpLXxLGjJ7DNATKBIBbVSnMTRlk5P/qU0HSn4AR0K7gcyaJXGAnWd5i5HjoMM
pqD9Da8w2lFncJ8rJtCCQjJgRdoeoGd7DcuNrCc2W2PDV6U8VDW+VeLYbL4OkVG/
hv7sB2UGGwwTu4evDDsjs+ZfMYAQ9Fxype/cIl4+1YXqdCd7kmA5CO4ufLKjRTG/
i5Dw73y87eQRV57rn90sl8ep4Iw8H3Z+V2dN5NghX88BnAhnQmrd1ckN72xCFCIh
Bf46vv7d9yexkhJmzg6oGMnOzQ48hRfJHWL50OuxTF8gCa+btLvdLU5aMDwu4riE
GJZ180w0LJHsJb6WXoWrDZbM3SsyLjk1ZgcbkEurVaT4poDgCUPwK+qs3oYCeA8z
Qt5SDOW/pxWbz5gUMZ4F6PjCaIPTmzsvMq1QT8L7hHY2Gfxs9rCt5etp3PpLbOAx
j8mq/FLah89MDupp4ZPxRjnERDtEyOjFdHZecEj5QTaC0K3NjW7XvB1Ljus6EZ9y
d0GIbVbBwmQs+wlprHlVtghz4MoNKkI/PjoiuKhFRCF5n1uqoSvtJD/AkphdiV1I
WcbxXblFTyGRfrl6TXTRuCa05dgH+oPkTeLxR3a8WS9eF6rZwApmycYDmTd5P03q
eB7qu6qroUiipP0bp49mZ1jwx1Xu4NI+FyX3yGfY5uqC3fGsY7O9YDk5NofY8kZb
C3dPwRBIz8PHbJKAyzYvr5HwirTMqJ9TtssKaokrX0BCxFp+xrNVIQYRGDX8KqQs
uh85LpD8Z9vwrrhiP8f1WvczHUUKLClTDWHIx+tBGN3GQa2cXBnr/M0ooPm+7+NX
DoWGG1H+jlodMaszcOXz9h5nhlGBLpc64LE2W8NfBtIIrSvdaxmFR99e2+nELwdj
PTjIj0ajIWXEvpetUF+qzN5CWMFBqiOE+l11NdUshBTwcx3ao7BNFTSjHu2Bg3/D
iI6qyKLuetNu6QZtbUVf1laO4Gj8lDAKE8oeQx/3YYq42BF7x7zNnUj1lChqNba/
ofafK080TjB8Wjrh4hTb0wfKKSGlhY7cAwMg7klK8AemVCdOU1ET4rr7W5KICk/a
y6mES1kFLE7URw2/rWTrSW7qns7dsHfOQhODoifFzMEY8SZ2ty5DBXKPlGJ8w054
PiTHK6D5P5NAw5/4icJCuzTeclmjcFaudOCTF3AjsLG0H6RPQ4iTIzmp+39ik7RB
ToANwVAAmfyR5rNoKdQ5ur7jfLw25fidkFTeyt5DEl5LD8MBUqqWjSMox7/IbglE
msOihXnL6LdiwFQeFFOHgp6FrUtWnksYXssRftUBf7tyh2LEFOYeYDhzM6wpXD3p
25wTXyRlCI2aCcMBgcCKCmOnf9Wf6G7mypruYYun2PfUHPvE+886DE1C8BgMLf8t
t2ij7NzsAdC2fHPYm0Df+nf6tXSYrPWpgAOObOmSJDts/WpBKO+QUk2U74oMzNzY
7nIMT77KTQ6Ohn4uOsPx229oyZFIo0zmJX3khNXY5Y0GsTyRy6sJx0E3qR37bKd/
8QCOG/JOWyIAbHhqsMZCWQqS8PH+MUigUaEkqsFwPJ9nBMc6/kU3nGFdXTecavoe
8kK79iB+k0bnHLYhBMPxSzJFHrSxebAzwidr+oq/8F6KRSRPFRonEkRpwDdnZkGI
LUsX0OAieX5uAaPtbPUH+cPR/1LvmJ806D5hox1Hr6XyNeql83SOwHA+5mG05gWZ
7lJOBIeBoIjyPKMBp3k/aPu9PmNXvabAeNVu3e2WWpmrg0IHp1Y/JzVZhq7d6Qka
1HMa8O8Ry/SYRBnMly/4+/KQSQjVkPUr6MtoA2dYo3P90Kn9c0siOiiEDmnqPQR2
3kcuLdNb+Vj2JFYql5GF3mMuUp0BizQyz5Lp5ZxYYVwBNdm4z+Or4VAzh8gUKpek
RaluU9Q/9bBVZ/dyRbYDTMnsVk2aZgeOGRyZwh+hJaubcdi7gxqaFlVLWyYJTxD/
oEKZMlMg2dVr4qFvIGr8Eej/OQzBGKuMBUKOluENf20bhrPISe8CAL47ZbTP729d
WKpak2fsZfpo/O13DPI0rE7/iHhPZtm1Ki/mC4InSNszTaC83w/Q5kqmKPsLOpPX
OujQX86hJ08rQXYfCmCUqHpcIa3J2lhKbatvaQbM0w1bakR5karqKIk47Sw3/PBv
DUgY3D/NbaYSPzRn+TqEBdgN8l81ZdY3vvD2p0r/WtStxZieqbp3hpGQnGE1ce6L
Xq9qe9lXU2bv5gyiunDjMYsEpwrfxnrO3xlr7OH1TD35HxigWrWuTtSoBYHBK9B4
C6kn7S1FlCd4a/olX3o3j+9C8Cu2FtCf5AKAadV1dRgenqViAWi2oTWyJQMFO+oZ
c9g4fZLjEyRQz9X7WdXF9Z39kwTG5Jg3Ji9+GRLLGUF+kVwtNTCCChsDJ9cgHqxD
9wh5UvK7r8btlaTJHeBokkzaX9yjkS9IpGsY5vR4qhNULABhQ7T/wIRE09fXH4lW
O12i0KJjtt++W14shuKx+AWbd5SMm/dDwhwmzYHe9GwyOisDEvufe8rb5zyGJiHl
CJ8xUCMejU9aTVymu79ySyr32SjOK/usMdrzm2HaVPnHgW4Dr3DBJ8iJCwWzVkIW
Wb/hGDByKnbkov7B/S4TWVOA2wWTIJ6JmATrYhr9BYs3KCAGrX1MLLFUychpOeUl
11yAKIV1qGVVMPHBF5X6UAGu5jmiTKKBCPeRdPiyYLVAlrBN9bCJFKM0rtD0PAE4
A5dITrD/+FutFwVq7XAWk8sU00o9jjKknBdDFE2rxuEJNEHFL1yKcaoHkZ51Rny2
WwmVvzarBJdMV/6/FchtoD5AvMEN0C/MGK1/38KyPEuKFNURxBaeFjEwnLk9qsjD
iiD3Px93BkvqOK4PcuFAwLG/Ub7tITR+sjT/rAwyBQ0bqiDRM1sPWsnt91hSTPO3
OTxT6QzoW7XPryqJ3ZDhl37ZEJP9p04bBwk03jPhq4J+KOUYF1rdHW478eYaYZtL
SZwh2UPUqi0H3gdBx1gF8+7NuQ6KurbcAkWLKysuFpp8psvOLqmlErjpiNZ9/NqU
Qyh3CxyEC6jGMQPdZmrWO/uaRDj9rtuxIckryt6XSXRL0gjS60tL3QOc1QA4+tEm
Aap/R015Vk9Y7WQgjbWCgPCI8ikS01KdbQASTeE2wODiFRusWgZ+O3vT+rM7yNn5
beua5HCoPZK7miO88QzVGW0ER0+AYpPGAbnH92hV7cZK88AryQkNZ7M1LILDeU9q
X6eyT5wrU+GvpFeMlZrj6GoZAwIza/Hd107FznpCrO9Y/6n1kpgR6RXt72hOTnr2
N0X5dMhqXDBQ/Ma60R/6gNZGwcCa1IN1AUi4Z5PY1eHP8wL82n258bDlErulcp8I
oGnrQ9SUhAdscTy0S6L1H+zCeT9nMdjKXkoXSoYVMKungMh7F82V7oAB6LE5naLI
Zs5SQEMI4epRLB0HSWLNDJk6qBinuhN202J09KhD4tsCqcpKkw2Q9xjZVVrXiawc
J+rxuzfZ6mmsRUwX1qaFVBONGLbEwiSDWTNfua4hewFAVOCgrMFOHq65DcHYzZla
FGFyZ6uMDTVNnQBpLbWvZ5NbyhgqNBxlxp9VV9BtHLl1m4mVX/dTDBanLhxDEISC
fDKlqvWRHmOwNzFEjRK9Km2o/SLiAgi9IcpDoU1tScapCFt5wV8otvTuGnGprnT4
7csLnwUG5JZEgLc4NDVHULZcDOggEpZHPTN8/cxy7zYoRyCgDD6qgUZcyP5SR1av
hEJw/0v5HwPyLdWz6erNxnlIJB/IjR8fd/HWKeZCPRdMrBHd3efimXgDXlVM5Fdi
SxiuLBUkUhB2d8d9fPsu482quF1LC//bIUwJMqVjbIjzbIlkGzWNRMsTr6py53Tr
j/XBKG7Bvnz9c3AXkrNTgg==
`protect END_PROTECTED
