`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cw2oD38dvvBYq8HNbVUru/MLX6LPpXVR4h8SMQOKxU8AZDxpcjkxQLpMHr/ti2OT
SwjbppA9DgwzAj8qBfsAaSwE9i0KktWBWJ6f2zjT7gImaFRlgKhTQuAQL9VwCA5y
O/WGkXg0sH0CVGHojwOaamgEgVgIDZk1VbUilK6ZtjUOAHcdDuEOIm84IxMh8y7U
RPHnuY6gnzQTw3AoHee5lJ+jDLJbzQEAhZR+G0hU/biXoco8dT63chQZpvd8JAQl
tKpZ614MPPkdkBjVWUc9hSR8OTxOb5aInN8nCZkzKlvJS+NjP7x6bQJzUnqrY0hL
HwyLXvwbaX9K4PmeNKN9mf+9/lWGPCmK8WxHZyRnZVkA8U1yvHgIKWrTVD7BPhO9
DRv2RxwKh/TVaYnIURiB1bIFOelJDLfsNVGz3R/SEr8TzYATiAM6xOzOLWBCSsw1
CtvptWFOCj7sIjWdhnCMC/94Rzkt1/tq0I3hvFFMwBV9x/koqDhrMwwsyTCjwzQQ
qgeGW9BH6/FzMi53PXleTnJd615brXegBleyif802o3yTR2LA44UWByZz4dzaWYT
GF8LB1EvD/aQmpaVLzPf8lBmiM/j8roLnNaW20PujT1IooLwuOa14zfW5cIevfAF
9KenSII8QpC3Rbjfk1R0d9NW3bR2PVKIYXvAPVIZiNL9JEX4pR1OygP0Vy7/zM6k
9wPTiTdcN/7ZudFnvSTQoB7Iwa4hfn0BhCYZ3nOycXYI3Oah0LqUbSfxqdgX5p2X
`protect END_PROTECTED
