`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rfanqVcCAZAGTmSfdGVlTaMaRM4OvbI+Z+YZXvL8TpGtKGsggEoeshZGBiJGPSu8
g/wt5wK7m3z+vpTEkKG10ZWqeS72zqCA5CuUPlyB6DuJ1SuKpv19ZEqS5WDekAvG
52bW0HBHOnUKSoE8JoiKFByyjx9WypH6vGCTb6TGDW99oLoTQ1zpjPqHkMTeh+6y
n6SnffgbcHQtQ5XC1A6Ia5FYAdvAH4vEoVhjIEwMsFiEjGWNdyHswvVwNvq2jKl0
tR7YbHzwKH6lr3a2QTbJ4ZY8g63TLOjdmgXB1KRzG5rrvFB/NEcHEknYZUAAcMpr
wZF0b3fQ+AjCfrDnOWx7k4kVdzwJbkqqaK+xonNbiUynzWOAmD0DzWcah6gjVxhj
zlR8kFioPdYdMgUJjFCKjzOnBeh2NIE5xVHa1PJUXglwqajzs80FoKdoP4XpwNRn
mpksb/oeVFmaUmYxrAn9x74T5V47q29TL3eci+JCNz0kuQgx2r1zNPZZdq5DT34u
BFgvj3uPIUPwjt5S8zQ6tHJ4OSVj5D+GbIDL+/sDZ+TIgr/IUTNfPJbSRW+h+T35
h6V98wd/MUtV4l/0TAaTXS4aE7ZRKocGDa9QTeV7q6H25hm0AsHfx99oDzkcUL+c
EpUKTIPpF2b1KO4qdehmpDGiX6Hk6npCW+c3DA6Z5JsTQQ1JEs5y2rr4HabGfiI1
8QJGFaGezU5H747JIN9h5j4tw3YKqeuoswz57rjspErqX7Jdf1KCf1EZ4NV0ZCof
Y1R+mBbyzMFM4YPdf/y1cJ/3DmjKetru3gUl8oGmZ3jHnxy9Pj1xpCWRFxD8yp4F
9M2uGi0gXElf6aCWBIFgtaWEPyOu161MmCFgf859phG11y3PxCZLwcwby6Ijia7A
v/LyLIYV7qszmEoHHm6XKb5o/S29pSvQTc9tm9H235jUNyiI438UUN+fhaHvpUWN
UyRsVRelP6PTU8sXtpTcJK3fsV5ItM48HN5L3RjeJvtvCuiTkZunfVxosrURNXj5
rOX54vLSK1hXYYMhbSpdTIDHmNGTs7KRsjabbZs0xm0JghuQGTXZDpL9HU24v8PC
4MwrP/zUMVR2Q9WKiXvjrIFewJW9GOg35eoJ1ATg+m9b5GF9n3Ptx5drfZiHETPj
eyMwWCK7ZgtnTqY19fD4uOE4+R7jo8ti5p6s2DMeScKGAfnEKe0Hj9QelUWQmC+b
ABZ+UjcU3q1APQ5MujtB/rJyJXfpDheU7oVn7xkYR9KL4HmyLAx8R9on34sXJPkx
nywHqW6BRikpGslXnbo2x6U7XWa5dE2wsrnvcEU3wcdNQcxtv9ixmuDJ3YjcO2Co
s/9QiI7vBDcH0pF46zv0Hkqr8Hk7PDcVR09rQZodgrXvhzS99C6ykuxfT+AC7GvH
Y9CE5+6jswvwVl26HfVpwZ8EGSy3gRmEVdUFNNfAtc/h+dZPNd+nD+Us7enczWv0
ZRqSrqnHRYMg3LqEfArC6Hxmavjq4LgVauqK6834me+WbMvgoDTcP3aKzXQ04Iej
UjwzZU7SST+45Dm8XmXHJz4Kes6W/Ha0nZDtnU3TV5m4JaSka8AG3xWLLeLHgAMp
2cNG00kCPi96ctM1JCCAu5VJ38gPzXl1iDAb/cnHzjqFjxKeMuJwgCi4yTtwjHf2
r8CLRC1AtGj+QknWH+RIXAjVUlPBltGUh/Z4qMjMg2Rduha/lhCLXuvpqy6drEjW
n6JiDveQbMhuw4gKkmFHE2M4CbNsXfUo9sjAvo0kqhjYM4P97hqhvuy2AZdwCv9M
QmUn2hmK8ciW8y1DltYiBG6zgr/uGvgdkCyC0R1WF70sqlV9ZCZafXn+X2g5mzmw
mcaqCeY6TH+zsXtj+fbfUICOCXDCotm7rbid+McrsnePDVNNsXh472Y/4cBidXu3
0m1xNJ7RTefCqXSIc0l4UfWzokzVDP39kTVoTN0FOMcd+3WOQbeAUFjw6VAOW1l3
c+HDVte5ZOkPUacD5ftP97LeR6KfUOCy4C42gRNHvTmA8Q6kgwFKOZWuHq+4bwZc
W+v7lBoV0pvODk6xV8xg8GGsEo8+Kdj/h/ClhHWYXfpRK+tU9eeYcZLZn/3zQ2n/
g2DYnpN0eGfTYBrepvPzI7IcZYvNMveonh+69IVarXj5iPjwuJDstZ6ViK7UQC2S
Rr30xqjnT2+BLsi7nVWWy4Cwd5zP7rSSg8bjJPNPdgHsYTfm+TyGRSix/ZXT8Zb2
mC9zWYGoKOn8DFkKukuZ+bNkTL8Ddi/d2fn0lBtcbDt6t+1O5YRSzFxo/ayDH8ui
u3OQ5QJwEFyq8F3CO/VP0X6Qt3kBG2p6gs1BQIWVk+9+PrOjjvNB2auI6AtaG3gw
oswW/a7FJW01C+ehcZEp+Q+5EXFo0eQB9tFYNXcv+bkLDsILAerj3M4Qc9wsrHLU
j4tnW4kwIDyXLWYSpbbMoJNVZCaID/9rb/XBxzO9fAiOdLE3Jdq4ekYe+xMy/RnK
R5shI7S9xjHKt6QfnQZjzpXZGqw5Xzb4R/luc/UuzxFgyYOgC2LCHDMEeHUiZQmW
39Ug/KQzmPIMSEtvWWslo4OZD1NgrE9ZREsn0Q1jLLVvbxSsKYoc5s02dpsEYeu9
7A3ACg3u33dsd0XM8pprVGttxqv5Th4HJ53ydrqf7YbinakvnpmTjgI0itvdTWZM
Nr2uV0lNb87yA1bLnfYFYfm5e04uu5Fx90sBRZJTKY1fv/V1vP7idM1NHc1ZlLzl
MUuYE+Ya9EFcEUCXJuPZoZGaK73vRaXs+69OcJv6q0ogWDZ2OuO9L1GVVjsWJHK2
MYgB7bfJrgXbXwOdaL17/R6aqrRrrxXWHAB9v1QbDP0P8J11VxY2RaurFzw1q5wn
shbBFzPTQvsfSjduGpkJ1hIPFuqvgRYRu6PihUS64FthC1+UG/a+fHzl0XivlKCA
w1210BHIfANI1Wq2SQBFW92XF/onNDXrVA10Ov6Jj45n+BHZY3MySKeCLjzoaSfn
D7sa25j3txLbhJkOjtxN+wH2718qtS9OjYxRITwnwyKj35ccFOrT9FzfPtUdDg3O
wGOzapcoleH+WGXR/isaSWIiAeohHeOPqVdiXFWTkKdDGnHybGt+dQSkA+Mo80UT
7fsPL1aoVlmAc3Re3D8FASGR/y1jKy4PpEO8q8+e06neHg5GRhjyfvvwtPsQ7J5g
7RnGHMQK+nAed9Ut52A1hOJ7DD84qMqcZHYJpO84z3XbqtsCjGK3pmXvsMUsY8Se
ut1rp/oXH2oNAzhlueMwqHBa62RJ3u3Ff5DFDjoo29ar6qS0AGmO7b/jTYtP1dIW
7Cw/uqq1JbezXcAFt1DZpMvv1dUEWV9AlPqipMRzz1f3ULQrABwwQ7GxE6YGyuGB
iIosEWQnsF8PBc+++81KMRHvFOeoBAnBUzrxaHBYTpaHDc+O1QoDjzRkzGK87FDG
K+VEcKwAn5k1fw1zaSVo2JN9D9ldMd9NutrR3NMObsz1MIc1DV5iurtV21J4w0vm
SBs10snzNUDFXcSf7CQ/iE4Ko7gvsHPIUFd12PgZWvk1Zey9dnOU7T1wa9NlsOF+
2G0EQgNN7IAPjEAvK2kGHNFiq1zbEDCLzhXUomFCpA9NmF70kJThxUK6+vnq3Hls
OUYj+B2JZILwzK+RJ/lk1TqRq2DSmBDaa6I3eyJsvcLi0p2l5HCErCUmfNEb/rSo
9XknjoN/6OIn/Eld8sOPfdgrAPdv5Nf3QApVXbpLSW9TUt6b8Qd3zVvsbwn2Vxrl
I2b8s1Zb9I22qd86J8czwQUKnxP/3A4q4b3cPXa2yLLz+jiPj4TJgvsZBMg23bY3
7TOlLsfFAdnavvImrtXf2bSpNh9Kw7rbmvH6w5DohOYlfBu9eR31M7ziZHSxPP4S
2YkcwYnEBJKta4IQ/BTuCjMEWRkTjeia2d8HH5j/GHw6K2K9l0eyru38dG3RkVYV
fz4KNv/HCBnP8ilwTdIRs+I/E4zyJyulaMzj35EivlQxCO+bsonBNZEeFMukM2Ut
MZ2lJzcAJ24ubXwh9L+hb4bEbT3ERQUBUU5rGmSYbAKa88Rg4ZR4ssy+Aq62NpDh
9gpMHHCXbTkRfC8oZtxZ6YlehD+aimtIyOSLijkE9IxlWu7xtqeJr/H9TIfpHjt+
u7FaE/zdQ0cE++FJuacj+XQW6el5MXkO2gKQ80rIcMsl7PeKm3sMxS+vCltT841B
tvosHrRcn6H5visYxlGqe8HJdDOSOsrOfQTwASY/ZFrFYJZnXYOpETVFMuFPOQLD
053xYf0A/NV6otp8uWlIeB3alHRteXDIWeQPfQ1noT64L+TwAwSlCRNZVZt7usNO
rtGTLVkk+AK+Rbwb4o6usYSQlrqk1YFyja+3zTY51/ndUFYts7NLoT+ehETNshtb
4ic7wDst2Hke7+eVl7wMSlZQxua3j7f4BIdd+2B+zAFRhiZqVnuQji5hK5DLOCmC
PQM9vg1aJHBxh3LlVj8im8uwXKLDl9h7Y5TL+6RkBgE6rwe1kX1HVXZuJXDwujkx
slEssPq5o7+okhMZ+jTfUlI75WtroWksMQdj8wdlfSUVCJ78tgGwUV+arBtLvxYU
g0ten6BVA3v0QYu4IjHBHcDmeD7XvtW91VV8rrz/plc68c4Kw7gju73OTVBirYxy
yQgJ/ioexqm4Wkvw2xczEp9sJ6y9+BSdvYrMLjr/ktRHajYt5OqNYHfG5hq31oX5
cMmmjCJqeGqonap4b6+h5Hf6cTdqgIsKZBy37y+kX5lQRBCI0BObfqCfSyvYmNJb
zm/EWdUu4XjAqk6l8KaH4qT54DyqIixmZTufey7H+HnB3/Cbq8M1U/4NZMfM4pZX
0VEp4mYTgevIruAmL0cqRIq9Xsv6hzdfQdFKLQc/Pzjhcwc6GTwpeSL5+kX1KVQ4
FPdTuypp72Y8CLddHQ3rKAZTOc6FtdtKngJexd2dpWx9tsn2p1TVceHQ0kBMnzE5
cwzWQ9EuLS1BZf8vIlCdITp7sYCKiQcOlehhO5m37GDTC+ZsNaaJk8UMAOq9gfjT
N4rwvSrfnKKZNXHXE8D/oA==
`protect END_PROTECTED
