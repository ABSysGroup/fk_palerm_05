`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s6sIHEDXnzwckCia2hxBRq4L2oTUAiE3wCc7d6dNZ3XZNxkfNIWIYn9gVrAo8W7s
/5WMWyW6DgVIqsscSbk8klY+V0ZydLZvh2TvUMVHZ7c8PjZKG7VcWr5uZzohjUXr
Lm4UtV3KnlsmWF4ARUmU6yLmjxVtQ/i5RaxdRxp316iF/gteiVSqHzaaQOByLBQa
bo2fhJdhmaqLcfWn2Q+zyPzPSwFBYbJg7p6RFOdPfR4jjXXgIuppLfQtrP3s0wtJ
TxoL9Qzfwknv6DAY62esT5NjA7R+HHbAvc9rVE/caOoeAD1+5+gBnLNrxCMczlXM
hcuX1s37+Ah13SDkJR0rye8Arq9CHWiwEy8wgGGT/4Hblp+InagW45+7t9UC8bgz
7hwL0/q8rt8oNvXhQd3QWkGX2St6CuzVH6fhoENnC6W2roFRA5ydNz+2OJxhbSQx
dkN1lPOAhrS/HeCWD3MfKjfxi9dL8N7Gcw75RQYqEnU=
`protect END_PROTECTED
