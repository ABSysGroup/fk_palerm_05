`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LPiPaD9z49iP+XOSqPwL2GoItbkP49O0F81y6siRTMfXpK4w/ZivuiagrDT8Y94y
3KP2DRUhBdwDMl6wUJC4Ft5/U1GS1hctHRVxyzyxCcBbiw7ZZafLKmyfmnGP6VG6
M5Ai1Lq7VfITmzgZvAGRFkdtQZJiWl62ebZlM6HrsYDJj9YjyPsp8x4aL9MJDawv
WReHIP0Xcjvxnx/tHBDBjGbGJJbjnP2IlJzFJp6LObCt0gEjPyXxQ/8CGuvrGvkb
zvg8UEpWVGCzFbJFJt602FgDqSWOOlAzF1JghuXpRYWgWSIIG1mKPTq2SgeyjNnV
9+lE32OM2VV/FXq6P6rS1lAWMxpUkctoacW2me2eUYMacCI9ofObf5AgEkxDm/rr
0CWgtnJ8iLrzfBSQxsr/AzYjQ9JIL+auzQe8dO+Y2SB4ISS0IJ9+GYn+f5+4k74H
kdRxLA2ib+j0uPWQM9ZQekHwc4M9PkINIL6wfa5mF+oesyskpyD0VvpIAnIm0Ies
kZU856jTVXgoom6pLc32ET1va3zDj3YsOqTHGYWeihWh5Rog9SijnwPBYDlAlgwv
FteKPuXvVeKyc9IOLnB+WAget4xApiBhb7l4cZvQlay9YShURO/QDbj/wh5jnTBS
ZNVUP0+SxvHj3d9YFx2MDkKYDNitB/J0Op8fawCSlFz6Pdosu7JmzhAvGZq/tmcy
HslaaSXq/zRteMmXQgaN8phatRAJoRc9MvD2+onwaIOcxVjMfPQr6Wq+i3s3E3R+
Pq3IvphQITRtcjBKfgUubRJz8zujxf0boOtn1+RrZngm9J3Gv7+DG0xdaeY/AzkW
Kg0K8vt6grxPBBu7RrkKPPkawfz5PS6urIIdtDdhQIME8xB3jm9MzRwzcEm2swqR
ZgaKwsAy+VJEVfBatWjehSqguDySwoM2Kdwe5dMF95lS0kyZlGmlK3O+RZi9g1e5
/QBAtdCV25zmAnuKYExiIA==
`protect END_PROTECTED
