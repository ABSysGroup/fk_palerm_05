`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
beH0gzmMCEPiA2RW6mKlCuajGjL2XwFlN4EtW/QIUj1uqjBfv0T97mz28AgIrTjm
WFAX0pZfgTODJOmJxFSf5Bgehs9KDeZJPr88fn7J/pM1ZQL0JGRwl/jHqOhOTF1G
D48tq0KYxey1EDR36pq7q7P79JRdiQXYF76Q8lJ1Gcdj0yTAvrMH4HO/GkrfYLRd
wILgR1yLsANoARvfFjCevCsDZwhR53cTzhwmgRxZcJIbvBPBIn4HcdsH3hOUH9Ji
H7HnMOZ03gRyhoEQZcFYVUm2XDB6xpQIf+mirWyviLr4WsjLGnMaEVsgQXI821qr
jvOv/sB4Zt5+jv7TgNcID/BASzBMGDCOy7TV1yNAxwzyNOBXz5cv0BfDqZ7NYoRm
pA/oVcfkjCDLyYX32h+GVPG6/tfVO6xrH9ogBgHtCvZL4bU9pc1T6LQ964GwEMt4
1meAGfGwrH2o/4c5yWTfBDlXEURYD/GMEweVvip+4svs8f3vfqfEDkL0CQLF7FP5
PXTv1UjCSDbYkfrz82Y0YeWetAaP+3xpT0R2760vtZmYZ0m0nQqdO03+2FmH1XcV
xNEFSqfUAG4YjyZ4sOidhZ4IOn7tz4yrMF+2RdtNB1phppYwigfRcyLe+6SSzf9U
Fq5vrY7IAH5ygdFyw84PMxpDIPyQPbC3vTr1kRmp/7EK+zQtNBIJEdudnXQBOy0Q
VFvkiwfKRQWBxAQcgAN4KipgGnsPnoqcVEdJWXWWHsVL+MOQC6rpbtpBGb52v9W8
QzxfrD7L+VynuYlrv6iMXPtc5dSLefF6yt/XlgiGQyD1pO25bEst2m9i7i2DpYsw
LfBPCbxDvSUguXrAUUTzQfA/3tuIs0JdLriYpKw4yydwtbyBEPc4L3kMQX25BVDf
i9NiqP1cLvY1YWTwovHB0+vJuCf/7SP34nVcI3WFv0XHPnNF57PD0o2uNp7adneZ
hcRuSReYqvAbstKjsHNIdLTF8aKq1fh+cRKJZq8k430lN5Cv7VLob+2u9g+El64q
op2qyQkf8bDZHm36y1O0OIJ3+E72G6NyuwizyNDUZ4g1c+r3RrmHsNrWiBjLMqMH
Wo3r/Y0mLBO5O+pJklP7sYqbhNxMtPE/bEDzvpKfxd8YhldqGoAbc5O9J7vbKRnG
GUaNxGuoPUHUE7WPNm0DoQ==
`protect END_PROTECTED
