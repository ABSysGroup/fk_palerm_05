`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UaKeN5YDfNJgSVwo/909d0RZX3Rn/YjDAk3nqMpkaJ5/veGm0cL2E4GZ1jMK5pfM
NhNql6SFPYr9NBhNa3MmnzBqTymdBZ0+mO5zPJeZxUFV+10dljuRZqynucMe1cM4
7KDTnk4fmAe4FNJj7wz8hRg3fkCWJjdmtSC9Mt+IFNrq+gT0OcCkEAny8g5sv615
4hK7bYuY+/ESQWIH3/4W9/J24mEynsyfNTrO0CySZMDLSkmb9wDK8oskiKLb/OMc
+Sz+Co6gr4ruYUHulsrgOKYTD88993C0zthkN4lMLbgIP1BVvClViDh7CQ3hd8gR
ZOQUITv5l0mmEP9lu03vIwbAyhCVtfzaF0+UoWFStvrZaVceD07h7mRQuXeIzsAQ
y9Pyvk88GNxy54l/HNVMTggGK7pIYZibZYWzO1cWktM8D3KpaDWlB4ANZF12lkUY
EYYpmO+LIYjrfljldceLqBKlY0Em2D1CO+eOkH+bpkpO/fySg/5ku4oFmcn+tnbN
58hLyo4PczV3JCxpuDbSloeLl97iZ+pw03N1jr8x/4c=
`protect END_PROTECTED
