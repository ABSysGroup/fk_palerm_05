`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RmCHhQic1jY9uYDo4Nj7M61QMoLFCn7ZGz9REq1a+z9epMg92xGt1KxPrtqbTK2S
MrSAHAqs5foBG2WNv+jh0/bwnwKCdcrFw/rUFySNVUsCf3HJSPcGcrbTwLLpSjvS
TV3xqOgAWhNokedCA6DVEpsnQ4v7t7o2QTySDCQJ+bpuqWTC3jtQ3B+lLEb/FPTR
IR3zqu16DNKC4Ri6g/Th5za0hkRKHJJ4qY+kfGMxJxDqVVEKB2l/69MgccsGWhlX
w64c3j443uFrmXqCdfQOrA==
`protect END_PROTECTED
