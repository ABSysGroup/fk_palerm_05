`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bJoDBHGL3Ljm/SViARGFzKyoKO9hq215liNu7Sm83b25LrR32U0Tu0khtghOeTgz
3o9PjB3+qx0Qp/SZhl8aHD1Sat+NHe25F6ypRDywY2o8KRCy1QYfV+c7bcFzT8pc
z9315iprKEmUy1/GeypdVqT4fmcfhHVPCRKuMYnCOtoeqHpT4+dubmmyjeGgfrnE
0P3tWulGkrhWx4CrRBGEHqGpR6CNu2QzznFZV012I4CFV+m0k5cL57Ew2RSvIrVJ
ibti+c5avvWXDdCCke3L2T0aCHQDa4ESSZDHsLSpCpUpHSwFXMsBnlnX+2umGGjs
JFt6zrDBqk1GZxufCg960AxVcz9akqy5xT+n4bR9sCiTqmYnO5YtZGt6n7hkjTW9
0acPMXmxEtexNHTFwxYxBlYhv1+rl8nsUWbC9WQ4WgVDLbVHtp674cjrJXw+lhSo
jQNGJHS4Ewb8+GvH9ImftSo2uq09zwhDNvaiIyMYCUUQLpvdkdlXR1Kb+FisbHZ2
UqeQx7862VQJFfqB7Qvvor3GvF0vkIy5yG+O92r/5HVge4pM1PH1kxdB1U9vreYS
a0X9MPGomdMpDEYKQLUL1w==
`protect END_PROTECTED
