`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QWGGFSw5eequjspk+tV3wiKqOhl0/e0CwgwnuGLplfIEgG98FuIRPaTcSeKA6agq
O/tb+8Wu7bn4Xainn3RWkxSURgfHcPTeTKJi+ONmUSJz2Fvm9JrX5a7X+U1bs4K7
sTwwUBOA7e5Et8n3lXkF8ufwaDlz6DtemqONZ5ZmdLZrlGbzZgbmjWltq0u+Oqf0
ooJbmlrnjVwLhZFERaHyKWSHdIPYzdkrLlTkRZMLH6ZkYwZd61R5M2c96I0h0/WZ
uzwaO3Y/C8oZAYMmge9FY9MEnJ7LS6X0wkPF4tOKItkVyhz++7dg9eJeRVgsLgzr
VDxu8692fTjeg3IxJM8BjAjgyie2nKEgxagu+ZK+deFf47uDf6br8mUcAhZHTkMi
l+mjSO/S3VzySlSykfPZjmyfqoNxMQOrVhNljDS1e+k7gysb8R7riqs71aHLPXX2
zojfeCKc83w2QS0+i8USbw==
`protect END_PROTECTED
