`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P0Q1gJfxFHxp9rmeFhHeB0KZQZDIO6mW3FfVhp13kSqmkaKKZJyQI/ML9p6aW7XA
/iA4/VpKqQHWXNJ2sk/8YYnWe23Qt5QqzPxWrW/2+rTlYbXSWEYKjntedla7ioeR
/3mZaI67iS+zVf0jEdb5EVn1zIuG3/68+UNPkHZTpgo92RcOU0MYuLyENmSf+CZ7
4kkuo0BjmTFcECq8tqeJcFKDVnRikfpaXXwxOroTZMYq8hwj5AMhaDUl8BCzqm3G
25zpIrdo7ku1GxEalv2rU0dIowTPkpm73eGBj+YvmHmwa+IUZXv4fz3HAzgot5d5
KHYzd6H0L47indz0oR3SjLHVRd1iXJ1afF6T8A1CMlJoJGsHVG2cNxpw3vUplTUb
nWgXOGAJ3mCDfO4BSvEE8khuzAkDIQn9EDpphlvjAgz1bzCEkqmqkG66cBPnlnU2
hU2JE8nl8qpuQLcjDsZL2xHUFcLXS7/kwHrc3S/wtU6cxWI7jcIDIM9RfAM8FyXs
qM0YhUtGXOX43weNsSp5kgHzVZT/2QWB/iW8CMyvkplnr9B3ZpSiiDsf8J8USwBK
CDS0+rWfS1/dGAQhfauLGn4B1I5Z8OG0E3lCiGVx/YTW9QJvPnfrC0kRVxxoCTRi
S3J2RqAytUdqzpYT78t89CP/3FMjwWRc2GV/jmYUhjTPhzoEw/kBDCV1SUFfS4kd
oNgfvBQbXxo+CYogphOJMBuj3Q9lZDinIn9AK6dmxFQ=
`protect END_PROTECTED
