`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GRa9ycwJRTy30Hvz/eyvvn+YoRGuy02uxzxLpa5+TOXDBTFSe7XFgggQdCZKES3o
CxVhyYgL4ltI6uHfKRwCd0gybelLLtyM8o16JITdGb8FpyILLxBejq3CXG7erJkN
6+P8jsAY+CstUeSNapU6BrsXlOyxdbx3YDJZuVvEeMn1cECWckPli0rOofbjy0TQ
t1flg93ElhhQ6t0DCamI+5Hv5xwTHr+HsZk8irN95YCzRcAoUN3IaehO5VnsTt7p
K2+iWlsAOgMokhVEWx/5fmLjcJ1+9u0LlB1bnL0/fcfYF40e4twmTByHvc6bt9ru
8kAYmF0GwpiBDc5FFfSoU3FMDelfypcZfs86bsp+d7LZhQOaPJ14ZoTIoD9qv6LL
fFc3gICWeGsHAipZU2UWz2DfCTIt6x5EoJ8lbIW9WQY21niPq+l1rh6MDL6aDt6h
TbHikLoOE1skK3UBPchF3sbi3VH9fXyTxqwP/FbwYNclVJZvDIwygWoVKDqUP7QR
LQ/cPHj4DltpNU79GT/x6WUvtvW57ca1N78xu24KIZHz/KMWcCjO/jD0bFmeh4Bh
C1CZQ/bg/WzC+kVIz/eSp8T7lPJYh5eELTT5h/2tQPPtsLlxA5K6q/URlphUAsRL
yl5+iv7kF1PS+rietxqde6kTxNT7dbrTOUSlxwzs8gimgeOfe3d3C4ygl7v00SQp
9KDI1S6YB1S65RL1SJU9NXN68Iv7ee8IyscofNEcM7uD1ghC75Zqf+txS52jMc5t
GAR984SyGgmpMxrtrhcNEApV1PdeFH2/nQx5gr65viWBBWxIsFfC8eayi2F6OIGn
dUoZCHiWgrhBXZbJRoAKxcZ56AqWQM3S+sobpe502QQBCZpC59bnUMkgabBYBwP3
WyGu7Y3COQkHxxrJiumnvdGSxIzH3tWcNwokdCcxAHma3VcfhVnwt9nnDF2H11ut
C50+pBSedmmDg9MIw86P6YJJ5PLSxyJfzuFJgqTJSqo=
`protect END_PROTECTED
