`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BnY54E9SWSNgA7+TDmiYPS5QHVbzmMe8r7k5Sqq0y5lDCu7O5I1ZLCqG1ThUkNsK
IZTuFQMydGPxfm3BH1JZS1E60WyuaIvEJ35zRsxtaMBEYrLE1r2bfnISPSlHSslX
Tlpbnwl9cTJLgUGTRymXdAmB3TFWXuPXkfhO341vQxMHYKMLDlVpT+6Zrms/wO3X
2h2eebYzQIHoDWcYOKtPzkEbqIUGLV1XcjqRV6TnI7+ZPWfYBD13hPuyl5uVSPE0
U1KDfyHukYUNAO1J66h80PILAoUr8tjJL87ORTto3H+0CksWoxU8Xzask+mit0zs
aq/X/XKu9hCV+ja0BFjiqT6B172begeMNiDhha0qnD2mFkRhJMAE8HA/7897mR5k
g/jzvy566o+R6jN4RK1Ju6OFXGPs4bt7Rw2bRBhkhKMQP10GMJ6TTqB0UI6r30TC
3ztmGrcbWkrU7XsEjeQidJ/RLwS/8ELYo+LCP0jTAkq/Gd1qQKW0XgLJ+juSvNsF
h8hiLRt8cKzmJ8dg4mIEyxYlEo1upBeyJmStFa8rDa47Z3aIiurBP39vYtEQbuPe
S5MYl+17R4MLgciGv4mCkksICFebiqC9jLFPyjDO6zoVBQFqDAyDIK0CMTVtbDe6
QBbr6aV9zLVe5DIXQ9Pw7NbvDtGoLupj/QYBEluNxg/WFRv7EzAyc3NfbCkl+wf3
AwcVA2MINycCIEFHMPmfzld24q6ORUpXwjFfSeqj4FDHuFzAI7A725P/x1VMNpPd
K3LdLZeNffy28gmD3wbi0gv5qPLsrABUKPewzzT0I9WLJnB+ppxDvKbNxfTfCCtS
Fvbc+x0tqJ98XlYGTfGdoU6HheotIDJ1IBpH4ktwEpDPlZlOsRuJHKIqNLBBCuko
qNznieNYRDkVd7nBPH9dNUML56x8R6cw8T93I2PCE6O6oKbQSzueAD1GO+YUoSUe
4nwZOJ22tcPXOiO7iRoV4jmcI2aiCijZiMuHwnwhNGRmO0WNbIsUZDBjO9M1nnDF
xlNbfYZDrmiJMsb/yUnobVtqvH693YfMSr9Jbq5aYkI=
`protect END_PROTECTED
