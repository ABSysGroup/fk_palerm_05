`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XYeyvjsbfIBrCm038aPyJJ7OhAY5hxkT8a9OX6u5/J0S7uzo2pC1IRM8miEwft8t
YS13v6ZtTM4v4n+tL7lR1mqNWieD4H7ZK7Dczbka89hGx84DItO1x10OdPHKrKDU
9FVDuueWXwjnvkY5N3i4AxKdQ4G7+KrvOUCcL4COnXeOb08G8X5sb5rFDWrzboeE
a9VLtl861voi01S6Sy+uzFsCUDidvruZupJIdIdoDNRJHk4M2JZxcn9XtDvLw9Do
k5333jl3WGbnvGj9tek2VCHZ/AKcJ9iFcSNMwuAuFhpTpxKeB7UE9f+l6q+2BkW8
vFhfuGy0jzw00j/0Ai+qMDac3ZqB6chfSeY9uxAtl8ZclvxtJaG/vrGB5TcMhkre
ob5VEmNNjWTtzatfDCtNy5bbqS89FyQCjpqzOYQ3l90fadTUAa1VF7AHM7X6DKBo
1ZwvBxWR2ULXC7LWWH5YiNZk5K1GJ/tKLAUixCVnZfOmLm0IW9+GfvdcyAu41Sul
`protect END_PROTECTED
