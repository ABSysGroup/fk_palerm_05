`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dUM8rgc0RXvYzg8uuKH9TqAc98Ozqtb57RO8VU199mghKEhUxMCmeWMNEyd4etVV
YWHoszsXmnLC1XgNuU8es+WpPCMknXDLboLOQ8libTV2FbyTJUUT50DldTO4rRD6
2jxj7n5PPngqP6aeeuuK+CQE8wTbbHfrShDeJSRzBy/ba8N7gLd1s3/YRvm2CJd2
BhIy6DJjYYtpkEzGNEc3E3f1cY3Hrb6ZCl7ySO3rodSkc6yI5rBz5mmrEAF7Z6IL
0nrBLV1cgVhqg+tWt6Io4gIHpotw2Z36afsdlMrefnUhVU33D1aasSj9BTZRYNON
jhp8mR9cr6ysipO7i7xPRHcbfSXL7dUlA+FHJ9/4gnucrIClbC+mk3W54HkN8sWL
wOIDkz9xcJZPRiwQhtbFviZrlRXGsYKtIaqy2SbAYxfDUSKulrb6ytw5MMSUfVTj
lXJzCklDcMzJ4inyixdsJWUUDv3vvlSIbDP1tgKLLyOUaT8vDM1VB6c27X73aZGp
GlEdpcd1hJJyzZX4o33BBS4iCzCt05ip3o6HtbSogiUJLC5hdaZqDkHAGB9U7XlH
Bdlx3aNjFeATyr6nwZILerKmBOrxJHHMent08H30aGH/DJG4z92AQJJpGJl3dXKy
8HGIakEJ5pmPOuXPoNp7niPnAe3wsauZ6OC+pwPqhVJcClXWpzRbVpdm3Mopveil
Vk3QjyJcLLXysYWyEOBJqMDchNnZIiLgg2NuUssOFVX6ElV7F62XHOMdETZRXXmI
1sQP/8mdlhSySFPTPzb5zMDW98H0d/+i6exxTHN895f2e6+pXNyC83AqLu5rDh5U
WxN50JRIrEgyzLiwNSx2UraXhTFTwQXpq27Z7lIzQw6T0s6ZUwCnVfn863jhYUV/
wiXyYCqcsIv3exLvZmSG68ARDjslh21QlWfTROoS1cnVvb6bbXWLY7Ve9eATBxFW
mppT4j5zLJvJ+eCVrM6k0VxnpmsiKzJgaBqcGroN35p/dsPlWHqgWq4howhRHmwn
4Q0labrdwx7UY+rJv/liYEvuxykFd3gj0/pAzvRb6pzQ2SpT0RTBaIa7uPR5TvYl
VnO7lir4JRJb0O4KC0upG9Ped4Swpl9i5TTHfP2gkuIAXDB0v5aUpp3IOCnqA0QO
7Fpk5jmj5VKvJ3JsmxZuDtXV9rNmtMMizCHdPkkIPFDSkkMZVZXhkLxRsdXCkB4t
AnSatZ2y6pGxOsXpmVftoNuBkLkyB8mS4bEZA0IdYeWFhRYInfkQuCwfL4kttXag
vCU8L7WBWNlDnDV398Xsxp8JrfrC+FGpB7BfsJjsrTntFZKSYn0tIkBnQTKxQk9G
FGajGpI4FZ39u5Ji8GRwNlGT/knNa5pXLo0N3Z+3iWV2XEns0lwSxTOA7y/1PPtc
LqF0aCWznTfRvWcfUSbpRRDiHPi7jj+/jOcDOlwMlRM=
`protect END_PROTECTED
