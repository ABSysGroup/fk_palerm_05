`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6jQWj89k3K8TcoLqnvrD65ruinBJitvkcKDCkk02pAdXAIsMTHBW7CV0gUoc0JGX
BXnPSWJYwQiUxwYuA+p198T/wmivfzy03srCT0753qiSn81njj/q+vfTIdwDosew
tqsdxtP7fau697ARxJW32WPSO3JvULPzWORA3DWsnlZuLbxjNmZSfBC67NY7kO1v
lZsArA8bw2c6foZRtb6X/gxCdrUag9dWB4dgTF/Ouoq9ay5PTMSBmdlDAUOJFEFf
BPxjji7OslwQ4h0XyUNRo6bvkf35/IM+Q1xzV+3R0Dj9Cbko+MLyRPWPswquBx8J
AjGUQ5J6agPIg/xJ7tmMdG4qTejh5ZohYVJxi6tbjvnEVOd+aqwN5QORZmn9hAtz
BqtYRmFG3sjXBkrvrJQBnJkYEQ5XMa/nGUlasjj7epKdtQzaO2aHMhonfbWFEWAN
goSfhKUlsJQjhjmUkGcr5TGulpTXe1tFQsqNgAmvCM9IwPK0LAhxMw5Db6k/EaX9
QgM0hf15wW0ceTW+UUHhuci+or1e1sP9VzFR58bp/ejsyuTQ6Jq6qa6jvg6ppaeG
OxA7HdFCEV9tiAdNltyh6HREJEVDsphxwxOdU2DBalIk/40DrtK7C0dB9YVVLCks
Qv2N+tohZ4DhwvlEGLIcVH58lbUoFc+vVd9LT4+DI+JcoRUdwAqGmxQs/tihpGaM
nfAN4jbCcffFT+pCWrt+SG28bCkbcbJHRu10+ygLj/Je0FKtyRI3sYW+marCwvyh
R4p86Yvt13edkiUHWgzBu5d9HkxOTDjDhA8vDXpydj9/3s4V/b4ylWXlzFW5PDao
S8j6WsZSK0Q8acZQP+Ooz/B53BNTxuH2Ivft0h3tJabI4ERTqc4GjjR9Zs1UhbqA
sktx095OEindnGoOVtWAq7/9GkQQwk0P7UoI8GjY6GyU+bEZ57e5+pRFZg/M6gB0
H5V8SXNtlnz1XYMx4FfN8Z/p98sybVQ2XyOuj6RoIn+qYA44QqgS1w/4gmNt9Jv7
JV/qABI1q1PNBemWIPynNe5ppWVhBHjoifsW8Bk+nmA31H3eXmz6//+Dpzl32Hxy
YTWKhJ1yYpiPViduGyyV9kRqoBcAmBP5nhSoe+eGZ4WYDmgD/VTC+to86XsCqknS
bTHrlWQHMISKl0KqheJNJ2Q3yXKtjaaytmkGkNJ6tDswLcxal/MllPjp+YXQCLOF
DQG3x8ognLLuVSx7qC7q7zyVVSwgbBjlZQpiYn4+neFQi16g5sxVk4ZHE4Nl4RCx
GJAdqQQIiJ9PV3bUK4QnppJuv5BWcg9Jn6/no+oJ3QfhP9/mCevWA5wC2L0MUXHg
QA2BLOPfxZbttrd+lLPsorsM/jbY6fsL1aRjUArGdjWkfctKxQi3fCWFipiMbaiA
GnO6eB+XoX9plswFeoisGmpeAJ8jGqdyUlaY5qYrMjhvU3JIyHtkkifPWrldVqc5
fWE8Begu8qdz+BwWIyQ6mP/TPnNHThVv6wYBd10bY5JGpmw0yvY2IEU4K7Zb1DWG
OKRjc1wdxr2f4CID9LVGn1GHC8wsCiCdVoaA3qjk4jbk8qCYopho0TUbZpSvIWS1
vCguNjKemikmGsuEOLQmlxQ9lNGqGq0TS79wN4vL+NyxyOaNYVDvUOclaKl7DDnW
FCWCCgDtzONhbceNvoCDYEaI5f/UgyXqpsRI6vBmngfIrN/X4wG0JBL/Ceb2JfHl
soLZVfXN4IgyjQvu95CNFtpmWT7lU8VttnhiSkOlPGqplSbepnKhUGv6PpHCUFhm
gwuYOQxRGMMMOEjEMNXsUAcArj7Om7kMQHOfOdJ3Pkk4Aa/2XtpyzT8wWjvIGgbX
/wEjIjRsWxloBdjq5bR7qwOctiPDDIzcROve2wO2UaVLG5KpeIteaQgYMbO5D+OR
/+sv8nlcrmQ8aPKcrNRFjSgOXC12I4zzVcxBD9qG/e+FVHQhEAFNZ6yD9jWYe6GA
m1SbEWdygVUxXReIEFlZOzk5322vV165WMVRRXl9nayQr7q2QbX6TCEnzUWkXWzs
i9sZE3k3Ej24Y8naRQ/yphjJu34yuf/VETujl1TxeLuK7d6ME6CJo/R+u8i3awsb
SP7PYomRcIzQ+Nwpa4Jx9SGqKtlp+AxUbyMkSUIaHBymssOwFXKTXorkzr3J/p1S
QwAqleuBxpfdMvQnnEkfkY9wUO3Ou0RCGEUTxKMo8AKZd+M5bOTEU+rKUkcc6aJq
7y564aBL8tQzMyLbYH1pr1be17YaX2gbv0w2IPatMU2AZEsJERByATY11eGpr+oi
VwceiVW/Qo3Kt84g6mLVpfW/KKLdoTP3F4glNsAe0Uafr42EKKSoPSCQ5GjB2uKF
VbRfe0QkvHfixTZoqbb35LA8Yn3gXtPIx/TlzEs82cJJ2czsnpoxbr+KULY4CcgH
1Oj9CR2QkoV4By0A96uWzE3Vn6xp3yjVP3+u9VYs+6iiXuouLo9KcOnlrOBK3205
V2D+grJzH7ewM/SWSlFRJ9FNHeCLipsHw/K7/JSHxxRiBTt8FjtnSpN83qFM3Lf2
Mh4RAxyLb691uWxJrs00D/KCeY4QWuUcqJtHoHepryWU5MY7EIL6++vF86fbDFgE
OrLrWDmZV7LEmQrEY0MwaZIwSv1aCoky7qHEf+Is2HEWEP3Ryf8EIu9dcV6KtP1H
ACAV49Jfb0Rg/y1PMEWSEA==
`protect END_PROTECTED
