`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HyeOWoIOyDQhBIlb/qOlbZCgOdtRWRHicudi2vF+4foJLLrd7O98c2+VGG60HHTS
mYbE6s8fe6CXpKn8+HW+8348rSrjAUWq3ldQkozMmU5ckyTmGm287vh29pjT7mQz
H8DuYbe+Zzw5Mq3kk/ZVMrhh5FdzAk3NpJyNLifXiRpSrFrJo+QljMxC8INCqUNA
SKJEqGd7zmb6qq0tPbyxrmK8Q64Ot94q56jHMr0I0Wu09o3dpFC8YFk4Kosl65+S
xqT0bFYMGYXge+H/nYt1MmqTb/wdj0KWOrMIF1fMNoVK8TkTQkbdiGmZf+r2r/x/
iAOjhNLI4zwUaUi4qVI3ZaQjPU54nEyldSF+ELvN6WkbPh2dA1HUI7Ib9Ycy/Bh/
1pRA9wOPkjbacGrJz1g+jsjgfvxtyxEZ3p5Z9Y57RG9IXDQUqNQv8tUlYP6Wh6dz
ARQHiWsU/yYyUIDTpzACtjdIekWrV2fEQID0Ueum8XXgMAPx37quhehvfTo46/zZ
nbOBzSQ/SXJRDUXAjihXvUkw4UK9xZEvy+naLjuHx9l4vv17ohL1eaAZBxcZ2yD2
TVnS2bNRWWgJfzXJn7WOKxBjRUq6irFbY2kAiFoEr9IHm4PyS8PBuiytpUXmSln6
eWBM/JQ6RpBw7Uqa2Ua61Egy349QYWzccMw+9X82lYBXzQ2Bl9qXaj0w5BQ2GwAm
QRJFRZH+ibw8mNRxtAOYO/xglTgTilb+KaHh+zfMgv1nyJ831YSCONPZTjZUCwy7
7N7cTDK17MuD1pQW+rX+BYEUiQqqf7OzlI5JRL8Bsjr+4F8Pt3ylfN8ZihhNWGss
970tswV8C3gVcyBlHGTflj2QKe4O+Rug/yzEPwpoo/Xh4Exae/QBhw+6EJepihtw
`protect END_PROTECTED
