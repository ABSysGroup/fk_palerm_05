`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x+KniTw/FOTksiJBbGCF2OYQaz2bqXwh5wBJlexNpLuOYy6YJz2JFw4r0Ic55zIY
KI7pW9fBgWuyEaF9c3gw51gTFAMg+BUGNhHQ5Kw678vZ/v4C+kxAEte4hx1b7lPA
iNCWi2UDgCMFPSZKkI9HkN5urnHP2J2vgU/vq17AwXhkPrLI3nEmIDh5SF90h0Is
/wbDYJWMQO16/YRyOWG01Lpbo8HF0Y4Ur0bXuvR8yqQmviIPaetUuTV05Mqq4y1S
CgvGvfk5D2f7gKAEMcrus7wwGWPteRk/MROl1+eUdEXVYscaddA9V5oNjPBtda1r
vwCbYDUjf84T22oMnThylgIZdY4xOZrA9B5LQlbc1jduyQLkgNHcVzsY+Jyzp9ko
Vf08UTxgIIhc2QO3pa+PI5dBFlm49+E5rBipcQ566pJZU+HYepBXEpT2e51TIQua
J4N/X4mSx7iuHv1RTEzaS4y0KQyt3W/mnfdiplSufkFb+OPTDsKmWSDDOxiNg8SB
8N57FRXaR+NbGDQ0qrPWBU3NI4eyOmkowgZaK4JucaVcJQgoKWjsPWF3vA5f4bij
+M4ipRZ+TGSUIX8twr0H2lKEY133US/+dK+N2zJ/AZA=
`protect END_PROTECTED
