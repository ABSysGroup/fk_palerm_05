`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vf8In4/JKQohtV6akqauCv57W6AvEuElKMPAGWKFYHMAHjNtj8o6NnZHF/hQX/DJ
63GAmRf/ugiDVXQd5I+HMnqFJzopxSzfPHgCJmk5GTYbpul4kn3rp79tS1dkinFC
rzlQeUDEJkt30YjiuVB8E1MK32mz99unJrXAB8KLL9a0fTnEh/rcb4ZaHeDw/cdJ
/PkbPg54snE4s2L7w6OM8bICvFF0/9mx7hOQ0podB7R6WDMxZ4Rvfz57gQzseE6p
WWqFWVOByVQ2NJwRJ5a7tm4EGpUh0hNA4yXRWyv5bea8HJEa/YGmdZZ+OQxK/ahv
eeRj21PfLO1Q+BFwwLWodEGS4wI4A1Py/aPOSRutwpubVt6U1X9XG3gI2swdBH7V
0UxB3v+8TNysdDXExsQcamyq5/cGL55pcnWRu57XXrP6XBfh03SVMuHV+cJJVr1R
3fslDYovfpKINFHcJdVE0JRDdpiVTPaTx9mjq/qMSfFIOPXyNrLkeETjORnOrqv9
by7sPf0tQIdi2HtIQQ/PqSuLbO+sJXb2yVQ5gWvRyqjAcSa0golDwPUU7hxPa5QB
XHVmhSYOUh4htr+YK0jvwaPPV2JjgZboHoS2QxdS1vuMgGUYhwTQTgImuD4EgBUm
uq+8bSs88svLGBC96O63NQ==
`protect END_PROTECTED
