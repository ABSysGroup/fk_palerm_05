`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BVUtaxyVzPavbKnHrl7KxHeSeLozrOUT1h6Z5AFV+CY3RSwZllogjTgwH7baEopS
iiDz5ntsg+c4UGJ2oq/B+XWtE3BJSL/7g/8ERJR+17tMa6P4FfySFQahReOPj3Dp
RA53V0JM4psIS/ZBeYMStKmDOxXZAyVhCIRdpapaVy5ZhpkfOrT6CRDH0wDRuM6n
4nCRUjSYpK/wiESVhoHwd+5mQ+Z4vag6EbygyVLqEMLv3e/JKqozDv5BC1CC/HVD
MEjp6Z9AWYOB9qayHEaSRhHyaYgl7GvLXOWkmM7ZQ5L7+sKDw8YFLFN6TUw23tHJ
YDnyhBBQaPuQY/j+9H/NueOh/ifz+eY6QNOn/weJPgh6jTNkpXGqZjNXsq551dYS
y/WmvuhM6haMp7gLEQIL4paO5JgteRs7K9Hp4ttRQeEM4fet38Tk688X/0+RqYtt
oZs74Ig887bdLiexlt4xrz16KKY9rfM2GYSG8z0wDvHEIDEDSzoDILYoR+brsjVi
vganG381e1v3HK+SSbQiGHa9C+fu/+epSdM3s8xkw3pvKtcJoo/9qlLSLPZhLE9n
`protect END_PROTECTED
