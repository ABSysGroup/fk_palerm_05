`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lkv4VAyG44MTdxMWsmoB3IfAT1iKjHhQI4iE5XsQtRMmKI+/W6vFI2Tbq/MenDdq
3T2PVLuoeqdpyaoA2Euh2hwMgezaPMxH17al8/Tebqi0LJGTzj0RWU0Hk0J4qLaT
fbfgM0z8Wu+iC448nC0wmpxtGvtoa+1T3Ylm80oQS8WlC3uVu/ahfuVEttpcp/3u
gBzbZFvAyBgrzaWrjU04WlSxB3aVaqLzzCDzb+ht9Cz/1+f88kBDHLI4QzusRS/2
+fd2+mr7dca0ECwb9BBHAV+Ggwn4q+0d0xHBwkC80a34atG/NZmEf6T4X+4/ao4d
H/0t+qBdCe8lSpr/lKd27lEc2zsemyY2bUpv+hlqI2bPbubhL0RVweXsuF6ImXDI
5M3w3de+09RW3yjDsgE/8tKq6L3Tk/voMROluHr1JY78ihwG2peAWCdlEO9EwJQo
EAAmMmpoUREcyqoTFf9Cd3opbh+EnMybTnQkogawEdqNOYiqeuFqufASfDbzay1Z
QYe9laioGXOe1OZ61iHdGIY08+IuC7RbofVASGaI6gsX9420YpyvWxUnvqPy5MxI
rngpWj8XnZiqcbjDzYKaK7OcJgK+cQtPenFAB9IhSrqFgO99w0GJBhFtct2QVCMR
nBZz9iVMmQBS7HQzq2mpszTGuI2tAhGpOkq7KeQJBYwp5sDIKLbnxyShrjvW6X59
D/T2dhd6nhYanLCa1Iyr6XowRGcVluVaNAXfxwRvyQvquLrE0qedQ8RnxOZDcgy9
NSzJXEr9HgkH6tIcYxLfxCA/GDdtgWTBb6asl33prlMQ3TdQ9NYLg90dMbxb+gcB
/brQfvCH2B1HmCS72yMq9H7UPODbAhWEg4uOF1i/9O/K+YpfIIMb8XgwZglaTTt/
h0FNDGQTChFzrmS0MIjRyQl8EtMOGeTFMWe4dlRQvpWfhinzW1pZIH9kgijQsuXz
gU6z+cRGBdeZB+jO7l7jprzH3ms0JtG734T8NbhG5HVKcGSSwdFIrS4uPVABgeoN
UXOiLpXRTzk0Hfg8d5l74vruUt4CMzuXLb8X/c7/1l1sqwxKqLdgQfJbj1eO1CrZ
WfyuRJaTzfu2J/jxYbbeVMEn4ke5RFRAf/lTHsuYKviPpWLsz/dO7sbEXM6/CohZ
IWXrlvll3/uYzERRRV01Wed6mzAMBN+nXfFnjAABxIbjHngyMYsU7uFV6V8MMWyN
qkAtpLYNlurCWUBg8Y2Ap85OtfmABA41wmxLqGWUEuse5XWMlVbCfqQc77dzRGWU
qL7KXnmKUjBNJpzyH7S41m/PjvQqNyOrshk7b3FTXoGBZlMeXWRf4KUmagw7BI9b
oPZOLulU2lZMe69lfL3QNW0+mSYSDkLm7l9Ds0Vab3YldvtRYOJxwpPPvCIM0AgL
G3W0wCXVHkmFDrCS134F37wojfK0GzuCApEs+/MRHxBkxf6tw4hkidu1ZhM7QXbb
8sTLOXtyXuoEO69rlAOPoBPc5JdSCsHeFWPWdYGBfb8l36h8C4VaYzy1Xt0FGQ4d
eGl8RmmSQOgyAsZkrZxn4TXslpD9UHrXKGZ+5Mz1jd3TZAPDnQcvnJIhFMzME6Ej
+ZbK2JL8V0vifxG0K3yzFB67+Q9jwTRzSHQYXlFzdcCX/dpHTmsD+qoo3oYeGuC4
4xTCM94HwW4vkif02bkn0v1rc/nOxn7B9FsXwaqJzKkeOAozv6gv6ITfM+EAhb0C
XnvMm3VRWKnarg2jNzyma6+ZECfdf3bvK4SedjFu6iHCOTBap9LdwYg3rj2QQ19S
7TF8wvEkYp+uwBQkU6Qm4r/1ZCnWyzfQMaaJq1QrBcMyG6kQfLQAM41BIj4bq2wG
EdBqbmtc1VWV28NqAUDqfdAC9zQCPoAYgke7mP+IWu0ZexGPHRHbHSpEOINUwGam
vLxLgAPDdcM20Gus2RCENWn0Ib4/ZVAPIWbnK4qKjw/JsMkP8DGQOh+zAGyCnXiT
LCfkdgTZPpskPm/Q/sETkwrVMU6Xjfx7WLeZmN9BE7JFJv6C/urwga3ed1S1fz3G
fHL8+v/aVtTCsGW325Cu+YDiWf//0ZA647YfknGagXSDNbnu/2XhNU9bAtxH9Ruh
SX8c2xl1YdxHvjLsmKd9p26i9nFP8PT96t5WttlCxweD09sV7myunNS8iGVEtLsR
6vDrKPF6rE4FLVER6Aa/5hGIuTaPTiJEV3kCDFwQGmg/dwcJerc3A2MDQdAr9XnO
qquLFDeRBXHuNSFDrIEEdXJPkUeClgbs646L4arIdM7tfKb6y6YjQYZwe5ctlfHI
pSlaH+uHOOqRRkwN4zMJW+oni2dmgoexb3aWFvPIsfcKvidC0ShkHXAUd/+3lLHL
RDOEIB4+o4IR5KPqVRxj01ldUqUt6QuDKrVL4viKypXFgDvkua+Ffag+Cb1e3UYC
ACEcAXsbpsR3zjjDxAm/L0f8DBpPcSMDQZmQUpVaKr4xmXB4ovyvyl2HJdkA2UTY
kOPgZvFCCIaY+/WkWCUqE6N+sIO6nDrZUdX+s9nuyDMmhB1kRMI0lTHkoM0bu3fI
+ZpZIPxKj4vUZ+sEU/7tHEPGo4MyHoXsQaLLq79XgHuGv9hSSotI56gYXbMWkGcc
Y27nK0loQWO8VVH5hFvsidBzveqnHtp3SgP0MwUb4CSmM/0bEQGrKfCMnRH56NTk
UPb2eJebEXs++0dwXusIErAZ5lhVP23n6TN0WMX90uZ3aAhjZGtQNIs0ILdL7xwc
YNGI91pWnfc2IKEs7/AGoofUyS3915VoIxpUPKVj0CRLh2/f9I16MBsebvNHPi6r
XxLFbdjm0fYjIEsoCzEHyBd4NiT+cGUIETU19ZVwqY9zhXLiqbaYtTPcD+2h1faX
zBP4RnP85AoC7sPiAwQAeepGH5IFyhik7pqGBQ8yC6APKDZ4xEpXJCT/T5ZhE4UP
MwdFQjoaX9HK4K67WQ7IdShYRMYUwL/3v+HR1CEvC2gCPeS9YymffViLJ3aZZDIM
eCzZ2OiHT1o85TOT7GygWoQ7k6nQ497UREfErHncVOKahtU67k/7LqjwFN4WetZ1
8uJj+ROoNC1ClUdIRnYx6wJa6AMkk+PFHVWhDRPXcCmAe1zW7GwZ8HCMdugksOGA
MV7mi8Xk7tTfDBq6PDWwQrSkegcRNQPKeVZyIT1IKnEqhWSy0E7HRe99yGXgjUZZ
mbtk+8WlpdPFqYrNlkR4SpB5VBNB9olOONWuTs+GvnH2ts27VN1RJBgoTA5li4zT
kF+hPv8G4koWokteqrvCN+ar7RTTodh6DOJc+1J9cXnqu1yIYcW34XEg4SwJ9eJ/
ICoI0e5raqPUnApyLYfLkEjEFa78sFS7HnNFsRMFNZts1EylTPm2QV3cNRar7tdi
fFdMQQZYgJsi9zROyXTuv2ybBFJb8Y8eYmXC9at4RUL0PBBDpjXEqxLfGFt7C/rW
PA2ZwwNRLEwCi59NtUv46fzKMceWEmuwbnOnE/nEGWFnIUCpd/rTB770aRBFf1R3
sj8qHzKRLXJhdYEdIKIyQ3KFCDTH2fKNWeMizu+uXRQ5rlNBG51Igf9f5pQIlipE
hosMNMVnYnyxQdiZUTAtmStXz2E8KG5cSdTA1mO3lckvSerR+av9wXlkY1QwJLoJ
mnvRY3oqcQt2U4NX6owwuNZGKWIJ4GnAR99YkPb6wAdWc10kukXgPXKAU+s6nhk3
wnird6kc3rxOA/0tioV8bQNXx0zVVH/2wn0mfKh9ZmNSeWc0aVR1Rljps7BaXC8L
UCA+BuvBVqFVrGJV2pTzbM1g9GtzJSHa8JeSWOi8YbzOOWlHYESqlmrZnWMwybcU
FUiu3LrGSdvSbfSlUt0KfHX0z15pJDCG6sjc3AdTGfnl7uBb8MYhbECGG5q9WXOE
Jn/jgFtqnyp3pSY30DiD2kah9bQ8saundsQfFQqAaBSUexZhkBytwMQwJ62NW3YX
sBiC+WLXCSDN/AOTTPzCmzo/sQMb4lr5Eomd915krkAIKRIg6ORgG9Aaw1wiXRTb
lckf2ePLNgF3Ypluyv9Dac/D3sN/BxLk9WpD9Xt7s69Mft6VGke1AhZNTubyR0CU
S8g7mT1fOM+TrShHMom1xXmNp+KUzExW9n2R93vROHNCjJaf5HnWv7TI4cOsyaF+
qEUXTz4BiUzXpSAjAAK9V1KOwy0MggHZhjIZo7phVJx9arg3XXR7oEmm6I3/Zhrz
sP5nthnTAIwEqidj0VkygB9CryH+cVurtA1Cs/my6gYIvmFwuIg5r/WCVLEAVnJb
Tpw1pVztWYmI/qeab0EvkmyIdO6d3DFmcNA9FMM+vLTyj23O2XrX2mxVbRZ5+LER
JEyiKnrALRe/g9vHE3EEsPL3ZipE9RyHdrbDTJzpBOiB7Ubif8oGdZ9kNpHgBPyP
jDfw657aFfaIa62cphKDOkvLZ1UkSR1Sx4y7zZqB5JU=
`protect END_PROTECTED
