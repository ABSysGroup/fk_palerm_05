`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OoHlWTpKiP4RAJtzhalTc78qmVUPxEiarDJrpeDAlEB2tAF94EZIg9m3gSZX3zTQ
1iKUjPpzxeQsIWRNv1f6x6I0UjPV51Q0OX7mRE5DMpqwrXqRykNfFfuTLR7GKLiF
Hk/W6NEBC+lHSAeGdPe2Xv6FkukmE2FpYy6L0zAPmlUPpKjszV0n9dDVOOSrzpqE
lRaPa9Zc8X9nGKeEfSnzYVRlFlO36d2gR0FycWyhYJa0XJHTVCnimg/u6mzmLm9o
1cvzRMw+EVMiz5YGmLvPgnzj+ttqf5tJQF588Puyd7s1kct07OInV7bCk5j9eXGj
r5UbtmFW+Lgkl3SwH45RMiubpxPPRzUH0rZG3rX4ifXsBoTNKPxRtDSvDB7YdvQs
SCn4UDnZU7qjF7TrzalObLpvMSF28200+5yI2+KyJrx3HAAfOeEyTeK9SfQwKHjK
SlheNlrasaBdbhvHhZZ3KmUQrG+LkTxsjAurmLm4WG1PKW9r+JELtJ6XuxjGJgma
fmGkvT2ag0EGjBZB+VRzS+37caiqqF5Tk/7PvCV1rqvokOK6I3B2SGLfaFYJuFqO
QyQEgmflBDUlUb47I+OUnO+4ewNjqPTG4YnGvUlnvXWBfiQf2AgUKeUqGmtk4A+y
/2pLwGjd0euXc604Q1/hBjfYea/Kk/0Lc07wKld3KX8hVa6XT1RccPKFbyxrdENZ
e2eyC8WCYVGpF4MoZhDv9MYqKJulyN5w2eLzPiHmGqv+/ehAvp1CT29vy9n2ugRM
1sJgu8lVZ7x70N2FkvAObK/HtEnm0k9zybSDEtKHIaVLqz+Tbl+nSoO0C/ny+vIo
xrLkSsDKnkgnSvaEPP3SDdbmluWiqLkaq+BSylbep1+IJOi+csRhwwacBDCTR044
bKax6Pq/iJs/uqMI1NBM67Hs7ndcxFr2NGvwdvbIwRDSflkCohYBCdBFqLn4LG5Q
`protect END_PROTECTED
