`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tYWq8BCAkrdJWJ5G8+AfkXdFo9PtIu/TxdJhzNiqC0eLpl5MgpifbzyLUhrWQ+KL
2MbzQtDleuiuFo9BE76UtbV9WR+pEvizLsRlv1ANm2HFFcP8uelxG/cqLl67+Tmo
vji0oqiBcAk5vpkMwdabQBTpM9G72Xi8WVyVydiDvkhaZWohbcE/e+PuTMwRCH81
VI4U4niV/eA8O2UOdYMC5MgSkZHXVhYXS1txvu7nlpJtGaBrBuZonXCKKaGm+9Yo
35OoC+1nEhMCQq8ZTX8NVZFM0VFxzdfTJ7VfhTn3iN3mdt6LnV86VdLwEsLQjV2X
0Q39oniQqbAav1fEN6SfHPguo7SB/XB9zmHRgtP2uu70mVf6t0Devr6M+Gxggj2W
LeGg1yNHCPb7xmqPEQMRW1LI7LpbFJEw/knokXuRafLcr3hgRBaYwWIHsvTtULMl
6nX2H5WOTQ5POVkEX/zojSncB9qUzhx46Bi0RQukgV6KnLr240ZBAmGyTOIkqw07
WoveyCFiKOo6Jak6GvgEYFX5M6nN80CxeVtQwCCpKYzsLeQoy8Pomrd64EWrKg7Q
rHm+Q+zXbjNxSG9ebrRunf7v+Q8Aeufpt0iPADHcy5DuW8u7JUoNBW75iHHyjQAc
GA9z3EBinTaDeNxHuRYWxOtoiSWPLedcPhdHQ8Ak5en8Y4OnIKvvLiYwgNC9N37G
xgmd5tb2O1BiM6oUM1Ew5lk1mD7p/x7huW37ielsSaA8SazVCddYtZmwcKGpBasF
wF5CFbRvrd6fDzZlcNNtgNKQgyeioePu2bqzsL3Uc5sffp4DqNIzVmSryeJVJIa8
x5MUfhwRQMclqgJlvvQxGpIT+AEqNXmrieB5FO9JROVHVnCTT5UWYKkQ1O5LA3qJ
RulyXD25poJJeYsiRS1n3AUgwUoKZIkkGMxoaX8FhUIQjXzpPjzaLnFT0N35sM07
ffHaVc0fvGmJ+a8EBOuXHbi1fByekOcaDUvgVTdBh+Gb7PazBuR0HAICVSpbIC0o
/sdB5b0SIIVXMe8ra60ugjWCeENzbdMCWxE5G271wclSkjyTRvjdopKRnXjICDhF
CQVAh/p12V9PJB/d8eGSIGEAsr5oaeJ+fnYX4Cfkmp/YOvXIJYXv7Om5ukfb4KA9
UlaZA0gncJ9KM9oTCNSj/ukV+5VDOiwWOyCzZfTruN8cc5QaG3gfp/ULLyDAmGzj
qTouTLtMLrlpPEx/4r30I5WM+CTUL/9BI5fhZ5KjjMdWK82cdj0r4GAjCtYRNwDD
`protect END_PROTECTED
