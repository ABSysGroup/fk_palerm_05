`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uYIngdNF5FHosUT3QLoPKICyBjNiHTX7zW/NJ4rd1jePnEs871BcKppRT2KY9Y0c
FAytmlxqB00tE1kxIyruUTy+6umAaMYSXUxMCl3U/co7dThb1lG9jXb6MohUJdIo
w5A3sJURTasQH0+tq1yqV/xFKuwbMUElG2Qqfabiveu+mB5nTltr8hxr9CBaWVnh
0mgVkhDH61d2rd5e2+blAh28o2aAwjvmvY2b1EAFeFYKKN1Vmh3CUXOjGU1x2nFy
IJC/lV8P/gAr4+3D4iX3cKL3Fb+3Lh/sW9GnJY2UYKjb52J0mlQsW+sXrVKqaowM
AsPMM2g9gLCSghKShHWbmm3HuQ2JWoWpzhQbMMJ15Vb/CHURz0HW0iWpY2JQbnDw
3CLt9fBrej3uWZHBmrhy81M6lhmErMU6y9R6qaMg/cjNIvVggbvBWC68Dtiu6aYG
LweLtz/Mv1AH+r2FPqh4ynmNcaWXqRFh89tyg7l4rxOAIgsjSv+K3GV+v2uflwE1
dYL/e0pzgBjOvN5kLfh2hNscQJkjAeWxRx7S3yVNAs2VpRJLhjFj6rQTIart4pW0
4X5GIh01n2VMLvbGO3LWTXoGki9eVUbvIQ+BEhhWcqk=
`protect END_PROTECTED
