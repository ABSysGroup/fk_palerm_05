`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a1wPC9o4ShmxTfvmfOn/VUo6XzpnSjuNq1ZfhSYlEuoyVd7aE1zcNNm9sMQABFU5
J2G54ed/Wl4B9mSgoNYV/6aBWA5oMpwAQJa4Dm5AV598o0nIgGYdw+bmkNsgCAup
SPbDsGeYc/RiADtpWgRLi6PfHakpfk+cZrVkcdKRhgKLeWLMKQC3ucIWKOqX8u8H
cmpvde31VRG30hbIkuBAQFMDS13/q1vH3SbgzyPbi4xPvBqLKGUHzJ2UcZZ3JMWP
zbzXVd7b/miBggFN1amzVGotiYxa7bk3A+O0b4CJv5OtYgy4eRiAGtvF6mz4gMVU
5a/ZPzcjy33FUzHrKP7jiXMFqJiQ1FO5v9L9YpLc1JC0FP20jHfK+hco9sGuYCrc
6ctLuwYHmwHJTJlwyAlbvPQaxU3YMnwAc84pgID0s/92sFaYtxtekwpFIiJQNLa1
u74y7m8zvw/nZncyjH0D6repCCbcl1qdsBI36wsB/lciWE2ubI0bak+IK2qMyBmQ
Kv8Yb5V0MhUCQy7VGhE0gCFDfhUsKPzVGAJEa9mn5Fi63weJLVeg70WmyWC09jRY
yg2tzMvhqEO6kIhiEkFXX7sP9kNb6gXSTl5PdXSzq02V/MK266jZ46mqh5tRHoct
1DEGtEI4Rxb7kPEUI0zzyj2YlucctVlw47g7yIeFoOcR15YHXoCTDZZIiz2JipVS
Gs3GU3hbLygUjgQzeBW0PgDKcD28XHFfkcCW1tgGmyFT+JweKLV5oZ1Hl98iLzdE
EVrxuLIBR4HsjsAi7lWCFhYjXVOfLMPZckAFVHjQO+2QK+zTMzRWx/i29kXd3JlL
UVk5ym25MLyjoi6C9wzy7e/H6FBnpDUPzGfEEuoU1tw5AAtgzHTK1JZyMJAoP/Y7
9hIAGHTOReOUafDslEgx7OiQVA4KwJgkkNeskwwHq5cxw7FtgGo+bGXX4yVuCeG8
6XAaIUGCTPiHWEz9ogU5zlykJ6vm+MSJwVInaiYtaX++luFzmDe8ytI2EXyCT8oZ
t9XdAnpodGsUBlyoTZ0wNswrUjNWFrxAb/0sUWx1GkT10WSd8paUcaZ/DL7nZ6hW
Oe9jkeYiVgx9CpfN4YPWZhbz2/EMopVqVH3CtgZc3cPYPp4JFIdqNjNrVBgXXGAU
fUEUGcog3YoR7SDHarZVDXg59g5fVSk3r6dq6KU2mZzDmD1cwy18TjroOdYwzZqV
YKNk7rFArT1lO26MFo1VAMg4XUHnjiJFUBAFzzoQzqrBglSoBVZxYfD2R5ojGtQj
qICn/1FyZP8fDXdOrBAdIIK5RRQpbPYVHLz7C+K71hW/hQygUFT/9K+tEOw0MmUi
sKrMppRpJjwdAEJ4GHkhrhk+ly23g8nNHwafWYbVgwtduQfWkohPW67P7wq3SZXW
axOPkNy4G5YtWhxhBJXqzatS4tg3Z0G4dVGONAUr+Z5TALh9Y3B9PpcTlrjAl0Pf
W/tdXiRQNZ+eRp5oTfRDs/YNra8lD2Fn1A4bvrZ7svtJD3reTsJxc2w9gs/SYHwA
yPcfJcVdBBgCSkWDT95u2Bqkzc7pnMmLdw5C4OvhS1k3Yi4qdhkUFGl9/zB6+UUR
gTH3ZfVLb/CUATYwLDNbFs846IGr95jev4RMhukKFvCAMu+fHbPslaV5KkniK3oQ
9dm536SsLKCvEle2+WODEpSEfSNtqDRZbrGyH8OyRJoETFKsBz3NCyxrJBZS8xxy
R7/aEX0n/rdICB3+bbF+n/kKQSjl+JW4O8IAhldssfbm4pbthtbtVYYBuN6YHIXU
XxerA6tETCaOcaPkz8Rc8x7xI62N8hUBE+ja8shS60CkI199bvwsWkPqf5Ui/EXP
NNpDffNXdaXrXJxXAcRUXHCn2qL1q9YFFpmlwEPwcF5fH9djPagxYmlJG9QkZVYK
NeygTRSSfAADyUsAPEp1VexjDXoAQASkO8N5i501pn0NHNIKIejhJRp3+yTYTMbQ
T5JvRFQG4ePUzWl50d7o9EQZ9Ddh3nvOV0wDfzKvvYZ5FO+tNqC7LXABj9ZPa5dK
tkGQIK4ZY8r/uqDLQT1Pfcn8BDBX9uJZckvt+NsI+pqVkx9G3ZbKyeCnFLoq3rcE
5KTPvILfXXNSsu/N2UweLdPF8Uk4BVyZGF3KEsu1Zg7ToWQWppTY26T7n6SrtLoc
4EdccJ/h0m6JLF7RmJ+9ow==
`protect END_PROTECTED
