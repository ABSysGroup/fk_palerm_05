`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0QdnOUvbKTO64NNzZiei7SR4VsFcR3ADlDkwXl9hW/vFeGn/Gd4Ep1vfH8jI9ca7
9EByTYz42W7gqWAGFyCOhZdaAJbE4JKwSddoiKmHMCd2sIAl5MrjuO5Lu2bb2SGD
rcaycJk6M5c5zzhbxh54ZdDh/QUdPnll8ZlsD9j6pCSlmvF5BOx51nGpgdt69A0F
eM3xRoXChDHbIz37+awYbJ0ExOP4svrr64ecHlBX7CmYh2AMzXJlZ3pW59tOr9ln
`protect END_PROTECTED
