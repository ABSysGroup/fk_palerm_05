`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zl7RShttWp48YsZ4cDO949LpTiL+Hw6Um/KM7ZF4OChY8D9OWogBwEiz37kLlTxU
mLVLZjTQjnaDqjTMjWAj9NIsU7VuX0iSVeTlxxqwlHCmcJKsigv/3Mnl0EcDLxSm
Ild8qvHsmCpklRIUrcSD3Qh2t5z9iYsN4owZhRHd6lhu/a1CHqPoK/ZOd528y9BQ
UDwCIWF9dWJfBhwnG5cla7uAUq7bI3grjJalsjsbpvj/ChTmx/yL7puCyg6fdx+0
2lYLZ8dShP+ohJt0lR20JyZpp5GdzvW8Y72u0wdkHLFyuvzqfu3cmIUCotGbT/g8
V5lK1h5qTvgrw9yuhsZfVGVItfduN38vEWI10WYRYQEhcUFLNQ41wSONzVJpj1HS
2tctcclMLs2+i25sLiZPS4o++yEMVavro5E3m+NIwwzp5SedvBN2g92BPNEJhHO9
K0arWywzcMdNK5Qtvr+s5/xN0v04/5GyRyVY2mhoxeuID8QsQfnfo84QfSX5lYI0
3KRpMKkiaFmofbBDYOJdJiBTxaUPt4Cb+nhtgmSdnB6h3pIB70VAT32U6To4kmgu
8wEw6N4z/ZtGABlm/fjDflk5ONXuFdGgiz9+HjW0468rV/R76njulGg9iJygvdpR
CkJG0Ez7ofu9lsMTWH+j06iUdiJMb1L2uGYOsEqTYYdIta2PMZO+7Ocar6MU+2hv
2zgnshAjuZ+ZMnDv5v03Abe7GNS755vLmsNYUoibRpSz++ZB+//rat9NftyyGICe
DRvOFM2rPlA4uN2xLESSVPXv/Yf3WkP+DOnt4fHgx4aKxIAddCLgvRSTUxm69yaZ
9m+CfetgEZywlHdagHVWL8OvVhTUE3rIVO/fl4sh4F9VMcW3K+wj1Ds0fLY4nnQm
LLGE16T6tFg+sJapp3g0jKZLV4LIxXsTB8NfwgKjDWc/YPfDQW2hnpzv+C1bxyUa
`protect END_PROTECTED
