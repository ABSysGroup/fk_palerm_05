`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/V+6OkM0Xs5syhFwTy9UQVW6buP3fqWRSxAvbSN97/YlR2OTioK4aD4J/RCprb5R
pINfORq3fiBKpUAEwVx5CV21rMjEWynU3QXZxVcsVdZCGNu2W4+sy9d3qsrl599m
/vwIAHGcUmSgYgop70KUDoyxPg79AY0UZRh6JBtgbQzued+mTAbMfu5VTjTFbqIh
j54b9iwn1CKdjPBi0A1SYOqSkDZY+rC5ek1Erd509lXlvWsL/qw9ArmaAHT5szDT
Aerno+jQ4HflZAtjpMBBZ/fWDb+WruKdkYcg4xfA3qVsuSG94/e+XaF4wgeByTkS
qMa6knVo9bvKr2Ga6DjBBkuGrlveqK08iMnldDUlJ8qetD3tGc9UMzaEFAAvi70T
/Mq1y1PecUVrDtcCWNfz5bjrLJ6XsVL+EOzQT39VS4V4q9qVYjASsB3Fe+//plP1
CKGOQaXv+CMGc90gU0A5XpE2U6HOLtWTxvGc+FNEl3PzBC9TL78AV66ATzzogvGS
C0C4zwjezDKZGYkymZXVrMQNPwe/tivM1zWYkR2dJhqOeB8Ht4M6x+4vPCTHTeRe
`protect END_PROTECTED
