`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aSldEthxAGTxUUbwWP0K3zheRYUDbYOpU9I8LlaXbVPpXVnTC95HcWhyPLgY9l5m
O/eKgwqKetQEqPQFrw/nxSWpegw8HMrcRx922gT+BraaSRtIt1/mCAhQvbj+DYht
CtzAD+ScPgJqBcyH0x3821TlXY7d/nAwuJlBiz37vgbWnhSszUG3QK74t5rP/yhT
LRyWgHTHyBnBzDeOiIORp0YvskeSVFvRN5C1mvGBUipVMGygpCDp0LRi342ZH7kG
Slk4Pm/Yv7R5Z3LCe5L15tDtuJXD76Q8v/J6nPDy9HA2fxwib8Fd6+s2Y4wk5oZ7
4iVdJSRYoVHhE3/JpkUeCw==
`protect END_PROTECTED
