`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dC+GIQtlu428lXqbS42ocbcudG++anBIprv9mXCBcs29mJTZOOWFLpC7SZ/sr2ko
IqFMi4YPJZM0w+WEt2f05D8paq3ERm6gyFiBCsd9/FvrTh85hmRPg2wLmq+ZUf3S
rnHij6PN7NQVxs99a0STo546ixKX2VLoDY4IiwcDAZU++qq7Bhijx3dLAuutShad
GioJ0TLnglCXGhlMvDNMNWBPs4DQsMprLNNIB8ZI0I8l89K+5vw5959qdGYEakX/
3AD/eDbi/DyiX6KQupYjzoghvhXho+X6eCQOXn8qgybj4fQqDZrJ3+ksntekm1lG
YVOYeB9SgKqXepBJniS6rkICX75MYp10+ifaq58JCn/2nZnC0SbIufFkJyHj2RNN
IxZPmPTAzZROBZAWQEt5b5bVOJpfDq0hWZyGfvoEmDhGZBD0ESj1minxRgC4WfTO
KXk6g64/0gkOlHnfCwiFj2zRvt7nxqC7dzbrIVQHjmKgdRHUJuXgIvxhTr59qBzj
8pccRD7/8fa7VCSCSJfdSTrn31GIAcw4gipZWQ6NmaSd+SJ/F3fhaXZakBkIVl7E
RFvY1cYGYTMhwTGb3limyF/SY6CGYm0Y6UTZHaJpwg1jxeLoze5T/llIFG2V6Y0f
cp0ZxsG4NTEHsmNSgCGZO8MA5STTEqmVOziv9/N2Iwt5hurdEMW/PM4olSygfexq
pOLooXxC23NrQOKn08vpRPrJPNw5YFpfAG1zp93c1rpc8MuxVIgbB+XdEON+FTWV
Z/cwSE++8EiGbvgyD8OJXGdOxvqdMbDzlAyMudP1CKZBmKWAIQNmLJNquxeaPYoJ
QtpcPJGLcXPYcuquTPhhhfQ5vA8lQNOWjqtke7UR0vA=
`protect END_PROTECTED
