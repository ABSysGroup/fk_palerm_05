`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IjSX8upZFrO/KaxpoImOcb82uwp+Co+/c3YWe2+dnnfrj2jkOZSpv6wAwiUKxZ8G
C9q0Wx+oWpAOIObfj9mQkP91jYt68bhzB9Otdh3TtHDukjUq406Lqt3GrAhQBVD7
0wjEeV7a5wc0jNR2JynDer+ZP2aevkDbuRsbTtRGf0MbJ55Qe/1r3W/BfQu/GEmm
cDm0YDcWrlitZVyQ3rOgTIgBX6FYLbiJv5+BAPGBAqOR5WXb0CHZZiXbTH8By+bV
sqzkLctDZw0tCMLk2JQRqbDdn3v66wTD7rf3oqncU3K5gLmAVLXQaBDCMhU7VH7R
rwM+Ym3YQvRvbuII+M7sgdzX/+N378+TMKtx0UUjtpKxUZC8w+5/mOZPWcSVQSxV
6UG7T6L3D76qi7vw1l+7Kn4J1qtWuNL9AzBrQXXys2WQts7j9F4dSufGEw1DU+Nb
z/F9cowHNefUvunoVaDpmwXdsJxXhTAhg0jUUdA1wiZ8ZEZC9pFgVL4PeygRm1Ze
7ZHmHR8bdEbmYXp80UGZ6seSuaSIpsANXYNq/Jt11OPJmo65XydAGjAIU3U5ikF7
UO31ECEgMHamy5bWgVLonQL3jLVD9r6RcwOdpvtdeu8sQCNCtQjOblxpUuUHi1Gp
be4CxbfWmN84YWlsStiQeHJbZedzC0MIx22cAAPTIxu7FuOMElapNKoxRq47VIcg
1FTjbLsewNRMTR/0vSpE7clJXno5P1EUs0gHK6esORxtPB7vE4fcNc+tTzcyVnnJ
l8nZu+SutANAglwOsh7wTfhlzYECs6opC35UaUavoNgefzlF7WvU5iK0lp8W6IX+
GxgxnkRuFbZnUA+yTO8N3G2bX212jB6cdeWdvhr30Bl+cZjj4MJDee/GQtj/PBtk
9Ln7JKr9gDcQU+JY6DLrpmajb06KPHATHLBQBgWWJvxq5kfgQgidVpJTq7usckJU
Lx7Evep7ouwdhEESrzLUItaS1K2PWg4lBBj6S1gG/t55csUPRgUaiek71dHLz12O
11r4gkYJ8iF7J1czyaWdPFgZzsuHIRD4jIOiBSI8txkCwgOgzOQn76nnjje+ibJm
6ipi8ap1Ygrx6WY/DA0vjL7AriyTP0R/UT4r0uXyV/Qi2GW5gdoIuPZq8GtFfDGB
4Ba173sh2bg7cf2XfatO63TdpiyWoG3RPfLHz/0hHoUBF+3er04jAhi35acPe8UI
vg7QkBvpNDba70nXHav98imTV0A1SIh1jqUWKmA52RcQjeZlCuaytQLOjGx1AKTQ
xLPQvCbVIBjEbsc7hz/J5XiFxKg+nLkXpNksIYlKCdWt0/mLieyYxja0uNKJqdEn
bBzNFn8a86ORtqIocG6xkZajgPofYvzNjk1BadftaotKHEGGLHlQinIhvwg9rNz4
hFN/nD7zJcM9gB7EHnzT0sSKMxzdHSmJTHv9N57EVQyoysuVQmX0lkXgWZKnUB3O
Rpu8G5nOQMq+JAvts4BcyrjeHVlTlMM0m3IMImlXEwne9dxPxyRoTtNHDZIxYQkx
JliI669yHeVFoVKfYhh13kDKf0AiXg0sg6o/zale2fYsiHDIiPoHr8r/G5s0Z4yP
/381Iz5UuBFbiVzM60CBSZgblQzb628mL2/dvP5WUqRRZzv9TJSZpUlucasWSqnU
47ZG7eLKcbrQ2moeuJEhZAammk6ZYt852rZSSoHPYPXS6jxJ+S4XiL+TNCR5RXxF
lfDc7+tVKUF+wzkBJ2J8kIp4GJrEQcB6EcxXmQSBfHXJTdKDqEStrtcXlYCKL9fe
cqZG218HN6PmTghXtPBTnC9nV0C4RcGa3k7+M/b4w3U=
`protect END_PROTECTED
