`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lo+GOpKiRFllHqvwj5hOings2kjv6GlFYpDlrwS7tb4Y/a2+YkF8cdIj1oTm2EoR
jZmNnxLSmrg0CQoXfxO2qqoLcstMJxmUXvjyq2aeHXcVRMAsRKUB2DW3YkStl1Cz
Z7tZy9rXm8HeKTUMUHfPg9NbjdH0MYmFVBtJYQOnBEscK/Hak+TGVb5XuTHNQEbv
GGO6V8bnU2jJjqtsVbGvWBxvgsY0DhxvkyT/C4JHFw6x+yXedxW8ONhaPM40nf33
cxrn/ywatfV2MoLXIMmZ1wa4VR2GkRqFQEQult9CIRU/bsTwZOWBmtf6tEiF6iEL
jfnLj9BpMP/IRv12I6fpKAGiJFMH2T+p19LikBL1To58NOmua6Fc0Qezo+hFsaIo
y3VqNaj6hvjJe5PLaNu0gfGEsr4O5B/TGgM1W6XcKkVig9ny0DaCUKV5UjhY1w2q
lLg4dV1+ceVwpObuZ4rtIlqnkGGwW+JNZHUWawErOu5DupC9Ovj2Z2sivLGKbnN+
UzrXA8xx2+7SiJAoNQd8TJTimulz3OhF7gQfrNWz5JprsyCEfD01G5Z1bRV7xodZ
/aPfd0YoF69t4AmuL38xpZlHOF6h5R5PL3RtuH3snWpb8IH9J7UxQTItPMAK+v6O
yERXfeJMz3yqpbVtEFWNyu8/XV13lUiQt1alEx7NaMzrE6D7XolZ/Jh7mXyCghEv
mgsyqucJrEXRmBl93euYR0LZsVDGCJ+7UNwWEmxR8EPjWdODEIKGWBaBtrHGpTCM
gI9FzRlQypGtr9TBI3pOoGoY/38Ag5qYp2jqo2j7+KSAKzmNyeAivnZ6/3dNtiV/
Gu9bUAzT42PrC2qCGCWFM97VVyem/q0p10TLpTFbKgSFRKHc439lS6RSm8EvzCm2
pSwBNfSZ1YECcWLIS0iM2U1DZWuvxrURiKkgP2U4jAAkKIyn8Lmx1iWOK9AF+6L1
U74afsCvavxAi1HAov9Ox+X0dRizW/fm4+LvIT0NJB2bg7ESq2dNqb96obacGtj7
UKQCUSIRzEe5N4KX9SJmkQRm5F3Fi/Hw2ExLyJJ7LABGclc7Kc8HtvCxv0+h0faK
jVt7iposcThRRTwlnV/21xIfgXjdZWvRv704YkkCuUgiKp8fP3FLVcxbs4A3maV9
66FFYR/bE0pTPxFgWMZQXL66SnYk/eJbkY3S2eAwW8ASA1UtHfKs93IRsLDICd54
o46f1OXBfEAMdDFC2EmLnmIgtrhlPqtwj9NS/qJTz+AxxZOs5WCF4GcHJ7kXEQhs
FTvXFnuKZ2QHDXmlAZzCbAX/NsmrImYC1QLNY4dCtWNYDz29SBLme0pzmqFKpZIo
q+hXGTbNSzm/APKvKwoJuNnkJK1CNi6ehwAdvd2oiKcLQUWQ8RNXOP0yi8UYFz8K
GSvbzPg2azgSj4wWmhGX9VKgQ5sCKI+ewT5703b7IgH1o4a6dDvIfYhyPDuY9uG+
jAQIgB22WHZ/+sUtFzXZK5O4Q446nVrO4UB6R3UgekVkPRayLPLVnRn3syJF3wek
1j2aU7PJ1LNFciNLG4cgX6+QbYGKuAMzkrj17Pptsi8xH0eOP1tFq9zLJnEUe4yq
Wrr2iyWDu+rkxjcL4vZIFwTTVdz1RmZObsON7oW1oQNLLrjjKLh0E70cpkVI7EXR
ETRIo76fVfGCRm+7xTS1gYlZseFwJ/bp/S4wq4tY8JAozFu7343frtU+cEJ9YmWC
nswZrSdx+8xT/w3slY7sd7zaUgMrHwxbGZ36d76mWMnndxScB2LfDLYFh/+A1p+P
tDXQ5rwWgqoCQ8dMCRuvRfBdLUStkiNPHbdAv6IuMrkvRbsp68DtN31D5edaOt5P
n2dptwLGtjlLbhT16lQKsfkrub19+Gnd+LB0dXm0xoLPd7pmM1C7CnSIBmucxCmh
7UuI6A+j+GRkzSZMyErz1lJdJOY+zKVxHumAc82HBaQlw9/eqMQqUX17wks9w0Yn
4+vgvMkKtTpRKb1r3K3efocrVHrMkDW1geZUlSWO3rv+/512FC8p/ZIUITKp3n7g
+Qttt2KRO7fovBU/YOPP3ZHWvcJFIQ5hpyPFM3f8Lzh588/LiyFbGSmmWXSbugqM
EkGE1OzbGDh47JrpxQWIdFz78pMwceKIwRNbjdz1/k2Xz4Q14CEYDbd5/tBUxSty
pmwElLM6iPXZi4BPL5wSqd1ScQVUFngRRZKfeqG/e7HbezVYE4SKMkhM3LRfghJK
2czVhEQXxgD2uUCymkZ0EYYD/tuMpDTkmZYwNBKKmog0wX/u/ZvTMRZqMcLLH6+3
h6P0J2YhtjUdr2ECt5Q+08Wag05mWLtv2c6QC7g8UqBp1GFthegnPdBOZfthbgl4
rLY+5yynQoHu9uphWf1qiTiDDjKmUBVOuhNvCM9IysZVU0eJ1mRetig0kzVkz1Ol
9E2CduwQyUqIewxIwSHql9kMVpWqb20JUgffMf327yTVKgzHRxu52N2Lk9CmWSNn
ATZvVgY4QKH8QCC5eUp1YEzfWKrVxnMiJsJX2Ts6uRP5xPkjPPd9j+dUwwbwxWzq
mt4/Ums9y/mEHkASC93FAuDkEtni0WOsGq+hIWOTRr5RdYW0BLX/FlSSITXOsFiD
a+hV8YVpfy63NFt7czurPrsk+j1Ye1bKuSN/HlZeNbZY8KEenJSwGcV7BQleubLy
4xZEPWRoAK2EIUZKhOAy63cMo3MUpHazfP0+JYpugEEmiuN/dKQ/VpZ60q6D4nhw
qtSpIyvBq/F/KSBwvi2ydggD5k9ouZoQzooZzNRfnnWL4EWc+ociuy+u4kf6AFCo
4oiE3C5tw/x1sKT7idcByYA4BnE7GPq6K+/K/K+LvLPvD7TvCcJ+T5P4vFB1G7Mf
a9c2wTfm+6YabmWNb0XWMt3s6GLdmvyQUze+78WAB5X7GQ2AdnXbWpWN7/46f0do
aeoUvaGVOu+IDs+MgWVvIqdgyvC4I1q8ZFGMQNit51xKDIvIRMolWGnvdbi+UB35
eEXaCsVfKm2TUSw5OxSKyzbbMGbxnSxHw4st3CtRskMovEt4WEQt0JhlKptFkH2Y
sz6083q9thvi8kjMeQ24AV0v3VvJ7AxnROsELnAR9xK5bjNY/Jyt0D9SPYzFjSB8
RwcwvoTwKznenvhiFnrqZNHBEs84jXogX6X5cAUHp4jJ/E8uKwInx94z9o6YsZTK
LsluGM5WRi2zWjJWJv7cRZECZfJanK+i/C2jE54irhQVREqKsmHssdEVwNTlP2Ua
T1Q/ocDii27Z5holnC3iGmMGmnWZTeWXr3+WZzFyeQMqhTxS9v05gOLZULS2A66I
f0RGh2idwLg5/fDWgiwwJgnWv1ew56r9NUT6CTzdnHyjVPjGL6WZOnoHa8KhXhMq
Jo+tD7YFwaX8Fn5YsG1RCHGRV7qkgz2LvvniDxUsHzbIiRy1tgUxWCm0jbU25JV1
oc4P8Hm2/TClaVY6lkHfvp26cSwlBAl1XoyV/4o+6fg06BNN0L745RbZoywgEMeX
iB8Mq0WzSfE2yEHjp6E+2mqvs6PPrP/tfQlVxdi9ggd35JpJLYQWtqhkh9l9WWhl
TB5X8NFq+dLWAJwFiTs5sOnkWt9rPhgp6eOiQTiXVtvKAncrqbpgDavBQauVQyax
6SWZJ+M4SyDU6bdIQtO63qaqp9RWD6NUJJ5mUgAfTfsrNYowmPzRybLYjbkSa1yH
3sP9Q59xCRflyKHnUi+/UiIvWAXISyiTfHp4wBbmHD8hXsf61O9vvp9HImTqWDGt
z60buoaGmAIbaRhh53DslA==
`protect END_PROTECTED
