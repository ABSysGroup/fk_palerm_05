`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6485/o+wAFJ62pfJngNCqhUFLolU7so7WvyMd3y1fX5Hslr5aaOf8MQvDPYq3dyS
/yeuXPtwLVtYYFeWxBqS0Sd3SwzAPN1XjBxDM6AszIphKtu3p4fcbBsPdTVKNzMq
B270hwbbXf2pP2EsIsSLgfAi31PYkQP9qxwVAfWFxAolfsa4m/v2YkjlaMhvND8u
PwoyXh46ShP6d0xvn+2abvZMXGFGN8ymgF2vN3C4fXG/CG5cs1cdanc5njgSoqTl
jaVfdG3TqBeT6RpcXDo99XBq7UfAmeZn81FmVbrEPLwRk/i+7WHHP1I3zH0+N8Jr
s+NIkpUDtCxMaY1YGunmmX/8rgZS7gsN1Ytk1RviySHiVPa00eMFw0ubN7RS45uM
nzGZ5d4zqtdFMDmQi6HcB2ePpXk2OqAHuMuIyJqSFWi3DQMCQuFVWrKS/vZYQLTl
1ecJsWuLWR9VdoaXBV4YKnE+DTaA6gp/CafzWsbs/punvkpGcaM3gMeAcNzmqzt6
JiWRllZhwntfdquy+ZByQ3aHlPncCBm9ECsFwvE9gfjIInrd/byDtyu8RPTk5L88
iNOLD5juxio2OJnwVcabU8f88iCoTs9BtX7xEJ12EgS2lnoYfoZXVP0MJoobNLGp
MTPOhmTc8WuqNhFndNyGpw==
`protect END_PROTECTED
