`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+JMOz/mVqa/HpWUYP0xYZFHmYsReRtIKA0bvVGYmPlHrAIAhc6jIZUxvZtREgrLR
eumjUBnpkCrcAeakLLc8FFSxaPYRtgfVZrQF43HYvA8bD5gce7uOPNBSER9R/FfI
cfQq6p2bvBGvdfnCbTihdMGihxZj2FAqAzn6xSdYwPyDiMti8Y0ScgWVJ2wjxlyA
KVKkXqJSr0+bMRlgfoyKR+8Ykhq1FINTqrWhRMpzKc9WLfWXRZAkXRID8DbFAtAz
Au0sRaejuUQ66XRh+pbW36mPzjmsaDVpOPlC+xXk58jJIq7+gXLPHNsYhArjaJtl
6xiIaSoFMo6/2Wq+YmTfU826vT04dOXvhf1Z2zXNlzCV4/+1+g6lnoWVLSVBhuK4
s2YkDxTmufWVX/F4yq56EPeMXNpDQDkhp3Snu7KSYPm7Gjias+z/oT/DvfhU2Jqa
`protect END_PROTECTED
