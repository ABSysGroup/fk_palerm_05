`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gSUTHthRBaTJZLJw/sF4lZLwMso/j0My+DmKTekN8zpqbaa4JzSJrzhlnItHCFcW
RfouaN1cDS69MEQftK0uxK5+7E58LKRMbFJOC8HNpsjsQDGmNsAf6ZJbPbnX45lg
rHQbdcdaHbIm9IndZ4mrMY/zbd1b0dgwvSMG8S6TAgFXYv9bWiXv7/XcyoGZNHT8
K1Qk7012ygJ2YlBKYJ7NWyABamYv3zBI/KRrS/8UqoaD9yDuEveLtc/NFbmJLjk8
VBvy0UZH8bbx08CwD6wnmfEzpP1r1iV7gWr/EIqaXu0iSU4da8qbXRx44rQ1f6dB
U97oO2XdZzGlqBnBYH9t+q8pMAg7IKmjM5hxpCYkZjaFo4Amj0NWKORuipIhn9FL
9FMlZvTiLLeJMWF7MJjuNYrECgYVWdRRQ+CVwNHlDgt2Su/QnWhnBJd+DA0qCHr/
A0nXu2fTWZll0o72wfS3kw==
`protect END_PROTECTED
