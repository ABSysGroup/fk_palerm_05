`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dRE2eSRL3a2ke3zlSx9/5O3o3DiZyTWFvl7Tu48dW/FMtWuZ6rnAkYooZiFl72Ci
8vzlkneA5F0eKoV957vAppngP8Q76hg60h91/U0QZ+7Xy45vJXBcwnAMJZdyBUzU
NXHKYn4k1DmKOCQMmzqzXQ5Q3u+mrpgWwMdtbcAZWA8WK9dt0zYeEL9XbNIIlSj8
JlxzIm5sczjDV6El9cO7nqgkZycIgpyFNXDyqWS2RM7qLpiMGIpuwNedaa388XBi
2qfTl2JCkFMmC57FV1uESwPGLZr/D9xfCqLz0GQyH3K1zuoMoUuwpkomYHlCKUg6
k2Mbee5ibLTbfYGQDs6pNMD+fpUCuZ2GDIGCE9po9Qwms/0sunKvD8s53D6dPaxB
ZArVt4KZs1OAK0G5xtotGEyoXid/S9b6l8GjMGUVirZHqqVxkYM/9H04vSuYdLGw
8/lJ/UHXQ12Q61APVKQYSdfPDTG0HN6aD1DeMCSMK7Sbrg/eBBi9JMj78VLX+bde
p0DjSg63OPTm2IvgndhEafVBkj5eOvClR4Uz7Oiv4XIT8Dy8/Po6moKzeQqvfmBk
7tyNpzFvShrVpaBCNoci8kvEnHB2XOraKfmjNSDTGUURyIRvryPVf0zJBNAkTmhp
L56YxUwjeWyE9uQ+ErRzOAR5Ej2VO2BT19IKITIGNslijaapiClEawoBDoycN5Yp
wUi2RpB7yArACLNMKKvEAs9LgSv0t6gfZC4hLg0Leoh5nql/QzhtBeX2PVgCREtG
vz6DpjbEjs42lQGV+g2m6t3R7UTAQ7/vcldmk0qetRUpXXVfKjNFmSAoQqnT/3we
61OhgY+Ye7TNRnuohMs7LlmUTU8WrYPHtNcylfjkAuJ+okj+SAiOYVqFSx3EzY/o
GvRZ97ixwTHJi/5n/DLDUMGNW4Cxaj/29iIIx1C7YE7R422CBw/J1TSbApImslPc
BGjl2iX6oSAbSrO/VFOBCaYdBdNndAmXz5mfPi+VldWCCt4nOD79lQ1KzZjFP0Tt
PrF0syxhR48hch0m74Ok70iVYv95EgbX7uSxgZ/Bqd/ujJrWl1FQ7LZE5Qvu9HGA
R8Lh+KEjaPWPmR96c+HSZkzTODUIFYntAn6wmnh4VKgrKAbEqllXMuI2kr2aFwY6
mWlZlfX7bJaUmKuThgsrcuhog3bQvnNbeaRPrTmjS4oVr4O0Jzli+rqjg7pUNwzw
El4MiESRcxz02KemqLdzxRNrBD772EJnPWTHwCeEOO0zKnCXumVDu6nvZAhtjbNE
0MJscwtllel7miw9JXiE0yBhM6ai13aDM1/wYQXNmpRF1G4OhcZH66B2ck8lHkG8
ExJSsRl39TOgqzzUJbG+53r1u6SOaXLWV66v6LnXSx7vOYyeCg4h/HmYfCOMclYh
wNe7UOMaYBi+F+c+OeDBQtHNE0zUC5FV2+8FbBxFLiQ3IgVk74G2BBbvOz02m/JQ
Qij9iTP+WX2zqR8Bi/Q8ATLqbxg+GXbRhU3LtJhFgLrRGgnZdXXaOk7kzd6ZxCqg
6/+lJKT2Y/aY6DQezz/zKDfQfnb74D/B8DtLorxHDcGNasCKWlLy5TvKJv7FO6Pl
9+PJOtgVtu21aggYN7oqvdLU0PIuBoL4c6hF1zTKwDc0WKrtrYlUUUFyFuUqQD27
9AnwR5h0JM2BsosVm7cfc+zLRwEQNgxgLFk/svH1VaZlO6EmYIDo1zBoJCzmwfm0
JVDzFNuniYEVUD2ny73L24YpltX9chvqLqBLnIJ0h+N7Lf5qZKmUA+QNaMZAEIDV
ZX6WfmbhQrtWcOmvmn5oJDz3sX8hfxz2nADQkTlIE9rKs6weKqiRxcPe+AL6csQ6
S8S+yV676xrx12c7QIU2zZH5UDGfzOun8KBRL1sMSMdysmTRrQmJO/6dEQ4MLvB9
ldcoQ/ScaTVxN2GNCYI7xgdQjLaMne8wCZPL+6dwoLY+ulnxtKGioCSw0qCrrnvf
0gvnEnCOEuwqbEyAhmVvr91DL/WiwghBtZwTyqSspr3GsgCcAxryLWvgdiE9xAh6
aIXag8NvuI3KpwtseCC0A0Ycw98tSsqRniJW5krulGAMaX7YMZqzZ+3uoa1RA9MZ
MppAZHxCpISVaBUlHj8P7NVks/BkXrXBmQGOzB17c5SxF5PEIqHVxRPWHedbnO3h
jbOk4Iklqi0Wvxt8I1sbP9vdmKIdc4PMxmoZiYbpac2hiihQaY2WlIFNYYCrjy8C
6qnJrMeKQHacWsfB9b1unt5Sr/aUsJRsSOGv2P2o/sCuKMZEQramHKzvQKkjxWPO
0zJn85V3vVIcLV04pmLUPcOI0eyg4PbSM62xukxHeHgOk5UK73RlRHNGrdHWyDmZ
8OjNaIqgh5OXOpq0XeYOPoTx2wl/0X8sjKQ5knMPoZf3KKnJwIWRiSrnRff5MgK1
TOo/PHzaEphUtfUBxeztefV2T2iNB0ZBsnD4XjHH3ex9z/G8XDjELe6Dji1ijmUP
TcDQR0YtwIERQSImM/Ep43d1GUpHdB+oOcmFgMwcARtwgvbm32ccRr1ateZrQ0v0
wkHn0HWRAxAMF0pvuzvWieM/ltO6oYBE4y0eCCxcjAHqoBuxGSG4eK1rqNXFbmK0
CgqWHGNs7yLwVZLxzyrav0mpbVg2waFmJ1Z5M+wZ0Ya6IFc8km0NSzWV/xMGXaoI
Ms/DZBlNpWCxTwmQ/bjaczf9BaxhOVMJ5SJb9BiwGHXJPcFDgy2vPZssPjKlYX5w
sl0O+xCCddkrteYkbr4+6JEhvnqR12t8sKoMPuCvE2UGX+OkLapb4xEZlvhajSoW
qTZsnAYEksGoPE6SUMTtFf48IIEpBU8s00ywoQqZdz04hucBMlYk/HTyAtyGDzHZ
2mMYv8Dd3rpR1i+qmOwX4MODw3L/Foh2Qmtz5EVcjqPLsiPw9ZFKIgc9AR3N2psr
0FuX7gUJz7mqWO2cO2R/DXMk0odUyXwwG8ReR4IiRnj2n65OVTE6NuiCuRoGqDrS
9z0r+k/U+SDKma4CuBFMuyK3Wb0170/bRkDb5EYRrLYoDJ9HQvN6FwogdSfy+gyJ
WiJTTShK2OwqsItwbGj8qEFS8I+IzqPeXoxhbYgJKI6vDJ41fjjRSudZ6BVAARb+
rk0k8Zub4M5zeZr2K4fYuOr8wXALWij5PGTYxvPe5XptHkLf0oWFAZLsp/HndET2
F7coYxEJMwLuSlW6J3tHDNxfP0Y7kxT1OyHU5MyWoKGlgJKCbBjJOhRr6kECcxE4
eKu2qrs31dmmZE5QUiBfRcoRkMf5uSKmSt34Fsbp9F5aB1qvcA3M4tagpunnCrDo
E3VleBJ9QQpZMVFWOHkiGDk49TkSJwMcHcpXWjZsR9tj+c5w0h/1AKKgAyrnb6yM
nnxuZsHNZM+RP6DpamBRRFegmqFfgcCHJ5Cu4+aOGZVwPTM5g4CGImuZVScPFFPp
blsjlvWpSAalwHIANulSRKpZmIbbBbgGcw7sAP1zJtnTtqCHhjwcBvy2hx08/zXc
RuHnLwxG8Q6xlXcDMJck7uDJZ00DEwR/6iArsraCKO87Obd6FfwFIHh75nIWCLx3
E+M8a8a4ewcqTSTYp6yBM1pyUuy5F+IiPtkGwrmSwFI=
`protect END_PROTECTED
