`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RXuRpFT2rWFNoBDhMcbwI3JrYCwk4RkouIfXidPWf194FC1M/zr83IJTYcS62K7h
sCMO46LIyhUm10Js1d1+Q1yYXyIV61QBAcj/qaaNxjJEsHIT+DYwfXHneK2yXpuL
gnjC+pOTPzoK0L+AuhO+stKqbJSQ/2josEAeNC7iqwwkmRTwDrZmHLrrVM5qHRP3
ulBaMbcWbQjD39PWbGwlXUo4hmukqfKvq7xHbrz2RhscVa2O1IZauN59gv+AEDk4
e+HaavavZ6HIeewxtut+lNyRnEUlNFEwaMLWkL94tkRgQO4z94w0AAex6A3jV0Y9
9leCvKd7af0VgjHeQozgMNvCNviIDkwjrUa6rxpL7Lrn1+ZZxIzjpbW4ZkVwNhKj
JOyVYszm1Y9maQoYPFfAULOmB4xO+h0QO0lepgfriuEcAASNonbDq+83GfCsrRaJ
`protect END_PROTECTED
