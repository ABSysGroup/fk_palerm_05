`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oATp/AeKH6Kehp7EFJmrj6bPi9mtKAEh0Tr9v5NbvuHTPnPQYnXG2NaErMLBwPO5
J7HcokyDxodr2fOtP854K4jjCUVHL9yudc6IVTvyIRSU5XEroWH7APapVn7HFGtf
kDjZZo/5yf1b6dPkD7y2y+HT6/Hk4o6W/sFf+dyP0Q7qIs6GjCyyVcvMP5iTNyRu
Nlfd30rPeFgzhSZ2g8iALh3v3HmoeZrjYQ3iutsfJbaNKHfd+BQclAPNaCsihQUo
OilYCgbtYVwB0dWNWN3bk2mSo2jv/FQ9WzixIJF1NiZSf+Pm03Tss8PDHHprV6dE
Di81hF8DatJvZ3WpKf8n8+Pdk3ztKlPEdtoonm0fEKaU5joNsBI97JB/9crJ6AFt
tO6viD3KSHtoI/NbZSGpsezBkB/oKokMqOFBOSKzyEJEEw4PNFRsumvJ/n3WllF6
`protect END_PROTECTED
