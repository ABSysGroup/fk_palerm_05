`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WNmn9iuE47BRF1J8wOM+1mfXm0ztfIbUNfObCYXq9itKOw7Lh6RqB77m+BoHrckj
Mi8goWqcIH2EXNqq0eMQmSST6Jrqy6wYNiO9m8uUniB9zk8fHcHmjhQwKNpYb5GH
X5DxUaLyFsEImZS1ZfWevRkkw+4HDqKTMRyjc0ZSt5Z2l3Rph2pRKBcqzhv+tH0k
fbAe/06tVMJ2uVCeitt8PP1wlRuYWzr60rm6gXr6JYAGcBTEpW4zKFXwC0Q9GTo4
733nttZ5DP46tWqXws049od4Ho+7wkUuLkngRJ7VxWLnCl+83mj0sFBH12YZaga8
BQhO+WE8uAbehN1ejuFa6nR44ROl2VdoQnWy1HFAR+UjV3cjhYt5dLSC0YfHa3oo
yFx5Vz5wGCnqPec3mItdwEOXHqsD0zC9RWovuwxBYoTdVz5/Bz44jkZPxXxxO0MI
IbP9Gi1GIa2FN046BWfSlKOxUfulQjN7FWwj8IK0moHbl0pbv7cYCa0Z2hL8WfIo
ypD25thhdj/2ylh3SW/xi8D2ry2B/TwRZmQFaHh9yRWLckmk3JawGvqzAiZaIxgY
0Fkl9USy37JMGFzqxe14EXLt+QEbie7yJHLmDxnxqQiC1+33w5f8zgiuKX9LFthf
QMDXvhUsZxWIHtEfv36Si8QadbSVn9J00z23e5IId74x69GzjX+YP+J8V6AgtCGh
o0ZqbunL1r4ngDUPu5umBpx/5eqglGNuoqXc/IBUY6tlzjYZ33jpURFWyeocREEy
nGmVyJN0khuXnH9Vl9RN6gcmvbcpj44RZLWxzTZqisZhWdf4Tog90N5is6lcPzEc
Q72K/C0o2Uv0g1ecqvThXdN5+HWXHYoYncmHWD6bW7d+MuKgrf/zIVsaz2X/yUo9
ooSf7Zntu+buI/Fb7sG28ntSYP8nC4h5RfyJhgClPPmOI2+D+UNtfXWdvXd2Lqk7
s4fDkGcIapHPYiicknHavL/4HmJEFRXccxQcBGWHfvWlwdVIOtPI/6u0c4UR9twi
LKkMLodh38M2LyMhglR+hHlpvg3Vv9IwfwoUMrzRqcfyEx81wq6qugnk9PiMQaCe
IpGbD/Nvpj+WPdB8wUMrUCLKG9rJ+m+QOgmtfszzWbYgkMuVQs/tY2TovQ85cZPq
hmOK8aM/K8J9T1vExIG0l6lBPQGjRP70+N3eoSfS2JMjqbm6fRFLz0IsOoQaVxUN
z6+Evt/5galKtxqwnX9igVtwcaLTv9AkMnH3trUdMfDBaKQJkB3KtC/9XLFvFQ0P
bj0ndOKqVL1/38dxfKxsbd6WKWYJlfGa+oilD7S82K+z/QjoWOCGlLl22pitE5qy
x1V/Vps5A5T5Ua/bM9k8+46CoNx14NVMvur3JuMtjfJUjYdwmP6BTea69WH3v6tn
FNuY6LDKRUiKR7cUW+Zt2g==
`protect END_PROTECTED
