`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ayIvFrFiYFRSsVqYNbh5Spok+cn69uekVr6RuVzOZkyIyKuEl3p7y8XztSEm3iBt
FIFBXQSHI2FlUMIosvvPLjFY/i29TSZ2VoaUJGUPp9u+AhmbA1KKI7TdloTUkOal
hz4rihy+URbA1zSJAdqVDGFgr3Lxl+gOi0kCRvcRsVNrcUk8qk7tE86az2Au1uK1
IM8FSVyeVnCmBKVkQRdluSS3ewidvGJ5VYDdymvtWsEUeemlwAWxnklJw7WKBNz+
0wmbMNad21kPwGji2x5IadCsrR6uHad5yM5SzGTAxLi80rvsJI6d/fXrbNVQDeTE
l1x0/rgfjHQ7P4Aid2eDAg==
`protect END_PROTECTED
