`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b1y8bDoB+HxXgh2kMpb8cyfkgfw2zkrXnO12MomEdRTAocjekxkxWYUFWRiVvY/g
m5dmJ/lhIwnt4nzBfzIl/Ph8P64upu2iVGqrtBDFYvTsUf09rZ8fXTbIhfQi8VVl
v+Q4T40nPFlXsfzehSEN7hMlMeISfE/6rSPDCgMtmbEeFvuzUmHiwRrpi9zkt/Sw
vXUhuDw8cKzfsDB1sMNtZbkJKuN75+7Qct7hNwpkUqVhVVuium8YNAYrOgQR/OHc
NB+JMTZ5MJE8biXF7eC5dP49RoQKZZp1puHLuApt6epc+R724/h1SR13K2gGJdDu
acfnItCqMqqymRVU8SKi2TlgD6EBwTtBAFYPTjYXrDcsX+5MHjoSVADCzrdDk5zq
qnzXu3w6rTqbAKcXJJlfMDT49makt74/xEV9pFJt11PUl42ZZlTnRtYVIucZXQt4
uTADfRH1SL1IrEFrlMmTyZ0wKwBtxTNk+LYwKLuzFsPTQL73gwf3Luq/QLHwYpgq
PejPq+UIHwjyZhlRu855wXicuNckbpExqBpTZamIjqz0kIuSgibNP4U2oY07VdrH
ee9H4K42v0uxQuwV0gviL4FpQfP7HiiGpbREXni68/OjRy0yQmNqcECr+oH1sH+J
OvN1E9xNaD6zvwzg3YlQtg==
`protect END_PROTECTED
