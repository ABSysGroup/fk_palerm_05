`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nP/D5jgO/y5uLhY4bLVBdaQ9LthrgtKIu5F+O8tvQ+NQP54LVk8cHhHwDoQUTYEK
Jyh2rpYRjCivf9NIJ4L0Al3J6xBEQKa6N01Trxpk2cqfm5kddm4KEY4f78YB+qBB
q5slb+seEtYUwUYK42nnXeWparC1AseD5hsHIYvIbdK+Sn3U9tbkkeQaTJrjSa1X
cc4FrS9xVihVrZLra1ILrYNMqRVYexGTy3FILoe0b4XJ2IggIkmDFfTvXqAJWROf
KwEICg6tc/uZUGdlbU2WcqUzMOlCi9qOYkhWZnBJG9WmiInkjXwHlFvrTDRtKMEL
3hAk284FHfrNuadsL+fUNmXyv++2bYFeftv4GkOQmKzFlF6xQ/R+SI1dxAcmWqHp
+imEHIxIsKhGEMGiPAxmlzD183Vr/LmkFDPfNH0g8Ic8n9zPl2bBbKvIpWhYFCK+
Bf8Z8XO20ZFsLWjdlBqazBpfhm7ApuOaYl94qpwkmsTvxtVitsz7LgpYoYK8fQ8J
otG16NezTk7RNeULT/XJ5VjAFYC1Vd1VBfTpo/RrFO4NranLty7i5Nn5kymLfs2x
bjbijFZ0eRVQGi4rviLezCQEgAP9E1dtyYQZo2quNEc7oX8uzsTgSqUzq1CGkTR2
sCVWre7pFUnbD8BmPxC3j02vtbTLMx9d1eVfvqdMO0lDn5secjehM5GSlWtdI/1A
aQg8O6kWubET4I2zLMUp1YQRSfSxL6+jnQkPT6q+zT4JCBXYPD3/5CYeJo4N6Vkl
Po1L4pnl6tiz2OtQGGbQ648aDqWqnHh1xicVpEscZ91t5uQZZ0kYsrhmoFhsNFpu
1KeVkPetmP0fJIWn/PMqeiaO9yWX2/UoOpVJfcoWCDtwYaj2oDaLuSArhpWwTMUB
8tmWLwwJuY+rOuP4t2Ju/Oi5vDZ+xQX5drEHU4CnlS7nDKhS67IEuIC128i99SGp
CdAboal1uSHrtYq3br0Y3GdpAk1gKRdgiq95LG+KBgRFbQArtEjcWoL5QsLDdDjo
`protect END_PROTECTED
