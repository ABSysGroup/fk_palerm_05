`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D80q0wmWePEhaxftb3pvL3Zn9GK1umQn5jVwkzCNv7dHjZeJTrHpGAvWKEyOAwXl
yP3pnI5ENYQO7i+miNFFOSvGANT9unEITAX0fnRxUot12HQ/tNqw1xXQU7Z4yyfx
SLZJMuR/eSSFEh6nClLMt4I1tSlLTWfO5k6wnhesb0tnCNFiZp6z3mpeEwzs6+E7
rMMasEKZ4DgNwNk0jGlT0F9az0tR9mez1VOAsG3L6Ba7/VFwTb8IleXSHj2EeldH
zO7iyp1P5MoQI8d7Tgy5LHtMy8mrffCOm8rIGKfPXDPNzn6krHaDTo0dk56lTId0
`protect END_PROTECTED
