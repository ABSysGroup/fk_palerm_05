`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2VfC+envrfMcfBAJqhnvYh3HTw5kt3iMJVqsbcVC37grQajyX8jih8GAc4vf3zmJ
Ec8A55omf8ZfFY60603SAem3v6vxWlYjScyQR2vymsQ9wm1TLiqIUgXZwWygNdF7
s0oCqDp1e5C4lhP84YXZ6y/EH45LRLiwcjzu9NMERWDqpXLThEeepL6UgJlVqk8p
UnOPav13ptO+sUo1SMZyfbZBoDqaSq+WV/cQtqAv8c0AHWH2C2Y/blHxV7NEaijt
+2NLqsVgcHRiLN62aR9uAQWtOSkj9U3peNWOijqB7lSgpwrZ05ypzZtD4lZqfKfz
ML004BMO4HFzM6ju+k4jGg==
`protect END_PROTECTED
