`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fZIrXdaCZROOYWX0bVTCOpQ0wsiZbv11CWs7egvIZRdsuH3KT09RkGRjLTA6bGFS
BtjOswQkNnrUsOWvOJHOO2z8uij0IvsIcwwQHEsa2NkOelaCBAPbKD1PF3T9+Rgc
C2+wDM4udChz1jKhnu691DpUaPzQyqh8/Uw3zpxbo4Aws29aC6mJU9OihsSPxSkI
yhk0mZBGmJJ7cG+DNgdxEjhiPO5qSaVfCzTw9uiASrfEcvxgaP2AcQkKtWw+xblB
AAll6P08VG+oSRx5GT4qNXoBWj9XLXdGQmHS+5GxYZGcq0n4g+vxFTW27zFMbcs6
f/u1MbI2BVLFM6ktekYAxI25l7AC7a5ujdN94cHz4ZYqLVsibOiaNT8Jj0gPz8xw
ciNOJvCj5d0UFBwFUNBlanknMZy0X9P4TlEpDUrepGKlkKW2jotj/u1zTN7z6P2S
zF9ykcj/YsRmzqpfTY2jX/IH+PQIgX2UBGKasIgu6C1xHmaZRTy9l4PhRKw1caMf
7vDFSWkFzJQvDObD3IhnScsLKj1RNfuwIc/NPLevFyy0Ba6Ixnpg33FNV48xNy7o
9XhCZ24FUXajFILuadUOciQ+VNgTIIj2a43Zn3to9lsb4ihAUiwGUgenQRKhiqS8
WaCjmrT5mHkuzu+Rn8jlewOCdrt/DyBZ0SIyrEZ2UJh0bBgyE8nmN9OKa6dWek8T
7497gKSMRcevyKntTfUDqlBbGiTq1MBpE8NQ0l9o1F9iBQliSxJc3xkQUtafM64E
MJuDSTQV3iIfXVc//uFXn+rtDicHTTcUoZ7v8duqIW/HE6Psl6ZGCWMB16JYXCTv
rlTMKiXXVI1KRQ5tFA+IyfwbmPiu8931i6tGKMpLnpxSiLZa8BIRVTPcpNOHoITz
P90mm6TKTMpvcCr9Q9Af/G9v8vWg1OM1wKHsyVN6ozwnekHKqMAdyqf2bBH39mT0
Xf3bWs1vCDxLkUzJxdjriulLggoKods8min59NeawkO/2kJlAODVq7ryt91JzkvG
zlQlrUODBwWz+fVn0Uk3Z+FpVanxP5TdFHQvkKTXcT2v12TmLIOnhv7N85HA2SmA
PetnP1/YFP5iaT69Vxw1TT/6t2VvgcVyJT5fWaUTpJ9ghgz5TPvRxWv2gBzcX/Mx
UolQkkVuu9CQYO0/lk/4/5PKDu8bbWvVDtxgbFY1x/YVmoXSXskvRqofjzXVPZ4F
ZmnEB7tgUNoFIuB0DtscPA8P0hy4wzC2RdZD07pKOmHWXb3f2ntZqWS7zSyRMy0u
skDW1/dIFF5W5VBSBCI3iaKtMwCQV45gGwNC7Wt5Dd99VSXJNjN3/zWtUVwLEdA2
DwtBrurlR9liYGFpxZ1EyF6chBydinRZqmuDmzOtlzYln52EIaN127v/suGh2mCe
P57g3IfAGwnylQ/CghGGRXPpFE+7UtnWgpe6ZAx1hFWqnSH/FcC7G7zAsPu/Eqws
Dgx3tJApJF4renhM4aFemDnnT7qxkbHt28l4uUlnn57z+LZLEdT1d0hZRlCWjhZu
Iu/c9lUPjsSLVu+0cSjhbb2X7JMMkVCMI3DPcqxMvDDSlxqWxBqhRG/Jo0RI1RGM
X0uF2WYBdP9vRIlV3Hu20JMm59+I0pxtPsyWcdrRa1ZDnOvRjT0aq3rRg5uK/gw9
GqiG3XQZRyRUQHkGo+c7YywGGwK+SLVxraKVjiG+XPX99TuDPqpcaUn6b5nB2e+e
nTTV+/sQrFOH5zGqpX2hAA==
`protect END_PROTECTED
