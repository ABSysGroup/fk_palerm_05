`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fw4F2lqwuoXDOBBvgWqNg/5KakHtmlirzD/ShKGOKdX8JGfviJ1TMuZV0MABIWF6
p4+PikAhrTCvyoH3D+7ouUe4nHlUBDewM2d/f94eEzECbt14cTX59+XhoJrDKaBI
9Lu3Pfi3DrhQqHh15JyIWBCf/XOTbtIUCrJ8Onvv/8Yx6mxHEjDsjZ+AJ8jgbZbQ
14q3hrzXLpnpFqs3lj+5CkekvRYLExrHoIRN3IP+qlJgnSPtT+6NjDyoHewmK0Vk
rNAt+RgvkUOpGxBBy+covBxnSbCTSDc4zgecqeMvW+dLc5hCcfGWw4AAejbCYi3r
EB9lQRK1VuPNMmM3c0ajqw==
`protect END_PROTECTED
