`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YYvPoUUtPV2mfmPY9dfttNmDAxamPBZ8hX47LhZDsfn/zoT4y60NpLYmmedHb4an
6ys+jxjI4p4DpB/hwkyHpjba4kyRC/a71frLxm1sKcrQCgZNZtICyrWyPBF50PKS
B7C3SGF9Fwylj/FcmS9K2VYmX3MODJ0aa2CthexMQg4PVS5QbMRTHc3CwE0p/jEw
V8lkxHcDYMlpilVQnXbroz7cGYaRDLv0KyNqAwFTwhLNFGkWzuTTsHKB4uDXQ7V9
j2H5aDUzJ8tU7gBW5kuA5vcxusN0Rqu/2rwpCsKywIziam4B7NEe9K5bLaHN9ATZ
UdFcgxxTyxmQRcDYORi9tg==
`protect END_PROTECTED
