`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SQVgTw1oJvh5k7/xNEhZy3AcBIouiIf5R+r2rI+raGOPZy0DFFOY0aQ127d/7y3G
KnKuiVoljHKW9SiZcZV8GXJoGcjEJ1t7I6uVtIgOypbYTvVsUgIa8x9OK9fn0Mdt
+fLdOC//a3j0eCLb1bqaexaY9xs5FeOm3vO5w6FDSy008mwwINL3kLP9F1DJ/L2+
2SnKnGCeLF55xdPwIJZ/bndFwjAIMqEtnQo/tUVaYly224gqW3OJi9dErHiN29qh
PGjWkjuIJ4PIm/VwLXY7+ZCDRmEne+9xjbKV0tK7djfafPeZvBvE2VuKimlCGy00
CiD5mnhwRI79V3iMPvg5XGW6r9kd1p8uj21YR/vWFCoLqOM8WazQb53bF2lkokfD
oiZZYr8xy3UVYUCy12tbEVgM20OaIv8+AhBkOnn232vuNUIo44R0vuDKErfPhM27
cQpqBOrEHk3w+Ye19uVehJQd5bAJw1EWm2P0NJQ4Cjm4QPxYhV4/KxMEv6Cy0/Hb
aNsl3rjM4T8ZuFhfjvMvQ+XRBXDC452lE2/B/GWh3j4=
`protect END_PROTECTED
