`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I/YAlYY8BKYiDR+lZM9dn2i0SEQdkMB6ebqAnT4fCo3298FEPKWYjU/c0ZM2GlMq
ebIn8kXeEqWOJ0jzBu88Nd1eSK1/vQHhHiAZst0yVvRYsSYvwdXWj1WQzTKvPywG
+Zb+TjajsCEDlna1UHGqI+hhYYwfYAu1LvqdEc6ZTt0wRoVsEQRu7gDepPTS6pLA
ijmBFPqjDYh/jMnpuNl3cCTEldqZLqaTRtRaEJxEwkNCgre5QjPsUDlh091EGL1A
afvG9LXPbRzoscaeVdeeXhXkuUb1RmlBhu66Vf63SB1bYuY9F6pXXfQ0LzjNroK+
Y3kARZ7cwm8npKqjPeqgS+HFFn/yJEaSer5cq21w7GYA6m+9F+E0kLPq1BBRHGRZ
sehqlOOJvA1nIUVW5saW0dhfR606AKh6hIkO51lRD9kf2rWGIDf+fM1JojeNyBNv
jIhxco198c5wPvoPELCQWO7J6i1qxtOGRJcls5ledON/kHrdRpHupH5mz1qUFzX9
3kGprdW1Q6xb23Fx3oHeTro/LaxNKUQkGkVOuaSEGDCV8+bv0KbkEVfiYvKi8iFD
PBDKUAGXBA2s9XyQNqq4vfEVBqLs5eYsXVGhD2zXdb+warW7qjU66yKkfUAbBzw/
0Erqg3ncx5lvdACJreXlZuRlTp6EJAvNeOWNmkasxOQn5JSXCf4oAGPX280UzCGW
jK6B1lXthT05yA9LTbAOX1ywdXS0Syjosvwfj9y8ZXOIJrcrHH8FAw5Ij4PtJGqJ
i13XBtCVINAR9SrbwfH+N/xyMAdIz6t0mzW83gmQjP/6eXdOu6GrdvONrc9ks3Oh
02PgLqqrx4GFPXM1+sJ1sbcxA/umTu5P1UNaGb+w1xVs+YPVbHFIUCwhWZXpQEwo
`protect END_PROTECTED
