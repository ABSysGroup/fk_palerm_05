`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FUXcED9eU7N2TnflnRQ9kMk2RYLtC65GIBwtSFKVgeixlKLG8hPkJpIhpUM3TCCw
ym8dx0mRayJyDCj4/u+O8jMTUHzlAJu/M9Fn+ZM0JsePMMAeVpi1WORxGYiCTBKU
YUb8Vi5fjJ+/CIFBsDTt0HFmyd6RygvMJbd7RwsqkymcdxysG8ecd/BS1UbondjY
vUn8fAus5kzdW2WdF3Ed2lAIAVGPA6zRbv3Skvbs75CB4O9FjSfgZLZT/soHeIhC
JvCVUevEGllfxIRxa4EC/6NMPjTAjVkkgvt0mL3SfS8OuUJLxkDyPImQcDtIam8j
tiWyN8HAGvd75ciX11nz1DyZbzAQIQjLDcL6CDUc2L1H+sSgPCW/NeI7jpYP3ye9
YakForl9ZaAGxkOJRbmLX8Pj7cTCEug6Cpa9PksCdFvVw14HC+UGlOAlCDSENDVa
Ci9TGYa26WtaFL00mEToVHLknkeNbm3KLMw7S4OD2V+MKRjudjG3PbgIMCydrS/w
MuL8VzJRn3TdBZWxn9q0/bCnfDGenL4NDpKZyZFovOfpysQTDQzCLOXK55zEWTnf
MWvfPYHZF4o1uYkx4LdX5MmaASqZJc69ct1COn7cOKPcMHURGUeWb+jUiRm2t1gR
sCkZcds+2g8arIDbE6BgwzA81jHKP02gS2Ewck8onYU=
`protect END_PROTECTED
