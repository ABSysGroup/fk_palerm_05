`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GApUB8B3A8urHpEnYywdCtHnVXWMVGh4hkTb9nUfV4HQ5R8sCeqaOqZOSImTxoUK
0Ylj1RBwkhaRgLNeZLATTbBjVsmqZPojwYzEzXBaclcMrVzAdALM9GjqNk6sLKt7
u2nWGNOxf88jxjbTObkj3X5cwwNbnnlViDg38OYcgoyC55wWcTfU2LmJ07WdXS1y
WMfNvUjV1fqj0JQ8vPqCU1cQaESxAwytqsZfzZw26ZnlycMi/tEwV7t6pG84bTp8
HCWzsmz0Hb9zbrux5TB64IWzN5UgDyP92xcdiDyBlMD48C1gKFDrUXpcc08x2WCx
C6TRi3ZlnsbAc+a+vO/39w==
`protect END_PROTECTED
