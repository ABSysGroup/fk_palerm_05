`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ac70b/99gir+TunWJK/0SfCxquYvMO2gi8lUMkr0lHwd/km2m+2gKiYAoHeJV/Su
smlwDK9dsfCJaev12w35IS5ma5Z577vfiNX+dH7wGhUrcLxuazG9MiLdLp0zy0Ta
PjTgdJK1kJvzJOyK8VZqbpfs5PVOXyly2az2JkSTgSgLAeeHbou40zCx7C3O2vAk
l0GLaW/uTD+jtlRMwtawxPHwBssEPcFLj4tNu3bjX5pa4FS6l6SY/JpGIoYVsgJY
mXb3TflhjtLCTSM7CG9iUMFi2A2r29yuEheUqdN/Jzm3B1ILttDDqtBfz0d0kQh3
Tnkh301oT5tDuJLKenf/ZcowQoT2a1dnP1NrYlHCZTYYJ23PFgcHuTTiYuBdgvfO
0QeRFwFT//mKq7Qplie2PNDMz8krqQ1j8BVvctycy4Ibe56wX2vFc9P8ZpTDQMWY
nXDbLDHa4OmZ2+r69WQtB/1zZhZJWl73IsTZvyvokBW9g89bydZCtGjXW5Tgrrgs
aJqdWp7Qy/Lfozoc0Rtxa6MOaznYbzNBsedQ8hJv4v5lMz4+sJMY3qiG7kcrZNZJ
60E+EmA+klWsOQhcuEnX0WObCjDSF3F8lqiDw4meGhIOKFIOCPrhlPt49nz6Acc9
QpdYqBbWT4HKcrPmzePP9WmwRjcgyS94btQ+SpyYYpU6k3akAjtY4Y9COg6KAjjD
/5dxALrnQ6syvmIuZMisbinhExYs+j7U4Cz0gfKmtmKA1pbfSXY/uchfWGSlOw5U
0Z1fqzxIx2a2UeQxYVBZCR6+tp4KppNRkeDA/0QHHIwrb1ddpPFoZdYqA92C2PRC
Ha31BEv7wVlkg1p5tKcy17MA8EhDpxmKryfUPn5j3Nx1E+ZeCfPbIDOdQk2icQxm
E+4zqa+1nR4XYeWFiXwAfOUQpGESEYGONSx6iKK/1MUlcjrORiC2JFk+2hkSb6RY
sG66xP9GNDjearI4PIaNf5S2C0Eg9XgHJcxJktWASoQTW2wPnwQLTDX8DFHbXECW
v77hSqsqjbQkFqd2I96ItA/GoqI1YKRPOGSxyqDsdiVnVxgOtCTtjEFcA1uulIiL
pe/Ew6r53iSWgJSAfafKLsLhXHaAK/D2hyATnczeLnq5ZVvNmSZWmaKed1o+xrsf
/RVRNdbOWmYnT48ZhfsStDIsUwam8tfABBXzkNYAd4cVGIEXnJJ22S/MLdx0Pa/Z
gq+DscaaB9UFfiH0gtJHrAkpdiPpQeUyzhTKu66U7DhpQweqRu4RrYvlNHUdXbAe
E4XTUSoRg0qP5mcT7chYbntqKh00JpV+4SSkQ3uZDuGp/Ulz/3UnNKyPoUrTKXQW
Q/OhmMKzP3HtWki6tYxM8w==
`protect END_PROTECTED
