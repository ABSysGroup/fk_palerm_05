`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T/8yFV0Bf/r5kNIJdusHJF7ytB8yyKq05pfb9XlxLXrXU5WrvPVCnfnh6AYE3plJ
b2rbUbaAud3d6ymeHg1HUjR6SpZMkpVanvYdpmSUSj5O+hIx1+dvDnT3WiwA9CLC
SdUmp9hQDpdrz79KmltgcY+Opb9Fah5kzqpXrtbjIi7r9r1BuOVeiq3twshRtRlW
nDQsejSMkhjuvT4CCx0zNyAShgbZhS0AKSXbY9C2NnIVJR2+rYDVxTKE4S1HlmlE
aqXxDW8pY20MCV16Y2OgJPfP7EbKV37wp+2N4522NTKMwArge+ln8TPLgSdLiOEu
5+AKhFOfv6Slr9WStjjTVAaEensO9N5FV3GueI23Pyq9cZRHbAwhL9qs9i64q/8G
sUFIW2Hn+7HcAXNWz/R30INVA/6ERbrdkuP9QKuNTIQxB/MI6Yk0BBT32tRD6bVZ
4h1nmxNWR61/DTcarqaoGC++nAGsFmToFvC3+/NFh+HafraaxknnnYUNKy/qTURU
WkS5i7ghrBdY4Yz1IoUsvm1+Zb7HPBlpbGFrmvNsjJQ3bseLZ8EP1sTOsC+RiXz/
N5DRgyH8elpxx0PI56+86OufD5nL3G0g9RO9L8GumDk=
`protect END_PROTECTED
