`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q551stg7meEymFEW+U3O1irZ0s1B1kdC4fytvY3hDm0/bq99PSrNimdN2eFp3Bk2
lnc7vNCC6X8mKIq/O7ZauWFkYy1bAabGLvWoiMzOAD1NRxQdEbOh1mqG0O6HDePD
skAuTzGBfb8oxGZh7oTVFiFAvx2AMNKdgx9G0+//PDQgrewXTBK8L48KPhkXKM9n
Gnk6W9nOdo1HapcflIWqrM6we7XgRjYEISYUZIyuxNQXCDpGsDPv64wVXPFHjlQy
uo50pyKxaqbR7uijvWCUj+c0lv/3auSkXDDoFUgojpqU/iUw0bc7SxRrwtl9ejaC
n5knBCt3QF9gK5JJMloHSSKDZDUPW6kBI10J7tB+lM1bZzbHKlzzNptLLxq2xUOF
QL4AsXUZBmnDj2NfzOdBlR+VjEM9BAHpFRnWOxpv0yXfI2v+j5asg/AV7zfoiQpm
ZR5QXO7+SkTB2UXjr2BCRn8hRdctu2zGAv+TNCGlT0TYz7RMRqB2oiJYnzgI6oDG
uRz3NhX4s7mWIZ8ate6lgvVh2ZzykyLaQlkOVv1Thct6FG/RtN2ZF4/i5K9kMzE1
/RLim6NeAV4+pVe3INoeHZ3LnU8BBRNB3lwIU4Jv5TcT/YA57e/OARiwGpbKJOas
+aaomq09s0kRimVgrTi5bTBBuf1sbXclHBxXcbrQqw5gWIWm2SRsgQ6PifJETCqp
wt5u3jfrUhBvQkMWeOwtiZFSp5Qahvd8ro81rOlBxZvD992XFVv7EqkYCadjgKu/
hrB5xPufdaFlEbh2r9D/Yb05RnfM1FjLb2dCwzyV++VQ3jkvmkmElVCmRoldhTRT
QUyjnWSCXrGEga1285Rff2WReAFAK3fgqEy7JfNsXLHx80dUC24MbphX3hCtwPiQ
6i2UHTr5z4rD+MPaPb3XQcSR2RYEnz9vN+/BgamQmRsOKj/f6CZqmjuKX6vK2MgP
xtMbTHcLg9e5wbgMdaAGcKeKMK0cbUPROF+SgvYHrlrWkknzFnUOnqyg0n8lkN3J
TVs87T7lBK5WcXkjp0xdUrvTvjVKmXh4U5DMGSp3MBmoCNXKSmkJPGgNljwvHUEw
zL9LdmUFHou0X0jw85Y32UBRg8bjEDqCvF4kN5y6r8Cd+UeJF4lBW+0ozrsmxqhK
372oo/D9dVALRNWpCnNSwOjfPYwWoeoeEjPLlY4bAW1pqs6t+po12MZ4HsvxH5Mc
`protect END_PROTECTED
