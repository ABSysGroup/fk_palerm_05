`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wWyk1hXyhAIm33B0wsRt3n8MhTAhxmc4EXp+U4i/BCLWGG2K1Mg4WerNWVUdVd1p
tzq1HaMqpOPw+VQZ7j2ccK15IOWHUYbyj94Nj56Z1va0NyIBzaGDhwjqWs0P8x2t
/L2mWHVr+78CIRRwekur9H/8d1+uuMtlG961m4pjcx2PsG0MQErhBXw1/zAXcubV
0v5CwTtZ3G5Sb1or+0FmYfrjb5AypUZWsv029csx0lJDoHujLe16+HxPjpSrc/Om
4K3MdJ+0Pr5ySX9CeLCFKH74pSINDQztBFuX2vzrCMOL3Ya6wTORDWRDZWTNhjjU
62qJn9mrfO7jJ6vlK5yhjHejG3GgH4AorXg+fdKGhl6a6gu7h+ZVtw/I4+uFp+Bi
4r/iqT3lLC2lkB9l6QwJTYevqNQM9ou6DU0UbMGBm+ZDdGtUVyn7a3btf6Azw/P+
CJWDgzZ9aTIeMWgMscdPeHGWTo5ff0knShIbTD1ywePaSvMd/sb8STsVaAC57Thr
8lknl7c3koj313/AGwCcXmZELlZ0Pe0mOTE7NBVgdSy1shCfKnneTkO4D7U1sMPe
7BBpMgccAaqZhdEokb/gq93uywsZwFXPBtbHwObLWnSTKz/RXZxHZX3+voAtsrAH
yR9HHE9fwJhcl8plnRLIml1pqJJ0qmcUC+IyBj/VDhlORSpW8YcHDF7iAObbbYZq
+ag6FCOgk6JzqLz2YpGzi57rIcQaj0riWwDsxzx1EYouRhBouMyLEZwtlaSrGrMm
xdW31pENzx4oMrXel/f3WL89aDIiMQQNEQd+45spj6VxikmzgZBE5nAVCCx+CwBk
E16QbVDQFT65k75E1uGaFX2M4IU4W1Dw01hRakK1sBifRK1OfXjxdR27grUO5naL
DggBrcmpylUw7kSHphp3fq4rbrVYnEEjlyUyn6cyjdLcfLR9Ds5hEoGnraVveJ2C
04clkc6HoBYOhrHdqMPQIwJIMr13bBXkbYiyi0IFDchT0lrVR4uKwHOTKjwCEGEt
kMWNCzhRMGwokAjnKyo4dsElZJVY49/GYDDBf6qeXVzoNzXhORoQyHlmoKshgdbv
X1askWlY1N6PpG0kU7f+rgf852IFvrVb/3JGlyoXNGg+cf1d8HOe449Q73aDt2zA
Hi2DLB0ceYVtfQqBU9FLdqL/HOphbnfFVxmWPLM80T5IhH7JZEPVD83VGZryrJoL
Lud7WTCw0YoivcEi0MCByynq6fT8EnHmMOh4jQpFnq28ptXhKrsf1LXQJpkVOBcY
5VBU24VNoMSYtm7NY3pzfCE2bj+21hfvLk+8+VnHGwSTBFpGImmfLBh2OpJ8TsqC
bzJd6AGOwjs/i62yghKJXcB8+7yBFMku1hLq6wfzsY82wbhWcszSkbcR8KNG2Gu5
2T/fbEMEa4CeiXm12lJZKuEF9Dag81ouJ6+BtB6WWK5defOLVnQPDNf8dHOExbRU
yxJlOTT9ibWBfi1TNRX+Vs2/3Q5WsiWwIVbEys4yZCd4r8IGSR57nPGcPqV/g42F
GTIqu/rgloMMaafBxX6XphwfpBZz8WjfYC6/5rYBIwA802OgsMdWbWhHY8tqgCGz
qcZYyt93Wfpo1ZLTAEaoLYnYJIqF4BeLh7IOLFIC/EoereisG8KIFbOuLPrREyft
spDUpKKUnaKo+w7cb9cMdhWiFYrM2rGZ+eQo/+eiQL3wX9fHtul7pmH+jL0+VWwM
TX3EnyOJpxZBTC8Hj5Hh02HVKzxkxXHIgqtfSX/Ib8fyoaFrTRdf2DO7JH3IEuHE
L0a4fRUZkKYhtcOzC00WayR707h125Cs/bV0lEbepVhC9B9/ff84GEyfQP8vFaZk
mboWWd4Abxd7FdSXUT2qUuMrbR27BhWjhQcaRuICNCvVbH7lvmcjIv+9XWlB65c8
+rQ+Yj6Q984HweTccF159krEXWVLs2vUvwjDriLGwrU1hGzyHRUCBM6sXKM8pGIk
OOQVnMslc5T/4ckIpLZgXR6apQtETR5Sj+METmM638ukzbGOlkbYD9RFtRwoU4cv
sQWWP8DhD7I1GkvB98HBOOoleVeIPuV6Ol8UfQxrSqXxGd3pF3BoYYCkgFfhrK3H
Wj35zXipkezdbL4fG9visfhjs5JXPYhg+uGGeD+5LcWnDdTQU3HfUtU2Nmn213sy
a9N34kzfSbjInzgyyn5HjnwwuJJh54H0r7toQinGzKzVqCmwQ3843XPxqVazFhPe
p9JBwbGDS2z7mHcllmM7kwrD5pdgKTuwJv/OycR4qV4/cixi9VswQHwcrcwiHze8
9obuym/w8+5NALnA82/gNuP8cQIYSNMoU3CpfKkhB7WhJRHTyYOM7W0LX39Uh1G/
jwnUi2mknJNxfYTTi1IBm1astDwnvgowZx0ricjeJM2XgiyBPGMKx+gFL7ipA3IP
0y1P+ERM0GmpJ8Hg6ifkVSjw4bQle8aSG8+JSzrzWDFbwhp7yWvm4zsw4GOw8iKd
rlLsbRh15+HZUL2jp7qGOykF36lbkSq3y0RhW78ZrQOmGllCBUcvHWaCYRbFg1GV
CMjLK4uMH7ZnRN7CcZ3n2i6MzN0XR8w18r00HpeXHl5j/qyVCyuOQ8jqcRmghpZ7
wSWTRZ2lhq/Gdquu3p8IuvXzF43Q0YSL1UprLwndIkMtvtfbur1wHeeJSO/SyUHs
VeKxwsfLLq/nX558Mkeuacnisre7fxqbwjVOqBJIXlA1/FAw8/ayRJXFdOEzKOp5
AAAd/uOhTBn5QdlQFcDjO8MNx71bAQ1uJNwWI0Y+iQ0Art1vLxweEk2sFqKl5KkW
gFpVj2rEsytOnb/IeD7BlZujwnLTtEf4bHq/EZ+YWgzU/O6CEu3QuvUV8vD59rDO
bKIT196+AcFV6xwVjtuWHEyhpgq++DmPU4+IhGEccpyeMlMQYO0eTi93r5YRG2gU
1v2FAf7of594X8f2BTTos+Yj3f87vePw1yorjp7wRAUEK0PFNL3sFCVNC/UchJIT
7hHnOvuoZP/jn4GxNwv+raAeVGn4avneNehTB6dMb5/bluNz4LsEVgnY7whopYvg
NSqget41ngQdxnyw415Fqr0nIsu5CUrGgtCi6q4DzpOxddTl8SLpCk0GR5Oyo3sq
BGE3fNKe8RC4ySSxx94hWVrYk8kEOaY4w3Eb55Xxf4PqC43AX8ReYQS9bnb5ERbo
8zW6lflTHC63lQILiTrijsWlKFH0CzZYSBuZGnex0/ZVZqkXMbY7K+7DcrC//MfT
vJuOmw8tCQtOe5ai5K7Qgl5AhhWbhv9PmvhkvWnLP5QGasw7uudxheLrPU/3B6sh
rl35J430a+vCzHDK02uZQFLpaVRxHL4cpYJR+X/JbNG75i2lLIuGaCRRgCNtPDMm
4c62EzBEmbW0YEcHsKkeruXz7ifvlLQv7mar7fgX3pMSgUGpFIwGq/IcCgJJ2IX/
PGzU/A1yw32DOaeUhSdWq4KBUblROc1X0JuGKKGPWvtC4zHYcqe+YD1rvkEm1EQn
dYJF0bTtsgk1dapPalxgmb5UJk52F0nOwXjbQj2uHQVK5dTbVz34pfX5PXNHxFVu
1mv0rAatMNkdrhD1jJFR2GeEZ55Ej9K9+IFdSqR70FY2WSsu13hxmJiaN/AhDIFj
gOkADdAmVLBx/akajkV8eKO0MUJqFj3ZrX6x+YsROoLTBpP7gfUqGm2N8g1zL3Zr
cjnsbLOR37InX0K4hodVsSUU7KQWGvtkj8b1Tc0tsgBi5+sRG0QgURyFNE88Oswm
t+2hJZX+Ss3rXxHW6mgJEYE5gooSfCjBUbuHHfNFqncL/1Gxr2pfbgefUVjygCyH
789qhbn34BZ/RdFD/RC8ujLXdkC+feJPnLnQVHXP+v+epJP5zEwkHvHL3+kYUo50
TekUs3yLxTEE+0JVnAhNdUBsfq7DqpLZWWrnFc1/cRC331wmzGMG6kRQ0qAd7HU/
eHeqGTZGVcYHS4bYH/9bKQgKfjDCKkCxC9oQ37QI71bj9xFVUtLvP4+aqFi/NZQR
T+OKE+s57xqzcyGbj1dor9qOvV7NgdkhnVoTJW8ZitDaslSlGM9ZLMkGD6UmLn14
OHXMFVG3rsXfBetWVWHs3wzlPayWFcytPHmuuygu2VaYqDiHtTxMVAUAYCf2O0at
qiZz3cXlbqq9Lu7NUDRADiA/Tq7XSby6I49DnakQUemOwezxw71QC6ZpZEOK/d0J
PfhKlXKUM+Ujir8U9oHl8cBMs6pF1R95aroT0NmWpYFLXM1qoXmPz0qkObIMQdi0
aRJCFCJTd7Um4uW2Kg40tKLNyxVbvdAnDuskzbeMRML9CwyB3XJCKBMVWPZGtA20
AZ+csBEea9TjuSNyO8JlTj5rOWKBSMNFNuC+2daXnd/ngyERJZWsfOvX28ZuuWxE
skBwVrVu9VKW8q/pYWLUnB3zdg+ACE6oozlt5wh6DHFUSKu4WnUoJWpCmCl17QWQ
1kZscqM3BxFkSUW9KKNDgyq+vjSjd4X9n1uM08t2OqxrObjWB7uiohBV2h4IXBtL
UMMIfSJBwsgw7fvfIVXeYuJOyHW4Dhul0C5O3bsOImKMb2tWOaUavyuBu18OHFW5
ofqHVc6B0NnbY68CzQxACoWCBh9Su0rcrupKEH+2CdUOYRUjcTb1c0u+RX4zAoOx
B41NrFhG06bjA0ytddT7L342YbBK8EqcPdyW/utuRpk+5pi5578s7e+l24XOsEZR
GnTOaBjE0jBTdAO6/gS3SevWUMjiO40RO+B+zSaBEoyWDoEVcE54F5mqzksKWNuj
0GjBbgVkhK82KDYgcC9FWnrYFMwcY49cdxz/VJA1iuLAWIzughzWahJXRt8m0e9j
t/Ku+bSw3v8zwvf89WpYXCJRWh5M7XpAdNvKRelHwcV7nG763gxsVzq7Z5mPxA+V
6uImwev2pWwq9KqdwUbSIKf5xl+3pq02Jd85Qi75GWhepomdZTM6doH5TEIIeEyO
B5bASrXcw3B6ISeM4/6HMllUIxg+QTt142TVGWxTE1mkbtmsQvxABsD8NaLC/Is6
nahlXM9xebr/pQ+/mghl7eVocBKhlm3ddBJA6OjjEXeOi3JuXub7D1L6bdUyAZwa
g6zgx9foPeHefs9xwmbrw8lkBmGsZ4R7Ey0qKyBY9xEM4dPlOohxiqEwyqK45da2
zfd8P1z8Xr4ZfggppZnNPlVoBHUU7TioPjfKabVgFi9T78TqgiP32aWDk/gyM3xf
xhdUoQO7XFPBeTLXAexXOtiUeJm+/jf10GLOcNrXwes7r4sK588UlFjqrsyqoN4M
S0YBwfvlT7dXhWI+CCIC6alb0fd0+pyndMdT7mZCjGvlI41nZepLtib+c9q/1Gt5
Q7bcKKjV1aJgV3PGzHRQtotSs/iJVEIG/oqWEc7e2fhBgAT/gTDAGptSpbJrJpyk
qtdWJdmDqrPd30jNPxHQIfNnXH+phHed4zu2vx03KXZzFwaSV8xExgQX9UvCgsJh
HQ7NpPbJcO/HmgiOk/8BAmTmCn7O7sD+KYVO+HKUyaIwNkKJdBSPa60l5TEHaRc/
1MG0tIuwt+G/ksQkMyJiz2AFGcS5e2v0mW2mGn+IMgkYCENFavZ5YQAPragegvK5
6C8DVINc46O6IvYVp8/oJowMG/IXTZfroll0zw8he5w1xAH6zGPZk5qep19q0qRt
z7psp7wvU/d381vSsko4+dzv6GNOD35LFmBZOcNlDty3yEj90j1+FUUUGJXdolBK
W8rvXVKsgOAM5AcDha00Vmg0Y30L5lBnjlP8toU8fNbYXm1vpIN+G+08+fmDVsr+
5ZzqelLbkQenYH555baTNiHpIp1/xCFmi3nhqmqMrJbK4ho2HIGkQPo4Z7M+HBcG
EY1c14O6/9iyWsgqegndK3qtoxJk+hWo5sglQRM5ecVbLFz88Q2l4WzALfqK12oh
1ZajWvuFy0fWnur5+oRrbVRbQOVcRJiemOj6AxaXkU0HA8o0VXf+Dw6xf9GgcgAE
851LvqaWfXu4gWQG/VZmdt5E6T5fHg3YchrS1ZSEUSPAZb0gapYIudg0MeexbAom
zD97DHvg0iZeR5klkEB0TSsUb86WBaJe9kguow/kY5Vubx7TA79E9razxtq/14DI
mNn1Id+tGHQOtpRPWNq+wCSvynUvOM9w9jIO2IP+HshZfYVvjzV74QglFuQZL4Gl
XILXLfMepq3/b+PZBQR9x7j5Z6XoGneym6OOrAA4xPoDj5dOMBC7rMzVnOmOFBPy
1EdesGlYdg81DJ3XFVf1NHct0tPIZaqMrm/73qNMN/snZVFNEV/GLsclOB46KVW4
4mua/zGn1n5QDKKl4JHPp3eQjr9SGrZP0hVDvaSb+v5YxokcJcsAjkednJGNpe3f
MgiYp864kIhlW450ywlRf4q2jrVLzeFQb9NyJSh37eFxSdcWkMiXL+yNCM+8EhdV
930zXNRp31TM7ls5y6zmRINRZb9zAlQ2EmvHqz/0zoulUxQM1PzuH1AK9v1nkWLN
JIPu66BVW82RjWNvto8SY2famSkazwZM8ncthL+aC+NTatmrTXN0cL7405i+M7Vm
u3wcxSQIhJU/KEs7OjVzvhUtHpCTZdwRnXcDvaEMMuG4PYYk6crhWr4MFt6L2OiW
gllDo3TW2L1HWfPhY5L+u70RoQdZJXat+vKPWyhSSxVsRjSeLTHnbPqkVrZFGjrv
4U3joqeUC8lYwkG9ZUSxyzxj7bfHfgr3kKcNp8esZTgrnLBoWMh2/ri0dasbB393
CbLB+DWmfzPptLhC6LJghdY5Nm6qVXAGDf5JhWyy3PHMl3q+03v4EO47/4nGr11K
J6nxN2tWKg0JrU/4JMQYdeLlVKCx3pRZK8+TBC4gyL2Dhr4LJb4L28VX3w4ohYEx
7wgil1xE4L1snSYWtTyF6GDpuLtMHb6nEh6sJdZZhsT5tBL6N7e3lIUmZj+HRhVw
Hhbwr1lqGUAaypexDD/5oIrDj4FMf+lRTBOaGzEeBm7sowJ1+k20cWVfL9NHL91K
69H6JJ8xrt9ZLc0Uiupk5JXtPVWG3HcXwHAZj3rLVf306JdIzVScbKGVg2bdX7kW
a37MR7QKKAa+Rw1cLr/G+zbjHxLINeBG3AMbatPwUgCX+KIc99ykQRnxHB4peogs
BO30UrlzgG/IijTSyXLuTtcbP7LsPl8IDuDQ+C2LZiZJm93PAi8pjm6+JuO/7cOE
CcolNdwGkoStdZmE1wPEuCGbGhYEPqtuUoqNq2607AER7PztXUK7KmOf9LEWB1mt
5I+KvCnax5JOzqPRYaTdy4ibmzM2cJ1QGBPwVXdLDJNdPeP45aZKjonXtHhU+IP0
0OVlkgNzyztcMIjzRxNpwFOlj8kxMryc2na9/o7+RZh2pfvL8YwRd6AFtoY/Sk/I
lCtUQL20UwzsVgAhE/xj55I7jUnU/BOvDvwBm3Msb+6bB2HhKg5Aa2QG++CF1h0S
nO7s1t5sFC0SLPVHC9Ybq6af2ndxH25jXnV+dkWx2H36rsGV9RLv+DLFXG6L7wzv
5w63klBDBuvcGXzLvzw83+dO2H/b3ccJQ+E25wnUsHfXUKVjeqZvIQRpg4ZiXWoG
umEY3auq8Jq620Xvm1sGIQ3j5H0rJOnX342BVsVcPIAtYR+wSHkS+//yT8PKQyp8
JZgN3YFf3HSEZATNpHopw6ZAtWg7IwbTq3mnY94AoCyjyCu3NLhZflK5zAthQxiG
HPreZq9bELsir9DXoFTtGEx9zFZ02p0uSc4L1njVTvOTH9Jyt8dJNc5HPiSSIH2n
oF+mfuWoFHac5J2ZZoi7dgt+yGT649hq87jVYDZ0dLLDeHoLnzY/8l9JG/+cZD6o
tq49gPAbt7vEgQ4aAY2Sua73u604YOXUI+UcHZnOpTkFDPKFBbSBS5idXrIuWib0
wVv7BGtQLQy5bMT43vT08dWmBOGfoGlIE9RfYEpgf/OmbC0vc0TkEvw8PXJ2ubJ1
uIG1T8xiwtkHCtIQuoVsQjGM6bPEvv6eag6Uh4wRODhJSsm0oExkJdTORUNkc+xb
6yPUPettHnx90JA0eiYKUumAVSTyxGAayi9crCJ7hUyUT2bNxQ3EQVhusQBOGrer
PyxIOzDw5zJGAA/gCLNI0scyCV/iKEw1/JgG/llQeXvykBJPMzjREMvrpK+3Pl8t
tS620aDuz13zm475hAANnRXV5Zpr3YpYyHo2FaGOTxmHUPCmFy74VZkaM2xMDtO8
mOFcDqB1odZfAvnwVgLhIEsPNlnyxeWCJ6T0PYmDyHEkAvMSOPkRun2wWts/aVi/
8oqC/JBCcynHgkWaADyO6sU44h1wYhdN+78qmxNU/4sOZT5LjmsgENrlRxg5zJaA
lKB/OwUzVkLya0O8xCM4444lESdmU+9CV7/vSAeoAUdRL20fuslTIDF6CQLS/LWA
CwEvfqg1FjDCRJEGf25lFV5nTKK0D6Lb1Hh0L42OusF5wMRmbBffrqapB6AL7yOy
29ILxxmrfEYLekge3tcSbZwp9rjrXLVVLGkbMw5KHFBskpQSajkJ7joM1m/TPDtg
+5k322tQJpSmWrYjhNX+EKCAGgpuVHfmp364hkFK2X26YXKiF0DY5YbdAeZYgwrA
idT2yGcdUozsSjWPZG95NC1WmcGBVn6OEUoamGJI7RFjC9jJi2XWtPpIyb7PiZ0P
BaavCO99Obt4BP2W1i+yLg9HHEfcFNcEhlc9rLk+ZyAv+EKLDQfe0XWAwIugpBAp
JjR3Gwk3YzMtm98YNZUa3BxdOplum4mO+eCwb/iaU5Etpg9HDlmhVSjQ2WFc6emU
K6TlrtbzSvD98a5mBJT+B0fAL1OSRfReOFs/KCTHkNn6wQq0hIwaUFyTUHnQKZT0
EKAg2pS2qhc2bjyOhiZfRpPJpJuCMfP5ayeIwM93H0smYCp3KJHF5F+Stb7jTUrv
OhChUhoHxlULeOy86gf8iHNElqEiZbgEFL4myp3iXFa8WwFTSFkYZGb5WH8cxQXJ
8PUUmMpsUIJgcjHfFFCJXD/EP1mDEHSrgoWsM3pGHfYP3/YP08t8XO2UnnskIka0
JT63We4BuUhUzkn8yWtQ+9w46oDYZ3BHthtoubRmmFod90KnTMlhZKKar7W6FvPg
kQOTIXgvJBdl1YEcWhxp5DDTOYd/YyYKgisblDlDOwWR79pqKBsJLQJWt+Sp9pCt
plE2GS4998TrqUJJmvYRO9avGx5j34fu9iyy7m8KA/56tNuXpVv6FooRO+fdDjVG
iX+sH95DYiBLXLyHZvALHJF8f6yuc+xwCmQpp2MbR44SrewMInJmDCo1jjyPVhuv
qE05ujp+UjZQTMRx+GFcIHPCboW9xdEPS5/WO+cYKi3lK9Q+Y1zSXBkm+EbooBHo
ky1Xyno6CxoxCxozPLrvorm+okA4A6QPCRjxjTlGw/e9vWfY/+Ipn2h8Dr8XhyrD
vM3t4TgiEJyFUOQVzFb40weKwrZNzSCpBEtQOy+qKve4BXUZ+hwLAcx5MRSaxkR0
UeF6tA6UrLI8G6TZwoAhSA91afh13vhxvsGYWCGQjcSXM30R2WdOCIrB5hSwxzrV
EuNHdUgyY7Agf6RtNVGmfVUfcC3tLKwNPXrzOyFUFvRx3W+ADBe57bOkD2lyRVqz
tKXnEz1r/i1wScKj7uOzmzfJrT9ufryNN4gf7vo0VkypIFSdDfjjBIfRAMkpyeh9
55Y9tBf3c+gml3vsVWDbA7C+90aW/y9/0fENt0h6vHeA1UCC0ZsHqZal0wzRyVuY
Bkk5ToXzW7eGmP8AvORN3Prz245rU6RYmKxkqJpjuiyM7HHlHweut5I/7OrQkzLh
scHLWTDG4An6UtEYjiaACDv0d8rbqhXwZPUN+zL20ikF4jIyHOUpoASWkGHcRNmF
zk5eQvBUu3Vf+k+3EIgvUjyIYVFLVGhfN9NyqiRQEzuPQrDF1UmQjcf8TkvvZcDV
WwcuSB8iXFsnPsVetHh6WMfoYRQPEyII5wbqAOvCpiZRSV8m0Y7sgN0zOr/Pz9Dv
CAXoxzE2zpoScVVa42/P1Fgk5Kf+z2YBWspR1pqQzO2KRc0bTri6CnKW/NPFOXur
1a6ZB82qDXcm3tnAfNfYexiwAAUkXagWE1NSIzazKrXv3XqdfyFzEmpaUQ50NdrF
WTRkamFe2p/Jse8n5fC/UQo4W3jCTbMCXnG4EsV48xsrMYe4fgTy2pZxLJhkMeI+
J9kZJtuhodvuxhBr7JwNqpv1y1mtmHaJkuhNUEuN2VXCYO/LObIAjsBGCy+EiXAI
VUWqXceZp5I2DTMPe85PdbX5YFcU2AHph58ZeGoVV8CAPZb5jmBfJNA1GNAgFcdx
ImStppx8T4ox5b5Cg4ctzfLb/8dGMCUCNTwadJkUUO23YFeTL6AVu7oKjg0Guh81
F9qqkBmIMerRbSGBnVQPWCIe7eSdGLV3pvkN2it2Rp1LWZzQP7blSkTk81TFh+Pf
PzW1kwt7el3BfVRd78QIicJrfUFmUW7YDsgymGYnbbmQQSa/8hToey2GUvAN+3rb
MYlpiJe9W/dYzDjfSZxAD9GYWtc/qaQNyJmVQ0hnU47JikZdjc8ShHXPzsEH8Asl
f1K3ncU+/YQrNZoFi8ApjTAqKfFWgrjDHyPsQJjqjBFs6ZH+oKt1t9OIXmFVu360
PbXXmA1DjsGgC+Ayqu43eCb38sDSlb2bLLEdfA5XSUUTuoDm8HkeHZJaivz45Hez
uCGOT7gAMAhZ578sj5WoM8sH+0Y0LwdIo8NrcPXgz0JDqWGe+Ut6DMxSgySwjblF
IAqlGztK98MnNtPzSDGKCvxAC3BLK12S6dn/PvQmjtPPh9XU/eukxrkhrzowvDxm
rD02SEBjTw+8K8Nn0qXSG955zdR0CQUa9RfxvzkrmQzrSBeA8rjXPPX4irByZPDH
bqyMWF9Kcq1UguxcFH1iHMQUcflca4/OCU/mpdVRCCqpGDnyojkIBVMoZo7fuY8o
Uq3Zqci0Bp+KGhTIYdkrhE1SG03Y9MdJtaWjnDg1Ec5kiAzFCz8Kagrj95jgvI2E
cTMEsRPW3bRV/BBXztwTvJYimHZjlVctSd5On2K37FyCmbbVZgmZp2C2QqX2Oy87
7uowGrzd+f/QYTZzhZPThAJL8v1rM0llXvbMGNlpDfHpdMuWr2EoFqvGlUzLcmgv
Pr3hhyiIXy2JF0rLH4zBnhtTC8vMQxii9JDmgfXx6IlDLdGwV2zgY9vqgE28iPlX
yJhpDFM2LvxNLVTtENIltMZG47z/WFl4Jl+/tXDlep9EH+9HiM02WLizdAmELmLa
D3HEhxeiqfgUwqNJXJFTrNkdMIUkCAxwQvaM3HA4fPrwIxAbfw/vE6gLkLrrp/iB
ZpXnO7n2ddvNJ8tzaxWoW2/b0tKQ0clBL0Scro9G0uGTlByWpPXprVepgbRKv7GH
zD8FQrUUoBsFLVUmJWYZXLXpn/PowVMk++X3tVuUWIE9gPUX0HMkLMpaD5QMTVLE
RW0ppiKbBfDNSrh1wrY4vSDurhKiIJjgBrxOFdHAdO56KxstVn/HeXRFxMuZ1X5q
Re+BU65taHt/dt3CTcYSy0GZd0PK1Nj9TnpTSkn4b5glKa1kfuUZULSnnA8PyV9S
SvQicjvQm8pH4V/JUzzaigOmot0KEBwwNbMB4HzoICa3yGl8SUU/iYIL6L2daf5g
hKHoEj4GhsxnmQImqMpCQQ4kfJCsAeKliLm8DSvJeiaaWe66puiiL95Vv96JImKL
Kx4quGIleIfzGJFAkfzx/doCRFyGP34fUF0H3o1HDn+qCKTN/7WN2pnEkw4138nM
zzhsYIqB4xB5P9If2Z09cqSmWaDSCeHNK2sY+/xP8+Z6lkJppUTeVzyR4jTJaJbI
7L1ywUqNK2CN+G498WTSm9iDMJVjpFnnzh0t3h0f3gxcvSlg5pt4ARAE6lmJ4rRp
nPCsWLNxMsi96W+aj0zQT9My1p1zX4sKei6ZGj4Y7ZVlZr0jlL8sqjuBFN1FjtuM
sqxhvO9G5nJWpCNCjx448Esm+aFKvVrdB7NU4/qQ6yNC+pg9bkngUkgWe5an9tuV
T3yhgE7TmQWdVAwGTL/L5ON7f0wSXKkV12XS1/9aBbCEMcmCn5/kds261/5yAuS4
jg8cP6Y3cDs9WTE9UIKhSTQcHFj5Ve7bQYlux1BZjrX1f1DxNYdp/gpi75hbn8yH
h4Du/jZn0mT1zRJTqiWSK3TU++fpR15Kdgjg0sxwhO/wC5/ctOizE3jo44MfybA2
3PSuMYwiiQkJdt9Yh9hdNB94SraF3LXdOcMh8DZ44J1/LWYHjDS3sNRg2j9CrU9+
DtzTkuhHNp7zzMye69RBmVnCj+VBMc1gHB+of2ZAvvaXUdJMzAN++zgwWMNWcf08
XjEI4MAncb18NyjFKEzeN696UfXGXmdc0eyZn+axaTLiRIrKwF+mRVY9KZG4UVdf
q+9ElEBSkI9MN6oAq7A3gf5+g3Yg4dSQM2v4PapU5YLNJ9PtAYVqmWyqKkZx6ONK
+y2GdK8dA2ijkysWUVNpPfkGq8Jc2Wm7GpRhcU9Fuwur/yh1M+DoJaiVWGLBqAwt
4E0DQpqLN0R6z35FLAY4IIhUEOuClrOKmVIOGC4oJkKe3TCYfVIP2gPg6nXk7YBR
5Z3qHyuKfVHGaBglcdkZXVOk+n7Nu7uGyWIy+txh0/2SDua8OZCnRDDIn53Wtkba
aEiOmoKcZOh1EwQn57z6I0G7MD0OAZasiguo+c+lZiZR+AMbamxZXe9mmmE/ro6d
ygsAxQP+s0iY5OMVCqmNBKaaPwaLt5wkVKnhuYIRD2e62jXMeSTiOsBsCEnIKqAi
COIWNgnIdk1X70P0A1KSrFZaPPI+lXoEmjY4o7fQbjU/WFFrO947qd29aMBJL8Do
XXxl58coE1Kla40q0fYTKwHi8Wc82x2cL38Hj/Ivx7lTbBdJFimD5gIOiu/IRKPB
upX+xVQ4dZ7SWP/J2fBHsJPf3o5XpNFLaR/RSMqWobnKe8ET2WsdCQBmUlc6gYeq
ZChmvXpLk16pwvzLsvvOPXLw/sPj5Zl7KktZiYJ/2vU5vtjhUR7rHxyDDHkHPfwH
ZfM/VFbhIN/3U+Xbzd5oo7uZvI4azK7YYUOQ+JTRQQkft/3RPkBG0q2Nx/sYh9Zb
OiUOMsDqq0P5M3nERa34pgMJTk/qKoSrrrouMKWSdtHNO0+aIcyUoMgSPMn1eYp6
mDCXsjyDOXw9Uzgo905q8rIfNz1XCSjEjX+zd2NGPzKYHbuTVfRkMb7QhcCGYcEV
xsBfitfn6NGj6XjG3LMi/n8JXFltWkA3ZNY19qTxdj+eowqNhvzMji6JDLi6mUOS
y5bv6mZbXLVzLuLWq/J8WzB8r93enEk4kKBAFM94Y1Tzv45OeuOpAOePYGjIvQ1g
ADz2D6nJzJSCOk2NKdCcohMWChlSqsQhNs3s5fxKnCzchaiqNxQ/Te3+3xjdmRKm
tfEwY8KQnfOT9MHIYtRgEHZD2l7/luh5BqUnNWy1rt6GVjYIyotG+dbsUVFlKsxK
FMroE3L89QDkJ/VtLc3WS+yHZhIakAADS6H3dYfsh1QxHjCg9N9f8goY+zzoRlnK
XyJEECaXzGphwKjfEFKX4GDpeHN8wqhmgp2kxI8xfKo+eHo65qC/XscnwMdE3JcW
MXlvWHvmRxLjFqTYpaavLZ82B4yXTrJFx3Z6IXOR6mMO0Gt5HyM7JNkUKs0Z1ErL
c73qkiH3WtiZUQS1rfiVTPJisB6MlOmeZCUagr+dK4brneWl6ydp745LqF80yqKC
T1pvqQ+uLnEzfUw1PjT6LPrdNeJ4iMyZUzhcSWn8vL5EwYNRtxgpCNxdMc3rz062
0RzSRuLkgKq9QBGAWrxolJYARPlbpoMKrQXq17XuKgJaoQE0cNVzBNaj4uKchv5h
1duwLz7L4tqW4SfFwCM9tdxmLnDbjsjW2u6gsAaTHneUoKytEl7XM3PsZGWrhokd
5ybVKiluoezieqD3oJ7WilIDuEnQWkmk+5pPcMr/kmEx+3fQ2lvN2ruuwVNZZxZm
7xV/E+2i4ie2FzmfYeYvgVAD4Mq4inOVf2XvG2sE89LgzTKdACHp2+IVTc4fHJ6B
HUTrwHvjACr2QHFg8wDlbU7gRUr0fU6C7CeqO6xIPYFOtnLQycClIWUJ6gTwWURT
I9QVYB1n52HMOhgr0pqlccCrcJhFGlOhUVnAstaQCZevY9aijJ8ms/OOlS4l0I8U
rIMaymClqTrcE+3A9UFyf6d34i0tXUGCSxmO+x4M3sik3w+QJy29GAAntkQol7yF
eJqxIeu2Rq8vkiFCrYzUDRSwNItNu4/1JTOufQFTHaSKebIoQv7Ae0MugxOQmGua
DzquqaITUsoNDzfV8ihr4V0FxbdHgZhr1tDzTSA4797A8vt1XdotetI7mo/mqBBv
2GlylM4W2mNfNOk1nZolhvfqzdMMYkv2+0AGhXCEaQm8uuy5aRy3+eVrvn5jjFlL
sIceo3AjX2aRuU1KarEqUsUZtwN0wgbeSLu/SiZNBIBZ0Eok51eZaeypBQ9sSbG4
Xa5pHSgbKwx976CCrOx7iwfNaT3aUypAFCWttboB75TyZPbRiMkNvyOIWeOKEtpT
qqkFNYnl2bkuNU9DcjhvobrR/iuQKI2KS+bJiHcM/Ju4pwu7yWh0CVVanPE6Dh05
0I94KHAg9nkCe4JI0UYGRGNR1p6rDt0AELn3x+twkh7g0s+JIoTbDi6i4PZn7TdC
Ay3JNS7xBscfUKCA3ce6EzxkLeb36Ygwj+vgy1a5EPyk+7kBlA0aaoqVUZ4IMsXF
UpvDRbX4LaGmntUY9Wq3YS9Y9c7QpgTV4An1Ulwh/Np4uilfes7V6lKKXjbRwMmJ
lnlzcinF6DeR55awpG1gS5Feeamu8pNP3k+JX8oLs5FJbtIrUUVf7hxSKDr7/zMa
BP6/D3H+mtRzPvJjat1siXZSG8Ydhpw7Vcm/JgLnatujsOUJZLhVT86z2pVSJV0K
Jbb6bRRMlsh2VVxgiwKLGail+WjT7EEmMVuo8oIIrn8rWrLquD5WIk7A5bMSeaXW
uP3dW/rhwQNXgtFVS/6iqdzl1nsWLgXGSH1wt2x7BFYucM+fJ1/rXt3G+2iBq+tq
68kqcjoa19yai6JJyQridEoKQC3LCJMli86D+fuDh3YgIzbGZYHfGmnWS3JzK4mx
/zxGQqXPfjzU9mWd1MHs00jYH+XOtreZUvLo6/DujvGO7Lte5ca8qZa1fWBCPPsl
27KpjJswU40ICPWpz5qtrFLkSZmfUQbl4dhmTl8C+BG4W3j/F9sctoHnG5InRKtB
fkK0BUHaPaVAdEhDhHSB0K+f/sJYWK1eToM2F2u800zHV6RHXhq/kC/iyCxQ0HHs
0soLaKTr2GVNileBlKWCxmXOOjys8OJjK5RfRbs9iB7maOEJ3waAKB7e+RFH3bG0
24/uAhQAfcE8R2cYKZ7Nwv1bbWIx3EvuiR1NUX/vZfIHHaKttkCLCTfwwiyWY7AQ
5NMJ9sev3ZIHOKd/jYcZk3ZEYJ860OJncOd0QiAaixN2duru+q849MoJB7of7tKx
P6HW4DxMtVPcV18Ow+9qcfP5axGvKLQFWJMQCoMqyqv3/retTNP2lTHVNVHASkrw
bUpgT45DpKAVYNGTDKEiJErOj8FMVms4Q6CzQMBukhkjO/9S+ttnFFSVo32sm5+I
s2yhHe8cv5vPNuHKOE/zXlJNSEj8YqaBY10VMXDCsy+cGh8f2i/acVfWb07kuzJv
aPWqp/FDAsR7woWqUtcGg+6OOptAr4ct9cMyUitzI8DU7MhUKN1Yomgev6Zyk/rK
pAfeam3s9ITsOq2TgVvsP4lugOSyCk0fXUWvuZVLuLn/kUVO7AFrY30FRVcmuKnz
+lSwR6Hjaee0UypqAHikRK9ev5T4jcgV2G1c6ZGKbpqcscX0F7C8ijuE9bayo1gB
yyWQjcjb21by7OVqzgXeCVbgkF1xTKvBY6JQel6C9pBH+2r88ztP2KoO55PlQuRd
bpiqB+WPrJpHuuBTsitkeN8lAm3xVTx0eQdgxAGiDkLoaUcPHmEniaJQb49lu/ip
0EVUENWMJTuNq4QFnV5gHCnogf0ymWugacerwbwTZo3DFsOB3dy55JxIS1CbmIDp
btZa7C/n9lXcj5IfsHu9QV7N47A47NtZxFNjxbBiYlAt1pahCws2CTRxaZe9DUQC
jSFvk0tpb5XCCCs5B6LaOUJXA8ndRkC0WKYs4c+1nk0AnPvTfdkWXN3drvXVT+fi
KALaIHsYzZZiMc/w4GYoJs9dG9V80LiCYqZbABp191P/B9xawFfcdg+n22XdyfQp
In06UPMoMQXJJ65R7COxrVTB6+gSd/x9OF/jO58xSIOa3HpGO7y0wp2W4DpGQCWF
COWls8Af/3/Pjp85jl71A94L/JjsJjjkJaJxtauwe6iUtFkiyNT7vYYg1M2NqCV6
/k+xlbrilK8J0q9gzHmSN+/aDig1SS75orOfn2QiXYNZ7+S634ccBOlLCuIAp2nF
JOzuBuqTspcNGAfClCmWZY4374lFDokeGXAr1TVEVvMh9nJ8AuSWvB35oEuArYn2
fUwRuMh5Lp2PBmUU/H9t0TebYKkmUpsdWq0bUH+IV6KrftTxnybCHbDGxeVCT1oo
NN63kMZ/MVD4TCH+HBdCES/pGsn/cSluhLIUKnlHxPXeicvBBCre28Yg1aJL5H6w
zJe/rXvg6n6O9vxwheQC8RE5SVJtdjn19h/VnSDFInTkg+bUiQRuNC4ULvU47TL8
35XS+rViosCphFROERKYqDuvTrY/yvGNhQye6u7vY/aDh/RJt5p1bR32CIdWQNB5
X7knnAJfEjNgc2FsdPDWOT5AkJpScQjIqHZSTaNO2d0zktAtqt1COpveJQ3WIZOc
yj9guI8x4VcY4DNtFJDGpSpROQmdQohGk8b1vMGLXNZswTTNz6uWVqOnzG6PjITQ
E2OZAVyuVx3BF8Z75bq3REIhlnIpOfE5PYASoIo7dD8GSxMLNd7Hh2YncimviyCK
HLDa/EBSycMM51L3Y2st9KNXx6EHpjHwjul+Lzk1r276LOjHuKl6roFpvHZDatLF
sQLeB9sc1vr9ODnVtz0huw2PA3EAlQXsJDjDM4p2dTCQhKjdA84xSov7D4mANvTO
E04DcE7rww/TLbpDRbexh8yhWlLRGHV6uc9+4gmcBdY63ErI8owqSe/CD/iCwmi8
G6IxlPi12ZKExxoqlTzkVpXerHYToYBPe3ghzOJBvYjU1uykxW0BsihY9OOFUy1Y
m2v1GdHt/v19+Wz0v97C9NDej+kG7rhfhd1oTJsjoHfUNonW9pZTyD5PUy+tmuzE
DCkgYVoVmBke8B0ctCSYizB2Pm0PJXngn6nxsJoMa5xQhLpip7Joa7MllHyCqdBm
vTc/RoMB+GlAzYlFUg0+iIuLr8gA5O4W1IkxNBINvNqNu8HKabouStLHDToD9Jpn
g2AxX4xfWlCnTPhA55pMs8TPQKAAbwYpd/VclXrT9SalyFsHUqhFRCJE5uEN5Ccd
DBnodO8I4yeXPZdD5iDkuVVuN3hw9oBi3clzCTLoIAZdtnG69AHxN8f/xgkUvMC1
qbUJKmXITa34iuXi0lsI3ak+hIhnje+Hp1n9v/OqsNbKeoP4rGzOzglBxEYt0GHH
Ivun/qoLnlswOMsoUgrY+CyUKQP30DuJQw4PMAVBOWzbS6o/dxtSwUmQjltzdPe8
S4Yv2Wnh6WHfHy0o3tUbuYDrfC43l1qLAdmbtZ5O3j0CZrSaCGpGRZSgjzC/ksGE
3+K2M+XDB0NL37+qzwW4uwTEE6mv70pTnoe8AtOuaqPZM0KdUvWz2k/0UcC4nc9m
wuB24jshCtZzXgCYbLY/7bRcVdwtPV7ol0aY/d+DUqAB6PBfvR2pThndLl1PHNWb
mUxuAVyIGyf4wxFEUe87RxcS2YSR0gSOT7mPJdntZTmS9snDJr6VD4xwnF/ukNAZ
LJjQn4q0ilhGnQeOuVlQyixeKPKXy2ZbYkewJsprYM9z11oHizvjM0mWaPy96PZz
9DXZZsTshU6piOdMyNLdJPNbBriK1T0sng644dpYcawF7Z78gwFGdf9wxCkrJv6v
G1boYhNrtXIEIlf5nnK058GZCDCDtDhMqYkXm/VJRuyoayBOSIGMef0652H/lCtX
A2zjcujwGQzoakGw8SBQ1m9dKfUsUeN6oB4YINzzfvNANBfySSa5k1ofVPGGpwWf
anFNQwpXjXVJAEGdss1BlQ0xYECLF65tOt2DrTYwHxZbkpWXSqnWWs7ntzKf5UUB
CIa41Vg2lfhWsa/cYkjAADdlThmTd1BEllBhSYrBQueMYG+K8+Sa48xan3FEKpLc
mrsymBDGKYv+EpmlQzBrDTxTG0DpOkc5UMlN6TXfzCzfZTZzXrgpxyackWsmV10V
M2raC43M/MM5XNfzai3FOIM1dtsuQULUrUCfiK1KfOX2918anyUc6dyWfkln8JGo
6AwioCGLL2HzE/fgUdH3TJ3Zhq95hCtf/YIWoLYt5cqnaREAmhQ1QMUr/UbPqWOO
jyEfjEMCAf4g2fZHsKEVMaews/cc5JPgy/bh2GOGZSkb2RmR23QpCTwVOfcSWsU4
Ayv5/qe+FfqGpyDWEmbbZtLSPhG7N8G3sUkd9GGcq1bzrqQ729jeuNeOV9eiZ6BH
3pnWF3inw1oAYX3htvA8fwwceXBbBHTWgGAfCkAWTiqFvh7r9VWs3nt6no98IQVN
uJOE7vQ62VmApiJAYvq5bbfBMmjdeEWddprwknN5UwKV+pEt/orek/tK7Ogv4fqH
K6/cpJjZP2SIlgXlcS05OlZyasMsyYGYFIrs/3ey5u1owGBPBWYiNfYrM44BPvco
Ukf06q1iMtD1YtBiZ9hIa96ktTsFqeRVg5THiwtn/qZ2A7eac23fmdLhH71Xvutl
EcmN7TnZGoQQiteo8PSZHjDyTyhQ18dimvjFpHk1a29Wf9seXNQlO25zi/rF9L6q
wABaQAmoPagX/7yoehZloVFFvAZN1NpyjUHJE9xRHJolGfollXV4uk/UWQZ4Poi1
u8kvFugyTaPT4kMc1ApgQJNqoLBUFQIWXwZWXgPT9o1FXX5KE6f4VDjRlhxz+zt6
E9QbqDUQ8wzgqEGJ0VALeW/37WbB1SsYn9nBX3vC6EweStMWjcUyZx78shK9tJUw
W2FYfr9rAMwqrXNp/WItmoj1Q9oPLJ9XeFo+NTj2ioaEcrfSaY/ADy0O7OvCBEod
5/ovkUPSoWo0XzMLhnPKveGywq8n24x3cCTsopwx2hb25ikWbbN2+3LMX6RkrGUC
bFPBgz2Prc/rI3UcaD7jVW5nVcebvsq1KzqnTL3Viq/tvLJPyhw8wqpE3yAtuTuy
ekfYBkKPZDEKxxd6eg+lVnujQ8YpxKBDQRgx01FQ5iL/UvPtOVKZfTsoi5DdbQNL
wXK3DAOoOKuF0umZJCbI6RExI1pUBI6i39UdDgpq1BlUNu6R4nffLAZ/EK7DWV2r
tbhDJvfQI+yVTF4xMFAnpQx6BRMrCrwGVkeBanNM9Xzc67zqUxY2AvIyUcAgD8dc
CYwEDXmRYZiyhEX4Ytv9g4/ERq2pE4bkX508Eopnx8K3Ycyly8MpjsBGHCNWW3LZ
30e/WLjFmU3fm7eGWQC4gNKa8UjUMyermVzeyT4q33zZrG0ydfAOw3jrtp+cidIU
Q+WxxXof1HYc3Vu1IpJ+26oPC1+tQUKBw4s+spuni0yJv8a7+84yY7zqB1oMHgrC
zT9wTJNfm8WUlsKF6aUkRUifiy1RbQQAI5kGi5bNUq1xFvx/02HU4765omHLYlyR
Kqg30k0Vc+GLfb/f0LHI1kBF30x0IZNGyWLTqVl01eK929Dd1jaoMSavls+uoorE
KzuPki3NDZfNHBQYNmbB+KrZbYVyvHFihkze2bPsNo13m9nKWsXzvIQTMCdPwRNV
NAd0qwNDMZVxCscQuzA+oV6TjYWygK+xxz+dM6maqjFeOJPCZEXBDiDB5i+jsIMs
dKD5/m8zUdNwD6+15lCh1zuoH/MpC9emvS4KwfH25CtREBsM10mlKs8nPWHYHsZm
4bhE/LI2k3yaQz1d6nMrUM0l1FmWuignz/2AAOl0mAosxUoECzhCRd4Ai14ItQWB
zmHI+9fxzRnBdOuI7KmjeL0Zu3BBJ7YXxPETI6QoI5yuYkRIG4buWgd/WZz9Col0
XCNQ7zwk1+0GJo1kDjFtTP8gvRiDRBGZtzm8r+26EdmiqxIE7QSOOdozt6M2MEFL
LmAHPExN7g82Zw90xegnUl4Y7fXWLx63d8QIhp5n+p5B7uCYe9n5FOzBHmSSwOjd
xonsaTGlZlN9JYTJ9s2Vg67Q995irQrqk9OGFttD+A18ymU5c0EZsWHXVay12k7L
lFQqB9NR8XIwPRXo/MGs4aeldDpZhxgQUOR8a2Ng6ppboQiGJXXQ3KjNo95KSR7x
r41GPmmt9hde1ojtKWNn0xUDveAJFrvpDtPiov9KP2rW+UM6CyDZJk9Vbr0MiMCw
ThrFJukBqZyqIPuG9TRDjEM6eu2BG6GvoCoFOdRvIPzyWh45bIX3zu2v7ncbZXnx
rqBVp+dIMwoHBg+VYjMZ/DFKr04ez78OwtsnvDtxMtSCOKdXCDnDZ6PJeT1xlquD
/ZEbvV+jGXSYWCgOxfoV1C6L00esfYAIGpWvltF+k2HyE1BHsKnG0IaQ58puAxmU
/3LkS5OQdNqNbIJlXiXUcJvogIpcubIU6j4RGjeve5RInOaxV0SUiLf91CzLsoyW
TFR0Ggdr/75+b114jk5aifxKpqLK78NCMpXRNls+dt6KAsug2EjtTQizU0LyHTsS
HvtV1pc5s0f1o+IymaGOjkGCPJ8vv9AOZcid7E8XiNSSVMA7v3Q7sw65KRx1rpl8
A5iF8HMAMCoYegQWpIS3YPoaRNgFT4lQMbBpL/NhR+zguxHQl0sIgvizdVMWs5ho
N3fDWj3Z4iKOG1dCFmXpwKREIEXNXSZL10H3d/S/QJvP8ecIIBetWZEFca7YECOL
S4uxwTWZChLA+9mdFnTT6sTQOjIeWWZ7YKSboEwENuGLw+Wt8qTOnlZUcpof3am0
rkFA2Hg+EvqBvko0BcfSqXZFKXYfeG0s2ioIDSvmfwgmuMq7S11unV8BsZsIKYWy
/jNhGMWwHou/9X02VVSrx405vdl1LJtAMe6sM+kI65mCC3WpkErwGMjV229mJSid
f6HMb4uur7brTIpGAA7MvQv5wUpTBq21NmM5a+dp53HeiKnin+29o/jeYbQtUpn+
5kO0fj/v5dj7VpuvUu6JydZfWU7YfzzplAqznIJtngitjBNHGKlA8Z409BRqWcKw
CEOabYdiifWKYn/I8lipySa4PXhc4QVRaWsclXla6/Q4zyk5Omvy+yvwvIuSRyGE
2KCA/b3kNF05y8G5l2f05o6+q+yeUWtj8iFn93ID3TN3m71izLBe7rcKGcCboSg0
C1E3cWkaGutdrXBznonSlYaYjbO8ejHQBoCIHETgME+kniJ22ol9a1qu2lqxBmgK
yBNNqVrTbYuJlPNvOzZIaxTvcKFTECxSsIBxz5j22rBDOWvajM3AmvKBRqC0qDdq
wxHzhM+ICWreJikflAdO4GifroX3vDzX5cKobdeihpOx65ugek6NmdoYqKkI4qz3
Jt8BRrLdbNsIBBYO6JR/dHZV/35KOY9eFic8Z4Yw7NZRMMHP4JWKb5IKbum0qXmd
F3kW/Fsm4WJN1cV3Lo7PvKIwofdk472o84mbl9ujvH4cLjr44vqIwh/sfTx/tiw7
5tikOgeU3fQLWmgdvrsEMfhMN9Jd2p4uriedd8wqRE2eUg04dn4m3/zbCiAIF82l
Ati3nSh3nxSi8R4zw9qHDGEhnd7Nj/skG/Bje46DukiYrGpexbnnr/I4rnjkru+1
jGl+/Qe8tUAozLqaku3aVvqUUwG5whtc/XLPRJRCezyDV5g7CuBBkNAbsa5zVpxm
2OMA32X591eLtX63JNyFCMCQZNOqhoN7RYF7mrN9Xj5u8UChsUjmwGtGmTfPrlgy
mCDDSAqXs7pc9RHPFdYSgbEyh26eB5yAdEf9V1ATail2FcQOeSR3uuO8JVYzHOk+
rTINtEdUmpQ3xhzAT9YsMMNs6+NBkjYUEET4Atet/+ZFz5MElujMBD8c+RtHJHPP
m/W/Ulz5vaFw79yX16epOI3D8zP4PnnsOdMlfufesTiOfQZ07D1zPfyzaNAqyojj
LK5RrKX90+S7whOFrHuNEosIN0IqzrCajckTFI03Z3BTeJfwWe2wVmx/3366/kF4
wDQaLwpzpxMdH4/jjuU6HT88wfqibMBApFN8/3eNlhmCT08fazopWocllcqm6JSF
2wlH8Gu5dzX5ZYK3dcHtzeLWw6g1wup92xSADGPW/WuQG9pyrkPXhOsJR4qsxZjv
6GU3fQs6xJ9Okd/KX27n/nNwT8NPvXAlhewE2MohqO6cVIDzavmydKeG+8++xupp
bg8NuN2ozLrZ7OWC6fK1dgBMYcD4aULxjcNy96NqFokQAdGm3IlC1Uir2FA/O25R
p43zSmRDBAlFFisVwTu12b5WQJheyx383UmxNTjZjDxK6mtImvqN1blpyMEESnxm
486YCE0jIAvJWa8A4Im7WtJwKvRghvDRDlyMhOWfDEZdDDJwZNatcsxBuTFqiYFQ
MwA/uT65T0Qq10f8xQ7wojgN7q1OjbTNTmqoBrKUnq7Gytvxl8lWzYxSB7rkev4G
ODRfW4SSp5BU7LmT98L6ZK2FZErZXlXrYuyT7nNbVpYBI/wh5cyDkIO4APfMWS33
690z9xv/ak+8SDzI4xCUZgQhwE8GLAWk/biu9Yul8qoqw3GBlbP4637u5c7yVc0W
Js+PhZf2yKIgkx8zqIWXY7Vn953YH8q4Dg5kZTS+PLnkfKQTWT9dtEZOKrHFhKbJ
LnET09XZ9PBzMecLwbSpz5R+MRD5fY3mscQTTv3RQWp2w4lYXXCndAPozMvEHyqo
iDDAwFptzk8Yn1uDHJWN4c0AY5K5ww3nA7ngLpVFvY1eRoQW8apd+tkC1AbSTWAj
nWe1LBVEaWxg/9uXwWVGm+nFgzmeLSRqG58C0AA0Y8v1Tho2R2xJgrCDD+WPivmq
NTG9qVBzkPrwqhFo4czpaT2bZcNxIXnRe/Wg3j7PRfbPpXlatxtTRO+IMO3PZwzS
RQnpANZggnNkKLf9F0vGBzg2VQo0h188tFy4fEzKqT4cquWGCs7uNktMvlCk0XGH
YOFIynZlfE1Ru/8WUz4yt95NOu95fVIVHSCTrWV4ZRvxH5i6GrJ1LT5WznLXQFWY
OfNMNMTxFxX0501Goviq4YiUHudVRe5sgpXsyuerDdl4v6RawAStP/YAx3o/STYr
TB4Oem0ZCleGsodbuGzu5T6+O3DTBlnJxXGy3ZxybQfYlGn95DULac4QizvCtFAD
vLg9HYEF8CWAU511TOWiBt2vhNlHrvsZFoLFnIGWxabsQcEme3T3/tS+BRmhJNAp
/eyFKEgC6ZEvO40SApeOUf4baTXVJHxOphYCPLgpISRxFOiaJhwklR/BeVIgTSZE
+5pOprKLXvmafmiq5UYEyJqQZbeOiHkDs6a2jW53lCmEiQLzcGrOEbbOAgP9HQ6G
0d+BSTKYJCqMk4vCS326NPpvSTdNjjf3joa5TW3ARfnJB0ZtZkDR8ywl5uCEsoMC
G+UARppGYqHchu/I8uDHUli38T2oox43KXAtTpNDdspzAh7QWGaE+FHb56YLOwzs
70WVurD+4n02jLXRgqlap80lJJBOR2lVzjkZSAHjqqmQkuF5vIss3uMUBus/PxxC
xlNAqvHONwdc7VlfmvzEWPVNCp4TTPJFyYjACfU9QveaiZU2773ij9RdnJvva7jw
V6V5dZ83Nystr6JKKEg2YbE+TojJokCH6m9GigEVE0a4bNcx7VoNqodkuOUzjr2I
qWdrdlIMpqcGaG4eQLKxJ/jFLRue1RAQrcljqjHZLItExJpFsiFaLOafP9IgjGxl
Hrad44ucm3OC5r+w2+2Kdix3dlV+CNI/LL4i5zXb7JNS/xdezGUB++xb3uJooB0c
UQow1yEfiEVd3TCZdw6ZT7s9Q8WxHSkznY0d/ODlLg82yObXMd8eBLulCdzImJcb
2vjW0tzwu6uk8vqk0K7GAOGGrlr/4RzZEqGaCxeTorMQqdKb2g8Y+WW5S1mW8Cg8
zCeUJMGC71yob8V9b/Rm2n2FY5TsVMOgjrH9pRULRJTm6PissGVoD8pgk+AajQ6Z
pzUUeRCwkFwbrdX0cBvLrpgMbLNUs3C1SkV9myNOXlNEhlG4/3kQ/cjc6Na0odHr
c2VFKoKY21cPKTYVRkIYY/7MoP69XucUaMTX2WnzGq4qIp2g4RDoYopECE7BMlhA
EtVhyGCI/UueBq3bg+qwkqRg0ANyi2Mlo1bP/Egcv/tHlkrboFw3dJYtzX70P3Dq
pp3Ub3qwtv3DW77Bx1MO7PphGq8Gcq1v33u9/WK40SN9siOvNzPziOZf++HnGvZU
+xCSDQyp1zvnmuYVwFX6AzXVaqpq/7A0ndoWPwiBOcrF04pkL36Go1MBFqC7TsjI
KPtWs4HewD1JEhUn4QZ3FZBNVRAbeORf5KP6eTWQfMyhCqULNkl2fwcpCAehFrpc
m8WfA+EYsHkKlo5j4CPKUxgLkLuGLlYWq8aPCb+fxMUNyK5WRlMupfsHaVZD13LU
VNGHp4cWWzzHjQUcjA6FRd+3s7xQOF+NccBuHaqyzUIU31ACirmQzkrAwvycYcPd
W0nL/mt9dPaSki3gWDT0i5EiE8bVfNnQUBINSVuwMVt2ZpPhJ0CJ2tExxUWiSS1f
eFZL37yayhRV4/cLou6qDxa95qMJwqeWeLrW3kDHTO1chRtUCNjTDUJ6Q09lG3VK
0RkVnMMYF+UdgE070we/YwA6kqGv7QgIYJD7ln/R6WHJqswoYp9/rALuq+11SRU6
MikNpcnNkSMIL1NXrGIeT89cAs9qJ5e4qzLw2r4JdzWVdu86VDjR8v2dtywzf1rE
m722gJygcvY+htejB6/YT72DlYgT1OyaBt3UMZL/uoYn5b+XXHBpE+si096xvHFv
iC1jvPMtST7t0znCBNuxOCyPeCT4E25EF3jrNPEu/gKIhFV3rXANZFL/GeiHvKAE
01FBr83xbll805FEdPzPnNe+wMEp1bunMwZzfkfudQd8lu00ejX85JnTQe2cwGxH
ReCrGw83/QeEyHuQzM6pDIw96jAHVTSQ0KfOVCF4mr55n4yde9cSHrYt1LP1l3d2
1w7R35WGElVRQjC550Lw2LYSxT9abnHE5ELcna0kv2ci51a/4MMcaNzgke9akIko
OTCncLCrKdyWTktoQ9nycc0ACANUGPyjqD0vc/0etdWKqqhmNUcK+YJf3bjYB3x9
Oa+YAcvg6YK+UF2uVEL996sSJUupKNT6ucO98L2f6LJG01ckHoKMqjkyu/u6Dyxb
hW43xmwVjeAYaNFW6w+2yIcOqT4NttkY2A6PoT+GUmNNo6Ea97dtjCnf46m+cf+D
FUQyVYB5Vd2pBMimAcZe6yYO6T3orkvxmtKpiV8hlQ6ii2/broJPwst7TtttpXv/
MHhLjoNV7Jpgr6xAxARCd4ku9yPEaAb+raQMlUaZTiPBKf/Bdl59SbxHkZGnqeed
1tCLytO+e/zyLJx6HpeOu4qs058yHoI4jGjYPFLuSNC+6iceR92ohoNWl/xrVgJ2
syoHoEMiNk+fMHoNlJYmvGI7V+j9kQyiG0Wwa2QKKvKdB3R2UlWRKJ5pNF9V/dSQ
QSnkMwm7P2YxFrJawIzTBtidfqWINND789Ke1mj8LSC59yq7/cbQgp8Ear8JIeiX
uGuj238uPAW8gk0nIOwoGwOf8ujl6YGXQeVlc3GOdcfNWfmORj+uR1esd+CqGOjc
7tNw4codlQOFzyC88mlkmdEWvb7IjRVOUNCWkZvRu3dTp5nC6oYU0aXDnTvJwtSj
EMzL9yElJ8v3ie7khOIjlPaq+IdTOyZDSggrvm9GhykIE1/0YZk0fHBsXm6y8EyA
E9H/vk3c+3CGq1DbYaZzFE8VyEeSk98+6JbU/W7N2cadlW2zLqoF0qK9Mih8T/Qt
rCQdsePBwB/f+/F1tctXOQnKq5h18uPgyMOW0MIBGQRjqp38CJjRyiNzXtZ/6XoZ
sh4tBmM4gT8p3yGXX5eeeoh8ZkmmzVWtE69MKYAdCbuPgErCI/+RNGPBNJsb05sB
0MnQqMlJ80c+yNF+sxYE/iw593cc1Uyl+pGC9YplbZTVMpEozksUfhQkjeaADnSJ
5awv+BfuhwzRloFMkoYLvwDllgUyWQq92/+fg91twwyoEnc1LZ/b+nmneCCHgW4L
0h7WHBOG2AtlweTy/+oE3fZUq8BR4GOrUtM9pAc5DaU4D6j4bP5APsVQR440P5k1
mPT0AnmTx3GkkW8PPI6dNVxHSEFPwimOw+ymngYzQSeGSBs5VlwMF29zgo94eQG5
F4RZoeoKGCMUmI+Jr2tS9Mmu7wJyjtc3U2rwQi7sbTfv3/eFzdNlNwgdIoSqZBsZ
dYkqnzkHrmAi+KD0phELlCfD45jNbJRjbGPltf24P5zQbtHn2RDLb06QCSxm6zNc
0vJkvPuKuBOtzm3l3YccaELiEYGMSi+3RvLhrmDBzWuESD2x4VDVQbI6XNCnFj96
7L/mgd1r7OqKlFhSpDzOKLbszucEAS4BL9wD5AjU0CvTG7wX/z0O0LyOcJDrqx3j
687o43fkyVKt5CzNABb/bmWMges8rAFoCwydP3z5hbxP4W8duzUPY0J9y75vGXaP
1iMM+t147JXv1AFsjHVp9O4g1/p0t+fC0cYHEkZluM4/FZ6BZHamTQpfTwLDC1ea
MkAnOfWfSTcU7wQACRJkQa+3Gfug2qKb926ZfohW3MxE6FX9QrTAeGX/2MlIqzlr
OoCjRk64WpkCfVjRrilIvZJHt5SbXaFbsUwEYPuQwU+GhvQqOYceOVO9JPLR6OT5
2JIqnbK7QVGwOy526cNjykhN2nb+ELQwG2AgmcpiH02BYCjS88s4jDsj/+24z4mT
gN0hvSnHaypWttTWYEuOmtW50jKh9NGAnct8DiH/1g5kbl+4FZrsQwyrZwBe1pcP
f/qGqcAtJWCI2yV/PSjIx9YTZIJ+pjPvpljS4InJtwoo1Dej6Eb3mOUCBLu/zKjv
B1vZy5MHx2ANHwiPS7dmjwp6hJruxSmkukUL/V9/nDQf0Ii5Ob7XpHUQRBjnL7wL
B69nSDQiv0zfduW3kuE6XQk6vtDzeOC/MAlY/JAwswHuoypg/S6Mx7t5CyFCtmQw
Mbuxj1bKuJJ0S9mnS6Zr12KtJTpXEegETUAIM6FKaifiTxtp+K3hrYRQwXdMdSGc
DVEkB/xGkoKVkt7lVI0FZebEmkOOhoNVVq3OVTERktBchAmZCXKCiN7UO/LEJJzV
/6vEN3WMFWY0aoFyX1WBMM+DkSjLagFD0LyfTLkkU4t0/OcVmH/aK7XkVKjZ2ogh
0jjKqGBCjbQTkK1T9ymFwZsNnV/RhKjKop+0UKTUmPsRjlKfcTBCfz4rXVFfGUwd
1D39mkGNxDY7vUX5ZHtueWKBZ7uobqbkrE2ei7Yy5qfhXpV1MTnW4OAdk5PObtog
RvC/FKtJoqZIB2boXL0VrntXDJSDg/tp8I8B1d6svyugqc+k5r2Kz2LUtlOSB8Bj
wUpwpjHFvB8B8YtbHZDk43nWBX87YnU79HA0yLLchkiGzs7nian+NySKIsJUV4Gs
zGJYUtuJ1AaYxKb85TEdZH1rje2JXxUWMsVhx6Go2xM7Q9gosN6lgErf7DdY8GKF
cuF4O91ZX7YbzSJ9j229mcUBVtpjZ6bxI4vbcNlv7SHeB53bcOTaUUKVJKrszumk
XN5qCqAnhHt9SG0nruwMoh/s/tKvrbOCM2vSwhHi9DOm0xT8zmZcDCGtesP/oPhr
xWf7Dm7oinkc3vZF+qjHvwl64VxnTG+otpwWvSyj/qttbg9JB9HBW/1DqcncCyna
UYmpTn0T08Slh/ZBGzHmsYhTkMKEG6ZWJUgD1rdlgF0JlQpPwN1wqYRdil5uoyrf
AcJc2WPMCk7j0esle7Tz06miotMzxHfWVD3YEx+PAM5mCmPgv2/OMb5NVZTmMhog
uot9gHQ7/dotVnyqWzlBrbVKFPQ4gXBFUrWlhZ4ScZY4vrvXe89zEcJsL5zI4UQr
sn+0Nxld2oZTfsA4AhsxQRnNhJErNEH/gYYkjvzq2mgFUMKjvEX35frkYYAi3GQS
ndyghS5b0dOEmjIBNeFJVyOhRAdSPWOGkmOsA+yv3S0=
`protect END_PROTECTED
