`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V5NsO32++Jc1rhXyInQtay6lHOSOxNSTLDj7dblyxXiT6clHsA4deMJqAZlxP+n3
Gn1OeJx/CLzUiPgt9AMq/V7rus+0adUU+ur1RgNf1Xyesz7WOXLbBdqyyHJb47aN
hcA+TBP52DxO5ykUGt4OzQR7Qsqh0zCVjYOMj18RwcBg6AemDNI53t9NdLRzELY1
DLLywaRlgBX1cFnvl3QgZmrmVOqu0FV968cj+tRMhMtEhqMrn04CXHBu3meFKDlz
kvsAHADGBlR8cPzX6Wi2zxiCLuaV8+/HkrQA0T2d6e5VO5hVeNDF5HUda5tY5lvw
pDHkmdxn1/FSTiRWwNzoictug46sduBHXSifAcKL+rnv8Jj4hD3Pm7t4R79Y4r9p
PaPQNrWz0w1MnhfHm+X+5dVb3TUHBUh9XI4JkvcyrCXnQv5Rxg38pxu/BNnHGXLJ
VFYtThuFBQQ/Qyh9Qr27Orl5nVJsp4pvXhNk6ofBLjeIKkRM9c9li85taCWKJ7vc
LjLvwJAkQbpQ5Yp3AzuzlmPqp4M6Ba5L7vA7o1ALHx0Wtr11EsmT7QaDElGnYZr4
x90RvG8Xe4mQvG+t6iRoLHk/IBqAbkanqIoC7lGSakOYhn5sRKNFXfT51cLx5gr6
RmE60Aanq1S7wVot80QEzKhACoT/d1iIRBheXUuT1uvQzbti1uZ0we6JlU6YdUyt
Dvuf7XgfqcaEvnW/xHOrlLpGRbm52xzyek10VnUuMIht0AvQtBdD4RHiY65D7mqW
Pz3aasj0s9R7BsJ8XUfIULil+94wiloPnTdQ6p3t2FTDrBvmr1tTXpks1PaWY517
GDacQmiVb78459ZGAacFk5/yXvyoEZCKht8tT1i9v3y7EfCw2CuszL1eAMNWG/rj
SQVpEHA6RYbHtZeu/Au16c0FOs7Bt2x0aa2P29KHU9oRHVOK4/cjz+XtJFC2a1YB
+8Ttw5bVf8ajYrH2Zdvhn2XUh7EA0Ms8sT1zu4qfjAIrITEaEUec3UCjEpKg519a
y2IZd3iHF9yk6CSr8Ne1oz7e5pVAo4dQmn9DWqvNN7opkFcYP+6v+Ph2NFILiTql
`protect END_PROTECTED
