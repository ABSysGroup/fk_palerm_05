`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V1Oy9OhYc1ZkApvSzgg1gQIK3bOADyY/7f5u/4gU+sB35IAzvZB9NVkKNSv+kC44
hGQmnVQzvQmchcq1EaniMwAe954CZlFHYE445jjrwzet1DYGp9pM2OjHooWin7ug
zv+qbVjXTSK/lWOD4wHPVgVBYV6TC9TmLSGFr1ZPWk12zusFgiN13CbXO46TmGeF
erlYJ0GeezNu5th/mGXRRl35HaL8Y3y27CSjC6L2qdFdq0SRJ4DsY9sAv+rjVwLP
WZSS+lrIDhZsIq0PNQOizmMh7DABBPazPrUWGTxiSSLKIGPxsg5UDQe0kow8i0CF
+uO+awjTC/DG6IJVfqEevQDHgOO9O00gszSswpXndar52XaUTEwdhMExcoINUTxX
xZHAuSe/la5vemUW1xhMoZLUG+F4seLvb23XMzeRcZ3iou4tCihAcahrKABMqCvb
z5JiiX+2n3eZ2oyFtQzIneKnofbtXZpr1nria4eY62JGugRvgvPKgdgxtMCLxbhJ
/R+YYyew/WkfxiJZSyE7Qdm+4w1Slvw9Jwiuu6tDxiN2q9YHWVB2B1LyzWUQrhIH
OlEBH0T1l4rsEh9Vhmj95YVTQr88f5n4ZJCCCeKeJph3vja/ijOFtdoU1ZFbw5fK
xLr2G9DZJdHWAY/yfLOMRw==
`protect END_PROTECTED
