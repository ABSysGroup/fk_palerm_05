`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dMuYkWwGVHLDH6EQ/wwDYBseInT2iMXcpArDOjRdQSO+keWcVPA62Z3Ow0jrRsY3
F5Z9qSYZxrGEiJ8BVXsdJUc+QWvKoqTzvDvwXV/m6VbtZbfvHmHs9KSjFEfE6Gnq
iXk5CbhjWnrxrvLF9u5wE07zWrKjMiK+dJ26jpn5MNWCu+TemAZXj6kmHBIHIXWT
Q7borbvbzkyPNcg60zHs1jWYwILn06SE11pZrHt6XmX2R6g00RDQlW8KkMNXc0Tu
zjKB/odcpHTnxCjdqU7czZifsUW4rXs9xuxXCMS/DhEDAG94L/rh8tP9l8Jfv77C
RDJp1nRh4jPVUmKzmvf92xGXVUnuC/BSyheqEsaNMpad7OGGJnK1JWwt8M4ytCQS
+Q++eyg0P2fidEMqnpjno/unvol+vyNPv3d/ydBGtcqvaA+07IJtiG17Cyp4sWiS
eAAIAwgenzY5tFgEHlYEVpIRGhXbWPv4R1rzG02LLU+lf87onJE8fAaZchTTUskH
WLW0VhJmauXA/bbgMy7HwOdO93wXoQd+cvegZw9Q4V2gdvuRm/UGqQmic/uNQ81f
fOYMuk9U9i6Nt73F0VoNl9KJUubFN0CB76OVzwyyd+P9AMcTBc8WX0cNGUGnWKWC
0XSJLCyM3KOBvSik21kNrrvzJZ89htsP4Y9kIDTlHgiV1RTzEXHNL6+RYIhnwQMa
rwk3utscxUehZ+LJtc0xRAG4K4uQOr4dF3HulyEWfmC0iKioS+s3jTDorhlOnzv5
0kx0NvySD/b3dQlC6uqabA==
`protect END_PROTECTED
