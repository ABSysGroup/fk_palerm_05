`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DxwzeLCTNuj+FK7VlY4/Kw5GHssc+7AOFnPxVqi5h3OSeIMYhcv4r3mi9MYER1iq
dN4CVjO7ZVe8NrxTbV1Z5X/Yp7BS02/IGReq557L8nXoKB+VkNzRz5JmJo/Smom2
N/ftpv3qL+LkvBB7h0mSed9LSND7FqdjfWxvuz+WA9LCesKVI78BDQQSSSU0JM76
vQ3sz2kICtkjOS7ZpBbY9jkOTcY1TQytp8cc1rSF9R9FnpfV75P69ZlFIIi5LkWs
uZSLrNbqqTGrHrjtmRD9kZlRV3czxD94O7km6Ka8uJbVZ8kxTo9H40gzfmqyvEdB
bIcRFnop6OU7SGIqN28MJfiieAnQLUy3rMhXlprKWi4c3FMao8C6JyBvlzrGDZiy
wC4uGBCTLVnfd+Om4UDD78rsqwFZbv8SS98vC3PvDbOu0KKfSxO5Il3qO/WEP8LG
`protect END_PROTECTED
