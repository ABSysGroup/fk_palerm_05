`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aMaLSTFoLkMxDbXjvtiji0qgxvpBFxSxDWM4d4Eo5863S06HplDwViZDJEAiMH63
OSOEsXVvuYqibWssJw41+d2DsEfuRfuU8jaLQ82E8nSkcF8zb+wlZDBEVyx7Bj2a
NGtrB1z34FgJByMybWq6pglVl8al+EaZNlh2waLiJROFw7k6xuVptlNJ7JETXVkg
t2oHrq05tn61REhZ5gOs9tu3iJRx84lNdvY9/AoZj8Rcc4KT2m+oAnMMfhmNzgwg
h1fRq810PvKTEBUAWR02cmL0M34S4CCDF1m9NwSY/kWGEJrKil3YVbPxdaDoFacG
qgQTbOBQG/gpZ/8Y4mFP1KIicOOV49kvtyZE9Exp/3ne8bvm5kvFXGpEwuVzVYXv
tPFcNoQlXAHD1fz5ErNmqVACxVosUqS3p0rUoN99M1xdU46UIO2kge5woWUiKLlp
UNlw/oKiSxI8EqjnBKpg47hUH/gVx+eJrxIuauJaghnQzY2Ls2W5oDSv7ZkOqS8e
2C9zF8IwoP1oyEApdpCO1VoA/3I+KaYc56QluFmMvp9Evnr1CAlLR/rWQ7Vm5ujy
YDzSxW+0PmJhdtmWkQgmckS4Ba6rZtKZPOysTIqdOtWG0OWSYI0s0t16+FBYHVvn
ilIMtURUmS4WdCF+yCFUcp/S994/LcxOc5da+JnK93+T3M3zoIodskAvFLr3tV7e
2FjEhQYv77mka6sm+bIUvEfHWFm9AbXLIrLOE4ayuz6OTKRp2tRikyRrfEBfz18n
r2oFWfM/dp7UxM+wgDIe29TMgKLMyk+IROh4uMguvDJniMRk/2ngtShEYNB6AKym
x4Vu6PO1iDaPaiZa0nTQdv3Aqv7PVHg6FYRaGNVSOcOxyVlg94XO0FsC5uGVVfrs
UMzT5rhIzqdpQbNuc1dBegAiH7Cm7ZWT0SX5vMLYqiliwDo7goNPJxwxCzAGV+2I
nwozghjf4uvyR//nFcPYD79Q1lYjJ0tPVlX3kl4hifkOWes7nZi0WDscnZb3vSpZ
+2c3eJRA4UVw0nopWDnyWO2+d7qpmPi2fXTLaEHn9lfpcu7Yxr9Jx3yK3lCQlQq6
W3mkfhFmv4JQm9Vw35wasuIt3SLq2xpzb/nsz6vT5Os3nILPTpG9w2/53dfpBriI
h+nfAEIycoF8oG8MvJZDNnCJUVPbjFUT3OXFfZZwYjN7HmfDCttUI73xM3mOkbXj
KiNqj7VeOQRyf+m+u59357WXHEsNADtP3xzJbT+c+okiIQZu2NB/hYrAcgGsLOo0
JzyxnXRYyAA5TbxEOaijcIfPpIsyXPLm5JVeoIKL7Mw/kK00QFFgzpMGHtkyrC4b
nPfxEQT9Vn9Zlg7luN4AIwfjKDNc2wZ41yl5OgLVk6kC4BpPOf99VHK2tt1NssJz
bW09HYQd2VzDPAfYVVf/ZIFY7q16edDHseYVWdLjoaWcbxN6/Aa+YGas8VQeQ76z
tlSxNOk/Am8g7KoMHjJobxDDcN3A+pEtZxk/00nJcP6goiQXMK6d+/vISl+NFdbV
URcNN47QqJgTmQVxRfyPczHamWWE6dNxzs5WBFDWRVuyNjn7JxRq9RbdM7ADAA2D
CteFkCeBZR+218uMc5fimSE/F/5oMwKoCYKPkFdRqKptEP/BLssWbiDA7qMOJs12
swNP5xflxJEqnNCN9PZkQPNMIHX+86JbXIgv1N1xR/b0leE9lHeRZlj6miWaBEJZ
Ky4K/xLCHHIKHnhRGl+KxAk5DuX30TKG2EbHzo5uJxrDQ3wzKoVjvFSjRf6I8D7W
TwkoBYwK3sC/JxX4K8TT70Kkv6Q7/sjGZ2km4Wxc1ZOb7C2d3H+be6i4b1baPb42
qFsB3TDlFqD4tx8DngpIh1JX4fRmJHTwe7AuuLujmv2E7FbWAvZH1hbI+6y46cd/
kqIXs0otf24DU0FEAst70Diz89BuvWvpcYd1tu2fZo+K+PU2y01WPniX4eGUWv8I
mNI2hTqUkcAk78q07sm3pljj1b0apYiGPkJzSg+hJXQHS8jFOOB1O+ZNgY1o0TxN
+e5xMXMHBu9BgAb16rPZDRN7V6PkLmU/aXHC1w8gl3gZ+TMSM8lRp7189rMAnjXK
fT4vF0Vunj5n6J3AdOGN9JapcZAy0Fg75nyZvrBLyMReMLo3pqaJ8rXmtlkJTA2F
NzTLIDitMZI5uvdOGq6O4I5Uy4f/VETSnjKawEJsP74Ew/J79bLmk3Ln/ztBlgRr
UvGrJ1HCq5jcp7ImlNCH9db+qXBTDjkb71j2EeSIYcvsepqQ0LQW1zZpmQNqDcfH
ICJQnX54obaqzWCZOuauFQedoKPFLSSW5Mol6lpsq50FXMtuLBzE814J9//IKMnG
VYSHWr5Svp0m+pIlkT4wOyFKtOwK1+3dHbe+i7yVMHpKQejwoWh0B+6GFJO9boqz
`protect END_PROTECTED
