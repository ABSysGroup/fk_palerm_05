`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eij877QJJG57+try9wBhkUHMnDKh0tiOdCXGhKrnHlCEnXAxrLj5X+0rv58OKvw4
hffKA5qciTSWhBLO1+pqFDLFTL0AkH6e5Bk2p8YPUlD5eysedUt4Hz/VPVJjJwF8
o138/olFcSAxWhKhxTBbA3wx0Ez0O40Ip7tEtuPixpPkv92NGKXAHJFKhFpevJr6
orpcbbf4CsXIE31mPsYJrmXCyfn28u4Emp+YXTI0UWRpL9X+Jm4d4QBnXtSwz5R4
V+KFMWQI2vzQGASvPC8y1cqp4K/RkuY4J4aobzFst5+jyZeICx9z+HIVGkd/trM0
b5MVFnKFt7wmZNdR7eOr5oKFFADoO2wCSclO2Hn7JjWCgwxxn9K9zg3hDf0Hdpmz
XTnwQMxV6K3oy5GXV5nqoJIxaCmSdtqcxCrRGK3C93SCuEVrTolwZYNSx4lbc01W
oB6kqMq1SociX9B7CwCyyE6CJ1u3sO2a3+sQ5vt0+jCHe4z4YD3HnK01U6g/Jup0
fElUTEXA0J7gplo/1x5aGVaWLmBeuCUjtTthPiPS+MAvL5w5kT7tQ+jYKQCvBSXu
rJM8iXcgAcxgLeFhF+1PgtUnjVMyLgoHlKxmNbSvhqa3VjOAJOH6Mg091wh8teFK
Uqilnl+nYYzfmRnppky7yT5uOXZp5b456Pxh9N3ipOGDud0AI5e2nmAlQMPGQ66Q
9OlcReHUWZOLYIk9w7rbvwPazvoV0kNy9U4qIgba5Fkymx100zA3ZpXksz2xtR4u
Ypuw/kOpm3VD+I7TbxC91yHc7w0mPlG54vC2kHO9KYuFDWpt6NKKLy82Iu1o+E3l
NwKdg2Vdu99dPF2ec9Egv0RPWwMETyg8rzpzBjDdw3E4cAAGLBe4XgHlkWaJMPg5
fZ3SV2fJilMzNH350SpMTefAIFANoPIZYU5rxXIlKJO4IldErMNrjJ9zVGEqfVXv
JiyRtc3TLeLrpjSNcVFFZ06gRPnOAozk1YW8ZCTQGzxZ0UBJtNHmJDbzKltjSY90
0z+yDWbze9H3nFYRkUUtwd3EHqI4b9ZKAPr+d3FLMMIKk/MpNfhLN7tdYIN2kynk
MORWGC9iVFVvneBDt4BGJX7Yu63czK4OAruWPX+CxSWKW8BN9wz/+PRB8/s6mf4h
mndHCU3Z1Lz63cGuBf1q6700BFyFtaqHNIpZvtTjg4zQSyZXQWO0DDbqDu1YFoQo
tz0FCBmsIpX2ggaz3h49JijYR0mhZuMuy6+2xCRKHnENGhwaOtuCq5m8BzAifMEd
MZOcwbIDshbFrgftJMSP9rTZzPC9WNB6aWwrBnuY0dyoKYw+qPC2tT2JyDF8PtWz
Y12fteWNp/TrrPvv9gFU3EdVUyUJHwdjGPTJZo7URLyv5+146+Mppq8Db5t6HmWd
m9gdjP7+18wQHWKJtoWmrJowXS1DWET2mVA0wr3++Os=
`protect END_PROTECTED
