`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1qrrl3dId96gbsxvB+Yi4SGHzsp7RZwjILFZCdTseXY1bo+sgnqdkMNU0WIjPGXd
491hsqX3BS4IGQEv39880XlmWp+yHScjUikv622425wPfmqGKlY57t/OVgO0mMX3
ZZemwwgrwaGaYGU7Sj43xUU7m0CNRt9rKFgN9hMWp64Ow1J+NrFwb/F/F3suy+0p
5C3MKxFDZz5Fbo8z+ZUQgVVtcDfaShuvF4s3i7PHSyoAJnyfZEdtH8gVej53xuBn
UU24WkDdoVOPraQ6pvjkeAvv4S0TdVITEqqUW47wmJJGfZt9Job7Z0zKxYPeRcrr
NtYidFXAtLj4CbISHg/75ni1EIy5xq+UJABk2dwAShFFmGm9yh7m41aNeJ4AbFUk
YCyDhTko/MoO23SJvvOwUBVzMS+QVFQaQU7dZ1HU/uG10LAkGOzqtGWR0WhulKxo
g934mRmcDHIx3ZOrToKHtGB1wpdMcYJJrYUjKV6WoD7NagjmqvaWRY/OpRe0wqwe
cWZTGHiUbcfFJD5cnZeIeNaCR1tYu4a3EY/K4LeQLR0gCD9Orh3r3am8rQmg7/Z2
f1JZ4Rgj3cHXYHCVxg03K7wWe+GusqTMe/mL1E38NFMJuDMwLJBDT9nqshWhN3WF
hIdZzUNvY21KywLzRdrGQJSL6zJlEGE6yV9Y8LCOsETOd5hQF4U8WA7k5fqALplj
SIgrqxO8XtAnYvQ2GLYfhRypHTdS5gkZpHFUvRsY+TKuDCWqRS21IWufSiMNd8Wy
Cu2hUtKOAfvHfsNa7SYIBR5dZJtyPQuUh+blkpodI/S0HTuByN0rTcNOEZSOQgqw
effroCt56mnGjsp+zApwSd5N4F4xCho/GUdp3/VURXKwkUGu4BfHIHxvEg2oQi/l
NkPERKBP5PFg1oLkBTXCdkFzQy0ETu9MKhuo0zIf3Z4ZNZiUWErD4tKHPeCWWIHE
fhlrWjxhwHE0Bj5+Lp93oFsN4q3AyUV/1w3sTkdvHk+MQ/Hw8OFooQ3PjdwJCAAk
vWz3lj79fcdY+NB+mN+UpRa1syQKk6ckaFah+z6J9QiYAnnIuKrOISiMwoPBive7
ffDzOUix1OJy6ICtN1UuJeUfAmb0LZ4BiZQmKAr3bwGhpfIo1bHvrY0vpkW0zTme
ShsG4Bdx1mLRxLSCmklMm3oBHLI+NTml/DCUc/2quxZs747+9F1yz7pn8gk1/wM6
LkTZISVYfil9XqEZRS5yHiJrlVi5dYDoCKZyrD+5mbIeFcqLpgkM95HRG2VzQsgY
vpmdQhoyN9/iYmrjF2rnz3+XrrXi8bLpJivlP/AlVRTqKBracijP/RMGyJXTCJJQ
x/kVjWdBwMG8EnZBY8vEzHqSUpenVk+FVcqqIrul2aE3PnKIq+OXINwQj8mb8qVu
No5ri7wCcBmsKrkRTLBuxx7vKo9Uil+O3oe/GZGIj350veI52iQ1KXrX4O9E+XSS
zzUGauLEQ7oquFaG24fGY7j+1bSYIwhmqmSsjnK5Dr7QY2jcqMcpE/K0/k+FVCb0
ps3+n6S/wqcUk8vi3smekz0LgxkQiW8xMnmHxOFyM+/Zm2S8Zdlp/XBhqFyxvsWc
8MS1fEhyXM/B1J25YdHblir9NeJO6XJ/NheOJ7HyyYR/ciY1Y0tZhQk4CkQSo7rj
y/l/Lbaz8RfDQxqABunivyERGfJtrKo5zhRrJDFwe9c7NcskwNg8cXTz4enSy7iV
SMFtXiVc0xdL90mmXCtMEy/Jkd4NA0oJmooXOcZIwjc=
`protect END_PROTECTED
