`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3VimcjbH60m3PK7iq1uc5EsfEZ4+q1JGnAlpVn/vXMo/Sr73RFhtPBq6qGLoLVgU
5HZ4twXMSaL1Q+YSxx4WlN1jsUIGbPKv5JWCi0NNVkRH1VBBFceYqC4+J2I1O9Wv
9S3RFCZCvCaTKcnNRiHsX8S7ZRWfSVdFioW6m4M8bRjK1ilbrwQnicdeI04O2yyO
5MQ7W+x0G/UBNLei6AOCU+qS/DqbC8JkdCDVFZPcyn45uxWYVuRKKTxpmi/wcz9F
EX+wsCmfqyhsY25kkMEs25EKkrmRSN5lc6mldQ7uTvY=
`protect END_PROTECTED
