`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pCaoM45Gv9mQgZ02lNfusecnzftEYUOE/BaRkwvrhSb1M17hD0GsQP8rd91SMris
GYy5yaV1EiMV92nsDpdru+dEOMz5f+RdJ/lKIGG5Uf7BZxBKiKNJ0uIyAqYTH3kF
H5DBwQyEGoVlMzXP1YGwAeq2Q8MDWU3Bdev6853axZO48fneXa1R0LKs2R/x0tkJ
sfNhlClzWee7gaLlzKlIBAHk0le7zFmHMevND8dLGvoJjtrcKjP6qkHL7YaVQ1RB
rQ+POytwtLVtYx51eejMjr19SFGHDqlDr3vk09PEwqvFyzthBUOA9d3lf+77Y2W4
tkJTJj3mMV1/0SqQzkikc69pkqA9YmLAfa6UP/sfJ6s+nVR7HNZeolWF9k4bX9Pt
AmIIEDLzGeepBa5GeOS3AUCh8uuinpyPatSYYJtOtidI7wj/Oid2T1U9ctsSCp+s
O2oyxEy8kHVy2aeO2zpqbUccjxzWMZWBysgzZXm2RkIPsPBYWOC99x98yCjIG8A+
4t4Y9OyAxYo6fIZu9mDPwN6GdUokZ+6Wq5Y/Ny8MPJbBLxIdjwsuATQIsr0GJ8yX
pMjzTInreQr/fECQLnkU/yVaYvaCT0QYPJ33XZvuNS8DRBM+VTD3+sk9Ji+lXXvn
Tmw2j/564TZi2KHnM2rt7c2anolAt1yx+rVQpZQ7u2FljDDGY6t/pB8c/ltWkz7I
`protect END_PROTECTED
