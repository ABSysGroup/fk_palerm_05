`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V+o+sQxQCkluwhJxNDNYF1ZcSUUPqRz76CYEwaCJC4Ai0fgpRY1RACm5ASt92rix
XaTYrAj2/6SJBB5Q13x6AUzdZ4E5urUoR1hKBz0InYdYEvQpT2rvlED15JTUJrGm
vU/YXtzDOca+3fXnyNI8OJy7zb3VGzr643cdAa3dT1KeZ4qHAukLp+80FNbMxdQa
4ut1ML67jC+ZEzacXkcbBwHheTORM9c8P54AKtwiQxXEC8J9v2Vf7z1+p6yud4SS
fcV/2F9FqEEU33XZBC8ilIkPzjMC3tx0hlJ4IHB+1tVlwg3kksEW3lH+n7BaHIOe
kUP+UyoHrKNyDuxsjyp/mLurfHFW4nEhFUFRCgy8B7LdjFdTEAYeb/bMCGCUTclD
40E8F1Q1H7KRWTQLz6qWgfN4PAzkRJU07GtTA6uGssENGyaJckugKtDYrUACEXXF
to+cm3rib8bEfaPgFyOiU1ft1kKikwGyFjBgUD1C8HH2DIipwqUTmPRb/zgeA27t
Rw1swiPdvKSVnknvS+jkxbmi2wy8kMEEeHKctTXtAbPcrLVFrB9OcH1l8TjXWK6r
Qwucruhy805bPVbzemH5cZ83t7XDcI2buk8MLNf25e0GQWUv18SV9ydbyGrjmiAf
/AhO+bF8lO2mBkhQgrD52Q6pNwnrAeHgE1mVWGRNM5/oPvDNJa0WHdf9FrLOjfnK
u1BXrqwlCxQOlIqHiAjl8HAS1QQ9ZUDqVxcAR4nn0xave4U4jm/51gAYLd5HmktQ
JInGbdpwva4RAWgpS8E7dlU3Ap5kMokWtvv5YhlOnWqwWcP6vzBmLJ6TsWxanN1t
fU+8z/bFN7CW+2szsfQAuUtXW4vfh0qNKWm3zgWJk+7SPICWw6GPYr5n7fX2EFTb
Pj5+3iKKbW4tr8hunc52DPF5MhZGtgK3h3XFsZJaBEl0O5JEXpAi818c6AKp1EWl
`protect END_PROTECTED
