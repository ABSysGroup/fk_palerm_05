`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PIQmDmY6HkyDEWFKc8FcHVJlRlGQv+MZM+ujOhLPlRbu/NsCvwjd+hk29Azk9wky
hyaq7Bt9IgMMapuGjlvV8QInw2MWcUnaAbYBLsb9duz401UBP5aBZswCzd21GGQo
4sBmlt9aS+DczuQPHKkH8dAKvrPB0i6URthz9zKR7+h3PuFewPZYJG+LYVhiyBto
EtZr5zXd0c4xO+q9ohMguOEcGNWJcbPv4At+uy78F3YW3dufYtSyUWmBLJU9HPdj
LIqKMJIS7o44BkmfizOw78HcdnvldQ3LPHkn0bH4wDYwbPjC1kRbUwg1HXyp+a7Q
uOujPlCAOZs/ebQM5C1DsA==
`protect END_PROTECTED
