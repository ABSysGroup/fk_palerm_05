`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+TTn4ibHEDqUJLCiVfVqeUhQkv7yFimx5M783Rb5cRzku/vhcw7e1OT1cCTd/txp
SvKiilqlqL7PPKojwulQwwIt+BFO5YkX00Fknb+5VPOdZnW5xMeVr/e9iQb01JzH
2JUSBaWJr9b1x9ezLvocVdoxucWCyladzsy2ps2Xw4/H2G+LKMOEFivLEXn71y6M
cHPzbikuESAbdEiByt+LtyAxzcPAiKZpR4TPg3scUi/IusrAbgl1/Y1gSg8mLLru
Rtj4x4CGjzDRaIxCSfqctAdyXpS65Gqc21nM+cb92swPmHYhnk+GWkJojeuVL0B4
1cyKoPp3OxOQLn8+5m3luJpi1uA5EKeoQviIT15CPgFY0iwr0qk+FFn8+AEi9HDT
eMEfImpuLGGk9Ny67o+MJSNgrJ6JqSrUi5xj0/BiKAafEoMFba2IDYaFnn7TUzGC
fBCNf51vFGhge/j90qlV7uMz7lUVVfIqr3dF/3uV2LqtlU3WMtBbpu2n4HMNAU7p
MHi8+yiOAt2ONLdlivmJSi7ZtAAT1hZaQmznKHt0f2wrM2t8Uv74itExZfoU/DXz
qlj7jE2PfPDfEjy5hoXama+JKviyNjAuDqnNPv0C1O6DT0UJU6z3D+cRh1sl8ril
Edyyay74Ffeha5gCNiyP28rIqTSUp5ngGx5c+g3h+qivnBw2xNZ1Wx3O0CIclgTW
whO1L7P0Tz26KSpf/n7S2Q0L0sjWghJlFYbuHytGWmYMGdbEkXm620bYe8rAhSgg
qJUC8d8F58e040BpFASC3hpbxGBSiPafam1Mzl5G+L7TeLyEToi4fr/yZVw22Zg+
ZnOtSy0e7MvUD0fjkPaHyWFTB7DMjoCIe5AMsg74mN5gBJNQEG3DaK9rPM+sr3ft
`protect END_PROTECTED
