`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J5EKkoMRPYefbUcx0kl2SbQDhMmZnIAfQHlLFJw17OYKBJCsCPKrcxUOAID5zfeQ
A37EhGvfGnjYDrNKmxFWMO+jxAzhaVPoeczCocFJksL3SibiKCK9BwKz/akBNhwi
Ptme4cycNkmajBty26fOrzSrHgY1j45TNzbCVlXSYH1gjtlCkdg55hNMQwXoSW9m
1Q9HBlPZhM/EOchhqLAqc1Redmchre5jg3RCxmm2kE9rQYH1Can+Y3KRi2GrI9/O
x3pUTreukvWPuB/Lww3IXiE7VYf9tDaUzCv0CP4TqNjzijKdyGPK1c2nlgHBfL8G
G9QYJL908eGDQNTAm7vMMA==
`protect END_PROTECTED
