`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
21lczeivIGt5ceG7rh6cf4NQyWxsTftJJpoSAib0nb5x9Oe92vWfSFz7tdeWSYap
hs8OuJTWoym0krVEkYHjsTBQukEudNZURG2diaPQ522ULDQQ8efeSE7n5DifO5gC
triY2hNIjjyPVOHdZddLniqQcT2nQAsp/5z4RnZtzjcmBMdF+6SaQSdDIlP0U1Y9
UBUtv9jVaaJgGdEqMKy3JRzhjC5U3oMaKn/tz7cSZbZyfxhucNGQZQifeZ9d9ouA
jS0wDFCeTD+mRMlHsXoW/48SHNg01oOQ7VnSOaAwAflc2t8u2lVe0JipZ8ZZ5+q6
p8+wFWkzq5e8SIbP6l9AzmdRGbjET7WJkda1nrZJOh54EJhhQR3U90NBhrBJFbiZ
Z2oOgwWMVCCsw1x12Az8X8vtVl2Fj3LhNT5vZPx2jMYLQr2hdms3tUhS4QIpPL3G
qPnqxoOqjBYZK0Q3GrhDsFask5ErZHuvBTLenaLEaXmuRVOASD2hdk6p+9Y41RRH
eOKA+ghZNMF/SCbFjOAId7AbwAAXpt5vyewcsMxPfRbpE5d4C0/r1WrEztuwQnU4
GRzHD2mhqr7VlXIMF8sHT902PLdBIdAQEBxA2n2OLzyuY1NLjszPuUTh6OSIpOjN
slFR1z0qcapIWV2LMWs5Gg==
`protect END_PROTECTED
