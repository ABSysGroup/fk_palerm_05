`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4eJ5Y3iekCpmAkm8Dyx+ze1e4B2RU/tK7gO3MAdaHGxjyDDhj9QH12jpRE5EGItf
xT4LF45jHFk80ffkHka0cXrbjbuis7weUZS+3qxPOUBEeUMX5bvisBW7AVzE9cM9
1vTn1M1XJMebP4f7hOCAhEPp67Hohz431df1pmZGB0Pzs6ztY1RfG76zIY4WqGwm
m1N7sT2XfKcvqs5pkrqfjmqdWMWhw5ROsWEVrJh5RNYlwan2xgvGHpwqjd+MtqYp
QkWmWCwO8ZQHRYnRM11XlAR8DEPouz8elsWWHGlODqBeJaCCPU+f/Q6ZF8azUQwn
pMrXHjXZRM8Ad/LIRBfR3sEyHIJxFgKWB1KzUepEviRL4w/jtpHjgVEjstV3jr0z
G3qjfLeabgxhzgKa9qq5QHUD5qKgf+kYWjwUBiSoP9zaBvMuMgkIlhVn02s4GDvw
IVgJqmrokULWctMom8I9Smj2wqPMjrfGgKNzYceWbU2NItfNR0Aj1A9nOT2Ea8nJ
5D8oJI/qHDdBDYOiVOuxxaLvlGlCzPPCbGJDdFDjMts4bOZpRAxDzgEGskgn0x2F
imKLQ4TD+TPhJtDRmDhdw3b261tP+ZVETP/juBE3fo2ONtUZOrP6UgkWI+lABQ96
1d0JGufsJly8ee7c7PVZF+jAdFgd2DhO6uzzg3+A2wy1tcG/CY4cdYZW3ReOyqu2
lvd4KAdI3qa/J+JW33URWeOVF77q23AZYtxA82bwbaetIe07sq4vWSFp/NP1+kq5
igKJw82ASnX2anvBwRp6sPNWmvkqLxOf2nhEEnFcOTdUOvTojJYQoInpGKoCPclW
30in60/eWZ5PH/oB4lReXwCQsm4YGVOF5W/+fimhAO5ZhpZ3lPS/VMTgoZrX7bKH
94E49btXvaBcKuSRmEapXH+S3spcJ2ex7pHRn+6t/eRsG0ylriPJi42V2yEALEHy
T4zqg0q+qK3V6rtWVKkz1gZ5dTj3LA5DpSWPRMVtKBNdXRZQkhJOJbqeIXLkk9kT
oNWbag58Hy6WmsvZxIWv9mGoi0MGsUFPvAlFn4vrLUPJDQ1AuskIS6blLo2fMlMU
5Tn8CrDiOSmeCeXW8PX9Jq+WBBTrbCmKzVoFGZY40Gc=
`protect END_PROTECTED
