`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M329Hysdtsb6jH82MZ2020MlLeks4w2SdI4eqPs1+CJKguVfyvarnCyT+YfAFZPk
oCrv03W8Eg5/4pi/ppwKMmznYS6JzN3NWOavpN7SW8l/kQgDgeg43315qX3XILXU
vt6zlSI+cDY4LrYVyMkbb6LTfY831pxASj3pgmDIWMyY2A3KjAVzKHuiJyuMe9Kp
n3Ub8JU+ekvgdpNAO4pGyKRj9CWMihRrU4RMMwTdPEkf84mRU4b3wRgOasaOl8Gy
JZccNXzG8LWu+aPITN8rPZE3VT7mXDifM9GYwLn7MOqtOxGqxHQF8JNBl33exKBx
9nfASgv8LRtU5+ntDhQLUKuOzfPdO9LNfdgvc+jvJyEJHovTH+O6GW0nIQ1Ho8kV
t+gI254UNY+pkJViV/K0lMfMoOV41VdfnVd/MIBTU3GzbOgXmDT++I3Lrt2Z/+Dl
5StkTT+EJXoyFcxRpEsuXcSsd49tk6RnjvWk3VhZhNgbTC2UhPeZsHZ84C0eBjxD
/cNFLsQ1sbGJGa8g0Rl4QeSC/mX9bwD3UdPNUkbSDtxKHmx2N7LvFkd/90b1xDGE
Sale+7h7rMMqTrcD1gDvGOW4JgYzoKsv2M0jL8PDGPlZ6juL0Ji2w+/wvKqeAN+7
pEznK8s0o+4k0PsMeeoNy/0rhjqtIUjUZAft8XwVhIYF2vNRRNXtg5QiPKQnbAvt
eacjI7nwoagBdhR2U5KojQZlHdIu92bTLDtyt8vVwYYxPtL3o7Qo8jbtfSyv59Do
bQj9d9VH6HtnBAZwKdLFuO+cFJoQJ5lxTqxH/K33J6pZlzAiWkfDQp8kUo1avpRn
sGjrUEtFDnaK0Qk+xvpvg+/Fka1ejGD4SxUN5qh+U+DfbYvBpqc36W1soN6h9X6y
TSjrVQWjN7yxC2cQ/R7Dh6PuMI2/Ek+5JUDTT8sDzBSaeqp+v5Wwy9aE9P0HOgam
`protect END_PROTECTED
