`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9QG+GDBpfHqf4BUcqNaEeh29rchRKoKMhd4AYQ20pm8B6MJOvbxe+iLwGunYqOpk
LXim3ZpIX5TdWLejuJCEJ50U/zMemx8ifhYG++yY2vidfGJ5o6ogeb/r9+dohSU3
d28zWHSNFr8DmKg+4xdR0pzxLIkm3ixXv2/ns5ou+NxK+bsSmGSFUGoFCmZDKXcq
hOsRnDCTtX2ZVNpzJ1m/V78WimJCYxMtC7w6TWLgeZatL7IZbpTORAXs/sYaIPq6
7mXujytfVJXG4MTziPyX1P2RtaHanFWZtmaw7zBlWc021I4F8X7a6Ny067c0iDBL
j2cEaGRRZaCBzJPX7iVZRXukMLXwQvjRf+gko1wNgEcF1ERpU4Thm3uXjtFksuuM
fGXw750bncokgoWgrAMj3EdqgqU5i4SXfzUxeOqYyBpM6Uy5wrq3axdY1gfFL1W+
AxkuZQj3DTi5VLelC7flbHsvcqhBlnCkXUncCVs5YHKPtnm+buYWfyAi4i3aLWQN
dG/ZpEgde1uokG3G1/0FhCNGt5glPNtWFhc8lcEAOSGajkDm7AcygZm2fWesCm/4
lGJcLzPAoQLL71SuFbKU66lnLEIM3WMRUAjdUq5v4lOM7kTkvayr7COJsHVJp0c3
RT7xrpak7zX0T/c3OH3ALxq4yDop6XL2+rvW21qaf+nGU2jDnkSFkYiJVw2VX2UT
W2ZwQmMR/YUsC8lnlqkWqGkHjssRLw9lIML7QbbkfX3UiIfEFIBDHHi6TcxuBZwE
fqPdpB5xcxy/Wjwos4SDupWL/aBIdJYyjzDkG6RbCZa2IJEArJOjrsO421qiBMDy
F8qYsExv+5+oOI4roMxxmgcMDfEtk8qyU8rA4WQ8jBkJZhsURFgtoamQ4DLfxK6r
2GdmcgABCWH6PfPYuvDjVYPkRBgBa14GVLggUgxBQTyP+PVzhz1+1ex2k0jNM1Xu
v0Yb7winH8UsuHg0Nq4KAZKUycWWUoZaYzWc7fqibHuf9px/sbej43JC5d1COC0j
kldU6bPR3Ex8gAZeh6YB1giJkO7xppnY2eyEWJkPLAlK7Er1bpSKcFdzFmm+rdLg
BGFKoPN3cgiMgE+KhjSvczXoVnQZ84/YV1o/p/Z+TVtW7p/y9qVExXSFhZaeWgEN
ji7KNVwIVyGtc4kRq0aYQ8KcH4e73gWb1Waof8bD1DvxcPQs5Yl3eptfUXwUKD4X
wpZOsI25j+q34UgeqU1MVpE4RoW8zJ9Tl1mC3z6sQDO1KZPsyn+WBrSXV/94GN2N
pFUUQodZkRNUwZK50psU8pwmCfXPBuw9jjG7gvp++TNg14e9AVTJ5bsnkzZ4UZRJ
XDAzAh2aWvTmBphbYKlMAjdxaRcUTvI8GqjhrikkKbnlUIwX0cGFhlT7lpy0uaEQ
75xyktEemlLA4RxVvYL6W/rtOyf0K+4LU94XQ3fzSjx6nsW0JqX+J0yKPus32S5Z
5Cd9X7LNbDZaWtfopj8iBmpqZuwGuWlN7H9+D3+5AqYxUFuGYYLggKQD9v9nPMIv
ClQ+lXp5STK/Pc6WdbffuDRZXjt/UBEd0v4fVnMj6GHJfpctMbLjOfnHLV4pcP23
/6hpikRA+1HlNacSNf/l1bV4duLNoBUaYqjkJpO8eeVVMoNYG0tmeisY6yjZG/Mb
otemt1NaYLQa/7MGSyq2Fd4aFQM2um3vtEPun5lI7BjRAGdrLxD6m0uKKkDvX4vh
eqSRkoaP+tiZ7YkGvRAtpZiL97GWc8dsCxRz1HhQZP+nkbCxUCKXH2sxvJtBZXYk
xl3Gd0JG5yu+LhLGPEn+1Ep0nunAk8LTO9Xu1oy3UNlvRJVBLwZCt4P+1ygyk7D0
VGJ6+LcWbdqBVi2n9bolJ2KAR4mTRLu9iIOYu83HugdIBk6tj5jpXGbvoBwYi7+1
O0hRBMbrKB9APjT+cOi9Fz4GvUnbGWUUIHj/tJtaXr+01iNadFki9ADeuQyPpE1L
G059ZJDa76o5+HBGla4Qu71PDZkmm4CCFKS4cGhNCZHJ4+x4f9cTgr1v69/Z8cAG
7kSIsDVXuK4uXE4euH2f1DMO3NnbOQYgnug5coMpRc+ohZLZK4p8TpD9bg7B+DJ2
G8S65yHiyBBWdoZ6zSMgkd9Zsj5mkVukyqhvMqSxNLuCmidZpVHKoCYRwpghY/M7
tOJEYXvFOmPu7r/2RGcOKQiKSjmIkj9XxD9z6VfcjHSEtFsCMs7sk0xlCoj8ndop
1mrAKYRwxbmnnINAKP3v+S5bl7OyPMTHzgovtCb82LbMrv3BL0DZJvl8UDDfaxiv
6jt0GDDaG67FebAavJ9ZM3K0vy4D5j9/W1IO0beBZeB0N+1QKFliun+Wvf/4OuNl
5CrHHeQXomgnN1kJzzjZ7e68+l0TU8b6CS13o1N+L4zqazBYwgBOL6zFrQqwAgfB
PZI52fdI26LJGh4T6MkIW/xvySpJkS9unkNa0UhQSpwDFoUqOAsbfdQ2w3ceAUBH
YMH2nYonSyKKq57myYEMpjsy4uMuv8o3IxyAVHSICsyY3XCeO7tMPZQwQ38YWxvo
9l76TQxbHOxtsAmCGj4ZeqSi7N0+h1NHoRGd27pGS8kQUKjsgYzpE2nWX8xHSFxL
MufSgwcNQpCMU/tZu7KkAQX0tX6V9wVlp3qFedSTFpLj0zrdLAcBZSWx2tQMbAFl
hK0131f3iVJHqs9YpRjgDBmQ+VlGOF4Q7sLVMRmVqra94juSrZxOHaJmOIYkF/6y
uAHU9uZsQ+owfN7OViissg54SSsfOvmuP2lVSiTxjdGqy41DuKj4iAUODwizB6NY
GJUP+1b+sLJYFVcY9SQUzFTL7KwR+CFTbXRyQfel/sG8RdXW9k8PrE84o5y3Y3fh
ZqbZysigsByTEjh7YjKZXY/4ZSdY+ij/QZJhCJtd2VLEVqSrzZGj/eFiGVfBbwCY
VpP9XVWJkFGBqQwoxhIwpXZmqp3eaZkAlPAJhmkW9Z3RhcqZVmA/Hmcdqcf47R2/
11UE+f94BVYPqi2rkEtDP0pRD06QWaMvlQL0PwvkzHi7KEgOG0/8a8+pFlO1IKMz
qGhn1FNaMzQViZNxYvwrPScH1OtsduR9P5zHVWe7jSTEMSFLPVdhRpk4Dq6A4e5w
sKYBddvsY6HV2FWSg1+DiqOxOBSBUQIIHUnh3T8RaoPL5YMdsJ1Gxn4qLSJMy9GM
TxsBP9R6oHxAUnKoOU9WPgIQXYKSnkuYXK41twiYfadT86fsTxjeb2N0mB9ceVfQ
BoOEpEk4LGxX16CxHSGbybhTmcch0YWS3UCbbssUSIMK5m9TYK1uAA8hnIr98iWF
zwuysJmebwCUqkrfvn1FRzQKsadObfNkIr5RNXKlUnm7m7fnidU3IA+7N31gzmNu
9cfGgENmG4kMDdUXh/Dync7qqfdlLl17FZLJ64zI36E2aUOM6cymQIH6sdW9KgPB
HXMWOKHOLmQrYisPxhteb3LcFFjjbG40S0Joge9vhxxBHbFIywm+dwBoH0mFtMKE
zsKROJHExPK1udwk2KEehZrCKMB1CvgA7PlhSnAPn5WP4qNbV+x5vBL44z7V1LGL
G29XGHQfZi/+kC9NGPwYfYszd1TcmYJXunXUUCyr85/sCRwnvCHltE5ruvD2T9BM
CMXIbTEEk+JcjGrbhKCo0ITLcnpqMhJrTFOYqiF+eOlABt21piQB+uBo5SqRDvOA
t0jQgpgUA9InJPmI6YBeqhYT4eoUd7qkUSX8oOvmO0NwAb1+V+fOwMzTkdboq/rN
208j9L9ZqZ3vQrmRJWLg5M1b8TARXD4aAaqByUnTdo3ojsdyHg6bV2JymhIvQ/fT
bzEqFqAAMD4hKkiDbDI4o+cf3kDC2MZCC9dha5119JUfjvD/9MHFmMnP5g6zKOEq
r1taCFTbaJNwg6gKR8+7+UgGcXbw9Bi4uIR3+PGdHd4/GaKFOriGX3pQWNVG7Mn6
ejyVUYumUrhrSLyB9u7pNZ+PkFpYL4yNTY/89XWbOAuLcYd2Y/4h5FyKGZOP18ic
mQwYMiPfTVdhjPr3+dwOHe5sjv5gcbDBNMl2nbJb7eWXMlwKPsgSZMPp8nB9PF9E
BCkQ0+yDAzIwT88D/JddmWifVzkqlDi32GB3dTLoJ52XGaRrPtlPqYHf6cETn1zF
Na5wWK8xjn3ZBh3mOLinzp8zyu1vUZHvn/+D55r4ngGP2dMn7kRXtIdqnynqiDcW
1guJMQIGGMTYtXtXB8qLQFmIgvok1YRsxGmB2NBYpXwOui7zWfMS/EIt1gIjUmu6
gh3rGaqAm8Uf8WG8lQ8RpWwzJZg09FAM07QdhXqifbTe9gpzlk6FV0rbSesAFItz
kloStSKaxeFyE1F/cIN8QfCWebb2aE3UeM/hSW10r/BCFhfYISakj+W+J0SkoQGJ
LXiG0Xvj8oID4wVCdQPeOApmXesy/eS2IMfgnmzQV1pVeqnhxaVV4l+YJkuUcEF3
zsmpc4wuWk3GmCx5RPvFIe87yriIO5ZDnUaRobvMO5meK5mjksHui70z7NbtlNPR
hDVrFBgJWdDF6mwZzIEz2LvtgkfNeQMvgi/nhPWLBRLDWYXlMRwKYtYgpvdAyvDy
DSyQID1VJLcSwoTsPRjobiyDZCSXzyVjMmuSqNQh4h6snfB6DcWk3LpeMRFDlsOw
KO2rx4APg37yUuF6E6rd3NEYc8lc+6mB0mbPxk3Tpt75wpAYlnz3eHm5FtquX/hw
jL+blqplhAw789O8RU/ZsgZfcWRmh/IByefsGtDjaLQCVv8HWXgF8nVPyqjI4GAO
PDZPbBvBaIAoSw3bytJkQnkr/94SL2OpcvI2U8xn6HHJfdGS8IbGskoKirHY3EGS
tkyc1mDFcR4Pz/SQ+pSq8pi8ApVwtgOMe5UbvrcKVIopmqafY/R24udMZN2rmdSp
orqGS86bE+VF34k0//1JDW+qIfghn8y/Cp4uBTfgSwemhpYJZpTI/Kd0BOvEB7eW
REds30u9vxkvZjw6l9RCt1YUeGBwa2qeeSZJYUFeqTJ8Gbpbw6i0c52Gu41Ki8ja
1jcLQAenH/XEkd/i9lqjydYU2cuCyXbxtRSScHXbxmVCY9lNt9J33R0yHmIrLPgX
kZ7r08Q3yPrzP4oKBS5MKnb0gTS5BjIpNiZu1BxMrE06rd1lexFSFRvQzsUdqmHj
YpJReFFFBCpmimkGpoKL+2mVyFpPAQIiSvmERCYdaMrhDL3/S2TBqtPjlXArHkNt
h/F3/rRFJVL6JdHoq3Q7/DnHp39QToz/6TBZFx32JC66AHaw0RZuMDD1UmVBI4Je
PYL+rjitacKZIxuKZ7gLATsqMUNV6U6lIpDlPj7ryxkuFaA3z+4GW/wqgWyzCGBL
lpPeQsBiMhBOg51RteRm7vITz5CuM+6ETRY6BHze8GvZfsepSNqQ3rhp7B6Sy/wl
oZsMRuX+XtubY5r0ky7uyTx9eVWtiTVgdBWhnq9TrpiWejKYrzyRy9ZNs/39A3Gf
YGjYYybuHKXK6gC7jxEWGrnd9wqqbCKgFt+hASrGxrFD5CFSwqucKoIyhQa0cG0E
K6Oa4vrsa3kttt7F9iMsllDTq/1924CjSJ21eAI0EF84yTtznlmrynYEyMuSMH+U
rnof+XUyQpPy/GDOMes1va5x7KdkNFYfVatduXUJQRgfZ4aLj6ektDloPUYPC9l5
TG8wJrnLlnGfGEWms1E3a/WeutNBJuSN5bxDXQhUYl07X+kcOic/1af4RB4dt46h
AmtbK7lcQxD+2D6jen6a8BJSV3HA5/1c+hTWXdXJhVY4PGOJC/bTJMKh52vfgLD0
R6NLwIskzLTtxMh6NAYkqQ63/KNPtXrFhJRGFASlYsQoY1IP9JQGgp8EL/kkAmQq
NCskLV+wPe9T8cBMzt63aj3+JlSY36kwfXQfT2Ci5wzTsjtwUpgt9Mtxalxa8B/X
d1XtZGho6PEWHnmz0cWLgbYltfUDqxL85ROSPTMMJae8olRAr6uzxE9hR6nwgaby
/7w5S+SRloInGrevlGBbWWlkLupUJ0SQLaAdet4auaAWZCwFJr1SW63D8TXjj4SK
mfurPvF7lii7ZGLdAgb1Bb6PsR0k66V0SGG2YZX6r3vt0D+1byeEUtW/3+KelQ06
3dfkh5Gdhv87QppmLoIFDNqV8qeRKu6sTe2h++Ion3ajELDZl5mSEnAyFlM9A7Ka
YpGGumQsPgvp4DBMzokLZXgPHY131rFTXDYKYkUakWe1HMxSkW/3UjTvT00lqJ2b
6XB6bPIezqfkDa99SUQ1AcDUthtkR1sqnS9SbbWk5Nq4iHmbO2nkWOZ6fvpq8qBi
Io0T6/qj0IeIKIayvGyhp7BtME+qeVrWoMPGPrpttTNtFoqJr0/g73VNWioWQoek
mA7pqKz564rCxS2Cn6GmkVuj0wVAewOryVh2cTFP3vffu4EwSEXayPn6Kz5RMGa4
5QbO5Wsony9YU9O3J8dTKzj922Xsnhl+z1vZRIt4YnamxdHOmPZ+og0dS/mAlAhk
KXGKKlaQTj5UbWx+6/f2Sa125jXWP7uY/GP4EbcrnhnAwhSWNEScjilKSTc3Ql0h
Vl3jIudTMVQ5WbSwLjmAbVVvyNIWPh2DV2cBbj8FJMyfiV9Iqk+NryI5lFT3MHSm
PliBKoiaDGx/TbS2rWRrCemGUusrW0DrgRuQc4bjAt1Bl1NwWceVEfqcZCAPaTWW
OqXL3gZiNlDwvNzhFV3AgiupNwG112EdbeWrs0PqkLY/w+fM3WjuLrVG9i/2zZnY
kx2HePNImgnwwd6CBWfxvolkGJy6fnr8oz0kpzmeuhPsHeR7GK1rgQfLbdY7IgB1
QXCh1muSAfLryghNu4JPcrnTrZV8xdPGrNpwqaeEOpauMP+woGR67k96k2ONutXv
mZivMXSkmICe8ZjLk19YYXTMMx6LEH+qNAK5+V7mzbTF2d4fgIOvfGNuRlVeqe28
ewIq35lIw9ecLaru8EykpRNCZXbPCX7ECrQ2QJHwMNuXxO2xaa77v6WSwvRdn1Me
E73xGbiKr8VXjF8+/Qid6ww007KExy1V4idDNllDijNd0ACHelozaTvZV8zimk9u
KenpPdpFtKoK2IJprhV+GfIUWEQQhZZ1O6pyWoETUQbW2TYdxRigIqc+rroxWkvj
TXIzFqsNGs9PEalhAhzm1yVbUgiD/Ko7DP4mmlIMXpmgFlQqAfVs7HpNonKTA6j9
fixHkQn3pEwr9AM4gvMi3D3IKkRtaGlraTpUosOESFRVKcRbUUAeK42fhK/48TXR
cFPQvmecvm1rOaI9oYepKNNPbO5qo0TRx8uB2t/jxZIebRBdGsXw6XT1NEzOr9HP
dQ9XnOKy0v+WyU+XNwdvvSexcL8fv09P0WKf5i6NjugsQGLw+tGW9G6pC2AWf+KA
tjRlFTFAVcziNT1V69ZNJW8mD5z1fsZ9r2toIArtTwZKsdPvft4btszbcZl9wGpE
0TWJHXuDqIPe3grpUvtRIcHEAiAo0rAbjZ/uJ3beHdB6Nqg7i0m8CUmLRMo4CvIG
racUXEo/gYp5KeXq01m8DwKA2voKPmNuHxXSx4XslvkuAyg1iKNUNU09kut51YVI
nFm+K+TaZ9IJ/bnw6r0o7yhkk8zcKT1FBo2A+u0lku2Gxab8709GQsGkXl4ss5ru
wwcqg71VHwBGMQ9ET5tzefXznRZ4KIQzw5Hz6L4G17CdaPOdzTaISdhhs8ttlEcz
CyyoEWVrxN14lP0xRrrPLVLc/eEBsVTMAgRicgusdt0m+iai1vUfgBcHzq7ySVcg
Us+GRYtzVd3gfv8fvlXZITsmMzytvGzD57+zdb5Ju4hXGJZYgQRZWSdrNwy+UYRW
/WqWn9VsZwbm2tsgogXwbb1c+JEFKhEVODvLvjPrqtoRH1SocovgtaSc7WuDMuwb
4VnO0FgAjBUH/2pBCQ1QI7pr8hqFbRd8OuMl1ftbQl+XxRtpepLL1XDxvJicc+89
gzZyq7OcxQM9uL9z5Xu6GVG1KGvbk2TQwEUWPmDVENw7/LD2HeOLcS2DsQd2zmFr
90eEm0bsfidPWLn9SExaxyVHrh6kkqAqAuVX3Uqvbj1fyrBgqawtBsL79zTNBCZh
ObPNIxdxdLeGrjgd+0z2d8kTYbG6kdM/tbMHWDlO4Y8WKiWZHR5DGfA1Nb/9N/rw
7V3mDYNVXjwjEFBeTjbU98CNuGQ/Crt+56TANQrEkMTRJGEoXnwMtLDnkMmcspd6
D2tMQ2mAvCVOSkjqVRfDrTX+swrJOv5sTOA95fKUJyy1bbC97xdB3q+FC8wUaYLW
hvjAjP60AT7eOtA8ete0Jj7f77KFveyyGnTaytvWik/n3t++QUZA6A5/wF5q2Mub
W8BJdAr/nFu0OvR/iWM8Z6jHAhhOfY+Af1R69yKnwUKc/BfO52bCGFTi+CfHtMoX
BnadQA3FbHKdMUhwXKl/PLQjfidGW7WwFo8RIoefNs3yJuSpjj8Vz5KhOSswYVNE
WuIE3kN4wKecf8rLGM37/bjtpNayU0/vfc1iuSoimL5ckjS6/050tIVjrX1L/tmq
T4bBAPaTegvElCXU4SPabw+uYpZqnfQ2SeJ+WmcqngZVOkdcELHQs1KB102r4Hc0
2tYK22M3B1DAYmEekrOaH7xnxdajJ2Oj9Lfkl7Xnrdmm2ldI6lN2f8Cby2APlkaQ
4uEtBn/uCfSEZUjyA31K99VZ97uSJp7Yv5cG2IsSf4WDhQL+v1LjoWvM5oWNgh7d
AQfpGWcyaGVBUEbx0wi2plan8mlobOe7EybuHtkSN3WFEbDzfecrn1L/rs3zqzt/
dxsrhZBX8nhnOWZ/JtXf2LbSbD/n64/yEavMXFT9elz8gwuPGnGwy/kMIL0saugo
rx2UZ34QuT8rbwTmkPpxlKPFYpgq1knj+NI+8Ro5TnmwKoI7K/3MsojYlT7A2VtC
FAoVVvFah8FWZrJH5+NIhan2xggbkijowXfN1rQ4IypC0VSLgskd4jrFkeMARaH+
uSj+JIX99mvTHe/mcdnMQrv9eCiN+uS9gdYnp5SOIzaDG2KZuFwdmbHIk3Y4ZFRK
KdKVI+z7t1IWBOmLQey1tZUlWRIQW7OoCNWSosKfag/EqKe7TZfje6XQBRaCksPr
3JF9lv3GBTAo3iOIquvvSu6oL85gz1KFDsoD+hU0SkVAoT6X3z/FaWQdiYr/QQJX
mcsakoE0FZYUUhi51OI4ih+h7NmzZ/dnImjsH4ZG5ysWXw34OZooUPegIFasNtPL
mihymzZezV2Qcd87ft0eWf1dzmfaINWqCGXtw7dtPCI5zGXW/qcHat042Yv5KuUK
tDs+mv0Q69sSLfL+HQ1FSZk45C90VldeSw16dUrNebxaw+radE7mCzSR5XNYz5xJ
6yU6vVB52KnHG5Dno+xwzwN0rAolIwAXaxF+2z+WZCrYbapy6XlDGdMs16gT2tyK
miaw6yQtJLh/hEBNP2E1ymlXtZ0JlmPiC+wuLjvoBA98KG4O62ALLbrmkTdBIsFH
r8lPSlKQJu8h9nvD8kE2qCWRv3Q73Bb/xgxh7ySe4WfqM5J0q3T2Kso0Q7KrRZZc
lxFP/qyLXpdDxHc3489RMJIfIf/bXtEdUrXlXLVqs6K2hNMW+qmAizQHpbtKrTR/
/WGoTuLYEQFyN4JcBlh/NpyakWIDRC3WDlIqjfzWHtqSdp2D2XcuvoIH5kdAJbj+
3+BIolhRdMOKja7WWCEPUZ+tJwHI5X0PgwAccFArFwlOtwAhuJrCeuwsJq62Bw97
B7pI3UuXemFl+Cjp+ivgYRMwUx/KWXfsCQbzsKjpeFAtcmh70G1zw601gWaBRnEH
RvfD/txk47Irv3xpiQCNzG8os5dBJJU2JPGKaPG/B9ZNgdhMrPNTykpgCePPmhPQ
0TV1LnbAV/sHeFY9vGcdIeSpDdAacNmG8vaKhrMU5oh5GYBqiAd2zx5pyvRovLPG
7e8X0ivweO9wQ27478Wjps1BaXUyi17vyoUfhQlpoR2G1LKltzTYlG79pDRHnPDv
R4uA9eVKOVZ7oXLE4ioBfacU9UHJ8e0mKNCJno+4JjNMFEkZtoAtS1VXZE18XNwV
ey0wD0othgwPUOLIsBG1kciZxt0FPh+NOH2n2Kmo8MV18X605vzm5Wa0JPcm+OJw
BTJ7qb0akhIgrdPT3LeOXYk9AaJGJ4MGmIpzwrn+uaHYyFxXLoreh6O5nAfB8AIN
fNRSA5k3eYZrNY/M46LjEuZsVpKwxLfv3Vy2YZSF5QsJI4Ko3ZU3AuPVFOIwUdeQ
PXigK9p9h+HvwEFsIwbSBvTxhNeChqIzQBOJdXcieXQZlPS7SvOCsRoibCxzErUC
/Mwhw5W/NE1M4ptXCsTMk4zxO7JTX+9xeCTOMLQJSqbE+g5q0EuhkMnGrUF8xbJZ
aTQU1tw0y1nJO0MN4g2EolrmKqfLoyTsEiECd8/rvxMMjg6vL4lgIbn9e6P7BE1I
xQyQc7ROWEUS/Yz9NWko/XFpBx6lBPuXSo0ihUaFCFMdBjky9W44QqK0BngMUX/T
uVVqcxRNRWaQ/4V6kGU8Kd5okmLv4CO/AR+bvGUu65N6/xkF6SEIIU8VAqyPTcfP
vqcumo+g/3hynipTNeeQHx/yJ/lw7kUk8NJmEgIyIwYcHa3xubuWhT0bwEO0n9xT
DR8sgHuOvSQo5wj0Yyvy6EJvGWcownuf9fCaF+QZiLKSgIuqEhqHZeeOABMCHpQa
x1gDgxxUciw3noJ94b1YgibgAdOc7yzpr31WImaFn+lqnOQ2gKnaMSiyTTUTSMn1
ttEEtxoVJ+5fvCZ3ls0MV9SrucjCZxEqE2GFLpAnFtS80XZ8V3naQi3ay69A76QV
fbKBiNKJwHRbvcKjoViPUHh9w+khf/2u12yYGUGpSVL1JV0qkmBZh2zi2i81cMGP
xgQwTAkVB+NUxfTfsokbOjWpd+7PF7lWvRwu46pXv9M2AHlFYu0Le071zHcZupN3
dCDjKa6bHS0t+1RqlPIsELXh6qIYLi/nbIr4ihExci09PgUIJI6H99DKPtdGSvKR
p1KZPcnIPX+kvWKauE+TGlaTNULYYCgt8I7nwFjrrtlN6eSa9J2lnIN0QZEqMi84
FEO+bGOxqd4UiKHECTe9zHRc0yXiYvuTzd2B4k9cGUL7pfMPpS35pid7CuYaQu1F
6H3fq7WUyyXMz5ys2NKKJpzawYycDjg34f3CMH2mpZBZmt3Niiy9aDm8sUJK0Qu7
TW1B7I/VESv1QHQYXgfLBinP9vEwQKQu2rj/F3dQ90KLE+fW+C06XZ3TqdufPy/4
T3LDym5AMXNDVq5I67n4XB7ECnm5nERcUEB412pWHiS+VfqHLT5IvCXUmbibO1zC
DQozLeIsgNDdHe1iefGaTRORzHlpNyivWrWXo/k4XSFpr7pewAATmB3VU25O/9Be
wL39LeJwWwWVvPuyc71GmTW2UJuqpeCJNSTTM3okCyovSCc8LFWP0wgJE5/c3Vay
EoOT97tvCB0VNdMNPnxvzPEwO4/5UFy7dfoUJe480TrBXe4Ja8rBOBPnm6tCJjcc
jaghB2u0V4C+9cBYXalrsiuxHXWrr5CJqy/fDubUw0MUeYtOOrxAJvdytFkFMRN3
xJcFJ9DGcdxI3FYy1Z8UF4bcpxz4NsFr/lsUFWAFwg1U0kYL/PaQHU86lg2EGMQ/
ghVI5xFRJIWgNthtQ6WSFYV9xFbTKhTaRlSMHKqk2D1uQjmG9YaxU7u/EEuMMkFg
17NOgl9csloneI4Q3w5i12Ym11UfPVpEQFTOx35JhZGYdJspQETOd0cnOOq9LuKk
h5xi4TWTQ0Wsu6IjjBQz3RErGwjsqw5SCsZfO7tmY2EUAnmanD/a3Tx676d5dmUV
QzHLLUd+cye7St3yKOnkOXrMSZWOKdPMF1xc5+OLbB0kIi0Y5833dF79x12V9Y+4
0BjvQC5LSR/HGy0+0cZGgJly66iPG3FeKuQIaGRAFB3WP9Qo+QZTG2sBRL6hDbLe
nI+X0p/0R5KgFhy3i7wPYSyUDBnbsRTRvxP0CZ69CxPtEW7V5mz9zzGCGEfkTdCR
WfYUSDFxSHuSw+ngsRtfZcMGU4JhTduCpgp5n78TJku7al7W9EZ9uLfO2KcUrbDM
bOUxNXs8rjCK+0iAM/OTLyByqJhEnlwcRApf1MgyY2NKMNnFwX1RNK2jTmKpP3Z+
FamHEjP+PvnQaDh1PMzxQePv9M5MuvKykmmB4A3pJCK7zzb/8waxmkG3+/VD42gd
kmss6f4Fl4NY33oyz/P2ZqeG0y4SSQY6Rbxl6HF6q333fXgARUOnHFBWh9OmrRiC
pkOaL08JWu9MtqjtsJHpEjMpT82cw9Ngor+fewGRBBnM5pv1vawkIzvqo2Px6JA2
uJSZ63p5qrqRWwYY2dbOvGeXApAvwlvypwhkgJb60iuX6QwprNiwvQG+LNyZpphh
Wotr8SF5IfQOe6YUL9gaw8E3Jv3eZuPd1i5XpDPUO44t5bYHQ3RcBycD5TZ5knJj
VbPMSSKZlCQl5w6xnNJ7LkkFfszfw5FgFHxEkqQz6Hz0U7AabtGfiDBkCW8yqgrS
J9jphVtCfHg495UzTeZYjX1LOWfrJwpW3wbq1pGSa1xJ3BrTai5lKyqNSb6fSoR2
LyagnLsj0QsZJRFDf6E6TXoOw+FSfgmfGaRX5ZkdGSmPYhNsFpCD2XCtEunvwRfk
UDRcuBZEfXPL6bNysyPc2YIzLWhIry5YLd9ylsJyub7bH5aFnlrxNxG/DSENp+nC
nOElKKDk4QjGBA96mEIQN3v1o8t7h2xaHG1G5ZPl+8VI4vP1INRUsmY2yRrXSkiS
aWPoGxkUwBZFURXiAXBk5f4cIc5nB7WkqSqpVgtQNV6MlvwXLouvh0dOhKJCPTKB
vLJ2TKNcy1dCRBPL8vLAELBXg/Jp3DVZPMOICvmT9zqjRXSNM5wILwIFlvP9m9Fc
g3VsgJG7eR+tHw7fqV9eMx9GYpWW0lRpOEuAGTjZvCQzurdtd7lmoSGpBo/QVw1Z
F8hmPMgbAK89YDf8jKhLcR02JFLuobqL6JCJvdLz0livK1KyYcB+rmUITYiL8N3M
jOqiaRym6noBbWc6/dv623T0dW7yvu7W8xrAdQcWRQ7nqugGsOBWUhyF45ZNLqlI
fvug41HcakAitL87PzARZwwgiQkXqNWgDVNcp52s6IKvJ3SHJ/uEHcKqprAcO3v9
4BFd6zTMKN9xQZsjVCibN52rwWgulwSER5flBDk9joJvYCKCzkr3AJ4t8pKpFgpB
3dTIucP9Oa5lPjZDlqgMWuNRIJap975jQpq6jGIuwY+ec2YHytErBGlZg/QdGSkr
+6kqTnxwkQzS1n3D4oC2vrFBoSK0NkaJFc1jw8veReS3tLdvtPZ36RmIihMWb4+9
AqIPUbpqBLcvzuPVW937WzsCi09of7BpY5Y5ryLnLWOrEjpT5xmipt2euDHidsSM
7e1XGsJEs2wjqBOZ9k6oRM9oEfixKzu+4v2yvL14cGKAc/yJfaJt+K/6MRLjUiCy
KjEJsWX2ysaMpJqPDHuuA6cew5AYuBBbs1ujwNnQV+azluoYWCI5ndyIpIIB79LC
ujVYoUxuBbM2K/1v1/DY1hIDViC3qgdDwcJtvQMFEw3cB3Wd+GNLk+26sRprEJJ7
zLCp3/E9VU7wewwERxO050uVi35FujUe7LNhEImnS6t0l0hdDZeC4eNU4oppPhWo
xEsJ5X5Jb/QvZP1mr2+iSLrRzm2Ko9tXRz1QxuoE2PlzC3NzHx1W6Slaq5PMH8y2
Isvh51Wqt94H0EEXrQC7jNNAEOrUoM4KwYt3lyRfZ045MPKJtSmL7bxjENVknqDN
3DEGdjUDQTyQAlqWhSqsjfLapqYkdFfLxI3Im5Z7tSgvoT8L7pQqM5NFje/NLkVH
+jYppg8ZW6O89PzSE8RvChkSHOh+0UqKpAUtk/GNcRKs+hexit94+LmOGMTGYiVI
JJHrGo7QyHkPtundVIQCmqcgeqPknJmpX2nco2e4mIvOXHybBZlVpJg3ZUTw/BiS
YG5BDUzUserdfL8m7RgUegEO77D1qHPNHGf3U8DQDAxUdvv2HlhhKktc+4E/nXyi
i1IMdl1s6K/wmgV5fgT/PCuvj4Wj4kfTE8uFVYQjmcA0gPwctZtN5ZL3GIcCdLjh
B2a+Lz2kVbjsyyXJNVAAWPRYvEFxR4S2ZkVQ+Oizz1ONfXd9i+FszGmZdQQvTXtk
z+Lr75QsqWUHvnpifmVTgkBlMa8wNPPYvJu3aSErX4KVpeg5FoS8PTvBy6cdXffu
ti1FoYLl5DErQBaI9etI1veZAogWBGnsT2HESKTJva40Q0hP1mY0K55TiH4bD3ra
F/V7RflpyG70OCd7qwJstg8jc94830ctSMyFLZcmZ20XClFuEdQgFMmf8ml92k8t
drVR5SH32h0WcTYBx9cq+RR7lJz5enrYyq88Ewd1UMJT0EvG4BcI+ou6/0aP5lvw
6TQ+Bjy5NXvNp/t49W5HshdpLduNwttizetrCehmtneUxaZ6ZQLHVLWst2nwcGj8
R+Q2uT2dqK3yhmLXDeNLb7Zh9aUs+O/xZA/sUunC28dUPuQno5JDwxJ+O41fbcJp
UdgdO933sY8FW74K2eHMSf5PsEkWAeT7Rw1He3pEX08URAj9WiJ2LzVkIKjOsaJ3
l17IO1hSOEh24Dhmq2Rmo1lsckyibTEPJSzM0wznhH0iT35iq3tq3Vl9R5S3/Jjz
xU44rEyug4n3Hi0np46y4rn68GIZQjykVOyyE7qZ1aRydhz0YEz6kIG2t+SrsUFS
Tsg/OmpgaGwkX4+C1xa6XzUrNETq0xzhAXgiWVi5vr/w4fRdSnflZWlrsDzURbNz
rIQPlEnVniQfMSxX76myW73JKcGtngotEb7F2W+Q9NF0kjfTnpVrHF77wnwEqb/u
W62BCDkzQIBaxAZs8HWUYbQ4V/mfei2PYgxOyjxSc6clUzu3aHGj/rPlK7qw2rwC
mTwZBaPu/maTgTxKkSGAmOIfuPkeGlOMQa1Bpd3sSnysu2H3Zlb4WUy6BtekwX6O
WDOZVFe/mGhc48nHKiS9WiBqhTVb9sD0eQchaBbamqN1/5trtLI3Ldpn5HHmagcl
bum4BJ50vqOHkQGjYNSoH2kM29Jz6ObCnT2bFARpkweGOMifpkqN+lzuTQHmpOSO
sXhwths30wBdZDTaWCYBRWUfa2MMYlcZ0NY2sX6uLWmAX6NXkF52jMVg2PEmVTZq
vzYGxady3zmWugfLL46Zdy1vKsUf+r1UsRNjDhoSETS94sS9jQse5akZtPbGVq2d
cX2+aVHL0EglNZ+d6maqybOWKR+TuYMZx/9BLVPuKLFfD+dsrB57F6YiCv1M4Ddn
wlym3fmH71iHjOUURt7wxlO/Tu9KKO9/xp2pH2poIj7sLPvA8YHWINOlwRE9iiu9
z2sHk9TqQMUc9MVRDbhz1C2l7sdVkN3nJJaY6qk1/2nTtYLmJHlQmDW0zMpA9puy
QekGYMFSwjb4+d/th8Go/A7RJxLk5qcCIt6xVy0ykuOy0ymJFLQHuOtc+7IVnPLb
BpcyWsN0KFkPVTpg8iNEQPAqbJF8rGQvBZj/CAdgCgvjj6X2fFzMYQ3H+JXLUusL
l+9OMuj3f3SSiORD6t5SWrinHcvX8u+1HKNewaaBqCJ4aAHt451ikGO2Su1CQU31
ClZN3D2KRWv7Tk69GzIypADsGndjI91Gs1QLklBGzScrK8DbmX+Jr1Z8VZLTfCd2
U63DS8II/c8yQZy5iP67xt4T5RK22j04deaztQIXNFtfitM9p73gpl3SPa8J4Hcj
tqvochCdms1h9yHUpBbInEPy1tq47YhZaTsnM7/EHdkr1U7K/HWl5L19YFDOT46Q
CpTQ5c3f1CNixrxL8z/NaeKfcaZ4UUuhmoj9CNWyEsRUS7vb+CRZDFkTZd2dCWA1
3yD9H7X79GT9mErZNS2+cbT9y8aHCrTrsGdRUPUXNIrznQEtyqZcPO4k5VzJTbRO
OAQrO8m9MKPI4CG1sqEt4S7iqchJ5K6CuiV5OTEmFxoO2nGzCmg9xg1AAdAAiVWt
1QbFAc//WnTN9a776VgY1WoHRY4Yb2xsB5ZfaJ+iM/qqvnSTryKqLKSz/7w/2ynK
tx53WKD7Q0mr/XKRUwj9AL0vayOh92TV/s47CxM3FbIbPElEs5cdNb889TowBw9j
6jzQnr8UTeNDnDe4nQTQKnM+6LhlhNEYUpPqzqgbLxijV9q0s4yZqv86NbvU36yA
DITq5E7zq6HhD2Jkf7LI5irdIJvXK8NhPucP/h1Lb03yJTp+VEwb1WOLzdoNUHHC
9t623PDaaQcpsE8SJKl4emh8GjEIU89M41Y+OAjntqrTOGzdUbV52jWyEi+W3rU1
g6QMord/zr2r15o/+ioWh0/Z+2qeMifkG2FRXTsCgG4E+OOcIV2ZLe1vreQydxQV
H2cjuoKNNNG3tgBDUcBUSqr2PoIUybarmRl/ghiH+l0LS0VVyU2Yshhb27NWnbLy
YgMRD2jnB0ZAq0Ne3X3Y8f9fpimCxcujY2gDYt5pGHeazHKg8UQbGJA0tXUhM0R3
KmcQ0Kgy/ZCqPWxhSZ6KNDKHWaDqogsJ171skmqrir1mxKaqhAWc5OO1d3Zx3gPw
3BPrbkoR1MJacQjKpnCnnOCtKtPw3RRY9Rp2yGyH243dG/m9HzcXqB3ABTxBuCNb
7CsM1aOUJ2UfXuevLPztN0Zn9O7V5/raDN6tlf8s5aZQO4PLaeAd3lLLtk3nFLXv
TCJiaN9Ut3EuYQok7wDw8b4Ez3KBsBYt8AoFmbX7Wfsh29VFk0ZNAkktWwhT7Fn6
g8LlXcdcaCH25DSctOgt4d5JHf+JFujYzEmqdKCbkxP/3zUBj39KJ2raQdGkvN2m
32ocIt0o6vlRGrMRrGekTF1SrgZSBIAtLuVqu9uZY1MLJ86ax7F+y7zgNc+ry48h
lADP0RJJW3tPP0xb8D3/BMD8Lr6g4wZRPmQbQ3VS/pedhZbq8JCnQZ5qJBDNrduk
2mzg7dNuW78hHoGkrqeT9gnlTy3fiY8nWtAg4kALrmnmTHO3xPcB+0os/F/ZjllO
lPSENXhB04bXyTWdF7n2P4KdaW2qIgijBjWEGnKCXiYM+CPVj2xeOi3+tpAl4dh9
/btsyqVkCXjrpgAcVSR5tAL6+UEJrmqm0xSTjjWpBpBweq2dd1l9/dp3KXQ7ZdPB
R3eFiQKagsYA2n7LQHyncZIcgbbRJ95NeDgDbKDRoytwt4eiacaEtfcLEMO7IMxq
mYuTEVw5yLb8SLcOxpZ3egqPRyFNBeQqKj217sTBmMPonzMXEj5uKD9EdkmGSeVj
u4i9bIcDy4WYTGwd/Sp0ZAooTa95jzR1jOmWZx1l8m5ktOLQQeXNckO1YdA7khu/
/WXVzX4XxVspgEzE5Ic3pY9bHrP+sWnmphM1O13D/v7LDkptfDzIPiYpbyzijKcU
Tl5a2FPgnF4KFjtT2EEeMaYYiWFB+0M6LCPR0Yv6skNzwdmSuDCciZKlGlFzxx10
wZ8sf+JvmF+dlT9QXEaBKGJQ2CDeThLeKWHlYlgNyV08mNK944tE7//rayd/Rjvq
Xj9oenShUnfYakejeN4NLHr/guAsGuUjJ9Iq/rfTMsXBgx8oZ6P0TQP1wAX5U6YQ
J3UQfJgWXDhEfUiNfLH/B/2sTuCQpNi5TlRz60EnOWe7AP00CyCFlO9hzijSjCbS
bgtgX8g06kWCjWerFfDhnEiGgoUIJGSoHe+jSVbulFlk/tIyzh/qeB0yMlUgsoUW
McaG96UMKpb//uBPC4ninuc6OYtIHuJsHiS3TC1KJXZJ2kphMT9NI6QMj51bnqcg
3CHtj1sbbA/mLonnNBoG96TWr92u1OcxuH/n5qYTDYH8Acbg45LkluAkJLvXnBJY
BJ2LICv+ep1/RwG7yNhNKfSYjRf+nbHXDIt5F9eujhYPU3QXFUaVOthNk0zjvotp
Wa+zvKRgAskp/bd/jTKJReMgPQqeHIrhaWmQwP0BIY16hKiqqsn6PKDSNcsL9Chx
luHCKQjbc426lWGyuOViv9prKaiwzihOUJefvmzBPy/PVEzfVe4mW4lVYLpD2mmD
KzWysrEiHv/FLfObvdHtoB5TOoSwMomfBxtYEULiMO0kbUJoA1E5SjBdv/bEFj1f
0i/EqeVgc/u/0YhqhzrTevKTAgc38NQmQROhwWJgdA/y6M1nZNn6L9odfwKEaa8a
MGaWSHNnVkx96I5WA0+BmaveO+wVZiEdU1HEgnDhreoK6a1vd5UDiYICXsAcIquO
2u1sEEoEt/UygaA5B6OanBfSOPoqf5uoYtmuL1djo/2zZ7cLm06hsWsLO4PKhH/b
jpHF9m4vB0wvt0Z8grddQRi20g6E2xlrcytQ0VwC6BnOm9pLCn5ZVLJqGBAiBsHe
b9NAFz2uyE9TOiHhVxzbkin9XktiGgWNBBxgsIXKdM6LdGsXCNpvrruFxa0Z5IRY
ztGE9ZOysxXDSjE4UAieJeqtjSST6PduuH7Jf0l+A4cb25ewcFSzEqhU5HXJ2hq/
mbMayM8u3lgdd6QH/OcBYqAA2RAhC6cJy5Tult0uN0fFgg7LMH6DCJ1ep6gCaSe2
z/ql4eDgGXUGWUvjiKm0l9oX6xeYlwvkL52JUp78pqsiTNa0u2E0UZ9dy6v7zUCg
uz6yeuEqR3/a23q6roxSXxBpTCQBsfkPssn1uC8SA4XvIdNGZk3Yg75sWgz7hzPE
VWdx3qg0T6MKtXSr8ZFlm/sLz8h3qS0pFMuzTLmHa8Onm2tz9epxiWd0sq1RerO4
l7qs4mkTliM3G/nAqgQta0ZpO9khx+M/rT8XGam0Tc9pCN8/k4HtSH1cwKnTtHuw
Zfms45o613LaVD07fMYZ+IFNR4+vE/3uc3gHMVl+ylZ5KMZQKP5mVqC+/p2TUGYw
1YEJTYY17xf6STTuozEhElJtockYrGIHzl66fDK21JFhCInuaNzMyR2DLz0BE56Q
DA+JQrZ/UK1GWe/tnTidGnGfh0IjQCOhg54PaEbLtudfVbtvk1QrxfM4C7mDOQvA
bR9SRpwWIotg26RD8F5pGkywzmS2olS1GmaPYmXnSKNezrLQfKuF46v+4sDa00wT
TWJXp6ywLHiMirfdcgiQrxUcQAJsPV9K4OS8H5MQOexnaTRN3JnzlEmaHQWC0oUY
XKdNEgZdYwbUIfZTiDDH72+wruKGSQMnVqszfBZ7+ZBRjZEHNe0zjnVW5Ky3caFf
gNRc6k5ZbaXBPol33whXz52KoVw7RQmtEdnqbq37z6BSOT4hobkaom56l7028PH9
YkZGTmyy+FZEe8KoHKnKa1QnkJxvIqEc2s1uLQAzn0AC2no94CCeCxA6zH6vFioN
77dJV1t5w/f/HPJDwNatAXOnqxns1sm4G2132k35r0gzmV1VUts63iWH7LL1BgUq
bzvHuKoFYCT96o+MoCvjEAjromC8uuJMgWXg4gr+bujkKaYsG6LvwXRC962rY2c7
2Sr5cZEMX49OQ+lCy7SaB8yMqR6dl7y5LItcCsUHUqn/Oj7ZY83i1fnLqGwp9caQ
Qpz0+yG7xN30bK/PzXhBT+2WXIpwG8Vu+D2jX18cZuZqZ/uu/sv8U7NXzBtMlrb9
IlTotdv8uCTiw72uWRdJBG4/xzqvmYRHlo2vzfKRZiKDQzQ0t448ZC4cNh22AhED
VgiMmx3mFZ3F7rkYGv4Ji5xniWXqAAJZiVcKiskj4nIvBWb/iW/2zFu4i/0+RRKC
c3wbyAbmyxOiCF+9IzLimRdH919a1Rk7uwC5n9eYmGkIXUXkSRrcosZW3a4fdy5U
fd9UZHGngInoHPe3+j9ieYA9nNvlej72iK/DP4GwP2ido/xbsTVyOjpdFlC0b56I
MjBSdOs5tEo4BWy9SBJOYR4mbWlNFVUkdzDBv+8QAJpGZpDWQ9IG0TyPyYjmZ94h
VHJxzV2MnX0SBNrWxV9zYoOVaAAeY7UW2RHULzDvXXe3WGfRO2euDNwl9Vy5t4DV
G13q4qja2Dy9o9YG0hz8bfvMCNns9E4qbWNKaGDwgiqFFG34m+2cQUsGnLKH40W7
HKfIIreeW6UF3cnkamko6uA0/fVPzSV21Rq7EFtXs5u/T0TTLhkQv3iC3lYfNaP2
+P4BMgNG+HpTxSNiKSnMVVDKVLZf/23wm4VSjmS6MqL5O57G6TeFovOm3BRO5iuq
//OYsqxL5sFLj6NR/Dk3Bm+DiW7Uesyn5wTgAFTCcKvZTILqjFa7dkg1JMyUs2Q3
dZGHBEIYqmawkHO7Gjfg5RTxDVzU0mNhf8LeOqTchvLdG47C66++6h9s3maLCGYS
Vr1oLBTeRGEg+boGneZBIcuKUJP4f7Ia/lynXJlj3A7XLw1zYA6LGA9+GVVPMms2
TDXEQQSicSH+mbpajOv2aj3n9m7g96R8fZ2h0j/mMMvKQLJ7FCRfqBo0/QnWoCmV
YMvh9t4ms1I0pzReHvtM7slU05GPffbkXQlSXYCaHDODUmSXm9EY+aCdODscIeXZ
IyNdDxUr80ZREYkGyhKHHieF+ieAJqoPVPEFtY1BF01QHqERNdB96VggSexREsLj
k8/wieKZUhE6VzfblfYoWK1nF7XN8H5TvlGfrT/6kU0wH//oj6dgjWt1ZKOshl7F
lk6l1JyFOg9/Hbwgk3tsjU/psv8v5AoU2nrZjLr8Gb9iNUajANjU0DB71lsk212w
ZL5UPF5pUxmdG4bezaUzYU2IeKhiSNpfoVb54KvZQjDeURxyPt1h/Y5fk8ck9dsq
6iuTE6DlTEsxt3ycZe8gyI3c+dZY+r4euMBM2AwLCsdZ/mq+jF14GJyfuXI9qrTG
poy+zrmDjmxGG9+vp6td/x/IxkuYw8jzoVW0FtUOt6rTEw4hY6sbsugQhcyxYtKA
mY1A/e+RDY+1XQuo124K3dajAo72wdGvJKjcODogQ4XmOlj6rLmmQu9PLvg4rrhf
maYXVsv29SVlZmINiCUMUXzIrBcw7no60rM7Ibduzp5eTN3NK7DJVW1QG87/Medf
jmN2rt09EmxskvQwUphqvwfuKBMPs1UWE6VfU7jJDx6KuuFAwgioVCj1kBqV4/Cj
UyrGpdUU1lxRosZyWaf/ZFjyKLzUQhpDIUQLpLU1nxgZiLHfYr0pcGx7iYhHNdbB
fxeh91Sl13KCDlY5/JnP0CzOqT6JKnlZVA9oEEiRjprXHUJ0lTUuirVV8a/dO7NX
bnOatJit4brwSVwiARTymcilv6wheZAGP0Wt9p8zQXzLfsGNSZjz6fm3HQfWVft6
/rkXaPmzATNLBehQvLjWd3BYoADO7QZEGM7HTJ1PGVwy3VsplqPgVFaIJqdkw5sZ
OXDc5x+9YVFNkPPCQiExrZOocEYKKh3ZrZG3aMFuF6D9tFxmZHDRC1S8A1anFslg
Ms6oap+Ftj5YZPn96lSDkSG9p8GCc/jj54r+VCMTGF5ilMfnmFfCn+1DeT22zTE5
81VnigiWoh8Rmi+fhvHfEo61h7o74B3ERDgutyF1HEmqWbAQGj79DiGIy9bABI+A
PGQRCleC1jgIH3GMzPv8Pofxpj7iP1kpsobiIwL9AhxzLNts7MbMy4K/IuHtuU45
Bbza3YuiidkTuI9Rm0jQgVSXp58LSdsgqb97mCANryvifGrG3x/oDN/pejYzfxxd
oqY/vIlh/f/emftqyxn9rlpJ1kT2j1ya3B4ezuEcpmck+AhvN4rDug8P5oRZ6d9l
PGdKZzRkuPeVo8DdjH9oFBXdbq4mKVu72GsiTsYGOw9/ctfI6e6P0YeFDjv4dRmF
ZUqClqtfIkaY+zE6v6ZT8jqBfVb/NViLs5PSEVyMDnQrGPASFkBXsLv5d3QXQHE8
eKYVKNhSygWjUybmMBPfAbpWcKJkhMNSY2TWTGb6HrrLv21tdJqTfoqnRUtIvV6V
nAkQyiEbpDcnuIiVI7uf1hWa1q/fv/d3mC8MwBC7v29C9i+0wQDM5WGJciarbaxc
nj58VwFV37kigm8cPEpGjMDcFMPjc4veKWlhyAKI8pVaNX+ZV8U/laoV/13bvnFF
DmPJapqOo7g42QHvlEGNYa2jwvt/cT3rqPh5HseIeNzVh/5Y+Q4u6VcyY0Aq8NRV
kwebFXjzTffRjHDZyf8wShPwZ+C9yoHCMqxSXFzpL32sIeYbw7kzM7vU5yI6Bqc6
mEWKRLks81bj6BMiLHLup7h5N3/rSLD6GKc3A3AmOHFbFlLFTX/PsaQ9DH9Tp7sJ
E6NztbAUV3YKXuTe0gqmuFJNEvmENFvSOIFHNoTexEwrSZjMTSId305UzMQCcei/
BzfJ+NribXiiTeA+pcclnQ73eDQGVr8Rut397LuzocqkEXvRdmn3bzz32LIP/iEB
Tou9Gsi90sPww+DcJkgO7vP9QP2XtdfytyTldus4wSqdGd/4E7j23ZfKTfsICJKr
G1O45HFkZRizRwkQOMWF+Ixl9np2A4DLDKf5JhSKrtcOnPqYm8sbEpbJRSI8e11n
P4jOlhx2jtIBWElXZbWNEPV0JA3Hm1lByzGLOrIBTHlgW5V0zGgDtMOBKKSlXBPP
/wF4S4Zru+xPRjgcHa6Qh3+Iaa+zo6w4Me67mezz12ru1bLCcJpCwBFx2QCIzFF3
+TRvT9OZlRoT7iYeU45gjNs6stR+ATm+swNDerDaW1Y/X0HuRmXvmyOsxsW9o/V0
E9thmeJ/RXjo7k6EamJZVjqHYYq6q0SsmhpRBX48XkWo3SDo86yx+3L3kEbztbuN
iO7qgSl6Wb53k1hHxKoBV+lANZQcAN+UVkvnu267aGeRfm2Y5XGWD93psRxQImbz
dYCsq4D17E250GLGg7+x9+fONdJu7kHuuZ96q2W6CH048Mxj9O811CQKW0gWjxJy
CaPHzArrK9+fZr0GR6GHCvyTUWjLeYIODfLQCVLbvShob4PmlI6lp2PpLYPDpCt+
04Vwq+8fWYVsuivwGAKE7JDfcaK07NlbYVQxWOdUMhI+X+RDKjZENlr0H/tsGEAL
HwcZF1e1kQ6zxlQOAtuZG46uL7UGsuLaC9APuQIJD1nRbI0rn3C4oWMnrESszuKY
Wf3P1wPLPZUuFZwJTfGmKTsE7iamPMGrViWWIe2o4WhktNaT8jeQkItkerKHjQTw
u3hAOLNJg8uUWoA9WdBffQA8NqwUajhp8PZ+ryUFx4iqUPXkgu4NSlYgARag8Qys
6dpNP+ctD3Jx/OvSnHKviqLFRcZzRCjiXiiIg0bDN8ykc/ZmwJcs7gRfdNpqSBjG
/rruPmZop52qZC0sg3+Weqh3U3VGS75fQtfHiA5oSMxCxdKQTAc/sWzj7Zbk6bTv
rhLFjkAizvlhHlDPFRS3WSgvJFDJBYt73IJ2+TXClgvQpP55tpvBRbj+Eo6O1uGt
E2TDohGWtw+9m5ifbV9BlX6lVo8uKWTxBe86OPAsv+V0VN2G5t+CVK/AWNsS6FFM
2XT/n5yrrJH+LuiFe7JzzJcoAFHaX2mrbnExHv0YUoW5bbDVSjJRbYsG1OHRBX2S
UXLaDJNJExlUzL2NJ7YXXStNQtpVtbgmoTkR2ZbY5JNba3b5FnddPOJdT9PT61z4
/XKMsYubRU/PQ+GzSf3bnA4hY7vANreDJZBPK8Ve7XL29qA+bNZwPCUyEqFqgxum
oxDY3tq2OYrSuMEz9v/8orbbDDE8H7dfMDNS3E0fsz5Z7qKq6CeTBT6rARRhJzeE
+mvz96WahSXYYuKQ/k46SLC1529BEE06Sg/sbS8x/mr5zXeI9VW7fPyRAgtxMgyM
b1BBwllD0iYOtOZa+ShGvCgRmtJavIoAjtWEbcxlKT+ir+24h+7z6aVVi5bx0y1a
XCw1Ei3eCQHU+Uf+ESXavgtJxjSZ0KFKAJ85CPtCdu4H98kAk3Cvcm1abyJotb1e
Ey1r1Df88Jcd23tZxU7R7uBLFYMNJmEtS1x6TX/uA28ROna2I8gQuU2zmHQ2tcHI
2vzj2DbS6VfQ1Ua048Mwt6bJ/+djKBSDfKoWi9Wwce7/zZA9putAGFn4tDolTIXt
JCPRZR71MGjPb/EDX9Cd4L/vIOK8TZVlpFPDek7GCt59Tde3tGVztSfZ4tRugC/4
EsBOD+t8s2rbLvOEtwvi7Ud8G43FXb98wLXu8X7cycBBcj10MRh5rUT4vRCI1rJO
S62+aWfM4KKuvQgxmv53AWtcfAYr/37iXSuZCS3wPKmZtbZ47qHP7EYRXyOnv9dg
yPmRr+XkFkJVXVZvVFiLEotcoIFPd4rEr4KdxQFYhf0R9+A85Aec4CKV0Ij6EwO+
JTDG1HmYgxRvB0IYg0NZXwhDH9b2MPIEYOQDgW5Fyie8CaIQyzX+7+uTNbQTwJqj
kjzC0B+UAbE4KD16WEWf9t+DVZiUok+zMMvc7T028UjBCg+4USrhTrI5/p4IyHPv
mq76DDuapsE0s6R8XvQBzJ5iZT87gTF2JD/hUiPcglvW7zcMrG2Z/BEu0p3zp6t7
mzXNzgojZxV9KDz/t1XI+iHyybq96IHxUc0kwegLaRTAEhyHdSiv/kqsb8aim+ob
XqGm0MSO95uD3lf7SsqqOTLGrh/lZrY/yaRAolFRgc2J+FmUe9TosWaFBFlzpHQp
Jz6nL6hr/N3Jr0mrdeD21o0nHkhds1kzaRtZmlbMlicqro8/vBbredvMvQgBz4my
OVjAH2DmnFbLrN38w4lVTiELIncFmkJKIAD31XeQLMEalY5z5NxnrT4gqVSMx4sY
xPe9ngp8budpC3UItZyuIf7J755deviMJfst7d5226qzVPlvm7gy9eIDI5UvAbrh
ZumsG24gUaI8SIuR/PHRQmmjOlHlqzvMlJwiQmNnlH5nwPiLTX/0Pgne6M4S+oML
DxwyhKPn6fmeC1sfYhrJBX0HOhLJ2tKGkKiinj246asA2Pw9/p8y2a28XDcEFnKZ
MlCsbUa7q5QOov/dl1OsBCOKfjBmAd1okcg3lhnk2TPaSgKhHRr5+OpmowcqRZUx
aL0mmL2uf38erjc1XMBVFk3cxBz+i4J2msoyjPhFnbUV0cbsn0eV8eUE8DCW3FgS
3aj/Wntdli8IS6Bbepv7ez0x8abVCgnr8KM9xE0kiXILxC2x/y8N/NEnqzZvJ+bQ
Zzoug5NG2va4TCtZyAUdupocN2wIxNHQ4zI+wqkO00PcV+9OFWYNeSQhZG3NTUku
/OaAxVfR3bSYFP0vgKBrXfuGSRLbUi0fsBt2QiKd+rk/pl6L2/GuDN3r6GNaDVB3
uYDKmc+1JwkKYDPVwU+23HUbyyqvye5QyqbaQOJbmRGIHr+tzUJiiFWFbrTu+apW
W6N0pQAzL1A+VyNUn60tBqCCHBP/zV7nQMQuWBMZ9gHifk5eHe25OyY2854qjWdA
nY6VWP96a6Z26rqQDSBcKHf/ByZxwqMmDV/fVgk+nXMD9IWtkWwYdXjBraEZRuOL
cdjJSNNPeO6hHNR872MNxS77HUA2d/DPtdQETZm1Ttj002by77u+v8PTbClTrZgp
lhBowUoxyBl3AmX5hUdMcsTb/awv+JoqSXair7R/+Ez4r9xhCCvjYTHc0OTxWhMG
8X64vNYf6SYJd00KgqdYGtbMIG8gYRo0Lpv5mD8BKyvOWmLyQWEy+zWt9TpypUut
MtfcRHdZa63ESd2w3g333YcHMOFcp84PJqEJKrfBaHsj+wsHRJBsresnpJWFsXYe
lBUT4+yD+9zT3j0p+IyQxkFS6SQubqm1gBykBix/nvLmnwmGCYxhE6mU3N25SrEe
SsOuQ3P9U6lb10rrUsxdHtFcTeLDmAQS+gf8xFHMgg/Po/q+MZXjpTn0ABF+Z1ng
33EeNpjfzdlVrjaqofRgGonXphMsN/DH12PDNV09A7suyQxaWGEIvkQ18U28UjYa
HQn4JXgM7DT4Ua9YsWeU7noReR8zcbfj6LyQK1cda53Y/9HUaoHVxVRE+0yjSrIa
QnBriPTfYFSJKTSSGjDO2LIpM95JPTz/KMcsj9IGIo+XOs7tbDXYKykMCGkpZU7Z
XOoHHx21ocYHKQB0DoTDQRYTtBFrah2MUsP6orT4Jx+/kUOWUacLb/GPYRIjWpxt
G6kD0aCyHRGXEJOr2KmWGY+nGxk/l26iUaVuy7bQLg4mJqUH1cyHZ6SaerKvQyLc
Q2HRDCsCNVnKm0H5fHqMv/EyGQiG7LoRWPlBieE1euOflXm6gZvBQit4Vtc0RRB/
rQukB1KsOBmH+7GByW6pRN45aPXmzv8AEV4Ij1K3uQoaIWZitGB98TJ4RMjLPG+t
dwZGh/LDqrsrkPIW2GGhzhBzozXprYHTn8SxyZI2WEgO7NUTZ5hwBBAbBVmYp81e
1yFd3+Gxe4SeT2ZfOyk349LJwuuRIjtfhoYvVOJKTjNXad2wmmPD8UhVNBSLLOWF
v6izTByW/Nd7/zpZaubaoiwEssW1Lu7HOXtjVW0vlXx4HURFhp5nvM3r60Ox351h
B9iWk+leaQw4J1tXA4+0en7BIwXyvFFi4VWQI8H+GCGJHHDYI6hUEu3TuH7zZAae
gf0t62s9LO7x37whQPmkWlgwDiTjJWCNVwxUVWfK+TV6qcKW13sy2x4FXuDW7x8Y
kc7rtjINfveNNJ3Po39eUvymi7t3bYnoK/P4kOE/auFJ7iRyjQqzEUovo8ZhZE+z
t7bh5gVFxvisyPfU48eWhzd1/Xqlwl2nmyHeExounGWt4AEWO33dEVb7QTKqVUId
peo+CxdtiOE9NbwU0KBClF1E4XFmL+1QWEU4FSDPQS6NjQavEVIQx36O8K6eDmpS
dmAq+8lxsS+uHtlow2J0+sIAVPV/JWyyU7VkSx8pu4ogLs4bWQTWGo/gcku8Dl14
FWbdMor/VGeUGarv/bzX1yg4WncH3fERp/n1DSOmrWPpJB2IoxC5GNOMuYqTwOHI
oII9/o08ECZ//j04D4ufrtapTeIBNf+dg9I/FvNrqxznOv7tfvZ7xkRHyKrNA2+x
iD1GaZSlQeW0jqw9DOsUTa6yV4mFpvc0tUJW5PB066Qt5GG4+6iogzpfy9Vvethw
0op8m28WxXWAco/uz1AZ44EjlfJRLhOjuslzUxJI8V2tKkpbp3OxuKWCSUNsNP+Z
/4Lnuk5V1stO5VjDn+/piz2bBg+kcqBc4zn2GpmeJbKCELMjH/g/PMTsrMQfAbb5
tsmie5EXAGrmQ+mDdoKF+a+Yi8TlhNHIpm53Xw5LiO+66QsY+/e2Mytsk0gdTj9M
XE6P7uCMdSGli3uJwsKUMLypaFZB0jgQOjmy3p5jKqbLSaIHzTkWmitpb9CbFK98
xRSd6X+AaEHV6RZM2PK/Hh93jWE6mdnb7jaTWQeNVnAReK9CVpTZbnQDHKezq5Jy
sJdMAKUFYNPPggM+mbrhJh3UvPkczGcTO8heeHkzNaAUrQQL2bnhmb85knEzr2D4
tegiqeiUSRPBq1nmEMZn+mv3ezFzSn7/w+PdQ75BBc3+OWHmIt0qyWjO+cW6FSoA
TCM7j5SjlwdWcNdlD4fUbfoDXUIYQVg1G4ETlTc2mZaJtE2nTj9tnoSq1JzSpogD
+FBH/XTgu190L/nNOPUo9gLBCnSgyInxt34oEgnEZVlAkfKAXqIzwyJ6aXWRkJ/n
IP1u6KIZmZtEQ+6e1yKhEesQNjvzdgHuUpzbFRrRrCezrMazMEb/XjZ1Lcu5ovFY
W5NhuH/VPomxzlcbOpTMKi7GTCIhuD/dCazgJOpkY9nTmrwO5H1t3LQB9I2lVsag
d+iXKeG90LpXqtZ7wnwgK8StMorihEQg4+k96OD+JQSAbc8O+a+lkkXf/F2YuwHx
K0cQfL4GwHHNUHBurK6KNC6I37yZDUprBbeHfaAcQcqKB9hXtLRY5RkWDY25ZVh3
8ezsGQnVcSEmZEPTO++cITANzkIm96CNmmbot8t/WCa3u+mobUhGCWUs2e6kDPbc
opXnmIfUp4JKAs8iEvO1+4HMpavXHkOgYJ534dJu7wC0z2rMHQl6AsmkR//IoMNU
8JcD/28DOnk7h2snZhcz4yCuzcKPgALYhCxEeKirKkui4PD5kKiCv0kX2dbJe7yF
F1Cwfj+m7K9xKkIornn6Nq9WOdrVS/x0E9Ou2Ao9XAd6wm9kFcYZ34mGPOhRsfZc
+ommDK07oMXV6vY2L67Sm3kbDXkMMKkqOPYEgXgeKqdFVp/oo8Fl15TJBFuysdY0
ZZdSYjHt1tNaNkZZ5crN9EfSW+uYPV6JSZmlTye+jjwdSjcSyGfPkwCfmlaOKKJ4
3WMYa1z0xqt549JDyVZQicAkRhQnIhAjcJfRIsp9ELP6BBtHoLeKYmfgbsjF+SZB
JaGYp4EcAu+4yEBDl/4EpZ5Gto5JnVW+P19Vo81ji2yaLMyo4TMnODR3pzVtu4k8
LmUsGBse10w6tKtRN8Q4/9XPZD9R30mxdGygVNVrObS7t1l10SAKQgqsX2SWQk6w
vAZx5EF2yn1wTCF6h0pTF8aeRHMHj1YmBZCwze4xUaDCcMG1FvqX85m19Bl7QEIz
0LH3gWvsyHF/mpKXovSf94srEgeCYwgNxqLtA2ymGxR+Ig6MTV0y4a5BzLc3Yoq1
sIXzOsdHWUamcbgTDLJUFDPlT8QQWYmNGx6yhzCVM2tqR0nYvr5F03G882zv5G2p
xWqGQuIMWbUwkE7IkN2uP8AS0qyw1qOOW5F2jVrU97XzKblj/yPUVn0725ozUsuM
Hoqiq9sJggc+HVoMZesSOEBVYyzja3h2WFFu5gSbslrve+cM3g/XV/e+IzreYb6z
LhOQrvrAq82Mhyl+Z6OCqU0icAETCXIswRfAL6kv+icE3OkAY9OSaFpi8V+r8pUV
GmCab0pb/8UZHqYrcUjqRbpfS8sWH98OV7FLv3zGf0SA2RLzfs/RjDJSnRH3YZOs
y9ln0LFJp3s8QITdcG21Gxrq+QFqSX+re4axvGSexzdGEhKkZxlDWUy2tT0QeNeN
NPzVMJZTmGDEVIV0zCq3grETRG8aqtxRiZ/lGEhOFDCrJuKNIT30C4EGp+5xpWLb
qi3aggNfc/SjecS/FS7KgfJo20+Y3fbg7D5wOOOd0XqsULNpvy7Xd22zeUz/TmTY
XhAfeSoTEvmu3bDV872LgOIjaAMDlM+uCPIq1YjGcGxFp5xC1avdAUD31TdKyd1+
1NbxO9IPEIUGeCdyYMiryYOb6Db9QQfROvzhdz7Fe5HgLpEgfKPJsjx0fwbBDHXv
JSHt37xSxLzsaAKggjOqxy4Hc/aknwunLjxWMuZv/JaC4ysAKNBoiCaqozwN3Zt/
HuDy+B7Q8ellpWNhVc7t8rLwIwvqFsvuqZZ8JRoB6oC4DTMaddNms5O4xG7Au2EC
LUZMQlonK4VgKNuA+Znnh/FffHVojSBGZSq2QtxnpiGFNu8voBIgmvawWzrjR2sp
yGwdyah8NZHwfTbiVUa/rQ==
`protect END_PROTECTED
