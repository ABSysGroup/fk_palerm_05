`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WgHIVnF1ysI1MthGPlac0Y2hQAE2iOMxNw+e2F2V5dEnXBPzqqBtS0yDbzO8LPTg
ckpcGiWZA/11M5MFiwg1Kl5KNtjxZ90j4Z+Sclwr35RJ/0HiMqQjr1Mb8oVcA2nj
Enp0IdUmL7kmzNnkT2giiT4IwOpMvOBqQOXOFqE4smEa5Um+qNSDrO9/9GR4MzFL
r0XYHsR+gubI8bSrorTuU8ElzOyHhWhzXA2DF8IrFOhT3g6N+RH66/BeFVcixINc
scomz39OqNQbKeq9Wi78J+5iJ/ZmGiEqK+BjGgIjgA8RMaoIhP14ad6mZxYoqjZ7
GiLI9xc8AaBXo9Ncq6q9KrdsgBGieoBy750BYqr6bp11zBYAxATAsmiE0aYeXH5V
EMem7XKyUOVWl0smou/h9abU0py0RNKIB94hR7X1J4zb0JMqm9kp4EKElHKPbf+e
ZKGMbaVBERYdxtcVPPGS/yAbf4AUSZ8r8n3pat7o6qs10w0dZ96a/FtFSGF715Tc
gjWBjO39mUArzbunn2WGodoJZhLxxODQ6c42L5tbTeW3LJ3uE7zWQt+34TTQZZtb
Ki82wmhXgHrU2Gz52qF4xKrStkDDw2/ehquynPUwKxZUMe8DKxPH7dGl8u4wLj1k
l2nJ5EXsyyFCU8khjtQjfbZpMFWh/VCX0baOVPFs0us6iBeOwrO1Mq2H3IVmG92k
/oVYBBh7xxYdp8B6DjQfHzSvJ5XwXuSzaibminV10BZ97s7euK+A1pkO01v1Dfr6
tqSS/ivFv5aogpcf2hvAWTqbuY3PktMGHXB2w/jd5ZszM3nzakY4YdTbkXA2lKXa
IPBCSH5ExxCChhgO5JhGhKfBfi3iFWtBSXCYENsPjHxqBvdWmm+PlVysJfOTErG5
Ov9cQFYf9tkVKcz9/gZYttDfVSS617BxjjGnG86LrKfxmXO+ayc+xvyKtMhIBbC0
7mo+sPWym9/XdlLmpBwM7CHLruzINUaXuKS9DtXMbc2JyzDrRiQdkxhnjY/KplZ5
i88wdwIqvNqqs57w0JxPXjm2kXmrdLdOaN/pha67HBG3XFVVLakXrEQy6cvx5uRM
ZfEb1MgkpdmgFlyl1qJG4Bj8MUHDdB2icV6stRfuW20DFaFHHcVuscEKHI5LUvjW
Lse6yJu0HHiWetvhKjB05ZrgpnY6+uRYlHQr2vJLhXhL+MqiLj7W62m+qOkeyXlt
PuM5JF9wR0s/3UbVYT3blwyhABDP4c36QC5dDvfudMNBab1V4fQK05qXAb8a3elc
f5uvazy4cT15ysjwPjFR61ua3dgZ/7OeNTs0cUuvbo8RPGBwI7NhSrMRDvvyFTeT
44fXKIxiEaI++1sqaogQBOSoqbuylavmb4y2HiMln67pNqGwNlguy+ZBniJld4Ho
mgUVcopP4GWPYrBb8CJKCYgq2oSYwBr1xJYZ6m2+Hl02QH3IusvgmEjdOXg3GS/b
P5H18Y9VzKacZS7uLwB5yx12Knc1UbYvu8CYYBSNoLYri8jPEaGwXK7QztEBuIhe
sKCf7LArDZ4vwx3jHr6d5tjOET/g4A25BV1YcsNvMN6ModbOZkNtGv5pTxhKqNiR
ZxAe2JtivS9L0183JLLVjQTTMHEYP75Fcd3yIXLzC0CNIP38jdzseSGToThBbnrT
Ozqbc5YKlQOoUt9amRLAV5MMK/5FKpOhXcjPpcTRg6mNbaaH+Q6OzHVKUT1eFAL6
n+9QvUXruP/niiTp7r8Ab9akg/p2hVqr+SQMzI7NDD2npHqKoGKKBwGigpoazBbl
uuCaspYQGzpLwVmYh38zIhY3qE03N1LM/GTHK2bjSdYCpsBYgeUfzOKVpY+h6sN/
dr+TC2NveJVhj0tV+nTTdEWEDeQv5h7Bwo9HlvmnAc/94DjpZG8jz/VPQ0iajdDB
RQe/eGCd5zQ5+iwNaKyvYIy8fP197QAouGH9aG83ipLnUFW/mJTmLrje/DiY5Ie3
nCPFK36Jt3wh9x/mA4UoKEtyHdSby76h0BCnwzwvp5bHgks2HtGmAUYdz589yOYl
uIAR4I8shYTKPuq3Nu3hVKhHAUJNg3kErTdtw+RSKu2oeq6tKLSYU8DJpRKM7lrE
g0wM4aLeT06sd4Y6fzUaWLlz/9OEyHNhGkH9Z+tTa3eEk1s9o3yBhiZt6yXqSF34
uCkwQO3T0ZUrZcJuedkX8LtUAdhbhdCeR8/8WhvP+VSGc8J07sy2ABfyk4broqjx
//g2cQIL7FmFsv/wpOO5u2TuLzjHvMk22g+pxlXDHxnPciENLJChvhhtq3fc0JPA
i01/qg4kyHOi1U9pspyJG0Q3HA9V8otvL3ZNLIGR/2NlO7vFEvBSTpjeYwh8bZMB
K7fyuB+24UwCuOdyXINFIZEBkPOWOuMnkiT90QOrkTY/jC7YHGnqQaJ0BiHb9DtI
O/oFRq92M/kgMSBRebeR2BVHZTqVkDovWRE9IJcyKbBU4aj+K93nDgk5/2J3nTCR
Nzi+FpQ610/etFjbrWeExM1oorV5LzbUCXf6jSYlZ7LOZS/U7hSw11INrWvNzo6W
xJsyCPvJLybo+Dw45OREOmuMhYo9V/uFeet/8bSyybIBSoI8aqShX0r0MLtxQUVX
EQXqNoLmxJXj0lUl3RQ4rCDq6cwu5fmw4KXZhytswobIFxvdCgMUuH9N4fxpzz4z
3TqDBQ8MzkyObat8i13zwAya68385j6Vs69EBZg1SDFNg3qkE7UdJBSmrCipF4I0
5OPqnEUHxojGk5qrdIV+FwmY/8dxd2YgADJMjeCGwXvSlvQIlaaB6EU6Y6wlPl1b
dpbaHh9axaKhta8IiDr62TQoJLHaO7IPW9qM6LJYRwXySz70NNupmcH2/mAtVKt5
G2XXQaQfqFgsRGmMixarlLpcOByCdLrXcAWMe7uPEfLb2PfPhWIT11mQpRMklJlJ
KmCmzjEiqenfDeq1Ndym3ihIUoLpSuOUmD9mnR45lfI0p3U9rDBJJUOkFKIHci+E
lQI30ZfHFqkrOBMdFsbHzFz+4W04mcLQCD8wsJpltsKMl4dgxCbPPl7PhyNEI+tp
1SQEDxkGK9+bT4e/Bs8FlBBAj2pup/naHCBldTVZWHE0XzPjEKEiIs+44gXHp+fz
fqdLQQ6m2ydysh1Yg8S00ySp7KV7L8q5JINoQHwOBfSsbdjHF9xMiD+pVAz+avBG
KKLEGFkzywcK83JCNyyFHDAeTIzlBeQElnjwFMkQjN/CHJdvJVszkTB44fQfRacJ
usgcn/lvY0X0UaVvAygaslQcMC5qE5yNSd/W7AS/lIZ3qNFKOVCegOsNbFrCWLZ7
GBI6HN1P0A3l4FTwzD34K7TW2rFNQg6I4+chvIZbidFvp78afPzDdoUwgeltdYeM
85X9c6gWMrnSgls0MI/qbyCIelj3tryD1CHS1/xzVHsnKfb8q7UhUJiSroGGXDBu
+/xOtFrW5IrKuIHVaFkevPFa6QFoIuAAcZoAY4++8GJxsWhfTKB7COiIDc0lFrSj
p9umz64YUG3dwnoR1IHUgeGcsuacIBvgQ7sSzqIFP0xjJYS8QNvu4nE3UVZzOVmC
gGNklJiBXW5/4tz6nou8qw8DcoT8mU5dNmG4W3CXM40aT5eFA3R1/F6OjzSe1IaI
neyYtfdSaQpewMh8QoW4UGb2mG07K60L1R8nW3BKWQdjqzy4pKcuhFnvhZL2QjOu
q+ibtxfjvRUNwL9o6J1B8ozhwuBmbPuHMhXRi8TbDfYkXfocdnBC709WRY+Sh8L1
dsgxtly/NynFYlqeo/y8sao/Um/ywYA2G8d9J1dQ+e1K1u0e4MuVidLPvDxRoGlL
E9YW4T2X/GqlmcvsiAGtQ+GsmuyfJ+FIB2XQm61cWPO8dkcRpdd0R4WcbzVTkrJ8
60XmdBN4TJz8adKw0/t2z+frpMbc+w0us0W0Saavgq5ijKPOl9bzBIlaxx2SBD+g
qnbI9cqOkZMwGEuj4xVPQQ1jvFcAif+41WGu0qvmuPgS2GNCH8H0JMORU5khgYgk
NgeaNJB6zQLLwpA1ySenkAN6+J0394pYgcZ8U+aQ36dFOgQcNLA/fxPjvmokwfrj
Hrt2/0OCfhBB1vSVmqq1V0M6Pr090VYvHh4WxNwNV8G+SvWqVSVHcK9Q10DZyYb4
v5tZ825tCmA3qVZP1+48Iy45OScVba3nZ/AbV7or+2hjsaasesgE74xj1YKachOQ
ydPtmSs971O/x2Gi/Q/9Epo3e6OkvuTe7RMb489ZtA5idRt6sqCL4QAsQBJp8ZiZ
5qx+3XTQhZm7DmgmFWJ0VWeGdqmo9324yBfakMikxH8BG1mcD2agDhkfPKqQ7iio
cr+7S/sSeNkD7X31koGJTDsKOH24O7w9xvPsSCV+NdrkZEYAj/9ROpu2DIx2X7+r
6BnlU3AVCV5vUHUCMSsagwtFfrNLk88l4q8s2hCao7tNxIaxW1QeEB19DtOYGucW
vblXKofFdAGB0RVzH3/SAgusW7wk0UqUBLKtH6mAQYguoO1bkhkTyuHacS6JXbCG
4Gj1EvYi84WOIs56m1D51LeFrwX3sGRrfl3k3R3fk8DO3g6wKBIUqNDxQ/hpeXxZ
nKlYR0zGBjMQMI2+vjZs6DeW/ZWf3CPW/1cdHMm+sVf4A1KA71X/gtD04bOdyqVP
DiyJA9BQI3XdT30+hMpsIm29mn9tw+djb/tTOZviZAHXYiMxalpfSY9ZyiyhWOVZ
E52ukIuHEi1zrrNC7ZDcVEQwdQDiOoQdKz5kChhc5jzqcgQFEFOThnvJPv1/veTv
40mYIZCdxfs9j3hAfqq1hpctIKyGbY6og4isjczfBJYCtwrW3TAvC0sB10SzdrsF
iU4kR+3474JxPYclKEDAl5f4hvmrHmKf438TZ6ibUDSnrNWPF1HYEHtFJEqs7vQx
LX+L+vzcFELxg1zAJZ7UF6q3KBjiYEG/vLabRUxKjAfq07i/1kfBDUZw5kpy3Zxu
FGyj1pHv8ZYgcgaqHMXvHkgFPIti9cnB+mXJUQhQotnj3uRYn55yeFvPvuEzrHJI
IRohezr24zEW9ezBqQQfnz91e6h3XuYoj44VA7lZvdDBID39DIgI8sU5CzHZxRB0
w2vsLTXjnMrYlj3uvjitHthbf4CvanutsF1RTzl6D6EOtzqXE5Ge2QYZO330FjYT
spkIwVh6iBT6Wa4chgHio2Ig4iLpFoybrTnO7vt3zIBksKenHSqXAofSFkHGmohU
05IVdxIvLtUDn6q2XP2dr/DmY8HNS72n5nntW+J1BwE4WWTZI0XWp/3UvMDxQkas
uNOnSBgeBN7AHSs1di9AntvaZNmd2NKxreVdYjfbPXhHBBvR2KXOdhn50dCD5f3F
F1mA6eixsp0kLGXkZetJ7WejVAfY5ilKzxvU6/Lbg5Vg0+8eGr62D9LdyzLypL/h
lX0Qnh5aPmPGz7NNcJ8a1rIAaeHbdAX1b1PJB1TMdELBvdWgpEbnugz3d/k575XP
JMIP2+yvup2BGPRcAoiDCYtrvxznR6huWyMSikurTF+1O0FiIE6Q+H6MEcETismf
UrmSnb/uAxBwcI0OlfDHTg2JeS4wxXNch7cRPLI/65Q2pAWfNPRdbwC1mqXwv+Hy
DC/epP7/d7pyOkA2xfrexq4P8kJt/Oa99ctO9uq1i5IaVAPjWKdFsAvuoEtkX6qA
MPzUS+zgw90D5dkCkI/sQYLNLKbBU7SdeilVXexe4p9V1NOhZojOXJZO0UENWBm6
J2buloCVOHwehs0rgzMC+K/NXaLh+GEecXy864N6Q/higYTMhqD4W81OiitMIRxO
BQVfUyAPH20uXwriU5SFg4m2nAiBe9fG6KixAYPi9bnVWrxmtBOxw173PuKKk5p1
WrCjPBb05RN9jofXMKwtDvaAl9GqDD18XPuNpcbGCLqXbEoYubdfNoddJFKF1pbV
olI1agXkCQ58RRcbAOI72KTgGnnOEm9Oos4lamAELmWo1EOnosClJ1iSG3S/D6KY
4HGSYKsuZ1fO5T2HZJ9ijnzE8jb/iwzpJhpJ6PUf4ZEsPgmjHj1EGC2x7PTxzlbF
m2ImlRIOJlJ0VbivzgT80l4dH1raEHG0TdzOwMxnynKiW5orGpD1VrLOx1TsOoS6
a07MyZEZxDiWat+07wz4VCZu663s5qihvcn6SWlMUY1YQgsTlOMOFBatAqorzduf
/JzpOBDhra+3MrwbNpy3xYxl3Gs6Hlk2hdbHAclGy0cV9Cj6W7lR/pbo+bzweLkl
YUyNzGwu1BoIBChWu0x0GVSN5NL89z1j2z+DtHxbewNIyW/ULNhGHGnLWAzgxITM
KoDwum4lJ1LrmO50UijtY+L5EJwsSXrSzNOS0OWOCjZheg3ZTxm0RSQClQdxe5DR
7q3SvV2g/4b2pNMBGOOknXo5NoT0+1H7VetNhXkqDaWyyugsv7RQznyNenfTVS57
lOLLMj4tFt58RP7fNUC8bwZDL8kX6wf/O5FPB0k1FQb+czFJ/iHUObKN6+7C8hIb
Z+igJY2JdZNlhZOd9pEcUNWnHCdQXSEHG+MQc3E2fSF9a6MWQJIpJjKIgOXUu+UV
vdY/bVp21wQFEU8RsdlF/l1yFQlwhfKZyYF+1aUkkZEAuUpxrcY6eXyLe0DIEvSR
GIsd3es9eR/ekjGJmOAE4YrUErbyoJpioLOWgVUqe7krO5W2T75TjN5tR+ZbhYaR
HPOA1V7HvocAoqLFVO82KZm1pF3ncnF9XCqvejolt2ehDW8mDsN25e4S43VgEZ6Y
gFiWbW5okctdSvNgros5pM+Qm1cc2VuXRxlQmd1gPQmnEjlOp+SLZAacPGnvT+0c
ecTFNDmP2g3JLiDBCyoJY6vzrIE1HUK0Vop2boxNdzNbpoQ5dARldYdvsa2QsBds
u3w6aNzs6i02yztDdFPKNvY5IkvnQpE8x3cYBhcFX2P0igiikTawAAvhIoA0bIj/
YZgEOsNP+Fyyhl1y/m7hxTgDTHtwsESc5ELuN07YxttFBRvnPu0r6POzUrg153+J
z1h3jqyHDWUQoL0YzCQOZ8sHLHyc++kxGy70TZpUqPZBFtJAYBGGlIx/PdPifd+f
iDUKHcKlyyJoy6RQNZlbuwYRip/I5CqT5yl5RJgzmvRC5JQUdK83kMjXe9Zsw5kf
0BxJB1HQJe1GzU82oRBa3xJDUUBI358pN3CBZih0bpB15G3/wja7HMCLYVAZSwlr
pJzjIOHjvedFdo905V/7DHVo/3Ug6CYyWD1BgCr78U8QQlZV7gGojEgHxkiABNo2
g4S7Rc/uApaPIE8fU8T0Eauy6lp+stvrw7Dz7NzWK2vW5g7TwTMzsAgu9I4+64gB
6VAr8pWs26EFeK8iBleINRebKI0pOw+DNVUtHZOmbkfiPOFh+yzd8LgeFVDzM4Y+
0KKs2TYOu2cLNmGIQF2+jaycr4XgJ4SyKEsFLB8Q4X99nJ36bchXV6SN4jcp+jQo
hkb/LjMayzZaep+wN7mH9fPR7cK6zrA7TfIFKsMvOcGGsl5WFQz8i6q2b5yfDaUi
KsQkgnMfq+k3pFIGIFQOT0xIGT8kpgEFpN3dQtGZhYQQKfgW0RUSBi0egqTFuZiH
dbsPQ6Vy8zcPR3mFEqhD5sAbfpbsWfGpKT+Jcm1x0lx6Ka7MoN2VxapZ2c8qB763
gpEeIcPLNn/NN0aAtML/7udRUn9INfLXnCWzZrfkqGbhb2tdLF52AMJ2rcE5MoU5
5kQ15Jw/ffV3jK3/7Cdhh1Ndq7/ggb+1OtHv393bceA3CM5oI4pJDj7Wp2K4mdLi
sldUTaHoJqq3JbMmFQYdxCiqcqL3QjdxxXdynkaM0b5n2p/Ub29PRezDZfQ4QobQ
MBGbnukMEDD0/YhFJPB+BcA8/40vX3DiEo6bwUmUnffFDKejQj7RLcjSiTBiL8TA
l/Jd5lT0rWtNfANpFIOQL7AKwy/zd3NBMHGvqkiH/SNtzHUzOVHlzgxa4BYsNRav
L6LXB1T6sdP1DMKHxil6eR/gL7s2qcaxjJflPeu7uR8XP27L3P9wNLuHAwnDbhcI
ZNwFL5Tiz/mFhNYv9AC+7REG3YQWltHcfA0J7KJb66G6Zv7aVVrnDPmMTEYWimjM
QLcpp3+FKPVXUVBkyzshEudy28amGngk/SA6O9eCvLHDM8qd21BBa5p4dJpMJNUs
Okz7LSupuuL9zx0fBLN/m7xCmdRdFgNS25QTurIcVb88i8L+CSnpx+YIrKRwPUH0
7lljM0C0GmHdHZ/a5ijJL12Ip4ULJRi2TdYjoF2kgN/tcqW5rg3Q1FH8P2tNfGwU
FGariMr0c7gRd4eZiIKIcQj2QbaChzvjf8Ub50U1XR1F4CRFDO4gSYvbAOFCWb6q
ZMwDT4DWrMfA4KF7NPzwcUZbww2tWbSydAskpXk2BkiV2yj17vldWQSh+/HxQk74
0RsDLUmmaOVn5Cg8+LyBoVH7sBvY+1TtscKlZNtdVOZzl5RizvErnoCGENVybSVu
CIR9a8onGEAsRetRwBAoRkTmjWRwyHUJV7c2q8Pge2UdSMMnxt0YBfN0fQ1fkCqR
34Np9St5sfzJpGpP9P7xEoESySChrfZhmT7373poV6aDAFbKRaBgFdiGjgUyJkYt
bZRVMjyBOQlIxyfc46lCeuK2nNm9fTUErhfE/trAE75xuq2SLZMregd5SZkU/I07
ajKbIfAD+lW0Mcxn0OmoVIQEM1B+Ff4OoQIftLMw7Lc8TDq1fW/2UUG8WVzmXcUL
VbAk/s/P91dN8z3DDF7sLizStwbjlNZ8CITP8LH184DvtdIYVMB33Pk+VdQPiPCX
S9lXi/qf2UGphRTpnLhHalrTAEX5UsNG2beeCxArv25HTFMvADP8lBonHiLQaWya
nmucFk4EoQ8kGNdYJK09h1trv+lJjh6VLbg7AYfKIQVL/rMbMpOka7ljDDKVnxS2
lzIEMSCUoV4tvdyMgi6x+BgOrTpuwhKDIfQ4ImleDkipUDCN3G53ZhJlK6TxjJnr
IrgrmiSjVKN6ZA8NUF9xDue14PgTb4aMLlgYQWCswU9TyvdeimVzLhpVIf9z0tDu
3gfwua1zhvhRu3UOr9KgF5mbZKkijOzBeS2c0BfCQJuzuagxJCmfF7eWWu7PaZsJ
ObF0ANaiecUyB5ZmZOiFDsly7PwQpD9r8JdckmFIVkX794VBL9RV0vVd5mysoykX
1BT+zwr6E+XVTibwoUolJP1cXMqm17uOBmcg+qYlzEf0qcVmfKARjhYDEFUc3esa
ND+TFDRXSIPX50Z8nuSc4K4qVMP5MXeBzRk7s3UYokJl9/ihiaKuHuvT7oiljOuZ
E+uV3ka3Q7iGvCV+cUZ0TMXwYZGSiHcVDWO+GKNnc9GLnbcKeGDlNysSVnVnjbSk
bgI3yh3w9Laa6XBrNXHzNFL72HkNtGqsK7LvZrHdPu9FvgzZe5ZDLm1OSb6/5Lma
pA3k2qVrLK4DQ9u5bASy/9PnA0nJo1FOuzrf/0qtnVnVHLZQw7/jZTss+SbbDww5
OSZcJf6u2cT1AMSWCF9l0WiLy6nget/zRsR9ynNfNTMudl3XHOTwHCYQB71sCQPm
exxzaGU93clfN6CoZie/FyY53xFvVB6UhKuFc22sO2wKPSU+TwZCMT5/1JCUfRRo
1VlHqK9PJ/c2L0amw0FAC4QNQ+mE+32YsXWoXdFy4V2MejtFEWNJNHGxpMk8epc9
M9yrzqeflmbvqXlVIXG5nIHwVgWOq/1bdD/BHAxFtJ7gCaLwP7XRkbLhaH36iXCK
OmqZjo6OlBFq3nHItG9kjtK8SWvRM7Fp3pRYgPpTWyXc6R9SYRuU7/meueLtwiKJ
uEu5isTfucrMEFC01L7wPjqKSOPNMNxYA756tDiOHY5XCxXl9iFN4TQ9gO9hOlGS
Dknitvu5/b1v0yPNZ9TModCn8iGE8EUZrLFaJ/sV4L7JqP2Tv3iab6uDCRoaM0jE
xlVL2PpYqKvCoXy3Lih53YDOZDpIfB1+yMj0ulXdHT2bTrK6Fg0ezDEIzJslF5ri
jvqNVwlTP6YWc58VGZWYVgKFPzGq57gdKV3N1fN/1MPipbVSHHeed/Gr8OiY6Tqb
Gx6JuK5HA+Y+AHbzii4i2yLSWyU/0v6wjPofaEiX6FqbkAmTebPOTkQ/LT+ZxRLJ
4vJUbCikAdCKEXyeXMHyVkzHk/mL5Vm1v/ajZ5LHVxjryssd7ooVroAySPGvG+Wu
E/KoB8k0IfzF4mGeF1DjHNfP06nR5xcdcS5hfZ4alyLYXxHLAGznKF/2Y20UfXea
SoDLwW6iHanSrb3xxxu9Xjp0+74zxgi9Q03KwOb5UbN2Vsb0I9k4x4WMxCYFgBMP
u3+/KhOcTmLyWch1GRSUssBZss7mTQWCVA3pWQuvAqgozX+gomkDQLw7oO6yDsVk
wjusZwayFL6Hsa7We2sFr+y54W8vk5q7DRfG4JFYuB8G9sudYjoSGBBfYmUnQaMX
ckYE2dHQ1KZydDjgnx660zSYA3QJ2KaFvQsuHBoFcQGzvE+niPycSv8XYo37ChJ6
b82jxixVetVPpzcrFGS/dIlVaGk7J9n4kR7KehYq41GnXGDEuVeljnUVTU7iwixn
kTpqf5rEaJXDTw2XGPX67ucRyJiFPYbdW3kcvZIoQhGWuhR1JlGuQcCs33eGc2KN
X+ollUN4GqF3OCsrxqkhFYjh73GqHWccjpZNLoVoy7yrw/P8H3SFmK5awd/O36D/
jYjZ/BnRb9bZBBvp5vtTaKaP4HPFkz6HLih4/JW6WWt7ZNO8d5YhxJGuGBnuGfRN
Ni3/W8qXa367R/5HbRxUurVDcJ2Ab+AGjE0n8EhkPAUyzuCdW25QChhCU3PcF9m+
3SAlhKfmwIpQ9V/a4ZMXZqjBdhECathz/RPtt9TbeuT6fsNxjcuI5yuenUfLLVEa
uBOFLmjzJ8WONhwIDz60aw2c1sabIywsOsiRa7nBuBkbItw+Nb17lPgb+RavBl33
991tilBV7oR4FgF2O49MUJzD+/HCuZrenEm0iZIWjuXyzVKCRnvO3PyG9R4SZtDO
rIilHaYm8F+pqkiBuNynMsAS00CAwd3N0a6PLnB5fJX58rvfJlKmUOrKBrsSC5oZ
fJxIuTg3Idhmb7oPB31kRULus0ZCpVJJG2ovY0ZtYtiRsySnUC+T6PiXTHU4utzn
TQk+9QCdViE1AIYUYU92GeAy3dZqebCfYYwYArU1CrICNY+bcWCzOppnWN/uEIrZ
0z0N55WZwtCBwlaWErT4gh7sn43L3JY7OoHpnE+lxfoSVr3B0y/lxa4JBI/ks30E
4pBLVI94NfuVg6FaAv+zuLrFYASAlEJKvFkaf+P7cw6UFt48r4jKR9zv8dE4FEs8
KI5rUmM0dmx0YjP3MPzl5iVS8Ixjvksv6wv271T3JQEMq89PP+/Q2gePIfVA7oXI
0pc62a8fGYlk5zoitWisD8gU7UUA2DdBlduJSEFqPiNYUZ8/5hLP1i3U7tv3kruk
hc8IrXLfoSt292//JSEQc08j9F3RUNn0mPa6IRnzR0X4Hk6nJlE5fu0wwKRK8lR1
qnZM5OTKSVy/u5n3tfV5+JYPGTna3YI7OYCAOAwvNfS8V8HeUKLdVYdCD8VDUh1j
bQxox1+CHogyR4s0IKACprzFWHrdE3Aue3Oj2ufsLVQuWQgojQDHyiE8SJOW4KwL
B2L4n7ihfL80S7JIk4v2hH8xcuwvOB6UNO8Aw9FUESRxVPHksDh952Zvcvdxd1t/
JgvQ6Y9sDC0faaorH/dfHYFfwEVNUkUr3PESDNZhnp7p8oz9W5JNL9/VuEE6xwLs
XIY6CNp63tySLiovuh38ykNXaLv8wc9vrlc2IDvm98RjrpyiwtA9UVWb9nVkEIbG
60mltAZFiHSOTEClsLfVAerZWh4sYdAoZEeXOltytMKwcxOiXb/JFfEgAyaltCH2
ulqdXFqXEWazi4VagEwGHA2tGURgbsE0nMx8DQMU/Ctu6xfGKNI7PXHdYl7zXmJM
tvgTVlkZ3Ts8aZGbhvf7rCb1/KgLiOREJtYHbMZJlHxk349fesWICHiO3OoHqdj8
XRk0wy4aVhaZ+MfzCaKDsxO52J8LGMDjOa2Zcx4p7+UHmJ/N7j8jCcKceM4LKEzd
Un1V5AqxQrP56UJGC3nLxRYuKlMkktJvkLKaw+Tn6A5w7fuI8s5hxeI7uilktZvc
aW5hUSdwVpk2/RfS+SYadr00ZtmCT3z1QKte6kwd4ixBgI2g+92JhcAwyPMLGt6v
bsNpucsZP6GBotVQzqqoZmF/ru+bgjLZ9x2NTKN0HuswYIk6Xi9pbyIThZRiGYlL
WSWhEghZYVqTee0FLE+91jRxOS/ImJCOj2lf10MeGuLFxiGiiIRRskwq8L6YLZIC
eTqdAKO8EH6HFdS9QnkqkW1y824waC/oVYKvPusFr3OsT8l3JXs0Z+OgOT/V6du6
Zl0XtG0Zi59PZ8gaCpJ2I3LZu/ZuL/QiJE/okeQbvC5+6TtcvuTd2+BBHGEOwFi4
BU9CyOanO53pNsbg06O5eM7w67qoIbto6DpbzQHWCLhTcuIjHskj/difLlMemU8q
wZOgvXZxHqteijblHKvSuyUNi/aJiracvWkDkyRjwADid1LgoR/36gki/GRexxUv
9QwiFOw9409Pe0VvCzFwAVWbC9+mKYGZV1ZEoSVv6pabE0ZHodu60wd0Dl2iwjn/
y8fuBD/fYa+uGhE4tlAqbfMiWS4msk6AAvgN4JOrEp2Sh66wRpbvqgrBFYDYlpYa
TZSnZZ6OshOPx9VjOnVq9OCFdY/WL4gZnHwTkUiQL60rcirzVLGAnozviyA2YoO0
rsmGeSz6O/gYqEuIM3m4/wA61QAHY8rJ+fJqTZGaU/vQVWoUtOxix15vty9ahCLx
izOeFQmACOVn5XJRol4DLxNJ6vd/PSW+cME11DbYoHBcKMCcG+m7KWwfU6BSDwV4
3HvN3u+t6wcWCtJYfQfuIyydIjTOuVc9WYqkk8GMS/KQIWqEhIzslwG8fKlguDNJ
DpbAiuUjODFakZvq1/us+RbvMDSbwjaL/suoklDpKtqtOZ4ac9zd356mJFcania9
fh+XSnwcFpIWtf6qMkMceKpRZJR3BdsgBlOweXujl+CKdmsAnG5ncPG5CzieelQe
DHUjIytFTrm5AoIbSH0pMJ3OVN9mHwVF7vPJouoS2GuXgNPCmbDFdI4aSMuxEeE/
lYWdqJ5jsdzneRDI7zfcM+SdGKWqwQcb6O44HcbCAnOjvnHhD+9T1iKjs09Oiqv+
i0+XYnz9WwgxjGCTWL8ow/Za5G5teAHmO5GG/+9Mb8UWO1HI/oEZV/3xrOLzVgko
SJK2SkHt/GhQKwI3ODkU2RNZ2AqfN5U45HHyCnhz8fXyQHzbJgv0KjC1trJWIk3m
vmkKLu6AubixgzPzrozEIYuym3AfBqipYjmnGTdsDB+CCWlViagNGStB/kExLC56
lGcoLEyES+4/QUknkWNtCOlk8bt8eSDPlD1A501K6Gz2n4wvcsM8WDOfZIOrynjB
wdShpaXR3fGIOJ+wRrcMI0UF29ujjynMGGOVEjmK03Jy86y8e+NQQxC+gkoIT4ho
oNpwWX/M2ITN/LSRcMegrqTlZpfaeRLKYSH6UCr6OEujxdK9E6k201ILinqlOz+r
6tC1Jy3lsGF88MdmFFtz9ifMWLelnZdmShw0oDseCC9CdC25yb7dKfDTFmkUSmKL
nzYq8+syJHfJp3hncWRwWL3npxHcYYRhz9zuqACn6gmHC9yC4eRvV0dqrs6f4kau
2TlKs18Md8YE7dAp8iNyXXqDJBtTOlqQAUNgs4PPmbjB0H/JwoXHuz7u+1g9J4ub
Ut+egdZbrOz5ieKrMBqGtf9skV9GJzRqLVC8qMM7/zfb22pgloo7BPyu8ekDoLLO
zF71oJ/1cmQOgC808dq7WO3KQnHYq24WMtKaaUmJqYnk8khpWrukPUKfPeB/3TJl
75idS6+dWdqXsPQvm9a/zCTzdGuBdcdizFw1rONA4vy1SDL7C9NdTOA1R66yvNv8
MGiVv4+bSOZeipUONkGmwTrWrA5DPYFL0j1IvM0jnRnN0uxhuWZolJ+4ZUd9Oz1w
TQecyxAP/YP8OzGhdUmZ1twtc9dP2CzIqDLn6oI5BGjoJTrKKNxBWdIK3bJtdiCN
oIWqp3Ot4eA8ExPrqD8Wse10Aj3P3gcOo17xKG4hdUb8TgeHsIvVwDCxrxiXkzCd
1JYFTqbMyDq9cTOYnGXTABjjdEM/6NNN/udcXmbKk96Nmkiz30UurgPYv9CuCUhg
djoUqxIvFGJ05m9pOiJwMljdrN0f0F063auimuHzzbfrnM9qv0pJ3Tj/P+0Uo8cY
AiCU5wwJOvXmqx0+Nu28kLfgddrx+6GaBdf1IBJHMoi+M4pdYMTxc6e2IYl8P4XC
bj6Iygf3+e5vIN8ZRKY8PPN60Jp7NgVUt0Sx+R2betNgSNMliV8+MIH752fPCyjT
JezevfTtcY3U6kAcVERF32BI0QLIVEYGmsVp0jXEj731lGEu07w553THEf93IrHW
vLDoGIochmYPa/GScLwdQutweqTOC/1IA8VPraPJMIr2aLJJkIpvh8Y10LZ11XID
tBtSQUAZtQuzZJqFhHjFYHJwwo6OSeGv1Bj7wjdDYeUQqEPhdpTrg1wJw93m981l
S1lXMGm2cS0cLXS6n8VF4c0X5kZTGzXR4qpINGdxD7U7tmJdKaMSCMrNTu1zfr22
EveepZvHkW9FkR1cz1K1btLFJ3VyK7uGQYtD+PrnmAY4FUXOyo5txHVEAn6hzrdb
HxqtcPOh2hzGYTOK4KF2OrfoUgGObTxEfETvclHUWf2zlwasfHY7/VJhBnGY27mL
pZ42XA00pP6lpbUWybAjQRaPiP3tCQvnDH8Sevbtg22y/s+0t/7BJiTLQKQn93xv
xm7+O2rF8uiTeePy7Cnfw6YrkcdEUN06UVOOzqexKK7b2Nn4OlPIqQyXA8nQQlqS
NSk51VnPSvjOWJA9FsyQSnC0Odn2/q0VAvue0SXzJx3At9WEx/FU9yl4FiDofA7Y
0+z5oVlXlUMHKcd1FDD0Nt0uceElS6XoxklzunmflFWQznyzEcNSWCZdNWoocL/+
NluVEUZL1vamu1KUdU3wMcc2FLHVkAzsRnNPJ4JTwahAsiRe3BGnQ14eNa41qjso
9/bPgEwmByJERnv+PbgIo3YChKE4XizO3uWYhOyWVoEX9vCoprav7xHVPLjpD1Q3
WuLFVrwG5waPsFWNxiYFRWb9GvCuQsfMs67zLbPPJOpqkZIfNoE11K19tj1RL3cY
dbxS5qfQaXiadhCzZgJHOldcdlRFcaTGzwm0+/5JrhU6B2mkQqJXABZ6+6DxIa3E
TONja69CbTXktSkAO/jQiHIAL1+0N6dubWH3czJyssW4cBY3RswNB0B8/JYCdWam
GSjW1z4UVMSq4ICNxRbhVuMjSTD4psx7+T+R2pd6XSPpq5ao+Nx8x63vEdGZs00h
3kA+ouU5cM4+XUNVeoU4A0BSlsNAaeTtgdjfC5qoT/LDt6g8IvjyHhC/5y2y7H2N
tLObPVj0t5mU65aaijrz2LJdhsQbt7AdtK4rRh7yksD6p3GSylAWmuPh21Pn1YU1
PSDJyMyRPhZr7Qe7GiTZ3PVx0BRsNafkc/w1b3CPLXI1GxN7Zn27erDK22vcJOWP
kmstxNgrNNy3KISzofJBdNoqdY3wVXf20Ia6TN7VMvZQJpEtPNCEE13D4IyKJIHa
VCiPSwBy9U5CulMdfJQdh2CUaheAfYlXbfVafvdY1nmiQhGs97ij9L/5/zdUc+/W
cUomPKNPaqN/L2cF48oUKKJk94f0V0SPJEd5RX51EK9esiNWbrbkUX2GUe1vY0J/
7Pbxut+iLtrN5J1xzPLjdRggyQujGp+qT7Om/VdBwwdmLDRbh/f1qtVqZ76IsAUX
ULGLfx3TpzsiZCitFw0CHU0T/CNyt+bQIjTIbKcmu/Z4rK3FYpoKtn3rxg1/H6HE
TNsOgWenq4Nn69+L9VM76FNLIxodJGnqTGy2h/o7K6IvOR83idvzw0ZNQ4No2c/9
ZUh18dxWjqmraCGG+DzytqvgGDo6pxR3AzCSMqa+M7Wu/JW2BNh05TSqzz/aVAo7
zkPzx7frGXb2q2KcgUUon4iGyoDhhER/lbPljJ9NObeZZoUfet+7BDy/9nuphCHl
8cvCdQDiMy25P0yMG+VwV5w8OY46RaI0iGSFn9CqOxhleCtBzAEWbA8DDth/ESeu
T5/QL/F1qED/Rud5EjJThvqR8nCBWhD5jdIJam3EJZJ6dWGMlCLpkAhrQ0zQ7ZSD
aOkSp3ztm5+BUL2LBRQ/RXbT2H9RUV15kjpetcNSZUpagR5EVyzfQlQTjKs32rEq
6hXeDi4f2JpTWCkMMh2Me7vKaei6m5ENRvnplYS7g9oJh/j/hErlitz52MyqiLK5
tQp1lu5GErq9iof9sXFGdQszR8QzQ8ujgZpNuxQbCFPWpgvrnA2D3kcgQ3NyFeiV
KXAZ8alSurOrfTeifIRPiS9eILA+/lUJziXTdImyXmCJM6ZhQPYsDV4PWSG7mhIe
Oriw6FNhen7jMadcsK71TtdIaWiDNVhkFnhthnAYNBXY56jPyBkr/uWsGfI02Wcf
GL7oFcmlmVRoz2MTrzLXmN/zkliYlU9oR8puuc7tUyIcGMC0aEJg1LCsRJ5mjjM2
mkNRqnilp0xaqlhkonWsxqJaxrxoqhNfacjQTD3VNjliecdqhd0nKXXuR0HcmMcU
funkHqrF5cC5cF1DBPiW65EZsfXMjROg6OiZPb7HDlDYDF80sNIbqpMGTs+2WYEM
lIOqvCbB4ieL0y6TuGTgRkEfFR3wOcmuVmo7pNh1rfkgFdtQaHxTQCUpB7o0wewn
GJcdpOQiiRTlj8VxEKUXokj8xpP5gtSsTkxytyKu1/Wft8NQFUCBPp7E9o+CW3wJ
Wpv8eO0X630pfYVDuo08GxTGqR60kvjkQ3w76DeFWvfYnb2mYBNkH5GfMNXCUNFC
LDoKpUImjQPDcyx28NKmBw8y/DxdxxWlB59XwS1lAZWTQR4J2EnotoArkMJVFT5Q
s1fQnZjaOl7bsdrMKK8qlGMXow9bi/uPvhxXT/U64pF11SpWoY3o6BagCCX3YTkS
9YXKLPc8o+/qpvNJJqyLU1LvuuXkFKxAZRkd3s7QGDpjtjA8/T4L2dssdO7o7gSo
1OrKCcgdLiJR2yMbnsz+PTQMLVJwxFBhFY+lgQvkxGSvwj3QvBTmS6SddIj85YtI
iBSeYwkFuAZyhLfxprvR5icJCVHBIJlPLAOnLGZj7V08Xy9oW9g4w9MBEzHWe8Vm
Rh/TlvR3Go9TU/fGiSrMxEkx7xcLHHsEXHTUqqxDXUDR3uya3kBb1c33P3OoXyj7
Wi4jr2EyC/rEB/r3hK7orgQ2bLk/8Hv2GNd/judbsG++gqIe4u0yWDy87L7UFGQ1
iaFNIBlxSnn3VAFqSA8fA+lOvoY4iE/Ov3zTwsITuUaUFrRZ+o1oudgC2VB3R9BW
KF9QhsJs7N4po6Qi7pyTN3K9rBfN4wVRoKxVh81LY5U+yyO/M3K25nYvEHECdWrI
I4fZQsUmwDtpV2Kpc8rGbcOKabVLcdnuqn6hv8mAWwYKbLvE98iuQZO91QW/CsFr
sG1yjms302myl7jccruDkbB2uQhC+MNXscP0n0X0A3FAVBDIMVWLDf5ametGU9eV
iTGbpDiO/f0yrRgpBO4K+dRURdjPcYB02yOhFcbZsCRgI412IFJHSg+Amwv+jHDE
nsdmAQk2ysuiPvJfJ2V7ZBWOQru4ozc5gikg6z3i5gjDI0t5tBSMqECzBZEtC9FW
YAbs3MIgkNdHlqgB0Ys5fjWp9oXz2c5zwokjtk8sFzYUhX8gugcUMHZr7AKufume
YwdtY/AhkHA7ecRJLz/mCIcNo9ozw+jM6qWSxbjoHbakT7aoqpfuG22JZMjqZa+C
Afr03AUV34B3xy0d0JG07SMLq6Z62RyKv1CNbVdlZhooOTvXTxRQV/GB08SQGOtS
cXUgkoI1PdcGPGcF3bzjsomhYVx0Uh1qGKWjPJYJVsm/CK+4WtK25c3bYVuqaW1+
OSRVvX+2JHMzapwpjjtDcWtYnFJyGBgqvR/FSd6or/1VfWL0y7nQ/1aDm2NkTi2U
m5/pxd1pubUz0dCOOx6VJlnI9BAvxOeE5b8ef2nRdAaQiAmZTQSj3NQ7z71sXTfM
Lt83nn7VeqrcAw8fDZzzEtMvUOoHU0DBfgGT3WOklDrDR0W+Kgk4yF+D3itF5L5S
hmxDiezSSxFcgku7KgdqrgthJ5T7d4KOpNspYEbIXxd00HBcr127EvRejdtCzrpC
/e2Ync3Mrbp5DJs8tiXtnh639Tf0J1VuZndR7nW356TUXDNnmhleZi93vtnAZPyK
xXknEqyygREI1Xr8CqiIqiT9MlzDdYeiW7CoAnXdchlE0XlY71wXM9NNDPkMXl4W
sOeOHH/psD95vPApzp+rx0hqxxW1PhMsVdfTRFtLcdQFo5PRdcV9Iygo3+fw2iJh
gF/ta3N9W79DPPdRimjPE2vKe9CXEPdxORGmEOqI/uErXd63BQ71+ELbmu9k3gvv
M+dgSa3z1xMHWr6Hi0Ee2c5u5OtGQESm1aOBhmOy9bDAnxC1TdMRaaJ0iyXPtJDn
V3zeGpk2kwpwnImnfJ16GOv2BJ8kb8orQTn6VKVJUOSlAlXuISp3JU9KEdiw5v5Y
4Wa3dPZ72Q16uVcQiq9pLKAP63j+jmSzTbT2+4dclk9Vl4/20rmQNvsAbzUozDsw
Ai9/sVtEc3GTDYC85WFgMql0WhCGacLeja8LAGVRE5ETEEIo8r1j1dfCMOazc+Wp
qRCQtNOgMDXc7++1DiEhDAfxyTKfxfKz1YMvsAnUAtkbaWPL0p+xyMUqp9ReHRCB
etiQ4XZQg57N0Xp4GLEHZjvJIKc4g9ruBNNCMyWr2Bjf06zxdIn9nwjXRme1bTAb
1PHfifrfES0EEJFbMr2uC2M8P1YkdgxlbWVe0K79zjBQlXxHMshNGijQxhWFnV83
xXZnYhRajI+BNkNhd9eWGPG8t9xCD5dSWO5m4UgGvU7nMDJpY+17rkPMVziL5eF9
/x6s+zTi2+3kk+LrcgCZMZnh2gSSsDuEXWEqqGqLVkvJpbMQ6Kc0cB+1wtU4S4xK
rixv6lCwrgdeCjzXY83y/vkEITJlM5sgUGxzwOs+whYXmJRCwKlirt0CkF7fdg96
Lr+3l8LAs/DF0UqmhLyzz5/F9DHIcrc7PaMNYOzk5Kh9TW6Ht0/J0s04sm3O2Ujh
9iFhUxxiBKl2mVi0Xkw6LDTfG8jWf4qY0MELIXaNWbmt8sMDoVrJ6z6QMV7Nw6/H
pthd03PGuLAHEZGaTxWXa5PPm0Bco0vbrV5QufDyhDFLh6tKDvinMO4pUl2pSvRo
pxFWPH9AN0h3YlCo8h7MyEm/w0KYBC+vzKwtG7oZdxUVpe1C3OYBbnIHhvqIcK7d
7e3FieuwAnbTJEGgBT6XqQORWvht6z6dsPN7LUJW4sMPyFrVRr2deno1WM7Rdco/
hMk/llOtz9sBiM/MJbbMqXplHv4Z7wjVUt6Qas90ZYlgccg33NIZ7FiB2aYTu1tJ
mI15JVaJakDFfqak8tpPJ789Bch280Pp9TeSKWoji03+ZgsYFdpisXEfK4wZQi75
0J8WB23zhHMBPnVjEfjrIcWq6z70tWV6ZRXmdS0GQ+u3E9JcW+mks/R+k2ewuRXy
u6W06nnQhdFQ+XCKSxWyTbws2bhccYnOjw5Qm4kTAkc3SL3mVwEe+F7KzmvOBh0S
5N3f0k64HPFfgpIPR/jrQOKRPlrSDcEVg2wmhxvk2GotoRgB0weA4uvL3k7Pqqlu
VUXgWtLoHIh6BTjbnENw6iYk222+QDSUtody8gS3rqcq31C2rJzvlkIv6O//mBwK
YUFSdKFvfI6dL6PWlomxgZ4sX8A/cM/+j1iGg9WPdc5JbFsvF+DTLJnD2p3AHT/N
EFDc8QgGaEvi/7+q57mBGa0Bx7gu7IDA6ALPOCauoDXn7MwY2iA6Jx+jZkuPoswE
S3VuFpZqyR1So0lDAz3RmZDrJCa0YtxsEH0E5we3q/zHU4Ionv7QHlLOdlIQVxTP
AFCKLExNwpJavfLh9nO6nR51E+7Yb5vaeG2J0bHVSH0mIKpKUgfjjVtyPCJatF0G
ekaObfEU3f6gJ1ZzS7Uk3ECoQtNEY/jI16wCzDJiVeu+pC8EgxsG4pMLMOcy8XMm
bcopU6e67e+IMXOw1WIIjKuJzHyH1OYHcH5olMxxDFOiRTrh/3T2YrOSYP1LQb5e
g+c60MgRq6e/1yqVlOviq4C6Fz4+hvm3KzxOz23OJJud5nWFYqldad6Hf2dHchIt
PiiyN2HJ7QGUw22xHjKo+SBCUZ3aNtFZpQ3NgLMKRlY9xVCG88gZUplMzux53+yH
4jPK2wH9lxA3OU1UWCRLQw==
`protect END_PROTECTED
