`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lkK03PKOtwMf0iE9/3V3IcMCI2E2pybhk7L6h0D0+5VrvblgDtEQu0GrOFy0PAZZ
hDdCDGVRo4slzOnaFZb/tSjGpjxvSPiOGTWNpxJBIWFWl7tI/laRSP9+n2aU4KVP
0naX9KKw1+8zE6I2DYGtVC9AuIFr/uDbah+DnUKmZy6gpfzgFnsYQCiRkccAvT1Q
RzToBdn/kWSo2vbQ4kJhSJDWbaV66kqkcQeSuI1WPlyNajx+suomTOJziYRq4M90
BEL9OtLhzPxPQIf/kR7klkaahiYHeYNMLJWUvayFhrurAB7h/ROMfHMccegMpJ/z
NzL9I0wGBpgZ0N/b+iD+OyENJOglPCKcQ/jYPVZWCb6uoSCCxg8ySPKiqgo+uM8G
qy3dQ12mGl/C+7Z8VGTqkTif6cxAtboQMkzrELZkI0NkjmO6x12OwyT6et+k7++N
1g6hPw/+9knXPMrtnvoAsYIfJifVCuQQEil7jf8Oj0tA+iYKcUs27XQwylOWooGj
EKst2qGEdMReEWFCE+Mv7221Nyp6c5WY9Z61Q3L7sCxDhdRzVVyz1Tvu7He/F3rT
lnN7G8SH15VNoMayIaFJaK3T5knhtKl9u0Vd7Lk1lfWYpG5+iLRcRwaqmS6wyMMt
Cp0crC5UkjDRiWEku1z038JdbtAKFkurnFH68XHllNZ3a0K71PR+C7xY0g4pJyBp
dsUWZcqd0G+kIllr1WDXxsopY1WfY2FPds8y+t1Sj7OpiCgxGRtulU2pqlRSFKC3
hKSAprgk37nY1jgOZZOwFNkIteZgtdW7zatqM7G3VdMRfOIZGjfxMPuJkSZWn93F
gSZ/6GVRzuJxWzpl+l79iIfIecb/1DtgIcy4asMdSHDsYSGT2Rt/upryXWeTsnh6
q4R32M2MdpHq44sHSm/zwGi03cUULh26LNZU4zACzH6rEEkbLD681xMkxAaepKys
2zFFObPcC1d846WUs9bALkAEvh6Uj7vH9u6iuvLZNZZo+egyAw/Z9w39TNTclsQa
io7dNfOCqL+8STKsU12y8nYa/cDX2wgNlwmot/QA074rYxa0foapU7/L2MBO6yco
16VeK0ZawVuxYV+zlxEE/rtUH8n8RGIRzOUw9wZCxvDpq5uOIlP8HHYC1gYunKXv
Yu0PUDb8uAW00M6cz9i1NcD6hR77OluHF640dVezekp/32rqG9rtUCZdWjHELSRJ
2s0dhl54jotonT+6kn+fyN1AKevUW80oTBWgcoYRkYlivwPYZuyfA4Vzj3OXw/g5
QYPo9o5FbCRpXd11NSUZ1IWWwhXgYob5ixkIqqGHkSsxtBeMy5ERVHIKd3K2J0VO
JJPcqMK4ECIMVYI5bC0aw1XvsdgtJszN+6L0zjrRE2KaqCGA7oslWltrHz7rxqep
LpRoNHUQvpzUd7JH9BAI4a48KIRpskhHMG2062gV15+sxmG3sXiKoFsXgrf5Pva7
`protect END_PROTECTED
