`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uKH3FTte0d8vZGd3pH4s7o+1uUMTMZyPVF1zUYxHbRuEkxXMLpWhLecDv3+4Hxut
u8QkeNGeYP9xd2tGRSrP8CxqCtgDR5o3y3aDkzTIef2PYRUUwY+6FzvJ1QRSEWkU
hwn97EvM4DxMC/Ia1z2ruriixim6q+iVzozhw5jHnTfZ0/lvsWjDI9+mR74W/QnM
FR1MgPi3+4J2h9856yelk2SU/0usfuaoBo6Q9YSRl5+WHwfy2MztPtDd1hmCCrnK
`protect END_PROTECTED
