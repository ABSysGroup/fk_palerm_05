`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
18mQwxl86CKcVMFgfHWP6CmGeyKK25zE389MA+tm55MUqDyI3XxPACXIqSOUZeH4
xesh+M0NOZVVp2ua6+2/sKceJGS5VCbpLlmWY0ci16gA0vFmSKP4EpbYL95P9qCA
nxg1gU3OrsTOPGc95LUfIJe2Brgw6ND7Cl6UotNpb+zEStbr8EV2grwTWDsg+Yv6
tT0hTFJrJtH77PdmvoXL1kkmlcDDby2EXk41QeXgqcgzVlNnGgFHK7JSYEgljKRD
NlFY5+5hL6cQ10t6LxOeb5KzHlFEJpNG/60BWwP4nlHnJ0cnWte70uFQ0LCT6JI/
sMRs2ezUbdAu5YTn63G5RW0pelDO+w9lxI3RC6UJ6ApbW95kMsXwDTbZS1dSe9Jg
`protect END_PROTECTED
