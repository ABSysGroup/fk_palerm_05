`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9KFkOchI2F778UjbOFewV5ZLC1uyod8X75DUwwMUQoNrRUWDaAz8FMkLjExI9Ry0
snaMA/CTMp8onI55+Fot2VYntEfjWytcsDWcuN8bn4We4hbULj1pYfs3tshV8Kgq
G4KeTPU45xeOZmF9ZlMSLR1tlIwzL0uXXuFDk/KBjF0HqQryHMp3O05MiABdtJEL
/2yk6K1PeRIze57YPUIW7ivslgHuMPcJ0dS2+fJSDeGb8Iqc2m7rosMqkjGwVTQ8
9foFLGiMZvAVSJ5KWvACf/rVTCK0l7S3ASjd3BRp6tXCRBpYS8FERDhUVuOIkt9A
q1obBpoJvoTXflFvY/cZQg==
`protect END_PROTECTED
