`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nONzZy+7vO+W/e/C4PwzqauMsu3YVQHk93w0AICcjlP0TL2SiKLddrvxK48AAdxE
Dg1QDHF50eTpxaYGaa6pjd/U3ctvj2SJlL7yrPZSbueT2xJT2xCb7AK8xVr3TzK7
rY+ylcBO2Zw2UM3RSwMOR5IP+t+FToR5OGpqdEUyo5zFbtm8hDtNmUMXolg5jD8r
P5yy/XE39nDpyww8jNuLmEnpQY8g4+HCt+VflhwkMf0NxVqGlCrL2TKwhbNSRTCx
`protect END_PROTECTED
