`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0aMn4egHcGKDdR9NTEbE6rZlkUM7cTLklkSrNdbPqmNFEWaQDKp6rZ5S8STr+ow1
AW/ZpCvzJS5d5+dqfFk+mMV+ptzOYZkm7pbYehCgtL7Vu1qT8bi3ai4C9GmuxpXq
XdAdIlg+a79g0O9dKVwXbmikheQuHLDvcAprhHU7H3sTNhPhwW7ocvDdvD0VR8I8
qIYEfJmSgI8s1ndBn/m7+tsQaBfoPnn8PoEa/dc0c/RBzfbpgL9xBR7S8QYzA++f
OWEAWcfI7dslLlHhKZUAr9vrR7+v2fzfMfGXElG+X0Z2uk/1MgInmYyIvrgoGlIn
H8ml6fVY1SBELCSEyMmw80vXVjRuPCKeReX3YOoof9k50IV1zP4Q/VOEIfiGJnin
cndTYRNefyniucTpMtWrVaMScEQ51+7NBVDMNKOEnO54+gxGbjGnMUiRoXep8Jg0
mRNWq6CRQhfZ3YKMqF5PwXSA9vCdeoAaclWBVDQGAa3+GLQTk4Pk4BvJyqLqNG5b
TuDJHf7H2tXCartr8gupNtw+xiiWifY7erazhZNECVYg53FhojcloaLrPS4FEUSR
WT3Uwe9KTlg7c99eyQzuinVhGFv1RSa6G4AMr9Ym2mXK4cSok6zClShh+ComRwZX
a9TjRMiv7wHtPJjc9rEI9rSVEYfOM2nEJfVjECrxTxubHg1xmzihMcMOhgKXfhgo
CUJfE4K/EYzwYknPC0FLYEwdFpo+7HAihppY7GxnSowHx5v3na0m79w3qy1V719q
gSfFAAWiWHHbmv1FWmoE40oOYf0Ubre3iHyrRzI2bxQas2a+/I/CH/JlOe9fUKy4
MRSvviGwXsVvJWIF28Rn9Z3yxlzvJ8M0sY8lUFKS5Yi8ywpkLAU18ezqPu5k5hNf
AoS6R4GmBHeNbYIQ/y5cKXdVLhBFCYAaqDDUSKigjcDjWGD3ejwzrZnN1ynD7/JD
KxiM80tNOTFx2j2c4Fl25vjHjR8XAWBcBJrSfpDJL1i2ogvzDn2YfzNQcW0YrRxf
ekEK2nGCBuiWbV1opwUhbQ==
`protect END_PROTECTED
