`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xbKfr5UFvXxI0D10ihhzi5u/rJmwvLQ1wMPYle5scSaIcSv5tY4y4IrH6k2KzMQk
VFjNPshcAdv4NrOAvtx2dmBmvPZW2hEg+PDVwCouCf1m67BL9RNRFOm//Fo8SQxG
WgAQsw7siEResVDs53tNddqxjCnac5yiwyu+na+ffFcdSt1rt7/h2SQ7Qzrz9ORR
Lk5CSVEc5AaCJLvpNw02riRSA6oDqhs6pA02XisTJ3UuUDGDQIoev+2uB0aXpaTw
FRJIeDj2uKrSkMHVrxJM4JKWqbZgXSKl6P8ISjKQZQ+wSLj5IPc8I+Oa2GRMv/H1
b5aK11bLGo4BGPTuv4qx5ZE0fVa75YdqMqsBq29tcaiBTqNGwDKpC5tunxou+jrF
aNHzZvRpCD5J9cnNu67ponnzHxIvvdJc07ET2ahirum0DmMvPBQk3XkMKYm5WxW5
RqOy9qm2QQqDX2PMy1aGzuM+9txlC+SywtmX7z/FA5je/fV0XdoqtO+LK8uZU+ya
J25TyJeGTJFx0Ov37JEn03Z71lq9t7yUhekoinvnqOnKyHQzxcXkixga8GfL6cG0
hAA/9ZUrdID2Np7jCWpg1p00Y4EtCc7Ubz8jCAd0kQ0IcxoMmEmAoTC1vdg5KWhQ
Y0mgwyELkitpHe96XPO2Jq7FRV2PoMV6TrXIxnqDD5pFoVfUyHS+kroeX9NVYsv9
EQSIrmtHK5yQadoAnxMtKpev1HzkUJ/0bH5XPFjelkTs26K7F4mNG0/BqNUH5RFy
vDb/EUxLXFg6KFE79b3Kkkw4+/aWdgmAwWqFovjOL1rj/gw2tokqDXc3vzKcjVKv
ATOqjAqQVpE5SQcUTtbByQGE1GG0A5JJlSLgJp1VQZQrdyzPk1TQrC6CWSkeIEhH
q8s/AHBZKiabyow8/oZ418OH7DcqxgH1mA/e4HNwXEudLWSH8wG04IvBBT/7o8oE
eJ7/sX/qKrRFg6SNfmCEufV52bjRU4NOec8dPRMyPfBFGAv5aFlkGJkajNXOgLt1
9761G3E/E32/xAbm+L4HFTiVvyksavwH8dfKPlU5vkUrWW40/Bv6dULixrQStQZL
ZO39w7mvUKmBgmjruxdsMGB1GNBJNplkgrPt9wseOetyb708fQxkUAihDtf6dPtA
Py7MCkIjWx0SkUUducaU75lJWbZkH84mA3NfTntr+xldtVjoJjYwsDaRFKNvnaTm
BwFkFfMwYUy0QK3oUPrsSnaDCIzLnNY+bXJyeXOZ8nLlGWCDXm68JSoUhhRoHIHn
bs9T/EJy1qm/LPvrOu/sKzoj8w+5wfaub1sVd3CZCqLukZXb3Ndhcj0EF+D9JmIW
POWUqNMsRniREWgpfiVouPbHbh8/FMDM7HOZPKpgGPubCCNyE5aokwEckQyOkXYf
G2LWobUE58rJ+bUChi2eAgKmPekWawxBeprn/MoxLXNWcv3ObYvvNeuRelI1bfOE
1LCnJ2TR8MrJiOz0opd48l0ogdRZ6BGRIUGG/ffxRICdTqfsJ3/aDWlXgvAVevX8
PsPugdVjkpGomfoaCpDJtQcNdzWjqutcGaauJFzXtppwQTYTOY3UofQ7U+GL/mip
7v2U914bYK92uQ0t9azSW6uhn/bR9AEeq6YY6cFMWdygq4v+RmmdEAT2fj0aWTyi
JUhbsX23vNm76MVEXuQjk47M27gEBO3nBBrg8fYdGe0zWtsZvGeGmfDMw2xfok71
3UZZekXy7Xh0AB5JWWsve3hTVKoL33AC7GSIx4aN55Hy+/CsZdn74NPiIQhDCry6
J1Rq51+wVgfadrH9nxXKSENKfXBI8uSW8YMvErQkjxYSBo2xRDMbEIynkGI2DqJp
WgaAl6D2pmHlQvMnylxOG6FJuqOYvkto/FWZSSvctPHEib15wMJ2s2bXKA8vkGUB
yG6l4D/pJ23kIL8t2Oimet5MTfvdpTzrxMkvYEQC9y3YJxCGZzwxZpyEHuXI/foq
41NN2ClQwmQT9+VGOK65+y8R+NRVJiL+elJhhgCuDemCmshJ7qIjDDWiBPqJatd2
XL+72UekF2akjOmEzHobyd07keHMtSJTOfGW9skzUKtbBq2Jbb+9qx/O/d24Qfv4
ogGhafcn1FEPPeJNHV2Q2Mk1T6hh9LEfZ+JVIeM30cdC6Sk4trklOB0z1RwKRUh7
lIr98wrgTYW1A7QwyKz9bvUAlPAYnzrnkWKx4BgHqtXvjgosIUax599JDCxWmgBx
hOjda74tcU4ewnfQQcg6gkkIIzVeNJD66+lYQjtuYrCc6fVffzHJqwtlXUi+/1LD
C7WdKDBLlLF3yLceW5UblIlBWu+6xRXCazMW3F6xb+tCbiP9RcOWKNxaV1hre0co
vwco6qY74aQ4RABSp+JKQaxFSJedlHmZZhXOlIClNt4UJNCmNVzh1YZTaHvG/BcF
UjXkZ971SVTrEQs5FJHG8fZQ++EeqXZKu+xBBcmV+lr7FUI3HRiytX4QAADkDQ6N
CTHFrIC54txO/cpI9ogQIcGa/HZWZxQusuqTvY0QaonC+LXdDO/2wzbrOXsLEx5e
Vun48jPProzWoHYPpkpFMg/jJ95Sqsh+Dfjiu4x5gY0BdI5YDVyVSVW+Wmtqr+pm
02pW/TaNEuq3b8Wl942Rgbv5ifmQuyabgZesnsZmh8uHYGd8tm2GoAvCNX+wt8GQ
jNeJUXCEVjXHAac06+vnXp98Ys+r1WMIOYLP7T7uvA9hVQfjKsLfYKSADTMtcFok
fvgoPLQNgOmbc2NkosXrgrzfUojRl5oOsDOosPBoM7U7+Ja4TQsP4wpaEXa/qTP4
6GRjoNlzL5mw7BmqkzkZ9GU9Q/7HZJAp8eSlzsEmdMChhlwpYmT0vAfg6AT8s1jH
3lRrREmuImhrCeSMglUGzLF12xpxsBtdXC0kdq4NqARfblv6DOuGKOJYnQ58gucm
DTpiDV+UqaeKR99elvmumheKKWHhD8xBY7VmEIt2u1prmo8ZkHZwONTK+NmjyZO3
acr5LCLRE1JvczQymlR0F/Fb53EZfgXVS5tF7VLVncH23QodhaR7J77zp4SK4PFf
kwVKqLYoXdBPREbcLcMZrKgZv9n56VvLejhj0nuZWLQePoU3KW00ZHDVcqEzdNSW
clH2g3kE6zCFGZt11cQEX+Uy1lk1pIETpzeay1ImfH91BU431a+PqlGV9orjNfes
eEd6yb449/ukoyi0MU6Q4d+tt5fi2Tk5A6NcS21TfQaiZff4UO80SMT0BU33/vsV
ZmPr+ZrlJtW7seV99c7ii9Yrs3GDQfT5RS9TN7Ip12oiOGrUBqOLTK22ALNzrhAA
CIb7DUuOdJts2Ca1iIjNlSZ9t8PSuy9C1hhUVRndXmfUdJThugBk2tceJrzIaFVa
0B3wGvH5nW2TNlCPwaBvj0UFRhqBUXfyxbLswbCaSBF1wnCIovFdArBtPuXo0mOR
JOZejw3JXqH5XWDcNH/19Bi00woKIhGLbac8mCjZvM1Ek98q2Qcg4fgrgiyQyor/
Rtilw8POHZzptrlxLJRUsVVnlxKfxaNGldXZDBn749ENDnj/fC9Md25QFIW/4bLD
kA/MKTWPFog0rINBCC2bRxIpQx/HqsIs2fEeyHQ/9DbX+w2D8gLY88MUFXP2tOUE
xV+T5Ifdi54l6GDl6iI5UuMb+ZX4KIF+zgq7ccAg9vuChKthGTvWF3oMyBc4Al6U
aYKxPRbwYnAwORCR7qN7uy8Hf2nnqZYnxPcm7YBuIh4AKOC+yqI5/qMHdIwysFR7
a6pSoVOXtTfXVkl0sjnKIi9cAEjM7eUY6gFYx5tPyqBV5NaXyscgsiUMc2Nq8TjQ
g6+Ty4SXG0zhfmkMTJ5NnREZv/C50p+cGLlNoimB92z+lYzi4ET48jOTAz1vDq4O
dxj85FWoijjuelRK6wUXZKECotHsRA0oJa5u9st+y+hqrNbytJG3A4UTMJRTFppm
TVfWcJtr6WQaPKCHNKal90BCMrgvJD8rC9dGlhb68W7fFeEWJisXpQ8KITapOfMF
mV1H1ifY43FXnyvlNJZb7O9mDFxwZ/g9YEDBxwTsCuED6SJNH2oJVGma/LsJVNqc
`protect END_PROTECTED
