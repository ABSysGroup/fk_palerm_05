`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T8qhijXWnovXKKNzLQVrJdHRdVVKbET5kvE+8mTZZTpbvdakOrxBwiFXfnYDqYxB
Dl2+yRhiM2sjLwNCPDQXkqK3sIIHaP7CP3KDNptBnQc99iqs0J3KTAGnddGWGKYp
I/jIBn00SR7YeE2Z5PR1vrNDjfcWYqw5DTbX9rNdT0w8iViFWDVDxR8Gg16a5j+O
QQbvjZg9K4BZmrkS+UJNx27jKI1n9agaNNtOuGyJBfB04iOJepgXV9Kc97mxDoPz
NTKAQnSqL0IWaol+ahCruQbphZiPAhC6WrcAiM+yJxK8UMiipSVKsL7TfeqRPtzM
ol0N9AF1JykcaQbB04Gc3G5d/pIB0OwrM+toZe8vqjuCpuN28rR6clwtrPnDBr3r
2Z8CmaSxpjxSEWuvjAWpwiTx6tbpf2asGlQiEanz2ALgvWfwkTOcM0bsoPxo3Cvv
rNDPE6AOkaWRkoZ+gsHuTXF1vhU9WoWNkEB4X6Ut9OeNXMOuFKI9RKg6Dpekh9Lo
2rg5lmNMoIEGSiZHEZIawwcZ3HUaFxRqmker8X7raondhEPpNgbxfRMjMYsURb+P
JFK4CdqrCHOk28JLjI8jVPRgkjO2SU4yfGgJN2fzO6NZyuIeBmol0KqqEjU+YeH2
+C7/WFVSyX9SR+P+sGySETZ/n8kBWBQMXhM+9FJKj6Yp0dIkYIQhdJr/NDTZIwUT
xzP/O3wAPACUgUC2UauajRKHCTk4X4uS7wc1KppXZ5/uBqWo7Dk4a3xo8fQEBa27
cT+HfYE6PwMttJSxSmT4qvLpyZpAA/cx94KpQvWas5oxUuMYGJdMwcfhBfbqMzGD
NTjttc1NGwvnuRdfaZOeVM7GqHAPxUU4HbumORwEKvyA3tbPGBR0E/fj0bqYNBag
FYIZs+WU5fde6qidRYVhMJNdXyezZDukmR+1h30/Gy3oKGCCiZIgeZVWsr/zCV1s
nDxN9ltcbiD461J2yukZJ4uiPU6l34QVdIdIUwt3T4xUtb10E2OmBjaDLYTTTIYU
V9CQrDWYYjivwx5NO9EKPBt7jZn3QnYeCajQgcUp3Iz0P1LwqHb19X72o0spvZhC
3luw2QT3Vwx8zk7lOSCf/zlj53/lIhkymGC1lmXM9W/gGucvRiOaBgep8QoXcw+L
x0DZUa/HwGxHvHzg+CWtNQEunkc8CP3ACQAE62D5jhFZFz+Atm0pFbg8+KK6sxW2
GdQD2vnKOaGp2q8UNIGA2Qsyi0zbuPR/tbQ4meUOQPjWr3e4u8l5dijIE5iX6gXS
iCajV2/amZx8oJwv366uHaHsi0fwLTYFKxGSe06gH3ESQ9WYotkyx5uZjyZCEpxE
5/Qc6DqTcI429V9HAhkMziP4GKYu0yU0myy/7ymuCq35Xfmuj52GvkC9D4C5Nftn
YAePLNAoUaGI6/pasnaLh14KOQo5Gklie2Mz0qGfpW6dEQxjYR3zj0Hxr6UKv4jp
zTsMl0VSpBBiBgSYzNBEpjgKIQwparIzraKIsb2pMQPMuzLvfE1ky6H+QTnJIEio
XcHCBFnnK7WkWHToa3BHGnkOu4ThJ6OrvK/dWhGsZ9Qoc6ktMteKus5S/yOJeoGi
PjbReyCAmveFVyEwQVdb/pJyTkjgNywlYvt1o/ALj4LT+hIYh1pQzyYuFM6lg+dE
sqI4xx0ywqzhQ+lfCLivhg8Ff/gaYcGRUhv0LaXdSNxAXoJ542L35LLlRmzVsLl4
8ERKbVWDP3FjvNeCXid67AHrZ5GbIeickRyL9MpNbHtMy58ojZKcjMEbHncgFJH3
59RMBSF2C5mGl8apeC9I9cZOyScmg3scwuMAhfJyf+bxFOI+jxbC/Lv6xwbjtpyM
iWy9/oNFPTEbe5lYzCQXQUaoZkP7ocJqmedBiGegKZRGwIp2T4X8Pv3KHLqnvUTy
/yZAqdavBaTFOMSBYR86gwWmSgKroacXv6oju+Hijxz1Swda+zgbiUSN55m/f7K4
hNziJAUnpNJKMWUXIMsZt4CZkJbAdMWfvb7jYm+RlHzFjpK83cov6l33E/s6/PoJ
4T4eUoJW+7L/pEz43k8wiusHeoP78l9ZXIHQlsD8HEqi7bDwV97A0xnspt7UycZL
A/zF1XW40rNJdRn6icW5jdNPTALVPRvw7WddilCmSzBz3WUaB563yGB1ItoS5Six
mAGwq0mZaKxXlFI4RbQtx/h+m+GISa+/ZoCf5JX25WrjzDxf1ymk/MP6AjvCAlqk
qODjqbChj5oaUk3eHPYknKjgp3awEc/GLrFyOScczYISkOYM2eSPY6HMWnDZliPx
dNnPz32o21eD9c4/+z0jqjPxGBCRYU4fSgAZD3FB2kbO/wx8ZDAKkpAhVFiq0Vpk
dFCjMKAa3sSpJlAI5ZEC2xTWXNKYgx0YLK4vvHksKeL2mO0tcQ5agHiHFSt+XS90
CQYTHYXCuM1EaL/Z0awh27qXZbLn/UvTjlsVNA/htKSwYOGCG0Mqy8INXX6IdmON
dFaLALdHFJfnFmL2uYEYe8E4L1qBkry7qrKVWdfQ6xWcTK5kh5w9BQJ1fdi2LkJC
uad1w7HyEBNvignVKNRu25mEFKQLeXW/TeUuLcGBa0qQ93mBblyE2oZfBeTXfrzH
G616h38jbW8iNW1oCWTAdMpfDHGycp/bDXiO9oPKgL2PQjn8tbVtMzec8oMo9Ugz
Q6FSlBFZu2xmIEmLBUHonEq5h+aBiLWaklNGLbcQ1aYPvO5lEFTRRmvkTu4FBtam
2IyUxC+X2YNk6SnBOr+we5abJQikNe9w5TPckDcGeDldUwz3lhTR9hAS/6AZ9tti
GaZ/gNMGqYFFI6QSgEctqnmEA8ZndNJtrU7HOVrrljasHqRph++DMSrNxi8Ilspb
etVwBpxdoAjKPxmOfhJqR0sv3gjEClI1rsJPuhnw/fVpPWe13aLjwoEUViCFVZBS
Gd7VTihodLqYNnrviIgSe/symPP9LT5ppfi1tqcFEmNOVPy3nXf+9EM+6WxFErPp
e1TC+akgXcqmPCSU1Fg4Dbgk7jpTPf0ZWW2FmvkMkoX/ljcSddIO7oSaASdqw62t
Xaxc5oUNt1FcPNH2JZqUI51G6s/DWH2iKQ5BDkmU9IqMs+BNPExTlGYWGArzSYDc
4kfAR22hpqwTvEeN6VXOQBAoauvN5fnpuzQTdvxSN5ju3t75jJhL2wBlgN9CQSRn
oSxT0oTD5oZijdkCcoYaDN3kepWk3U1jkM+lWddwPfAjt79AgKXi201s37w546Rc
ILMtmenNmQWgT4wgOswDaYH/6WerCvdG+HOPLCb85IWWx5ue4E0ph5P42I1vGNEv
`protect END_PROTECTED
