`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BRtsGBvR6vo+b0rHBmuTlonu1l7Njn7fHVoqK5LxBWe9/6cEuUc6pJoFKgtKLTIE
t11CBZwYR11vc5CYbXkCyYqlwaaTJ3rAX1inwrdDjIHAlPRxqytZif/PSdQdzbSU
RyNVbbWzGuzCix1SXAtRQk8l1r6WaWUYtLkkuYSkG+J/jHMEq7uRB9S/vOxWXazf
pJgfvck2en2YfUlJo9JKhedkqlER3ApA9p+yAMjzexFtUtcBRRmLrmZ6yhA+J3fj
nCbY6owYfuXKpLLXDLIg0A==
`protect END_PROTECTED
