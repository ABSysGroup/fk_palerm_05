`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ewo92x+4uTjwmaDEnfFfw1gRKGCKprI2bPTUvltJ5tM2byoD2ZT5EkwrIaAW/JdF
s7UhjhClhBEa8apBAUj7dO2gYQPKy/wBnlDxdYQqmtcOZDfk5sRDQWuT5SQT1fmc
Ik6LkGTxTUwl85Iv4nwxRoGuDm/V+T89nN2kS2iUyjBLQLYT+eLL82vaFy5a5oYi
pGHD0pvkQRRNqoFctJZ+k9oRS0bxlluCfvsY/LhcuexQ9Uaob0BjJQ4vUuBkaNqI
rFixA2ZS+OaCRFjHsEZsH0pEDlzeRzqmxn9rhr3fVTWCv1XI2FUMExCpnjbFb13h
f9II6tO8Siy/5HgEtgwewbTXYVea3fsbhjf+NpHBMkUHTvLn62hU71plMng04SRn
CFlCS+rNh7HaC51KN9D8DTwDfy9dHMNTlq35ZwRkI3eKMF1jrDGGyuaKYkjWwaSu
Pjc7Y3xDTsoKApa02WBHv0qdChQSTbLS6XGQzav5FSbBYK878vX4IxQ3j00vRySa
ikFiKcH23v60cckFfrJDvfLY1alQYu+tv1XgBiAGB1ADRiOsK4ZTIfSb+ShG5eJr
jYglytqZwAEpd/MA8hqrQ58ISr5QpLvKnsatzGeq4Pg5VCBlA6KaUxfCRC2WxrxP
G+Ul4m0SkZN9qgSdfQvhT0yUrLEmxUq361KyTtfJRcS3n2TtNgHskJ+1a/gH6lHs
iid4UdskiAaTSRX/ZgcV2MdHHgK1qPedgEOg4uDNfug=
`protect END_PROTECTED
