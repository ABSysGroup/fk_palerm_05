`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
asAC1vvF0AnRKzIGS3G9siRzBUPzYJ+AYEoYxZs4CzWz4fWmts69nqaScvuNVHrF
OsHhsV8C6suHhOrGZF97unGXZrvDakgPPNQJxpg7tZc7KsZ1y0p56W8qvQTSKzqW
GEYfjduuEAp934StlZktr/L1anR1gV6M8e1Ue3M73biIn+EaOI+hMyGK+md3k+x7
7CTUUQQMaKFRZmxJmsnF9+zx81iIc9hhHWxXgE14lNzlvdaVGcEH83MkzDWPRF8O
f83bhcyjuncyIUDimGejrRa5zifQjSHIpj02gAAIx/rUgQ6S5FEzV+v8MblbivJf
q3nG/EQIdXSY3O6TAa2Kh7Unz3tFeHOOK8XABq/Jf7t05+ZAhlMMwtCqjjXKMSVk
Qef2Pgljzhf/3ITQ1dxxRtfOfSLZa01nuJHHIbhSiYvz6D4nGuEf1TvgteJylldK
YQG1oVMVfJfPwr71rIemhyKBkSIh/kAoYraIGMlbgGT79CoWeYi3dSwfRmrkdpVM
UnZb5owS5b+4+ggGSLy4b6tyhxu6iAGYHU7ktj2+D8arqJgEUoWYMLraM7kNJqNZ
hZ48I33ZlicotsFvVblXFwOmI7Pzd6aV/i2G1INE04k=
`protect END_PROTECTED
