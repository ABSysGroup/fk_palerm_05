`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2THrF6MPEbZysffrdLWICoqEnLPs3qQf9k3QRACRTCcpmR6woNVjSriqX7BQz92h
GbRDS6YbWHx5hU6/lJIMgXBj5DNwSTCwH5MJB8C/2hqE4cxQKvTFGqSkkDZkPBPW
d3sPAUGZwA05CsWfVBp0ysNZFCKnjirlG3Y8x1e07KsCbEOYV02glrwatm+Tzcah
rR5S0W1MhTW9b2/mTW2ToFVpTgSDSV4+g3aHZIXOAVCMro+ECCJTuRkRvpK5/A1b
8eVC9CQdy4zfl0NOL4s/Lr6Dlx+d/hv3GMfGO0RKtAkbYUi8DE4Y2SkHXhVZIX1b
27mGWWc9fOpIX0WpHsbw2N5MGN2EvDm74dU0zUbgNObwG8T1dX760f9V19KPZ8IV
GlslTVLnY36nZS2P7J/LommRKgzuvpNE/Qj/7ePh+P71IwoAPfqNiBvmH7MVHYV/
dXgj/Dh02rUCbPq/p25bxDbNPuAWe0jZiASRY+4k6HYFmnW4wzt1SwBgG0hhW3yQ
RPxHE5L7J9N1y/MuOumOHsVwSGcQmf//1mCLY1JXHipuw9lrM0iUhqt2OBIJC8nH
RssqIndrGZ0Kb5U3icYDr1RFzV9LnihsaxpH9xMeYjJ8PA/cYgJTEmosAVmc8elZ
Q8NL4rxkeJEBIt/sgTGQFs7s7sXp4DGxSfWag88PmcA3sSwlIrHZPc5TWBABWlxv
0e2RdcGBu90f5D4gT/S5kybOO9RsQ5t5/iCVIuB+Hyn8QZDQr+/kzSJBDyeZGLNC
YWj71IGhhKusMr8X/9xYLomn1Zs1FQ1LbbdP2muSwMeDKoN3Vwpxh03FqD9O/IvK
WTXv6o3erUC/+aRyH3axiYXoFOQorqCoj4p6bfZUMCa9IYpyIPR5rpDgMxMqdjDO
JDzzgW3ZHmEpRD07SnwkjuIydoqzcACLeiR4z7nLng4rdIZRWaEeAZ6craqiUnCs
Ch43jtxnRIYVyditDsxilLosKfnAYonnHJIUTsfxVZaLco01H/T2k4t2GdA3XtFy
QpcVSlgB1WoO3ZvjVvdeNCd7gIutJcOPzcScDx084P9XzeDRvhYnwEGO4M97fekF
w7Gke2zFprL74t5PZUvTrSrn539zmeTuBhV+g8ZKF203+VpLVFcBxYmvSGRmI3NN
LbAiCbEMijxp5nWahtfc3LFMToireQWTIKBHNsKgjldmz3iOMOBR4wnL2GfWZZAP
cHFLd28oAbF/Xc2YtN5QwUBD2B1lx8RTfdnNFSxQkI6AqHUD/jcawPulJ3e0ZtnP
ieTKo31OgLeIm2BdHwMFSrEHInx8bS8TJonDfG6bxqbTRVV1BcNCQJvwsKoNFwhi
`protect END_PROTECTED
