`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
78SoHNMuA+4Z/qZd0Cwy+W5fTBbLnVuAXKY8CgIw62/L3xBQBQkQjGLfwVglnAWk
qmAMT9y9zdmV01sp1IPo6RZp3GNX0R+/K0xZpC+MoEKsZq1R1YUE78D064GXt6+V
X3iLrIG2Mgb9cA/2G0INEBNRfLWzm3zt0VDZ6ccV4Ce8Mh4iVjQmcxWm/Ci+AH/m
w5bMNRlxDzGE0l0BhW+Gh4K6b1dXroIzDYQh9P6Iuy/Jk4kiJE4kVy88eboCM1iV
QW/7XvxXE5lZPB2vckTmqP0LMLkMXcTf7Bt9+/IIure7g0I5lucY/YCtRjY4bDi3
huGYWHRQ8E1LVTlFAcUQVmXUeJNvqxFgRsFQrIeKEz+gt54w9eZXmSDnw8Y4spay
gmvEz5MfvUWlJ3j+kTIKxfV4PFMwZW8tXWJZrq5xfBqfJoAzlUFU6TDvzsFVYZhi
jRTiO6tmvt3ayRCY87e3k9a+0qQgvFtfCtFI3/j9lcC5MNpd7yBSevm7psW9QtD/
wQoRj0UZVpe/rEMmmlXht9NNpdzk47Djp/y+BxT69kzAEACaSE5bkjiABJ3dAaJS
z5tsTyw/i/d30liqwYizGNGL1BoimdthMWTNTSFjxbdv2cbekDeLIxSBiXkXVT0w
LgMH7RdP+Tv45rBPtnrkNj2FmzDWPhPOvjJ25Wtj/Xj4Cr7SYxyS6FVBelu5PRZT
HczvKp63TefaBvLrmpyCirGxavgXXdxjquNlT+VzK1mScwGUfj0XcMziwfLPOGnI
l8pXGZtGIi6vLqEmewZi255dRj/LHoKNSj4jsXPcyDktPmWRWJjPlTgStFrXD3sv
fYd4gJRo1AKPuOLw8BQMW9qYQUC5W9D7vqYKaxJBVAjOzW5B4sHPSt2ekA4p7+tI
ZQQXK9nkDHcmb3DpaJKU34RBOFM+dOKCgMH91s8U26P8IVMHnJc/YARz3eT36Pe2
V/3hk77Q6oqsagA4YD+T/s78e03jJ+6leXDQfkbA8n/V7qHoM7DYhSJ5zot/YHia
Xxy9zsst/MlD8hD2Xeb5SlbrSMx4ZaHpAaxiJYVy/ScpomLo6Nr50mRS1UMXxy6C
AI5+8MavNhDL2GHQB7OsOE/hyB41hd+Qtlr96lM26r5t3qR7xbjaqdKIJs6HT3G7
ryKvMLsT5q5q6d8YktppbssIOYd8Px+5jaY7Up0dS34E6XNn5Tucmy4yFQC7nz86
cLvTWkwUCrXgqdwwLZUm92k3nGpbQY1PC7XJsGaxnFxrFToQDShjUEOuO9+mJWmR
Ckz1pW3QXiz8Y00duPCivxxAhqmXpM5GsqZVX9q0R16T07pcyXTXU7ZFSuq8euIV
QGjMKm0/ktbm200xOzBYGXrNYU/0x/jbiKjrnXHz4U6gC7NEi2v/B+2oyHni4y7I
sh59hpaeHP6KylBot3nKYCQjPigNCCsu4DSaBnt8BHlxs1R5D38hYVnSuKtVqhuS
kGVZPb2Zip6BYVxJmI5vO8pkIGsG3n80S6rdGJ07FUhBdrrDVdWP53+gfbQguQpq
eggzEgfcscf+2QIbtN90+eyqFFX/863IJgF3vZTmnxfbT3RiAVpsq9GO+OWjOXBg
rGw2tO7evvSIwsuUFhh3oy8iyK1DM1Aa8ET6QVohwZI9M8KM5LlBzUJhPGydIKTK
E915ITfdgogQ1doeXfWZ9OxEM078QVg35F/6hnCRYveLFOXXWmqRHxV+UEfAxg6E
J1TZOXFJuUV/fR+e+6GpB31rXAlSTl37buF2eIcBrJfmFkLHv4VD3doUa5Cxw9Pp
eNpO29ShXVS4jg2bMexRW+Rpa9q+vF0zYAv0vTpYygr67JOBVkBA2MX5B63YAux9
OtFIgliqgUmTlHKwP81r99X1WrUCjX38z0YKRTcTR+DAlLOtiimWlEcmnja0GOVr
JHKfrcThAaxdPbpWXh10lH3+RI44qkNuvx6xmuS0hXbRFxyu18t/FwxMkUk87L2k
4jUtfmCntHrydEuDdvzzpzbFvyPTdRL0yB9wJ9VfEIP7sUlb6iVt9u84SzN7NvSB
JU9kWGX7va78HNUvFJ2J6Eeovis1fNfp+kymWm0a545I/ZjbjoMu6OQF4tFtoDdj
2TGtQeWnCmiMlUlgtaXBwRrEjyVBxj13K4HsyRjKDemVkjiQ4CLjg+NYBNmxrCDy
6X4gxpVPYMS0up4raCzc9BH/rKR8KVZT06N8oCDrdHlg6prSFztEt/yM0Psmwau0
Jy5efllFYlpUoKDX3AiLiR/rRyvqMXL8RmTWmTyv5pUz5SEDxwG5+zDGCwtVRwH8
PV26NJr7A5Cdo9iBtLs4y53rKsR4U0qnu80BdAzzaLwv0JhW1h+VjU40nRFEb3Gy
W8YYthTLW/xDPnCMqR2JyI+Q82HqGu8kRudu/Prsui9+lIuhu0G2iu1pp/0fo61e
WijIsn3l6XHvguNAsicSi/i+Sr4KWeUBf6LNQa4+EXtO4NfZ8gUTy4eS2euCXiq4
EO2//D8feeqVqbcOw8fSlNnMlOf9uKkbKj7DS5SE7SivtMaZkL75aVGVsuXacTZo
9z1cB7PIav7EuuqVErurRTas1BfoYxYvtj0Y0dqwmY8mDZR5b0vGL7xxGY4PX7C8
VQSPwA6KfpV15LvHhTcWgs7SwIVd5fNqs5wpC+ChTnFk+XeIJ+fg38CUrSbZmtIx
qufCD+rI8mXDtmSDvpvkYr9v0n/prPj7G+F0lcBhEBhjJeg63smYabWZ6+hD0IYm
fwK+sU6nvNnnUcDf4KIErIDOONlL522q28tpc63Nhp8iaXM5UAyyLy+2cUK+PmUR
oovgLWWvGO7GsFYqKlBh7mwPON4Dvm7EdJyWKbHooz1R7kEppz4Il+Y2aO1A1SJs
lxCqKv0OjDpwsKilbNLn4XpC0t4pblVnw+3MBUn79N0Q+8HZtpzb8L8F7fru4iHX
PsMHAIq/Q7UR5j5ohFPHGDvSHOYXzG1tgOCcBg0c3LlJUaUenPW0b0sGbDsq7fsW
bVnrWoNoVlG5nMWSWfMOFU/q5jGEeQKlq0BGp4y9moRIsi7nCcQ0IeTFH1qNoVna
fdw0mzo4fcngq/pHGNwQdwBXLrclr7eyr4C2U9rIo2h/r+yfc/xqvtNM1OJF7Bkg
xfMGay/wZYMsdOO9puHuCNhf7CFy8nCI2KV7oTsyWRvv11gsDivzgejqW8AcGHQc
hZXW5FdyLCJHJzRX2HCEBGRPFzlE2YvGEx6+/OMW/Thn3yK3I+saifb94DVrCRCr
21ZknC3t410IvC6RX+koit/zxdGcu50vvzugFt+5EufZApPtj8Go4efSckUq3tJ2
hyLpWDkX61F9K+vW3a+G3VJdp4pYcSCETk9VonkPJlmBqbB16n3ngwH8yNQPU5fI
UlIuzvGMqTCeWnNRbMaEaq95Bx7Wj5Xu8RMD+NEMq/Og4q44Vi4dKBbPdj/d4Xmq
c8G9nHni5+x7Yq6yrPrVw3ouJxuDqpJjxYPSzevhapliAabSmd/5FlId+29lhokD
rEz+QQx/1TOwbsM+0qm6+FLPzCySiCoZTL4FITi4sPUhI4bdBTdKFYrQQZMffJZ6
0ZFefUQ+DXN6nsrBH09Tebp36rqpJV/6xSGO5Dw/gZR0mf09h/9yMDWPEzYl7hRL
URK6VDYBU9dj6IzdIWitBiH1wkn0uftymh7oy97EwDzNoB3ewNHhCGysJdUQ9g9U
xyDC62bX8dn0oYuraJ6KbdOOoLg/nw3mXPQUQqmgGa2j2Ek7Dn4g/+wURyHQvc5L
HbRKGowYAu+NsOhAyr8WJQvBNnhxRccPEE2Q+0mr3GofAgCOqDL4dLFetzIzSI+r
KDOC9xNxsnGbjW/HIrYAVIKsKjsp777O2dtce0BePeB12ndppbM+2XLZrHzjVBFC
JOQa/Mrl3WjfWTvGmOQ30Xkzm1dGKgJSxFIYv2/2zzZlyvqr2zqdCfZ0Am8Ovy2h
1s3z4YBIq7I25uAZzsRRKxQy6a+WxameL5cphhTnBSUVg7B3vR5+255izqtKW4QX
i9G99nZVNjpc1AP/4y8yZYpcBnhnJuBc4PogGOmKElHAT/iwk0s7GgVz8AFlOsWI
KLbbKyT1cLEy2y/+WDraFjf3COdIAYnyhutLurRVIkG0SYtr5LLaxEK+Kto9jKDx
CXb8pLtS8JApOpK72pmoBQ2aVZMdrYUNM7XLHCO/INFQaNHN/C0n0TGuw7vV0bkJ
OLg6H+gB7QzkavVCqZk2rj1NytU6mWEjMRm+eZzFNjVw/SrSrDTwtNJVeHN+wmKx
VZx1sGjtoS86EYJXVwxP1PHoL7tt5xPB+Q00dwGhypkME510HGfSPvnTb71BP7+9
GXVjSVOxeSgld0BuppUFffGqH1XK+i+g9Jh8ewyXoxZy7ExjU4oSngaQXYlaNBKk
4XEmG7meOAi+LBCtI0v2KiZVhbZXPk6p5yhbc3vEJDR9i1NtBwOzL4qcdHEUluJh
HqpmWQiPzo85q6zZ1JA09aCphCjCVCadq/MqrOEfWbSMukcdjWEHlo/ks8NgO4f0
8ia4ccfBezhNcUcbLf53pNExtEL+8a4kgE5GRXmoSHakVTeu4x0E5/oUZrPccL7s
wgWPZY0gbbmcFFJGEwnr8o4ibcZ+oDNq5T9XebUdsXLsz795xzDxjr3q/JeBNcWN
F0U2ivnPmCsKpbsyi6G259OVDQ4KG5kcFnPg9cjW8CNe/nFgYcZcQhLyaULzqBtS
kkUSv0L5gVsGi5Asrd1BMfusZTKu80CsnEwCQR1nzIQr8kNWkhP6a3cgZkP0Ibcw
1au/3MydMcwfN6B8hRt391Rdu/xalqcNb+pqTWjTUcDlvte8lfgVaXHJ0/QQ4gWj
2qGVbv/CW96FyEA9L664hLBstAnkIjI/5M3v4Bji8stVfGz0bzbVwt2z7AC9TE5e
vme2rwUc44MHqTkyOj426gskvIDQd8iYPdXl/8EVy8K4lDxVksD1KpXqgMb26A7g
VHIbhhuobUh/fl8UgpAKc88A+s2FHZheHClrXxbze1baDD/tZCcGR7ED1lWYGMUi
vdvsF2K9TCSdk8yXYYX6SB9KcRE2aWejEP/igQr3byl6tFnoohFAT5BtjoD8UnSS
oTT4se9iFyaRyb/69oQgtTFeo07QKuuNFJ/BU/9CgDrwaIXpmmaozxVzBk+UGSNo
LsBrv+Wq5VDdeQ08d/FrmBDB6ryehLlRhU1YZagyjRnrSW9JRikZHvbmnj2/ShAm
C/EKPsgO0OyiRa3+2ioZ/21i3q7Wq5VnCec+Oj7K4LSGHqHxPSOzbJVXytBdrL3v
30Abp0O9kqafPWuqd717B7UN2L5jOrJWVkxujhd5FgyMqlCCoj00xWQNLJuXd2in
owAYq0H38Q/CzSLkwKUfJWfZ/VNJZzn9frX5ddubRPxuQEAlFnZxAyCL7bbo+pf1
w/jXOljSkOwYdw5B0HrkOSCjOT3BSXiwgWFxCF5qtajk/KNzVdR8rtXF+Tevbojn
CaxIH66mT5/8VFjkNSuA5b7giiNJB5pAuCWsMrJA8gQ=
`protect END_PROTECTED
