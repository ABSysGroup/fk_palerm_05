`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rCBNYEP/QfrSHyF908v3W43VGWaFoUoSopZBJCcHb7es389ccB3gpuqwgbZ2emsj
EaRUCda1yehfWXZboLootSbKcT5QEaBfUfzrLLeLuQPEV3Kwexz1ktC+uG1F1gGG
uJ2kNNersyeU97JGt0wRgDPdPOyqZWnVnWagBzEQv8bXNAxhQeMOdgkz4vpgcUNK
T+YQSTZIGOxAy6frPrWhNlF/WBAIRqNiL6rAukrENOW62R26zMdDQUV7+ap7Q82S
Lnoz0d3MyQl7L/Y9NqCb/t8YeJLIl3pZ9KVMrxgMYX3fGSou9AUQH1LOHyqvPexK
GG/8spUHF3LF/3l6Z/xUWA==
`protect END_PROTECTED
