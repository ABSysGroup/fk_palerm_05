`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xPuAovZEuq5xG9PwAMyma0QpjVf+ou2QFFBV8XD4BNnIkl9iCyqODnHWk6RfckU9
jAUvmS3dCkm6P1iM+HEkpC2bu2WpaxCC0NeZLD+ImqhJz+UhToUtkTdHzeVQuwvO
CMqFpL1NNTCs6vepgjwjDvnUKkq9JeLTFSwF1pDJB5U0QAk9hACvp1Nszuxwz8Rc
Wqqf7SE7bcv3sGXRV2wKwhMpx8G6s4GQprgR+nkgd/DLZVmfn6ml8Nw1wqJdZhjR
E6y7X1t7AhZX/DDa4pzOe6x41diGmgIEsK7y1rK9b/e20PGChFoIwLdShiqlv+2U
TIwATHRKjS4GzA/EngjLLQXEUXk56OIv+S8/bclV20ctAwO8nxSjKIk8GBaWAdYm
HHi8/OsgVAttIrcvdlPo4DF60RRIDIpemMmgH2TBul5PLNSwxmM7Lrh3Ea93VO8O
IhVjJfecR0MHht5Yp0lCKYGsA2kkFWJJDkILF0gf5/JYe99bFI414irp8ESlHagy
eZsj14IDF95mfaNAH3x8QXZyM/R2NlraSZ2pli78tlF6TEKwP3YPG4nrOK8NDaje
Z5uAWc6FRgusFjXSKjMC0jkHr0ScTLRmdHsFcrRoHJIXa1Dd51KrBcodDWelzcfu
4krrnowZ6ncWo8LpEiSNuhmIDHHY4hZJSXb6f2S7RUGZDHYWIHw9DkeuUC3Mrue0
eNHN6+gN5GEUUI/dfTTV+BjXWNDO2SG26YZ5sd6HvobfJQqnoUfTq6Yp8/HZDa+d
u8XIZATG/bRnzW4Rk0aLdk/57zx4pjlx+h2MMgyYBMKnMKKJkY/jdMy2pNZErmZ1
04L61+CgvykjZF+MSstBK95cG1IfL2JQLJK5yOSkUkMUf7LnZEjc0hztYx12+1A8
/A63slt6CEyc6gpKi5sbt6k6aS4//Yl5+mL1Bt9/H2gx0mwWqFVaSRJXw4t1PwL8
8ZpT4PJjC5X/t7mlb8Q8mES34Mdd5Qge7w5n7Vp5p37QR1jlDubAxHJy8xsqHTgH
ZwlSvrdQlZMVStIKX8e8KDTIl7ckPM9v/YdYjzlDob+PulxIqJoiSPzi3W9yRJDg
vp3hfepgEChoZZJkh7OtIIkiFpet3VrvT5OnaoxxI7dMVE9AZhgK4TOzbG5FCIrY
ijk4FiL4hm1lUONNNY/ZQ5Hh7jjxrpd/g4mY+p+H6TCDKhtpERyIKlmLiXu1NItA
g9cZNYS5B0EwZ3mCjshtd4q5geBDQEgvtkthNprkwBdowhuljyOMqxCgIeFwvIV7
7zOJ5mWlYMyeM26G4ynt4KPdsTrgbWHPrO4o1838Z2Wce2723F7FEDj7uK8Qy5js
ONfhes8sH123I0LfFu19YHnkGBPtlTtlEACThz8e7L7EKfa5iBjU0FyepSfXTpQU
4J2ErEGuIK7Nwk4WFQKihbtmH9G7CCRMXu+9fqVdzyU3g4xG+0Vx9BiQCM2ZjJym
W3j/qybXsGshR9hwdLiIoGsLpEktnL6y38od3ej/5Sm4DgxmWaCxy3ldIQAuXLK0
JdOOk0WZ8bPtpILWFRWG9fWOGlbfzLX1jYk2YTg+1t+SEzPKB75KlFumhHrxlP/p
RaZMS5X4pXBc0ygn2yFP48FLLmSbTdXAin/L6SschqvnRiZQ2uJ3wLYemCHh6HId
0LN6R5OPg/jktpIFBKt1Y66GmfkVH2jIB8xHI6kaazV9SM0u2kq6XgBtc4Sejdoe
mVr7QfnHugGxuZEyuJBO8uC0w8Mc7MrUkICOrxIu9qcVAB4Msb4Izrdiyxkfx4nz
o6ASDi+49qKJyNY5bh9eltybuu7xD389LCNCfxcFsmDm1dH8f5jCm5w2DxZnnX0p
FTwccySbkZl3BKqyoj84kSuQulYfQUKkBtbnJFDa+6DHrtSyqA4GdcXn6ReEoHFi
cHvGEbbxv+Mam1lLDhen5SkDcrLlr8A1QcgDWRi7HQCbWjnad7nOakhMi8jj8u38
BJzFhMhygeMCcTrXMyBnKUA3sSmQNjXajRQ7s2oMv1z3R/Sv7jiNNN46g/wKvsp3
S7YeStIP6bH9Z6JS2aEO23jArYnytVyf33UT+GPGz4wEDo5c0aIH8WTAJgatgxqW
F0OAr6+lo3PK5MqHTVbK8xOmW5/SFwce85KgqZxUhecCGPMzGFk0E1tH01lvY9UV
IPeFExuxsTiyLMYDEoFmGPKusVeNquvyLZoHp0+2P0ZWQlOA847Jh4ZwakBwCrsQ
dAiPH0mYm8YvgnVTb2qr/o39pNJq1d7hDR2hTCCkEnAyNoKHRAyzgjVn187cMNHQ
aVH6HyJ474eMRGIgS4OAHaBcuzI7a6xh0Ay1syOy98QoQnnt5NSjqbAtPXOahu1a
RAfv1RVwQlZAiU+z2J/e4Jna2Nlm3NbrmM6A0tZpR7Sb7rzK0/3Xbr9INAVLOyt5
jZyjwRNwkYcbjKXhKGETov10BJ0HvKhYSINUZgKWtaQOTbH8yKrvkY0a7zNwy1yV
afjXyRg4aquygSrKs8bIN+GzBUJzxZOcisafhtjJWKYQELVJB86SxEgPCgM5LHhu
evYey1Ujg2VMLmlncvrxWiijll0BZK3evwdoMC5rTyT/XojPmudWqjjDxPIpZWLd
Ufq1Jn/RHzOVxSfwILf8RdGyEJZT/1hTR55vUJ4mi16ohS9XSf4NVoF7FU9N27nR
mK6eTxguIg4cWYLEoHgmP3bSEC17cR4R/aU18N1Vw9ttC2snPT0JmqX9iY8K1lmL
5k4vHqyaxNqbp2sKg0yEUEtitRSlqFXBVg5guZrDVVVnZeXseMVk+CLJfiQYp1BV
mH9OYRCNNHqd35nnN1YRRI7e4hAsYmZ7s+uvFPEMu/efv0gUHvmIPYcc3K3ZKPeZ
flSqSgrhTMI2UZV5VZ3oF3r2qfvQbXDjQBBSKI5nMpsY8PYcUmdn2svt+2rI+LKT
4nKDNbKB+lgAwldBknxca+Sq4eYz3pyq2cpnV2Vv7R949pkt2WqtJ6BBbKTvpNNS
tVfeLgqHftZxrJlGpth5CeLhc89Adz8sOO2oJ+Mz/ws0kCuBQ3TkVie4XZ8TAzqa
gDcIsRf2UXN5GEoXieTEcLBQJcWW/jw9kzKQ72YYE5qtyaic/nh6x3rJso+yDvQs
3QiDR2wS5DibH1cR2nlDzFQn1JZ1k45mAssuZg3fvlohNclcBzr4il+QZ+KeRt2M
H5PLQ8F5W1C/NlUz//RzqKLhX3vwx7jh960ePx5IkcurloyXhs3IHD3HaCtalb0+
w0MUG5Jrf+su/MbL/3yzG81jGLx27dLqaIBbSZARpU2Ma+fjITp7MOYoDqAkSwWG
Ue4XHCriRyJeyY2rFCu9xHcNHXkWr9e0k5U3f+b/9iNVzFB3DKhjHkVyVSsKvkr2
vGmwx+NhqgH+xE6aWITsKyjqkA8iJAuDCUN6mRkYGfm8mcrl59jM9Y0D7bfGaCKu
u6Ylc5W11/2ItJKjye1Hh5g6BkzuyTxMjm1k5Rh3f5x4WuMpiUeMvJeqy2iBHI56
Wdv7inSRZGHXN7l4EtNLfpwrC9v3JPiTNBWojzOc+Cb9kfgieNVIvVNz92ew3QRa
ieMYQ8ud2b5sVJRBpNH4XcC0k/gXr9sKrp+PZd1WiCeJ/bC0TMhiyB6BqlnH4JBC
E7K19wZLt8KAR26wcu+UmNZle/0i8KKgdgA00lD+irldc46vfTotXt6iWBqX93RW
041dtfFi7SWlCEiXjjgwXtio/LUj8LeHluhc94pi7r8o3/igekM6W3nEJiA3vDOo
E8KA4AnQvJ4ADg6fro457bzkzkZpq2Yjdaqz7MuzW0c/9lZKAmyoH0ELGVhoBUoT
MXlGywoRnY8miReS2BJjHJQCwVXPT/maSZ3DRe40A3O6LSugkuQq0nd07S568CnB
XTDpv9wwojzZnOYLCITa7OCKFJiM4rCZiBfabu8MBOqcIYOyI/gglbIfQju6J5VX
pIwPZtSN8hd7Cv2nlTQQg9BGWof7pNvhf98SeBlVF77s0b788Nf7NLmT/k8ritbe
scv3XIDDdV8bwZBNBRFuyV73k+USae4CQFBUszQCR7XnL+zZ0hvxeZN/A3Y2V5Oi
fKqWUXWoK2CPmb9d7cHAMEEvUrhzNLG6HkqcOgbJzxlSsYsZKbQ0CAxlbav0+QK2
JqoWbyDPwdoSRXmECemlf5mnPHKZfNCquF5KstGHkkyxQKHnyQUVzegKO1AXKO9/
Rw0vULWREdGvAWhvfBo2zKy2HOxoi35pVv++0VCC/W+JK5OuvHSuzpY66QUp8R2U
UDnu7m8YQpx/pP1TEsbMmqiZLgJemOi+gD/937qe7ACNt6pR8d5ZPms1iUEOrh4S
8cXhq7jofsox/8ASeIK+Gx1Fq+8YzmVIh9n01su9uwiv31uaceaOXHak42L35XhT
s5SIC7aLwfW9vNEu0vKOuHK7LKlbKUaUrn4mMiPsVz4ZkPp2QyIZywPzI8Or5Mry
b2blZyVWfs9jQLtjhh5fAvcZ33UAIAfB60mBWpKGjRjCAxMA+152VhxH3rOwr4AG
RL/YLMytBuLulN+ngCABuX5xN2eiTYuMoG1nfpwjBz2/wA7s9xPxTnZn7Sm50Md+
75Lgvj51Z3N3uRmMH/S1g6nG79Ln7oN7mBX+5ZBATws5U4cjewl/mOGkW8IRlYnA
ki9o5LWTI0fOZf9MI0u9GafnSKdfftX2BjN/sCKr4l0tTPlj2u4NL/sfL36xO8O1
yP1qWBoUzDk8b//Xbhz6Xct9wN4X0Q1uTEulwdxSCtfXHf8/Xg6/dgAjzlKuSXaw
fVnmrT/dxqieVbnT7UX3SoMHMb4RGNGH8U75HDU+V1okiSaIP/eEDf+WmKxbwynF
qN3F5/h6dRKxswfReOaB75wTLD4q9Zm4n66D5jS5CedgKsF/3e4n/qk2xdl+NMb/
QvMy5+u5f+G/kfE6gCVQLYkvoQUC4m8z4sv8XQ+vJpkxiM2AxAuJcXa1LFrEehFQ
5PPkKtmRfmpFurtoccVyEbz6flNAYOB/SqUWz74jmLoniFmUAh7CViAPGOpjAhlo
XRpcq1TycedjNQZl6DiocwCv3BE9mgKKl/XBoon3PYs59sJ7XhwJ/QHmrataEh6/
rE7ZdnzW4U3y6HY1GRcxZrvA3a2PQfXyMDz4aWCFHsxTsTofoudTExnSE5q/LqcC
bzbjTtG85CGBP53ucjbiBAf9qzSSfY1aHvMHO3cjy+rHvJ4s/6+TwE11GdiC1f3V
PJtmfuz+itApCH6TF6NmTXZuLAXOq5iEQDK6stX+IY6wmluKMfcWwKVP0MugbBVv
rjmkgEOrNbCeMbGxhL3pEnK4tDAscOOpoV6tDnpumEVgPrN5OYRAnh7F0T0s146r
IV5ktykM8JZxRaJpkIC48cosw9eSEA3t/YUJvKB3athlgB2KDdUWDnmeU6lHfIo9
njTh9kAsDYyykPsAH5wG8I1wdjJPV2Zh6K8AZekiR6/ibAKtjoV60T8T7ju7whJL
+ALEqWAUgWys5hmG5ca0TFtluMjRx9eGccUstaAvO8hgJQP2CLyS12Kdwoo1EKSf
JaHDXeXeY9GYlNOqPQjdOx9PdaBz/QHgEklAgfpXlgP3a1q8R75L9ryfnwxJJXfG
nyL7QTJB1c3Uu5z10m9PPXooHHWsdibkEzwmdKF/RAtrQFCsnj2Rb1hBtPvT14Jm
QFxj0NuOYQl3w7fMWTzALd/NmJrqmxR+7vB526HwQe0clon/m+mGflLMO+8Y20VB
ULjSgODS1aE5BJYtLM7aem3YLrSC6XvBEPD1ecRQKYVCCbDsPu3Mb7mUzSy0EMDq
umfwryuKyhUPb54rkPm5togI+ouNj940m3z1kS9gxsWSG5HbkNUrO4hyehYonS4S
sO1GKaAu+4vmG3JHy5uuVSTJj22l0DqhSOICA966AiBwFF2YDzrScct/kqE+Meqx
QuBnShMKq5SLG9EQ309F+8Y7A8m7s30zDu84A9PBjFO5s0oSh21Ojb+rOolFZhwq
PnWG5FpDQaODN+oSr1qyBA==
`protect END_PROTECTED
