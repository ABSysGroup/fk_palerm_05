`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1O59oQAnHfyIBe3rgzJAfukEbRRvKE/PVazX3S432XovoBP0Rut+syCrZqK6koxA
Fl6GpguTVBMUAFhfxB1fApXKxFnJcUuJgwNeS/9i3P+/n0UwZaaCz6jTxXkHT6ju
y9JnmCNmNVR20YGqJQjfWUW90hOjT9Jp2QDfVbz9jQowEY4/n+cfzcCsX6qu37at
I3L1Du3+ZZ1PQGxj572pTeTaEEud6U2wbdYSex3CvvA/CDec5k4TyHB6v78cT+Va
vBXOZqSsy8996qJTclVavmUz8vw6x3jS4ZUR0xcNcUNAJJMcbQaOjR8lrmzBemVL
/b4miF757jLHJbeL0X82kwRVGvGJZUmAxP//6hTw4stVkql5Ss/j52OLaPLTTyUR
wiHJmwoXsrq2qnP+fqrC7A==
`protect END_PROTECTED
