`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
36hAigLH9/vM9qTaW05+zWYHkoNQmjuXVH49SyKzp8TIieGG7Hjao9awpjdHc0zO
easc5tBCGsSPX2Z0YjPUpSumT/OjpIJ/gJuIG+M3tIk33cdcuAJYd9eYcSYLXe/x
dsBnSVkU+CGS2KiQQ9r0ChLVwHn7XLZX+yvcg3QwGGjmGZ71qvzpPvgf3FsyuZJY
1Q2g52uiYzH9jE5CP0vYJu0SB1SpoQoE0LiFQ06QfhzbALRmK9CbT/EroIjZtc1B
6+xtGRvoeECBQKES3WR/jjnD2BGeFIIGlQ88hOKGAgnIJR6wPL2ge1xK5OUHRJEB
rxCSPVCnOSZJ3+jys8hbHw==
`protect END_PROTECTED
