`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sK04gBxoe1mc3H9pkopAvXRGmwEMe1+g8lqNxSvbx5R9PR+yLVfDTBs9biYnsMzv
8VPFA3bKVKgH4NVghHrigA+MLAXhKGXGI+gclZvF5IyoNEN+ASG6rgZpc0VHJK6u
GT/wRoY7BaAzZnk4CKsSQ53ogpHvW2Fa7QbmlpvEp0PGBSVvG3gJ4fuLqslWLyEF
quX8XqTw/+fp0CM/ILHBcPYVZ15sHxVN5+guPFFGzOv4MKhZEVAUWmevxDqPjGgf
36FSh+BR9Qj6pdDUgQZnhPG15KlCPMuSbkL4Y+C3JTRMF6GcN3oagoABTG8G3i7P
oAW3PgPrrQEQPvS0K8NUq4Bsjtw7eaCxuaB0OKM4pkk/9j0BF//Cn3eg5Hf2LYTw
POKrFPLNM3kVyXYvABsIut08fQvCkCF4k0OLJVI7LB/CRGPp9MDax0IFFpBwHfFv
kjj7kt7kXHHnTAjevS6bE5NWwbDFlJrV10YjV274+zY=
`protect END_PROTECTED
