`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zTxeg/AbIH9L7/yvwBFFFtpWRtG5bv8YAdDArrE091O2lkf/EPm3gcJ8upjpia8u
d+Pwc3RE9fWLjIqykH4mEBInN+Mvn0vijz9Q/PFpjLT3pKn/J3uA//LJCF6MpMc6
7x99HxsaYF8+uYIZ2lyCZN/ogdk4UxXpdOzrqxA8gzHo/PK3M237WQm3Y/riAMUq
pIZHwgsiDAdoBF/ycrK9cS0mxJtwmRcomeR85Kmw25HWqa1NYZwRBcFFTl3EoOnO
m3hNCqw1J/uJBwAIbf2Gp/AWr4o2Vf3QEBKqteZqM0lk8eDVjIqjBnm42+aocT7e
5IuNCv0QMF/JAHj5qbkR4ZWf1NMsY5LSmzpnrx5j6yw5Tphki+L1IURcaef85WAr
PIAsVIB9mn7az8ToFW2bKZR7/LMIG4NljViM0pM2buKUe7vumbTLDYa9w7895/Iu
SwFNpzui7F4VyyNRUxVLPPwTlGH7YVlio+kJU/2s06qGvXBk4esCesJHrh+G47la
6DZKc+h2AIcITA3lFnk4fHW8gY71ctvsH0vVJhUpdX963D+kQMtX6q9SGcj8qb/J
w00aONsO2GT5VsPIsmb0Ml/7EMO7M5P4WGzCFV6qOXMlOrhfEo0i5zp3KZur5hSg
qgRRETwJf0HO6AqyIwZqSP456PdrDfE55N+qzWg6SmYfSEE0nm2PEick6bKNoWm+
m74TXTKwApE9+CiKdQi8K5YEjUlGXNYzpjaZ45WKcd9EgOfo7nbaYNXs7cfVl32J
dzWM2Y8hBMSzeMvsozYdVtgG3VIVSh3PXAfRU7n7aOc2TDwlHoowXyLo5hE7JgDR
vLfXBk60kFINlltcR7IP3e9RzUmu9qFDrfTCU9udLmmX0gKKBMx4ey6nhRwxDTxY
eThgPW4C9VrKO6U+9qf7RWAaxX3L1E6Zcii4M7/7cSjkaDa0FHiA2LHSUfhNZRPw
CRQz6BE0MaHjhkQTl6KX8RxnAvVdyt2ILXjpjQKZ9GypWFgt91UFGbdyU8LeQfJz
`protect END_PROTECTED
