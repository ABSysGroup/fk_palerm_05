`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bemYX2xtcULeB9Oj03OWCIETbhN+/cJLAP4ySBXzrL2Edp7mjkhrftSEAYY8QLZG
GhOlPp9/SmU+11++bVqSeSbSSrob/ON4ogqvAwRJWH7lMDUb6D0xU/k4uukOVo6Y
sIPcS9KYT5lLwd7es+stXeGgSe3tCchFg6wb8eDeiLkliF5CL2mDhOgrjtTFx9h6
2u4CJUDVtZ2ICI6weGCEsB57HDnwHCKSlGe83rF1DRrFVXnjavwqxCxLw6DFKFL3
53NPnJrnnrSIjlfC9B/YjAhvhIrmVD7XeFZUapJRbsJhF6gerjfcyx0GAfXPFLAs
DvG0HT3xDVshUd0Rwr2g1j4dHKf42uwFtab+QYt+pfo51c39xkgU0hFw+NIILBP8
D1DC3E5BtilybsKYtkMU1JnpdEuxm6DQ3zr1QZyT1a3lYwIw4AV1CC+Iupt2qRhD
dT1OKECj9+LwGchRIeElIAVF3/jSAFoLYXc/9lUJv2JHu3/q7xesQqEbWHgo476V
CPCoUuFMW4foHOniOmg0m/PkgUPSUTpgznJbMoYfBhCQkB3sZfPwhn8XMK5i0tF6
eTYQ/D3E10k/8QLDOIJL6iXNJnFOCHwJtv63mAGBhjtYVxvz0JGIhxGsycalBJwA
J8vPRjUDFj1AF5Gccak/7MUl9VtixjAF3+C3WYnlgVKpMm0bqccnimYRpbPAQPOW
mMPSxgUuFQ9yNFPk2yGPK4BjX1KW2kxeQiIyIXQt9+bRNZtDdzaZXjYtGW79lZv0
ryRfwmWFC3UOxlSyt7qZm741ifqeTCRgZSZw0wU2magQmCywrczAiOwSi9Y2z+f9
mPBTmkjtU+f3vTOdvVjbmvH0BVWpXQbq8rGyJIwhDSa1zX1q4hr8phBjWmYhLwLh
3dELzn6Vpo91M+bl285mC1GackWRhLii5WBgAYaDMGsBk6zdKMwjgReW6Rhz7k6G
VqJ39hF+PZE6Ju/YFNu0wrCuzKgsRlUol2MxmqCOn1NiJRzqKMrKza8mKsQ1iFxs
O8zXTAHM+YkGGZlx/wyYdwlTzjR9I0aGMABy7qqKrOBtLcRqbxhIzlUEaYoX1BUD
usaVxpmMNEs+kwM3hR+tFEfU811pFonxP6zGiHLE0XvaItvTuVg9j94a9E2yGSc0
eukot3pl5EfoXqo8r/TWn33fA+Wp9X4x+ILgfOxMJEpLBVL1oDIOFMKRjwSjELqF
XZfk4zybbFOxjxvll2DpfHpDR1EAxHyN9tX7ne39YuKioZbhlX2MWWpQbZHsRmFq
H7ZIhUEsVady4LB2u+JKz8pXxqhNeBdAkEZ4DyO5gDXtwIYuNOl9fwynL8kHMtVm
wxQav5roEJkFlgrw+seH0Yu2BlxRSWuILxISBpNxLVHbPUlZi9XUkfxp9tOzQsSc
6iuqaVv2o9idmAQUtaSzoecl0396iE2PIxlLNU4F5XPTu2/czeKR87iZDlA7ZjYX
v6k1C5bMlQyS0tewvIcu2zdPLnH9h23PEdM2iRoJm/l891fZjlSn04rV0TVbPZRa
csYwwxOVrN0kXOsub5HJvzBH0RxPGm22fxP1CCURgNUqB3vXXrw7/u0O4FX14U0Z
kvGdPKcuOZCB/19gySa/87kVKNGo9PSuMB8Y/dLeghcZFBJIG1JIc63e0OGIU/el
IxB58W/RFdAJG6jlXigIDMxCtQpB0ZmQ3f+JgwfsREoDx525mPGPZYdbgEognfpA
JT+pHLU8zDNQyTBf0FMHTuc/vvIagPj+fWZzCRNzfMEjas0mcjvpdHHYLNKcxT9X
RP6B4d7/DX4+Sqn3fGPlyO5884oS01c0/eM1bN9cWq22DR+sdFdq/RvSAOJAb6Og
3nEfo/+G4Cl/xZ2R4EYXpD5NKe16pasvxQ37+1snY5x5op+09ny7cr7BIk+riFkl
KvJz7LDOW6BRHkxpjlZRKJpuaigLYmpbeydmeb56Lk9lJpjyBOH6fNFZtGQCm2cx
6mO3wVxu8x3MEiaq1qlLKH0cGrqBh0D0Ls/oML/38zxoFc+XOn5fLdZVmarXMqbA
fVuMIxsVpIc8fNUF0mMDGF9ERKGU6+qNfS9v4skVzebvgvoxCOKM/JrUC6MWbRJS
QU8ThT9+nwh392rfdznthUAch1T5Z/QRohU+gtR5uGXhzoyLZ6HgR9mvG1PrKgye
YLjJFpeWmk82HH57I6qpjOATreZB7FKGm9S7Vb5mRo3x4t4H7ViSfNdlL4izcnjb
2eQkqIjeB0HC2YGcSO/HYt82vha+BoMT5T17gi7GnK0hoAeDHKlufWIH1TOX+jdH
EtfEkyw63Kvfx7kDCxUCKh+BBXjtKwRWnBMw9UkCJWMvgLk0y2DPXco7kz+8T6ez
psHAOsz8qe8412WkTCwV27S0bcONgmI3Vg3sJKqWSEzefPzngAm2dNeNCSQ3aEOZ
FrHi9L05uk2IRJ/ki71j/mp+b8s1tSMn1otnvgnPD1JdHVZ1MTG1qMx1sD/7EaWx
yD/++Y/4g+EEviOcRRHh5JE78Xi1tGMDSpGZoqq2VZ/YC59B1i1uDrIeGJqhlSgA
cPor4ahKsvHCccKZwGxCCxXN/iY+f6WKEqVcteufsb+c9LQtev9UvXtBLIvh3zU+
yrDryQw54Mt4NEWMVrT05+ChSHwGo05V3i0fBaBtDFU2E8coxZtQCq6E4j9JJ7Gu
7QvrzlWdBno8tabx1YzpcjOr3nY3fVBn07oPm3zGtYSOINpZOasrVTQBeCSE7sLx
9dcLAGEamh09U1tNJhAeKI7BxmUXowqCq8FcSJTYtB0sgzqg/GxEniR1GvLx5NKV
lG/9M93LfueAQR2WkRLuypr4JLXk7BZxho1+BRjZpOKSdZlaSCu3wgOgKNJC/t6K
3C0mx9AicMzqEyZhUXJ6oQMGkiZ1R6h5ZnS9GJl96v6yx0setCjpwSZ5prk0sm1f
p78bN0PUFc9HRD5T3agoRK0gBkKhvgYWb+A5ky1/LVLf6d1Rc80vA7Lv4pMqxLeY
Z4pMrmkERQJapAl85J+mwfzgSwJQlfyCpvYq88b19w7tq5nuvjxsghpkc2vKG+77
j2jrGMX2F9Rv4Xxx4du/v+cdKHsZE7HNr8vunOuOS13HMLXsvL3+7OYaE5HjASfW
coMjK63J51xTQxPdG3E/3Nj0M4/ACHSsHpUx0Vrz16p8fLOWH60hflQoCxMjWzl4
739q4jf386l2qhnN5lXeNQabaYtjLQYN+ez9yiPtmWj/Mr18lJjWrKoK9BlIcibZ
B80WYG/aADCmAwUcoGJE+tf2/QdNA7u0prug5jrzD56rlJh7pK1/ptIUhTz1aY7z
i1WzixephEERd0P+rK+ym7t57vU+6oFYGesqibGDHPHbcxrFG2AKU/7QEpfyy7Ht
cjiVqlK8nqBXbO0MGJc8L/BV1emc+Y+cEvKxf5o/ZRgvAReul2OQjiYOpZqg6b2j
8qjiNpwR4FXgTXXmR27oPukhydS3ngWhYt/LE+QlzOeL4Ukf89ltBS2D9lFETnn9
qvauyhHoIRYDoSBqdoWhPxecd+nV8BSG3j8Kwf73lYrvfph/1zY1KnoWoRmUgwjC
6/rbFwXwl2eWtvfUvDj7KVWcQLxmYkpDdbHgIwSAmc5Zt/znAP9sV1t6lrEHRdCN
f/Y7JvLNjZEgphPBxTlu8A6J1m2yLl5kSotOSESKHEu6jCVmRfwMKOz0w7YYhJ1N
QajBNEQNzC196vG++Ya3QNcaTQgS2/7OzBiXvW0iz/NJ3IvQt9GIYhob7SXSCqEG
wdGABmwqcQs7TaHw7IVYZZK/0qIDV0adNiFEFh13bXbwQ+BRZRsb2LiW00X6F9M3
Lt2WNjoUaCeLkM+piLW1UtVI2DU33e4IXzixCt+00vqSpkdrHqRDJMNbMwKOK2hq
bLs/7dBLyl9ufeqqhDx4HBkksrAizm00MWDUSPYbbjcyfvrbbeznO5Rk+92EZuhB
Cd+PJ6J6Yz/1dUDPAJz5HI88E/uMqIUgfSiKARXygWDcG6rAayw+H920JzRfmsbq
jpR/GGH8gfP+F1FM6aHceG1hY5b/z9NphL7DdUUf2rHcbRzB3PCiv3pHg0ODE50z
3UQ9cIKDtD2794NoPox8Eu/XlLtVWxRnX3hCH1CHr7UbJFBGgeZqC6vvNtGIAcZB
AY9vZif4TIxAfrz6+WYjG2Ph4zMg4nQM9pV96FIWUr22RbBIq5l+orfWBoj5LBnt
3MqrW8sKEjvQfL5AKZ1f9e8NkyEsduZgBxaP++gl/Jwqoh00bU9kwb0ogBSkfFza
ekCymFl+Wsz7ZdvsagPsH3bAusBgktjOK3oiFo4Oo9fNnfoauWjOLVWgJVEs3mSL
0Uw0OB2T26ZdH040TqZB1iTAQFooeavaGIYfQ0E5EyfIPdCHIY23lVuD1mDRFh9G
vdIa0BmCy5dzop6nESsznk3cgXVED4NqyA0exVet9kMbMiG7h+QN1is+yAeoIWOM
m+AP33ijp+afRC+M573qUdJz3CVjpdZi4bqjJgGS5zwz3yFIZGUtR0Iva0baBAxo
LYEvCAjAr1PGtFvQzM7j7rN2/YpDxVABwvu+m/iwYijAQ3RNR1q0QNM2F6eslNT+
F8Bv45UkAyhae+pm1eJzJ/+MBcNmIN6Pffy4JIYwd+0M9i4whrotUuzN8AOdF0MV
us8W3C6Dhho46jMieJDg2//WrUY9QPDzkwwU4gjeNjR7lrBqFDKKDcerocQks1QR
1avI7zeQbtaVtZIf3IqY2ljyYZIHw+2kChR+VyVuHv1hbqgg8JmnUU/rIWhLJPIP
nfx8VfSbcUbXPGEDlxGj20YLRISyenmO6tNgpFR6j2ZjxhDaEk43u/3hv9O4WXPp
8M7ck8PvBxu9DGttNmMZ6wvYF04bjM+TExSmPszl5jdOs4r7odxVovtBvTy8JJSr
El3K8Bf2PKJ1gPXr0aQ8+v80RKcMKQ+B2Vyw81HGBbA3L8aqB9Rgo4pW6U5X5Wp9
w6sI0K1SLfOtAgeQDHT72scp469GUEEO1BbjE7JlpuyWcC6yc8Ae80WyCBLEbuav
XVoyRpUArk8LvH9P2pa7+3KW6bC4Ssa2Vp4/QTZLNr71z+kUvXpUgVahyDZtlECq
BYiy+hRvW6N6093Oky1MjV+vDbxiP/3iIrcxqIjYxGGMiXFUS3A7QCVObkkBC4hq
Yc6EUbwvhHSO6+EdPwq14azmSHyiF32uf6nDstlsgIJLfZit0e6Wv0gfXkLguYMP
7qM1v4L4yCLih4QeIjU3SqEEiKHCE03YPGHBga9mBnwjHZKSdblqLna1PJReUCOd
uWRnV09HNsYTfny44wPm6Smr/bX55nN7khVflCLFKRcZ9iJQNjFz/4dOs79YHN0P
8C62OdZG9hJBnYLd6aUXk0vPFKd8FEcUoNADBLNviUhHDPllEYXMDQVG7rar1+nu
UoDy5MBADMvtl+lZULsyS8R9HbeN53+Ze0pWGkSZ0JaR/eRgiqmQMJto57K4MGuW
1Zyo+n5GlwXkN2GEtBrU4GCfd/iuw87QDAr9KJZb/qzCuZE6CpsJcEImf2LLpmci
PitSuAvXHS1UcC3x55rp7dTpFqPZjJs6SUILapz65eDlctpvlo9/EIplfGUnKUfq
g8oz+IHugF1LY5v5xvPiS/BV4StWjgW+KoAHRDg5dp8KKeysnf3cGgOgMK4jxBn9
3PULFcNBexOzaSo/sxqzo8gunFA/sAVWmr6r7gFtKdPuagliayD1OsPUTMlaTOnE
4BOc0VhfZHD9BxQQgxDMe8k0OGVGjVQWoolt5a6itZBzLRYXVW45pNjYzS/BJ9V4
pY2pdevavN5EcNsqkCtJQ3N3nFwC6Uyoeku5QhhHcnU7ICz3OSeaa8cMzh9KW+Mz
z8beBp4I7og1Kemw57vP/m8t+Bt69JBno2xGHIIgt96HxHjJMYC/8rB9vQZ7X6ME
Bcxvj+R4jSJiVb+hYT3h8LYLF8/R2XAHp/q1E3DYwcvw8xN4zrKwdN3H1yZgnXoP
5pv3OwMoSvlJmcJJIR4NymmJ0dH61XiT3g2POFDYG75zkM3OVUBDhSMWbqQYytG9
YtaSD0eFumf/w4gUBH0QZI+giuo82phKR0CSkuGP5q/OQlu1h4759wKPOKn2ayiP
zIVAxwekLcPOvnMC4f/ziq1pRAJV1pu8M14BpA/14q+RsL7rC5POY6U2CY7RwZDJ
+m1QB0zjkanvaxc9/cGtF2sUawxBaR3swvicgSG4KwDSaPLzN+kCtFKFdbg/USS2
Wl3NvV33K+RjPoHg43C3OA2QFDWD97OIED93IpReOUDBc9MeeKhGKb+N26cBXJpB
LR8QpT0TMHAeAUMthONG9EtYFH01fC06O8AYmZl2lfT63E9zzYGIPdD4sPFgkjM4
r3huQV+4B6n58MbrKWgw+oyQJ83MRk2EvBsmN3tcKDbuFclDuUVZl3VJL47mWYyg
CRpErgcOKlEcBh7Tbh06z40FxB3Bm5aVvb1yLoIebAt9F2GqVnlvHb3Oi1DCodue
btWe+O7YIIFBb8d0XLQLHzHdsgrHRxibWVBilB/+dk3UlsQl9BMX2S8b8knw07Y3
YssQ7zx3fSNo0T3McBR0CgOiJtgETM2Q4P2bXmApCvaCWRUd6erU1kZXxbILiOiC
9Z/07eEoIrkmhrKqEIkV7YnMSspZrc306MgEXlWtPmQ/LFhrrKb+cO9/35p9Px3W
DIMlmmvJYdm72bYftubZ1zbecK5vpvjPMKuQuyC8Jh7+KIpXmOIBslm1VWyXjZpT
4ZkSHxLL4qgltjHY4bC5jbanZDQxlaGKlg4B+Lc06nGGBaPpQoxIxOBT4tOdVFCy
q0wsVsSbtkMowG/v5433TwjC3zmwiW4DUu8v1OOzscWpXIthABnrz6ZESIPVnDMq
v7SlBkUGD6sRUNw5+A0mg8JlQ14QfYFR4gWCO1JcYdALL+EO3U6kdY2CZ6iPNMXD
cgViFDhBtUlfpM9qK705NSObX7rzjHhFn3QydEu8OGqNJtvzHsepwgC1F67tNftw
CUgJmfW5/hfBx8ofUSM822EQ3rrYvF1B9USLZs6cDsvaDc+l57mAhf9HIPmPzZfE
uy+pp3n06GUGCurXbGbvhBEMrpgN6NMOPRSfg7/zXxdbsBCc6iveorwn50FLDqHq
FGsAJK5w+nT6Ovdbq9gewVxEOP/iJS1oOVYHfrjxs8u2SxgF17LCO9Wu7SizGGQn
LE+JUgaTzgjHOqZyk1ZKNff1D08Yb5S746dQqVuUf6b47pO9i0dYWUXnwq4jnysS
`protect END_PROTECTED
