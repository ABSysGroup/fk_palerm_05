`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EIGow60f7NVSuRc594S6d44p8yybo+/d5hp54PrF03TVS8OjHAxG7l9EmhhTWKfU
V940ymqddJm3GNSFro8VCilgCkT2hzl3Xr9uetVquEjOlvKAdStv6ucPEGyl77Jo
tpTlecqH7at8UqD9Rx4w/YOF+Of8G6evBw3L7y0n0pkOH5/acNqzGVxofm1+AZA1
Nt7k2N3qFj5wgTp4JZAi1kYiZ1fLdV71ZWFQxDZXTLzoASiA/R9Sj0jXB+yjC5ri
fglI9nTO+YY0lNXyMpX8IafBY9nY5cB5KvkE/NnIrnUYSBEyt4/oiOJnzqTUMYRS
fkGN9tBUv86y1EhBwZlLDr3Zfq+5qPU3GRk0DDx50x7jOgOXH6HfhPyvjAaeRb7e
rYhCVlP3Rt9xzgD/4765QHuEZU8XoKcP+FDYKTYqB7I=
`protect END_PROTECTED
