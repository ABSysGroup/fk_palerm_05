`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ziAepL4XfoJpzfpBbkw3kipzfg9qLmNDmzNKQo5F7T/nwyuLB8aOdUbrtI2rI4AK
OaF+lF9IoilEfhEg5ZRmvhQTVVKn6gsnMa9J8/SMeR+fa9WDE1F/A6LGiEAJlpDI
LpWqc+CCYYvb/Z2v4N9vJICBcKQbQGgZtKluSigVPVGZQrXNNSta2lZ48lv7YOQb
5tElCBPJdD36G+2sSk3trTpamK0QeA/BVGHpDQOLRok45DPK3pxIy/RL6CC904dR
dhdqacaJCP4Uo9JXq2Q7t3gN2WWB78C9vHgHiqH9PeDa3HdW7o0mQ+RuxpGSRoot
cwzRUOi29K0gcp2KIfxvpNzRWJjIgl5eN8lXfi4zTNMJhHEync99eWTSrEqQOO9g
8aja4IFT2tJrjNjzbhWisb6LlIAbjuCdZaZw7+C9T1CUxXfC5Ks8RIEeZkCnytsM
w4xlv885uhjEmdEEzFtL8bIk06lQb50wtk5Ra3agGOPbVeBRxhmaVXkGjhhaj7Z0
Ut5RnpFt71H/DuFBkxwjcX7TFSJpJjh1eD/tPz8HGadBXDcBdkyapbPGdFuBOu9H
Sz4cf5yDPcUM4KhWwXPLXUJfvIUSSswXNRUniwJ/THgSWiB5YqarHgHXhXagSIP7
lZKoNwQaR0igewfd39vDa23TTQUK279guBI91loTuMLpYgT26ZMpew/FxoLnqr3c
uHxIf1Y+J0QIe4hchrMLi8lomyoK+8RA2biOjAK/ht20I5PKMbXR4/se83UM2o+l
gW/VwdoApSv833QovRyVz2g+eEdQI5K3MI0h30mqn+VjN8uYPQtgUZ+LiIaUZX7V
xTwhoBBoK5brIMi6e5xKlp4gCBy20Qm6eHBgzjvRd2k1/vSdUc5fvfvqkWQ1ZSXa
9iSWeMpXVPzDSTh5fMKgHiLyLY0LJmJeN52CpGtCv/8ZHQGmV75K7rLXhlg0E8JD
wMehXs7THe4n5FclnkXsbYR3eyJUGIMZ+lfwm8cQ2E36EFoQOIzE4Vb1zvkXUG7C
y6jlzzg+Y4bzpdAm6OzzkXkDdGEoZhL7sxe2Np7GxtnycVV12NI0hKpzxPdd9tPY
8QpEcyUbcaSxcub2cQ1nxpanQ39Vsmn4XpAjjzyJgS++oHSBcUv4D+0QDREYKc+B
Dkgm9jNj4elNaMfeqp7FqewAJXLkIwr5biOEqHuc7X3OFR8zcfHZJTiq2b63IeNI
tevjJIXVLy6L/e5UazzxqKVMIRa9/W+m6arQaqMbTMy7iO1IG0AOYPPFEkoqKC1n
d+24PN6rg3bWQRpVSJyZwSXAQfwv3k5/nMzcEji1CWsFk54/tF+GS269TDVOzHe6
mlliuDiGWkgHAXNX8Swu3BGps06r5N1g24hmrT7BvLT06rctcxAtcScF5gFyvB+3
UE5zlXLPeXOO3UHnTlngBKxHsveFbYbguTohEwdMlg9XlEM4wwkVhJe0A8rFC4DO
b+e3AAXn6qgQy8i52wqBuw==
`protect END_PROTECTED
