`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ocaf7LF42Eup0zq0bL/9ZbJKB70h3lG7kLqc84SodgsGNCNBwC0xgR7ceDym0nFX
Fs1aJlcRkUeb8H37AztuVipTjTKARU0VQNMMDZSoKuQYHkzuUDLpolDDxa4YuNLi
hGDUimrZyuzDqttrl2U17MJm6BWYfj/nrzdhIPILUZJRu449EHDD3lG1ntMiK0Ah
Ywut2qGBNg+YD6JGp2u7VTEICxjZ9RECC7ucrd5sPsEKejK4MFb66ruYFnFKO3tV
kiejwAe0HVcK7cSPdrk2Lw==
`protect END_PROTECTED
