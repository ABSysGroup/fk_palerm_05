`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xZ3ZdDNLYP/DYUpeYhYs3Wit3eboEYPz9x+laox5hOHiFZOnLQj4t53w00fUQ72r
HeJN7CZFlXuidfe+xU6ZVTetDEh81hJbI5dtXat6ugkZzUwgFAWtB9Z1fDU84ktW
6Wg/Be4sKJscSkQCUJblhD29POpOsFthkNMey2Ay/Gt0k8ly9q9Whxp5oV0Y71P5
PYxYc6Rnu6RCwnTRgzaVS67NagGc4YKoDWNgAFG0gY+11vzmJg8D0EquvKXv/zZa
1NTMgN03HSlcVcaPosVLhOrcHXebjzToKTn+Mdf35ji6Ee5dZ6TCpsTjl7TGpCLj
mIyatDKjMJzbJZfJIvN8NdhNhwUZaobeUJB3nCfYQl+dCWmMC2git5stE2lX/Tcv
zcWNfX+tFOqFK3nUh81vZCV2NkQi9SG5Tx4vXiUP68w=
`protect END_PROTECTED
