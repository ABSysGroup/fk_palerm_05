`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+stKT4gRLm52rES3JSLp7pyrvoArtfmwj745puQj9J/0MIqpPAO/M/NkJWI9CqZ3
2e4cpSytVQq+vm2pkKrKVBYm8KC7oUJ/XgSCBkkotKxh5918UsarQ+MNz0N4zl82
+XJhkI0KqsbP3L4C+1N8a5hqSvX2kR12/2a+55KZmAVfbjGmNhrPku3zm5Ngw3mz
HRyloLzApNv2OoLxyxBY4iCdmANR1aEYIx+aNbe0ien177Y4iajcBDvXiO++5YCx
uLLLacdvDhEZL2Kq1umwHdwPGmN87F3tLe7zaft9P4GOwBoedJy+oQ8NlM1pCIlD
tu9z97ZhNTir5UYcdRb9RPrbt8lDWAEv5GbqOG+gGJ35m1vTiYD9CzAbNZWjjm9j
uS32qWEYS7d9z/5ldj+2s0bfz9dSQTcaaRmnrBWxuzlzrTUEsV+x41QK5C5QTdpn
MRCPE/e7A/i3cNJWD1OpnWXN9c3ggKcq20b8MVVAuui+DLV5+WsNZz2o1HhIyouc
RjRfOOYyLN4R+Q49nGUpaDeGFOUMWT/hk/f97oAHApobURPb/h76kLSZiOwAP8fy
jG5HaIYj1xaUgW+es5Qe9S52QRhTL2Cae41S0DRtWz5OSvMnobJQGf+bT9HJSIEO
1dV4WXmRgVyuw9uYAfhoAvB3OxLcnDOFfX5BnJPgN8Fn7WePP9isAq2xT1zivvhP
PNCPHQ4pEuBbjY5mncuowA==
`protect END_PROTECTED
