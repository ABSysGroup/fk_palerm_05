`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W1xUH5Iy55+jcFWNdsdMtSOW0GhXjdQcgy8DugeMCvZ+UNFQ4/Oa002LrHiCyYhq
O1Am3JiE/UeH7zt14DKJpPCOMf4omcDpCb3BM4u52KMX5AUcw5uPQnsK4ip409gV
9vZIFk0rge4JcGacD2hp3Pok6/bTC7/kb7I9JPqrbxyIPxbQdYiX15dWtruX3EZa
D1sWWMxPGyMvtof/3jdrWb10ZUnCz8U2jA2EOTPnkPzOXNgglDhG4CO4coNW2NHJ
tw3AbUYLMk2DBOToUi5fz8PK4ILhRvJhovhC657gSaZRTcTC5JuwvMQ2eXA8TrMP
/KCMsJ/koNxeOX3WQTpyCi7nyNo6gS4kWcUET+cG4vBFwveqaX+SWJVu/X0/9Nj0
NPZ8yHPjuanUbR5Z/frIioOpGAq/YMwoEIBd8KETvUrlWDuLFJnjM2c/5EP9H9J4
GYxBt6Z/PohURP8gAgEAdJAfJmvBFK33n5Mkb1Ner14BXT+niSu7jhdD0Jd+dh3Q
l/KA76UBFT89x94lnTRPggm2tjPjkOEFo8KzMRZYAXZYSx8l0T7vxAWzVF4hwWYM
0oMRp+7rrHXyFjtIuPKgNU9MQVJNE+ljSuJcmlWmqciGTnbCpz7aC+tOXosBlyHa
f2pX+GkaILFzzZTmknkDYsNEWFQ4cOzuIDRWtmrTQCQwXlrRgm5hug1hGtLL8NIO
8SlZcQdmLCE9EZmeqyKQMqDe4HVhLSPB+Y5dqM22JQXgGj1ETePMLlodGn/sU9k1
iJboDjmuHCFjCAPa8C26AlPoBGVSl1sbVH1gbYkHTib77OxwZCBKxOqVfleF9iny
vnRch+uyOux595hR8M6GxejYEGfay4TOL64HiXDvR0fVaW/cSxXSUF+FqXuJvpjh
/8aw+u6C8F8skdCK0P8E7B1lH2pHZalbNQL9SJsiqtk7uDxLI9slC06DKOHVkKwb
VkTtokLVMaxzUV9dVpknmA==
`protect END_PROTECTED
