`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QesVe/uvdPgdBwVj9K7vCR0z1hXiKMRLm9fjU5M3Iz+2Pp0W6szFLN1ExtZd6l1l
m50j3DCbY+OYjnXipU8fI4cHhq5SnnSobWXfon1mMr39zwETNIH+JH1yjPDRJ3Sa
80yXTkZcsGhJMQawzLJ08OBP/yhxlJzJ2cxX6BXGLN5w9rkoUsR9TZu1rkbAqxWa
PIsjRSQCOc5/i0UBdPOsHXjFUwYUhNtZRpwfoxm7P2yPn1IJWpnqWT7G84JAesCv
wdLUr/18TG7r7nXw7eiG2g==
`protect END_PROTECTED
