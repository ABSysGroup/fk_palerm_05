`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+HTHYTzGokgFKmDVLn5DSd+EpSiuiaLALGlxJf/zHIJPi41GpfKOGzowDTwxMwQ+
qEQWmYBJ2gvtKblifX6KoJdTOd1m1wzR63WIQ9RGB7flI5NlR50KghHH5FRV8A4U
velfmIGc4pTUQNCs39YSzagns4WmqZXp7P0U69XfOAAbZhg63hAiPZPeagQQEVEy
HWStzF14KbSglSczQhsWeDGgaS5gzjHeLeJCF0mCrlUB3WFhG/Y3d+wUx2yEN4wB
f7FBezYc1U1PXM8DiANKPVBfw8LGmEI4xwmiUTIWjECjhm9YVwS1utCQFAx07oc/
l5uWZg5vcXxEkRkSLRp3K7UOHmz28LxlcRHg2+Sh+1HGW+5v6DjiMTCEuSjKB6wl
BMKxJ2DcKaC8wDQAOq8D1LqPoiEOVEqgmts2CZqLBnPz1dXtqGbOoZIGuJ2FDhXj
+AbGG+uTkKvI5zbtsXEU2z5fIbxkqXpwGJPUiml9Vjcxh2vZwD9g/pgKL/xBirxg
yoRg7qz2YS4wNhqp+1wm9iNZQzqMVsMwb7RMsEPOgbnx/jkGS/5l1A1zVxVPuWcm
6/qdnLMSAt/ULDQ/9XrjbN7FuX4hGzvXU4ZMSxlZatr+obyCxkvPpzIdOA//ohy2
vjESD/2VvHih9KSdVrV2ugAW4spT01BM7EoillgBFQJnAeO06PT744m06zG16VJX
+skDSuk9nb0CD9SNxERyG1FXAtrxpA+9lVc/8Y9rUOs5a0U2CeyPQqy1R7SYTxmO
aSN4W44Krfjj0aXhUlvnIw==
`protect END_PROTECTED
