`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
26vTkTWK1kOYSylBH4504FYL67JAA2JVqyLmKs/84wnHysmK5yK1GUvgVCY1q5Vp
rcU6qpexcSHpRPa8wf03M0g7es7vVhjkRWcXzGCSKtKS3vie2j0uchUptTxB40Xz
yYuSWjT2PB63R00oPAzkBgAlZpHWRfUA72fLQobVca9zvxDzd+rtSvXQIVSgwpcT
guTiq9ckFqGI5efxNVAfwCZu1yLyu2ibeYeMnWtJYpcKolyLgh4iC/ek5L7roWTr
o9c1njw/4BcPPDiE8hRhThb6vCuCBnjkWhO6sUM1e9s14uRRY/eWNxkC3nZma78X
y/FuMa/L3mxIbSYh2jm/0KYv4+4uCOvKqE3JAV6JIGzKgNiDgpdgGt+qiQxts5mv
jvjDwBe9elgxrors7OWWjWS2HG5a+FvtLbeFwqgdd65YWmKE4mrW9Y4nAUyt4UcD
5U+hbrQtlqr+reibo/Oxe7jI3jjM4Bv5jlxGv0es36+ZQ2Yrkh8tKRo0HieOHXYN
GOhWATHOM1i3pcTYDxLkGFEo/ZEC3QOHCtqcTdjWLpZFVNc1Kd5SaoDfh4uAJiVC
IThy93RN34HQOT0euQ1AAxTQCmNJD6OTlwjsZTQb54ODuLG47l+UegzX1gUp0MXr
Ks3oP7h/AffGa4Hgx3Zfsbug0dltMS5XJW9zLkZMB8JU45lCLtAyCU+5Q/q8JBG6
dZv/qJsnskD2SDb2MrP4tDeamuqxXPcJJhsetDWScjWrxx2/YfKENcoOw5bFJ6k8
Z6ydhqGQqZe2mEX41vf3tbvOYqutriDAAEiOJZF/6/jofjCPsjMPUqbQ+upJTe72
5Bs3iPuTcjSSmUekB+xhyQ==
`protect END_PROTECTED
