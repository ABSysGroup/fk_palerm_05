`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/xmBpMuW++SC7tUIQSUROx4yz5c91hfnXDqmSrGbw/Q0eEavGbIKzVV3cEhUMwhl
9/kmKNR5reeb6aYKdw+LZfUNOVTjRjAlznHahcioseUGHWyLdi8EYlo7wL7WuRl/
QwjVcg39FkPpFz5NpxmAfYWiraIOaaAdsN0kPHJwyNpqpcE94vruOBt2KPp2qdqf
DPm4l66Nu6kJYm0nE6jpxOfhPEx29b6gdyWdI/NrpOhdu+/GdovUUBLq75Tr5ZAM
pH2wc3jmsZpZf7OIcraq/g==
`protect END_PROTECTED
