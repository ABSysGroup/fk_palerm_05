`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oQs4MVSdKZ77UUT4ZLNOtxsyislbJzfYF2NDBX8z6vqZ3Ql7Uv4FYEjR8bSMyIeX
byiSgPXQG53R/E2PqYPskIK4weJxrGw8hFhZG5szuAKXm1P+KdxoCWFjAe8Vk+ok
Y05Gs9JYo/Z9WrFsgJ6lmW32CJdNmD7hpw824/TNLIITBChPMv7q2OcQhoLh0sUM
BpJx1Dk6BwcDacLw+9gVtCs8x9SpUWd62z6jiHjateWYLjqQkFJD3iNd6rPWGXiM
u0DNi7alLrfqeZqdHD204I3MkNK5mEGdzybdHbD5wgJ5oGV9+FAOVKbp1I7slTFH
U8mv/kWVcmnQ8M4LfrRgWCr+jpNCT8p+8qlEWsBUqHOa4u5rIk9xAeTM1/x5awKS
uc8SVy/IIuQ0y5diMw7pACpLq/l2CXwZnZ/YtCtwoArZU040+MCkkpAM+ZDADIA6
OzPPCTq7n2vtfsm8JwAprjGSq+keXoCaYwFD9Tjbc6KBNg6WFIzfM3SeVwmW63qm
iqJ9H7tzOe5WtbzdqE3fAO6BsyhFuVkP5o4HHB+Oo/sLsH2+zU400UemrqRFEW3L
7YAAKcEFBfwS4Fr3M4Io1hD96PR3d/xIfH6UVy2TtD7W6da8iaWDmJvNoL4phIn0
gXvmBthTSUFmHNNG9qSOWV0e9D6bLFNvBggJKVUcP+mncGnbLExngbC0CMLgTR1N
jHi1m8xXeMPbqUuRK8/shaFFNvznZd3yDmd6I6s9hjoaPlXwdZTxaGIoZZ8MSPk0
dYSR6r+DdFTFZ4nFPRZl7WEyO/YzbfW5TdEVLPG7NxK9iMzSd1bBB2NVh1rrCJTf
S6hZB6tKyl6gGfM3UupD0RGUBNuFt4vPgIVNODTKYtD0Ezw3+gf044ndElAL5mBM
bUOw56HmoEseFw2+6AyZNFZjUWQ1vg1vaRgBJ4AEUlE4wy53FbuA62GAmx+siANv
H70O1JoUnuVaH/hB89ZD4haQmlMZBfu1XQVIvpeGX8ENr5KV6sCeIo8Kq8U3Eorq
A0UgP5i4eEoJJMscUyCmGTU2QHwUMleCQXoGAfa71K0vdAi3mrx3DLomeW311D+N
7uqWIX5y0/+SCmPJWtlEyY57TZQqOvRvL4Oo0qd2sMdyTP6vVPLr0iB0y4sSts6B
t4hEklgVxxijvte2vdf/sxRyPluMEKs0OiAjWUAvwP0DqCVsvAj6ig1kYQZOG0Y/
j6/ywhG6scNLo9sI9d73XnuiF1cE1Pfemh/FHoMfxZYKQ+SnmRO2IO9b5DqgL3/5
SekQOJRNvmGs3gFzDTfrO2NC9hX2ddTWxHMH7S84F8Zuqore3jOrL2cATaGkmcbY
ujc3eKqcKKnPWwbBy0e69nRDSinbf/yw+pPTDDnxaMFqfDoNDe9T07bNC7sblDmM
Vt8sugqHEe3UY8q1f8DTmbEM+Np+FVWYDAnz+7ywvJgPSCOX97Q/RRB3zwSLwvlX
AjCLIb+333q1L4kSUjAuIeEO8/4J/gg9hC4Pd+5eqBUtWgLbiWETwrBUpxSiIbAD
anXKIECPs07UsXmaFDl/pJIdEDzVQCh9wwzuxY65aeTyVt6aF2yHDVs43DcwFPRz
Vn/bcHk5EuR/5bbk9+hboYd90dvGOhbdwa+3Al9ELNUVyv6d+roZRkCPPuRzxlXG
H/NUb+qp4BXRSTGjh0bs08TFW1nFjkDkx4Wb2eIf7jID8me8vWbM3XtvjoBUuVeA
FOiPFXcPldAiluFspJmUd6EAr7YcpsrxpI8FJFy33nyTsPXpxVZCB9OGx98IX7wF
K4iZYXE3sDhzzb0KkfvLknc+lq4YAIgCyv988ZoWlLY32i/keH+/doFP00GhROXm
R8KCqNVtzI8QzjaARBs11uscNtz13J3B3KgsIfmKPZNFicHv0U4AasuOUObn+urC
MIvjEUu5Y3jPpDkdQvIdln6y2HqUERmvPSULfstPP4Oo7TXih+7pD5saphJgJqcX
DL9RUQUneGIcdBuD+jtH9cq4pKyXYoUFlOi7nCquLdsgRyDARS8A1pIA1dXKzWdW
yu75oVn60TX8qbbjeNoGTQ==
`protect END_PROTECTED
