`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RuNxCZ6Em7eoyQ5N6/p2zAhyjN7iy4SbjbhFya+s3CWOSPUSqhsfs1bu3aZKKMMR
Y65aThAvcjj9R5QJshivr2wIAehNoiIxJDwwB/fT1cGjggwR0RtbkeWHOybMU0X1
dFwq2OpKDNCtpL89V8sI1/H/9VnKYwyyfzL42JDQm5csmWBk7eKw9SwFy7JbyvYh
UA1sX0KgwbcsuhZ8roejb1xygj62It/sNNUccQZ350NO/HTYNweOlR3Sa9JASd1j
yRVOZdZp5fG9IFLt5KpZk8TtlthyMnOlpc6sn6jSbOWRV7TGbdM0lAS5MpowHiFL
Gng7LXuMZ9Rnz8gCWaw51MH3/PDO9OkFtmKKE2yDyIdrCp2CEe1T/IQDNGfWweso
HlBluDqiS1KMw6M5l6n7Th26+SWmA8xceoB7G2/pAG0l656wfXaovnUIX6qOhHtr
NJdO+Ez+QerooSJot+j3BKuZq9d5pfiG/zYJjz1CqM2XaAhlfZH4FGL+XDLvWpeB
y+X/ggch/JwHexihyvBvNNq47NWMiXcrKZRRyFuQOVwUIerEoUxArJ1Jvpqrf/2J
CiprSeSbNRuS3c6U1stnL42vCfNL/Qm1wlTytNqomePBJyFUdNZThBoDFpxA8dA3
KF59Y1fXXrLq5fwnFyu1Xkg7WhS2dWeFRzq1UPwDaDV2rJSAWs4l4/2xqcYK6VmN
nXBD8YmAIC1PvdlxM7qk1jpIMrQS4+qx2tLg0S9AtdUepOd7AYDFQMeKXGsae3a/
TZHK7+jtW/lE7hHwrP37A3yYDxQUdvL7lHBU7vtK74K9Qayjw15pMFr9iJEHCehG
3Z3Up3HpXkleIl0+PGG2UBeohIOhk7THZoLybhIF4XOiaHOe/9lZn29Q2ovGv7XZ
mKni+sxjRdg9yzDtGcGF7Db0748THp242G7GKZjVcDxiwmb6H5FkR3yDCxYUH1+7
yzCcIpm5YK81mNhAtWf0cRpEwwi+YAxs7EYDTfO90ym+62CyVO1RlyCNfq5RbhCE
SCBhYUzyKhsnkwzsohTvwf0TRD62iZOYe99Xcm7xn15R3Tdb45MVQgQ2pEX/fyWT
c9zbVcL8lUCYYIckWQORjudR5ORkJMPRVZ3kMjgKg+8JQU7RNpscyP7xgyQLZh+x
hpmOkFi9NUzfdyn+6zpoBt/YZ0yr4loZvTJEqsScM1xRM970qOwU8mAjtWJLUsY6
jb0O37vVbHBzuMrICbuwiEmsnS8zW4dQ62zs4VFh/y5k91CmEGuDVPeOrQbAYw41
A+NTQBdrW7e5RnfJ4p+7MflF2R+fik8/SxNzCE8wlKnD5a4Y6waMN8I/4J3JuJER
V6D6wVt3t4Zs97gCwMl/8rOY9EaWVWBpqjB3KGBHPCf+K7aunSxRg+UmSIWl+YrX
PecLMJ4ZD0BESGAcFlI8ylWtKozWkw7b2xmL0/j01KEWFCgTIbe6oMcOWRzRmRu5
/Wpf4/IYaZobf3/aAiqrw7frI3qSMqC/NzAeQ3Zcqaefm86EYYki89RCFvanXgE1
MCoZ+mGrNgmPmvzOMNphV+sd0qcSfJyU08BKAdUjRxQTv4NJUvBgECphDW4cx7nw
K/VUicXMEeDJewyhP80mshFLHDghPVTr6JiQoewaImFq8hxUMGLMjlApLK4cFREZ
K9/Fh3SDtRTdL6vwSYzOiJGic2ilbYari4jpphhKmlXCcp8TbB4Pg5wusJf9uV6q
QSBOd3A3jPBMxRY/LZjGAsmMGEagBg2ijG40yU8FSMxJU2US09YAGyruWN3yPQa5
+GIgPgMUYOhSHcKtSoQmEeNLqZZ+bFR/f4/k9n64IHNhT4Bul5QsSEctLreUygPf
AEJqsUi8CsCDToRPgP/rZ9wi77aqZCl9JrgBOcyfY4uInv+i6jk0PXjqRUYdmopC
3dJkY5KP0GZafgIGMtP7W91a/besxku6kN2zhiTIwyyKid3pCMQpjekKj7gAaFF8
scvjJebioEkFwPY9dAxQmBR+7MKTxbn4tHa/MPNsGPwo7L+02E6V/Q6blzLviFNO
rd0O2VBiu1K6wAxMOuHZQ95EfSlIkDimty86I7R8o45zNPZ+ksZh3kMzl28vXF6P
SnQlAKIF4TuEvYybUFfESUFdrwdcdHYVvmnHOHAYl8tvykiCyyL7x7JrcXI/dPL/
duMlYX7NTKVJtn1xrvW2TfVGmGfDbg52n3OhBHEtuBpL0FB/Y1RYz328AyG28l26
v658n31VZ47btrp2BtOz77gRUUz11JFBWzdEy7bVKxd58RfnwlSK0sV80Aq3xEri
Qnz0lQ0pWGolqhCGbMZPDvmrxflrZFq5N1GB/ErQTyOI4i/dtIVKx3rHsol+AJE0
yHENmw75aDEa0gfNdChovgCoEx3lbVX7wFqKrxrFZ2fgR4HoPHuOcPEmRqjc0iRw
Xdr59dqF3BXwmGs+xJW8MUgS+P1vuFM4hf1FRh6HW9XIVWwfY1sxM3vaiPyO1IUc
0REIFXO62C4H57AW+vW2q51heTBsn6zO+I+rDYFOhR82mICgCJg4EPuDPqosz76j
4Nj2cC6wskk9p0bGNA5USj388fSFdsVwvTr9YHipSUfgQ9du2Ze3xhWXvqzqFbG2
0EJ8QuuaWzMX2SpTEQrO2jGkgYz0Y8sj/mNqyWdvvusqTHBSgJ2x4X21Vh5h/k+b
7QAmdnv7Nqpvr90d29LCpNXzWJSuiQ/8e74PM/F5TunEYmnfkZBLC8JTYQjrQvLK
5LmPVUmbaOGhYT18w89891Fq5ZTyucEIjEGhEmc074tdqQSaiLMLuf4jUpChF8Kb
tAf9iTKdLX+OcanEPji40WoPzvV7AchMLAoIeWyL8S51+CwFksZm2y4Izt67bGvD
W3XhhGJvyLzBHIqUphOp8RLQtLpq7/5doDd4Y3rOs9V10BzukPP/iCyYLt1X9SJM
yyVxVx8lGvkw5tfh8sb2VD0qiuW1UXfmbhWk8PqaUgYBh38ofGx4tSF9qtzSz6qG
9OjFJy6koEO389huHN9Tb2A57YQPyfOcXe8bpDHmbWLi1oQ6xw61Lyxv5baHQFGl
wuf27+wkX3zhLSu2f7tTkGwKg1EpvVF6eZqeCxhQUdMfzcFP+ow7yHYKeimQw2uF
KhrLi6NvUjd7T2i59j1E/E0Umcex5/N2P+DgXly/HdY5/oIKK+4GN3hN9YUVkl35
Om5xfF1C5CLKnAt6VvKvOGHZfsN38lDDyfX7RFPMivWZotLcvY8Ptx3inget5Nhm
3hG6BsP3LUqSc3A+4g+kuiLqz80ZAbpDSizNFt1GYzQn+TTwd5AhPWxWPg+7ojJR
8bBhX9bfxz7qW4CPY8hl2JRZhrbX3Uk6lrdWkzaKkofdCGvhERznTthzeX+Sfail
j99nGaasQh4gKMeHn2OO3fHjXFkZQN7SbIuhF4FlNOeyv20sGb3fgbZDWdpBkUfH
jVMIZdt3FK5X62TcgoATGI8MJf2Ia8qW+ib96NvXm9x8LFVufySKn1G2PH8r9KJh
Fhv5Ks4jhw0B8Db9Qb564j5umgInHo3ofd0fKkD+CEstHAVHyh7sOGGWPO9Xz5QH
MFX3a3FGzJpvK23W4QrjifZMkyYVTGVgJWj1fRBfi3k7uxG3qrtK6/HhIa3kkbUG
RY4YseEnrtGXfGXQfo4PLyCHU916XbatZnDsRMpGqgLDWD9/vLYkqbRnfzuS+7pX
AUluo6QrlUMw1D5iG1epXPLfmHVhhBH8/xZRtQ+zDPRrY2ZZrJypaw4pwLD8gcGB
L+ZWbslgo/TX4RvpMqYPF45g3jRXKEGO2aaml3Vu4iRvElH/ebElCavy+k4lq/Wl
M0K/MuatSQvsXxVzBS+TOtREmTS6zYk3WlViewM2AbnEvS0KBsqV72p1Hi3Rs+Et
hyFLCvLbbfERtQt9cvH+B/POPT4Z600kGo2SdfLPNt8ZkmSveSkYUJqJDNQqI1SS
3XM0Ps0fNomZaAlgSFcwtqrlLsEKjNiiYNc6K2wSEffo5uyZ9QDmYFoNcrFzzgc5
NL+EFEPYQT/Wxh4LP3/AQCMoRX5vEgHLjdiqAo/XI05bGmTvG7ADFugPp+BDsOBZ
mLVvd2TAS0Wrxqx5reHg9zrIJxgcPHdlTmykY3a9jkQ5hIU6kBOPX/HyeFW9g9ZA
UD+A9nHoDhU9sRe+Fakpgw60goQFQjbjWKZZUvZSAbLz+PQLmEpBFGoz098Ss+S2
OljCNttMTyRVl1ubsInhwHFM+HcJFVnG1Im3KI0sEBgAXpvELenVJhykSfj0Guw0
cai4/2c9DBjqOzd8Er257w7wv1AYXwNlUlxPdrzk0BvSLzzy6OdrM0GzWFpJ8gL1
fInV7AXgRsFw8MIIbENqVLujHEbnnLJ4jOlsLK9J40I722CWTfKY0NG2cdz62QJY
oHCLoi/3wEFD3SG0FKfX+5FPQcWu/4VlKwkn+SpNH/us0KjhWRNqneo9dIMYPPD4
//tWMAZAWqoXiFRHP4SBLdYS6Qzg98lZcIAKdb78w9IvlAQgZmDshQcldqQVPpc2
n1MVYPn4vvZvjBEyIKg8cISxAaaffUmL+RG0k7qu8Mear4j7m0L/gGF3SgsFA1Au
NEjamsXqE7XzoeMbpFLBYlRhWm7Q/fAc31VYf5F8owzQL74GMX2ioWc+hBrGvfIJ
I7AUK9p6zcf8ZjCD329j9M8TPeQsfHUt/2VFiQri3fW2CprX/ZYYp5TCJXeU20W+
88vVXQckzX15VfJyCe58axdUVCNDuDXNVWnUb1qslOfp5u40os7HWu38ojBFWTRH
h5PnoD6EUkgIYv+3p9lcIWs/W61jOCcKTm7Y5/A9aQt9RNmFnPIWbYWrhP199O8x
2oASPT0ABaeSmVtIZYP+Nk8qj/ZP+to3FpPmUdVW1XShscYcyquJO5KlojI7uIvb
9WA+fj7Sg4FW/1MFgIZkCRiesGya07f2Wvk2PWtTKdqmoy+8rA7FNq48T5tby2Zw
wa1Jw+eNcBiApvKuBD5NpsAF6mObRaq8mjXu4iA9pL65iEweEQ7ms3FG4jt9sZQ5
yPIU3YJ5z1CYQgGzSvzaaCZcwm6srFe75ST0cy6dHnG4bhpXIJGOfqZ4QJFBavY7
zhqD2Q3ngVx/l/M1W6nfCZ0T0o3tsC641F3D7ehs5/6afTlHiIQwpSvhZCjnZRRh
TPmv4Tft5lvQHhtVTguke4Rl9v4if/0T7IZDz77sYhct9YyniQBc5X7FUsipasE0
Qt14IPzSPkEaILPipAGDQxtFVpH8QE4YeXPovYGOvgYfwvhxZ+lPyE5cNfoGe6Nv
J2cuZSRDvfzBQGrPZ2yz3w5vVlPEorstGxHwlHZbsEOsh2jhaA6deWN81jfeaT95
PYR8DPosLjOpIZ/MxtA+zRa8YeXbl76uMeQqebylsgMyIV5V9hv+Y95jGbf49V78
2EetZQ4MJ/AGhn6vNucT8TdHinfF9QYjka6Q5Pbz/8Xquz6MGOke0vZRzlIDG5f5
wxI+XhctcldcbP1dnZO7Kz0g2RPW3uF/TN0NoyW57vs3ImclIwGVCCGpSBquViLx
8cFMwOyTyAorixyi8COmRJl0OLEmfJYDEVaMoibzAiVpXNy3VLXVJ6uSIMNFgRil
iuIIFzynfNwccKMwfOYOLHQmc378knNOBaCG6UgHEYyFYZQgakVQ7q0ENbQ6wRXe
ksGmj6xn1SNzQGI1Hgzk9LO3UNGiPIMnd/ku3hHNRNfpt7bY5u8NsWYzoesCNVh+
2SRUnfj0t6o/hNeVBklPYyMRg2kxQYV7VolpMK2IELG0/5tgYB/12Ws3u+q2n0mf
9R3VmAD0QtLq0NdCjdR9J2XHY9ACKazbz48sPdJ6o5KMcylkxUr8UMvky/5CPzNa
Dz+g6BhWW9t0klafrfzddkyTaxaIZjSxP7rPPRo1ZKP6985fs6ebOZE290L4+51M
lj+AnONHnvAgLRrwiHuY8luUOWV+ldgdyfYRwfbn0IOYFXFYlLJEc/l/n5Fv7XxA
vCgIXrwkOwvT9dluGFs7Qp+Ww6uiuiBnrLpjCbjDp5O0mHGYnKjIcPGfLxEDWIIG
hYZqvsExYTCC25YVjfIrtKvdAA/ONfgXa3eE8XPn040dB43BkpuXkbcntU1eCqeC
TJNXmP1a5FttfA+GB4ge01bYN8Ug9ZoxaM8CPBCM5Qcl/Hh6a26LgSFRoXqJP2S8
eJ/mwoEWZvpAte27LABRkZxypajxKWX3TFa6wG+ymvtWCVcsuRJpIW4fI7LRHqgP
YncY/NLVy/OOUd+SUyEZwL1iHGP9+2bItooyMWZ64bY=
`protect END_PROTECTED
