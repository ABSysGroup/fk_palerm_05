`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HlvvmihXYJ+SY6EmMEXkXfQqt0CQf9ti9Pa/blWzjqU1d1z33kzMEgmvl0UAbL8t
/dt/s6FKZTksiQIcxQ7rynF3FLz8tn+5dRXQD6vObSEeEnbsOn6WB8Bp4ZlQFlac
b5OyLRhs4cmBR4/SCC2oojrMluVJED5ivBO0KTMfOowXUOo0+FflFNZg/F8MUAdl
WTkHYXM/xNbA1AMWXhYxqPzacS0RMnY3GqflrlhFgDlRsWTbGYuF3LB6LnfShz7H
1iOHp9YfBPPCrJli1aVMhOZrEbPgG8eMHHOZLCmKuNegK3zOUutSC0d/cih+CMzs
XWw4KpaMQ8KFZZBUfJ6Oc8TFBkLVijG0BZo7G+31YUXgD/ZFdKAR6qwx+Svob0BB
gS/xgk7SxO8eFdHO6Vzo9q+RZO9TZtMUizUMrnW4W7zMedCOEp+nl3at7X4SqPtw
1YblzCJJhSgtzEA20JUu8gtTHhreEm2qW0Y6HGWgERowkXP8Ro+ii4L7w0OgUo+H
`protect END_PROTECTED
