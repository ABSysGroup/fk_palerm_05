`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E8BqVsMXFmCR4ejAgnvk1N89aTriiJ2ubLpeD3zRQllK9SmjfrUhzZgnZrmZW5/p
P2bK1VpE0tVm1KxUqIAgOQPy3Whs0aDrEVHaCFXCCHHERglmKIYHaoJ+0tzl5rzf
KQf4W8h3eBD9H3zqCPtGg1YWoaKAXq8LR4Y6I5U8P3SAtI7TJX9ppDkd67zizzxk
S0PmM0fQYhCeR89dyy/pJozo+LwCNYaD9RPXzkr++sa4NQKvEExGGsTyWOKkBJD7
GTFZv84CfM9x94sVrpAzoMbs1cVxNp4T+arQx9Ztk2eDqY/OvjqxVibOCa1E4aqB
nZcX82WYJ2fcngXLWTnfPLc7jTcJt2thiUzC4QCDKb++t+VXEarKH8kn9lEzYmJg
u430MU/abHxDKo6jt57gAq3PaWggK2YvbFdKRqgOhtlu1bVl9yjjYd2UTbfbWVzl
6xy23BHCoXgtzmrAFPSOia/yCcwhIYWjTERqISot9mascF//G3z62AuIa6/LkFsH
Pf472HzIoyiMNJ4Yen/Nmiji6/tLeMOyTyZUzYuQ97U6M+aJGXYttJd316IjLrxi
93FT91StqjTepZ2tyZVc4qpAXTgo213NgPHE46ND8k6UuYwgiN7JP023H9xTfIK+
IxwHybJqgJsQ2aVM/gGGbZ6azrw5MHkouZgiDflmweVeUYZMyzhcRi5PexslcT4t
fVwT4XCzW9BglmZY8ckOR2LbYp80jw1qqsXLEzIMbielz9A24a30uUKoJ+rWIMjP
1R24nm4hAWCixcgxB0eKX40Ccn8Xplit4aoCaVKa3kupld+wQoIDLN44G4g4vCXe
ZrutZJAdPu7pnAw5J5x25JSdDrgc25gC5AvRHHNHVFKgk0fiV0hKAfXz73b4c3g/
+S9a6tzhoG4dSC/KheBfs9DUcDql7LZn7RbRM2xyQK3aSSoi9I8iFzV55vvd8LpA
pEGsz7+4OW9AH7HicsG9Z07awxInepPvwJQk3fynfQtdJJ8NyowvKojy52NTJZvI
rZi/QFf2d28LxeD3eB/gSu8+++oFDE0UEKX6lYKt3mtC0R8/1N7P3BKbkpPRvqrk
c3LHIv4+tDdPvCv3jFwnqmQc1wsqkZjrLNdYdqA/atQ0rZUTMUpT4LMeQiu8rki2
mimGkya/IXstoYsiQ5EI0coQ51YBlWLmHZiIq4InAouucXsNXYWZ1mC2kAmeGQUf
3eFofFDQ+LtvIM71afO63V/pWfRYtyJFLnLtKt56qzyXAOLOcPle/b4e3nN51t9s
JZCmycIdE6JkVUA/0heJqdfDcw7u8mxr06XUyxweBZEPe0Yt2UgL4aKzjXfOFiUE
k9MfsSSDlKyC12JYVS51pQD7sOHQXmfqtHHq3n7XAL0Jdx1moUyD3Ufqc1fC2Oz3
PLRGflfE62n6Qb5BMOeKkRfu3hwmAB7uHFY3NM0QO3KmhgJkqNJL5eRNWiVk+Ak1
yQkMiiraU5bcrT6dt366zg==
`protect END_PROTECTED
