`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IV8htAqN5jHlDNoPm+5hjKM8VcGvHDpbBUamQvkCoFVZAX7+Jfb7LcvjpaPlkL5x
ooDTCq2srv2wLxmS+sH09XjOWUxpNC2EfA9LE6R18TX7K+ePsGa95yxYLWJ4TGNx
2dcYS0ixQKIe2/WmoqD77Z716C9DOVGhWUtAx7EsAyqaPBGEhMIicwvp3prAG4jM
TAXfR/byBX8Iot3ROnzHf9QI3Rv1Q/TsgxEONQ43K8J96ic/7vLJeX0PzWIPzP2x
jM7oeWfy1NRzsD8WIIec2FFSnF6/LGq1XefSSuKsmiU0PMFL1H/XUEVjDN5VKYqb
Po++Bov/e6SbsGAMB2WZWiKpRukK1t+P/xtayuGGoNNfmYZPLrR9PKuCVrNVNInl
`protect END_PROTECTED
