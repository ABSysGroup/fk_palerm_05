`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vcJT+9uWG79smtn6Yik9wWnk6cWPX9BdqhuBrwUvT2sXTi9T3WctXe42k9AyPHUJ
eyj1AI8p3ytrurbynmVQB4F/AqbxfZ76RiSWrxKZw0oy3YRsy5vGG7QgT5ATihk1
t4maINYOv+QkiNYqcWl7L0BpBFhTqDXD2w0kFB2MTf5ObjxV3sifDiy8OB36GyCs
yEMpzm4OfJWIHGlbut7alWC4+e/B4UxWv/BgEVoiPZrmMmahfLly4jiMI84vihfI
JAokH6rZ+5KeL57PGfGr4Sq/ZlKzWZHFYVs2pJKmQBwNyujtRzCdUWTE3K8s26VQ
+XwApzz50S/xrGvXcMpKA8o4ynIxlQzkQw8S6tz4g2dqVjwNm6GtK1xl9oPFRns0
MseAla5jNm8wiWwgOUQIlOCjbHpsiGA3zao+E96lS4Zb3EZ/hwH1nhj6to74k170
8In6PnvWhCpjv4MLjOvlvixtMr1Uy+YIwIluotU/F5CfZ47rO2yDNbLaQamvKn3V
pgc0pH3+VOdwfrwtfCMZFR8KgADB5gfDjxEpQGZbYjyuU4SyzypRFy5Duex8ZdiX
hc+LWRWlbduQLKPTk5kHIIZfELOHBuWkYtWRdPQrRhQsLdFTjn3P/DzDj22acDzN
V9pkH4l2wtNeXAcqLtC2Autgz+Xel1lZmjK/R5fRC6YWUk2pSWWQTH2Swm1w9yNM
wVeRJKeLiPsL8mM9PeWM7460GFPZC+QOXzFR9nTeSH0UZjVqT2EGAI6b+DQFDCME
B+dBiA+zQb7MRPQqj4w4W71CV1BADc7JHCkeBfkrD/p2AMpx7zGGTasFX74UnFAm
j6E50E55AQJlSjhV18cqCQQSxQuod83bOkQWHb+Qp5zCfFQjA9dg+NaE4tNrPp2C
7jOUWWQ5rSDEYmKG5QFfsQ==
`protect END_PROTECTED
