`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GngCAxmNgxqwXRbNR0Mcc47ddBaEFB+WGfH6DF4PAx+e9nP4pDEUCcZHAHOjpBey
hSXTmTv2l9rZLjbWWGCGyjY27WDAqrVnIrkKcWeDSG7I382g07m+waxufGYbVHxQ
+8y6miRAHv9d6EDIpdhH13pfh0pNoZdECB3vrsQQvm+EJQOWNDxtEDkv9WEFz+8e
gABuYfiD5baZ3NeYDy5rtmsLYmcoAuZDpW3kKNvSdFTvMFfYT5RXTENYt9eUYMQs
i4Kq0XeRidoJ85GVwKDbNfLv8xNdSjSG2Y+ODnnyR/PE7fpw2k/1uQgOgzyMr2fm
ydhcza9WHdeDoo59bqBuy1PRXZ2yk3kiIvRMXXzFtJvFKa+1lJ9CaZhBuN6bFFxT
utTUidh1AcCTDIMDGIfgEA==
`protect END_PROTECTED
