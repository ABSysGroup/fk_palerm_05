`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W1A1ze9RBKGYlojpJeE8CV/AhL2ffE8AMyLxQbbSBqL2Q9xc1sZHMZZrrFZfoB+G
dKWJHqOnoJsiuETJ1wyedzDeKVVT+bKeX0It5vPN75rFh6fj9UBftts++k5fQWBj
6REnvwGqT0xnf9oNSKwyV/BGpTKXqH6eJMuBVPfBoDsCwhkc1DUghNo1yRc/V0Jp
yAbg1xajeppcwR7XDisrjAwPsdzXzXNP5i66JDYU9gmRPWPROV5o5uJwm/xpSUXk
c/NgT6FeFfU8YWkJSQojmw==
`protect END_PROTECTED
