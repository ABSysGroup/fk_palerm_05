`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OEBs+L+0on0hof01a+Z0e87WzCEGXRsY9NNkSpi3Cv/jEd6dI42Dv0Ft+oRuv+s4
kF4SnTUZxYtj+LZubJ03DQONzr0Q9GAKrJLW3c4lVo75aWCVqoQDXpUd9ee5SKFa
/nI/rMzmEEZefhEr64ys72B2i3JpJmSwoRTbnwFBW1sNSeyutpb8TXtpXWrGelPK
zYaEbsoMkUp1gdHayiSIg2u3jzMotjkjO7Fvlvmgpl5nx2Lllz/p4QujyDkEKWWW
BmgzFfQdFZWboHEFCxYAyR52gvinCBpATyPgrEIkWFiLyYW5tI9OEx+uQlHjoE1/
flLDsoTWz3p9vFvjnP0njeMO8qwJjrzcc2NDD0BFibko/OQ/4BlnHt2+ytOCUinF
M3A8qcvzS4peNz7dtvoE+LTiVWi7NpngbG0uX/s7nb8=
`protect END_PROTECTED
