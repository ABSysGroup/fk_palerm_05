`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T9ei93BwrRQmaKQnSaN+n+emr9Vp7lsnP/H3RjNr5c9EglOFbcfg09IDWF2psMeI
5uvcLlZFHMUXfGwvfUYtVXgOdCk5XOyzF5oTwgfZGJmKhwmsKAJ1jjcnwnri2hvW
m2TgnMnyMePMsPDSU58mDegdNNgmgoaOnCyKRMqwcPDivbKneEzhCMugqOm+HbtG
keASly+HEX18fBZbj6U/i9mL1ApohDtdUHJUS9i88hXT8cUCoOIhg9fckbKhiF9a
2QmfUWI8HnSyRfRCbLWcL/r+eHEnw2pWfdYwdByCOLceLTZTom/vEdg4rqua3zv1
+wpYMfZK7JBCzUFppgLt1x3tiZN+6pfpI5mwJ7dR7tHSkj2+9S73gpj6dVpLGhVM
g+ZOdzVwALBOiJ20OljEKyVTXalWLvgSm4XJ8Dcx21UGfM+JxV1goVdV+xRNWbh8
jZ78CwYMVIURLRSEPMLEv7nBp39GfpsXLncoE428K0wS/Y2+rZUZW3KP+yZr2EEp
MVz4G0fMTHCFw77kUq8/lMySt09xGchj0ibTjXWO3RmbG1aH6CL6ZO/D4oqKZH/N
4grdFsBWXwceYud+FCJyfQ5J/cYjnjN/Aqq+jjsbSQ3cKjjj9Opa0gL+0JLt9b7B
PDAMMpNRR+Fjxj9GovShn4OoBbQ4/4PlcBb+1kQ5iw+DMya5C8q/1l6eLUnP2IvZ
smdZNvBYBTKWFU6jPwjj1o15sS+CZcsXj2Al8jMf3HO/Ny/Jv5g/HrfoeZGkBYjk
irSIMQ8aiVicAul/N39Y7fiL0YWDkXiGi1xpFfqIP4qIzVWfJurauZbm+65hkAu1
kyOYF5DU/hPaTIqv3YrhBwvqtxm7pwtPmM63Irr4YTzNXpp1zHvhSb41xj+6X1XU
XdUDmvF9r5wkmKUdL11uUkKRb4IY/wKtsltth+DE71Rusm51kfk8Ij9MDWvq5xg9
Ku9kcwEtbkDSJBOoOgg9hXz/W6jsLXLgPAmHp+Dfwq7lT8zQSfHr0HSNNMsr3z52
u/onJ7OiP5e2DQy1ucQNeQkgDsilBwZuS2Pl58u9KIfPEaUVoDpCdfRwBkhx2ynR
4YtTONxs7R+KW1XpoViA2cvxQ6EgUlJQiivSsDOd1CUoWfKLmttDxkrIUtEJhZtp
iPD+kxucedV6mBEP/xWfiZD9zrFVFKvTCWOHsQZt7LOI6IvMud9pZDLer/Cv4yh5
J4d7ybd2Y0R9/XRRIhikz+fp7j5nqaaMSHFRsxrIUlCITZdAB/QpLXn9q6sSS+cC
Oiskp+Ox1z471JP05nrheEij7+gaEeNJXXjN/eqAUCXfIn2D7ChKsBkTS4hQh2+o
IcAWkhSpCM5aLKfgTuzBIq9fjGpUA3yFKU+k/0qH7E+1IL7StIjeTjsvIgB1Ugae
sqPv9pX/XVnZ6dHMdHD4bvOhwKYYd6ROZKuZ+tPY3P8bNSZ+CkLQwkFMwnshzE10
V24q/y8MCUDZ8QesRa6dZb7xFk7AYT3VfxUVRhRaYdVnYSFGJQ3bP0RmHm+zKUBr
YS5DtwESoPa69BJIQUY9G2D5EZBeL5XMgGkrpKKwV1ufiEVkwWM7I46NPPgeUavF
RE2RLBh/Nab3etsr0lymIgqokzzFSVrZSLFmvLiFNFJey4VaCfMlwpBNpSPVrMFX
a0SJ9rDXUGWzzZ0RbCbusxu2WqdcCDEjSh6Ui/CPcA3Gsj9JWq3/NRSZVWxXTRkd
`protect END_PROTECTED
