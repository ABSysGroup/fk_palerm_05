`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GGjZ4Q4it4ixshjqgtUKwvTYHZvdWeGJn5PrReNl50hbG4G0vNLaBudqwdB5S/S0
s92Pk0DQPrGAYDdiGcV3wD0tGuVXyj6FUlxQA+bBV/MbTSN6DlhXgF0B2FoNwZCd
0w08YjYLpvuocMFYNV0JrSd6W4/My/4jm4+bqSclB+eXb6iQT8wYUuoyDb9z3zpp
lCsRuIj5vzA62YEt76ZQSo7Et4V4IEoiqLR5f10AY5qVk1q1DkUV2yqlIqzwa7iK
8U+HENFLo5fYnWVsHraIEGKXCQI52pbdhX5FZxRw5GQpKwmncx1cfq62fBXRkX5p
30w3gzuISiRz2hW8PAxVgZSpwjI0weiGws1I017huyAkUuSSTDloAnH0a6iseObg
AYZW7h89UrLqYzat/2svEQ==
`protect END_PROTECTED
