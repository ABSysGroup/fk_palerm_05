`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
blKaIf5tBP57tyC+FmruIEePRWQsFcXev2TkA6G8UxpQvrJncEgmyMWmEKT8RaoL
JBtuqV3kjCVPaRRCH+30NJgitbz1p85w/PCj4l6AeNuVSK1cvzQPdDcr/8cjFQwv
46epBksUhv2LJg+5wEC34XBa/zl52+PFIM6DlNUedh7Yn8W/CpI2vajdKLBVvhOT
cR1c+vsegmtXKmnaZSNr0qx300NX3rrRr7Gd+cPrlKnVAhJHy4RsttyNcW8S20nQ
tl4GJ2unc6Imk2a1B5+uxFPZGj4XJU2yBgwk9Obo52IuPNle8zIfn/b5663x/MB5
4L0B0mG04KIwG94Ss9yyf23k3QYHkKA/vg7HQGsSngXqfa5/jt2jPl3nqr8JAU09
cCb4WE/XKgoXrp+S0qH09SbFVUtT5JNGpm3/jx/Wh80Z5BrpBeRBZTWcnK2I9y+T
9C+VJFtvthVUqbsV3M6OM4WiJJ87wmIPlQ+Oam26cROfLQST19tnHK3f0YwobtU7
S0K72THadlGp0HTUkCpoivMVZxP9AVfGx0BP3S0T3TCj2mRopBCjy65wE3Nh3And
o0SvA73kqxCznDHvJI69rnQC1CA84ZC5+7GIo812u5Q2ja9eO/3I20YuW/aob72q
MrZ/omgw1Y9jZYcfT8tofA9RqikmDt9RWqqhy1KG0EinL8haLuGKA/b9+nl2yN6h
h3+UT6Zi1tOJ+0PxVFoHDZz4Otu5GrfN2oEtcIvrX4q//TQpot2omS47/O8xafeI
a2L2/MlsklXns9/qxf1+u+1JIxHirPRH9AHmsBrhyhydkDE87jOAMLPpGPBAHD8F
iLHbe83wUDwqcStfH6jI2YdOXprmLfKBl72Q3drAzs8bm9RWP2sTtQFCNxHy+yIR
elPSwz0t10LPzRz+893o50xx2gRCsSoNCTTupJBs9gim1Z6gpHVseavE09QLpr9z
ZNjCMFJPD2bef6eGHhce+IcajEcLezXgDkVhsvaqgSacl94Fc974paGFUtJUz8hF
kKn6qo/otHmfGAlS+gzrHgB/BIyu6IfTjxY17kgqwd7IQs3IYZLS7IKQRKNcxkKJ
azQOYvTcJjqTJf/Q5OdZcxy7f1cXFw2e0nD0W5rXFLk4YE1eNPgU0LQUyewGvXmX
YIituwDTX4B8tYuGKbjLzSvBROyeckWSRWafTWaSNbexchYTbldRlvKjfXjRGK7g
Aq2ZWtM394LpdFTaJ3Fl2gS7EV2/4Sgk4rgZ/FeZ/bWGPgXvw8bwrEvSSey3pZKp
THndBaSZZ4Ppb+zXMEq5Kb4iXlLKKZdljJp0ANVcFEsQGYXusssA8xafAfFsQxYn
oBqQXlskmqgcShSNukey2TVNcXSnVHT37IbufED78DSFW7vNHcLn77wAk8W8GK55
7aVCfmIcqnS7MnigZK2SNBvu6UaLZ6iayAyslPWt613mAkWs/S77Wth3bQflcos3
tfyn8yFYQTw9MMbUcdx9PAm1opTSZbKOKzFmvPrvN4gaTho6fDz6K3179b+kYKUf
vml7yxTAbBwPJpi7IOtj93uZMOmhl7ONyFA5vwmVrx5p2BAMAbuACO/ZQcEImtSY
oUfr0tId6XV+PYGePfwReL8LVxNqNqEZ/HR4hfph99ySZvVv14xYBHU6EQRyj2us
5WzGVPUv+AVJhEu9B73i9K2EIAc7C0DPX6LcZYwUxl1Y10ptq2U70HM6st2ETstj
oQVEbJuw1zlqCZpQM1pEbQI99uxI8A9J2PBvAUc6oumaCEO12kh0inMRyf0SNJ6E
zXLrXPyAIoHfm7k6kRxOsA7mbOBR0KbiUNr7JAwm+Fy8djqgDXWzCCW3gHCVubQ5
9kSVTaq5Gp7uKko/z5zCmaOeVn7FwfnE508z1Of8dAkBtRMMYjM1D1pQe4J+s+eR
O0iawy0qV6/nDoqVAmmL1s8PLsis/NQV2MJnzoZ8sbsqJTVT85gxwzoMG0QXR7GT
+fiHUbLoeKGixPkY/8D1Ega5cxz0LYfuEvnlnpcR+3NpHUUTNtCs+6hEreL7Z0yL
e74aJkFJyg+2vW0Y2C65Tp4uMFOkPjuitPW8AMCWd25Kq0vIT51SB3+xqQXtVHpd
VLT/ZEuaSxQrQvg+jbicU+ZDR4/WtYsLG9XnHh3ECKc3MQunH92ayNkCRILhr3Nl
zTRDdqeGoKSZ/rGPtE1bHqG6tlum2JHkr2Ofk6eqgpjYW1UsDfzPdkJUPPJPUsuX
Oq0KpC/N+YrV/NH5et95FRA9FgrjK4/bOTfe6MmU98BDzK+Z7pUnZa5UK4dGGYoe
4EovK9hnB+GynHtSjMVrzzmC8AnKgOXIfVsa0aulw2WOHFlC7bCfpNZLz7amhneH
kfuVpBBL/uk2HKkTfw6B+/Pl5B9FDV91lHoqOyqVgIkFrw3wqA6ez84Fl8ApT6zb
hK2F5THHpkg/7or3xmVp0wzEuA1XBZJvlqrjoEFuJRosf+KY66caI7c6S/o99VqL
TH3cAEiIF4MSw/xss55IvuSH9DnxTPyejoUSQB9lLWKwqU8C1UfQORMB+PTPg+Uh
OW2tcQyiIH/EPtl/huLNtAnIGHX1OSqB+cCtpkG2znN7ZhOFkWJjK8J7HD/E/vf/
LEVeX7E/yVu5UiHFZUpFB1R3de8y88j0VtSvxz8aULQwPg6ejZNEgm6eok2OXDHx
zAU6QDoUnxYSBrH3MCmlAyvU4IoBqHhaKTQb3mNDA5/OfX3LvgMqD+KfMA+MWoQd
`protect END_PROTECTED
