`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k63TOGPOhhnb6oLwur2lI48cZPmBdIohCqLPr/t5BxlaE4UE1bhrS41UkCXlMODL
eptc59ph/BgB34k5DTvT/f3pazpEl1E4nRiKBxIWSKQwxuWNDlmOaTAaZDaAKxeG
jURwiKP9VgQcdwDFy+XWVaralFlSN3jesrrt3DpNd3itEgfHF1c2oltGO5FNoukG
Mhg0qDzxI9+eaEsHsvxT27dtZWbmf96zdbkWKDvfN2kshgO+GEdcP/p8qyfLQmeu
1/sD+NIs/e/FmGtwrEpH8QYf/bR5dyGzkRA5h8F0PsTC2lxU6UzghO6Xz4XPEjRE
Azs06G6F/Sx/Y2q7k5j1+JszYT2iHszjtKeJXkxPtDmJDcIa3Zmw+Nqe3Omm8Bt0
FA6mHlLp1tfoKx3c6XuiUQnd4IQkVwRbTteqKeaOW4A=
`protect END_PROTECTED
