`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fTjho/sO9KxO4we/mmzAQ5gsxKxGeUpE+R7ca2ITi7AxqZMXA/ZVPG59EQr4o2hH
ADfeksekD/b3KeMa9cWOvxHyLpyhlSpeOuGubyp6RELJDt2Hm39MSRNGnFq9IQbx
8Q604oAkXRxiyIaJ32IIl4QmfzmnnBpQf/4CJQ2EpLu0L9k4EqiYn+GXTD9kmc1+
9K8kqxGVsTv8HEnlYCMrmDu4F7QTI09lCK3QHY7JwUllL7OeR9cp7Uq/NGvucjZQ
uGXYWOS0bHWNjyYjJ6wiFTuPyl5xGz15HcJtWPevvr+8ff7shD2BAZp0Tx1NmrMH
bj4TiQZhBRn1dbC7c9fSTCIfByB1WQ2V9chZcccYnH4MADQqIQ19ZlAkeRECUXc9
z7KilehUA+tkNt0i1BvtIRXVzdrnzMsvGwTRtJYplI8oSZTxMePrO5L5R5eoBCLg
CnYy3PDuA7AW9Xxpkf2xxjuocAKBFlOy2084dqiql9CaAikCe69UDgqahLm240XF
HWuK+Ll/b8ZF0wK97UMhUGqIYjvdI3cAVgmZumMbFkioz4NimjiAOGJQ8ofyvINQ
Ta/DbTfM9scXVLy5HV1kvBlTwGIRjYSpsnNLH9ukvvYK4ZGRQfmCAipMzISX8gYt
3JKt75n0PDdhwb2vwSg3eA==
`protect END_PROTECTED
