`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5tw/hZdWFmR9GKlFnyQqe10Ofcc7PcH+U4W9wnI72iAKlEp0XI6Z6aS1/C4fCGzp
fS5j28pjOyxztpt2BR1ICHUlZmzb3mLUY/3D68D5To+S/SBQpfbkMaAmsOaWd0vx
N6IVy+D+m0rOqpTDXyE28UjSnG7zl2UJ+7ivNT3WK2AK7Y07Oe0p2gclA3qTfAf5
BwDoMAVn4FwTTC0fdd+JgkFL0SFUaJmToqp+CtGeBobUPI2hHPo5H71KZQXpyiYj
sXuviDFtjgRj0ZMejcyYWQGdzYKiOwEJ6cVzRXMvUDAAOqAt1ORp0yI9g+d4lfk1
tM17+x35BObjcEapmipFsgyLiHgQCk/B+tZTbY957YR/LrYySvZW2YR00ssDdUxo
lxgCETJyfEbj4rt4JgFQfKRnQsQiu4yeXFcTaBGNlMCf5GOz02u4oH2fSlO/Mh3z
iJpbxrvofbjujkXa+W7GQLq/hwGv0M6ZtTW/LhsvnXyh8KtEyI3ZnkiBoyP0PcDh
yTf07P7nO5Np0OKhcGI8gsGR/30iLTSESAB30ZBnm6805pcc7kj5C4j0l/g5S2fX
M7yYDO5ucigwUA1uMsAm0tkB2pWY7coVJu1SJHPAqdtO4Tv3e7woYiWu/NM0W58E
xXcMcPR5lnrdhC2LN8iTsm/2StxjlDWUmF/ycLdMLBZB6RgVmYigdYTfGFBWsWuo
BGEigz3fPKNukm3D+EvwSUC8ZlCCDSfIvUQiPLxIpjfj/ib1adYGe7Kl56669KfN
JNhbAnhr/7qKSG4tKFc/JV1MQJt4lfzBVlFWpsvuWV+7cteikyxqlMi23BQEEAc4
03TlmhG5nrDJN9Qmape4Rpb/8Kr03uE01B/0COwmMVb+fPYXlRPBTYH+Nfz7XJzq
Oa3kbUvMNNlZbuBAwRzOqRTw0OsjEyNrMB5EgFMoOfm8OU+DIQqBE5XcfD34yql8
gSEZ8snGrvODgIi0RUGL/PmRvaigL+ADftxmt3bPczlS+d1CY556vZabFJg5Z6CN
+3BX8JOa7LpELYw3MCdS0lSi1R1nkFN5HIvahJWhCvwNzhTQrEjgFvh/SYNoyIN/
5zgL/vNU3xEa29yeZpeATXeE8vcoGcSxaV9nPYFSQBh2Ba8ln3Df0kee06DGiW+g
ssc0shimWJc8fmPLogGDI+k9VCrziJtWHZ6zDG1VcmQ7UvvAu46+uKWSWiXAdX5R
45vi5cp5Dr0TgAPH+X+KVgEeNOjw1mX8LhF7iqYpARNyP4EZcXV2033Kw62dc0Wr
9UybZYQG7HS9MbqQTdmp/XzX7llcs4Vwh9s0sFXsPNObZnzIf62SfWgyonujXsGV
Qc5TqYTsizE+0b23Q5IKDMkQnDVpedBjlW5Qbdr2Ps1K+szb2YiUXUNzqeHwN32Q
nyLdMwM6edK8gTWck8zAO9h23tHK/e0gYw+R94wFWju20JxHIU97Or54kdunR6GS
um7oBWRepCFXgRTRgeOVApvOgDjjFMnsd1GaasfhPyFXr09FJyO2vHWTOquMG5k7
yyj0b6J+vPQxCKlFd2qjxoeLkT+I4UWUHygIBkJ+gtN4uv/azW8tzv6lm0fsMrDj
WLyWDugRrC7liLwD/5m3WBTJHc8+ADfHe+8sMZh60/3ZkoiXbdveichbWVprywEq
fL4/X1MBYFTMLcEHBVVpuqHPyzIOqnyqhJUimpHLBZdX1SM84DrPVskpEK2ct6ia
le4NftqnwuJTLyDjhArwXZ16qnrI2KyUnpVS2Q4KB9fgPeta0CNd2nT2w8ML08re
aiVc/k6IZDQHX+J/sNr+BrVUXFjWkz0rfoZ8ifKVh4vF7AeRAIhBcSRDXvuTCvk9
Xaw4jkADWxYrmw4LVMJI4faxRe8S5FjS5VUCFKN9U1CYrislPcz0FwmHVhzRDkLY
JBqxoDrpZ19ulYcDIUmatfXUCZCcrYatgpTbigZR2HvL9AX/DYtEhkrqDzoVGhCb
rikCsED8k7yr2zRQxjLRe6YeU+AMDwaY1Q5DvYpkcS1jkfrJSszHX+3Ifk12ujik
ZbOsVFS2RLFSaJqRrDGgGKDgzMKSXXThC/31/GtHnpfOe847muL0gpZESTPuvaXn
mef+wHNOVE23f/sNmIbivauhmltCjz8sVRM8KFaZo4+80GSD8fOYZYltO6/AAPBs
pRy41Xwwb999s0gl27ja0Im0excrWHXgHn7x7ghw3zj7AD5evAKD3/8nNrLGSSBW
deqLaGDu+kh3cK5SHhvV+4ZQoJu73x3ssM0Sse5UxW8Iar+UGsevqHr8mbZvSv+4
mN/NpPfFf/TA3Hq4ctfID/uW/2xKW1DSqYms+X7uXaz+4mGgERQRqgQXQpZNXfnZ
romsQ29FVgCHPiOiutdIwR5fPmspl9Im0HR04GX3Jw9pCnNZ0Ll2fBVfmQfnibpl
C0h/ndUhHxK3ViDahAFvEl43eLB255XNjW0K5w6Py2OQGFcsj6SPzW450kwt6Vmm
6Mucoci0ia7N2+XJAs3JUGwUaQHdHd9ADdBZWlopyPwZXGR/eAS3zMbpBc19sR8K
koV6W7js/elFBL+biBPIZaM9YnI6JCUs5BdOyOp4ivGYR6fXaQUemrHVha1oFojx
YPSafqE4c7RuqzW3/Ww0IqUCc8UD0lGld4Xm5vx7vaPPeACgNR6qCv1bWGTki8Yt
Uf/kX1J0yaRYmxjitkib4Nr7WULb5x7aQliIWTUXN94weRCnH4uUyVv/oPuFVdVl
lVvW07d9LdQ52rszVvSndUbPuOsNQDmkvGGjNYtjNZ3p6dzugbR4Wfv5A1r1q8vQ
Uxr1ODCYIlS9r32BsokgbmYoUx/uFA3oyxuxWKgTl0t9KFi36KinPvzHuasQ8oDZ
TQkKZqoRooyzi/PHHx8Ki/UPCD5ooPEL7Myqn9YOALYQZLZqRag7T1ePDdiM5k/w
F2VzSjryhuwVF6dd0nCCbbWPmaKtMdL9/6GLGCx2xDHZ3T2pUUk8Sd0Tc39z782B
ckWhSKgazImP8JFlJNYnFuj76oxs2A2QvajJDDt4lbZmdGqc1BM69CV03umL/6pd
Z8qvalqu7aTD3/IMgZYhTPK/5gF6O0jkW66advIm5tBnK/anP9D0JlEeLQyEqOqM
5kVWm7QbT0qPwOIoD0uN8UUxsFAr33OBP07aGdHc5r0rc+2+N5Rz9DqStL2cD/LO
DOgbFSgXb4xqWsWBJClasXUkmnodH2Chb9Lp1kQN45JPFe9DRNjE3UuI3lHD7tST
ZBIFk5eSDYmYEa23zKITthKTkD4MWShKTg4NTry4XW2Pp9zHBEC7FT/y05k6e012
zTLyhw/XUFkWaFKdX6yidiLeZJ5wS2c1p8oiSaJ3KGRybSztJh82kWYZcYZRXewW
qUQLS5LuqjVJ4aBFgtvurZwyg9r/2x9NlihWRiNDxdI2h7EusCGSdFwvNsuTroXH
xVFgTNK8+giHI8Hp+kcv1yP4n5icRCIPQPXOBfBQYwJ6NCtIm4UNIPj24OOG2Pen
srMJO74gE1aoN4+aL8ZJipjkEb9NRdfCttA2GgkTP2u5aFsfiKB1a+n5YSOAVuAH
zn94SX+mC//MzrkmLXPopUrv8y7eARrH/NRqzQjKBY5Dees9FD1P4HMzYeuaiVZM
c1BPnjh5q9uUM/ObSmMTpYxYfXGAr5Hc71G29qAuUeqJJ9LKM+GeDFX91wdoU4Cs
`protect END_PROTECTED
