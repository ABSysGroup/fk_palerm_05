`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
79UyiCaAkzql9LDQ/txbVtLbaY3cmkm6QHVOqx9rKY6MAO9UKAzy8Jr8BpTtmIzf
d5Lbt/NZ8UFMKEox2ucGQxmptqI+SPVjrEFpHzoDL5PDOxpFwtW4QuJdVxwwaF3d
U6wV5DE3zVYxbMgyIJHLRFpBUzOdr0yTOfkyDh6i+7G2cjiMfGgxU3f1ki8exUBy
eE0wHjsS25IsUwr44nKjlIQWAzn7FNhoMua/+3NRMohTh+u/tpsMyhFBwCDgVFHM
3LuB2ACDtj/nLCCFI2bEeIIe3ZqCpw/aYqyjqVNGd3DEyKZ/pqo44FD6HA72cq86
ZQsGCzoFbgWnNz1El4E6+b99R1eDx3UOtfyjM36glSn48bsN9Jw+yiLSQbKU6amJ
`protect END_PROTECTED
