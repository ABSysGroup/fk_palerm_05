`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DAspgjm4wlEXXHNQeoFixcgSCsVO6ejXOFPE2aI6WVCd+c3BI+YzoFjAxxJKX7eX
rJrDAhxocGdaYD4LFuFqVz0eVFthaTRBRqBSCDIz2cqIBWIxqLfRc+1KscN82A9v
h4fkxrmagzYqUNPqlGalfTGZ7PQu+niaFnnbd1pV1UezJy0dm0WgZkgsQy0Cn07Q
WI/Hh3Ru2yo4Wb+0GtJVwo2MQ2UxzT8gplxhRqW+UPl5GNxf4vc7k2PgZb7fVnaU
muEiuSocYNdiDKjaGIL0kbHT6HOjfCsmlxcdSB7dyf3TqxCZWZdHMfxtyaoZxSYS
qAVzn/nNKYwz9cG6Lrp81ZvciurbEwU6TCpe6WAMhlXBSiDRUnw9JO0cj/6+vYTW
RUTGaSktQ4yX3PmZiMYZesSWyx+Rp4aF0bih4shcwNXT/r5+oYdPf1aemWbUWjwi
Vb7xfNy0tD+0dRPo4E4uBWBFTo8+1+NAG8SyF46zA+zryrl7NJJN6ZCHOPwWVZOm
pBTJ9g8IgY2ePuv51cW+33TtoNqOV++cSRzaOhztSKeG6BDzDeUGKkmy+3HTo1Vc
fEL+3fud64/Dz2qvs0oLtxB5VzhtMNv5w45ch4q7z2K9W3dkfXszvqxaoZi1rx5E
YaZxMObJzTMeYOqyxAZx366oY34aaHIprrgNYwvKwULr1kbI1w8efmHwQnzbMCNT
cxsVVHfpRQjphYYYrH+tlIZFQJ6t/+iisCeKuR0MleIfjtgjZT3Z4Xj8Sn979Z8S
zlaXLpADvfnKwiOwFH3QQPsK+fUMxwd8iFVzjcQu7hgUXT/0rI2YHzYzp1M92+K6
QmyyJyPSWJ1TeLmYrO4mHFzw5WIsfiQDp5QljjYkYrduKaAly7043lw0GPE/B18F
CFbXph5BH7MGBcr4ho4wPJWwhfYVM6u7z4QmP1BDkOSjCBLNblDfn51NH50m3mpb
OIIcEBTI1Za9AR/xJ3OjiF6w3ZswteMR/fn1TMedgHrGPU6neeJZv7g70TMsVguu
jwqzxN0PA38m2TxR8lEAwuQ+7PQXZ4/sw1DJmE270/CyGgmhtfj/fSY3HOWe2Fh8
pDDewwbVkWF20js92Y5f3F8SO7s5+Iea26gQsoAlA1F2XYdMt4/gH8S+5ax4WLah
lPpB7/cH/1DshIDxdV1K7+o1noSMGDha2mT6v0wLTmTl+DeAFg8yBy/F9va0h6aR
RI/lpp1b6Iz7zt4Zu4cd+kAIVw43L4rzrjinzdDdwiNXV7Rxf8J3AHjXf5g0LI9Q
5vJpSOIvYUIJrN41C2MwD2PLqPgvu4iUqIBD/oawr9C8IQ4KigYiJJCXHVS8/Wmz
559wD1F1JnntUzAtEsZ3IxnU8ZNY4pmVuGpRz3A3ttR4NQ2Fwk7wRz/b0OTrIDLE
+ihPt7UAUnBTvkFGt1ogxf7USMRgCSTp1QG4a2U1EicGKukTDXeDt5KfiKQ2QL8Q
EEaiRZ673kKCa9sTyVEPCM9kiQzSwUP7XIsIKU/WwZZTxZBgB86rqpkWfwd0Nhos
hSijbeAgt6SHWcF89KdHRiLY6OUyA7OIr/jVGTTFyyjymQY6r/zbpgzBPekBmFTi
cs9Yo4ma145E2VEcbanwqozmiIIT0AZtc4CuoUIEOhdRyaokmxlj31cvJ+mWIHRP
Tb9Slx68IWqU1q0OrcE3NM81mjw1Ui/agDJNSQ4JeE2Hue7Zg8NkPgrZX5gPNP25
e4xzZvOlVyWWlVOnvDG9v89RW6xRSCUSMyfHvHbl10XusF/z1Z+y7Uq2nV+vD0HL
+IMjZ0+x1004uMmamgf9SBIlTEDPoMui/6570tZm/jQ4jRvurWKl5Ss0ACm/5cAt
LmzsWwX0b4hfSK7WwMbsKDdqPU4HGnNOwf6I7s+SOHWz/FMy8DXcxZllE1jYyRst
N8IGbGaSkvbcYGCzcohh9pNUfSR9Se9VJaIgy63neGmGtm5fP4fGXKXRgorfwVvU
cbQfj9vq1AYU/fC8GmCzaXVdZ5fqy3UNfVeon7pXGABXaRdasA1CFIYCJ66T5Yco
8WZlYTd9em1ecbMH6eohqlrOT5+zgKWilQZXy/a7gW9W/nmG9iWkw2vWe3P5IOYZ
MP/LmLWPbqQAAMRr3fGomTxZ7/1aPoxVSddgWwwtobV02a38yRvQmxLcBo8QAqmI
xMz4MTGLEu8ApgaNejy/1IppTr6s/SccNIk3uLL8HE4wwfkMyRSorxRJk0W9FNxS
Si21teBqUCoIMFJoa96BdOJ6xegSaacmlcRPemZV6jjKGGoAEmqOdesfI3f0JxP+
6itDrr6rU7MZB/lZtV4hqYHceCaRdzqwpoI5mk6bYbJJhvuYIX8UGYeGryow13W4
U2NVdyzk0rhJPCL6EbrWNHnLLkaYk2bj9bhQZJoNp7YurfaaLM5ZIQa98XqkBSOG
7zbKsABJBVSd449/xkfjsqcTxfDtiJMqicdB1lkdGAx3UybZLVI1GbwsGgogsxG/
TNNQ67ZesHPSih73PdPm7b7EN+yfgttlF/dvtSe1bO5fMKwAh2xaDbd+kmauQEVa
WQFINFvIW2q5ytVHjs2pAfr6YdDliZOv39nSKasA3KR7T0SxgKjnDscVAUQ+B6hD
QXO+wPFf/SrSfiLrSNvmizJ/FAsxtzDd++4/mYwJLP+lemakdeTdPHoyGT0wCWl0
0M5YKB7rQWrdN/WurR7Yp/CYC0Knv5Resn4SizRMtuv2LyU3uRw39oApDI14ipqg
F2OlpgfEvcVV2m+6TUL12iw4vh5ZGvLBs8IIeLIkwXDWxaHrB0x/Ki/+aXfqfgjd
8U0Z47zsNK9IEOrw+YiZLGOjGPTJAZhIyArkS5wRou76ScAcErhdnk+TrrBSBIav
zbzz3YVA78LjEtbYITaSu9Onxww+FY9F206ziI2c1Jv+2uVmhErHfLFnVjMRAbnh
fq+bI66yIwwfNN8u4AvltgwutOhSQbL8tf77pVbr9zrWCGmILKu32wkWlNI0m7M6
16S8Z6eYtEzHLPOfqhXNZiLuVRemzfQrSRPAMc45XNAqC8DwVpxBwiftxJP4zu5q
GQdjsyOMlpgKO3dVK7YfgEkDrPJrdrmf+c0PCnHN6/OIPxAWLnG1x2hX69BYFGS6
F2V++G6DstquRenk1MOBIBurN0DzX2/QY3SCKMsiNQLFoMZjIeUauMa1Y+d1Lnbq
IMZhXxVtM2Vg9uGOxLkKAE3tAus3lHtGtdxtEAFpBLlZlTYOjUF3WxWP4lwG6Wf7
7OnfVF14mpfLdxzbDHY1ykUqRe5dt7XAKtE9lqbWVQTTJM+jBDA0GE3POh+jLEl+
gwmeaSJZb3nIOyXKP233J1ebadvYV93kWVZkqT5f1OPsrpQkCSfgQJjay2BK/das
fT4FLxGYEIfalwVj5gbhte0KTE30NlhOIddbnXUXksP7PE+2PxzMFvLKSZhAgLUa
gK4l/MQbAo8mmyI3Nno4NEIh6pTo6+ehf/Q/L7xKuaHkqysrJj/iRnwIYX+VkWqS
8arQEk7pFr8gQIAncnQkb04hQ1p6ko22uYPAHaCy6nYMrfcTalQqsUrq7wwTT3i/
5Qiw+6x/xFpk2hfCYIe8O1qeSIhbWjtkO/CH5M1EmdCUSe2jlUa2klZgj+B+KAf6
v4fype4p+F5D2gzHQLCd5qGmL8f0Jx/NnJIlB7drgVD3OZh2sSQRELYoObr6xTIk
s0Hg0rPD74l4VQJyI0tbu46JcjRerwEV+ho+hwTUQz3gSu0L/LCTAFt8HPaZDhKb
ehTNjdzqO+JZe3VAsO51tQf+sbHi1MGeiqUyoFWgzNUdJS745BU7YAl3b2HyjEUC
w9hXNXIYsxD47gdGSThvRZ30VY1sKApfCIOFjxMsnfh8XJfwGkeIa0jTp27sjNnw
E0UHS7Li9jAg3vKEWeSYMqxhCYhCdRUyA1uQKNe+854xfNqD1dWeqz/8SCFHcNiT
X0Mb3MBmR/rIEHvW6rfeAV/Hh7iq0nfya2HDIZTRAR53q7wDv+BcgySM49fGdCyM
KGmUidrBAmN/XGl6bL+OfXpL+Nbi89D5I69qZgWv50syKlwBFFl0xcjPG+IDw5ar
0mMSVQFMDWXpIlDfI0ea+EqbfnPkSLhVOmOd/jKBhG6O5/LuP0Z3ZuWyavTOlrBX
vhGKartBzYYOAz5kFzUsEhbdGuEMpYWO9EPtlz1McjxX/zgPmCaWBAviMTEGeByb
AHqa0eiyteISwk5cd8v9zSe4l6CM0Ljm0w0SAE16VpU7G33NLftH5Rj1l3Ly9o7t
6aAE1iUE8j2V4/rgxoFcgKBHocHP8kq02HW8GI/tAui9p3+UOwTevg4mDcoQh0T7
jwRmp9Ste9gYBQR2k+rbhldxqahfMSpRxpZ/Mtd0A8pY270OybLU+GlPw92B26ff
IQP0OZW6DRgqj0ApRFNvTw7vd3vsrVWx3DAVSaBNN4yArfkurdXNqddLbxrzloXs
z9stwiKimo5OEdqApHfGBg5c8Q8ajp1iVIUNZihIH7r+KiZwuc8CGq/qAn2Mj3P+
n4t/ze/P5BHPQB4T7ygIGR8thzV0RaZTSlF3jjF1AAHFKAj+92+XlV9YbsKxEEjS
+wmPanNHyc4j+FL7pES+xcifMcwanHEUhnA0EUTqvOrTp7eqhI+YvDdNhDhHpekq
AlTGMgE2iUW5I4yQmlpEoFmduNtAcn9BUm8URHQnlpJ44qi14RfLpDJyXvhVS1J9
baNr8RyXxUyPC96tr54wWNfWeB2Bq8tTxv2wqgCBXstFDYWUpkitpnAku9F+H391
wiQdlHttnEpoOuMb9i8//AiFsRfpv2JYm576Fv3jJjgYg25nQ4AdpH+CqUGsaX/Z
ArK6JE88MSO0EIVLuR3Lle58NTXXp1aJUDkybKh7aEhFJsWsmRGjhdQjsno/3am1
vgauvUd0qyE9OUTWAitlalwtK6Jqlh9O0aCdxDrQ0KwA4F7wUaiUllSng09N1lTO
HOOMZzG9UYt3AsvzT6gIXV9MzhRwkR1p4nSWInyyjke9W4/DZ6OP+2auZLWRugaB
LRIDDEbraIfBGO26FOTwP/xA62XD1Ezmhd8PyajnAo2uXNGZj6ZVbyaywQrOMaiJ
mpEPEQet2fDwom0nEN8MfGUUtjSyzPPg5VoWADqTrM+cD57yruTfMReLGkhTHOAw
stwzmDA3YFv7S5GmFpSb9sBmitGl8qwF8QsiCMy4qV858L2Mmp0iizTNkkZSESRj
vbVl+68UjpObVTuDUoFQhV2DU16Nymwxd9s1N8MtRvBTlkoEQlTVA45JOcu07ddf
1u///GeXzhyIC2p4EZZEsNZvT+dsno9dL7JZXHo3Cv4oKHdxSD734LuYeEuw64Z6
9N1733XgNewQOvxh9A64bzPBmPfkwAKPg7wZ6473/ZYlsBUVzRPwEUmwxPPDKhGx
neWoP+wf71aVWLcf6oKS4aUk4dSs81HGvaCWRkKydVNzLfBE6+FiyyrgIAO1aTB0
hZbJwibX+ixGDMz46AhERgVbshFbEFsgBJw8KRCPfHUxLB3sFYwQ4ZEWqw6+n8Sv
SdATEym3z59lvMy9+3tVka4Wzqz8nbdPmSgZgkUWQWsiC+1wNXERaqeatOTcpjrB
GQTpdw4MPJBnHrk7pHjS9FAqTERRb1Mr371MFnz7sAcEg9fcc8hDbEj1qkhzo7Mq
FTl0+ywwQkbuQ+tlozus8uQ0vcsYSXvj9PGsjoHpuqgDD8BbuyEuoGdIrFW2iSsZ
L6SuvJE1qc4UjQONm5EozqjvC3/ylQCmtpRK0DJRWEDPEqW8PoKzjCNBoJe3io9Z
1NooMF995vQrHRc9pc5KdGQfK5zbiJOiBZJruiQdCdfv6XqSRg1ExrYLxefh9fci
NN/RHWPZfKQbLphPQ4c0u8dbmAOKiqABzpeJMUMPPvH4tNjTdGVrZdP/Kw1HpxCl
z28GNG7AY8dPxb7M24eqM2EHDXAXdp3t3SRrsv6mIWUJ51CHvdEwieiprKLo8fZi
W4gGqKqS5tl9qCUkb3u7salhaRXdH6b1fANzVBKlks3YAyZQOdx/sT+dpNDUBqF7
erOMWF/LmRXfVlk+EMPMVmBCf35KU/e9uy/sPGiF5Aj4YR7oRR7NRiEIeHcFG7br
9FIW+QMLHnx4g7SL+c71k55I3s0vMRyy9uFsU3VpYVyYNYaU/IFpQGoB8ykYPxmm
Coqs2LVcLa0eMv8Gk6RLK19IQvgzms6OW2IhodgapBt87TYGxhdFJIEBwDFYAq0U
/4WUrkcEvviP9VQztgp5vJhVTuN101+5gtBn1gnYfIfOPTUEcko24vzsNautAziD
wMQ5OhEwylPIFjYIAoyIjKX1DaAlj/B6ikZoEgQMF5JdNSrn6JF0IDvibO1Qwptn
e/d/+Fd/b4cfbIDwyMbBx2V0zR28CEv6ns+wZVWCJMmLnuBOy/3ZWj5wgGDCnS9I
mvD2opoTLyCoYIqFcA8KnsQcXUgDXVhGvm03CW4zXJ/vUoob1axdf3C6ecRoFcmh
eawxX4R/10zTXtRhhYQSEytDP2QqumTwl1LxCuMBwX3FQ08FNdCNQqSMMsTuSGFf
89K3f02Hc1YNE6M3FNGdKgiHu+ivL5Lh3jgknK5f57mFufGhmE3pW5gCf7MXO03B
aYqP3c72EpPR2p/QFvdkeZX/Dvgrtc3AwublqHzOqFA+JucMEdFU8oR/ihVdciAo
PwncgvhGZcnrHuYEcLlWitzj+vo/ZUnYqMdia+CucBcLPfC8Lm4gLZOj3DRANraR
2E5+LBYbQaeCV8SYlqq1s2LZ4819e9s8iCg4urS6WwA4XgpBBTfJzWjtYw3UalnH
ogSA6TLWctpaFw1VnqeWcbapz8AJsjeN5TwKUHy0/ccnCATCiSJiuRGB97Fmb2Ix
LPbzKFwx8/nCUzDuyjm4voJjSiIXXo1BSNszTsN1e9QzuypsbE8B0AmVujC0Ftdd
+miCpFgFHQBLni09W/Knk3sPo6GKksrQKxrtbr7tNZStRtibkxg7oBBxITq15n5w
laARQvmkhMh8YXEdt91Nqen2s//0NWItnVwD152bg+WGdjqVjsCuqK4NzMrogCUy
0/j/ddVgfDqlG9XnBzjFxbEwemnIxIOmsWFEF5QKwaN3Mm7uxSCKvi0l2C07J0lA
czUv2jWuzlZOF2Pq5kbykFhpyQ/+zSB1zyy902r5fPTWtxqFxmkykp3bLgR0mqeK
pT4kbnUvjdqbXA7RkyM5KBeWpJjVN6lJ+rBLFFIuD71D5n0GSPJUQlM7EMDaxJlC
fhYFqx03viz7sY7wGB5M7nWEl9fsjWT98Bcd3SjICLkhimEBXY+TPjTlENB/QYsK
93WjDSniUMcuHaAON4G8SWGmwCMT2+YjQfLvldLRpJp9oNmKszj6j8eiWZUx9gg6
4AboaAXUgsjEGYVIsgflYIsblGmAkwaLa4nXMh4BejXZL0jLE7rkVf5Urt/3uF1Z
VweyoeU6vHcBBNypuiJFutcncg1g2LBnlZwDWiFiI+BtN6qGyNvmKWJaGTrJBWib
b+ECc9NseEtrvktLx89lXkpNtzJhno12zAbkhdj0Trb9uwQFjQhzoE4dghTF8qCF
0//PgpbfJjZBFlNHXJQUwqeJAPuBPoZyS6/0006QNejlhENSUSFfvWqBu4T7/5k8
1nlzQnvdNRFmx/cDxPyuGmdEn3BlTj+3JnvjH5nVW8eeGpcsRLZMRpB4O6W0Rluy
q+IsU4Nf40yOlBK5CHuVBSa56Ni9n9WLKkpLKDTcx5vSk1SghwvJCUwbztLXcWXv
B6j+dhFFbeL3NaG6MrsM5NMujFw+1uiFPAst6G0sSW9kV/CFFdJwEEm7yDowZW8B
U9kuU0hIwaawZG7iWHhmaREZPWSlVDdYzO0CrCk6iMTt4VoVz072OPW+1g62yCBr
JMCK/zecQAaJCsZVT8LSHr8LkyM3UeFHuklrM8agr2Wt0WVz2yDqjbQH3PdYgZBI
BSnv+/eOgfYKHTyq6ixXDnTLZiIRLI2jtk1JbTmJSz2nnwUVJYBto85SnMR6DnrC
BIe6lcTisfrZDmBuSVBopKG1NW20mhowCEs1cweNMinfUCfZm8p4u1rKQx5Uk4C2
fSlVkTxGxorOcrTGqLvcZOS0wHJ0i/dN+togeskhc7QvZORNJ8cTXEluzNUvud72
vmSuqNskZNpfXjpoUWqgMnPg5UQxiPX/WREUoiMkP6+f2EPUdfka67OdH+Iaim7k
4+Ot6UaASQrjFM4GVBonTVCsScbjmhHCuIDjhyJU64vk5huAC5EmUimxtgxG0x5X
tFuPGvT7tIU6uo23tZyz20A0AvDHNro+4bV0t5EeZG2UG5Qi8psO/lfzKJBxPxQj
9Voe2O8HKXbaGPEYg5zUiwe3aiQzH3K8YmkhWr/W1yt4N/5mY6vC21upckg0i9zo
p4kIp+pAIDbplKAdC+kS9s1+WZLCRcdBy4jTUufyIGYUcyIieAl1VE+p8rSAAby0
yepSAH3iKnLvCNaZDLmFZOtcZfRrpRKyecSGTO3qwaV1bNszrv7qhcH17c+Hm0hK
l1fqzGiJWXsr89+VXFaNNqJDplmcpSLytZZMwkKbOeuC70xpv2FcMNCNL4109QJf
I64oAMoCecPYRIu996EdxWyork8/tsMkXHLOu+zneMprLb1YPWKr3Gzua+uefR8y
rn6VRC+uNSMtuGAF09J4eQWJ4h86JMzOF9jXJEQnCW6ghDA2YRfZk0Jy65qWjWcD
pz+Rxj0Cg140Hp97SBOqQux6V3dB0B/xZfl7QY+hixMFVwYrxZA7WkPHHjEfrGXr
qT6snY6N0cXJ5mDlms4Zm3ADkpJ+4m/iQdvNgR3uOXi6a3RAXugnchUzvgDy5H5q
iQMjH4V0HfxWGIRwHzS2mArgp51qToBQbB05up7ZI5PsWssMSiqWu5Oi1KdldDFU
pgCNN1Y5r96jjOG/HGePYXtfDapGbGDbut1jheoKka1ANNdUNFNjVREz3yKQPGHw
aZ0kmY6kBE0A2A8C4A7ZLZszRtpBm8d0hdkAmSNtBkcXgHsQqR2hm0SB2xqfzA2t
1my3iQkU3rv5NTRXtv4uoww4CfJvJyBTENLLK21pAOzYS/XPi+t2tUlD2AswI8xf
RPrbL4B/3mPB9iQUbqBfjIQDjtuQpLNzPxOsc2igKUt7u9eEWsvPyvceKKXeUvfs
LYWyskslIpjsH4WJzwLIjsA2ENKE5CxNgRjfwqfY/PIlhxIDELShz7LnH3Uei31U
S6Wgul4HZoccmUw83szlBR/NRYYxocASLxhAHU2squbOc5bsRT/GrrzYyU6BbQLf
SjG9v7g+qCIEmLoQjKmQIk7DDPRZLHKozjT4lj0XMD24EF0jOoGXu04YDaBPHOF3
eIRux/xZzdnNmx/Zqqst8z4te5vMXUh+I6anuSAxHD/1H8t1E3jhbiOCMVtJhKt4
O7YvY2fWb/nWNG+mDW1lkEsmi5bDM/vXN9LmY8gnQZ9QDiO0oLFrWhRMAIEvqW0p
ivpXDzFpildaBSsqiOjVWLUNKEkMY3TQ6n7xzvMCGVsdeRvsQcdDJBNce261kl7k
JWWOsXt85fianjTDMOCSbItOHzUvLwAtTEJBCkgX8aq7N3Fa/om3g8fTkm35OVuz
6GjEPhzgrTwx0gkrOHJb3QH14C4y2pmxAZi26oKzJM2QaJUETIyShj4fFEl8fp/L
6QbiNKSNxlJmIR39PW27uhfXOmDhU3cCrI2ZC38PuJY23sBzu8veIHLxXSjSmRGo
6Mi9lHmNCvVXgKGktSKpeR2NazmSI4WOPrN1RIO2JN1n1rD/rA+bw2Y8tTrVtyso
67dMWRohZA9mdrDLF064OgvmBuh5dgHuc49zcrEgy3MuRKLT+chvcuD0gCzoORnA
EC4RC5fzXCOGJaINB0GgClN9+1I54ON9E4qN34EN30l3No4Dy2brv7IiWzNNVMaf
2EGBKtz5XjHZ06WRcrSkUle9cFYERYzADvSCKklzU1vAuisAU6Mn7tb6Naea+BV7
CdQSdElRACjgt9SWV0C5nsIW741Xw6goon0oq0SfhpUl7afEQmxMDEtKcazB0xqb
8siirfHT3E3u5fcmqwusLEt+ADwDtaLxQlDu0Jgf0khTTIy/Q0d/m89Zn1BJxzan
HquKxOQPEUsIXKAOcnZwOAeeWZTb4VCjWoFZ7UMBtwVeqxnnH3OrR2hGZ4XyP6Sh
yZCMDEk8qxfnKH0IyP+RsuTjBM1DmCm9qMEeU98grwE0ahOVrgajSQvMjYqUMCNU
MWyz9RlJOdwceZlioS9P8yBxVp7VLD2/dwqx9a3UmJ9LLczeub9DjpHsfW5ljglg
0gUihPcq2glU4TOl7YymseJ+z1Z9w7aKrK1xWZR1WMmiKUtPQ8MexNbnYvJVTh5f
1HSg2qK9N95f7hI1iZwpqYabAeRB2nnEdANryjGUTK2tkcsJgxdxDLH4aXt0YwR4
L0WbQgmjGJKmBqIxxCG+k/HFPPrC3h39/d0Q5bs4/vsjQvac5uLwtzUH3lO2/o9I
LSy8udyXSH+wqjycLqC3M6FPOg+ZoRsc7TwpSiFAel8Cv3a3rjKUzQUf/hm7tAHG
APaiftNHs922uytoefrzKAFFjAIydn3UnPW4QZ2MTMzvkjwOESp4HCCCT14qpRaO
zEIZKOsnCSBpV1WTmlMlYdWEg0P2W6A5bID1fXu/Gwv0sjOdFOHX7DQ4AmEVVJ1Z
yTAznbMUShDl6A3deTH7tlsVyXH6TUMO49wxY/PY2d7pNsAZgayq3pdrtjVRISFy
agzBLpKT58LeNP/XV9F9Wwe425GwbCWmRebsglUEB3fS+BzWoSqML7SNQCP5Ne6j
WujsoBAStHZqmsxYqmnkISrbX/VLhETjAWEuRzb0wF6/bf6qwXmtOIWeDpZtHHPZ
FL5OpLpeba+1BsZAXsRkYwo2t/h5NAk/b9oH8nkH3m2nrKTU1Q7HRrP+Dr9Ky6ob
NVFSLPdqVl6aq7d+eCkfn4Mm35+6fynn4tIbkPiPLR/sY4QRlTDPvcAynFHmwWa/
q3Dn1RIJJgAdlXFKE4B1vzUUTNSbkUF6XNCXX0uyNm+9zz3MFLyHM3DSly3k3b93
1UA9UqKpPePieA8YFeIE6L8kN0ur2z5/T9BHsmgl+W3zcw7iKIwuayEY69a5nq3V
ubbCpMBGkF3uKLLW125Kh/QENtaxnSgkuvxm961HKk1n5Yvpxqho/A24p9qCPO2n
3TL+XU05h96Y9X6GykIRcse1ghfRObxEYH9L9QXbZSdBHybFUiGUJemkiqPFBo8n
TrFGYPXhlKMOXWTn69BolwfpkTvpJxNMRbeTJqGjL4o3+xNqVsbS7899FTs+2GiU
uyc/iafsvXfmHhTH+zoioaw09nR5yTyA4IyV+38v1stAPPAIAlxmznOwwD3KK4BB
Innh5dubf5rKZ9dMQPC/3ULdgzDdTkCfiXcPdfCtbBNIJlnG62GDK1EoLPo0VzYX
EHWrQAZAL0r7FOsron+DogcVgYexKAxLfzivnoP7CDeWJmDShBPtGetEbR9ZvfyE
wT+e4FU/iuQGRW7HNdgBTEP4VwUPs2zeuo1qnlJCfsqNrX9JsjSFC7cxcNpn2IsO
4K0IUZCHA5x68p+InBMVNslGS5PUxFoYPbLE8VnFvZKOBpAImnTNwzImdoMKICLA
xFwHxN2m1px+evpHo8QGsu5qj9/vzo5elIxGKXl0m30Rxizk/b9h36xnLtG9VHku
O1dOZ5z1J/yUWyEQonDEd02A6oTtxqCJuUAgW3oEKo6uW9EbZPsnszEBOZfkWX7u
UqtYeyS2ZYDNemOcDwTHz2nAdbltB2TjRZgkpqdr5aI/cSGpvGNEGcwfiEJx7sZh
Jn9RBknrafsjBqMrZFb1+Tyo6H/PZNJqL21RRVaHcP0C9pXElWCIMqzrz46ct5Ft
/SwEfRD0zMIfpUnqYnvPqFEar1tSBOGYf1qR32JM9Moy3vwkHZHCtgqK0i5sR+WW
TiuHDUHC9YGU7UpXNnlqyVTUK+xBysWP6sygiBOapvdH6fBFVbgq1FnuNcn+izD4
hoXyq9SCxHf1Co/S4URU7o/CH5znpaXnZWdkKl+jhJiRRVDcXBvts0i33tAtkpcJ
J7BVWuY7X8iIDqfmfBIl/5GDvI+624FzfO6IIr0YC8L35BChZ7SR5yHJJZ5gLYfe
2a2FRDxrz/HidW6+CWCIGZN3XZaUzHystl5JpkxfC93ATEzf/YJbmnjpcHPv8wD7
rRr722+CaLhlgUMq7JpeFgFOGJmk0Xvv9ARnVj9dJ+f94OQLkT0CtZPLwJ6+tAa3
KpRsEGA9f0SF/eHsrEpPNb/6oZqC98ovy2IBBHBta/fMh95k1w1+3eYfRn9KZ8hM
Uf/DkpLp0lHQVbLOP4GEotDbSxTZ+e/sErXaviFe/BxKld42i/vA1mHlsWd61WBG
prKdy+7AtmnF3KfHZd0iADV7HAbKm2FCOn4MHaI5p7urAGL+wlRcV+3pZItaozR9
ETk28HAhGIXzPf+pdPT9V2X6Tw5b8o+vNOMXlkr2YUIWyfIwUUOUZqqbwc1cvBJq
/D0RWscZjj9wBz2kTlGDizGooLocr6a6tkubExjc4usHqcZ5a5+tpNJxnOv12LBs
Lfvq9LqLRBzd3f3bMDaXersdamZEyeO3U/SVBV/4Mxrs5k6t/gHzQo1wES65FCe6
w6GSi8bV7Nj0tB3utXTniNxgs0urBkdEZueJ4yEqexrFEkn+qkMHK90hbOlT+f5f
mHSY9UmypKpTc9HSBlKF9pATQVEOIQj6mfgN0Q1v9q3paiNE3/fJ5t3DZKx3X84a
LPG0trc9VM8XKlFte4rGAqyYAcRURZ5jtH1YsnpMFVaHaVtp/NCF1jgQelf9zAkT
ZVYHi4aTAi7AsJTuLN0YQk+ipueQ+fBWnGpM5ryOdEfGqmfLo88ZDt+LFsYV9wZy
a0Zy4ee8F0cnqBmQGM9uZ72nJ4RhajKKub633+ol0tB43y9lyGq3mfEqfTet0ooN
E2oaug8MF8EXqXEHdlQIzN/4yKvXNgdmLKzFa1vT9dgKUc+NuZ5tiAGRkPKJal5i
1A1MvcceSa+UA3AqzoJUDwrSy4QWKJOgLgV8+XwYKZkavqi5u6gRAQErpi4sIEjl
NU+Gegsv8KJV4HQ/hOx/z//BHe6BgvD+tuIqNxKv5rrLUzKRJz7XYBFb4RyGY7oI
4Bqz9pIn2SoAjQHqsC2o2Xgr4MoQpoDy6IZHDExM3U5LUAHG6CXd+zTF2QXdfFNL
NeuL3WpotB6BnLv9zCxCLUG4V0hj0+2ydnLSCiiyPgsbubEIKCmrKeqeIQKv3AMB
v/Hge2cryIG0xTxvNcUklNIW3HHJseiAkbcihRFxzPblcsSRoRsmTRgIiMMxh3lp
sjCviE7av3g2Iipy8ZW0nC59Qjbgfgz9GgkhBM9h56vd//NC/Y5XqwiQgBTZCnKL
K6Wmcy/1MOwrx52k8boa7HYTklwByVVb8rtKxWGezier6JRPGnLynLkbfvHfnpVw
7+8+l/I/2F+CFPzZP0kRgqm4nTmouC0yH5+tdegrh5UEFVCAgvEbh1cj3II7/+H7
J347EVb9PWVHMlwNyEDRmxXZNeRV59FD5uReoxwEPpyavB8/pFw64vuBLDsQOKfD
uS1GE5U3na6L5pp+nP/NWUJt9mjMNehAoXkgSvQgJADl+deuS6lNByErXBKgWf/7
A/EcdrIZnEMd5PpoKZVKOiBQTsYWXWZXJwIdyeOcGkCqDcRCXhhyNaUZ5Y2ydU4H
PycdPTW/w2qmN3qlXuSn6uxfTE02TveCX73w1GFu5j4AqHW/jj+MNQuB+HXiIwmL
TKnk2dMcf8MHOsoPP8gl+QCTTL68PZIQkzykVEdUajln5Qeo8pdSlt5keMkpmdox
`protect END_PROTECTED
