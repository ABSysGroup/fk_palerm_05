`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lN6TEthMp5nuIHFUw87tJip2RcGVfHI1oHSrtFN3aSeqJJ9rSJI7P4SScxhiYJRM
XFsfF+mY/4LM9J4U4xd0RksGfSsaUBPxu55DbgSvSOwEno8PtwslC51CghHM8c+U
uy2zruAJTxZSzwexMMQmMkKlZaznfcAMiR3pNcrUd71PLZy8sckBdZBvB6ZvG2Yk
doBdA6ixwZdZxHYQ211/2N1ypGTNR0vcdkCZLh3RNguDBBIOrx8qfvathvFXE8GE
/lf9In6tcV3UG7l7m9PftmIr28b0qJ7n1IxgHmpSiNdcQ1fFZl0kSB1Wcn3fydlt
NLydCYO5xCY5r31nkaerbSRRqZwT2Rv/Nl4IarOi5/QImfZKPGGu62BsJqi5MiT0
zoBpXZmHKax0oRxNVsQuKwOvJShOrmND7hri6ckhdc/nTHOXGDywtRc8Jk/rt4tM
pDiNEMon97+EgmFg1FbSUoyFJoYoObEYszMNhNBardMxHV6d3PAQSS4pwu6Ftd/F
iqLmdbz1lKIkFaqr4UhKKgk1phLDbWl9mrpqKVMuLGpPJOws8t7RUwW0JHQWPeYP
4KisEUX5/LxlkuzGFNuTt47ywFevozA14bA50wzD2r9fc3o8R4SniFOp0rv+z6dP
450JgDqvetjWcn1EvZE3fSkd+y2mSSG50Fcn5iny1tYjVTEYTTqR2mjhAzPVNbKO
jZtTfTTyJ1xODxuUhs1uEAQdBvyek1cVJuGAKEyfE4nbVVkCQHocjTTHU1nvQePj
UHSohuEu9WQMB0KZkirCE8+UOQQhUKziUvAVXM9gKlCEWqWVrWnbM7yAwZEzJFnS
DuyEH7HEdDx3l0aieQHP7B0GSK7kG+yPJQWtsGkjfPwJZ8DQftQP0JzELR66psfY
u5bPEmAwR2eVuJtKWB79LmiQ2dTERxwQyK50W7MposbTIjZNZLCKNUKubntxccyj
zdUXtiyGMEql1ycueOccdpX2fqkaXfw9g6RKBm50/WGuzCF6a9Ee6vwmHH7j9fko
WdUgUyd8b3Fh1otr/nKrmw/mipkDx6kgQij+En8aMTZ8QJn6JsSijweOyRLmupKd
EZQ2mVRdBJzCrA7taSvyBQYmRUkaSgMtmfr2QPvw11tHUFV+CDix6WVhDYU8lVuA
nWSplJez031S7uNyjshFJQ==
`protect END_PROTECTED
