`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ARM8HZJsIjZVho26un/BceHKp4ExqL6Gs7IFZSIcfZ8HJNpfQ5x4zEOIRjLQe6ZB
EIs1G+o4OspVPkzSDELDyfQhfFmRKoCqUd06YuGW6o0T0vP33zN3U854G2VfPxm/
NS5SS8+h5k/btQa4tOjvc1FO52cDGv6q9cBU4v3yFRMxcZKZEwJPTjpdUWHmxXGx
Avhno7GonY7bKAMSzvuAQKn9P2opUfVzx/faPEltJpt9Xc/AFmkunAIGmE5uB+pY
UhBw6nlr/fJk5yvmmURBepyEP9lo2FGB+zSdYDWeFSOv5kF15w0WXFmYgIRT/Wzj
kO757EHNtSsHESiFpE45O6MwOrkqO6u3tmHMlJZWUR5PQ7LE90/Ffal9e2e86n1v
CPFMUW0nT8Fd4blSd6nhlfu/6j3x2EbtQhtcUL5BYyHSVOiLv+zoWFi1zmcXgGmx
NYzND5kPKMaQDqsF4iBQZJhDUcFY+lDhoOxLmcDjKKat+b9UtOwjVeAn6xAp1A5e
FJ/51/Y4v+dRsf5U0lcBT3qHRmLP9l5I0HzNSlpoQCzTHVY3Om1yHVdTlS0b1GBr
EIQbGSmDNpcXNxrHYoeIxoN7dRgq4raBNKSQSenB3yNZY6GSL8hM0xTg1Rl5Fu3k
nCLn6vwhtvBgUMJByOrAio89ZI82AzYJxkY3i55LQEkMhDd+5Fppvr9uLkA7HmmP
sZqIdwW5augklqup6zGNvGmA28+57uxsBr8VCYj91/oVZfe+yO+XCg/ieqeNBlR6
lPuMTUcNvLdzkMGZdwR3zTtznox4mG1Do82CvLRdsDeqQ9eOQDxJFsxaEgHP7mK9
P2sDUSUu3CW2KguBXluYbOq1RbuYqflm7HUguJGG3AtspKR2Ks+XALf/LcFMG3TQ
NPHi4Dlj28Aom7xz0Hd5q4jkFLz4F9PDrt1M5CkczwgdJez22Q+le5l4oFPXv5q0
saTc7SL6naN4Vg9l6maGp8MJl+YCu/g12DrxLsmPi9REnW1hQ00Kes9m9QZB2Sy1
bV2inbHjPoJNta4noDi9qbhhpsGENGqaBM/HDx8VgFImq5MmW3o4tTRCXqFxEv0A
4zAkEF1CW+2d3vPmCP9pT2ZrifyR8oOFWgLT7Rsm3qlRUnEh772qZwSXIIxWnMTe
dhC4o/LEISK6gpdR7Z8UFEqcqyByL7dan38W7tjc4K1GBpv4lSgXeW8F9XI23mtu
F9xYQD3Cs6PIr2LaQK+o5/qtNp4yvwsVcF4JnWFIYcET3SqcPFMpuKf40+lOUMAH
mg+8qDgsiS4bBk7pqOZmaj0HJEPlcQUcBElJuM2O7Za++c5xJIxuMxoXAVi15SST
OUMM2dqk1uD3O/S5V2diRHq0Dzkx3d29+XaxTcoS01IMRhccBamxKsAf8m3nCeCH
LOdUL7Uof6BSJva95iAKLZSc7nuShbVurh0dO1uU5dp8PGUx5OoQkY5UurNkOVDN
7+rtxvTMwOZL9hVbwibrmgNJXR3K5v57nMjEehjF04vsMhImEbTnWJ/UI9x2D2pv
hrbJysvMtRvIS5Fl9F0fDaMNOY5ZEw1OB6CZNt0glhOsiQgnuEhGSVcJNTKfdwyD
aE9jAqTPoVQXxC0P4awQyxiBSvlMgSo3p5LSawixHCN14fubqiAbB9bLWfpL/B81
HQWlsefW3ApiQKoGEjsjNr6juYJiR1JgEImelCLoEfkagNTtdsrBpZ8WNHp6axGO
mIsrG+5vl2y2uuu0hU/eL+vL/BOSh8PIrd2B1vKHYPCWpLIF2zM8Hlx9kr4Gm6iI
zi9xtOB4UdiAVY7RVXEYoYxqFIRcH9EcaVe+2suC4Qpbf3voE8gxO92AoPiCPjyr
zwo2N0EJmVHDS0Fnwc04Lem0ssdX1L/j+IyijcBM05XiPmYMST10iqX3bZ5GEdHe
igxXI3Tj4AhiRvp6MKeM5lqPRk2K55J2nL+XMkkOlW+AXsIb8t6HnDlxmKMBBZJl
ncBhO2d8hX8s5O9IfL/kHg==
`protect END_PROTECTED
