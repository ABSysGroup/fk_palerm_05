`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IGpCO042daKN3ZaQGl4SLSK1/0zUNxbN8iIYRESwM9bhzWS/yflefLoF8b8wSxUL
zyF8AwQc83qjsdslkbrvnwR8r4MaAOPWdyxLgWKcc4VY7+HXEbZ5xdUIREtcoK01
1AkEVPjD7ZmpjfETCJpN8rsro+gpZCP/1sXNSjPhfPjEUHxUO5m8s5Ebn/h/cglw
mkf9a6z49g6MNpeTGcjp0eOatnIznMfId2EPuVNdhVe1svzU7NmvxnkeztoUyQsF
EVagBWS5F0hemLYtCqMy3AVMywkenTOXhEXkpiuQ8aEJ/vlmH9KDAyL+2Umq5rok
rUVoKiUqGGnZXd0JLEDtCxAYIPcRqRD0qBl9odsFNORQD1UmNmcOrGh54UwdKxP/
pShuCnGqZQRfRT7LqMFW7FnLICz04vqfQXikZYNL4ue/F1wFwbuP93BX7CahEviU
aRmcRlgj5/KjhyUYT4YTUx5FuWiRxEsXlwX1DPUQip6+ougkVgVtv4CGGKqU8ObW
lJBTlQW7x4zAelr0c4KY8MnK0BsYf0B+kYTT/Fn6Wbp82IcgPH5yoUERtDzAJbxB
eu9uCImp165+SEw9GVupoFa64mWDN2Mtch8LC2iU0GvyLLGbcnb8VKFHgybHAW59
5FLvSKrE46stHUynkhrTSkZFUYs5TuWCrTkFha56d+xrWmYa4SJZTGdRxwDWHB/e
t6Lw1ljS5w4BNx/iTx1LOlJwKMbJBSqKOG8ewvE5817KXl5/heKWV54xRttwsk1n
JxWqgrTgRwswKJeBnErhlPLmEgSKXwEcacA0muLIWs4=
`protect END_PROTECTED
