`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CWbROJNZdSI0aamm2kVg/J3fmWE3l2n4vgu0L8DH8oCbcC0AYgggApNqf7cWeXJ6
veqv5t3kULPvDEG5mdjQWgyBL8KP9QFGDCOGMGoC9ywYWX1DQ/4nMnNafHhNqyLZ
VBqs861Lni7HdmpjJJScsnqOVJjWDXeQPNVM/hZYaE0VhDawmKdqAxBHCX+40EPb
iOYHCsjfuEhSw+G0YpOLzfXJn/+pSgdLSxgJt+RvH8IHRYhrvy3osmvxhY74FqRC
bxjZM3Dq75Iv2fKvS3V8hqcfKCI8VnzIgVIfqhNi2kD+qLud76Zmcbi9RyDYx4CR
9s03boN5tMcgatgQmCfqznXqVd+6xvuVy9nYDIc9h8GegXsS+EAqci2DCnKX+ryF
`protect END_PROTECTED
