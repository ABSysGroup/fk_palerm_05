`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VGVZ82cMiHJX61nfCs4takrhlUm5vHMn1pXAdfGT28OwVEH5B7VVFpMs8iOlPQ9m
USC/as/z2xlGCz9GTQBKk1Wm9cCv+f75wKSKynn4xwRe876LLa6UwXM6EUw66317
kS/rBI/YA0N+YX3YIL4FElwjlXSVNxMztsbWJyEUxGdqAwswjWV4hsSeQ8lQILt1
U/Z0YwRuxYXYwyEel+A7cjhgT8BeHb4KEbG79qxnQVOLWW92teW4KrdgcZ4aDHTV
`protect END_PROTECTED
