`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
26ntB2IA6J6yVAZG7VMbLTMwnOZKlY72v261lxr7VFF4/AKxMsl+lnaxYHIM6RPb
0nCYitLrWbq0Txd0fa+tf0a4Ic31Etdcl+LHgqGhqf2++5X8E8EQuPC5CIlhddvd
/ydc4sQa7j2sUjoLmChmBvVhRftQMRP3lcLSTe0NxvjlCVvAeTiCuR2Du+473E6p
+wDNd9eHayZctLwxyzQhf28M8fczed2zYxxezjhpD3KsbbNK7rVxtjRuWoDIkfGQ
5iPBC0yVMwZZKdz6P/9KGkWYsiUZLfGb/na9E1pKt2hxsR6ODw/48xyRLujUyW1p
i8TLP72nOx+S7o044kB5kxI25gKKLmG7cKiBc94zt5WT2C/sI5tKRRGR+FiY4b60
qF1xHuhRUdiPjpb0aSKtO+XOrPf99zWlzigrq6htVHI0Iled6cHx6DHC+0SfzRvS
FCnYfMRzl3U8CJNypzyP68JjwcqfcXzNEwV/PdKMh+fP1g7AJlp2duHcQ9+gVpWU
EYaHkjeHwJXGQA+hRFF/CnQM4q5Y+1wZjGtfJaJf1OICoHJL6XxPiOn4V7yciZnU
K8oI+4KaGEyMdysPisgkqarP3TOHYqkKRqZEUOcvDlbPf4dZDD/tYQlIO/FS6cMo
Zc+dtZLla+FmZaz+FiWJ8e8viLH6O6ONopq35IeMq3nHt0u1WO1ylroby3gqvXka
Gvbsb4f+CY6cKWt0IooQ1fOfjw/FqmnoLCwFUpsWKS5FR7BQK/l8c9NXgs92yrww
xM41iXPsZcn748Dl+KoqLjQwOjsM83qrm51vfCtGPgYJzr5PEjONgiyqzc7Nhgch
4qXaBi6wh5taQoQttU+gs+7xHA90Ss6BAbVGT0tgjcyKO6un9yciMG82L9Cr6SQL
x03ZcmQb4wjCozURSbUAkEnjFQDpXdhBRKj7w5tfZlZSsc6Rg2pFNESTOHZHgTPQ
ES15e1yBp/Ko8810aI1CG4P6nm65Fu0a9Q7d9nSP6jo=
`protect END_PROTECTED
