`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P77vKrVhLEYFr2iGZvd+Iyafa+oK+M/Y5+LPunP2XYsqLMXZwOUlqs++f0kj30tV
pYbLtEZYFtK6uxdSLb33Hg+oCLtIVQ6vDPf/d5ZmXpnxxhPCa0BYpGjcsse8a6aG
fcFn7zz7LfzZeBHxLsrh1geU14QCdOylPFQBVEY3C4wKsMM8gE9MlcKvYdHGwMBT
vds/0KvtJ9OuBr3/ZsDZYiou/1zMsgySCLFQYECGeshLuuR0Yt5o6KbCBNhEY+Cz
TTA7aAiYK5tSYai2Wuvtrkq9k/TOfDhuWdmm0RtCf8TTC1RFVzcFIkfVVNQdWXEd
OjgE5tvF6QN50H5c8T+Gc1FMASf3FW0a7N2EEZQu4WDdWEYBOf8JiuAeowpfyFSU
z2hIPgMmHfu/cdNPVnVMjUhiYuPKpDar0HJ41oqp+IBQL6W8BrLL/uB4h5fHq6cs
FExqrBulfkKiuLNNLIFYKPWZMst0zM/ui5D/4QFCKgABDi6shYhckDUojXiB8STh
VxE4DNmV2Q8pMGGVRvaLlsaYqfvxv2oaw8GZtGjMHu/3Bhm4hYr8aEWFEfgM5bi7
iDgIVBgGC40tZPDHdWpBXTGXpu+iHeRNyu1M2h4DXSUOMClxSwlAJYR02UZtJDpQ
M1RBUeRZtGNf1bf75Pt2hN91qSCoZ/QbTGE4eurtPV7eU7MFDgCm3siPqJ8sIS5I
heTGHpEthN/wE4Yj8ovszbFCP0Bb7xrpWeZe9j5mkfDcKvAxBXa8R0cExjnTyEae
dRAepgIufCptsVk8+YsMojd4uk3ragBBxejnPOlcCB7q723XvU5RG1nOLcxUGl5F
Tx4Qz1FOtJ6UnqpGk+C+AkEC2VXXDGvKQriCmxctxRZnPlBPJRxNhbCGg4hs8Mkx
eHglZP0i979kzqq8kplJZfKaySzpDSVvC2WMJGOsvOP2WPumqfRPOrSFJsBOkaWr
JQqt0i8jiSak+8YYwLatNfUDmIOpUG9Lmh20hIBWHq29RleLLop2nyYiq3qg8KsK
NFQYSnJN0JcHIJhukgBZ35tvS0s78Ha0K5o1yGTLeo0y2JsrPg3Cs9fIP76aDkIs
6cVrv5IskZuED23+WON8wZ731UinmDLBz119GWJeiHDioDVBd21hln08L74U52yA
1yVsyIWrSo3psYJCQAWIoWz8VxaNvVz2qhcvgSkyoVSWA4JR7K0YmMRqC9kgYEc7
VcBuH7WWIZdmdC4hUTLYE9FA+TU0OKYHBF/jsv83q/gFM8e2GjGJpiJi9Myqtyb4
iwsqAnCZww2IOxpoj2a0ahxfp4quEhse9HBMS/+pH8touiTN8BjzMpEOmdTCi7mu
oQsanrOphHm4hJRkBDoLliurucuDtq2d57/hx4H8FS/5/HEs0WQ5F58Yj+1nh6X6
LuGJBNWjoPGvUgT0AHcjKSuQmnDIosoj8LjsSO2gZV4lDghsOQuHAmRzaYO1D2k/
lZ5W92vwaFXqAJhznfOc0LGW0rYVbk5dlXbif6bGJ7pDP3mCmjT8wWuHacPXDN9r
K5liFsFnSk6ggJYcW/Pc5MFQT5ufwcfA2hLxolP/1OFh4IraJPjM/BkBU3NlH15Y
6jTDrCq/h254oLAmwyeLooUX/hDqyoMF0pnKkyGdeVbAcajfoN5f2vI1sUOBI/j5
3Qjb2AQCy92Gpqy+isxIqA+WPl39YZqKDpf9h2objBJ1PAc7oKop9B6gMYymEWE9
GSD3QW+X1TUZtV76/DYcyyNAx4hqoTkKt9Lcha3UA+W7KXiWoNn4/vGq7v8Zvfvq
8A3HyfutopMhx5wlIyu55G1+9axXHQwKvYElakkXnUWLynrvgpalfm5kvFoydKPV
l+r9A/P+GcmfuOhN6hCKkdChpS8etf18ajdui5pMxlGNMSAP/ipEviWWH7wyX0AN
L4Gtt3AKDuyD5LhvOqCBg+UH9i3m1Bpj4xUh1t4d9Qo8K/T7vq6sPZQI6EYbunRV
xQb/XfDny2Zt4hkDLFdr8Q/KkH2CpCDJrEvON7/LqTyhH3h7xX+eyf8lMkwjx1OM
twYnIGoac3z19fc9bkoJc7FsyMv3DWxx9KiqgIIWJcmmVdVoNsuXB166P+MZTuNF
7A5DMDZclQpLpLNcRT8TETwoDakPTWJqc0W3jiaxCi1zN7bJdPi4Mv887jdXrS63
SGa9Xrf0gRMtIH4Pp9/DCPVKKu2NkHab9aXWhaLJB/oQsHCnl7eL7R8nvsOp9gB6
fr1710hq6BWtTjM4kTJHfHQvP22EkCJqhAtGxkiIOjbY9X4IhcA2H48HzHpt6X7V
B/xriFQUashyIsVOI4ryYFWdtkXech/HgadQk51DhN3glTadC376D1e+bFo2/oaD
78rWSxcWhD8f4Y7a0maHGa7Jo2IbUoAxTzdabjB/dsSkoibryuS85mYLQ9dSkCp5
W9h21Ud11skfn6yyxKByrqJco89+XVBvphswZgQgfRSx0Tl+l8sS6RxQ5hH711Ap
SIqqb9O/FptVHEZriGbLAbaKyT0IDhp58m1eX7f6JI5En8l9SWOXGItJGOSmNT7E
A4HWgX2Yw17F72AfnrXem3E9wMvNHIvljCgiK/nSQxsglTwUniFRkH4MpS5ykikx
SSUVDvbppdchxYKmWCPcWmKY3ZzvOC+6E5X4VG1S144Yk/6NvcFKs0SEKXqYS9sW
AfkSQiMj8GqOSNhnUpXpD62h+KE4e3j+F9Hc9vPw8MF4gZEDWvhUTYRQWBy1QEAM
AIGBhzf1ULBYLyZrqA1Vw43hdVb+qOBMKeCVgLSG5pB2BJvoCbI+IzNnnGJGukF9
F/oFhrnMF4z4Zf0t2PjYVarVIBI65gl8Cjx9abchblrJUuOVVkDvwHdqpNnL1ZRl
fV6yiMgerOO2Yb9JIAU9xVNwx0Vp7mubnLQVB1KHew6ZUH1d1qToN9aqqiBeBuAB
IJblogwbrK9bOZumaqDX7WwsAGnz+CYZHLd5u8qli0oNH6gfT1OOp2G8r6nAtWC4
XRljBbhsTSpRI/qu9/2UpNmrwp3znHDvIW3akTGPhIJOXq3prMjx9a0W0jR35EKR
gKhdA1q9uYPEh8NB7YrUt7n3jd7Q9vHyKMlAimyOjmQXMFRz7dG3xWm6BvGB8RPM
bDOPO9Shd/lTOnfCj3Ur6rzfHRiSpwmWual+Y2Ym8210oH/qqRuUZ9dQ9AagQOwB
qXqD4PP+W/cpgKVk72Yh60+xqjNV4kX3PnsKYSAcL44kKF/HtVz4ZEQ36WCLCSa+
fD7JMychNG1fxcs6MQClwp5Yix7sBpVFbu4qR2g6jicfh893yMY9aEdBkknBAgO6
geJy56ckgm9qicycp3U5+1zGtIn4T//ZM4rMX8TPOecBcjFU9i4aNaurIhek5zr/
QxNW76RaoxfKXb1+dpZ0YiiL32pEEdlYX8fDYokvaB276sgkYtYBZqJAkE04A8OZ
TDzOvZjFtqIsEDV99dCg0pTPSoNKn90ABDli9xG2H396DnuO08UTS2VN3EZkewZp
PLDlOf8iLT1VLAavA01DUSKiRNqaJYv8pJmmgEk7J7tESqV5hKZBpTGeX2w8hnC0
XeaDE4f5kn0+Oe8n2kGX1y+97TJMDvI1b4QTPhhI0PahD0PneKFxV4udS6nbKewd
nvJGUWyuZCD/atAZq4v+N4u8aj2qS/3YlDHhvGE73UgKwZTOxZUWjngy0G9TYGXY
2LEz4ZZi79RXOaK8rOflAqACgPOXexBWzwxsTrvfo+JHnoJJSqzcERdDXRg95PHA
pEjAAnmZCH+ZohjHBpeXgjyKMmGMFuUDpWFLfAdCg6wvl9wqiW6AgO0xtOKOcbeM
Q6gtCuiDUMMRr7m0yQd9GRHY8VTUqkIH2ykk7Ww0U5rcKKoeIa7KNiRFd9delegh
6m5u0ybYHs66HL+laFr1/8sjlwlVIp6Ui9/vG27T0xWNNg53zGcmKNi+KcuQZQ7J
L4ET5kwakUUJ5taq7Hc+nTw4Mcc0a66FagZaQ2FseI9PWnJ5FOQxt1IMR0I3R31V
7qo1vHW4NsHpWTNOWQg6+0E7RRxxY2DTFhUxZQ+PfCD4ezzi6ADdL2yV6k4sAZnk
h3ZX5tUV5JAfwTIyFofRSB6h+Ee+nYnGYznIdD3iuJugaoMGbtPeiWef0HJ18Pph
ZLTQi3eRccTg/aXS0ylmCPM0++cqy583bBjEdK5rM8/W9tmbQt6T5Ge/MYTkUNUX
ICB5qHg9EwY8NDfaII5RWRaJ0Hi+TzGjwHrx7VmwVRINrQeOX4VpkOleweJ8N8ox
Xzwfa/tqMYQ0PWh1OOix2wedeZBS83bK8q4+8W+5KaSwr3vd6WB9nJXmEb4cnyFL
H87Mm3M8pBjeiU/rmYW2a9q2TzeBKGCbZP56aEGofpTDk70diQp2Pyeli/WHAKaI
NvbPCEWW5zchEW5s2y1CbVBDFpyUDaYYT8qDa3d+5xClfd4pqOHTVQsquHyVOCWF
7c7h9ZW3KO+9VeNfI6zeziF39MrqK/mlRj4dP329EoHrPKsrb75g2jzju9hfSo4p
mkHo0N8fYh2Z31qkEXQWiJpzUmUbYhCySvLLPLzNC/Iv4iIHXsckV1FdZ+AQmg3G
c7B/ouRYbBM0uJj6fdXMsnJ8bTQrrfq+WG917aed0ILb+i3H3UbzjdwdoWgeGRS+
oAyUfzRfxka81m3bY18ZsrMHZZFabHSh8npCtundqpdWv6Bd9i+ZtyVxnCxQvLDe
HT5C7kqISs7rd9ikp0JooQ2snWdLUoMDDWDA4WW5LVPY2zuUIOc5HGmy1/cPKlYg
O1PbxKENjukowrInzJjwcQXrMTF2FFc0XRSQ4tWdieO2uUvCOB1BDmxXmLXA8UCR
4zYrvRbt01Zm3peZTYskjj0CtXjDq2ybSny/Zen6eIfIQ/ypnj3ULAm5/1EoQ7aE
z8FbLS4d31401g0W7+1wa5C4fEctKlJewKje3MZGshb/m6T7fdJX15zPY+LzouB/
gmt4Cc+vSN6d3CStDhfuWGkcaNvCevvaToiyN3xUeFJe7yd1EnZCk1wOhwjFQkM6
Z9CuHYT0q1R6rqiVpURQKOGckhfcVjy5sv+TF5T1hWetogH1JcYWDY11pscnyBfY
Lic4mHPukhK9OfMnI+OBuYkjHxXAVtRyiiF+xrAlaWYUTD3Q+MAE33XJ5SGVm1Ry
z5f634qbmcbvaURHzjA35XuCITc/fUvejokVeUNTo/4n2KXmYv1is+Onx+i+W5L1
aaS35wvDOkrAnqTv/b2ULZNvEBuJL93Ix8gkn+3aseoMq2ZoJmvL4fQVggpu0Jhm
WxxEDItb0kF+B4W2n2B47ZBVAFupiEYWBsK1zsryzhUEw+bccW4vYTMexl2nwwae
Yu3YlXRmH+c4jTGGhwFOu49wc8iPmW7x7D4M7CJWx+9IXNjEJdsIzqJa4iYT2Txf
OBhiF4+4xUh3rGsdN4wnabo97E4dOJ9mtQFwXKkXuZA=
`protect END_PROTECTED
