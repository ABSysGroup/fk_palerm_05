`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E8QxL+OLxpfkZQ56CIgatDxrT9yefvhQ0btd68lK9FiOccSNK+FmKwiJkkE2oE8z
9rhCw0xkOQywhqJ+QlU5WZl88Tdfvs3wJV2f73wyuwdelgpB5x5xX27012OS0VBk
OnxHQYGkK+0Y36fMmvfTfCfdydcgdTici/W7nVXGJczonsynCycFG4pDZpmdN74Y
hECak4oVrsX5dwXJFua5Cqd2uUtmQ7CaZCNiLr9YoT+5IwLVFLZUcxWC/8m4PlKL
VfTTYD0nApeMZy0vU1eCBvrEkAu1kWo7f7s0IrBNPDBryUPHxruym3x0TN1NBVcz
GRBSd3y45FQChmn45Yvktyj65LZVxEFovjo7UaupgHC+2YORe+NcBF2MekuMH5x3
jGPNAHER4W9Q68zvQQAh72AqZdCzO7AuhxQiXhGdMHXT5e0r0n+lmIWb9v3t7sBZ
rcnEHjU6Y/kt2W03SoUXA+5ooNMo02P18TafnP+sygfuid76tNdcbzO4nxstTM3Q
7LD4Mc0ONS9pUGHEj32EQUjGMhRKQJn2XZKFlVeJBGdpa9U0lStNvo0r1JKY2h/F
1yBiJWexrQhkRlYAmel7CmrgO/gfgzxSgdp2Wv6tG7jZGVpG5uSg4rr2jJy3bdhP
cwxGntAixAsr4bZMZZfn1/6OnSDRBSReDGNkyF6jXaZYnCQAENvEqJ6ohkJtIUd3
LSQ+P7ncB5rb3OzCuAF7+pdvD5pg1lh5jLovivJSx1Y9M+f48SKPB56BcfgUV3L5
vrK+/8/gq6Wryo8+TZIJtH7umxbKAWZgFShH/+rURTyz6VmoufIyItRn6Qdbb64+
yGolV/Y1+EycwrmxTkc15ESP7wmqg8DzjgHWrriZa80TkB9hgzEljOP6XMxRsBcW
rerFP/aIbdcA6y0RWazpws6mFbwviY3yskk2Q+IfDQ6DF519NEQsP0xoi0JJl6X/
IjZnzLljGRIOvBjey9Ms3HbK7nHcJiIbMVILASXQQQSk2ahIfJ6osmfblBGOyXqj
9/n9SphSYBLat3B2/1Zp6JRAiwCrLWNSzBtguFLZ7tEphlA9B5Yma2pWkNLTEU5D
fUxoVuX+MfKw2mUcS+Gk/xFxYGzWjSELuEzLbPg6oJgzx2o/MLjrbTnG5Q2VTQ5G
rYarmI2/pmsBlJ70ofwafHjf4ZY1JCZaAH2N60ZgvyP1Dgdie+4K6mcNXRwkfJag
+KUUWYewGTWscRJvutRkoCGqAs9HK0d428bV1CIY48UR9fBdUI/aEsbzCZRJnx26
5PJp4KQREgnDNATKHRXaYoHL1hS/26yVfi/BnVKuYizKmnjaTCFX/wU4l216qgTQ
n0ife69p/e6QJjoc4w+MdBCGAAp/k1ax/dWwQsMBEiSAg6wTq08IpGQ/qQHimycM
jYhtkdJ1saM5zZj4McmjMiz7iWENztJBX+c2Qnxpq4w1Smxs9hwFd5Fe/iEA9vU5
u17k/FSNXwZFxeX2yVtPFRjrLOYzA+cVNl1GWqZ8KJE=
`protect END_PROTECTED
