`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xw9UGEGskzKfNMlL/2I9Titj6w9TGf+3gsBU6SfyAfXhACawx6ivPFdLaEKMF0V/
p/d6CqfxpoI1TgkUgoX8Iamnh0QVNAoWJCtw8/48OQWGQKgS0mN/4Kp9Dd7uIrNU
KyR+bHwfiBmk3claihWLPZpmuWv18k5tcfJdD71NGV9WVFN10pe3bUHybBTbiwNW
b2OFAmubilaG1qbrWA8IYkYZWBzxNlIW7JHIWhU/83cTwlfiX0kNpQolBeoV/QB+
nA4rC/ikRLQkwiuH1B/6gRvhvepcygivQm8e5eMx8hfvLP+ifrw/ksPCFLuKTw4O
GPRBYuE9JlKaxiBvkqAmSOOGqQm2dkW2lOOZ1RlsmotmDCPFrFMTK3HQT/C1zJUi
XZmdEXEb5MXrKARdtCcNFKGsWTVR71sj3/uou5T+cLrcP40yENma2B5d5PFVLMry
hI4j06hAvE34+/P/qdOpzHbqhVmH7TqGAIUk1xZmW9qs5MxWCkggSCmvNQ1Oz5A4
vTtvUBr68RrAd+tXELkU9UswxRaTkHA47GCL3Zac4bHPRbQCb4HKfQrbRxwB1pj8
kUIbe0Fx0vq0kIYVOqkYY+XnM0EilZxGtdiVLTCyDzx5cdVGyooz1GFndX8ovRqL
eKlYpzMpkju4fdLoeSi8p5Cfd3gbnjCPdaf8N3tiZhz2BY+rW66pcd1Dg1gtTBY7
xXUBBMr+tUdSZ29jccUKgGnu0WC2z/JwbQEVoC+J0Ofac2xN8CjJ+u5aplJE6bvI
p7Sz+1CGtYCSfZ88KT02pTO4GHoqh13RgjHDaM1qpy3dWq3gJ3Cna8SF79gRC8xS
T4RtHiok7G/hFfuhQPOonj6kPVTWZajDdgBS23bJGGVH9OY8KkBSoYsn8sgwNND+
M9iLZofNz4CyoOlFPcnTFV6iQw5c+yFAIBJry9PzRyjxb++Uk8dT7ChVR5kqxGBd
fpUgoejqMz7ykS2Pui9DPAVn+gJM3BYlfEtE4S9IU8zkHmno7mvZkMZm3I1It/nH
/5p6xXmNNrIwPirkVoull+H9h87nUUk4TK/xfQtC9ZKPN5Nb9BAATMZpWIRNLO2O
xAnQzzybO2Ej2+6nWQ4GVch4Rau3mnygDXdqiO3QqMc=
`protect END_PROTECTED
