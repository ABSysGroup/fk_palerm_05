`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H9qF2mZ288QY+FKydum2cmbbRFHyQodVmoWtK5Bu/3TP8SdVIS1oJSplFMR27Xw6
Qr8IY1eS3do/URXXrvxYHSCX7lTRnKnukD7rWhuhK9KEjSUcipZlw9ZDWSKx0If8
fyX/sZvJ6GtyUVXEsZvFXt63a28uGljhHQ9U/ZFaCd8j7Ul0LGOszq2hnEp3fLHE
kgDPA8IiullBb+7+SqTCiaBPDegUZjQfNrFDonvM6224fpIKEov3iL5e0ua3u7dA
X8OcWiVLo876/yFZJuJFMLdQtGE9FNZp/BS4420qwCEm4tZt91vFv/awNbim8ErG
SOtyEEuIsHNdX5xDgKHmnulHNZ1GGonjD0g9CfIVVHV0SJSVlmkzJSIAhHZYs9Nq
/R7XstcgR49LXcNs19qfI2vKxLVYN8Cd90+nCbm3CMRpp5+JWphwJ/kQ3/s8ANbG
qtU/PR2TQqa+8KcveQ6Fq53QoJUjZPHZG9EACs7AbG6Y1SEE3KoDrpbyAV0b5a0Z
yMVxvBQGyJHu4S9JXf+7OBv0xJmWoDwsYRPyWUzB15JGcWMDyyMDnXBUreq8F68O
VnHtT03Gx6uJgWV3XIfuAiL7Z9ShURUdMx3tgs3DpVEACG5WJ++QuxaMiF9G28PJ
A2OJ5lfNsjMg+eBqhQ3iiITjczagj/9ZuuwZTvOZ4Oto+gVlNj3SKaVhAkRTDBAo
rDNnLEBSh0Hndoq/ZypAohxg+1T5xScAUp886bDG9txwMrQRQrKDYyb4rHeSyqeZ
jEQObHUIADYDTNdPzm8fLeAnr6jKS/5gyHKY2kUYvYWMVpHzGY6cm3yeR5aX7d0P
FgxsMMz1cRI7E+ttXUVKbzfxtc8Rj6+hC1vr+cH6SBoZiI2rim5d4KuS07pKAa+I
qI/Zoh57JCMF9yS1fQ3Axjz/vRw3CV6HJfpkjWcDj+c8PIHwzzj4DyBXKeHkWJqE
83kmbt84/HZCbRNrNAfYkRVXkmooZm+xKT9zmWHcclCmjzLJzAzoa1FP1JvpNfOx
Vz7rtwR6e6mhe89t0Sa2Eq8ssFatBM19yHSGobxe8WDi1b/gsrfB16uDkCL/HpSY
uxUOz7ksPXKylZ3fPEeHjR085RaYw3fqeC2+obNozfskCUrXNPTx+pIZGHIa93bc
zk7zMUkr3cFrYvES+F+vfmK32Q8mVLYJReFx3ucl7SlUTrO3+2y19x0T2xrJVjtF
bbqrLAVsz9my2fql7jp+7mwFFOLtCgYyHNoz2NbIsrbRhRtJAGsJyEN4RhU1NE3B
SLRu84EN1StZ1iJeOPhy6pzN7X5WqPdfVnE+rLpmzAruQd5SHHcG6uRuWeQLDLDt
jXI+AJaKA8Be7Nk3D+tYot7R+qzU4Aag/kE+tjW3QjE/JhUAmfCGO6H6F6+2jAbg
ybGDmoNTV6sc7u+E+KqYNZfrfgWdh1H7/RdXYUSCgZEUfbQhRpJdghaqWLvpO1/g
WTYFATd7Hs4R1LxtNNnuFesJNb2avBxeeA/UiWe0P80/p1NFkNwYukiDjA/lGXDA
MNX3sg0jpbnO/slQBXP/No2h091KjTVzNVQGzsspU7kEv0HVdTwrTDVa9AklI0h3
9eRVrSY5DJxAM+hGSMm8TvrAj70pCgZvi5LQ6igflUsO+bwKHyy/bnht8eolpi2Z
UNsgtFj+W4+7JV589cC7K2jQFshXQFbSkFH2yeLMtZy0MzV27AX9TiMgB75Q/q9M
iZC1KYg4hVf6VsDvUkWuGTNIrH0TH0fzwfzH0RrC8+wGZ/AhV+mGC0c1rx3Iyxm4
/1pZ/a4kcTpEgvMPs7vgsfMIYXNs0/Z+GPVhAPoxHm4idPhjBqdDgVqIF8Jil7AP
gqe6XeMlnWBD+eN4Wo5Tleh1DiU/0m3ikVssiNiD1bcXO3mV3QwQlma1AscVe/j4
IHmiaVoDglql0FurYimpm+a4Ih65LdenH9Snl6qct0DPXZT5iTtPuVTBQbo7UwQY
8YWvuXFsinGJf8hR8jzolmtgt9KdVtlqhc1uB3Obj4oqQTPFC5Qk86WpAowcF1tl
NjxLlg+2V/1iiMG8/2uIRfP+WlxtRf5zW20USeg6XPxpZzDr/fVzyYzVb/nY7yg4
yYjFzBjCmYVW9KGA9tC1qs3MoA8Jcm2S79VXFQrZiRhOmHCwfHTNpsiSIiKK/vYb
y7JCx+XHmSXj9hlsnmFJunuHK+KEvQERjZ+Q2i8IbqNaYsPJtuVJJrtJh3VsbFZc
fmMKnsc1pT7rGout+yOj1RbpktBkOueHYj4y7UqOVBakpzVXj8IuPLULbjUYbqc1
6k+alDjHpcimcg/gkN6Y5/dzCT3wyigLZXHxvKw2hKT1QKzVAG2MhNX2DVqxR9H5
XcyIvLnYDcDG65h6xOeJVwW/C454Um6RrynRuxKhkaEPrUro+h24EJQhgrrOE3t/
T/u7j6Xg8NygyDr92glEo15JZ+yHrywc1ZfPv23rhSZ1lZba09PD9OUIJ8mSUGTO
Ty9J/WT8gyPVvyA+yC+wSRo35qdY5Fb1L4kSZJlzCs1DZg6+2N3Ke3RUZE28EPUf
6D5SMDOQFKG2QYofzP3OuY9GnZCoJbfgJXnI/xig8zcyYB9UBjmjJKR93lHOyt9D
gfxuqUywwNGMlbM5+LzhQQg93sgg3DOK3+2NYEgxfRWidVF84UE2SlclSd2B4Ldj
2BX0hGNLkeYkbmXURJ9S5+Puca/l0IKm1HtLa92UJvmPtz3WO7XzL4iuzgNQmtDo
frmsxAXGLafJHuBYSpjvx8zom5IQ7Hfak8aM1jo06Q7kZQ0S1yxGyfXS9oIc7DwW
wcLLxgOArKqsuVW3Ak0MOZqjvc/iIDq7xWqJk1VX8e5hP2r/W1wLvCLIqqMeLa/h
Vyx4I85nEXZ1WT1MrCG1mw==
`protect END_PROTECTED
