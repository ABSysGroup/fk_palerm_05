`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v++Zy/uw40TwvdncOZQhTlMrQdhjCtewSVRyL9UMOlTwBnEu4TBge0aN0uD6DEaT
E7tgS2rmxvsbi4AKXgDLV9uZUFb6VMHX6fwXlXE5wo/7pGxE76ua6ZiQng5gXzP0
ayy3yoycXWZYRu0GzGIYvnh8Wyp2QZsHpl3yzthvwvhd1VtZ855nSOaEydLE4Ti5
qWw0vaQTwBCd7OVmns4BlsvtfJAze0PtdGRWRe+rrdoSsNa4wHWYPXGsQjLKvRh4
qRIV+yt41ujChNqo6YjQXX8f7Fvyez9wTC0lJsKUvRbCEcF3tkkWwwJU9azm36Bo
tN03/hnZb4OfO1Hl7fgoVtvuy6UsgM0NIZC6x01kfKW8sHJOirqnkV9+Sg97EXv0
cP8H+eFpDMVxgb0ItI/si0cRW7JxhMYivvTPeSYZeOdUzfDNd7WFm2+pCoI3Ryan
/4N1Cgrfskd4abL33UXNuPi0QUdozv+okwAucsua9bsVvraLyyBpDe6HuJN/KrQ3
yPW9AFIFwQHJCZ9afYpVG70Cpj/QO8SjcEzxQkIZmxp2BpO5Sscn5DOBfHGDVrjs
//+g6LxjT2sOJaoBAA/+HyOmVtdzYUDn5wgnxnRS3BpRoXRCFpjF68xE7RWCLxHt
/bkeazfc04xM++B4xqFJMB8aFXHsmkdrI5iGVst5Tn9ILqRiNzccvsBhjRM+BjC4
70waag1LmWIeeGFlfSl8/P6ywihQKw/L10CIteu5kYnA/1k0NNESJSfx1b5KT3mx
Wq+RdzSlKc1sLfYPxBKhU3mvteMOCVoJJTyF1KrcQ0YTprlLqHsps7nmSFVDQvSx
FGdOLexVQIDUsyLFFGWdztD21s8IUooXoZUmskKVaLf8SI6TkvBASNb00OPg/ISB
HZwxIg3ucK1XvF690/kFnD12wGhFHY/TbxEhxagMtdbnlZH9aD6XA3zosRqi4bhD
chNhm7dNhomJf+R0o26iFMj9m0VoxbvhMCJDRk1+QI7jULN9h1dLbPGhaWXKtnV+
OdjH0Pswd6rxSndy7ulVNa/OZN3OVaqWuhfYd1hdBzksSidqfcA5wCEvRaJ6ie0q
oceP/DYGJ5YVHF0p5+AoBPOZQlZjf4c37FoUpMlG6sZxMxV7M6jNE44HWyCTeYBq
n4LgW7GB/8k0cManVjQgfG/QJTvmWKL6ert9paEkWTmMmZimONEiGCdgKmyujy21
4COpMl66X8mey9gBsWpOR9jA0xThMpJexFTsvSHQ1dMDB0127uvD7akFDE5uaEEz
KXnY7lUZO4ouYbh60GQNXp70VKRvF+ZsZCxEoTIdyoxXvFIKqMUBoEDDC+ud3adT
OWK61vxQl3k8tyVAY5scDkKfUIvJHyr/b8w8GnJCjrCtP4tPEl+ZXowI8dKSst+R
p2A9YRnMr8X8rnGWr3sAXHnh0CvbrHwbCbk2ZB28XsUzAgv+QSsK8sxclnbx372H
z0XSRClOI/ndrPjAaPmtY5ZqksRmiJwF+4xABgirmA4j9rbDHQFIT0CiZbOK5qNb
LFHXKz3iTD68ur7bb20qX4E8DHHgpyZp5ledgeGVGrkWuOxrPwCynNTjn9IqD1y8
27cSjmFVGdyP2meaV0WTWGTGVgsIpJZBN2H6bfNwlhmLw64rpX0ZcqIchllGliGl
S07yQoRs8JiHpk1NW/JktQGACO4bz3YMu0pesXS3asklCoGZqJ039LBfVWBjAKYa
/Hs4UWrw1YXOVbEdduzESXg0FI5uRPAf17f1VER04K4euha3Kw+KEjI0uNYqnivC
XnyZDXDYy7Q+qi5PIR74XHv0qBCRGigG84Z92zzTVdoU2sBbZIcctHLQZTmk3uPR
zTWrYSQWU13ArVJ1wseh6ksSoeyQDphHlMhNI3tI0i39EQp5PO1TiM42ZE0OlBMe
`protect END_PROTECTED
