`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+OFKCRPLceLTWGZwyZMMMET8jLwgFuDhY9GSJoMqBYo+6Gsb9J69hOuKjagWeZ+t
Emtyr8uwvF85Xg89ChRh8WeWH8xm2/ikiT0XQUcu1xqcMUeAk9xPpTWauXz7TSV5
kDMm6YrcgZ6NYbC0z35bdW8PBuIH9WE5KOIU0z+uPKQGtC4aJdOnMnNtoLMq7W7A
52ui3BibhvuVcJ6oBY+GTzYNXnsde6ujme8jcFv0Z7Y/1ypVvzYH7992TbULGgDS
OObMfrb1d/dB07EM+DwWng2+Lvhkwh0ae5T6hjKJ2ns=
`protect END_PROTECTED
