`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d2g4aTOxnPUH+Bc9uoagT+moQ6aDrzaaQphk46pGfRgGQ4vYVe0JexqbDNmVts+C
ppJRi5dOV7eejWkPvxcBWUvlJClNfIJn/s7Lrmsz8i21I2vLmqGZ+HoYEhpUlT6v
RmKZQmADt3udRDHNiV52J0gFTg/lr2q/GNXI3ByPLWcHoWQUFAFsMXCCFcQqxj80
J74SNWeRqXkS3RnJA1DYCydxUdebpFh54Rvs7I911T0D5bsL3miLoMbOlaSvegR6
l2wLFIe2GreyHMIAZT01CWjvZ4kvTygKPJioG+dob1y1eTAChbkMU4j22UeKQJCE
P2E6XVYxVTZVx/ho5QKUdrVQP0bHE0RxV+tOqy9ArIRiLN33OZacKpbZ+vkghKkH
4nNwR0Mtwh0fCHvPMEftAVgTt+4LRxg6nGXvea/3E2w=
`protect END_PROTECTED
