`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gNodhK17WNVdJAsH4rpEwd0Jn4Ro9prSQL/mF41Awt84FSakY+hBuCtg8z7cJOV4
tcroUO3OeCmveTHfnZbxq+JlGXhARZ6IJnIiCuFKnEAB90hh/2OQxcqfd72pqHfa
3T9CC95MS7sJhBh93V1E1lnV1ta06I9M3k2foNgVw9LlBvh1H760MSgu3cC9BWUe
RK7wb0/QcHyJLSv46Z7rZloBHWghroeWTaQEZoVVwvxeHMzVUoIIiqpZ8Mz4TmuD
bF7XC4D51+UD/q8VJowdw2B90/uVGIR8BR23T9znSiHEIwa4n6uR/m0y/hB1UwJH
i+K5618u8pCTg6kRZn9J6zpN18iywVTpd9yA7zRGP67hzo7bFBqErpM83EYywd/Q
Vg6LTJB/IkcaTbxAVkb+G01o4LV8NQ5Qvush0H/B7sMOrMWxMOu5VzXP/O+RBEK4
eYNQUuFRGaX/dL/l+Iuqt+yXKJfox8GfNMBwdv4ZPEaY2gb85IThBUJsQh5Nnj9c
/dSfBSAOTHKsBerD/cYgm8izBQ2Kgrpw+XoTLu3wqfNWsyazysfY1di0dN0zaWHC
Sw+q9jY343cubxgiieV0GSkdsZVt7ZlyqMqxoKAuiVzfUgq8NKVo9jAyM/ey+qjq
FJ5fLyg34t94/PaS/II0sOTvvB5F4BaT9EQp4hrLVcT70hTHlJwO0ThrNFKiGXxz
nLyeN5GhJBOew73sRXVpsZOj5u4CCf+cEwIE1KW7K0YVu6DcanV0V9Bfc2Si7A65
1kI6UCGDlZH+EkBmXx9HYA18pxVrJF7Vq3iZS46dKNO1rbAlsfKJeKOXs7qFk/rG
P4BsNHj/ejoM4LHSo3DlFOot5TdEfxr7vfTTMc+YnCC+r0LhMJdEtGxkbe+OTH8z
Y1JbjdR0Jeh3uOGIC6hhIYMSkESbpj0WrBg+5fJSPZx6/wX5/XgzBW+f3Ublb5Cd
MppkMziAvlvJNyiyHUw/QxZtJhadyLX66AbP7rRxwtv1x3r/s3YIUPyr/IkkQT8/
K7j5/S+9xXZw5CjsXkXcos28qxNpN9WOm+Ho55OE4x4ORgVo8GSDUF6vPPEXaoZk
csj/3ulIPnqK79XPhIVtClZmv339kPLdpQKO/c2DsuHPa/AmuD3ejO+WBMgAOQc4
IvymbeUflK1qG89eZjesckTJ1aWuqK6kY3mhlhfIAseNdtoW9GfWPpYg1aYPs67f
xykyKJpqcrO6UP+swg5nPA==
`protect END_PROTECTED
