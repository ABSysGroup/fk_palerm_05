`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k7KcXC5DutixWoAG91HlNA96lFF1+YqiuS6Jj6IVGqFF2icGal6XbOw2x/LYOpub
i4VAJz+3qL00taHGnjXPRQ/i4HEzc3h5JWydPXw7fifiijpKmO8nZTOP1Sos69+F
0M1jlZCX3AJPDF4YwFF53FqUXiU2ItmWcmOHN+DCobjnuxrPRHmgoXPMFZNgDlAu
/PtIeiDZGomZkDkpamImPVZlsfZtTn9rjY29R76y0og3Z87yF7U3tgxUGMEunYh9
MwBhsVD0prNjD/3shia5nQ==
`protect END_PROTECTED
