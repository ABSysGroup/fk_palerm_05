`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AP5k4AJqkOfRw938e3zFrK7LZ4wVK0FKs/GoN+2LQpyZqlt27D5LxkE/8cb6N7jy
eOnYcaWOb9r3RtKYX7UlwC4GrvY+WpunzU4/Fxx1fCJSo2BIFMEZwDvuRfYNVMxl
/fcni/9/T1s5C81njsS+nCaD/h5AiMXRqx+Gen0HbjP2CGrKCkEO2BIezLlm71Uu
EMBJMapl1r/UXAbKZ0BwzG1wpo+9DRfo5VbHfJtmIn62Y24ezHAWYQOxmVwcxyHG
HaOwq6ObGNbXL7tlfhJVI6CaBXSjs+k24nc/OC34NCK4exhIiq558uc5kivnyPQ9
JlTqUpHf+9FzB0J6nwDI+NCH+JcZdz8p24qPwy4kCWPboFtZ3gV38uWNmHRqjOMc
PohuE8egwuch7S2+oNd3HFtq9KP4f7kwEwtcDVcE5ZirI8eL+o8gaArFYyhr+10b
oJSSCUjjWrsyVBLHt3trEYJHnvO94Ei6uFjdth6CA4b87yX5VX19++1VNmwZQyDb
UHO4EOKIeyjxNUsu0Rcof9DA80hCEOYt7LzF+SH/KTLsvzCdOrRGU5fhjJuFBl+b
93Rh/AUEXBcU7KG6JDyNJ8C6XLbzNFR4r5jJ/wCHDRFrwvbM470jcE+TKDBaqCgR
ifKxv1JKc/7FYd0WtoQlLZB2GdCfMovWByuJ980Lss4f1arbGClUpPOnAWn/5bA1
oGMyhy1/NhF0v8fFgijnoPV+E+yzw0pgjDWpm6FAVYO7F5xqUvV71zDBWz2RbQ3x
kYovtAbKJYtDoA8n0NJ2R//qRLd4OptbM+UfqqLtWlMf2dckIwDQ9TqeKU7RZWDx
Cr5z38ROtuVpXOFEaseQZU6snLyvkgONehvqZkfOc61AhtrJoF4zX3an4/a5YcYC
Fx5reF+qBYONEo5Yj31UdlxIMkRh7OCL+bJ/y5ePnHkqRFzvgapn2q/UtA0A4az8
sJp/BmTgHaOU0XU3oin2Bq/iZ41qzwuZ/SHd9wcyWdASH0Df9tUrXhmKfBGRRynj
`protect END_PROTECTED
