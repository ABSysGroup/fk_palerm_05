`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P12owb9lHivlrELJiVCFibvXntYWR1sGQF3NBx0mRCfDWzPDHK94UgBdWHg/o3Q7
9MPr0Vm0OjTYeZIec/HJzLlS4ffIE8zjfzi4Ga+LNgrg09ygQFYkAJiTlnXhAiiP
y1E2vhzyf78JDivWL6qVi4zwkJH/04P1pZocg2fXAf6GylND03c3Vf0iFeOSLBsA
5XZW2iKjHArGkbo4uGY7QnwKuYqXOH/xyeN+Ekg0ETDw2V55ngKXlvB8gZ2f+8Fd
v/iTXqydaDjJNogR1W7s+Kv9OPFMwBxGwlaEYS6phFrNYYUxfmTegg0Xot/FzMgt
NK6mJ1hGhSBeVBIqe213g8JPyI2i1uJtf7UKfBlzsAcES4qUIosX3emv4GXxTo6L
4PjJ0toCbiln7tOYwsHLlk+aeurqmAd986h8bKY6CBJWn8nzpyYKaEwmMJ4Ey2E2
mVDiyClLKwuZDlxXDBOGcEnvzGDVPMdmisC1XoSW8nExYabXjFY+7i7Ged8y3faY
h224p0pomqjZE36UA1gBvhGaXDuPsXs8UCoJG1XsJzx3rYrWcQD2wc1fs1WD2irK
YKHDMy7qXWz8E6/1NliiMZes7GafMU9nTxooNVQVgSGDD8XWO6ZmcvxnY4m34R2p
KpVnPz1HO9w3/ppLNsqBCCdkaDz9wjGk5heFpLSiQCg=
`protect END_PROTECTED
