`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Esrd9/Om40zWdyWHYcqdfUXd8KcfmXJI+o+5haTisj7DnA5oXVLODsotr+QkbmY
/rc9osuJJABO7XXOJZkRYgySNOjmzw0eb8gCmrSjEhiPV5QWNyeDMOzTj7PYDqcN
i+EUMM7csvkBtO5ZhMuFfHhrsVGhWRDzsscO5+EJ46YBaawfYqymrybBhoeRKRgF
AM66zYbTdVcJHiSSo6coyPXg/yLfZTQ8t0I1MOnkhaQkk52HJH73VUd9D8mWTQmw
rJ8qGzkDunSKDrynjr8NLY4VmcqAlXmc/+r93DhsPCrNVrZxPapYjcZk6CtkMzBE
`protect END_PROTECTED
