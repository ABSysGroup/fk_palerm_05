`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MEjuPDbcY7viApTCEbPB1Jwm/M4J4aF9hMmjf0us0XCTFWD5OoQNnakihAgub3kC
N0kofGEjzVT7USwVHNgw6ciGgkBbRJKqCe1TtXi/gDvMWT4FkrWHpraqJrPiQQ2H
k50G+wRUWbs4s/i/IyGoE+iWptDuEpQR5avItAWWYOQZWJlZlImWwRRShhD9GkEO
u3bc3mLnU4RPwiUaIRkWUK7ltdtndREy7kunn/wZWRRxtvSL3TPiYRyfdKHzATph
K0yIpbrm8SkgT93tlt3Emt4bC0/GKfchasu9g+OBMyu1ZiqMd+wjj0gbs6DLHRuC
Yt+REMcDf68sxUCfCWn0ElK0X6VnLTy40cAddxctBbzTf1Px6LIkUIG8aqFlLo0c
RwmlcfC5Qj0boS1UxgBnYurhR3t3meifgevGu5O0HYAfFnHCqFuc9AbpG0N3GJ2R
Z7bQX0cveyz66PMBIcVvAF5MH4pJQwacsnqqvyAQNA9bwi6iGao34OtfaNkPm5zI
AnHQfQKXTexOluJ0ObQJVlEGXFUh703MfEyY2z61BqjbC8/fczgdDb3oEJ5GhbJS
0cYcYwbaT2b4ZqNxwk8NMALv0L35s/6K6mM6eVkV4387b43PXRp617uXXBPYx/pH
jVhxE4AWBReqglTzRAhe8Wjr1Gez6ygTJvmNjTlQBrhHy7luMLeRe+O02O1atOZf
HZangFncJ6aQkyJitERJS/8QPPIJmPS5P5kOoS6K7uT9UWLnHIMDecoryrQ8AZ5x
9mWqx9Mv3c8Sw/Am6+H1IY3I4ngYH0WDZkjEWI6236Kky6izGk4UuoiExUyByKdQ
xFB1+tcdZWLLzuGBQEtRd7v5jHRTlQTfaHjwN7qXfRxmZh4EcYr55Ms2g6t0+x/8
7P28s64vrKO4BNRFgLtDFfWoJ6oy7VeFqn8GVTSPN90zQB8OuHpTFOMA435Bg5h/
`protect END_PROTECTED
