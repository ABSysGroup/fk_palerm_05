`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4MrMXDqgql65az04pfpyebZGDc4nAk+C73ju/4/fjPQJYkUO5xm6y24pdjRTnpg4
pjNfr2qexysUhX2uqcmbZJGJXhSyij7R8e5gOgYlZGZkIGxtp1EdbkNwDBRILnPk
/FpkCTUfKojWPA27ibErJn6YnNaLALlTxaBlpP3zOJOESsvSzDx7j2b6fP1Rq+nN
qkKP0pKeYoQICAFlWZ6U+oGo9CVaqW37A+mEpfFrtGldnAZ/VZLEQdVsWiE+OgpH
2lGhQX1INwnhunGpuSnRJeE7PBh85EzMxlQlAe1FlrPkhGsKvDYbXUIu9nF9VKdP
B7vP3rpYP2frzY+hGas9ds8n2tIGo5pCeT8dCrBRYTGC4PY01dY3jAQqKGx5U4yP
3wp+Yek0MtA6+nXKUH1CFU/3CFRaOIpJh+Yp4b0ZcP5WJBy4tyC+Iwcb9N5M+uds
08gQ5664NfU61PN3opluJF0DbY3CXPGJ/t6HX2dPBtS7Q4ro1/VokjNAKLmnD5wX
m3chHVROlEDJlVue2IOLpD780flVs3/1QJppH+3xAeqlK6DYUGfKxL+bBPArD6QX
LUVZ7T00al+ov1lf+9NEyNwZyoG8dWyuvkQ6G4JdVe7zWdhonqF1pb5x5yGE/OKe
wpVA6dptrm3HCzlfoCabj0Dk7qKnOMhOTOR0FZwy52gKkq1Ue4ZF/kxDOorMqYrg
vcWm3KP+OsITu63tHwoxx2uPY0Wl8Ogt4E1f4swCqvQyGpz3ztHrQ15N1VTn9F/a
2HZEkj8BtwGrIBfSvHi3wioMQgxzEgvGtCyhLKad2ds44WS7e77EGwMEFV/6zhyi
0UB9uD3mWboHUbMpMOCmFs2fVuwMeksR77F+2nm4Q7tgTMXynMFzxItsBDGMdMWD
rDq5c74os3dKna75Y5XTbXi51zX003Ro9lSSLysEy4UX28Wu3D2iSYVvdr3eP+CW
pt/NCgg7kwVzVifdJobEdvlJPaoZlLp57g+tQE15Od4XBt+KGFkyFBvVanlwxLW5
o+LtF6+WyVL24M29z8qp+HWafRnocRlBR72thmhYWvAO04mGav9SG3SR8SPS8Oqw
sEF+QLh+rupJKfTfHNfEy3LEGUxKzykGoYeRjHUaedCE/XlZ4UZLmRU4pS17D7z3
jhPqSqvyYt41jQc6jUhIGk3aOSYJr+2bb39e/ZjQLKiJYMRLdnrLYhE35NqocK0M
e/Mbv2tjMxJR7ya9DA988N646FpoMpTs7OmXsQxFuqgeVjN/B8e18O8TXbJ4KeoK
rwFs2gL2DGpz/4sceibES1yJo5feknmgdIddYBGuyNxSGHTzWjPTUtCJW87iGyVo
dNB/zoTNcMCl/NzaSzSUsOvcNKz0h+re4qQEVYBpXZ2fKy6GRx4s8Gdx6gdGEMeH
4JZ/pdIrNAs65E1zRbfguHYoOhJGkK2nIABlPd4f225ymjmxZ4w3QWqLzNvAfejm
H2OZ62xUjG9hw+8ng3guSEgCNUls6yeGCCkdmLNMTkX/U8BaFqw0VTrdIDaFRUFZ
RAVBtMfoOw84x6hBQvrWC3RcaNJetreqHncyRgoM50+8YzcbPktbJOF6/Z7wxzK3
EIcE5aKSw0FWgZ5hf1SSXGWuYuqYMbkFwy6jikgn/Vg2LhznEGw9UNK4EGykVI5/
CxFEzK25yyLndB1jggQIeov6Dv0baiu1QnllwV1QoE3PXDYx3sd7vQwr+fvNJtX9
kAdS0gfjYbe/3sRvD7Haqz9LsRQ0i0txxdvDXTO2gu4glO0Tgf7Q6IB6ql2fSWgM
SoP+hH6vgri4VKSU6foN0QFX5wPvfGzb3GqmRKHo6A5AiSTKTQlliQFPzfALSckb
dnL7MT6GwmlVGDFj/13Rs5zhqNhGPALBseFTzzTjwJMWJ3+lMU5MAt0hdUfsLN1E
mB5Rg5gA+y/+n3Msy0uVol+RkoBGYMjN4/0idSb1tOu6qI9ulGXppwD3pLpP80Su
E/VbmX5MdzuAM7NMpT/RKF+8as0KyyHkgw4XKMQ65rsG4JdOy5yMwMDUYXnf/osl
IN37oFrASjiW+lDWI5sCEIjLtE9FmrPVoUKlOySjPimgt9tVbpW1uLb4p6mshyhP
hHB2+wpIn2zL6+YZE50WtlZrK0+Jgk0PsN9mj1D4q0z0RruWZN+crv7cuGU66V3K
YgNrYmAzWaF+3bSXnAwWJMvsB7LnKBBJEgicw0ZDmdOFLtUn9cY23sSqYnEWgNj/
RxQWIq/waYowQCyUbf8MlsBex7bLdqsW1Qqx6AjRi6ORYUbT5IscTysNUras5Mr7
JgZXb0QvmLe4o19SgLRLIxlLIGKIxAmNvAJZKlFH8MtL5T1geD/26dURDZkFjff0
wAZK/969Eoqy33PiHwXsDDVzwvLrvW0+NfLunt2XCKVIoaMfCnrtu9EVaPDovdAt
jsT0Gt/YkWovEKEPNDpMLA==
`protect END_PROTECTED
