`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HdFnK8UseNZ+nSArtckLTXGUU1GMVVwqYoiJ13cDOZF3yByibHglC85ly1I9Rl7O
BzMuGBIOUIXHig/QJfLoGPbPp3wswQuqrbqBDF9ERVWGtwscAvMHEE0vFebnGi20
fT5gZIJrTPEFpN8MacBhAr2yMULnJ4+G86qY5pxKx0zG3z3DuHQ0uxhrt8kklnOa
MvnNywuIKKZURzZATRIAEn9DxSSmccsQNwqJnnc2ZQ/On4WvtDjOaU76U/mweP6Z
vLqjdApq284KTZMvq8fHqnkcAAijxlbWwoTJx0g7z9NCEdQcLRUzli61RJ8/DJHy
3nDgXZTek4QP/Bl/bRPRJ0b3RDDBKwq4s43nEqgW2XMnXDFuaMWENu6tEawmSGj1
+VeRmbild5C1+qEwj4hOD+bC/CyyYKVhcvzHchS+ppbM2C+g9U9IaPqAnP72zRev
b2LYON8cZlAp/zu5eQ9pJAT/mH33hvKeBm/6HEh7VS97NI7voRKY3Hc4v8VIXiPh
+lDsUEdlGDZlVTdvoi1t4bvESjPDMSrvStUZtTJiCdPNhSIUoDB4LyHfg9+tDxbV
vlJ4eslhqk6EqoycbMI/ChVeTDby3rfRa0S9tcAxMeKILeCgEuB5JL1QzRDAyUc0
sBldbQ9/HjOp95DnigIHSwYD8NzRDfyNehxPbxb70MDjRfVmQ5C8q5mZ4/u00nTH
3pgEVW/qDl6zfOH72QkOdzGATZTCvZtOdytBdBI6bP2mgTQncbIEEWHMTHmqRw/J
ekOn/vB9q+649oAEebrFR0rjzLFMOOJKW7I9YtIzWvHdOH3XGL3KrzGejNWK6AGQ
o5sYYwMZztYZDpvyQzfnXq6AOU2uBqKIIwEsZwhzmoFM/5TqKcwsSdCGw0p0iV4p
LSBiVfnkz5+jbAjxEMLH3cECCRj/6qY3IKPwdinBjWabXX+86ql5vdMCCtYmo9nY
cz3n9QtOfgCu282rwpuoNTWHWfhmcrgXONwu8ehrxX4gaRs7q4nZcYj9OFxAp8g8
S5/1KmFspG7ZOJaffq18pa08xPio50xy6khtOGD9aYWSYv4R+yIrxD8RiJLC5Tro
m1Aas3o0kAkaO3DFq2hbW2CgwvQ01XE3U9lOmmGaK3pJzLN1lKbDUAZhI/kXyZpf
UQZFk4ZblQ5PTqH66ofTqQYVK1Dj+/yAO3f43TkN28Uxml8U9Irh/J4f4ees2bHc
LzFLCTKEcscFkUZiUQ/eWvTJuxOs+zypsWVIkmG9ERR5iUqZH4/xduMUjgbAdBIs
qvDqhlwt4vsKL5/0sQ5DhH4QQDRFFkZRq104CST+8rAtSAQztBZ1V4MQlnKRIpua
edEc7aGfy8IpCyLjwAHuTdmqwnsFE4QCwkyVPzfJ65w=
`protect END_PROTECTED
