`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bvz70LNyA5iVCHAa/uUWCX1spk0JunfU5Es7Kjxbp3XyQFM/ilXhHzB1o9sSYYk3
NfBAsiDc2o000vaFfvD7LTBVHxlFK7+pbgTpGTs5sixlqmHM/pFKr1KG6usT9XoH
NVYtyWip/qpD+vJDwBmuZ7Egfp8LdI93DFml3dzgmYjgEFJ1xnU71fPbOHURKsob
qF/gRYzAezr4dnR8c38cNgaqJRoqkwH1ByEL1tikobMIct256jNFz4SxlIZmdOXw
/pHX/YMMDXSMHH1GUIRwpWfH1wN1pgKOUgWZfBLpmnR5gdMPVtAqWrGbP1v/tZKB
5U+WK6bkkUTqIZznjkQnn+gwvr+DxG8KokZSdjZOa/aMuIG9/l9nrsOl+WAvx0EO
drHRaXmgL20y6moiRFXkpejMEhPkI0MdH/WfvyBzlDUS8ecCZ9nwzPxxejS4BQ+R
O6MscyaexF5zFpPoGybENyDeRIYw18Jd20dqrxT95LO5BjzEGLuYm6USP6a6ebJe
0R57BJunfDV4zjOfrJ+HFpd2IwGOMnqbAzSmOAXTot050ZkGqjxcCU0D0HWVWw2J
mZZw0vFgS5plCxh4792auqGEhzFlxtV2ZRslvOx8I+BvlyWp81Q7yLdJpZObGLhX
qluzlxIn15UsCMriwmeOiQCC9iC9E/TNZ4g6W1gv01bUP2zD+/issm5NGzGQ+9bI
`protect END_PROTECTED
