`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xiIUflhFlOg9Dk9K9FRiaBEdjWoapGiqASAO8YV+nJL6pij/V/Dp0tb9Bx2nvqqK
OVEtyB8awhJr1mQWNJOWan65fpwxpl099WBzuz5hjC9MsYwuyPgJWvY0j/8zwxfb
jQahlMDVQSZB+o4vg/TjgI54UpR1yo8MMX2ZzWAsSL+eUsUrLRL3UPluhDw2ywHU
onEz4EyOyOMnPIdp4XOgTjNKhs/PtK2goqYGqVhm6DQOdwGKSCEt6/Fn2cfx+IP9
OYaCRwFnF3f3gRJBLl6D/++Lg9SPRzOvzyjjmgWeYCf02NAeL75Xnn8VFQ1KEoq7
6ydtiAWXyZ4CXhXP0LTTYuNuv2faEzubU3tbgxKdPn4JmFGMPZhmQxLBlVEWLFbS
N99XvH6lyfbBFMTOhcD/2fYgj/OF1uKNzvTZCczaVJg+aOxRwbtM1Llx3jaKuglm
RMxlWmJXmvl71Ao+6PoGjMPHp/7+wvJsnatDB2d/iV7Egs/g2mxQQyG0rcmzSbk2
Tuo0J8OZAUPKnQBAiOBCMGNREKTQhBAB5hmDc7bssh3XRIjvvy5o3WXRTBm9ZMeg
K+xIxNo+ibI2Yx350mbQWBM6kkkc8MEITx9s805+qyisB1ConLVXed11Ad3fqOwj
Gpt0OCv7kwVZO9alajbsiGtCT0GDXUXaOur2pqn3qfKzvqqHu5cAjkXFR00UhN6w
2HZmHCyCMgPj/mWULc4IkRiYKfp37T4NH8f7f240v7R5SK7gs9MCA1frJV3jFrYS
LaTYJYowe2WME59CKOMdvACoFPr0xfQY2EmaFZC7TcbNWmv8+XgbZC50LfUg2aIm
3+hVkVReSy//xKeV93zB1WTPIjWv0aWJz26vjdtBMzLDmiDv7qkTzNq4GhKubnZz
31nbVWPP72Fn2EgAAWRfPwqsF52qKHlFrt/eibykbQSXmCgsi6c2xYlmDIZ49b0A
wA439sC4feTmskKokTd3y2DMpuzJ+GCgFbcKjE/D/XNs4/1pGWtseKiWIQfx7nLw
GLNXubiWfbUvRc9PqcT5umUxEX7/20OSX5ZWOSLCcPx39wTiG0yJ7xlQ8MMBYLf8
IvS1af5fWfaLVYoRDoD+ak2P1JNQsuRdQ+mIJAJRSq8=
`protect END_PROTECTED
