`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mwNT0seWisoFRmsn8rhPyn0SU+sszbvE5PFd8Wvf0uKq3ZvBCdx4baf2Z46/JHrF
eDaWzjQqZkJG/g/dEr6l4zdydt6IguPNxQ52qflKLDxZuEBnKQh7FdfUcQMdTafK
3vOBizkl3+s1FOYbCRD3JYUeuYd2MKbmXTv6JS1JdmbTdZBjTHulc/f5E/Jg4nyu
szje31puF9xB1U78iGr4DmsC29YjkizLNAILuKnIcE9dPmEzuLeOjUcooHYiqkZC
LiohAK+FeA9lsDF6iMfAro9bf7KBSu705z9MzGuK5hEnW+WkHbKFoXcGNqsg31Oc
vyCsBRc9P26z1woKHM6mZtPPAAHDzDkPKfUCq1etAp+XkKllo5iFQVE+E34ONUrD
u5VRsuNsn/6xTcOZbUPv15S3H5g55xJQ59SGuApQzoHCwRW2fW1z86M3mp1fDTrd
`protect END_PROTECTED
