`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FDx/+wWyq7eyvmTg0Hl27/osZ+WzcuNNkuphVwicxT8S3/QS0TXKOJybzRgwlLqj
umS3IxNa82JlJS8UELOCypKob2mmmNj6iE/aHBW/DsurIdS1lkgodSmOhB/OxTtB
86TEds3Cf3GINCb//hQsCUNsdMnUEViNHK98WEVvQMdrDm0LIdcJagjoKTPVzKQK
BPiwZ7OTdQg/OFFSB+RUrvLAQ+kplbVt4FZcrguFk2JXAF0fE+ZHQ7U5jfo4e4E7
LZO/9ZymIWsVSwcl9sxws9AU1NkCP7m3sJ7Fn7ZglsV3CCwFPqoSpaYq2TIaoRju
daSKaU/VZkFfFb7Z+aA3y7KVvVzrGLtoBLHvo0Q8BmAFep/X+x2iZAa25SI3hfHT
1NlXNdoajPUSwjEyJI5OYBjHHg153K/ofrras7xLe/NZqU93kAhA1beFjdp3bZOl
QTN2yxOSeA6y5OW+XvPkCa2AWLpo2yXZhV8uCuknzdT/xTZt8o1ldFJJdnH68VcH
mTsKxWeQLtHQRz95nQHNjr4DYm4GG4dzZO8GW8OzjLOTK1CxWIbYtWA64h0VZFYF
NoBVlkeo0PJGrqOPglg0gvX+u7zZDHDxmZFe/Mp/Q3+aMSZ5RUfeVGQcDbsnJGTn
ZPTok/tZ5HYqfFjgne6Zmu54Xusn/W4lfKcTYKUz2yMa/P/8s3gO88V7RVqFmogv
gzOqfbViJwJwbsqFaKhVIbcS7t9mFyThPk4BNzgdRnZ0y4gcChAIaPx7oQ2qpA+5
Rr7qXJi8DXHGPVm+6ag0dBku772PEOHOsGrLkA9qdaeSKMFs2h3eYiPeFi7iqT0A
20CzKPLf4JnMSpUeXftYuy7cUe2SUJ4jDd+QtLB+g/4qQ72qQine2/VIOzxLaHaO
toKilzKVIGnW6KvjYtmp+pu0Cl2AvityVvl5kWrZW94H3y3pVzxm3RWqDzeSqU7y
KKR0Qkojz9QDIc4om+K6dxxL9LmefxutNtSwUgb1kVn0FMYFKiyVC3zRC2P9I4z7
4cZg5sHSCMXSwyvlrFayLztflax9RtiplIC5ssu1tBKrtsd/UULtvZN5Ielxrb1W
zrUXJG2v5psd6S6jF0g3QMcJugC0OF8TFjB83HINt10l8I1UBjqEMuy3FEjVoPTm
vIAo4Cr3pH5qHkVazvB2HpPVpcatqnGc7CsULtl8IInHYA8AOLe8mqgKKkmE/z0d
bfar7Vr3HY8jTQGuBZ2cMuoBVcWaJ5/9mPYzh1R+mDeUFFEJqEyD11Eo2fm4hecH
s9zopOxLWyEXEjof+pnmCoOqT7nPHSCZC5Qary66cmXMRoMUmzW+tH1q66jIHUSr
nvHdlzzSvGOeLeaUvdVgPc2Jekg36CtqwjnSu/CnFHLrpB3J85yfX/K/vRZmvyzO
9k5YdoYXQ3S52Icdw9cQpS0PJXsHqhryx9zZqi3CK3yLQ6n/rnmA6GOrI7MtcHOs
9Sfft9o3a31dYrb/afSX3eQAXmBP5Y215oonUUBiT23eUcgwFk3jFxQe0VC8O2ko
Oo5Z6jsme2DYxMcWhvxtG0iM/ryfomaf2Jfl19KT4OxymPvIU0NpfV6aD0PrcOiT
TPiBZocqqo9MG0geQEqTTMK9Ys3Ca334J/88gbL3xM8REAArjYTGMQ91Os/7EjTD
NuRxcthxgoJxsZDFP4ZQUhwNiendJWRlKQzgwBBo0KatMxh5BfruXOXrtm/zjJB0
B5rtAwCm2FDNtW6Pu3fSortKm0ImqqeB8X6jdl4FhFxFpIFpjhJKQmLsXGa22B0q
6XYlGeVTdJsNqSpZgqAWS6dNfVIABSDLWp+3FizRvTy+yCqi4MDC3dkW84Nb56Hk
wWdaQd8adljcX63CXdQBvXuTiULfjnk1AWlFGeS1rtPTDOAabWgDdRsyGvOcG2vB
ZDnn9ustOJ/CJzE5Q2LBjW3tvVTABjEUrN2CnWuyizP7QjXG5rX2t3/Dt7qG1jqV
JnWh2Fse38pJWA89U/6QU1MEDZOaCjusQyTgwKjogiY2+dBzTFHJRDsGBnvpdNZ1
MjX5kkFMElsO/9qsUj5ssR21vXq83aAOYWpEC7k0nmQVMYC/FcchzF7TJ5DOLYuL
8G9sDU7/X++3o0M7xY/I+XHBWZMOqB3laTZgVzPDXvwR6rzK7K7ig87N4QUsYxKA
+JextQDyiCoKSDRbcV1XZMq99b9hHC+fXhxk2sbq06+guHwRX1UaTvQ8qZvhFm4X
pmDUyUUMlZCdNvwPbdV+3cx8YsF+bZEOsMb33POSPpD6gSRfe1hdsZLM8Z1UHXvE
7BF9iCmZo+sAwt1uILe9oFdu/GMa1cW3Kzt+qwaKjCT3981jadCEJeFyngu8ol6U
dVUIcOq8tB9tZTmSyWozy1hkzIHy92VzcPWBRtb6EeQbguZwaXPXTqnx9ACrsfs+
U3mzAG2UPeIUa7+6eYhCVhxeDG3PnXQMh/1U4zZBcWMktANSsBMcbXlrwq4J5r8v
yzdfMMme/KTHN85bKlV4KB2fqV739vfGK1CuGOqPTN08CJH9HnWlpJutmMCtWzYd
5VFq+X6uMwRwaE38hLGCJcpSX0QSK74obO926SrEDB5+gcd4eShFXsfoZFdgMtXv
1Rqf0G+fOcvPK+V0c679FFQIbN9HelaLwaUhMjBU8geGTQFrCMNn6UYvTl5Z+bPN
vQw9Rfs5YwZ+2PCSGyLKnIIVjt95xT3iMHuaCIG22v8DD2w8L/Srv5oQLj73GvvP
Bq277bP6B1ldccksYXclatQ+TYWtpgZfusd0natzh4HPA0gUqx0EJ5NFe/ODXUHb
p2OEU2/Wte8t059+d+C962s2y1/E8UonwEWx2uQbDzDpPVE7eDiSsX8EvFLxKScV
nvoNZBsoUCw+qUvv9/Tn2M9EliDaEi0ViAFcJpKuOZcGrE9VRyDDFpSbBXMiQzUZ
zFyjFApH/j2+/fJB0znHMg==
`protect END_PROTECTED
