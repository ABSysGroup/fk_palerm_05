`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MxlUUGD5EI7vvD66toR5xSoP75S6CLhhs/W/8dNWGeJjlrk2TYgI8ApZa2j6kqyr
VCOIO5Y4O5G6H8cX55SLbaM5bxRNmzS/a/gyGJmplk6nALybHL0CdWnaTftFt/QB
9r7tzOEouFF595NZRmFAOxn3eEj99sreJRy2Ktb4RlmKizy+8wvSUwMY6I8qOcMC
zS1Yulzqt0a0buKwyUy5jHBnowe16ipk1tiXUP9+wtBpVp/yKuzmbCNEmsj3wxtx
2PQpL47wwTPpHPKg/MAEbC29J/uWerD0AZ633VE2vEzKFelGfTKcJeaGEMvwjmrp
LjFRs6F/Y0C7EqXOCNGVXWXDeA2iYxzAOnkn8zOmahXHqu9nRkHx0VXo/h5hM6AT
DaRsZvNfVRjgOFtTpSPJ5SNsfg8IyPF8rSPZioDfkuJ4mHL7Smd1KsttsN5wa/eh
CJ5dJ2KmX8l6onOXI6by5LyIraamdpVNEBlVr3uCmpd+0hNF2/YvuaCx6H6KRLjm
qr9Hbr7vHBDyLam5p6e7Lv0Pc5xf8YO1RdHY3Wsz7qaI292wXSknNG6YMW0K5ZSR
x1UCXKXK3aulvw7iN8rPwzJZBC5NL8j6CVZC8lpHz4x9heQ97TP3zEHELyacTU1x
1PscrmTZDqNuPUgQzxbfI8VVRs0zQqIOoVe6BokeGpo2CZdzmnB1ZFT4tsb8Zrkw
nmWYFe9SQ8A4e3vTrmnNXJTXcPi6anFVjPTYtmVRJvprc0j7bS0R43yxD7RKrA4a
t4q02Mtxy8+IkPyiOrfvZ5Hh+LznQpufdT5rIWMskJUOLK3f6oFH/8fTcYv6S9Hp
WDsti3g/R78Y27xevpwpWsQRabikw8dA82rlbo1yJinxxHf4sbbFAmCwfBs52xqS
uZEXzuL5K5k06VaAWdVxjWyhFQfJr8Wbb4YkQxcrglY7gvcpoMGUYKJPsUKz6zdd
HR7OYNSb0hUotlTX6BljKfRShRuKxRRqJgvXtHn5IiA/uIKQ1cIK+a7uY1S+ZYfJ
bfsX83MNKPnoS9Og/7XRQKDJrt51VY46YGOGJ2zibsFjING13xeNMNu+d5Zq+rHK
2SgUsnoqit6t39UIgmS4eN+hjbQ65DLs3ol1FuQzaUjLgNhkBQtBn39+BF/3UjQW
hz2yvqSZgX7UeM2MZlVdg55pK7ueH4Bzxt5GBbwx99NyzZ4pA9ktxh44669FKlOV
WaeCv1vAmYHaSy0nTjs4abA1CPrXTAuIJaLE81/ECERUtZkAJKoXlzRSykbnWj0z
QSG4MB/6q7Gs8+N8mybHdfXX38KMHOgMV0WPDfYPxbJ7xfUVsUznjZ3sm7nWxMxn
k5eCa5rphToK1pGIBHc+X9UsDRZLkoWe5BXYxigGBYuJjyvZG7wpC5l7FUDoEcnm
vhiRTcSykqekTdaLaqg5sU4lEPc6sFAKvhB0R3vCWGFPAAJMPUwFql+tP8RkVhw2
oA9t4IYU0DdNVzmsf8lax0NAVqOFyBQQzOhQeWTFa8UfRm+ULPCsBVF3gh4O8DpI
iayoDSXJq+mbEuRHjOGSwyDh8gNc6o6PxlGebdCz3/HFaH1+DPY1nRohfKBgbsmW
1/2VmMBd9KWZwHeUVJaiiQ4ZQgyU6B+zH1/1a08nNTtKqhrtu/J0qwyNK4Xo0JHg
aoip9A3/xItbj3Gv6laFC7hMW6AAAjhae+GfYnnhABV39yltU3ep+nv6QLLuNvRd
hvUV7VxcoMqfw8+gCSCV72rSLKwFeKH3+3/tV2YFyXVktIg93s5JC1pdrw+UZoYn
M8vSOxULKiSry2WBk6uUv2PTB6KmpB0VkjbfRGM6FpolmhXVCdH9XAIi1Pwnaz0s
mStdvb+PtOZn6jydYHfU0DhCATY9i3AsqNGeyBIngnsSl6IaFWOVmjkdaMBUTSoI
xEizGKOYumTO8kiR+hwXJ91KSlyyY8b1wta7NiPhTuRuuPM4dz6ITP/JR0iuz3Wp
RCK6Pi739V78CN6xjKO85M9zno8W6Z0UT9A22o2nXd1+oLikNSKyuYjJRCy1Ws00
OLqSAcrhZLtOuW6Qt79clwbcqv+DGvUmZsAyz8pSggVoxfJohrn4azIcd9zS2ogq
pCKy3lC9Jp6uatv4AAPDOkUhsonyL27r6Ucju33ARzGkh87lwxc+nbgt95yNCtYp
AHGrtidiUJhEYHHsTTfR2yl9dlnU9k+fUdCLFdq/lgPsk2XiBWr4gAsGYTCsnbkT
M+1LyZN3ZVbPHQVTKMTK8g==
`protect END_PROTECTED
