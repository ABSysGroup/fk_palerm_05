`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Z4vrTdZbKMu/MVeTzYjA6WRwY/b2nZBiIrYq9Ev5sV9DcurM13HXBvPR4uS6vvz
KcWkyE64uk5mAiCHOZxpRKktvu/3+ra++GFn+qG+giuPcXm5kC6lTCTzz1XYuotV
X/AjnWN3ojc2zIOVHFoHi92fTShuShe5ZqUM62S8DhNrGqp/UY+KFragzcw2Bzi4
4LKWsBlYKtXBskIiD60Zr1JUiODvPql+uC4PlldIMMjehrU8nWeqaSYj54ha6D/I
VAP87L/lvk5jsJada7VcmUY7MZAPeiundyTYCG9ihXvcOt6HMQXGZmR3opKbLrni
BfnXl4+K9xGtXwWw8HtHRRHKKuT/+yUakmw9fAhoAFJjBKSrxRdkEbEgkzejI6pD
Kpyg+gI6Dh/cYP9GISxwA7Q2PQB1rESlyn9nTzA6IGA5Any+Ka+DfmWdzXaykEIR
vIfiGAKq8dUdl7zPIAgCXaVMkMhF1aoqtKhU9bJc/xYoK0zoIIGrRu+PWHGEpeJy
oFdPTjJAM0/lbZDUrdFgUDnxowBZl+JgeBDhVHGdP8zO2dvHIEhtivkhUgbGd0iT
T1Lqw4mFT3kK69emg4uPR+LOXs9jwc64XpuL9E5CcjqWBgccIzVNh75XScDinxRU
1eUdNrQHjkYbg1cI8es2v4GV4c9VlOHPe0CbOM8YaiTqc5wizV9o7I96gF25dp9q
hmVLSkulPt4jL0gRqrQZ7LTQTmt2rQ9e/8i1kmkiZQI=
`protect END_PROTECTED
