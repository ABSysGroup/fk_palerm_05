`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vM0HB9T+rWciJ9Z/u3iwyoRVYrzztPbEaTap4FHopRrJE1idyhEQvaGOEjDs6Lhe
T0dj6F7+F3W9H6mu6cTdz5oyfNbZ7RtqOcG0c1mkCWaPyubkNvxSp0qhhX8BnrFl
iElI6VrsUczBsruJrMMw/SQIeZYqHFAZ+0ZXnCSqmSYrDklFQ32LLKbH3HNrZmFd
pNa5lfdj4+NyZLHQnBy292H52FlzWryH9EK++uiZPsVVOISyqhtmKcjPjvHJpuxB
eGd+vpl0wGXVm5MfHShDSGVgm7RmNWNZ2Sp93BJ6uTw46Ia/iXXPe4Npc0ocDy+W
iakU+EE8xt4ao1D4yr+37Re4J8gzFpBEsiK5fNZ1CZHgl4t6wI1IqkQpfUlqHe9B
/z17iOm64kC6cZjlkF94SpJ8qKLUjUcoG78IlKstUn2BEuvr3nKS61Dz6Ut1fBWe
RECAewdjN02YqWLTwOHcQhUC0pYSHklCOzpYVlM/x9cHtisv7Nwhs2mQ0IDAanpJ
n7ZaEhOeSF4CukIHNh6f2pxW1yE21x/asPsbKbmWzAE8UPQ7Xt6tu2qgXiWki+br
frYMJpraOPMkNNUsvyMGSOMI/qskmm9RAuHaltTNjjf25IqscU9RUoXO70HkmuWn
tsZ+B4AuxxUD8ODvKygOQj2vGihOZNOCc5OZJFl6JbFo1JVWk4fnpJxVeqfPjz7G
Q3+rB0DVATkk8/QR6SLqiaNxp3muyHoPiNolPihFj7+Ipxwz7NFDxJEIbocrBL8Y
i4nml7jAwL1CRMXDb0PSOEYgg4xpewHfjuMq9pjM1EN5Y4QdRfnKFH+4n0cABCip
rhboqBU/4vMSXSGf5pnQf3ZWq4Z6DS9rNvqjVNbJD4glNgQTODziHkWBBcz3jtp0
c0SJi2O0+q19C3YzKqigqU/u73KJsIBnYKen9WoJ4Px7AfJGtIvgVvEwgF0ec9v+
yQToOnIWKqZ1MSRfNU26nQgwK7gWLTjbK3PsnOCj2hTd9sLkfD90wJ+nY7Vx8svt
GelD/RVHzCH6SyEWP4glJWUQuqascmEKwpd/8KMAgvLxtoJ+dUojADJxmleux1Eb
pktRBd7mYK/paACKWX13vAkujgzZ3T4WVrPpcDayx78aRJB24HY23IhrsDJog9nI
gyUhswngFYgDyBx6h4yUBz0leKUwRmjWXJ1pedAO/oGRG5Vo06cWvL/TBqZekcNy
xg/rOQF2Df2lxffIi5GObt0tr+574SJUmOFuAd+ctuNWpzk4ScruaHAorMH9rHjG
wkLxixY05/Lz8iBpEfcs1YUapMDYdO8nY3xh94s7ixgxGXUGlrHnLm8lLxxW1LUd
3HEllNGOFtdgnv3LniId5XcLqt5c3UeXmPw/cVO40T8HLr+CiNGckOqKZ/Xd5Ozc
pu9y46GC1nmIeScYunOz4xXoTTtMNZdJiCSSNArGQTFDWmtpnlplnx+Gn7ARSBu1
CXJ8xl4D9lIrHTk7Zd1ZaaSoGfeD/bH8AMEM1SEwhFRogOawzgrYM4mStE+oB1vR
wZwgGoYkJ5FFPRfxDy/TaZNsmHpXfCs6h07PCfBlxN5w3aVI0lqromPQtf021rbK
Errm3ruZ9aYS7JUPYLK4FChFzpXrQrXzopaHvQHmyQP6XGqv6rTjNOtD/QP0+NDn
veWmrXSHm5F2IBT8ZJVktdd/Kzo/2SLRru1ACSDjRkysoEPvuH2sE1UpGy5Z9uK+
d28CdSzM0HqxaS5CQ9NkETY05csPEwTnWYysolfxyiz65O946RSxHgguqNfew/ct
ZWlzflUefZiUuhcvZz0n3HlDENG99jwD9fwBeaYaaS9+zjwaYM9qci7pdaALrY1t
j87vYMcXp6Go+r9lpXkuVzKnWRnc20X6nBmfMN1TGjDVJnNVUSx2dzCi2Z+Gkj7B
qz4HK6xuQHPteD6XKc/vxIdK+uRf0IFhwS4lUuzWptPo4iW5bU/gUGUBwXH4iMaV
llycQJzWTd3gdM1ifn0JBEWWY3dXmGhyBCFi16em2tvK/mq6GutNGzC6ViyEyaRq
HdafCoxZdwvG3PSgg3gzeBmIx8etIKpTqfbFwfY30sy0ODm/6RPLg/EyOZPCDv8A
RJ/ZJLxEPKGeQ8BjxZaYpNglIMCHjh44EI7bBfNQ61fFkqrPsHIKigZmSw52avzW
3an0ezoLfzpQvJHb9yrKnrdOGZdolRuShHpKPMWn2UKWfcExi5eax0OKpUucvP5Z
mlIXoyBEpt1OR/27z+m7OwChXj+Urf/mp+Ega0F11IAXc+BMNi4Dii+B+bgUT0Pd
pHztEt10oqUxfT4SpFcSVxk6MoJIXulj9n7D+IATwJn/bkYkOx7mbrCCJHuggFJP
WikbpHz7VGjEJk7UUfvi7SRVfYMAL026RUdLvdpA7HDtS8PQJpOY0xFLFrtoOcWH
D3/6MFBcVgR9uj98LPMY+E1SS5Y2y4HGz6TJEdlBmR3OH9jdL0y5tL3fGm9xytBs
HxKktTv7uu4R61bWy/h+QNQ2JKhp6X0Ra0L07SkD3RV9gcTf1y93YZRVZXmWuCCp
+/r7tNG1vGIW4QC0iw9CyarN+DdQb9N7HkSN2mcR5tRAK6a32RVXlVRjmK88zXbc
ab4wpsSXr9JDM5DfjshVzhLwmfAfypvq25m4QWKqgmk=
`protect END_PROTECTED
