`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4mYu2BqOYkcwbeVO29tTV6zAVlxM3yss+Yxf4KRXo7Q+5CEr3ZlL10soPcnUieqt
H2gBAuGho0G0TsjdPqiVfuh8fZSCW+zCbTy1PHcOzKObDp3QX57xi9w/XQ7EDI6j
xzY9BIkc2YdeBW7gydysHNEL3mDfeBYDsATEPuHmaXTz9PoSRl2CYJGdB9u7ilPt
3rgur3XxfIcgJftc5o56qj3Q+Y4YtjGiXbbk8qYp/qWbFu/zadxcGeioNjcqREW+
VkQc8WPVPWd04K2YZUhkNfIqWBWxKLcRnnfYDAYivz6LmieJ+CApxz8DDuVkZnEq
QGgQetWzqCN404uDPibdDnT7lI0hnDyoSj06RBWjhnPWWUnKzvwu08ipq5Ei7qLx
+ghhLUYptmPH2ZmHr+jvrdCuhFnaneaHLWNDwkqH7LdbMZfm+5VNCLSrCJeQEq7s
+x6Njuqd7s4Y4JqUspV9vQ==
`protect END_PROTECTED
