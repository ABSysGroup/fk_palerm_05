`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pCajcgGeH8CH+doKQ9YOTYLfO5jsOZtfcNXkyXrf9D2fdjG1lDnDu29QvEoAejRH
1rFH4mEEXNsLv3rznhGNOjTTTpNqdi1MOczn9wLJgBaAhj+4SwhtBn7NYBALrgMM
10z3OkxrWHWsVmO53qxmQltR6zcUyEC5sjRwcTTU2QPgFDpcUjvQ1empfuqm23lL
i/7fuX6tgpgg6TOFkl5W/8ttAN8s3hqgy4i0tRQm1wnBpLUijBOfno9SZK72ZFpN
EJ1dPzy5VwyZ4ARJdxxSlFNG9ubUP+GRUv/z3w1UqWpPEC23ajPhD7RicJChOuUF
w3aUUOSVDuOELKoyKbak7U0SQIpRHHZEsrjq0zj6Qq7vNbIHlAncEQVAfoIz10kC
5Heq4uvhbd4JQEwtw4qFENOmWp4IgjWX+N+78PhCfa7jYPRDG9OqBarxXOtnlz5n
78G5/vFcr7Zdu9ZXT+ljt3256q+v7P7jyF7tmxOGg+ellkqwxv2rT4CEBscyZdUQ
GnhNNqFnO778jFLqkagF28NvasXe6qG2kZglRCGSVypOXiQpcbNGfPsDMd7kjShP
TKS0OlsTWV6gbtxx7zJzyjmfDZxANixTDSXz7FwI1Sj2A+jyvTyMDaX2eiRDSZL3
IdUhddzO+Y362P23mibDmw==
`protect END_PROTECTED
