`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MFgEGMgX3gtZBRvtayJzv/Ssf6amDUYwuiKMeahBhe9MoR6tGSfugsRnkHtDK0V+
p6kw0nKf1mBxLUrwEYt5YebKDpdboTjS9ge2RzsqUToTR4xVFSQg6L5rVZQeb0MO
JFPMeAdmKUBiFIBRkkcGzPgjOdAPHSrIDURvuY7NjMuO71VbX5pchU3FdPG5dx/k
yxW7mpjnMTqfxjLQqFfVdoOII826ahMykJ2ksc7KicPwyzLyYEoky7t3hhqJyInp
ZI1yflaGCT3mbL+kXbnUfb0ICK+v9Vfrd8FcLLkioIZy6uO5GSvzAO/SlHdDVP3J
hqrAkk7dHund0MtGAwkgJw==
`protect END_PROTECTED
