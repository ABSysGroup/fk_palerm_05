`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i7gYXiCuwT/0VGbwAY7Hh1RrUnLQH8ZeSeBOJBH5y+7aKESRTQCcDCIsxMTpQCrt
UV38/B5Ar1NHgM61mIF0/VpGszy0OHdxvz0nyXNeZAHTXua0N5cdapXKoWVe6Arw
NUnJ0m1cn3+vQSebJ81Z30zoXwmVMzaQsU1tUuLoh5Qf2eo/xvfXlTg3aGx26k9L
b4g/E+wapLMUSiy247LDYHJwJEo5dWA6ng3sIH8XkGHxeMdKDe16eDeUsIb32oSF
doWZbRJRJgs/CbByF4zhGnmTM4ENyR21Hx7Xg1D/4heZqeutzJEMGHwOjWwW7E5f
doemyoPkEQmJTFnq9V5ukw==
`protect END_PROTECTED
