`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GXbIISH4BQgArjnx+tYEyncdhTbf6bXFgKdlFtnKqV3JBjia84KSvwDZ3UBf9ovB
TrDGsXNvt+Nkf5jYnzBES8vzOJh9lP4YDpuhvJwhjOkfejt1x4VQp4WL73ylx8YU
4TJdR0FUvtD2BK3T+Ch/nPl97xty2nqfsbqhyGI6x3W4DXPhJEZ6AZkMQ1r0sGH1
W1YuSDMgmwOcQXZfU1fcnMY0Kh5NUu+bJ9gTzxhxnn42hy/iS8rkvY83Fs8X/TWK
hYmkVvUhKEyQ4kd5rqrL8roo2sh6l5AqqgJkQtVEjrEv4ZMOO/Qknwv/WVICthLt
zWTRhq8XjznVjDDR0J5uDQ==
`protect END_PROTECTED
