`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mnEMKMU0u+a2c2FgQKqHorn4llF9rJIlY2nHkjPbuBkm6kr/AWaEUAuAimoFvFuL
LNa4bmCCDqbCQ3G0Q9Xrk34qSBDPXn0pjiaiIENiIobtJ/XZe4jaGDt/BOaRY25y
GiDQJm6Cen7qFGj2laFiT0iyS4JlOkCY2OCYiEaFu7FaQ5NiP6lsA3LtIxHXgeZg
VhZ/qEq3dc/djGB8/dxpWyusYmS9jQAKcKe93GSJZS9pSjF7pklxFz7ZAdlfjh8M
pReY7nZ4g1bGgXdt2e9T80BkkV0HVLyAE94Ke/tmr8yfv2HxVhcnxEq6HiofWpmV
r0/RYWt5Hz4BjsJ7VQwAswGcCzGVS7VLl6O3Stnb9gHdfI2GBfPumSqz5NHhXV6K
ChNGddh3Cz/8rk5o+ivQBiXJt9A4aDMv1O4pkh1C2UE4qMVDUsCGC9tg4Z8dpaN3
u52qGQTZNCTWrivJAg7PlTrIzZbVmNZy1yEzl9T1ltzwpCAZ5yOk6PbwtAYV3Nn8
sIvthXRAV0Ucckn419lP0Q==
`protect END_PROTECTED
