`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/z6U8GcQyPmsHn9NrGa2VXnveNOMebDllV+lsnBrY1GJ4SmFFkbWPxAwaLlVZXO0
lXK+49AFtXnqteYEYstavGj2SIU92nrZAzy7lib4PmKVd4p58Ya1s74xG8efU39P
uyyfA2CP1V/Vea28uFppww+DHTxeh/GdiB1sK7jT5xZ136YgLDmeIxr8CJB3myOX
AMWTlH1ZvZK++dxZFnmp/ObVVJWjb2AhnRS0UlToC11MknajhXqsDLdT0xOzndhf
AvlHzNwywqveonJVEeD+iBPoxz/0vLZavANMU+j47+gUwXphLRgwJv4Xm/8So+iP
O+hMIfmut/pHTwb//qq89lJE9a7/Yppm9dROiLHMFNiVxD1CU8PZWrJ7L1N0A//V
a42go3HuYd2RJnmL6lIaek2Wo7qfxrcoqnLO3q8DLKkUh6wdmJR868591jTXtR6Z
uBdpjycyVr1i+UXd3l7+rKmiTsClkRQAR5dp/XEdpvbIiXQKoVXhtsUhyi9GSfQW
9UCqNiKsuIH6POhEXijInsoEEMZBNPM2tOnAX9I0PiTPaZCvVgel+xsG4HR4efiY
mXmQmiQFIhO+kw0I8/VwNMorz1DxCn6lM3ywU0pfqOVXR1TSdaCmtvJ4c2fDiUyr
nsTBHHwm9513eKoFeCefRoUzI6QDtGZhMKsAwrkGhm4=
`protect END_PROTECTED
