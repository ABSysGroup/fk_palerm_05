`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uOQUVtJppsHY2d6w++quDDuDxjnS+wGvA5uDBiUd+x62LPJeTX6T7kYW+kA3D8iJ
EUjq3gw/29Za8L/42Xntk4FbFkxiQ1QEn/6fNoevlnBLH1LIns50IbAlSpjG7iHF
aXQVXpHHCSudx7tLAiHMcKLbDTl3yucr1sNaXVol0BxaixJfginuPXw7TRcx2W60
VLYDLIl/5j6/iMGJbsgsCGhGXSIpl57ibW08/Ma4LVDE0Wvx5CiXiZQdbPzXf0AE
c4NCMfZQ37Xjwker9KEFpsMJF2Jwj+ciJbktMqKgxGZBLGudMvFKX6JxdGdd0FdF
P5HYbiN27ICgtRgNJ7bI8qNRrRFlisA2vHMQbAB2iVXt77HKT324TP/KXI3JXR8m
Lh4nLwQi5CUd9sun8MryK/1dd2sxZnEDHZqed3yPTwK5BByJwSFOUspkS7La/cUX
JMR4GXUve4AL4Z6ADiK/FmdZn47rQI6FgSiwXqhopZ8lup858dwCq6t++yfCyUlF
+mIQeG1O0YTn6sahpHoaqwuFszULQm3CBHJPfXwvpV8qmCwb25t07qM1SYGDpbfi
LAVBvhRJ2LafN0gN+6Ht4dDusFuB9EC5jPl10r0AFLovePw968T5bVfFVf94jnUX
HPvDsS3042tDNgoukMiZ31k8xgHrL8RrXKcL9S67PqbSjeD/5Ira5q1fHd9OpWhR
fTBM6qKo7XJ5qLKxM2ahPJqPsQrWZ2TH2PH55q/l1fA5YfjqcDo46Tt7MncAOjUr
TIYIexYDIXXF9xJq19Z1vnSxeO8t2am/gspJQ5jgy3OibqP1M0stRqt6zDPEF9UP
x1UIV6eXaPq1fKn2rOMKMTkerPxtIRDKYxt+EZo4O6ZlwWdUEXQj3GY9qbwI7imD
n6ysIevTP6rlnCyYSFK3HAdppig3AzNYQ/UU16vi2fC3qwjkeJdYiip076dhJM6Q
JrpL+ev41Ke59xLTaI2KOQlLs6y+NZkZfdQF8K/CsX/9wqMG676dj3uD95Z7AvH/
z8GRf6wBfrNhNxRH0NEaf7pudDbr0IsjC+Mlh/mXIROzIfvRauky78W6cRXh1aDm
n+GYuVWv+VOwWeeA9lBpUBg1j8+WNK2clVXx4B24hucyJ61YsqAzcpLyGxNWB+iZ
b3W8wx+ZjxU24ECoYL08X0ja6VcPacFXuJep9pNdAOJcGUjjAZcxuo0KLIGtQi5j
vVMPUT27i7ETVbSeK+nqo4gDM/PdEou/gMjeULgQu1FChY/X1pMbECH240+dRQIN
m9QKKi9VtZvhL+/+ulI5IR5/NsuyQNiWgoLZC/qtawjEX12Oco6LU/eVl/XQZtcW
11q6AjxNOCYcXShLQQCI3kj2/SOD7a36u2tXM5xbXy/0l4gXciA5RNDUSKbihqXo
5m0iNzIrMj3bo1Znd9HmpwlUNZUgMG2WMT+EJT8KrKpdtdwB721oKP8y+NLEsrSG
HzCe3zTnYY7OYF+TZwCPHvHtXbCEKALCYdPXDeygLAdFUhabOwcx2HOiHSB++DTq
pQpG8PueVwkh5d9L3ngSh/+29eC71mzN6sTacaCpcgIe8BhS/uBe3hA15V2Ja9TE
CTsNwUlCaLDsjb36zfoTTixGCjYGSDAaFkERDvgjC+cKGTvrl6QipAXYa80X0ria
TzePSX0/wc+9GhaeOrTsLRzyH+sQApJHFlD2IbVWY7c+OIxplF4phhZR4PA1exKj
QzFgPzwg6yeTLDtZiqQmmUjPvZ8cCqm1EoodoCP48Hg6LYUEY7yhaoUQHByYC513
2g7xz2MYnFaV1/e8LVFiu1OKkZadaGr8THleeLbsqqJVIP/kvtzqtPOj3RgRLfSv
iwR2pbLF0dsW8TpW0+xlu8yVwWj9yWHdikSbOp8uD+tgHiqVnmLMLtHqGX6Vhdfh
dFuzsv3US8qCnSU5hhkYaSUijiUGA0OwBOfKcQVKdAElt5AkWB+s99RRQRhnvjzf
Pq2zgkVnfK1GDUpVUYcYzRxiIME1O/fwD4fbZcG3c/weOQVQ8hjynPSLuwSj5rEz
IkEa9ET0VUqKUR+7jLuKq8Hd3D1Tc3nFzUWDRQfk0eKrW9q760Rvk+sQmPLwhXA8
TtObnPgPMXjAtuMgozIToD+L6ft6+zTO7lXCvFYkLxDPS1ZICH8+xPoPT/Ya3Kl6
ZkUrQPTH86u9Rl49ci8UPor/rq2bj+Eby8egCKTqceGqHNz+dW3gq2kX+v+wHq56
xXTdgWH3sFJhPtkjUsW4bGT6gMTK/PjGw+N2Cl036nhkxLrpseyk5YPpiZwDq9ha
cfUbOJPt+9iRvQfxsNCuEWfgj3qsdf9xFqt7k7yLFj+TOG34SiLlkWoMRWtwBUuT
MA5/gpc8hciP2fOI+wQx+qgIFZsklI+NrGjcoH6ncdo/kiEtYkErsLoZUvUR4cBk
e52OVCaVy3sNkwtErsXCGfv0MMyb8Qe05I+0b3Kly6pWyYxEU0ovBqvjh6nbNcL7
nqLPYbOlmSck3/GglAoitA==
`protect END_PROTECTED
