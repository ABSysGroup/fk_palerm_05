`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vWJZIx33H2z6pHxHKvhc7NEWyB6EhCNRoqK7sOBB5yU5XnSvGcKickbqb9mrAFCr
lU4/fT6JAigkaRF54GflgM6RACXVkwNqEJbzSXKXGcF3T+AMehGdz25XbWssJjJL
1tmtpGVcvkOJoeWs4nmNVSMfda1h/Ov+UGHwQziy2zIK1CEZRkIrGwzlsUTGWRNu
uETVQ+97PblbhjkYSGdvw/9F82oYsLEiGNI9HQbhpoer104rNUTDpVakrZvSiyI3
PYc+Ngiw3T5U65mCVfs2YkQXRbGy31IZT6IQpS9z0BfLPP86RIrXEpKNwrXAodiG
1irGD3bXicu0yM3Fu5/WxqMC5nCmrTtkXLb1dM6xOleW9z6+JSJBNjv5d1QNUHdw
Uti96udUFRI16my2PxQdXTq18bFIjOhTMH4li9xsAttVSNdLmAx+Cwqah5oOqoQH
QPvFgouwTSXZkVwY4ZhJ+8LhJDvXN5WsxR70s8JvOV1+QAu4nmdmNl4WJV0EBVNN
fq6lQLg99RkaZBb6l6js/nOBzudbiI3Rdy0VZ5eluj5KoX9hOi9+2iKrwUdzw4dw
qh+2E9haVKF+Mxt7iQfWLcnHjScEFzy0JTV6Y8O9PNmB8BxZLjyADQwT4NBZnqI7
Ed7FSUp8ThM3mT6LA/ME27SaS9R6cMjhMvRimd0vYwfKohgV83HMCCh6umZEWK0U
`protect END_PROTECTED
