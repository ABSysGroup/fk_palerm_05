`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qNLRNE+KWzEAduMnOIAHVrppfKt59cOgCl5kSPN9xA9Dj/bWGntbow40UJc4ylqu
t/d8ucnmH98HMUGoXcCTfaMd51QjSs/GclDms7/oz9Q9UWY+eNoeFDQBV8+kcaIy
Ksimf9t/v+a6etasUdw6pYySyNNndxnKcqPSTBeuLpE/YyDUxFYQguVbdXMEUNWn
iK9nNqTvsnwAVLDmnHnciheM5iIHWn5Y0T+OvCIaFD2ROG/hav6w4fUz9h6b3VxR
L9Fi+JKZIFFKPfZOTCwWtMJOtX6aL8MNG0NRA5bqJiSVawYlhj4Lk7uRfiFE2oMf
HTOOBfEiQgqinfR5HvKzFT1jX2RtGDAtk60opwWOeaJau9+JXEykd+0V8WTm7GO7
+Yj8/ktp+Tyq8KaAe0KeX5sDAzpxGTTdTPF8Z5mNKtqbzI02cw0MtZ0VENVmxgSs
K0GSNfHyEGNqTQm29DDmQHFfocosqx5DbtYzHRicht3Z0xaOAS0kl2gBMpffqUvw
iPUZniUCxVyv92EhT9VcVCY3LXlzAS8uUITZNbhaVW0c4eAb/tcZ7Jznam+6Wgqp
AUhyygqgn14g0+AF+eQfZMZbNVe9U6LSPrKgZ3ftR1i8Z2xN/58MVYmhwhawWfjr
rdS+pe4AmzVuEY1upBziVg68BZgX6/cFs6uvNmCaGXlyujz+JJfNxXtrzKSO5NWS
IjxsiXjBA3BqABjh132HfCgBLEK9m/IIOI361zzB8J9eGGhWnQn2qdd0xT7dGftP
ZOLhcmlLZQ0/6krEA1NVDCEfufSjj1MioE/QSm8VwefNzkevzcAPU3oywK57XG+6
qFBYzrMLPAb1qbdD1cavJlvHgd+XSYYT6ICvEHRt3w+ZsKIXtLoVvNTPdrH1jevG
vG9qFSwPCp8EXDdGbvs5LV3Llc9hBuZqVPozqafNTmxyGXmBEMH5yTrU097N9JS1
`protect END_PROTECTED
