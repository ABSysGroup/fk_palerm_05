`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1RYD4IApEOK82BNNvAMsh0FatvEIc4mBOm6PjlHTmXJSirDlmfzTHVnCRMD5bz5f
tq1vRrx/jGQl9zOVicTaSW35UUlFNLlvGOGvHkhDZw5P4aMevogzJ+H9y7c33X1e
Zwt9tv7YKQuWeBoUFyajM9outtd2cBvHiiVeyiA1VPdvIdAiggXax+70khZxxJoJ
+6zs+ZTiBtWzvjcBA/Xzsz2ABknqWOKPIXftH5VsdlSF70vmwyQpfgkQmIwLMi95
tfWhgNcK8nrgBCgrZiOzj/qL/25VCVlZjcN/P9IQc5foLHOMvR2vYPcXRHcz/u7S
IqY2iyQpFfxjr72syN1SUnLdB2Z/XTz6ryF6E55l2yA=
`protect END_PROTECTED
