`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yfys/BPn3LfoWkTzmw2IPj7l00UrVxpMmtitROI7Rxst3WqElLuW+1qg1rfnPIk4
Ia0gvpm3Zo41hpBmGRZ06MWUKoucLy6bEAOYUGuofZ/3tGMSGXd3Gv6yZ9iUJeCN
Ei5dOh3Uhunm+KgoURksvXsgDvOc7Q++DWBMGR3SQPy1NYB5A3dEknTkjw3Xns0I
GCC1KOFTQMLqBIdMKcw7IohBO/w9Wwofav84BnACpq89UlWkfdMSL/s10xpWI9XO
L93KLGgbBB/7Bu1Jv1VuAwL0SEZRL23zXlKoefewJoqyZ366IV/wZaLkC+0pWFoN
M7LFngihS9lduFahY077RA==
`protect END_PROTECTED
