`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n+EyXJs/JiW35U7HajafXs6QY3B9ajOA1tgbkQ5Yn+fnHVMvdipW7VoKzofNcmKd
aPDP2pvmNv9UV3YPsp4Hv6DFLxNRjqC0QEtN7pNT1FYdbCeyvA3hk2yOabxnGydk
VWo3DE0HRdDgcqX3UlTB6NJjhG1iRgHTjwd3Y4ttE8C0eIDu/+WhR/nqZnYi9Rie
QfBgw7YoIz3ShPQnLxRpIfCsC6ocTSnC78CEtMhPXQVhkjFYYcHXQ96ZWWqrMkfl
gtCvYoCMigIx4HcVceEUVyWzg4Okif4wKGylkziH23zt6A7v+3kFA4ay7/8hTZGS
ypgtPt5PYulH5mdwgg5nMw==
`protect END_PROTECTED
