`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8i39xZrwWuhWbwGZ0Z2bydtLQX+vXP7/y6em6YKyX7Kqd3sUOP27wADHj9ovoORC
WhiaWWjXk5iDcP4YoSg2OJoq3YWul798DEBtU5LnWLjdJj6Na3IE8WAKagCD619r
VRfN1C9OtuWzxSTmOx9Tf3NkvQLDbU8Rp9ZsHbURr+4BMt+H7TxmZNzFN7TA8sju
09KLHMwoz2fzzn3gfPuE6jRo/iN2j/yNJIHZ/b/vwydwmSQSt3VRmhq9LM5Dg7gV
eQ330O/z75jh2TROH+++d0ZfRwp0YEmeINSx3SbVIiot2oFj7hKk1GvNXCtLGPyI
/bPims4xL6czz1VdIESEB9R5pyVAN5qiGCXPNEGQuTC5TGZ63KeBKx6kbb+bCzCe
7MtUMwn1jIR8ZCWbFHkHVA==
`protect END_PROTECTED
