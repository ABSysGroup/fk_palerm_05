`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dl13RyoBd1vjl0mbWoWCRivKwib63jmNPISH5DQbVMh3jMN8dZQZ1HiQUDN9tYRZ
owunxCEWawJDQBTIE/VBhoLDLM1nRG0Xzxd7DCnJ1qhwITTCu4NDsANvnKsvivwh
xT/2zY6Zo6hdiwAt7Y0LxE6aFn6qhWNJ5G9jF2w6oLde08zGUswu4JMjyOvorK5/
+xpmmBs2AwCEmQ5W7zoz7dzaYHI5mHsBgx2YKv9bPkoFmUobMuFel/qwUJ3aiX+B
C31uECuUCXT9OtHGHTpHuS7vW++XM9VOw1VwkzT79kSYrgFUUnZIiawgQRjSBfO0
3vG3RsfFVWClc45HFNi5auvVdpzYs2dvaMeZkLki/oIwwOG1vavBpfDmb4BMq2gq
QnQBIjFaVgIlhJxNe1U84A==
`protect END_PROTECTED
