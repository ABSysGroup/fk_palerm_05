`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dnHmXLU9peRVOtIfopTziybjJLtjdBVfm/BsnKMfxD7oLyHYJQd/ORq7OJWwXZ26
V7z4/DDE3E2sbEE3Ex860cuyuXh+PtHZ4ZEocAKOWb/bZAvchK7cBjZDYLPQGMJ9
yTRheih7XPOLL+4JJ2oR3ZP3+ulGrTw94WhK4yELD2g6dDx3IGpqo6ZpnVYJeXfj
zr3tNQ8RyqTe7aPLxdZVOXFcgS0mnWI7pP6/LMIHo2UUBB5liZh0fHV4nravsFp/
bUHg/VLsIjA3s31D3v4HkU6kUSkNyGlRt8phaGVtEEgxWuApkRt7SjXOfG8IaN/T
+rVXHOlzGVJSRUiqH6gCedBvRElk0b4tumeD7tDuCPu9gSax3eYfwYnkyB0+GOs/
umOq15aDVDK7QEdcUqqGtI+FcwYfL1eHeftrtVsVEDEviy4NGuWPBYeBhuA2Qymn
Gd7BMdhLrqwcPkSOEXd8Vr7evkKv2ZfBgXX2ACRHOR7tYWhv9UeGsEwoDksJ2bN/
s5OKgAGOGIP89ZhEfGsfZWc1VyUrgidu+zD9orIEYtGsGIZGvvNMNUjN+fJ/dUBa
Fve8Ls11adWNZnvxeDEiCMQKsCjSBL9hscObUB+20VveiE7bdrDiZTQeWE8FMSmW
sIQCh1c45vOibpGLzEp+p4KecQC1G7pJ9hvV1KEcDD0=
`protect END_PROTECTED
