`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TVx8+MTh0uFlVumvkdvRReF4gwQm9GvlYENjrcL2RmIJGMTWXlTcaa5CDZAmMyVX
DZuI37hpISTEFTNvoRg5jC0bDVTjlgQoxiIiQMStG+eefLdmRfcjZGc09AtjE/20
+gzJgVhnOpybNDYrsH5x4EFqAFRuUSIswSXvps+SFJErNcxBRow7mNHrfoSZth+1
gSKRSUVOq8oJhMDC4NJ5nNACCO6OQHuByEN0/ZfpvPUI1zXdropxFFVbkaR5M6YU
GsV0OTTXzPFPETmlF7iYuQziCGZ851qs55WJNMCENv7vdqKsc68KFEXrtzBOkxeN
QN5MUsKheWHfywoCyHi0tMJ0IqaJgyUAO+NQd8ugEZINtvDWFoGoS5eMs8aKiU1A
/y19tMVHtTDKkHoJ7pR27kSTY92I3PZ6g2EFZt/Zm4gvNw7MummV92mWQxIsrsYe
Z12x3wuLLWnHvVQd9CjQ8tlKLcT1Ppb42kgfm2N2t2xH/RlHPYQU44iMenZl2Dpn
xCdeIQcIn3bXYgTuJquSN+dxbaztwyeBI3OGZ8dJTw1imN/Fg8cTKpf70RpcZmc1
N4Ff2HAaevdIjcB9uylS3nu4T7YIiofdoc98ga6abv6N7lXTe2tB5nmCkrSsORJh
i+yVRNcwq+4IH+d90zMrw0htBuczbHi7OxcBJteoiQ+TpfWKoHMJ7AKQhVw66NRh
P+LKD6ivsmTHdWHuUAbLJzw5QMW17KeOEideN87L/Zin3iarY4QUzsOe7D48qrSD
upHQ4NXPW9rpZyE9PX2ukLYcR+CgTIg6aPqWDFVrUpH1ba77Q2yaExM/SPDYO3Bm
1241ySzhXw+DlDtkpPXTMqOpwTXLAH9Ccmw7PSJCQK+htEVeP5ETp+NqWaQra+jj
VBpWiPexwy8hVBAWa4z9hmuRXTGQwJNdq3qXr+acN6yH1ReiK8yeM033d1kDFu0M
bOiaoJV72jYsTandtHoUSMG4/imvMOujXG3y0GGRYyEUvMQ/2MZ6wFNnicYCm3ma
`protect END_PROTECTED
