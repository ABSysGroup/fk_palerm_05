`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oMwZfzt3QPHrv6lmh5UjSgygAqqLK9HEqKNVZZhMAAaDmMh2tMtT192YjmPR+c8Y
fl9WOO6LzELLhsKNaxFS+lfItS8mjZ+asuFaVeZCFbHNulWAUZt7EMjeKlvsCpM/
vYtvvBePo0DQ9XKdD/px3gaU5xSwULEeCzm+rfL2f05yt5lHaJ/EhJtQl0c9Wdzx
w7zvsD0dJekmxnAc749EQyg+fTeCif8hoRpou1LRWEYb/xPUps2gtc0CO1o2b9J+
qnV1REGU+d7u2+i9TX/4iJjdFHg9EVaikt2p7hXScfOScxPChSMa18ur6dX5Dxoh
ZbdtODVrT1WWrAVtZgclM9+eG6G5xE7lNnxS5x3jAHzTo1KItCNZILjRD5DIOuBb
rU6TZrSP+cvTMvF0PqJMp2Iv6lH5KoWkRfOPT4IjhLAZrswo0LPYlD7A7vwM2DOa
Pj+lWiDDQHf+7jyrqj6Y5b0bjBirzol9YOzxg7+rgSkg5eBuXMhO+FyUfiibTCkO
tMioS6uyBe7D9S0NqiCsdFW5M2oL3cKH/H9feqlGecKTHwBpNS/1sj12EwWFp5D6
zsUT0ZHPHYlgZoOfdyVsXET/+16SwGQF0FofAq/HKOuw5ei6CIY0U4MTjeX3NzPD
wh8T7kpo7CiYhXw2WEigFw==
`protect END_PROTECTED
