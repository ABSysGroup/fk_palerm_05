`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bGAkRcgkK5e1qO3QrisFZ+JcfQu8IEEY1HQ2S9XyKRG/jzjQDPANq0cU7cRcZRCo
Hs2xpUBvg0AGY4rJEnzeGv5f/39o+k43jAXkHsuhPE2XCp98g2dme/RcMRgvXGF/
c2AHjDiKK6aiUfZVuQTGqGqPev5nuRWTFqeeabgneNcq01dYlvsBUfo9MbS9ECPK
ys1rEHNdeQ73fLAOfggIVnP9CIESxX8dR1SA8NFu8NewQKcNcIoFCNQQWqrsjvgL
/A2UyyT68HMgSY7Uw3j2v5vMK6Lu/j18Jodhgpb69NdtwoSnm4UjYXiUVZcKCqHS
MHO8ty0IpUqDfhZ6Qb7Xu90USZqA79e/1cESecYRcevehjv2l6uKFgBfHM0MAqaw
EgGLh6CjRsEwoq91s8jzKOV4sGT60q5LzKLcJYl3J5o5lyLyPPSVO6cuPkjpST4E
7ohBL/NU9Pt7do2Rsr6G008KKL09s0doNBH4F6fipCiwQWTjjQ93CM3I2stToXKv
`protect END_PROTECTED
