`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vrze36bkhFffNhqNf4HA54ahkIrcV9mT12TNAmbrR6UkZAzZap3XRWf307CvOWA1
tLt+sW/HA46pcxywB6VMm1ZmQXqY8k1ZmzMO3mAAzTt4fko4Um/AQG1tPzJTzGrs
JoOH+/B1wZt+pf+DtQZmVs/EHop33TMbDiqthHAxfs5VU/H9qZw+ROcWQ3b0L8et
rPd0PiHX9TQmqTzMeebPfUkavcHay3xsYV8ZIAJemTA1OqnY9DIhBYiqoRvkUA9g
/AylxZTbYMrF0JnmfctCpm0FjpYBElJueZ1rbBHGJykYXVHeUmM9nHn++oo+xL5D
r4VrUBX/u3sdbNAy5Y13BvbW/soh65WfPuQj4EU9g2yploK44VLsBqoqf3Fr2lES
NOwellzG4akjv7tdBEjUbc9NVy6BK/oaPuvfJf68k+7Z0ZKYzrEDPj8f2LN0iE+4
hAulSwPHPkKDgmOdwYVxKIhyFvxzXhTen7o4WgoAnV+GH/l46GD6uoJkVtXqMJO8
HOhrZpK2bC7KL0FYZ8jy9DgbWXsuc7Zmjb/Sv58eXKmLUNLqc0E1anNMQcQ5Hwkl
yfXrMpop5UBRb2deeXE4hj38/blngl6IAktrvFQ6UjYr9CJr+cgzVFqaGo8MacYk
V8pxquZLXj03PwmSzcK1ew2TluY7PY9IGIC8A3LUcxi977lgmr766n4lKvswTYJm
pvg7dQxwhNDC1JbSIyw2gGYk8/qcNwU45MnpJ/WYdIVx5ufgeUBHqXMcCqVzHZC/
XVljuvfZ4Hu9oesqr35xJw==
`protect END_PROTECTED
