`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DxpJxM5t3dB1f8Qrc2heft0iL8g6S8S2IfUffdHaQ4GFEm82NbMFpaE+zeulL0AR
oRPIgUg0py4IWhE0K3DQbzj+rknTM34xkPexw2Un1jn3o6afoh0hF0qF+DKpNL61
9INKbrIuEcWog5W6QNnUNSKmA12nqJaY/tyDV3HtsPiIA2MMpTTtu++N5wQu5wxN
a/dhlg6uNDRnk4ZpXkA7ZU5i9dUUz9pkBVst4/jXP1c5LpMST10COHnY3jy5Pdo3
A6L86/E8iaxLQ6jPTv4VaBU7Oy079X/eVpAW9BcMe7vsE98Wd6EzClRfL8ijQ3xv
/z1aHzYnaLNhEMwfiiP+TWjDeDslSIGErPoo0HczPTA7NxCVicvM1mx9QELyVo7g
4wDkW2kd3hAfeBFlZhBFBb3wZDL3SxFxbT8VbrX7Mjpl1ve/RssGMT0dVQDMSuNX
ckElKrNVx+/Wii1N65TdQ99lcxGh413hNdc1mZnfSCs/opc0Q3SAwbb0Xbts5Eel
tys0A2rbgq9cZ+CZf8KwRVhEsh+G6LptEi20CwD9HLoZE6rYCeFULMyivOkPART2
MSzg7XZPh0AlM9Z81iNnK2uM91KzyYQTsSh0CSSUm03p9MsLQLGUBs1B20xqYsi7
MsgdMmr8xj55lcP//RsZ2qt1xDFuYHRsd7OO2omtU7MKTL5Ss54rRkF8DABAEJTW
E5gyKsaZEpajYxjXokOieQygX++utJkw4n2VhA+V2wZZ5eOyO5CAGNk6c7579UWu
Axn9gYJ7n4RluATlyH5OvtDBRY+PyalNv2JmZhNlxN59rJNvHAcN+xAXvZw7c+rD
Uo5JUOH9Qx9iXeqE6AgBmM5A8aDwsoLTpTLsUmye+ZU=
`protect END_PROTECTED
