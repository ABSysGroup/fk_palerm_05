`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7uSOhBWeFmRXtRKYZh/qpNiIsfWpj2PvDBgooz7rLsUqYdSZs1HWLYtPSD2W+4p5
zMa/gudcHxd28Y1DEHIqek+c/OpkWOnSFfp/7p2V+NwfgORctNYEOqK+q6JoBmGV
O8+6CeLD4qvurctKkVsYDjJTzbm1p8MDzGYw8eDLlE8YTbBlm7o7F42qEsXH6elK
pZFCclhj0egV7gZEAONHD5Hihq7BqJO5UlfJsbtEME4+OtP99VALDr2SDqAC0fNH
C++qJpjFajJBAJajyiNP1KcJSoZDQGKfcIIjjpRj2r0B4xR9cdQFOoZhLdVAbYH4
zjmO0ELLz8NyEhN0X5uiob0AIOsoRij5s5QcHhlOzsrMJdvtS7VUUEY4jVWyiurO
Iew2dHNqjWrLOI2UkM3HGsnLbFTurPKIxJee8fRB/CzxC5qWS0EbTqlOOUnSQUDw
9+cd0LFeL2aLE01xuvIEW29Nj459pc+/36vf0RmIH+z9cDrxpV/ZNTWGiHyy/cEg
bZBVTrWiLNe0URSFt3+VOPBYS2HfNASYwdU2YV4icNiOPpp2d2bcCa1vyZI/PYYX
3kQzXLBqKHgbdzkqKktcVQbTp5Vp/Scpu913BR2RWxVlEAOP0Pq93yI0bGSae9We
HXZ3+uIR1B5S9UgwIo4DxKYMOnQaWWpzdlsESalJjp1o0hJpWgWimsyJ749ij0xu
92sIhO5f/kvQj69nwOosT/XIimc1FsI51LKyruPxakGV0enIR4F8TYhY9Cfy19A5
pE/OeN/n2PoRnbZ3jntfytX/4v9ULuCfu/e7LyJE+oYH6PG7g4lO+jqc1acYuh5d
Ia4q1i+fbYwNG6cTJqWdBteoZq3YQBp48szMthD+gTJs4T5w483EAOCArNSukfbg
OvU9mSjVD5nhtiOCHKLwzxaoamzMkaR1qrXVwzD0XnwYzsq0+JOmq8gxev91DpUN
`protect END_PROTECTED
