`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xuoNla22TOUYiyXu8hT8DER5t8AvQcc1wn6z+8NWCklkenCaSlnXFEN1hS0Fc8R5
A+YlHQ+ugzkipWayYRooSJDUPMkXQezFuYHu50vbUttdh6h1+nu7PJm4M6TeRM+d
7ZbGFo1jSVNuq4hr/c5dtI16bAPPnyjSIaCEvy9WmM3VPj4tVOknKeDHEnvoiSJC
szbHBuIC2nuTH4tgFQbKeFG8g5aNVkoMtpgKMpPt2COqTAIiHOY37KAIf3mNmC+J
VhsTL2XhLjl+OAVnZiSOGgGuWEZPLNeX4WTOoZguRlot5rbikZa1r33i5NkPf+eF
vX8C452UUMDSI4rkjokxZnpNkGyoKeM3otKJtfWrhwHp/zc5gl2iQtcrca67MoBl
V9bhtCaHndaY+NIDLEGropD7/DL4XhYV3jlYLZom/UWN0TT9yPcuZEPpLZA2D5bZ
UOY1htWvjmBWMdmTDuaVuyHz79KuHQ3UOmy14Ybcq124DI4HUUthOkT6JYR6aNAq
68Mm3QX1rm0dzHy+6A6SWnYy1rywzsLBVsj/1u50grrugo7HiHL46aK2ZQFnOjBn
uSWpUB39t7e+FYheGwquRI062o1tF85OwkG/S4Qge8g7JfwlOLqenlU6soDim4ZM
3BRkuaeln9pphyrYCWW29GfsiFfY+bCHINSzEhTDtOU6bP6USkqYNDAnsX78/p+L
uE2/sKn+hKExEyZmALIS0SPsu8GT6O9URSaRfePIYGkOEbYj8JekKgXlCQ5/TBMN
7yIP4qLTngOp9X25mq6cWs5IDrfWni8NwKbOpEXJLaNELMU8ilOprcegUa27ZDf8
l5RYoMZnRCW0Sz4+k9vLikEpbSgZZFI1xmyQLxUvGLdHlvmXwqn7DCs3mVyDHVM4
gxDxhM4xh6zT5Zyl6q6x3p0I1VgwMGUY8xP+bQaW1sVuet3xBj2CCsrK2KMaOamr
PhIbiovlQ5KqZsLmz23gYSTEPkAtvWwgvp0IVU7n1kZiVwC1bKZ+gTwAQb+R0gos
aV00AqzdiRzVALB7mJIyFqdV0ioAAl6jJL6Kslsq0qP14F/UaPy/flRr5YimJSbE
Q08NBci9Uhb+GI3LgJdqM22lONAE2BbTmf/cbDG3AhuiLlnAKhMO72YRP2R5g5XT
3Pa8FA6knGd7fz2Yfc3il+O18M1TXiFcSU8K3kkBsS9OekYAEvizVqimYCKxmcSl
BAUrfoUKN5YUMgq6JlKMVTAqChC9xmkAqXPSJUtb9HoZoYTCPWYHaBk8YOnCLmI7
go/ah/qG3w1tLXGZh+XCItF9o67xfc86zXxAvTI/Wxx9MKx4aqhH9a2Lkrcd0zeG
TbY7YkzOhmpHaPbXhDWeqA==
`protect END_PROTECTED
