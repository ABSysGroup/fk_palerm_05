`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sqJamq3kAJF8nNFcwuoApHedFS1w2gtYROO86bsGADLLMWb8dRNxYUvITY7v35kU
lF9Dwvbyes6SEjk/X0aaGGmi0eKzIMq/HEWy3gHHBEzKIWiFY1AsIJ+F+C11Wem+
YMtrkor920EOfjZ36iq022v0vJOfrvMYPFZ/dTMPkZWs9TmPStKNRcLPbF6DP6Au
1ZHb2d4Sfyf1rLtMNXCKpx1nHjX+AYKAXzdkaiozm/dv4UmnnrBwRFPLj+C9/sjZ
vEYeYd9BE7tmnktq15M8enL6X9fxEmQSugiyZd2tNSGl2diu80ZQ2SGsGXctUv5D
ZyV8t16hhPx7+aMHayUuNjdznXBxkCc4tWt+E88C0cV0gqH3v1evABMe36aQOfD3
UwooH/z4L2QVtmw12B/6Tjl4EgmiiV3DeefWHza/RMXZH0RP38clzMFY4FNHXgIZ
H6j1feef7ZRoOxoPocGBuQ==
`protect END_PROTECTED
