`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FOfuZ2O/ywNc9yyA61y/O61IfW5yxl4bTNk6LVF+n93HMSZHbVcEJ7KdAwuF0nvg
QuBU3zqzRrb7z2XQVowkz3DRqWtZmCdwARXl5iVculHFrz9w27tTBvgbM/AnNez5
bxhUP5ZSsODdeiQWu5dw+pj9cajsgYsF2RK0DAz5XvETrqKCOXBA5fpB+0lz3sN5
5F9HvIacay0xv6kIzyIPo0GlFhv7Np0N2UTzL5TB/RAP5JHUd/jSR2YMcPhhambt
SNRVeqaJmaeKUvAOC/Mu6xZd/fJFznFEtTZ47/v+EcP5jVjDtEoF0Pn7TU4bDswi
B9lzT1Z2menbj4iQiWPFox4RF1ReZFn82bOQaZRJjd/Rg224ZXD87s2lKknMGGtH
rb5NGGbPNt4V4qxJDHvKi1i50AfJDpo4IvatdZkacmZoWF9oR7zA9Dng9eu/gZSc
98d3FWdOBYeXPinlOPljAiMfbpU/L4yELnoWSqi58PfjzVz9OvB6cSAE3Gj/djzd
9mk8HNdBaRSgjJFJsYC0/P8RdEEzpH6DubQ3UzWQ/di6OEuauF6W+snTmZzboDrN
VtyglIG1qk8bp7N30igW2DBJmD3ZV3ZA/BI1OXcf7To0AYOd8Jh6Hg/XwT1QzjaO
ocBM9YlTkWoJTiDbWsHNULhACSPcq/RpnTddjgWTMv652VhICZChr+oDUJ/gKj7c
9davA5Z3xqQHHynfarZ1nY6IvaVJ7JSSqgSnUu7POQz3UbazsXOepRWyoLf/wKVD
MbE2JetiekpW4lfNRO/q3aPNHrPdDpKVLRppIvVt46y/Pp/1xG+MVL7gDPBvYgaO
c/AmnZSKasTenOPnfaij5FOb6VH9rouLrIvymNdlQ+82MDMsxHiwwoyQmquyM9pC
GwzU85H4/3T37pW6u8Mer2tlJzGNZOwUnfcO0tDEpDEcEgs6jXE2sdQDJFK0HQdv
t40GjkXifghzWuid+rIppPoTBPWSmKQu7LiDFLFm+HpkZB03qAlgCHwra3b70ayz
a3xF/9hIVt4MCRB4zMQkVIom9/9132VUi92MNNkzAEuXDIKPr4jvIEOi6+IszPu/
`protect END_PROTECTED
