`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
axYZqP/ngPSi7AgDk/Ix8urLxIxJAjK86gVF+fjLkrm2Sf8Ey9HQu7m0BUZlICTH
JqkWQnCctD/1Rl0gKmfY5DkSHbjLfP6PNXeFLUZauqOgpDCBDIzfr2u8IpGAUaTn
jOhXX90KIi//BiMrLnKpg2L6I5OgXMYuLteJHAyFLG1eFwX5gy8zv/Pny9BUcYpx
HaILsuu0R9B8mkWWZ1eAMJHH5ItmEoUmiis0LJWZpoa4TcuC4+RQY9BTAoP8QKQ6
h9oYKXR+KXA0XJRcaUO2//nDdLm539GY/sF/nFwG7SKEW1XzTUcl4cvTL+/eRgRd
pduhl6/EJSBUhj+eLTv+OnyJzEh5I1/6uuFudWZAwY91COR/HHqg/mQVJCl4KVSS
J7VRmVEkVDA49ISl6JaZcENkAOtN32Cs28GtEgzKV9tfskOhyKZgDi5hVdi3oFmf
5ducdUsy2zriXrQB7rG5qoj0p3NwkQsCBNWbFhGnghFGlVZPEfBEhMcQq78cS2Ex
wnXU4n81wFMEEsQPJORe6m27/W5jx3/5IsdNLSEl5dgST+69SA06OjO1a/DOukZe
dbcx/RUtWAHW/wmf2P8ClVlSQNcGAHKpbkBgqykOEXJK4cpsOTBoet6u66FkpBEZ
dU3NXbXncRBWQ6kNnnZwyl9uJLNfolcSG6XjjL9kNaK81C16QwCC3LT209zcdXvZ
yXBFcjErCgKwF33gdfKsMQ+bGVbvq/v4DSsa9M60Qe7+VHxbYvY7mwZsLhfs+Psk
71UU+Ou7lWLGbxl7NsHnxollWQ9Jbg2rEIKoD2OKsEaRk1fmIb23WcfSJyBLT9kY
O47XM8ynelkOUZz/8Z7f1ShnEpIjGBlj7Yc35c14GZ+c/8IyNENK57B3q8e3DKRh
5Oyji5QlC8PqikNJOO7VAVxTrGDyHwfZqW2ajLAdoDZw91JdeBsm0npOI7NRGwxq
OD3Bwrb2acIz8urSAS2vrUlA18JzyL3L9t4XITz0HnJmQxhzYpHQjFtMWqe/k51m
OWAAGcTaNUtt+8/a/4jGy28B/bBA5cT6y69JcFhO+ZxbWDoqJQlCbxIHkN/H/wtu
7EF65yQ1y8BdEwT6PxfPqD1eujMbOid+gh3NTNEeLPjbhR1b46ixWjUp8fPMM9An
q5RiwiQrzuCt27FYrYCCuFkdbUDjdA/VJgTqHDo1n4fsVVFBePSJN70T+YA1lEGZ
2WDX9wS7oIS1WVgmiYH/BHrqTDNa74uHmuJUVCZzFoVxeQkklwE8Fu2an6GXNS/d
wwt77IoR6aFYJWHQvTjUcdX6metstrOgNp50Y33DW9ZWJZKphhZOk7BkvZrBRimw
58VUCc2TfTxQcIcn0JioiQcKI0FvEalt0nW2BocqHoxvxBKaWUZjAWUltH59hU0z
FzRo5+ycTviILzXfnJbm8OegwOKHULybVy0eYBim6PrXe8laiXTttykS6m/wUNTr
bMgm4uVEpJVJGra+rnFQAgaXz69yCiCXFCoDciPgKGRp7VkNnf/4eKmjcJmE2Ktl
IQX3nc2HklZF+7Jo/uS1qO3Gx0O9HViiYZGNTXDTWuZ8otn9CUlKA6OSlCvuPwQ5
9mq9JqyEFCxLojFz6y+kEo4hMe8A50GPa5ISzEnyb9QF+EP0ZFeYhAszA139Nnla
cazW0hNKSM/XORG8etM71bWDa9Pe0hteexFvIevtdOXLVvSN1ag6k7wtidChk/T2
i9gPcnX3ND4eCTezC2RHk8yxGkEaSP74D634IJCxRB+diYanRjA6PGFovBzWs8bx
TMdfYCBB+k736hUF0nMuPqNsqHKnEPq1Bj3m06xo7di9axcK1oVxuOZiy98besoK
REZoraZ2xV1UjUf6/rxXbx+3H6nusOnV9cv8XkRZ4ZT8l3z6hfgaRd+g6zKQ+h4R
tz1r8F1V/UVdyYY8quUMaxcb5y5SGGk1MRmKGMHvP7GZNpKvu4lSKLGKSO+WTOHK
SThPcQVbUjDYYwyhbjUq4cKrJXoHv7RolqAsRMfgAvPP6ABRit5NwG6nwvRJ9kNu
v5wisCidfB+ZPEyzZ3OQWdZa7yJdXrCd+Qrvpc/HJ1QYbeqW/EG1hmIFw/BUsHIS
vJi+y8JI5Uwfy3hHits8kkNS+Nni5+969QwZ2UJKmkQqT/QntB9JfGFRtHjfMY1u
o4mFVnuUVNK1cghV5UAfQorVMxXPATAgXWL3WBIJlhoPLP1VA1cTBLHzBiW/43bp
pr8JE+0jUbWGPiNU0UC+ZUSwSYLQV6NQBhnN3x41N4jR2OwhHdqn1UEa+F8tMnob
45nux3WgSEfikzSkG9KcewnoKHfCIEuvZjv+pWLBuVjU42kbAulmIJf2Fxopl8lO
KtJnK5s05TXiV8pv4Uzn2fxPlLdp+eTDb5qocjgq8QBJndq5wZOl8lTk1sU3a01d
YoHPs70f2bmfBgI8eLw33vQsDIQDqWAiYjUp1xYlTETXB3EN1cFssss3yBVwtqyQ
ohfmDl3D9cGXztzrusqwh7zHZJps5T3w9DXVU4q3fNBLlHKZniAQUaC1l3sZpN3c
ONU/8NFFkvXL3YcLaopmIEEeY8M9ZcS4iiEqi1hSFzPsvZlVtRwxV2gxSrQY+P3Q
GdYtSEYdvcRnbZ46lYgUhP7+EjGpkb7K0pSjFX7tuAWNRpM30R2ZQvDO6LWgqRQL
0lOBx1E88oMUhfWovIINkh0nNNlMtokKR1czCYNVJVB86puk41W0S+Xk09cByrQN
nXMFkJ4Ir39Ag34MixLMPckq4LrcEKJ9OXFCupK3nFJ4IAIgKIA7hwaA7Ztl6oYx
Mog/Twxgxc1FFL80lTOstCm2a8BL+G/4DqQJEk3UN2Y9KIHg11smc6GaWWWePgNP
6s2wQcCXtVJAFrCSHjs92aKQO4cxf74doG4EpuPs3euoqmC96xdDu2YQdN6Z/F5Y
PPp0QuNQ2+iX19YAtajZ8aiE6shH3scdv9a2iKdWV+NlSEA2Kgq3VnVaL/ny9+Kr
OAHPRAA3GFCvAzWCUQdXZgm2fPqjOt+t98RVypATv5+lWRd6FhrEZtTym19SiXXi
Huw8aHaKds7YdzF2WYFhYdB0Y6Viraj4HHLGealMMXu4QcUjeH+obKDffySaqShN
pB9JKn9cq3IcGv7NvvdUq/suWFHHzgsC7X0bHXytVIlJFgGsTw4K5/m+qmKREg66
9prS4OBaBtGEYmn+H8RYBXkcSJm16K+xhQCbMRK449B3DxvA9pSs6LszWkwZGPAP
Xh2okTqL7iNaVgGiIMGuXmQnEEyDsbMrghPlrm1a2OVwpuF35TmiIZgn9jrBXE7N
Qgpd1FmZLmtV/fZckZEhWA/C9UMJOLEKStzAm5sMMW7SX20Bbui0HQSYV8amQnXJ
6nJasgRiQcUH6laKk+dGPMebN0AMp2rRFX8d4KPBnyzqVBOx8npfOTszfebU+Z0Z
jyNP7U+siPXeQ+GncjTMOgnD3lS9gE6ZmjNlccJ/G83D1hp+ZC+OR4mUFXhiVEsQ
Sy9M76Pf7cfAwPgvdBgcLnd/ofneqjXoBSWYwfXIsnMcIboasD/WSzlVjvoECHSF
cw4BlcydkNkYtOIhGS4L9bo9jsb9Of1Tni4Vn2avJ7Vg5Oq98RfP0f26AJ6E1B9w
zw+yIL68GpqdF/wXioOgZnz6UPKrmtsQrdKUYdKtY86hQ9xUymL+3DlNLJGQ9h96
9z3fUiFtKwqvOHDQk1Uato+JOqjxd1SF1Zi2o5JcIZz6u31OmGr3q5KYYUWd2SHE
`protect END_PROTECTED
