`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/G2OcqKRaXXqrq285eAHfw6A4lAHlBglluObHBSLbzylCw1sXTRDB1KO4YU4xSHC
845hVMyZvEhnQwqQoVLFDvWHUmdZ9cyGzk+HhXScBGbMVCPiNxLq1Fkg7HZkL48I
8oC2UEneLoB0VFgraYo7JBBpwe73Yf8GVUdXadRW6VtEl2e/a4sxO5vgXNLokizL
qymIT/tg1knesib9mhyqVXHEYIx35GFc9fRX3JU4FL297y7OFrxVIm0SWUkVoLKa
e61YSnC2/jUaum1IhVcmxp8SQqfbD3re/hAwXpgLe8TBDD7NAKgLAzHyBeaWh12s
SFN+9Df5cnBDL5j21RVmnv+CKkFMytqWbMMqHPK8EbAkcoTmb2v8TmT3qc7kZiRp
ICG4Jusa0h5E2z88fhq1vQLHXCqjp8BhevW6uExdPCtUpge418k1FWSm5iXD5dii
5ZyZ1hJ74D+ljb/aRGxKZax13Xoicfb+rOAPNxBD2jDkNt4avTmB8uWsxln0nHA5
eYnPXN/eFESouM58lvzX5gP5dLoqvbxiR/GqhhwU28AeqN1xK+PW6UN28VyVOY6q
NbGhCmDDkEgYG9cCQZ0+juFenEU7nxhI2Y394YFWlk6WRaA636hH6bboerDhkXgL
Df6Lw9rQQfvKyg67rgjSc75a4asG60KhsU0iJ2Ij6/FjTpC+yqHjfUoxuzqrOpWS
TeTbBCpJry/mV7a56AD5Sw==
`protect END_PROTECTED
