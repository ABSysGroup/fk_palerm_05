`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u3V46MnIdxKb/mrK7ku4Zsgr1vOenMc5fRBagpip6FMRrDmYsp7NXW2XSGXgHNk9
AC8ss4uTOiO+HWG30ug8Awqk3Qi3Fd7fKM/ARy2OsfF/QFeh0gKebIpseeM0l5Ef
dZCQ23IIxkoYgogmWD5j7SrUeXiCICTYlir8VT16wXvWvx3G6O/JdeHAejWabjcJ
y2iI/mzYNBInukDlmVyL8wqevrO5HeEDGi2qWX1kud9/V+7yFO8CsrVBOv/JBg5T
CZB0ciKoZnj+4DPtcwP9IAwggvdJOUd1LD7nAMkcr6gW8X627KJXGGJP2wKvHU55
FBy3F2YikugrqK7uakMa7e7GlPyyIqnH19Jo9itjfQlm+bnGDn4L1+nqX/+yw3YK
SZHBYpUPyIaKSoLIWVzM+f1h+Xtyag3dS8ZrrXVYdONSP+sT0Pukms+MS6K/Ugu/
`protect END_PROTECTED
