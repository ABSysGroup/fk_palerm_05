`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mwZMA+4TZxx9L4YFluH+Pp9KoVCVfoioixMate2HIFZqU05pWxSznLufAI1Vu28F
4N9hyxFb7SejhFKZwDV3qtwUUioouyK3KcjzNV0Oe27rCSl4TAD9lC5r0lh+EM3/
2+w8a9Sae5+QmwVXJ9m4xv/fVuIXVN9fWdu2xuapHMjCfEAHgYKv5hj71H6dxm4k
Ecs+bULSc3TMOb+WQkzovkvwZs7z2eQPchZ93Zw6o6BcjYcAdq3LNdQN9KkIVW/P
0IEl/xJz05GXWgP8QTKNrhX0hSDhiwBVuem86PYYpvgSEjruEiGd50lLV6YsD1G+
FdSOB0nO+8cvg34T+aUyR6aqj8JjUpNdNAN1LQsWqkNkoa+tS1mHHj6jHESxYdCg
vGiQrIK2KVkMWyY0sZQuCjiuwqwiqZrGSunb8DfVq1tkzYozeS3N9r5sJaGFCtdO
jS78ZpTR/OIZutozWf3KQNP9Unhr1zO0oPfgb836UXyGdO1j47co4usKBLC4VFOl
GM95YjhWNg1WFTbHlNghqOkMYSJNhv5SyvIXQss5KZx2g6XY6unTrs/yXnRabEzb
fi+dDPez9ppQbSpylncKlYoQo8PVMxTOu0fGKwy6xVC9ZreMI/3EAniYIz2h5zZ6
8MrlnTCdFCIgz/yNXTg/KTxMWYIh6A2QjRcICDJYBpr9pQf0YgBVhdcKaaWLEJCa
mz9MB0V26xFB9TLobPKQAOj3vkW+8lnoY6O/1LzOcQfxjCfF7hgEkx6tTwnjmwH1
hsEqLjJc+Meh4b1GOL9LHhSSzzY66D6X1lHAXNYuTZanNdj0xz2QKAopc3d7+XbH
OT5z3LRQgkyL8zQbYeFnmAAof46NkZ5lPIyy/P+JezI=
`protect END_PROTECTED
