`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wf3zvWWT9OWys/hwBpRRubBpgJW1RitxHxexpOsbjpThozT8ZIONCjNq1cm3n0s3
rsqATHcST0bVhDQ3Kz6EQjYY0y0Z4ktdBI0WCTa699JIy0yhd7IBG5K5FGOFEh5n
nUUwNotiQeKppYdOECr40uft88/7LxRWotjyFFwhctmMKQgo1eVRmhEpt1MlybY9
QMpQxuk5FtV8wYpfJDDjqLdAEU9JB7Ye1k5y2QpEgI0V+dsCMuRTuWW2C08fBUTk
vX9ljyWqSgwyHxYS05IxM+eA0kodM+V4QhkMFg+T/bzI0cqO2p1OxoZo8wegDUlL
24H7bvqMs20j6V1wBOBim5+ugkrhfSF1xd4fjmjnapocOhW/j/fozupSWAKdJhcY
aRGtzGZZs+eI0H/4wj3O1easAO5fGK8r1SPZjMQg0IhKbXN/NTEy3fHIL+PZjGVk
bCo+pm8l57QgTYrk/DUhU3LUZBUVTtaoXF4lZ7Vm90TtSAKik0WxQFdYCOIp1KJl
ofPwxo1hqplAWhvktZXCMttBM8ZGPDMC4PuUkyoa84IFJTyi0E2shZXhwLvVvZMF
r+V7CeG82HKjc/U9YEuaoFHqrnLTxt6ya2PK5s3YD6Y5trtax09VfrSkfoNrFmnw
7xixyJzv3Br2a9f0X+YTPvkAm6oIOuK/cLNDFo1flbyrSGhzX7EHBqs6J3mydXBD
uoE23J8eHcqgyWS/0m17F7JPeFeNJxfJtdsGXZ6u6tJcV57qbVC6CdXjz4crUZY0
A9a/1wB9o0FUQ8LwZUadAeq80CULsognP0Cvnq5OtoV5AKwOuRCDnqzEVLP2LpM1
BfJ6ZxLxsf3jUAkVKWbXuTwiTrJnWjelbFQUfBcdr+WJh3CQ3JSwINYcxsPupLXm
NUnn1m9bthdcqRO16VJc5PL7RBfiiVM7csI7ibhps0QXV9z2Lfyb6bo42Z6K1do4
O/999VCt4DXaIRh/NxNkW2dxpwKH5fQi+rhRzixrCBHZ27zEIod+YxtnAfdRdEru
4LD2b7FUE0Di+AYDchO1G8Nnv+2QIci3nlIpaJ2RlJU9tfyU02Et1Q9xJIiNiEdt
GsozdvV92z2RiVw27z+z13t6qN2AcGle0HwzWCAknzV2QY2aD6rgAZ8jgy1trabx
QZwjbSvo879JNL7SbTYrLeenJbz5VSLtPqkxrs0tuQx56gPqqlDzybD87+u2Hu5h
VRhNXRufudZdZ5k9iMkwPmjiUb0RBmdzQTy/UIX+Yb0n2ngxsCh8H8JyJ71l/kOs
n7twL42UOCMlr6RiCfffNw==
`protect END_PROTECTED
