`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/jXYEI0zDctxrUBTQJURSpFMXk46raWUz6sk9C5OjPVgg8lJi35X5p0bStI2w99u
XG9XOIA/26ChN8vKtx0xsHFbFmTDpblMudSLrdXFivCt4X2c+XpO/gFmuY1cn5hO
bgd1tnyTMQZrf1W/hzds7B30iljCb79fudwBvKdj3M6E/8Bl5fdV83SSKFhdF2Qf
kB9ON6I7ATDxxrZd3NX/dOd8NYl2U/tvK57KkfNLhMtOxu4g/tjpPU29fNWekdFA
Au/Jr+QDPt2hVjWF2t26/qurP2/IF94Ho1IhMo2SruS1c3OHOPJugkURdbhesxqs
PjfsVe/UwtWbzx/1K7NnNbok5+V5JVABnTlJGZqgBGfJoxqj/chgmTRoHjFvPfgU
+x6dbbXoIzL6CtIph70uy469qqrIbq7H1iqD4IQNuki2tM+0kA+mUhc9xUkZ0u9Q
zVY2Qznqy1aIlBb3lEekI5KFexLe9ZEFq7Fv4q7AzFjTL7ntofFoeaqM63ZSII2A
PAEJFMZ483gxC7k6d0jv3s4IMksM+F2IHOH4y+qo8x7Ky6oHOzkHAYTSlDxcmbbe
4T0DVPyKjDtSfqyMsNO2JMyYSia6GHHHqeXogF2gfMCYMbiQXRNbWPHm8Ni27EHM
jf1hTUMu2EAMAi4nwVfQz5c+6iM1Oe2v5hdJ76eaErJ1MhB3mmaDlzRTWyNoW1l1
pkeiGAjoOKz4McJ7v6LbeqY7r133wa9eS/29LiN0oaKxrm7OVkP1xqPeZombzMnB
0ClOyyOWmCuABAe4L7Nc3Ac/z8iO0n0o1wtQ9x1inlh5fS0de+jbkejkB2Ikjujt
fDxrTL3aZiu6t9vNuxU0zV9UhmfVspxfoJavNj7eWhn9WKVY8kh0/vG38mU87vf1
G0bppASGe7XxTxggTUVGE05FIWZ4AnIuK2j3AfR9jConMSFwzPJ5fas5KIhsK9KA
`protect END_PROTECTED
