`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A/jVafW2K/oHh3pk1qW199i5GA5MJrw6syrpgKsXmJIxKOcod5ZHZkZXTQ5Kevfx
Xtfe0Led/epKBv3CEcB/L1fZlZd5Jb9LuNeqQbTNvgx04DAqeXMVQGCYjOROzyXI
mNJm+YUDL/STyrDjDgQUZ+IIbYAAm//ghePBP2aCABkonGy+xu2gLT06BF0HOKsX
NkvXo9swckEuNb9anRzSXl6Bv03cd7zh0DURwavubzj9GCyMPK8ixt3tS41tyG34
s7dK5N2Mhd42RUg4A6Yk1Q==
`protect END_PROTECTED
