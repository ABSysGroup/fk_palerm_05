`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A00GjxEPYlE07SWCRuqvLzJjjPJvt7MSVUulz2/TufPTkBdBGc6GkK9ubLOWRTgr
LLfTubvyYd8301iUkSMq3WbeMUHHTRWeIdzgCx4hcnikgJubVcmB+I7fd3GOw62K
JlfYMq7CGCSL6A4B5RDaUlL4wRTLf8ePOXwcbI1/upXlcCg0c1YKvN3v86/OUkIH
rmY2cGq3kdqap8QG0tQeOfvtn2GsXdbbz8DQcEjRE1r/501VvHZN+dL3EnpgaeqL
byizCDct5jbv9MJKrgXFPA==
`protect END_PROTECTED
