`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZboF0gtPepyRV2M7dNIVu3pUKvnBkaJ4z8qNMkr6M+YFdctY8SFgyeI0txjuAIB8
ibqcTB750TCcNWq5mAf50hIAecY9q6tFEs4wm7Vw8r76nib1i6poc5J70mqsZ+8B
sEHGMu4XSBgUEtl+SDxK7JA3dARsijcExTCqgz1dFufjL3jSz77a+ZJAMelCPIlr
V/iU6q3V2E9+Fw9EXiIX1G703z/whL6931ftdnTcB4GFQ4s/i+7y8hsJO7fZ1lo+
ZGebSROBeOUkFFfZSaqiFtcu6YH6Qqkvg7IECkXrVQxkKl/7Ap0rcc5hlqQ+TNGb
RVH0lR5Txnyah6+2sbpCEcOjUTK0AH6x9eKdv6K+ZktecAhYz4NFfYn7QQRoC52R
nMUcBxV6fi7JhJW5FTQpwktF7+U03U+O7VUC/JzUzgvb4a9M2kgU5jV7MoH4nAze
`protect END_PROTECTED
