`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6KyX08s9B6qQZZO+pCg60QJXnE7GRwonOtGjV5LgceINT0NvX5jX5Hf2nCQ4+tYp
iwlTntKlcHNgmgyaIBOf9QEezfp7kOMmZDcp4ZtxJ4Vm/jk+duHWTYfCVezYOiuQ
xWtjbyDMNtmzkTrsNN9/NYGntjgNNaB7kUR6dkss6oIaiyAZBi4lsrBIkMOFQ7e+
bixZYkBiNmh6EpJTTj1/5IF89AUgE3PfSEipOpuDSyqN1OOPsfWP5kvul1sc3Ghv
rI6sIsVSQKjL5U2IWlcxOylTjdY1KzzaWTyZ39d/kZS+nNCqCR+cNqbenvcAyxNv
LDHU4MUROFCDWzc28yEAooUp6vxJCriQLOpUE7Kx0jsDQyMJkreW7aL32npo/gvG
oF+qXAW7MJ8UqTbWyGMNogPkzvVkr2JUff2L0lZkYDFABZnQINSAHTrNURHsh+/m
iiElynD1IV5HdmexZdz3azG9eyzpMmqzPErFfXP4/VuppiH9DX/NBtVAG50yY8tK
4SDj3TSxbMOYwQYC9vn82EdBWEW4asT/WBwFzcMX43nhoVGZD4mqnAFrJ0s0GPr5
f+JwVAnhOwSd6CEnB5UrODAwlG759Ggzr0QZ7i11hz59WkcuVsbI++G5V9pSGyRQ
zxIeEEKiZ2cIuE4w9nSLeoYbjZs51G5WmPBIcyFlWANGLYQwg1S0O9k93IyfHace
MdrWVh1JYwhwJgjZBwA08SSLk+vBM3+9I+JxfN/sOgPyxDdr158FH9mM8LNkT/Uo
Ruap1KI/+dCjPSygTC4/CI+n1fFVYlJ+JOEoY8OGiEgO7q8SoKvu2B+6AfixHQ69
MnsFMrZUsN5KMrMhQB5gghXfQwXnYF2qzYSDE/vVlCuhOnkJFpt3GjdR/6iI7YLE
zy/5gvMKmvoQqmjFvQrfvgUKlZVgZFquxk8JPJDfAbgIPN40T2Iwy0KWB3OEPwjC
`protect END_PROTECTED
