`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GJLwcVHYlJ35sFzuNEnjSbhC4Y+LkOtZtjc5xCHCkZeVJ5FATrjIhXrxjcwTXfTq
67L2Ny9LfTi5kpLGhgnIXiFO0oG20cLM42ZSRRrK/p5lUVYERR6D4Gpcg/htkSMk
Ig00zsnElChPvvS45pb5hwitGsJyzJm6gH8R32b1DyRLd0WiZjSAWs6e5C+wptOe
o2LKTsXS8+PlAVjoEpAy8dFfY1gJB3YqhRGQ5Yixz3HTIDEMEOn9wHA37LSd7dpd
hRhInMDbdBhVOXFZPw+d0Gk46933cFb2fT1Jts+EK5cemXANgrPZZSOu9U/LN+JA
OyhT2lBxJDpmJxytHhXSyYsrONKHnujTtPdbeUtHsiCZRasXaehtWVibwSW7Km4x
UB8otsUcMXvflToSkLd9nYQOeb0oONS7mWvJ80mxdcqFkaQJP1IaiSZ6pD8Nzb7U
SVBCnpstXxJDNkF6k/hy2EG9HywJ6cTjb04GlHq6Bo8DvZh5d6nj7J27o0AKalba
ObYlEe01zFQBPFy/jB2N8nDtf0GhXERvHT1DVRYQykOZuYytwLkALZ9n6KoPzMGe
u7Z+Un2wiorXTKoU5XQLObxiq/cHuM+WWIXEuRAtoQfOZM5KV2Lmt19YpqNtKBQa
my5v7WpIunAd3IpEQE6l1UgwyyJ2f7ZKO7XYClhjLYQ=
`protect END_PROTECTED
