`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BGVvD4RVQGh6tuN7kyX8FFcDB/BhTU2ZtkFjHNsYwrnnAbPvOOcF5GUoZ3oFt4vY
w9vQg7q32hwr6jGj2KWsTzK8CrtkKSuEMMf62aMLh8QsXGw1+ZsqtYKEntDsu1ls
+UWnESjNn+ujX0jqPaOdHPamE0HRIkals+8+ja4DfjFUghe6pfF4EqxSeZ0vYDUI
BvE04PIy/o21DrpyK/exhUDXRBGxuqCXyYOHaIbvOAspqvLGJlLXXLQWO7zwgZlD
3QiNZi2/fVreXLNCKDvkVQ==
`protect END_PROTECTED
