`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rj/ZpUTJlMQXGEYQA3kZV2T82vr7QdV8D8/0W7kuH3DB8mqvHzS/7yOHZTLJmHpd
dYdasSPsRhyspTxzvmyJy4LpKECoddCL4N2IAMElioWlgDLXVDy49bM/FihdrOsH
6jZy2dDru8ZgHEorA7T5EGQ3gFEhBMNYKX8eGi80slijCQfPZIC3VzVuQJHxjX36
Dl1r+fEbqxn+2iCO7zhIy1PKPIxd2I7yEzyFEQQNO3/wZA0biizvvRZWKlGkgrii
2pCeCSrUBgPs9oX04lkH3OvLN0p+cHA7XH8mio2JfpzwBBNAh0dC0GxLMzdXTdxT
0ZPr1rhmF/o9Yc2dR8t0Pygdr5pewnEuas6nSzYE/GlC6VaimJnZbUD4c6mX5wuh
`protect END_PROTECTED
