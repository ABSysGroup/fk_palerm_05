`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mI+E6WqZVbZoRrWnbU6Zyht8irxZjPQKW7WJ1GkZw5Th1GL7Bd256a15sSRW0Xzx
2xNgKnwTq1CyqoAGNTYwKAePOH5L66dlzai8/rx0U06qToU/z0YSZYnGO8a0B9Im
s7MYiUYlMvfrtTpDtKGLyRSO5Xb8SfwIHkyWI0qVY94PzyL9qwHvec8q12ISVSkd
IalwAftWkOI/kadtwveuwSlG9UarS9Fsy+R+5q16hupnunoHKIPlTwa5dPYoTZVR
+VfQ2EulVc4R7V+qUaTL93aXIJUag/CWCsnJfb5LI2e4vMSjBlIJN5jaYgJf41yi
xvzIXCQlkWvTYbAO1XK2LOX2a+z95Ga8zjxri/vTe9tPziffVPswoHlejfhBWdWl
nSt+LdXyYyKfFBGX3Y8zUSJYg9f+WTaSHS+ZSD86jOVTwdAFn1tjjOFyU67RTmBe
4Ra+h6ruhyJGKEC9AQIK0jMHqj/e0EjOlOCKZ4pOQzdR9Z9A0PY6sBnPJxq5tZUx
aaWhID1ZhTzileDgJIMasEUXqmGqJPy5TG2QE5C/WQE6FQr6BJqJykr/Im38xUuf
EBsOOHq4RYqlh35NKbGb7e2Ulle9C33xFYdz5Xh+M2ktBpacDBRV/NDwO8CmmnW3
T2NExT0K3cwaPC2ShEwr3w==
`protect END_PROTECTED
