`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CqW/d6eogrmePq61/V1IyQVrNm/BxcvOT70RrsoE64cwr0izz3iejF/WYAfGPXc1
rNtEiOarRxZo6BGqSNx6e5M6jEn3ay9E0SuIx988csM+r4T4+KakOWub6zNPOkQA
g95VWdbjBJEXgIsDSsobPiOmfg2NfdCeVrrdAJiUrpglX4fDIixbxiOSXehWJCqx
zXHozjnha/zM4m3CRUKNP/6XXh8Wg/qURtQ+NI9NogoaVFM6nsF5utTSe1w5jqX4
xtQqiNSHup86GVtCpig0LIkPI4dvqAE//2Fzo+Sf2kxfL6zyHt0vaT2PxpYbjd3H
20/L6Ijwu3WuC0GUH01SMusidC5JUph5Tm0gWB7OumhL8LAxas1MfmTTR4WeGjXL
Nrs+oHkQB5oL27fCQOfN/8RMvnOtqS2E8eG4acGPqL5lOs5moeqlC2PF7Eq16eMI
VhE0+FjtclKCoSqRiDn8LZm16ga5/iCNgdiZD7HuVgk+TgwCbI30cCNtUAATINt8
FUn/Lt6Y3RZ7728sosa//ZD3nkD4h8rxwsWl8jrxunl5Zyk4Ah64cJZM5ZB7d59c
kFqNDyvN6aS72lPIEFYEnPxUp65oqLS4fcrZDevLo1KELjaT186V84EPT9fO6pFJ
L6qYbDu6k3jAKe++4Gr1vpDwL7bK++nhPlCHVo3Dr+UPgiJ3/rwWiaCEOgJ6L1Zc
MFhJPB4ltkVJFDnFuwxC9mfWhCt/gR/X7pfz6bi5gLzB8sRf9NJiWd95zO3oLfBv
VJAwnzw3urTuEEJXY7/xoQsx1NSVTBzc7T9DQ0RHQzmr/CgzW8j3A9xF5rc5v4OJ
y3g1hIVqhDR9b/v/GjInSqCiMsyr28uzO3v1edba1YNbHn0DKFcDv1/g1/lIn4Jv
+4S2m3vuOnMNm4lYi6Ks4hSXdoLSmo70x7x13hyjU5bzITLwPjsOrd6ImiQ7xlzd
2LqLkpZkkIDCTddYVXdb2iDsuLZiG91D2WwHWSrCtnS0vPjdGyXNayifw6COuBWf
uRbTrX1w2tMs9LhBhmTrVm3ZurWqkxRr0Mg6hPwsXBUU09FKXxbIC6TPqOnWZmcF
1Xyv9IfW7ObBJN1jzj0wKw==
`protect END_PROTECTED
