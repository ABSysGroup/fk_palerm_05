`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cqd10K5HTyVZr2ldQegT2J5osikfG7D71ynbtvCVQ0y5ZzzG3eUaU5OeEMHI8fV+
ktVUXAWy8U3+onFkD5pzeSeyBZ0brdg2oJuVHWxxMiA9fJnzAHj6iqG1HwyPtHxO
zIhllxYjj3B+krS79vRapI8FA12z6m9ILwbHstJSa2oTWkl4bTeUtqt4QDYaKOPY
9seS7gGi9RfbBgaUOqHEADGtDUQ+1HS9i+TNTnEbD32e7xLMabpg5jwi7NzeunoU
/NY7uLwTDdxhAK72xV0F2dy6FWenV0RAckCeEURlr7R/C1uj422+I+mn9QaTUgdU
e6IT9UEkMbCOAzIYc82BdQ/rBmxL+Jki2qxcwaMFfp3JylDzwfT00L756OuHrpX5
HV1L/bUPDNj/JZgzURe1dxuKUqP5hDj3blZqB4CKL9Z37pq1LDpYKHshmQ6M1ueC
bzHy1VkSmqlSil0ihmnhqYlD1z2lmeGAYihPE3y0U1edsjOG8tkLj2uxatCNSClk
yfWPeGIxLFOhVHtaAKcGV03yQzvH8LIT+R+EVN1E5lRpf3kHobch9SUQ+h150QRr
6AhQSIjBfH1Cx6EgexDcozlL1u+ZzbO1xvnqqmpKNrkbe/f5GyYr/WYMnKEUMT1r
1XM6JwFn7LdPHMM82EOLQg==
`protect END_PROTECTED
