`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y8MtXWoQRPn+o/kmnUqlox23aI8qzUlTbCySfBrxQ6u0b49BNr6i/dGlpjT3URpW
NHI0AbQjvJbx/lNzELEUPHgPZAWLSFJToPdLySc/ZZhEeAI7ZYQp15KBveesMqVF
uuJ2X6IAn8VlSGwbOtEdTMj3t7kIyuVcBQL3S+JmJx7rXVmSZ/G/TLrV5yPNqAzp
+WWb9R35F6XSXxslRhY7fBMMm8JEbwuR/abIHBkeCCzHy8aPhIw3MmWB8bFxW3d1
Q/Kn87DgRNe7bAlvAtPhbCRWtgUxQxukXz2PrVxPpwIOXkD1kY/SmfRA0XyHsFTI
FBdYPvMHliLnsiSVQA64IA==
`protect END_PROTECTED
