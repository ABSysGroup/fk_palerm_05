`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V+HLqIsVagEElba00yxDhZcpNeKhaKtdrzbiarZoX7CCAS/Cx4g+RCdh8krxjKED
4U6laWFSgPPHTwq+ANEDo4AsbXZIJG36FlvejxQA0VR+A/W8fcRxSI9YPrr1MGwD
pYXmJblWjOocBbAMwCIf1BvLupqyb3Z8K86HKxVSSCyTm+DV7IPeKphsf0OsDdAM
zDpMt8vLfQsFAX3at7UO11IjEabuKCGoDxyeROhcMeyizgiiFrsaPhanAdoTo2m/
erTIVGSdTez78HeifJGZmtzJAa+Hdepc6ppUSSYoTZmUQ3JWXe50HKMrh81u4qsg
uPEMSUO0i00ICo2LsvoUaaiDDcWZyXviUqURtQ/9z9rJwvp9qi34GSjofrJVjdNg
Xb9xbmeYJjQWiGkhtav94joVK6REOuVYymg873cowijkWSszL8OVGq78aFaUf2Zw
YLAaG0DqhIAtppI82tCVejuu0S0+duziZjLjAk47KkwbnrnCMG5ectOtmGZH7Eq2
JfHBHXBxHGB8xdIEXDObP7miCDncVEer0lKJEVipzGGVeMelvVYOKTJmaMgVfm3x
9BGeobXuUcGYIi5R9MkuMQxRM/GSp/yw2/NLDDdRSjWxTZoXUh09jkcW5WfV2Y62
uApg6CK5Z6Mcfq5f77gp4SiFm8eHXRw0o8L2Wh47r8loDiezeOzO1iRs5lzRzICu
gVo/HlNVikE4tJTj74Y1VxJdbM2IVOgG83SqrOn4DEacZrU/yxTXbL86zQ2UoCd5
HCQaY+Nm7Ma/OopPbuibK33mWY4Vf+JD76Zu13j0LdnuxBI0yOhva5PQiLp8wCem
fhioKxaq8iXTXP18w91zTDPB3bbl6nW6LMSoa7O3g58COr7xBOxx/h/WmAHMyrMJ
bFwcyju4O+eYEd0D91Wz2L5AHokssRs5D1YPaNGZRjSbiR/DqFzWdGsCgZ9lEE90
nUlFcNpYrwGS9+QDnrB2J7hJg0A6sM1CnMjnYf7d3YdLj76Q2TZ/coq0iEOXPWx/
0L1XCJU7/Q5SBbvbTbWPF5SIvb6vV7YAl/kfH5o1mkNDNF2iiiTQIKWxslhhLDV2
TojQM7S3oG42XyAezMOymMR+PBwaY9S/U5i2CZSG/vOwbAN+MrA6bunH4A7YPtz8
6F/L+CWPSs7upIZqMZrIe+1uZy7V3QySWyaN2WOKHKlT6XnwneByt0JWDP404V4H
+910V+YN0im/vNkPKKKQgZ+6PkoxUwV7vLyjwXe/9m6Bvi6+WrnCM4WogEoT/8+T
IXfDTq0bUxian04KKSrwB+lclquOukBG06WGPQORPYpTkK3fx701+EmYDHB1Y8Mg
fC5ZuJyrNAEW6kMc9xfDToIWwIvzFXpQoJkvBXLdP7UTPXQBQigYVBUHdLNJaobT
MFexP0dvKkhqy9d56HmSLSlMoU52JMBpVhyhql1Hs3z2LxSPbyN8pEmH2W+MYxmd
lrxUvo9Sk8kjbQ4EKj6zk1oFKLOjVt8hIfe+ol0tegVLmN9ORpDxbzacVKBml1gG
tc7GMLg073ipTHUOchEfG8ym/qnDch+lA22zBvgJQgjdV72NFtMWyzYCmXFSb8IZ
b/nCwjbbwFYgtA+btSfqL8JU0rj+XJi3raRThsvVdDH82ACtRPRHSDDH6mAd9Wjx
UFDhSCZFpnbaq5mZgkJu1e0/Lz3BsmyRQty3RpLEfVJt59qOfPLZnwtbWmaVw8gL
y1RewagetwKeJ04zK7iobSpx6rivCa+CWFwQ3ax/iRPWqp+YnmIiAUgHBwdAZEpU
6FSc9tc4KtBBMOnY2HvC+moL1/F9KB5ZL3AK6+jjWV6KjHu1qWSrEuP4ZKA0gg2U
NFXKQvMyGqReGBCdGai5nKeUvAic44nz0R9IcOwldwy8RtPsXm8K/yxgk6byUS5a
PA6YREQSXuc7dqtvI6ndyrxbe48F6pV3bf8DwoQMIeInbpMU5BebQHseKr8Geq4h
7cOskwRX3zNw/5Eh9BXOGZcpc4qveHJHp0gq1PI0ioC26qrRCTkftpAtXCClBsQZ
KWuWdcBJ+/JRBrv8rvTD+W4ndr8nEKMsJ2chnYQAjAZdDETfMqqW/FmFoIIlOb3P
dyZ8sx13r0tsqgXPssFPfH+QmFJgGNl9wuSrvP+1KPgCT4zuPscHmJ2wsFmtgCKa
eIx9ej33DqV+pmxRraLaSPXYDKPr9dnd9Ni+MBJWnOjvNUQSghdj9Inh/eZ5TNgA
kEFmR5OEUM5GnX6BVCs1oveQuFpXLBqHelAqt0adU70QsoFDWwyGTe2wSEEOxeJy
5LoqOgZppbvyrMfAZKtcqdNWMwbnoyrI2rsjMd+q5cCsecm/CP04Mk/ORhOhM9v8
AZiRrruFX6N3K5DSJQFn9dSuuKReNlsvDCVpCQz2QhtMsSHUXb5LJtec279NMmfy
oTANC0fpaM7QjIGnN47x/7SBrWryI4HehRG1Caid1z19BU6sGy5M7C1w+aNVV9Zs
Z9+fD6KyKN+pQUjp6q2YV7EZBUQw5+n4lK4es/RkiE9RFfNXNbd860DhAQWqV/lV
DgiZScLMF5qNq6Sr4n5p74Q/s835coev8QbTaqqvMvgErVBF//jUbK4AR2ZO8CZR
vfV5Cx0wEE7V0u48/+VmTqFnDOF+aQ45Z/Tx8uhSN2LHqBMHnvVhNVsaFMLm4LAi
B/4SbIvH+9wBS9buxetu1Vy+ynEA9UWQu/mxPbsLvqUFwJ3gHuYPz/5Z0O7kERQ3
FjAzSwg7gf1YarotL/wHBnyXZhSIVTPAwoHCB9xVw7V16nrV/Vh7Ui4yLdGXxYdc
g9GkuR1rWVMC4BH6l/C+xbwhOtuVfMGKdO2VnAuc7c4q8q25fbk8PKF6tnu5TtK+
JCCmLHKHWnIf/nfuJRZNLoF0gS1hWfo7+qh0qk9Vs8f5c0F1bLmvMkuBOj+MfbHy
21yAKaas7TKJHdd1NwI7beLdHA/N8G5Nw/lYcaETQulXpHsXzSmC9Iue6sePALUP
BPHh7HoxhvSeT72+EGGeUj897jr1TaH3uEexHcVf2okmzQwP4CY7uqwMNJ+xHbr7
ViPdWeKZTi8rvJ+nvf6Eui1f+aKDJ0ndqq9nsLaTr2w3S8SWoUP96pw5feoDa8oS
bOUh/8Buq+/rFJVMqHnWnhWJ/u7ms93nro/PzjIEOqR8vu4RB0KPemnewVksSqY6
i9q8D+BcROsvHFzocimBWZKgClz6GSPd3hy5YeuMeISO/5mdlRaXiJUEAs4qRbiA
OuB/vC9mstRXBf+PK3PLoA9xGPcI5EHENk0g0BsaPZBMwXdBeXvzX70Xx3UK8ltW
lgTxHTE/WYGCMx6VveuS0e62y00Rt88NxOn8g2F8LtIaM/FRNkSv0nTScBJICtYe
XowtimESz31HKbAZhvbEEqzNF/ypLdVnWkOw1+zaXcQ8RrYH8bqpEC6hDQBrIKKP
mEoPTiFF+2LAxs/OTDpqB2vGdn9OCYeDzpTzJ3iwqr1ultiCGpvz1hC6kc2cNi4P
f/0d9jBws+OShJfbvZ4wQoedS12VKkfN0rTZtiHLXUtrT4mW4CibjT/Z4Y5LI3Gd
1+NH70jThM+W1Zj/jH+lPnUhEvJaKihh7knedSJO+ThFZ1MMWStB8ByJsYJPGZvh
nhsqYqBXtJlTTHIrKmKZccUYk6x35N0nMxBn2vOFzr9/+wAVWF7JEBS9OAKHiwfj
7PQMRvUgX94Q5Eh8gO9rp9BhK81jSzwVFV7rPhugt5h2axJJu1QYv+l3+AMx0m+D
uSUMViS4UHvAeTBxCdSPSpmiSMARhQR2aBN91w9jYeTIEBG/8Pc4pdyyJU29fvnE
lJK13M8TFF0fgn/2hwwiya1vRdZyan881F+VM12bzyx9UPmsMwS4QqQbrWg2TYVZ
7UoEduiVeBtBMq1epQ1FpBiHx/8xgq32ptznvgm2JW5v8BOSvCwiy4bzYIs69RwW
vpJi6/43k1yrSZjs5mbpOvC+u7StKfTidPzbT7Mxhou833v7Cr9jvZI12V/LM2wr
swthbujAn6AwLjB1Mnxq7N4ZNtxeYA9rWq2yGYBRRTSp2xPOray86uxdniu3edZT
85ZGSZx5dG8+rlMqCD0pDDex36yLby8O2oTkEFRdBLna3JTl8iPQDndkV9FgDK58
K68egFQgHaKagi8QVlkzlcYGIUtwJC+vn2LR4Szs542pLy7l/vfuCL4zyKw332N2
GvGZ9ZbEZwETM3sRzUHvppab7pjEr3IU6gInws3OxmX3jX2/QQdpsCOn0RUtsMAd
YoieW3ab7czsF5vtTM50x39xtsi5TM97Nbq1/IevtzeH2ZYjKdqXFq/gos7dvTRA
HHD3ILhK/3rv7RWenW230LUoTNxJdEX+j4Y4RUMLLFgq3TUJkJ6bH5KLqcyJswS2
Pu06jY5LIdCHmBkBR6QzuFWr4YwfhT6e88L8obU4Fb/MSWVcvtHF0IDildfk2x9k
ZejR6sv3j9QXqfXbudek7mLAYavX58xbaADshVkqxROndKtNHIi95H+ECvqMrzfy
Vl4GVStYt+nNuH8ZbNxA8lAbTBzPXrqwJVDiIm6UidO8MYq3BpdhWZpgWFwI1jTN
L5scZIQqs8TZBrLn2UQo+BPh+E4R60K2EuPUnYPenjGTx3rgGzLqQPvNkGPD/Sgy
0EQMmK8yM+KJqy1vsav5TcbqQgAH8fobmcxoeM5lxOKE7rf1EJWaAlLXGOM6+1g4
XDU5qz956gjbmV+UC7w0TPdvB3XlLWVXXfxMImjkI0AFdJ5Bl+eCeqLA7hPbcxvy
Cdvlc5MO/u+bi/z3xNBgF4PfgQyzUvY2tR/yW9meBrE4AgcUbvV3TgB9Te4PwCX/
8SzE61GTgbwBLTFvLajeVocc3hIeXRlC2LIM+65HYPFzxUJyKN3FJHZ46RpPHFcH
coDwYQYRWIUETlkLr9v4+9WWy7D7Y/T6yyU8hkgB4HFBX+mpHKh0Piqco8Q7KJRC
sBZP9CSYKwAZDNMhAH1JkZikIvzEKpQRQSLUNB3BAmrbcjpPqJsAoyM1AgMypw/1
FumBkgCBDPVoG0nvq2WhiDa6/YTYnPIv2ZqS4bpcjjnCdAoXJC0q2HsZSr2rAM2H
xyZEIwWJ7ksvc3ghvmvQvBXCrk26cNe8bnTdPeLLai1T/JJmF9Khd2iX9SwSzlZW
aflAnsQC6ChF9FrpkH47+ADzxJKe97Cr4XsNmDfd6Ltx+o0YyayZVgMus1Ds8OGV
eXwNfBCN8iLP/34z684YEN9nCmnpbAhpa7tOikiuBz0Wf7pWjjszL3QW57j0A9vu
ywzfn1mWVFJbel8+kAPIgq9JNIYqvHQYoFDtQg/tkmc0h5dbTPnwLCN6DDJdPj7n
D9pjTdFb+8Qk8OAU7dHZ49qJO9J8bON4zzJHBxTON9MgVkI4XOiiSxthtqY1YdpY
Cca/WLLJ69gOyLsXfW+F+R7QYPI+ByB6meJ2nnowEbh4wAb548wrBt7aMcBRfXWn
4ta8ONqVzZyg2N8WebATzlZeACEvXD/t4EVrJhqslMA/J4pGxClujp1FSB3sY7/F
mdxRaRSN6jJn8KsFV4keYxMj8Q2ioBglFZ7bJLTyjghBVS+1DxxZ/JgzVQnhaIY4
89LrEbK8O0kZluWnpFyDoWNGeaMUJlMFipYrn3p6cpIYRz25m69bWaE/XqPIFRAH
jGpw39Mj41TEAn2hSipKeCtvOMEqd2K4d7NzmWaZhqhesxoEzYzJriBTHFxpRF1k
zCjh9I8etAgelD7oRRbYxm+LIcyb/dmIJu56Mj6ocr9NHcjKuMhBx8uNR5jOtFpB
g60JFP/Q+1HzbhSoG+TwCIhz92aJa+v6uX3iRJlpdtHkufmv1GEEk5JMYkuY7It0
e+IZmvjQQE2w8T/8kIoFq9kZAQfFy8JqlspMWKk6tNlOqKNrg3wlOhg29L121cI5
nxYbUS9KLtWlmTOyrFN2ESTS4tYpA+kDMo8uo7hSHERh+26LeMBP55PopO6SHoOo
+ze6KAZWpVR2NAOtSv/z5s5TmnNq1bp8zZb/Ubr5o3jw9sckRJHi659zaLB5ipWQ
NkekoW5/Rq7oWhu88KoZWWNU2DA+18e62QSWsOkYGBGJVXkObvIi0ksWOcDAPFad
OrV7DeCY1sfU/Pnqe4GnMXXL6XnfGMdCHa7/6ub+j+wo2wPnHZ2SIiW/QAphsTfD
zJLoogXVnqi4jeOl6e6qYS1gl33C4dOoTiuLyFAu190mDrUou6GwNW7yq3eNLGx+
8BfPT0LZI/iZ54Rd0GJKc3xnN7lNGmN0Y6J3igHYc9BpenJNhkvTq7Ng6pg5ffED
twKKfrldmGm2YGH4nHd768T/IgDNk2wf6GjWTEJZHnB2SEmKVAVqPNxMpQ7mQrsz
9AboD2+ttMIh83l5nHkhjB5BweWJOhQXIk0A55AbwkcbwjSA9F9DZuw4UDmlE43g
QnVu7GoP/LpONcMib/OaDvmoiCAEaKBQGmlK1VVLm2i5WavD4Sq5b5dJ0JLozF5R
FdRdJjuPFK7vj9Xjb3Pw4sFILdT/u2eAjhZtPoLkGUcPJL+/8Gb7KMTObId++G9l
gZqdWhQ6if9W+S2JTmZ1CD5Y83ORK7tEchhCqhwy9mwOIjyIdNARjvy6Vci48ihV
VjjBfU8SnufwTMZ0zwYTnPmwjyP/zbbTYE5mLvtB7sZwTwALkDP3Ai//LJPi08JX
cHwAyv6dJDU3yxzh4DQ4AflA23EvSApuXsdpnzpyJY+vltPcMRxaRxUm0ZtnsrkS
BsGDceRP8x63D4EH6dv1zrnJbAmI2SY3u0DYLe+vU+nmBBwcbRorAmDQfOoY7bzF
4KQK7aeMyAVUMenMAzXqk2ZfDnyJuRCkEqEIE5hcTTvy/Jamd8OLyoTjQG1ACZBj
j6doRR07Ce5deyPvWNbkAjVrwx6ZkdKxyKN8xQ+aSp+dH7AIVUo2aqNkmdCswU5m
B5L9GvQfTnfv4oNl0CH3wEHabCpIevZ9QpuQfALCrztSVf7t8TRA1m+yTqbLmhjn
PFjCPE1OAv8zk21uYjsd6sRxmRPPR4cExTDV7tKZ9s1LKrHBtmYP7RWZkcrqDd2s
HYJomYr5EeDp23fvBU2yVdlxJaY8MWDyhEJ6uuC06Lt6llABscHsmppewbH6t+vm
E4LrB7VLabwkOFygH0vsnEoso4BPLbM7Rj74Edk0sqCmKf908mHBNWr6bpvg8W4B
G4BGKMyb2crO90nmfjYFbDWK6RsYyJMAQ3QWqZ08sSAktsZOfK2ZlrTwuBzOAX9l
jTHOQILTivp84zU7b8N1DTq8R3lpfOm1u3MI4jwJUcJDaGW+/yiYZf0jZZ5ZOUap
nisCIMvM39XKoWQwHX+0Y9aLEqPQndpVYETU/Hj3lSjeP/gphoA22o8gJ4imWjn/
aoTC1PFRiCtVXO8Dv4zwDGtXFQUpavmErztRwbik8YuzRyE3YdeWP4BbE4IbTQaX
6dK/1ajV05GymbB0smuQOhCZFQgJPAURLg9y71itNoN5Enlak1XAmSFg18CJfH1K
EKLMjL0dc9mHp1N6c1sp7W2kGrhxX7iVq/Jd0Wtte8U5Ud2VzToyR50avgYzBLZt
lJlxckgzSHzm5i1bEfAlJQV8WTi26A10ovywc3rGCT5UQ5M+TLD/3pyMAu2jOWTb
4kJdAmJv8HM8rH/znyH+oCialDQ1+X4R5PLA/Mw0th48saNQGwCXHWkX3yq9Grie
iKNHXOT6G7QE1RiYpB2/7N6pXTPpDVN5QbesOZbSljGjg9iagOj9nLH8hSDpzcy+
FfFOOcKc1DQN19nlPUuh1SHJg0FZRL1oPXyAYDTOwDMMb2Euy8EcwQJFA/j/2ovk
2AxDrkRt7/Sk2ozBBLBOe6e6+mGN4NBGhcN//ZNJXA9c8QTiK9PoncJxDcv7TJjN
RLalyWCKBssjzNFvv7csTzDty1jQr5Hwkk0Xx1Xhc8J9iRqwxfiYSZex1CT9weM8
b2AFX8dOSZnoudQSqVakmpbLtg7O+KFw/Vx5sHSviWw07aJrGlbar+US62v8jOJI
BKetKKj+d51FJ1SnxuXiQcaoMNFO8fQ3lO4WXx+2RPhuOQI2k5lprZZquuzpMXui
wwOKTk/V/R1tnPqJY/ees0VZt5oGt1YxqRMDVhj9mRRZZlAr9Ol8juE14vovl++M
8uklSdX4KPriywB50qr+w3l57z8J4aFQ217tElFV+EBUyitwgfyt5gurttYa4X8+
nb9K7syOX32vobu9rNxEnX4ZPPeGFVKl5/PNuGyOdFcej38tS/Kfu036SBKbxlP7
X4E9sAfF1JjA0ALAoWR2DKV/vdNUHWpIphWm7yRtwNwoxj92Sd/G2bBYBZ9fXPXi
osn5SqXkesawDjkgmk+kVqykkDA/HYRtblEjW2OFqinYzu3bs2z6xSPfKlWHuMJ+
uj5GlMqAwHnZbKGWJ+Fkgw34r7pC4KUo1eBOd2RESEAcKLEz7XrkoocXRIIqHwPw
c/IIEqksgrYqkecf/QpG/dqaK3HSg7JitoGb8fiOcJInU/qlsKkBp0S3PCfQAcBx
aeDOOsOAmMNCZxb/JMwe3LCv252IQzjY9fSh8nlw8Klx7WVOZXYzB9OV79JPl5vU
JdFZCFVvWOoEp4bjuGXpE+2GVSFX3C09yFF3K4ZkcHEnxMqsxEm6VjRzLRbO/cRR
6vIreG6WJACAwxyqRy/mOH7wPjKr9jAlf4SfU5CVERC2fsM6554jAfsqoJmVWObl
JlgL49h+IYR4s/dho7QcAn+He2e7ISLKNmURumI/39DXf7wLF3qKB1I2BXsmehL6
1JJC7/ySZUBSi+Z264cubNmKiw+OW2LBSL+tQLv+8llhxHoBsREhOPeGA2GlAODJ
aZDKlP/5agn7sZTbH80tyOiJ0ZzTCKqZsCvVt1v1AJM+wbY8YpUKepeZOFxX0ur2
kJtEBlPBR6dOISOx1WqI2spM2dNBnqk/kXIEtObI1kyIkHsozn2Fn/uSa4tR/xQk
IGeQT0DQjH5NczVpKL6+FJUpAthqsAvju6cWAp7CIraZnENxW5xyi+EC4xC4zol9
4WM8Bkhsb0v3nQKwST5RyzM68C2EJV8BVbNogwf51/ycbur48+MFXdtCNgE/scXr
NCA4dlKz2QT93QYyvKIY538K7YyGpD9YFChXsTT6tcJyXNlNP5D2zSDLYOweSN4/
hAX/5eTWPZqAlWe5KAeOqKt2TuIPiI1DY+o0Q45xEa0jHx7PFHAsPsBzpTETnglx
WL0pgFoxq8aBFnPKlqu0wcl9+UAxi9vfy0cEtk4tBQbH7YpM8gozlDN5Q59af83D
AesI6PGhXZK1DmgBHOSd224wF+WIM5UQ+eTOj2kN2Xv0GEPrqB9uAXh6s7KygNLv
22mScVIHS9FnKPvxROejC4avhfjBrhekVVn+9NVwYRTDY+/Haug6WI7j1a5Jnlrh
5UuMrgeZ0N4OvsaZ/rPzkMJpHwUIlbJKXYxZJEbI24LBYbMu0JRanrU8f/4KGSdH
XNruogroRTU7z/xaP3y/kD0u0eNgt6aUeCFFI34MH+gHqzSN9gTZMYNF5qXkmdbz
gqAhtHtb3JFaYkHnriyd8mq1DotxRue8dbDoXEhHUg4Nyi1v8caGOXtoCd7f2t6v
Ve8KcbMF3zoDkdvegyuBlYlXgsjYEjj5HRIb2RDdmzPnswx0POUKc0tl7hjhjDGd
uqCiV0QpUX8XGbdhNPiDIDTi7HsvA+bRJJ5n3DZJnrCMp+jYsvHCWWJKbJoLtQqR
UgaLFlLVBd4d9z7UKUh5SC6BtPYzHZPYCPE/YICmxh1aCz/j1YRruyHXvmEuZpHi
FRh/ihvNSa1RMFe7AVnOfryFcRN3t1xHe44+LyOjW1RyhasXTjr5yjJeR/wr5VCu
dWgz+x42pFtuJmdFLDwMzgJ5EIAgaEYqLEBKmNlwXJCcrYkElnnbJKcArS4X6ovR
t+mH6ScUboJzyGfkzVr1LqLbC82kotpCQ404zwnHIKlmZ1i1oro4BYDo6zZkKBGJ
UUJZn1KFl/DEFMyclzmrDbDla7ldBEf0hbb52H5uAhaGCsDKvTbQbkT2MTLI4Cwd
1dku2O1G9X9FHkHP66repzhiQXxYn6MRqLqQIfu8XqCUiVesrutbWuiJauwXVZWh
+xeTbUFXDooK+aMleci7VTmXu/VnW8CvrUSps6T6IA4/XGbV9y9AJ/QgA2ty2e1y
ylxdU7vMdapwtAI9Yj5CFZrc3Ur6ycWvsRhedHuc1gQG0FTlPk5Ywk+rN/d7cRqM
kbnvT6kMu5LZ7wBIsdKk9vRHR2jZQ1nNiG3aOSq80e61uqaTjfcK2K/Alo4F7gkD
tN1S2yI+J2yky+izTp4g+BWPb1L18pneV5Lo+YWr/JG5M2gr46nBWVXY4hPwZA0e
pAoXTKwdR+nMqv+6fQDrTsAbQstt9QphWieIPQVMdw4VPOFZzD3kP16s7lrCmF1z
LFznVYxQ2hk3OTypj/LFIf4TUYVNOE2MkkWFYR0FYxc/Kz/XntU1Y4euS1+0M/Tf
rF1hEQLxlUJlJDEHonItlZ2nyLMljcyC2+DsrBHm42kURe6WZEW0DtZG2g2yO4iu
nz+hXQPfNPKSRjBvMjwxTtFPopeKylOR455dKkCz7DkOEu4ZWGEXeNAT6sXOOx1D
ifx2DO+bJQLJfg1z5aRyq6p4SNuUzDNvGcIcdmjE219GGNqDj2j3Jjo3Dj4H8wWH
zMawE1AxphF7t5KYtoIZjybh91WkXWkYLMrzDYWlGpkA6mkK0SiTyAbmImEDFb8T
KHtKU5vn2vkUIFEySmtDv3g5/hl3SDB3jnVxdsB/a6Y68L/96YvKXT6lV50dFpql
qNczyLllUlhisLdZgRmSQVoi9AdwYefx/jgC+mcxxTdCNkwAEDqHEKJkjSfRQ25k
XvPtRqyStLt5NY/1aKaMr08pXBFolsleSdkZRvC+DJDXMA62RjCGEXeoG6sUp7Jm
MDpOihaqUI0fY1lFcGbqbtqRCV9wyEgq2b3B4gUzkB3k04nW0tpVzbuS28fGolQn
sbB5KDFr5k+zhY9l18YB+iUL7Ri4gJZnCmhn410uIuMldN//DM1curRod9YjrDC1
l/HZ9FXv+5ukzX8sQWGG/4aI4WgrntaPEeoYDtPUNkCPg8jWcpLcLOnFH9HZ3TxK
OCaG3+iI+3YcvHCdUZGZn5774hCbjeXAL+seEcH4cvUbsLjM6m1O0YSCqKRzWvzh
Nnaa4tlx+OHpYunzFBiD/pvQ37rtABzfEQO8DzxGfLApkSjBdMQxI28CHSQDEVQd
sZtexg6LR6Ywr//ufr28Z1kY1kAHrB/KmkSMOcItOpIK4Enm8i789VIRuEvFrqyX
Si0VhtwQKb6oQKEK+EVvxpBxk6qa+Y9N+fOE7OfqG/rzcm6asHIG2AfFi4ee99C5
haAe1AUkEO/uWSt0qPH+bu/Mt9LMcgwJqhdpGgMa2qZlT4VjTmoOrKHgd8KAavs1
HTbnUd3WOl3YropIH5rzuov8lnZLNFXb5orXFN+RHIryvOwO66sqhTPeDu1/R3eK
UBXP01dJtkF07yKjYXDyC84cLrJvZiH3yf/Uaw8/A70nJfbHtnImGn+eWe/H4A6p
T+lHLwnXT/R1PLS9CeDEMdbTDos9P7Sh3YXZiJ5McZsTx+zSLkOw5PAy2tMX8uS+
zU3UTdjNG1dTXCcO2hOjt4GfOvzsTDgUEg4bctVtOizTR5B7QyJLJ9V23f+At+FV
Wyx2yWeBcTwTbbsFCvH9gCS8nOn126JASznuEszaajJ295YPuGazHacLKotiJ4GD
msWDl2hzcNK/HF8sqJDWNfaD+o9xYyn/iOe5LkiA1PlcX7dwyzzfZITVY5uN6mWD
CiWY3gDSu/4DzPRCM10xBnPBr6kQuo6dvc+nTlKNsvNMO54olz2lpP92zQdg0lLU
5phd+q3W2pvER4pyWblCjLHoyp8LSVkgIEfybCVsSXtV3FzYtte2tXSLsTY+StNZ
88t7VsQaWbRkRScusHPgvKmP1nel5XA7oCQqLgFhkc9+zF7fLfx9EOt2XH15sBJH
czHRy9taBX6VXK8BAtCfGQu93SSke2y7NhY64C+ulElzzEFRkpbr8wjW84msyWTj
kcRA8dKKKHnzrKCXDYdScOmeVLJiITVhQFtvyVl+XLBgP+1B+OKOZ/Q9rnKC2d5W
XV40CS2BVOHY9cxMyiZEaq7xIfNSetZcqke+PRwqh3ua1zSIVPtXhf/YcP04HYDi
MWNNdELB5AAoUtqHV16xZLSk7I1wQDpd70DuHi6IIbuMyYfsh7AE5l6s3eWrcl89
yo5wVBKjXJZnfzG38u2RtvMNOMxNwTQnXW3yk6f+mHQY0bdsPU8hNXcCeBnHnJ2P
loWzspYcirL72pNpCxICdDnm8mzGMN0yvaq6eAZvatH8Lbx6yXwCpSYdtC5JmpM9
JodfTqacoVCd0xM4LFyJeg4Jms0K7h00rXdmqlS6BjJPRuI0SXwCyj/NuXFfXRmi
d6ATSNcVIrzUfOHRhNqXRFhb4hBBq+seqMvY9GriyFP5gj0jGx/A4qEKYssjfnPh
a7AwRGAxjNihY/uHJLqg0DbIO2nNMLqDEg7T1wbFW/rtQ36nP2NNP4ZURRojc9PR
HO1xJUnaa0qXcKoHlNGwd+9BgrGQyy81/BVw5/a7Sl3t2/QWqehvdrmfIA7NLkb7
p+mRw4njEuBWC3+KWS4NKrJTF3qfljJzjLaBIz3/LIibraR8fxR/WFtxQr047erm
zalrQGiIwxbMX34DODcDXP79lajiXqyhVRAy5V9wY9fYO2+JF9Zu0EPrtOfrpw7p
dhYQUr+WQJAQ8ADUC+ViEul5dzxRkBE9qbk6FBuZdc9bSaEVWRzVeRmrHkb0R0Zu
eWw+DW43Fm/LMr1F6ohnwNPHo9zOgLkHG1CVDgI0gEKtXT1Z+Hseud2GT3jS9NpI
lCB/Goyo4jKujFmUhrRmt5WEh9lYXyHnwWFSSLPJNV2rmaZdWcvd4x1fD/3gncqL
rmb8f1yy0uUa/ud66i439/9ehOKZ03AGETWgTxdPFsBC14tDeX9oKRqWOXCJbDch
GS1YMg3syjT4JIK2wgXf76/wC6/qrO/fW8WewbzxnOEA0UBNz0oFdFr6uj+JT3//
8RX0Jrpr1cstapLFrVVRMhjZng/OWmpp8XRfjYr2Ct1x7tK/w9953+ALWueH3cox
vOw/Mvf9u32wKghluOt+E6ScsPxoiAd/IEAm3FFBC9AGFsHumw2qL7gc4mo4DG23
7HBmk/CAKv5bVu5aX9GqsQC0ZLs6HAKOqfdx1p1XFSr1r9RxIHVk3vBiDZGr40DN
SWXIEcqfgfWTDuveaQi1LbgITp90rMiZNdgJBQ81KCkOZK2we0eQ3vZREsXCRSjB
tTvPUXz0XXLGxeTwSrr+u+79KLCv8QqN31UqjrUMyCl5aNLl3uT+4+EGt+65YXh4
fCli3QGDEahwy0scjFocJftLchWoTu1Fs9FtiUFLQxVAp5xpDxiHQHCdl0PSjfku
Hu7GyyGgQ6ZeCSN31dN3h/l/upbaAmsYa6PrxJJ9O0vmJvha7lykEmDhN9jmfYys
KnsyZ5/jsRr6JanGy+uTJR/QG47EhAZXuuJN+3/66ZKskXXzGgPjC3KqEG38+8uS
kNAk5983En7X0nersqVQEM0P8u3ZwIccOzQHJM+M5aJqlg4sHXQ+ZgCOQL1csPci
zQgwRMtvK6p+sfu8jNUh5I/tfz5XyvzeXHWwocTfC4RhnLrfAoCgpOsuzbRI/hzd
eVIuVJtVuaxssUK7dOtHJvNMW+gIEWcKAJOo/zLJ/da2HbctiZtcswWtV3V3MBJl
0fdOGhShTvsbWJ187bjZ2Crk8ays4bkAG258EZCCJ1vwQ0CJzcXUQMIOsjCQPY8g
cDlMU3RT/iH1YYcCJs9HlP9hTg1J0WFJ4Ov9v1M0pIUd0pE4SAlp2OfPJJm8VA++
+cqVc2/lealv7CMibzFrI0uNQpu/J15HdosL0AXhUb9dDFoc3vpGGjc2tU9ngIMH
qAXmQCu4+a8qjMDhwThu4RhpZb3EIXcx0AehyPeoqJxpRs9elCiPHKazBAx18p8q
tPPI1ZpmtmMm2GCGLeGl11noQRR8pbQnxpq1sdKQW89wrnlGOxpaO8yZSytJgv0L
4quBSrJbfsX4VTrDAknJQio+nvVyHIG6RktaRB6IdTR1i7HqU+HMk+ePUkYg4fNr
UmXF4+BWS9zrlHh6NcR5Qq21TqqPqMma7d9woxKSAtpEIQnCjAok/qcSZCvhsjGi
oSJmBbY2047cqccgT4IcC7YV9Ke+KKXweMQ4/3ybdYx5LNK/xk+n2gabyywDy26T
vYiPzMXGitWwMFL6wm+YLUlj0qiXyBYRp1FxDxV8vDcixiDOcRTnU6poxYYw+rew
Gm0CqqgodGKD/buJpTpZSja1aHEMQif2GnrmaMtq/doJWagFMLGkcrk9k+k3aVEj
Yz7XsgZveNdeLLDDIMGew9PQTdBBW2emfxf8f0+aztHaXf7oy17pXUtIXBNCzyX1
YW4tIEtW3hEBNS7IOJmdUjbuBX9ZZJCbkH/vKoK2PNoYS4rAz1ZF2neFlqq0egzp
imACgCSSjcFIyAhEoVEOv1z1YBAeeA+pa1qJLdPcmbQAHzmtglhoLD2OFimspUQ/
h0luyZ+0rIEJJBaYrC0maF9xT5eLfGNEQZO85GMsHGw/OpRbhve8FWRd54XnL5wZ
jai3zzrYQIJRgsesZ2ZxOs4c2a31JijA0ghAJ/HVL4KMICwJhH4zfjdRu5FKeSV2
bDdOoUj2OmDUKsTaS0JkfANIpRLRLq7KRPsbKoFwVPHZVh4dDWuFpsE2EnZ6aRle
//HRryAdPcR4zQ3LzXzdLLqiJeP3Jvrqblu5GFNczMPqXRPiiPVV2VsZiyLCPHYR
7Gk2tKLvOV9OA7iXfSI+jooo/riAUv4QRNvqEdED9A12s2DGdw1RDK1zaWq2Yioc
1crRsQENuZ2eeTkE4BzVoKQGcJdtlFHLkWV6HuhqpVUlZ5bS380q8a48FPT3oe4c
CUYQCAage0iOw/BV7tz7P9zZQ5HTM1rWFkjB/iOs9WfADcXsnB9/d8hTO7G3i2GL
p/OyzTDJmJEhxmWKCFsQPrwRvugKYnQtbfqgviod8MULUqfU1k0R3bj7z0sOimzz
GQlEECIqHyRrV//8ueoq91sUBgv1RhN9mTmSKQ6FcbQmfihKBKcxKJUkceoApjZ6
ubaqNh84f7IkNdbOL8HrhnoATKtbKFvDkHmVzdnGDlI5OhLiWkPvlz94r/XGzPDk
7/K3+6Kw7uc35nE8Zjn560n1koawm6pNy8zI744aRfJqmYbmFTs8thN6hU+aAFSA
DRF693jeuX9mUhQqsSb7Z+pAs9/8TOGwlaHcH/1E4bwDkuTVYfU7aEUmCixwNS5Z
fRvLVf+kB8ZoU94p3BDHg5vlyJhBC93GDIAbXNGmwSHW1cko3Lx3ZaFEpqUIz+cP
+wj1i5WJKQZ8BvYB9CpIhg4r0SQ8cnQAQpqfeqJwCkNid/Bp9WFmpfB1ixammmhU
WDe4faEoxy5mFdmkJ/aZPa4KwdyCyTKsB9AppoDyQpq3KwvJlCZiTlOa/vM9rQ1L
XT/EAvrEV3LvGEmdhBkIvPO0SM/6jFckWtobc7FZSZQh7fDBM+cfmucZwmrtluQ2
BZsx5S8sosZrcHvfG28FF4+RsuiIAVLW1qL8E1wJxjkm5TecYMVz1KEmvQQFK4S4
EyhlLO0kkRBfcJ1KI9u59j8v6FGZCaurLezZhOVVbor3hf8O2jtFUmi5+aqn8O8o
4pW72ZazP7xPeBAs5i8352z08WLLsBLubeuVlGChGykXK7Xwc0aGRpwCCSEzMBjA
tGZnshhJa8AV4n4UIyEz30M0OW1KSDiTvBcZBo0+HzuoJZEUR5KpQXX8OFeo/yvt
h60kp0SSosW1IgckwPn5YSjZCWCmFBfW5WbgrbWEHcyWncPzHyXofF4gFrfnIWnc
im+1IycrqjQjuVoY/fj53rtarbwH2qqKkVlzVr6yAX7UknmjRp7nVacGp02C7l7v
4jrfhKNzWDWQCAtdDgkFhmYpi0aMwmQWIBfMjx2FYCKwPn+1TTLoMRd6e9/LV2V9
wW6qipakiVx/f5SAinIMn3sxTt0uND4StfzfNO0FEiKaHyvIuGsDy6no9P03g1jB
oXCtLJP5uh7tzw4vq+oI0Whlf2M+z8NE1NBTU5qVzw1//M0kU/JC4/eq7EfudQSW
Ts+YZuBmAPSszjOFfK79y7He7E1Hx2wLZe31Pbsz6QGFGOlMlu8T1NTxhmPTTBNY
tSaTC/2jl/BqCaOItL42CzsaxhLOk0cdF88FJpGa3FbnH3iJ3BWy7ZFHtrNRz1wi
/Ocd5JM+6JeHuzLFJiQy3L+wG7JfKBS4rPUEKi8JyhDlqPgYMUclI9uXTHA88FEH
owVYqabjetwgCHB8MTTf2Heaje9Q5GHatztaxum4lbxeliTPCkP1unj+ti3JnI5N
A4T4pv2VLwwi6vjuAPZdL4Sdef3oymyWZgZeHZMpUN74R5HA32minrv+IqTSLSjj
l+UsbC/X9qYEJd8Bcd+WOxm2YcDKqYj8XqLbEbUSK+bAOTYFcYIPuQ8Pm7VFpCuX
8PunxBxUYhEEBTqQZdY7HO3VAG/o5Z/zAZLvJS4pUeHXjMMlIDjYLc7V0isIqrSB
1TefHS1gmGCusSHZRNt2THI/BGb541azXX08qzXyCSFRYfVnRRJjUaZsiFCe4smD
RckwW35P3NN5tBezyLd5DwGRHYtaWb7qZS70/6Z4+zg8Da7nhLznpQTHRuMVj3EX
efCJQkB0/a8SMOQPLyt7uU+8mxHt4wZNm7t3pe0yzBUH0jEEk3I2aYsx6ckK/g/n
k0I9lLPRLDnesWepUarZ5aNUC8B/XcZ1Pxgiv2QpA0w2UfDXb7hpjQRja8KUkj9t
Evl8y2ERvn1gO9d2brDuGlyAlA+V/7Fw4Pyr5wJfE5JZKc0MYVk7K52A77HKuxkd
otg0hSaIMvp+MVgK3scrVbXPqbXlAonmtTYbLf7JnP1q2x6hdQsiLLcir4XkxAqo
q4MouNxdeVRjQS/XqCLQ0accgrjxDCR9gyKYzO46CnjIGJllHw3tirSaZpw6dYPT
jy/yqT0LWKCa2+k5TcnwEf5ziZyfQginMRp1EMheorKuvQfh0OvotwG/vAJy5c6R
+FEgU+d2meUqMiz0GOk33RwB7w16GrWpDrE6CSUCZHxtqp2EnsJS0HqUe2oSgbij
DKRe9DTZKSLACZpHKXPQscOQqm2p80crDoaiKLkOjUf5hvmYYHQ+LpC5cvcYsECc
2Xa6+Tn5PMK+LGE/AbwrUrnksTCPg5tfLkgndu6YO4T0kilHxecfXrnD88w5J0ps
0NW1RN5Ln+K/NVQQGd9IWbQm8EGVom6toGcAiPFZxy+vymmln5joI3jv77XisYMK
2pQhewff/x43qAijZNgpZh+bdxayu2lKQyuKHv/kdsTomS/1P4ZlhxHVdn68M68L
JDry5Au8ScozhL7cT2C7hZtkEE+DZt0hTluazXdrMHRzMdJkKKeFX/gps68qRvv4
S2SjrodQv7br/dkV8SV8jHxSNzrS+Cyrgd9Wud70rVM9Ij6KAM26TjIAM8dF/9J/
Uw9CNYK6I/K0HoVdo1rDteQJIwfIYr6o1VbKYdgvnceFZ16QO2mGPIr7zVCg2kuC
uNFNkHy+3Ncen1RuO13PAn5YIikJFcgz5UGwVJRjiUllhOoL7o6FHfbq0tE56mCy
Ccwa0W4OOM8v5UkGd2fcqmD5CfSFaBKWmI/8XpU496Eoe3HSv2h2wDchQrd+H4WC
rHPRc1AsH0g91mSSO79vC0dFynTyaRPiGkDFyziudWfgibvmHDa/omtU/P2+8wpQ
Rp0im1Ckpl2yhFBcz7tiBj3PVb20kh6miL0t+HeCa1zubQdgugGEliiTUCLupVZ3
c6OhRr2MjlQ5tftR51VFo2iYMI+60pyr1lYLxC+5s/Os5SfAh/NNz44WiQQJaYNr
Ca1x7Y5HskiXdL1VBrtVq9o0owjZAR1/MhGz/9Qv+GCGFx7MMqCRuX38kS4RPxj5
SZJ8uOvEI8o0qH4ZJ+GiAG/eSBum5JH8hGpWfPUHa5ou3AGMXMAh7PRhIMcV1l9G
KVNJFws26f9oVETRu/P8YN3I+a3Fqpkp2af/nD0rTRu0r4zYivBTqbfUpz5NaaAW
mfSdIha3xPBiyzlIoQbKz4WRtArp6AsogToGgmdcfBCXU9MbUZQZpqzPbj517wEL
F1A6F4iLwOHW8zDcLRt58TZ8GzBpfnGlWbfe0rdpAew19Q2pi0bcZJHweZg+ZEeW
4acC3RZrTSEC5/HZe7vYa8NG6QaFnKcK6Mam+JVE2VyArd7TJ3QPlpUVQ4j56Zb8
gr6ZCEjRhreVXmPgR1Yv1h+MLTUAIy0fvmwN0LKDvbU+AGCEjb2bgOCEdk+Ody3O
XTmNdN6DblQAAw5jU5aveSPyFSmtdZ3rKLRrex5sy+pqnrk1Cbe3x+yDRKCo77vo
03ZQ3y8hNTYGexnRjDLwGGhKdafq9e610Is5a2iM4IGvAt+6HuT1c1RjAHFRFjDu
epD1lvzrNoecgZhd4OaWsIEeSPWUMlMdCtrQfJl7h3+SNr/qW0mFv8LA7NHMEOOc
8HFZtOmRS8NjQRXmXuqKGY40qZ359JX4cXXg/BfKW5fNok4hkZvJ0EK4TA6KKWCY
U1YENjJRpjvjeo3cWalZggCK1MvpepGlSU7wHI6zzij2CoH0FRkZeZ3WRCiizXNx
BOONFdmawdnRJwT1Cr9RZ4SS5xGBQvTtHeu4rd9Eid2r9dlkgGJmNXMS9ReLgS4K
kUv6/U7u+0sztGgkuIxO3A0XSy4EdSSnbBFlhWUS5mCGyH70rZgmxOhamB5zeE1T
Uq5dHktbBni3yyWOVBdFOIO1dgxPOK/P9ORZ7uRVPbNR/H8sUmE3nLNC1kqd/5/o
ymtA+9h9coGHvsZ8ztaE8/bQBYQSlKclOnmhjF3yg/LMAmg4fTkDn/ESMVSByndu
Rkig2bDlIBc46w4sDsgYYXxS8lS6nNQNvsjBA9AUjR0Qu5osZqhoVmYeJApgbUW8
rG2hYEZNQJDRzviqS+DhTBjwsMmnYOHo57qICb7K7uylj0O0hmisFI/hzeH5YhH0
0Bc1ADSGcpinKJ33QZFxVayWQqr5sb317QL2eoYyB8tCTtToS8yAMvcgga9Gzv9h
BaBk6espP9CfnCjqXRLKtQRat8LCijnWUr/mcNBPGjI9s4MdzjBIUthJvFf7qv88
nXU9zy7VUKJn1hwLyUzsfKs+gdZZvAwfF435w6vHsELpxSqnooXrdxb/WledsWtf
aLHt6/PrJQOubiZ98dF9vALK76Vc/oyz+ma4KvnnZLk/CrGGPB6o/TL9+0DAPtlz
bimTunbPK4GnXjQ3CJ1Q9CwW693+QGMBkiHgVn2xjoi9GfGpZdhJVMUKqcA3vlVm
p018YGUm07qSv4nP0s22CZ/R5tzlcq5/wOIXttMSsXYMUV3d63AcV778uA0kJC5Y
XlsnM6uHAR4VPOYr7ADOzATQVNpSLrg0AfEKguzFxqEMx/2/HzZ2eSBbU3pePVsO
sdiP07imPxnh/eVXmwpS6naPjH+UhbNv6whoNnIsc4f4wzShOPeeU/70vaH6x/g6
3s+vZK7S0QDc4qqemzfbKWVkuHW9qNr119/f+IlTLYboZH8/XGfuODOZ0VL7iZ32
FhdOd3zTGCBVeQrPofv0R6DvECyrXMqJulWq5ItPfmbL/s6RCJSArigEOHRGTqIQ
g+MElElYtXHdyejpy+K6fTMpznZ6WG112VVRRvqKXTfhhjNrdqHZx3Ykoi0W8PT5
7rMtDP/aPHmCezP4Z/J66Der+tfer7y2kgncrcup8+MvdzHfY1bo3L8MtVAlx2yc
kO4wMuh/CNjdxYlOoLTCDawMSvK3h7c7QEu+Mh5/HUO/zZph483rQpRxb2o/RDdi
ujHkwSodjphOp/8H1ejzQtqFVrk6ehGC+9G6BdpqWS8Ohoj/s6SxVqnpzeaQ9k7c
CNroYy3s/jtjEEu8VJMRhfYxeiMB2oYso8hAzwMlg3Cc5EAHX2NZlMNnBJif2+ld
GO2sL+848MNIeFichlxlDZESMUkPSX7a1DeZFnjaaG4vQzaiwzrKWyk8Hy/T2xzo
xcHCapvKzU+R8KCOSDVtsdRLqYPa32yC+G2e9Fke7Iste2SQIajFW/5lHMdqurOv
TGBHsdXYRb/aVWuEEUs6O8Obn4joD+u5GRygQV78mBr4msl+j3zBdflTp33al03L
vL5c18dipbiuKmhr7KNSHVNuL3KvH+aDn1jEjOwx7DTl342+4xj1RGCoRzuE7RQj
PTjtCfkgkcBic57D8mKX13O2IqgG2swQnp96O8mS2nH+hQM1YO00bVhe4q1w4fpi
LH04QwILYn14CqiWAvWEXxkiAIhnsBB3IuwjuSq1EtxARPdV4dh1P153ueMtLJQ3
eFY5NbpKzEVcLDQUTWgNCFIhRwargZXxBaV6mDK8AjiDCO4NOKwId/dTZ5pII2JG
YNCzlkWW6Aea/ESpaM/BxOfIZK2ksv/8KHV4ZGkw/LLA232VjJKfTgP255bnbY0s
nxHGs3hVxJ3ht1wKA3OcQ0YXolQPnD94VN5apL0zRLbTbuf7+uBxYr/fpJNlxxVl
MJnFfl3MZWyRX0IpD/EQnGgmpdejwXjWyVDMpD75XfnLJG0jEquPFCZhsY4QDJJX
oB5NnxuWe4iMfVQaihId+/868coP27p/SziblXoFQ/m4wYyO5We8pxv6mwRiSCvU
6RDbraUpmzTCCgtM9oAIu79/bjfmuO9Y0N7nHmnjf2on257++pIUzMBq9h3fnRsz
nLnp26pRnxqoyro/b70//XoAM1F7//SGr/z2n8JDjFRTQXemw9B45wNfQWQm18EJ
atV8yjrB/X49BxAhWrsIfLRJKoaxw8/McVoiKxF+NXMrRKTUXW8smcYegZdWvjtS
2XdO/6rzmyfOA8uBvT7ehw7PESZ8WF5cafWBsKyIWpjlYSsOGYXcc2GLqJCX85Iy
z+5WOHxY227+/0xbJ//EE41pu1rUqX+cj7ywNLu8umbE3wQ+y3V/Ol3xrTBdTKaQ
SkCNT/cQW79g1PbmxZeolJG+8ZpfhYWjxUQ8fvXkv53GN6WtPBTtk3/35Ar3XSvq
u2CGhT+c6PoiPh5Atfw8OrqbAApiPlWoL1m7c8Qj80mz54YI/TWBLIJ+SB/m9z6L
FHmItWnYw7sRVJMdXQjtcPjh8ZI1bzgY8Dp9O7CZCXGLcl+ZbHDcjfEJH3D9bAGl
HRV6sozjC05DhF5muk5XKk1xb9cSRp6uUi6dEj9jEcuJEomFEoVIblvx5gYhWMOL
36fPJF7NPR/Ei94SePYn+pBPw+5UmahOtDIYVrzNQYNWHjuQXC3YAVq0BejPG3xE
F2OBqNFufDNR1aYIEKzMMrqaFRYwd/NMk3QsY4LLAneDW4hxYT1WP0RinZWF52aO
VxYaXNPXYsj0i9AVQl57UYZ3KxQVI14vwy2h+TbmEn5+6WjOwBUqyq2y5B4Nuvro
XNQ67ErArWHwNthq4WldfPuywzEcM5QwXsQmxEMWJugNR9HQQaY0S4FzrperKvBu
cBkFO1H3izHT2iCuUvxd+uecfuDIfnvY/07E4LHxIkKblbmgDPF9Yz8Ay/PBj5+t
4otfI9JPm5nUMN9BCYz6JINYOrx2ozzgA4HcvN3BjK4F3CH4Jv/Z+RaaHEzPDCWc
heK4tfiiJlFIftjgYO4XwThVFgcHMJ8kFMo9/NdfHpe7IQygmDHDamSw/yZB2ipJ
j9o9vdLimKdKnHMMI7pFzph2vYjbD5EB055v6CKTNhIbBKvfsTndzuAvM/DvZhgF
UwY6ElZB09LrrTYpMXJ7v4l8yIx7tGgBwPjvBTZRYrEQgaZrvhhb62br+klL8fUx
kEBm/I37wIITb4Pmccmf8YvP8mENfMZH5UbfSjxdachuI//t7Fqs8EeP0dLooROy
qVYOPOque0ZmA0UkBocFakr3DCoaw9XqC3cyru4rPMoXPANY/zW5Wui0nd5HcSyR
AhCG6b1HLIe0ZNnZE1ekzjbPwUZJzfxNfUgX8x3nVtjuGCC0Rm1TMwcDqcQ5LB2I
7PRinf/dFVU2zV6kq+Jnip42gFABQV+xTaZcsLN7WSbN7+OUGAYyk1FGXWSZ9ymh
xI6IF2LiDUWojNZhicirGl6o7TRHnjGCrVdCsxEWKvDZa5k1z0415QGd4AW+NpFj
G9NdYJMCjSspHXjHariftSMSSbtHF/0uUruc0hC3HwhOimt4j7wbLnYUPiujq3gC
qPLmX8bbwtd0qH5/Ub+5nnZIGnw628DweSAQ/noChiy6ZXXjEccmje8Kh6ZuA1+2
mmVAHT3yIrBK+dZZCZX2nWjxp3Sgwwnu3n3W3dylpt1gtJwOzi6A29Fo8mw3Id2Z
xhdlxdByGgHejF3S7oj+f++jq/Ze5vB+L6gDbuvURqJs4OnsdO+ngxekmxryHsJl
KxSdyStHYK4dR4/8F941wCKLI2MB0mpIllF5ryQTdb1hxnWvyyFGFk+LyrbiJXF3
mwMUQBiEp8Lua3/HFB9MlUV7VgCd1diJPkoOtLDPx7WTUyIU1LssZgbN8q0/JhyO
GwO/kYCuOySKDGxPRi6QhksdClgxzrp8f3bIUdn7VULtMi8UBxlvA7ADxzoNsm1W
gNLmb8KrvvEq/Ck+YpaOfAmWcuMWOTchH3eptfjGkjvTU+qNPNMfR5quEu0rKVRy
ZQKq3FtAcJ42p9XXMVuFxNAs8vr74cMwG/obZ1OlUW7qOdpbQBsFEbbw5v6LhrR8
MxVHsZiS7G1V+KUgoCaJk5/2km6rGpuMiMsTFGXCLtD+058niyRhV5K5NWTKN9w0
32z+8AJZxecCnHXpeEA7G+q0WOsDWyiZq4ZcxlNRqFTMeDgo/VJd07zYTUdkX+Pk
1OHRWnLgPhH6qTZG8FJ6krDhXpv/qANPekN5l7ydGIwtf+2901q9njt+sk10wdvF
zGVT/LB/vVLFZEbBwaF3DwWnM6gLG9Ux5v3jNXOwwLTkRlVJt5vfM6v1tXE2ZISv
0Z8y9K2EiAn1qD/E0IGK6IeUQTwd2g5ZrexLcCZxcTEZCZODd9XMHlq/8T4nxT3L
WB5xVS8/zFstm25N5WWIi1p+tnHBlgFwIx94MB6CbpU5LexlGJ4N1FBg3Y/vFDs8
yU5OqO8rgSL8YEyNCh89COxXweVcz2rYcVzLp0z1xDeOswPybE8w705ORWera3i+
hWSpn1j6nzVf1aWBmjGQiuWlmO7DeYA3Mki8IDYY/RpN6Twa6tHfQ2WOhryxV9Yd
naFMED0aooGgyMXm9+6ZBp3TU9AFORnrjGluS5fU5RahZK+3rlBIXJ7simpb2Bmv
wIfjvMKZS+hELaUcXo7fdgwHYsS3ZTex0jPo6xbRIceRuP4GG/vwHWg6uS6ZchgK
fzviCPMbARiXteBOUyaRRIzaPV6miJQjIAk3cCeS5c7W4bRmjTJkKPn5oNQjLv9M
sBgJ8GYbVrPXTiV/PI0SAzJVf84XXMHMovINoa1jIOeOVORlUNQjKI7k/+jpzozm
KRJt2YmUYScxKWC1/gah2rZ8yZK8bwcKSEGV9Ay+spZYiEDvioQSCBrAQSBlurqQ
bJ/pV45cZgC3uuZiuQYPav4Z6Ehe6naQ/fIK8ESbk+ZGZkny7EHl1gB/RZV6r0H8
zPeqCaHba4aFYXymGxYhlBlv/iQxD+OdJ+vQLLwbwNaP4saFruZgnWy6KFPOfxPj
5NFkAyPmpMQMZtACI8Vn/D5T8muZiu65xqcHiEf2h3Uj64F0WF46rE5uM3BPdb3X
EbVJ66s/FEjwEc9UXOdzFQbddSf6tbDpuS4s8vvFfe1bAfmUptDOTrnGMF9kE88x
YG1GWbwH86X7Z4bwbWP0D56ZIVMVRNeJlzUxSbnysoh/7aC9pwogze4fa/3WGebG
NTb2JUFBUnsygsfH47YiOOdlrN0xkUtvRRytrvzEJy3zGUSXgY3mHmnPEGbIdMzR
wIYCWtuOVlKOrodYfo9XooQx/TWj8IO7xZFd7vAyT25RayQe+19CSgSPExWLeE3K
kyTvC133sXL86Hx/Fz9xlp4dkhMA233TJ4QGPv41k2jo8Z/5WWklD5+CgBxVD/a+
6MIIzR8l3OG9v/n9SDoU7mqqWposcuQCrYjHqq76hn+etSn9LJbD/Zz6QK4UtNOz
Z9PhwfVs5CjqE0kYLV+a/tPCRHigF7jp75ay++0Ea8szxPZwOzIT2cSqwIkTeGPi
X4Ag9sn4p7bcLdS4OGZbTLNTvBbKAJR4IhkgAaLyHj3LSdFP+tSWBMbXjfyRSuig
TS9Mda64ySdeE9yOZxW8LRdSO1K/+vVrZt/2dxkOaERrUpkuHzPafBzO0tff5FBI
pl9kvrLyoAvK7ETYXkcZyhJo+ND9yBpsbtyG21fnlHjd/kmjSoVfBKmN/ouX3g6B
MPd5keMa5YQXTO+cabmXWBFtZDXvb7C44fuwqndFrHk=
`protect END_PROTECTED
