`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IhPx8uKBJcylwVEipzzEh4gauasnrih1E4nD/v2P/rbiW6WTf2691REqAsWMdoIH
r/4GWzlRLcHP3jQmZp1FxBatrlEf6YMPDej+qv2j3ujBqT4n698zfOssCJnRe+sG
aHeOdqGLwyrCIGJDoyy98Jn9s9X/7qXtzwFmIorXoVr8ZHNOwyBU29HXUB1mGRfX
PR+h0GYw9hPFcH5An2B9Nz856G7GIoDOE/RYGqYQ+coXF1govbYWrUTxrpd/5Hnv
z5XbIIakDT8bhAHvx7+qsNSXjzxROaM9vIvD8q1qfjHZD7aX558iO53hMAvrqqu8
r32ylrpeLjw16uCTbZLAAwJyrgszd+FyTRCe30nQb4C05r+T4ykT0MVIEjvjXVZT
kCJQYq0c7j+cSPh1J3n+iRv7QeLJmJGKAVehZhN7o6NjAmHQ7nlEIMXicWd6z7C1
dxQ8vFgAuan35LlKgU+Ijyi905NtctDhRC/jIbHm6vn3h3AdEgZgecv4nZcP05+q
eI9wCras8F2Tx1S5b4A5JuvpnJ349gUUUla/zkvQ1lec+IHoO41n6rYy5f6urivG
vxjWIqC9Pv7rt/+OWHnIbMqC1nKh6dAtfmBAAA49RNHZOQmDRXJdgmCas3lINW1S
5dQ2/LClhLdjgHz/XRvX/XQWCYCmIIYZqqJDSl2OvwNzPw6SScelqSihWZwvCJ0z
nzyh2QukDokDTGP/X4IHxeSm7iuTbvgVp+xG/sCvqZxD8Js3RuVJHdIdrO5gXjyA
5E4Iy3j8SDi2YVOuMSLJU6u2WsKmUFEbu7/PPy0dIowTOJKpcGcvhs9PPneQgJUv
0oN4W3gatXCaXB5ifVA6WKlGt0qGtzJxiMBQy5jbIljEDhswb3kgqxlDZwHQ938U
C/oJLlfi2+T6lgIRtRLgoJQ0v6MYbT1uvaVk+A6bdNYl3akbaZKbUbknlzMBeBPA
7rHVstc2mHt4xBmRTb4oqJdi2pcmekdbhvjfFlQSPA4MW6KB7oNoWuM0ch7sNDqs
ShFbaXOqOqslb8ualFa+pnuWuHyfSIUhHb7AoQ/RxiIAapxKQZMyLJXm1WEWM8tT
Ru3TZUO9E7dGHm/U8MNz86dUnoPuLZ1JjAGjY2+gCBlgFrOi+zPEK2fx++cTHzG7
KBZ4Jb9Hj18OVzelbE6xPjnbPGADXMJPQWSuNJNqKRH00lTW/al8syZbK83PQlS1
vHcH6tAaYYpHwramwW3ttH78cFu+beaFeUiVc3LZgJOQ0elrB/ntCDE1NIpOXkdy
dI11QypnQTguelHkjgM2/7DeRxBiCA3g7tIxbF07+BxSPYWw3gUS4NGOKWdQN0O7
iNfxCU1FDh3dx48DV8LymmiGhng0YlYhlXvo9NZ6OzBxuVpK6h6L4lh8OAEkh6sH
QxhFdugvtbsywX7HplDvcferSvi2KXQrQvjW0AGubEYRiZdgdjmNo+iI2U8bUIi1
fwAnnOjc+T6WaTkr0sCpRbXOypQEeHvKS6l1iGSmQ7XOGOXAHjBOA+utlClhpaIN
mxDI9zKenVFiXsPDQvpbb8FTtLsVkBzXmsxohaFYOV08+QUvGeEDgWkBCGAh9UA2
MoMh41fuxVgCKwyMLSoLWPfpJvq+XYi6mztIHV/33nuTUiMMADu9XbaW+5Kr1qao
KiPZpcfvQ1ACfdIdzTlN59hGUjuUxs4H+GENTaVywyJm/FfRzxhCUR9KPL+8eY06
sf5EfsjyUEWlvKdjrrOt8fUbZE2Xn5+EFNr5j8fByKuKvKC4epIaV3vWrTbwlZJ4
FdoM+wsBct7/pemmp1l/5IYVju2KB9s7+KkLPa9PQ2fvcWz+ErNs3Gw2WWRfAWD0
dlVLPewdZf1229DPISErnkB7oUhHzH1OFiArdeJzRvRleKURLt39xdliylaHWa4m
5N1yFyi3uGosXNu6H2uzebABMuLST76elmnOawGrCHe+byAuarhlZc9YQjvQi+Zd
aWgSa9Pwt4NZp9pUPyNoxiFf5tufrCRGo/ghqiAYXizNcPyD2jZms9gIaSCZhrD3
HaiyiTujQyB2vG93ylVnebgnQgQQIV5TDktvZDsjuA35V7E1lngub2mIQLSKmj6n
+RTest15m1ufSJFPVyy4V3RWCCNMx7DIeD0eRPGLmiglCTVUu9PTa/WTRYVyWyZQ
lylh24IzDrGEnfiMF8xKNIxAhEM1gVTYoSFL2vTm5KGyx0gSs+F7sbIURdlCZRaM
`protect END_PROTECTED
