`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gBk7qxbkqXmL0DA0FyH3cp+US3XCK3fvYlSuVfyUIhG2oGVkxsFiqWZ87xTaYngD
tub1ZkX7W/9cANRN1HoOjnVtQA/MxRpWlhmlTAeIcwfwW399ZZSfn+rgKlsc6YK0
dNAjjcA2kMwA9dtW2TAnV2+RReFhqFZk1xb/rtJETyaQGDBe4v4mlYnOaXVRe+Mx
F/4Tl/5lxBrL1fehdnJox1CoEiWlzQQYJ3ftVEse1uHYoOO4Qtp/GEaXOQPHmzkl
SoLQJ60JxwUlCy/Gf37s89FeKZBqE1waRDg+D3dn3dOfX0c9rgUMC0pl3HSfJKoY
WdtSRmvOGtwCjNdeMBwf8bNx+IXsu8Zo/hDHidNsWH/c/m4wTFuZA/vp8Ye7lt+3
BakfKg+w2TbEv5Y31165FviCmX6z7Py6Nb3sJDFHJlX1Mwb5eUJlp/7ZTPTwSVaI
iNfi0970yvkBTeSfabC090b8t1B5r+pgqy9umRmhzaJAqfYk+9EgZ0mGW/hIj6Kb
pauMyy3eShr+1tGw1cLzYSq7PyWhc0EbP3EWnqw5Hx2LAf+q+NvuSZwRZkOoKVAL
8rBlk7B/1e09/jfGrp1oUedYOCJ5rgyICwF4mjorcyhWDco++hDTNQPmbolfZGJf
1FDINeGA5eLx/gi7G9OnMBpYmD3E7TEyMvGIGbo2CSda/4etjDOgyhJi11T1ThlN
MUdjX7PORv5cUEEchYWg1HwkI8w6xq/rVPH04WXpv928r37XgNBufk2N+LS5e+5x
14ScRqcTo7Lt7YLw4j1nz5qy0T3ZDKBWD+7V+6je0U6vFkul1ff6ur4GioStUiUL
Bq7Qw0K529efAL5dm8TgdHq0xMK7v5mSxG/3uQaO9xaJ/Rh+M2NCm4YT06YxN/L8
L89uRmPqY6wVjn0/hmbP1qfsayXOE756HyHTypaqqKZcvLEYpdOtwGAYqDVdTuao
GmD9FxW7tnzCXRTiTCjPyox/oJX8IAfXDRsQ42A9SGVFXgdYdXGAvAM6L/LY0gm+
lQXca8829Vi41mjaI8V5jECaYg/oTRZ1a8bb8X14G3kvCN37vlatH79dxBAirL21
cQh3CohlwRjHtJ2VcQfliuDEykt9oCfF4f9ok+2IqM0TgNAzPi6afOEYm4cs/CDT
`protect END_PROTECTED
