`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y/aHS+6drNAqyilJ/oPev2lwoM8wflgCYrohu5xuyf9vyXHrHb/boxKiqfmZHfDJ
wOGxhbs/ISPAXODsUgw4jo3PKzSCTae2hluItEZ/IW2SksreFtTrk5i9H5di0pTe
lscZaHGKXG2cFz0fDj44XuLWQ6QeFxtQ1Lh5mQutDaDuHWIA5A6EqE8L9+tuQxDy
J5uO87z8us26dySMPxz5T6qpRwOHHdeDPaco9yQ4yfMSBMBoBvkiluk6q4AghCvB
f2MWb+vrTkpUStz5S4NEGOajobwOrQV+ryX1WCoXzNM0YtHZa57aAw9DNBuwjoWs
JS4wMvRdDYL9+Z75DJjBubi/Zlopwi+AzAQ8oLNypkuYdHTEFSs1yLHhRD0WLbow
/EGlKJ6UPfv2fgeBcrHn5pCdHSJszTdNpFbqVDoMyV7Pz8R5gib1sgbMVt5/vPbc
OEfUtjZcNCdzZ6rNULpzanf1JG8U0kflRQmulgQZoIh5yWEXPNtXSCZgwjNf/3Eu
C5Yh/d7H7G4CFcqi3ntii97LmOcL3MpEjUmJTMNUYmWlYqXNGayGcJfxoAP6X4iM
0hrcxxQ1M/bFke0UhTuHgg==
`protect END_PROTECTED
