`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RD14UH4OTMNaAWgpHqwirIZ7pSIGnAoBrT5OH2EPNOmsSdzPXTgT95A/a9Ta1/ei
mfd/b6cQpshfrhbXElrtNpAxHu10MYC1QwqAb4q2KRN5imCE45bJxR5dDxnxS23y
nMU/RdtEfBvYu/qdOvLtTez8o6ZIX1AKmTO405BcH25MHuLqo8mXQGCITbkIhcNW
q8qgHgX9SL+VZZJs6OV2srYWJFBteyiSiwBM2RlDyVzx8cVsHqhaqZPHb/nvO/xx
dv0nwxSLyOjWCQz7kb/eGIg8nBAKqPJYbSnTZOBDaFRxTKlUy8wkyN9mIcF1ZFPY
Weko4KA0fdr6JXYEk1XoOWXQ22VuMDyn5ksuSjeQkt7X+PQm/l/hpI2ODfpYHAQ1
Qb76lbnKTn8OrXprH+Kj5n5RRrpQ6NfVOrj28LfVjapqArLHWugGzvcskJehxhIn
zQN7KQNV971iztRpwNC+BX2L6oq1VkeIz2qNHD7bUJi6oomxV+g/g1Xt2HCIK03Y
BOq/6AggYg5jCHOEqnsgmQ23uL/23+roeqVo69izfklx2W+zzHTaHHg6jN8CQLgJ
TpZ51KDeZTu/or2ew7LF8tI+hT4ZYqpOpyBmlvP1rD0HfqbAUjP1Pat4ONZaohmY
kiefc55HwxTOGhrCTHACsWiJemikp5TXuDMdnaO//YEnwWhwvKY4X3ce12K9+nER
K3fGXO/4hIbho9KOF0OJ9LqYj2B06gmQYOHrPOU2kT/QUTImTFlvOAnX03Q7gSuf
J2tISdh5HYRQmP6wyR5mxzy9bLEevluqiF+Xr8phPYvJ4PRBjq8DUFonlGFWR/U5
cHJ7UB2V+km1BjyuPe1aynfnPikBV5+BC5dtmAkDfMLNCMdvZ6fEWcOiVxlJ3j9c
wmmWGxrn5Z0p1U1Rb4LGKS4UjNqTt8lJuLYpzUgsHyQREKmRcvK+zli8mF/YLwd6
k6Z2awPa8pF33SrQi9m4tIoGT3sWeC+3v/FGOzIQVgE3QECHcNw0goxSD30F34xC
evYDTl+Ip1fFte2mNL7dyjMiN1/UWHclmzwzT3AlhGgI9xw1M3VUvSDK1T+oDd4k
i1gIrHwqWEs9n0DcITmMaZCW/NpXNN3EsZPp0AQFm6Lzij1MKM/ABOa0XnhgVMRI
GV8K6+d8IMzatnUtET8qxtW1c91m/HUls6wdHBvHhwgOQOCnATYBPy44akuMUtMi
VLmUszHXthAnN+2RPvbm5LGiDqiipNaMW/GDes4XwkQeqn1N4ziyuXG09FirDbVu
S5HpxHwWNZ7ctV+FfKVSvIf/CssDNWdS6DiEZjiyfEeK1WyvCmBaEX0Hx19rfEiL
/mxdumZiSZKT83z3bGA3E7d+0ZqGCAemV+2sCNPsdU5zcnYNPmggsFSt9/iFQpxD
4MAmDq9+SMm5Jisb4rgL7plOLErbmksK0G6Hlot8hlz9zYLC2OVXVsRv4YJuSrKh
NN9HK9N12jqdQa0BCeEjayqlqbcLYMiOwgWVgxFlL/B6rjwJXYjzLP83dwIJXcXt
5d3lmT9EsaqijxWQmul4jhiiU7VULd1p/R4wNBk1Z/CEU086GwJVWhnLh/Q4iTj0
KR0s8Dzc9GAtzXb0JrdqXCPX1IoiBqnUCEyuDji9KzyseU0Zgrubjo1Hg14l6p6n
F17JAAtRKvkmXg88xnsCgmd6vwxvh+Q+jUANZl72jDUTS+SWK6/2QybsSl0vJtE2
G2NBdTV2q4ogZmlANj1ImaHn7uSxBFgiqbI6hAeOJl+yJa8CaBCEdIHA0AQeV8vk
c+Mj0wXHSmcHu/za7nBDF14nIU0aivqQMblRBApb2DH3t0mG/zrCIz/y2HOCpLld
44kFiGu+9XTb9Cz7Ra+b6PUzkSZ9eL63TAtpDIYBGgafdvRFnTUIbrys3VKwMMMO
dPdtBLbQ2LEjmksjtqZLrQ==
`protect END_PROTECTED
