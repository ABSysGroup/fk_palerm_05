`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NkCC8OPUTGOn1MU42M/W0/xiDwfRgK0v3d/DFQo6kwCGoQIj6PH4x/MgTVm/4gj7
dDmDURAeI9vqc/IuSc5jm7TshygDKiTyDcSsequQKhUyGwMQDiB150BdSp/OqBZq
aa7dVUNs1h4E7+7aSHh1zoRCqbgoiaZkdKMfXtEqE7+es80rJzehnC5JNoiamoYF
4y5pu+zRF92sOdIAYcHAkZtJUEHJ00JXBiAa6vxsETrgyBwZN1GqT05IASEK5CSc
HlrbAyZTO6dp8pijHacwblXq/8czxC6VA0ZFsKCYkbIEVwkMxL8j13GZuXrnYme6
nK+ZI4a8XjM/05Ezan76E1FRZELU+oPYuzRCjZ1O21XcQtfacHuGX351fi9gpECw
HMtEB8Md4tg6wWcgnZJjARAYBPcs9rQSS++av7Ph6sQoBZmx/wQjOIkcP4jLVxeL
V7vsS1fYxitl19vsKglJ/Q==
`protect END_PROTECTED
