`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U7S15ohX6FWIade+JwJOsT8ApICt8KLJ+4osIvwcF8DRdKqDbsd/8fxjW3qmBchT
qDcnvULqYIq+O+bpDil5j0UE0jGSXk9Z2ktumziUalJ6025sc1LnRRxArcV77A2e
zQo23z+ZM8lGa2AJbh4jKDrusKchhqo6Id3Jd3J9GFRyig2Av1NvCb4Qy99W8LLf
zeDQ2oWbKuUtR209/LTQ1q3a/TCvKsMIEprJX9Xo2OVvZ6P0jP4DdGQ0YJYIfmmH
Tm8Ss0dO1x/rGvDOHs37ORTWjbqmNRsxLPAHFhUBtcCzSbhUWa4gEvREi7geLPw8
t3OKjfxzi79p5fYsCtxlffvE+37c57+8TOxgM2zXNvCy8Uk7dvUL3GG4UcdYeBfa
ypd5j0B9whFgv0ys/jnYyRNCYau9EEBcWp5hltdpcYSlDSO9EHPwoV/tHo2G7SLO
KJDzljCwsaQCChPUz9GZqEQQWwKeJsJ0vjeGZumGoRUcOFsa68LKO27Gha4TW68g
H1KEK2+B92BIIyYgobDcKJwlgZEcjErqaFYLe42h4N1g9asmzb6/Io+U7jJoWVKM
hLi3KBVoGHPMbmd4d6jeBQWs/WlMgAVN6AZr78mG+owmpW5jwXu5Rx4+uL5aW34R
mWa42kWFAp4r4/VBmk9GkKcB3Seq5LK2qF5SnRTjpW4=
`protect END_PROTECTED
