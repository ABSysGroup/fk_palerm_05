`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZVcRzw+fRFC+gc5G5/H3cfepd/uvj6ngv01QbQxRTGAjyaJHjRWkqrYtt2KycX+C
W5cV8rNWpwW4x+w6cRNPk3RXw2KDDUjUM46yanA740g8+cVLSGbUd2VKKRnMEl1j
gEDqrcjwdMhzwJx655wfi2z3Q1gRifedLM9/HkMnTFS56CujMk50aBaKLDsVuoYy
EokEhmrRF4xM/BxuIGr2DrrgvQh5pt5QYRYN2+POLqrVdLmH7uJo/oMfw1SEvgBj
aTQ36HcPZuZfRkEqhNflVJ/TD8vk4PHhBlsSmusQCsm2DwWkSKrE5tDFP+BHCvJv
xfcsSUuGY726drIpd53kSX5JVmrrrSSDkgFwx0ROeXkYWt9qjSNOqBfzHcdXof7C
qBZdzNBuiBlQijl9XAfkYMXFMyQdoakOIj69xcvHTEwFGiH0J+TB8E4Q4ViC6dxg
+fN2lGmy7sYTxSN3iT57RSZlsFzBJEH5nMbQ0wUb1AfYV4TGHnr4FkVgZo8oxiZN
rwMDU/t0b0sHpmj/iBTghrlDKCOrmbezHZTmTccRtmqbRveTmZOLFbjoS5gWU9N8
`protect END_PROTECTED
