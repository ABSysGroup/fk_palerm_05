`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nZEHVf8N5Iwlccbef+KLbyNRBL5j0JbENJxLP4NSF4P9tLj6ytfLCHugWUFrc7bI
zDR/a9Mft5e5QAXdOg06GHVDtMDLPmI8zxTLOooFDCdryHqq80+GQ9rOloTD0FUB
ImNHlkWqvk8F6MP9Q2CaUCNZY8dHjVC2aIky/ZHHUKq4knwh3gzz7aCbIAVv0RTP
lIsphQAd7K/s8kVoBsiDI+6GjuFmaaNNrltObhneM2XiMY+wGmUZlMobyoJfKjz2
bbIATnx/cB23YlcFhg98+KYu/d9lOH5iFRvc5DilOFD/9kdeSNEy73Qn5e+5MR8/
JvnGHQoPe6SHNR11vBgky84//w0OGZcMCqMTaU4EagJaDuCW3zzGZKN9RiI9gy8V
3szLqJzDB2n+yHDAOjQ0To2UoGeFfMvKr7M2bsLh6uhzSvzLxsX5d4NMFkaLoHGN
yxbMzdYYb1xRqt01xkhKOP9adS8YAPv/kqmuHlspjPcEwV3968SgEXsWedCaIKW7
RHZuZ2ZSk1b2GB1XznM2CJTfgH3fvR/Zg/1TQi3b9bkpG4XS/8aCvJLCQmYAMyIx
UY3XRJAlKafDkh0TZQQOZk1Tx/9wviOUhFIpxSbFq0RVkSsq9yOnLjvlAUJm6kBK
Bc6pPJd0MDjmAVNSirBleJFTbFHIoGe4KRN4h5dhtVG0+yiq/rRnxx5fs+7MJYdT
ldyRVrgl9/Fjq+ZN9LKXOETBLJpaywGgb8NEoqfZMx4=
`protect END_PROTECTED
