`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ylP00UmxeHh119iYQKJvwo885uDyD/T+5wvGqBxj4BE/kO/tb5Rz/tNlfAsLl33g
bRJExZTnJN28nFtiOYqujCDOiEu9dDegIArLKyA2iY85hLNSaVxEMteMH2EJBybp
Q4EIkgDVmH+W2VKvnrdBU7/kSROkB3Lp9O7TsaDeMBQ/t0AO6cul08bMAkpJbafL
wnlAPOEaSt+haUpVzLDWbBnEGRozc2axyKjRQVbra7iJF/a7aDAf08jb92T6pVad
vqZzMJRQ/KpnG0/b3RgrYi2NT8S98n1GdL/4mI4O/wC2+6B5LdJP5jicrVyAVJeX
Z0uo8sbnJM9CqAAXlQgRoQ8aUAKCXPpE3Fma1fcrVtdsCo5pydLue2CnqdySomJX
yRgR4FOnbNxt5ADS1AOiyO4+497RnDVdAGKLAOq5xRc/TMH9TcNGePRxkvBwIcki
76CVvubUZsTP/ut/4Hx1/v7S3eQrD+uynniNILnm3/hgrMW4iJ1peZwdiK8qFD6f
08neoLVjVGwC86VgtN4Q2UD9inVOylRdyX7z89rPtitDj9mfoFMCMEf37F6zIlkb
P/OehJP5PCOYkUjIrfUNVwaJOgeTZRm7Fd77ueataSmFCugMcrRA6rEpgevDlyzP
Oroy07U49AFl0QzYN/YUXjZ+O/bFkPJx5QXJxA1O86FjQeAfiX8hDFncjim7YxMa
hlRW1aABSBTRAKIqs01o/cFJGTS5oHtSYAtSwIg5ljI4LOQq3LpUvUOqDisdKoEs
aoEHbNQ9PiX7IFz9k0sMIJ53SgAi5oKbEMcGY2d61u7u9AwgvLpV8AkF1X0PGzlm
1ApEqGQOW7gjFrooVpSluJDxnAh4rjfNRrCuypAoNEf0mlGREuq7g/ZgW8uMNsfV
vtm4XBgR3rEy3FsTTtXIL2yo+ZMjMaUX/Zc04YOvDvnKCzLovb1rXi3Mz4rtSXqJ
TLZZvq77sXA4zNHd3eRdKYLpp5uHlGVZg+fyDhDagg7tWsQD6jueA8gU2WoZp76m
zVLI66mZpBhxX6zErG2HWPDQvg7eKifNLC8cg1IWqTj1gHN5ll2QQXd3x99gY0QN
9eLJyDRkNR60BZkF0dT0lSwzUjySRO7umVN0Eb2879NHTC0r9rhhCL86fJnPU3tc
+yD9AjslPze3y/Ui1V9zYNuRmjcDfBz56ktpX2mAer6DIkfYc4UKSTiDCkQMAYIy
fb+buZ9vcNj9+Rd/z0TlEp8ogoj7gbpUsdbIs61rA00g8cB1W71U/Dz+WQkZbi1R
Myx3jnJ32LTPMsH1je6E1EnNFChSx6iaZFMIF5nWN0Hk4JMtGrpyaf/SZWHI4cSc
RzH3Rqqs1pF12dT3xY10qk55Fwf3lC/qbtbIXqxVYEofiGw2zW1fivqB1SF0rull
jBriHzPTJRsqvBOVFYseU2dTxBdFPMHDlcNgZ92AM05N2nYG5WKjAuQ4kP5czhz2
nwpKhTEjpG9motdyI2LEx8omZIdN207tJgiXFPX2mahjdk655jcJgQZghzxaCtKb
a8LuAZIsNpZr6r9nUCabqSKtqhieloVRbPGFi2qcftiLlDZptddfjXs3wAarqN9O
ouB6xLMk5yf1m45mo99Iv5ndGqIIHroRtF/sDIK6ZfJRFlDKyNhZsgXZqffpw0RG
Ah28M1IDOxaw57ovdVvbjRvcfhU9ALcIClQI7Id4L9d0mhOil4fEL26oPXd6TTub
6SAHIjiNwpnidVGL5TeyuuiFMce7Vp1QXKJFI4xa3bIxl3sW7khstkIMsxjGcIpw
qII7IoI+hAImBrlZ8libO10R+J6rsw9k/3A2HcZTkwjnD6UaKKswZiJljo1RteWE
DUJp3TMzEQLZFsZXkzMKfzkZgqzGW3296j8TQA3shmLXH2G+JLqoH+HO7x6GUEJZ
4Smw95TZTM4iyC+8+JEHodBW1iQFc5B+54sXgVKzSYN27NnFJRC33KuRtO1HvIJl
Cj9rw9ukpM0I5Vz41M86aD6K6+yOM14TlYlMCxfzhT4LCb92AOY47jrFXQdK68E3
aJ3DEe7T8FyciOtJggYXK9UpU+dhUHpygEp7dQRvh0YvbFoVwUt+AVeva86rgwsD
u5aU9lrc2XqatrMPC8+GP2rKxTxKGtqZixCSiWVOMHH9ocqfDi5NhABRq4vuu6kB
lw6TGNlsDnxwlc1f42bZonOQCs6fWAyYUDOy/ZgnQImotmNGNPAWMYnsd8BekXnX
koWyEsked7WpOVk1jEA8+8qAAUX2A/dACllUHjJY5oq50iBohEteP9Md191L1zie
sBBbGGwJZLBSAMqUOc7mPZKTYmBrSXjXNrNrcDHnujbkB7iH2xQDTmpHKh3qK3d3
PL+ho86bUoYhlZqhwrTvxhB1l98IssNXL+ELoJvmNOc6B+bfFZ80mirc+mi+irvA
Pp0X45OMscs01TefaudZs3OM/j3i/v2dbOQAKh0hQwrToEmMzVmD6RDxqHm8iFwB
zYNoxASLM85lhNY8fKnmQkVtD16LAT8fYgbfYFQhXgk5b4t/vrLhgeVJSeFq09D0
dm5Bv1Pw0njVauvulQTVo4HgodHgZu/T74K1WNL+/8GBU//S6Ndrvyebvmp23SGJ
LYUnjcF+ZPIZtGlt+hdzSpW1r9vCNmpea1+ejtc3DORqaa1w1/GEWm15AQy6QYxN
SC1efn9BGyw8WxnyJPmaOCI1+csh4MeKZJmXlZSdS9ZR/37Zvj2Dn1a+RAGX5R/4
cng8F2QX0Y6g4/8vHDJlnOkOKn2psVnv1iAH0f8G0AC7ixDhNIwpv4fGjwJee60w
BuJJSUNRe17Oef79t4sJ5h/3GIZfxp9cliUNuVdVZ5zSp7VqlXFhgbIZ/RcUdciW
Przg0OsOWv2gGW227NRjLi/YwS1mxEcB+pOfZW8bvOZYzUNeX3HCbrdiZLgH42S6
18/ygETPP95poLu0hnIAHEnovCeVDNZ4dyNBdiE47166UjTgBKpHhDgcCFoa+9Ru
OkVt7+jM8WHwybdvhSGLUQ==
`protect END_PROTECTED
