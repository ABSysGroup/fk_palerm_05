`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2p//7S9JC1ja/cyZDhXamA6a77JICOPAlZgcIaH7fDt/7wqYw02dEhfvcnEhSvcq
m/Z1mNQCQGcl3pGWpSvHg6nD6nwD3LVX83VAa9BlUsdfHgEOrBLgywp7lR4HPeJt
FvQZ13sTF+SWume77cXZ1DCHjetveuctQuEZLFaJivu/Ycq+lZ9v+ynriojo03Fu
IeBFwqS2xaaz+o5JQxtvDLYCcPqNx3S8aqH4XckozdnD5wpzX7CFeW6pCKR359DE
Hg5kpq9pFL8+tRylwXzptw387XDoiXC1btwft3vrZXqUbijYjXM6KD5wL/JKUyvu
Zm+nB5fx/10f3jcvppAokyEJnLqAYWEpzU2IxDRfIVQPo64xUCqAOF8mH/VWz0dX
tEsF5STWIiM17wpvzgYnud6nS0LtSmKtQcAn6aDwSccJ/UXJntP48HbchkQd2ci1
JeUF1d2wRgPDRfKOvNl9doczYxR9rHMUOpJC8eHVEcEPpIYMnb6yg/tus4SOz/Tu
3WWjKlstrMJAr7BaZpEEJ4Cl65egxRJpavNMeVUtoi51LF1/MNGysBcF7tbVlqEp
E4Gj1W7vazI1vaFfS1RDZhiGSv65wzvN1VtH8ZoukAo/MxZQa1c0KKV9sVwNEm5X
YUJQiNdl2VtPIBjYu2oezZoeSrEv13nxgPCZycj69imhDjTkpmcqT9Uxo9MxVSlo
yN3kKnpZt3ooQyakY1ARTJDYMNefYiUmbbhVVnazRoLeHh2+M3gPyn/axYXyXcZZ
ZeA9OX0LfTWPI7/IOWN9vD1aXOwvhjW/YeyB0shUEKM=
`protect END_PROTECTED
