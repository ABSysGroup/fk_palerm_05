`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VknWXh6vO6u03ybiiBn8/oueL7xgHnB9+bogcYxrKhjglvPodw5mNMgefLwZncz3
MxZrok4qwxfLPxAqfzMLaL6EX2zZ051lo0/QKtLxeXUgJv+Lb93moVui+luoAidW
4YARTmPnPTVm9Fe7OPE7QZI0pfJoGDo2uZHQJ1OV4093NdcOBqkRR3KjjZhEMGWs
jcAyb3JnRdSa4LY9oD5r89bF1hwSb7g/VmKm9OBZjXlSR9XLZcXfhonJ7JtfBT3U
Gwe9S8srAnkk7B4JyExc4iSBl++DxInxdVTuFX+B6bm20pV6d4CWV/1Szln9B0OK
667kJzM5i6VoqR4UTeXamYRbEqRvkE5kITudPXuQlfM9yqGJkvi9TBPCNhoYJxcK
xxTlBCsMSvLE/Zb4+dgW4bfz/mfnJITbczKhmc/fUC4zh+TNA7dommLxT6yTV77F
YqR23p3i3CNf88U3lY3SMtRwfgtOdGbInm3Z54gvFR/q4/uXcxND+5/GWUlLh39s
urd7zatMGVUuPxSW7mU9wHslS+tpHiYT+S5RAhqqpGriKGI+6XbEZWBI0KMaAbaN
UnaoAjA5+15ZnIyZ24RlAGJAKIZfXhTEg9rf7oZIhMqdVC2i4HRQ6mL0Tw5iHpJQ
vQoZut3w5dFxhYLwgfGHkUF2JLnuDIKkFp4vo0VWIXVLD+1nkTWSpeHt5AvP836b
MI3u+tZAnxMsQPUJmlxIxDAwsK2zlKRhbgVFRZ0VgsHaxxfZxZax2MZOVyaAzzQw
PXcZLbp+PmcwKDtuG9kGeKPDwFaXHNTbI2e6vncdbmm8SbrFdR2l/hKEfmEE+URA
bR00aTFotlVDE1OkeayArKTn6bNOrWXwmKnCkK9Ccl5wMbCAGIrLT2xxA9Hms7KG
qydCI86t3w4xb7ov6SpM6gu5FXe5SezqCd8Q95ccJEM6+Q8WUp/z2viFdm+KcMD+
BGgcvDIgCyXYImXZ94zOBJkjfH7uz1hnDqRduClZMIaeedwnNyRsNjHYlFxlScNk
BbASgXOD8phVMHW02UcLkuJvYKaqmTIODx+EJBgIdOKycADQIj4dQE6Dvw5TyrGD
YcpRXsqReHyiqU+v4ecF5ze88CaY69rYqWH7M6BFOVMX76J17wRataFqsVuhOtWm
kteNoMFDHSp80WLoYUJCxs/Vnn/unGcxqi4hxd+blPNI5K5TJgmQQwFglbjGP68D
9I8U9LwFPOMMWf47HG/2jZQB1XWR6ETNCSnDWUkELuaBxA+WVLRJltwZ+NtHNNFN
RTnCK+pAfmeZJ6fbvt3SodSJEdGTWbGMhLnYXU7MBHqZutqu0oxnVRWJmuWiG5/u
/aKtYN+YvKEDiQix2QqP7lD5Balml5eSdUpWLDQeGZ5FXGMub9ILq3uqRxv53Zif
l5pAthZU93mos47cLCKzAAoVYTzoBGqeq6vRjUOlArfSRZCzn1Dfta7owlb+/n1/
4a4yF+GlhWNd6tXKmW1ArXlnwghEgmYe/FA13WVzKpukdzjKVDSOwm5q5xQ3At5v
Q+A4WK8LbEBzsKLYK3/wNRN8uGvpo4ds/pPK7tLQDX+7CAPGyudsSLG0ob7pLJtS
izFYdz0mKWrtZztjKc4WvEhDZqc/WK8Bi8dAUwukovxmZckfyW6H8wktKxZdDFb+
eBlf0lwHPtbLyZPz9wFrh0lhYZNVRbRCRuWMdiGm8+Xs72W1Bu6QmId4xVk+RRc8
sRJqK6HJ3REB5DyVhdTwSTFYgUuseF4dyaUVTRzxrlo4NggpESFKW920Ynr8EAjk
`protect END_PROTECTED
