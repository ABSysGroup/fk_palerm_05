`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EFpYSPa728nhDTdaex5i14QNFwl3G2TXVgcHMQteI/psZdpwJqUb3obwe3pQioMS
yqnkZI2VTvIrQ/l65m2BaQKHScV2P7VFkYALSivJvbi3obOASOV7D9XZPpXFK0Wi
L/Jf0Rwca3D+vCtMAHL6vTkYHaL3gB75b9znkOkRe9l8quwxuULaf/87xlw5KUCz
6HCpkz1XNLvgnr6U7cMk/jqt5hb4WFT1mWG+OmtEKkYtC5uMVingLRIvZkjkuOG3
1SO2EggP6ZvD8wN27vYysUMycXucs2s0N+nsy2HcxuPI3OYgZ28S4Jt2zUjZVmdM
xYsrdvMLVnB37Yv7ClEeNRqeOI+hbBy2wy9FBOtVXVWWXhHiA3syvVgj7+SlWeXr
ty0Oe4MFuYjq/dHs6R3pfmmIVntF0KlQjD504Nq9q33Hf0oIjRuPyNxnNtd/NUHh
PJ3sQsGqOWGHXTG6ZOPhOgJtXNmjcTea6Wj3hHRgh1v2xdeBvkN8k8OLpKwE9+9+
JwvWyeLwqaujhUTURvvMv0qWGNt+Dfy9Z9BdlZwimxGAx/LjMMkMYpKyrgoAdACD
jbFc2Jfw887ZvF1aUy+2UdS6F9PZB12kMO4Cukm6LK0RS2mnWBrF3kjyekZccnxt
qevUYVyf/k6neeqJMqzyfNApJXPT/yQVFgIxyuOQc28hYiqPlw/jyBARw0uvSGIp
F5p27HpuNtH0CssKuajyWc5YGe0wSXgEAQPVpjSa9l/LV5VvHxvj3DD4sqN5WSKK
rQKJts0GELLdqvrJVypKjJJNDsqQvupuSPF76SCmv9o3g56Y53/Ft6UYxkB5g3Xp
+jPSXCfwgKj/cZyiObQ+1TY2GDJT3Ot33wMIYBhnVyX1ToVmwVs5bh8/6y1E4aSk
m3L5d1iJqxquwFx0WYP6Yc8Slxbn8WWxQeutZlDYx6GwH0gxU+LqYIxgBMrqn5Kb
0I1Tt+9S2lk0oQSeNW4MbcbcF7qFmS8dza3p50a5kRLGqOdQQ8WGJxYUx4g1ET16
48eINeI6oeop2edftbyxtFbwMnsBAYrRJcJgpCSgYGw7s7IA5ZmgulqUijVu8rqq
q5+1UEqfEef58bXHCwxi2DiHWGKVaSdrNo4r1QWoev+Aph29e1vQWpFq0VbglF89
UOuYRWd/ObVOe5XZnTp2EqsNEWaDGIWQ0s12qJrJ3h9Ehyz3axi79/+hbRk8FysP
ft6PFBfnX1c2l7Ah5r0oinTtUp1vPG7e8YLEdStYBeMpbwP7IP7apnbYP6opKbOF
hIcCZPP3Eq06whYEO+hs7PEhS95jO7sbhlZudf4NBglefIebV/iIts3btwP0aRGC
xInApgEpOGWARvbW7Tn0SpjNi3QqiyaRshKjbVe48ru+1k6bIJqDqtdj03x5oI1K
rE5Eg6J94aw4nPiZZCJRCmqFGDwFOBItZ1lDw8yr8x3DxcT+UB+H377bgofR+YKe
5Z2a6c7HTRrO9tX78JdEl0qUKrxDZdO57BOdPqaRyB0pcK8awuDcwyJ6chtFsNKL
A1DaC8XUQHt4p8Vxkdz4nCdBXgW15lChejSn2lbyWKQLQhhLsbNaUNtPhRxic5Q9
coVvDPWaQgCFOwC+HFmCJX6ibxEE8E30oubPvaJdD9745h/EYMDFeLd2EavVJ31u
ziXU/3AVTbz95hlONAUeaYteXXVhsr6YoBq9mVg0EBeQoZQOJHnLO2FCKoBxR+ih
6vIBfrnScdU3+MTGFT1W4O1lr+dJdvbgKTDy7DGshB5DY/cTxqH1vm/vMl9DYJ9W
bxwJv35Re06fZU++gMWRyp2AZdAjAqJ38W3kACl6PnCerumSM7xeaJxv3UgMlELP
xTY95zAkRW39TN9RKZwW4rGlAQqyMQqPvuEVFmE1U6s9NRD4KlkeUaXjo7/c00rd
XQ2wSCgbv8CwJFFDt3u9iIeJ2PD3OZPqBr0VHO/G5eG9K4NnokY6qeItA1NMVnQQ
FtRBf3kDgvN8SEflrpis+VZS1CvOqXLYaN9CyAgjajW9YMjSaUCpDvNgTPt2GA+u
x8ggi+eeYTqN4YR0+NwMDAtTkV4muuMU+PTNOwK9yAGl1OKJgSdc3FNTCZymSkNc
SgkJJBjSTAXv9O+wwP3wbB/VIokKC9rDtzbSEBn5Ux4/seUJumoNyhyhRAD3XIRD
ylorLVwAUzrx4btiECWEAcx5hkl2knwFer06zxF6I+ZAoUSu+1ul15wDhFPvGcuN
WpIAdn3v+XW1BwvhM9nJqMG/8sxsidQoa2LO8yuAueV9mdz0UZKQdkiqkCWF+WTE
SwKhNqoBfIXu+4aGob5S3MKx6e06TGPenFSPO26o++AMD9l/1AXlQ9LPNUpTr6uP
yX8yeKP03EKnJgtCSkhCliXHQ5T+vOunQOvn1sS8kZ13WuIkHqhwG6+e6J1e68T0
SVqQ3saGxLkExF8sRy7YV9ALG766rqKfE0rIClTHm/4Sg10ACge3QGJU7MjNyLFu
gwE+sgkESlfmaizxzqDT3iZe+c4f0ib4LFbEBcw+o/L2UwGhY7OS8nnMp1UuFpWX
tzMTpPKTl1F19R4LbbdrDftfL5od+/qRKZSIkMT9PgElzvgGWRDptO068IQM6aUZ
4xINJWJ0YYeD9bbYvGdRG5MsQ54xQecLfb0iUftw4v0rNzm9NNgtrHxes0LDgCwp
73/XFcBq61uz+1XYtmvN63zIXEEzM5EfKLIhTnPc79fXIyk4bEnpcBOtufAgYBoP
TEumg2BD4CnnQt0h663izhpxLL7T3A6RHXlCEk91T37Ciiz3RYIfb49MoxgVALIj
7N7ct1KWXSXRPqN+7NhynTX88iZHr1/kksF8Otkvlx6WuogGDc0V17Kzw0GNw+SV
Z3B9/e+gzRgXBMYQLEXWFrPYYi2YkRhLskgm/Q1hR0b8JhEoWkm9qtvqe3eHyfWg
KJjZgUTgQ2p0pLJPx87qYXAU2yuZ/VwT/wn7ZpUWdnK7sufBBRX+sXeAxoqT82mH
1nOO9pYfdiuMaA6WKEwVlyTHQYJU/OmarpqjsuEfe+RP48Jv1D/6oubH5RaWKH7C
Orxw3HgqEFflJDFeSCyADGcvTzgPg8E83HPEnoocVP5kWgDuG4oay1Zl22nMBoaA
ae7sz8DbdeHynduc+SLkKzqohKDCMxmIXODHjSjHii0rpojgdbSphYbTYp1erCI+
OzuV/zOow3EO1ehDqXgbe8tcPnC4hg1CoZry6KCrsXe7+BFuZAggwhtK4p7FHe76
OmlWWKiD2lSKA+jtgVOy9MZGWkp68FD+kl8e6X89+ppLqhXp7rzqwto/6/MV3Upf
rMxkRKzQzKXqEUowxoCpjbr01J0192dO0z2z/R2LqK0HceVwhrCnLuDIr/3QD8s/
hNEefGO2gUxPCxJ64UKiZOIb/DbeG2ezLPcOl3s8xqATw3KbEkfWhWL5I+2/faGN
BQx7883WzQBC3A9rV7x/psL6xPdgt5o4kNssMoAT8oGl78SGNiFwsTvLjfD8l3C2
NKrPrgeR9hu7pCWL1oIp7V0dGVl9JkgspTDmfi5doimObKoFFpSDEDwN9lGnbQgA
x4Y8XYBJY5onOS7Bm1ZYi2VWslvT0wgk99RpGtCLF39I2fWwu3bC0vsbRBiDVaug
b8RvmAq0sFtzFxhxXo+H12Avo/aoiKsXFW+RhXwkYrH+gBePQDujYyLZ76J9hlsG
lby4idMoHDwjmnJVBrGCcR1N2UsJUZy3FHXsDyPm3Wvm3q9kLWAOMfoe2xkLzVnt
`protect END_PROTECTED
