`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
18Kiyz28YLJ9IuEmvehpOJtaynI4I/eqwFqMR0Yk+E/B6TqwIW4cyuzYhGYcjm2w
4eiskf/rexQPP95BI/y049F6Nv7o7l7ZQB3aIVYYgWu36IliP8m/fIJJY3rrQYjj
M/1gLm/SjH4kl0FNqNHhh9GSvid31Be8dPQQ8j+PhjAorBvhK5Zg0wBMBme70tnb
MgBsqZ82DKg6qYscc8rjkXVOpsAitn5ic8IqoNK6JzgcTctWxHaaHPwLfMivL7Zv
Sd+Lw2pebw8VjvZF81NYDISSOZnEQgXY53spA/o51P2bJrdn6KfRurLRtqsUe0Cn
Id0e2ZK9IDeMcRowoXsCWZ2oPm6WMSsWxyY8b8H4X97QzTpJuIvRWkvHhDanFeED
9hp2J1DIKWJCIBz0DMAaauJpFiyuTW7M82GGYwT/c00LGxqKQXMv4VWcCr6qGEaF
v281UjUOxsb5dG9mK2YhidbK/tNmd73ZixsHb7DdRF0+U5E6qblQG5MkwaS3eK3l
32NDzI2m8fj/xfX3dWbqh2pSdYebES84be9QXVUu5aH1NUiCQK7zjuAlFuCynQT/
Yat8aGPnzRkdJ3hDWbHmb/FuF//rppN4Iu29hnRDU3mGsHnNsS+uuujYQJXPp9xx
PArjgQYrxhj8B39VA9SB+pMg2HvdeEeWPaPv/66cHEs=
`protect END_PROTECTED
