`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9iin3Fb7XjHdmWx5DeIbXESbttwqSeZmYPJMgRFLbtoyWC85nOK0aSKoekAOniHt
JBluTmSXGVSg+s7GUeh8GtChMDh0PX/VYY17g46xCLXyl5bebEHaIQi2+7IeinYE
EdKR5guj4LkpTx2IvADbq6zGJ7fzNJAbCPhSTjXsE2unKERn2niXsbBtflqX7MzV
yX7pDV9eptAP1cs/NGKRACZJSH6o0Yk0bxp8cXnlmDKHPAH/yfjFC8l8paB1UtDG
QzgkfHolaWTi0llfUMWZhSxztAglKfiUqouHp60FUJt4tWJozBoaRf5lvb48isje
hK4j21t0UwY44jEU2GDHN2Wu1ZncY33ElEFh9OaOqFdPx2P2s98RuvSnuaKJcxas
W6Dhh54VgvhTzUCcoqruDCs1GvLlyPxkLijQeFpg+IhwJrYce3JzVrPqHHksGo2L
JIPaHywkF5L3PBgPTphtSOW5Q7WdtEDbAzp34npgomnRZwvqkSTKB85chTHB5klD
m1P62rdKu5EJr06GOygXJpiW+oqmiGfpdRgPheg9zJDwcNxf/vjjFCpFXb3l8gPA
AijYOKAKcDcLRPwUGcrslqU9dGYb13xpVdtC57250k+6NAemecfCiCajS7teuyPX
EmIzo2/VUzPTjaOHKS8v2Hdl/nP+f9mFcL693NgnF0bCmRtqoS4qPFk8swVPWr8r
VttUPptaAkhcVgGYYcWG3Kt7zt9SgATPU2ddtiojbAeABVEyFmv3293KSYyhdcWv
EhjdAQEIpZRxF0ZMfW7p7jaiKaLeNFuSOrvorXSsyIaaV99YWDT3uo6DTawcFyzt
dTUTTCgPdPcNPlv6rHxCgupgapWMFVWmeI8daX7EbvpGjY+bdHTTZ763HeBbtAgW
f34cvhk/fdUHbFHms7JS2nIf2I1tiXGXB++Pol6MOGK+zJoGOQztxU1xFtIvzOYP
`protect END_PROTECTED
