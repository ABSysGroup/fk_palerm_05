`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5exN7m/i2uPICdkcBOfk4w6qwcDD2uXG8omEcsbqWaZFswLjz3Qu52U6VMSvt+nA
AmJlH9jm5m+MYBfMxQy6jCkHzCUPuW56XYFbRT1s2wGX3xVBBz7jJqUR0nDhSQO9
brSceRTE3bG1rWwGRU+cyERki2jI4aJWkHebI3ZaebMoQqOfM7my+IUo3+HPQ1FB
xz5AXSOrYUxmzBgMoYBidFd7k2SAbnksYGCPEwXYm7RjON+M6612aCEEPc7mEd+P
0N4FqTwXcoNtnxulUPT8TngQiNiVgA+Ct4NEL5Nihmt8y8DMq+CWHdA1FPTmuwyh
TVPB/UFTqLpvdR6xV7HhCiKw1hhd7N/2oCUxn1QIPk1knOb8IpxsU8KCRG/2ajw4
z/zhW1Auz6DMgimw25Gc0kjieztqnIK2Sw0uCudWw/tYRn2KacSjmTHfiSpLDos9
`protect END_PROTECTED
