`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w10oiqM7o8ILFONIeOnS6Xwf5BuRWeq+w0x/piQt2FXNcjg9LLlKkw8yHETo+RwH
RsHfkLfJUbP5JVuZObc5RIkS6DHCVJKCB8RjWTqzhAPGTKX6KxofDy37MQxOwze5
JJ57UEwBuYRHNR4l++4cvISxElcFqo1TYdgdxMwvHyQTgktsjcdyzTnn5xWQUkvF
uzb0vwdKT1p6O2ce6CI5D71UAcvW2fmY17q4kg5PYOOnCi5Do7s+QusDL68PEi2b
svf3tsXYB4PM49QkvsNoxOLGxZqxr88nNgBeRDc7dXv5IQEohaUui6ctAPLY5Jce
PcBQw7xjGYuolKdiR1+5+Q==
`protect END_PROTECTED
