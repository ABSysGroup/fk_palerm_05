`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F0soTmvAnRdKs+lTs5yJypleeis9ngASpzEb3zgcDDzawULyl40NAm+Xx4CQj8LB
Dl9+OqjyhvZkro+ixGaLGkLScx/7yLDwPd4xIDoNU0C54TREWpamDZJNthKyNcNR
vTObTbHQzXz/79tKeCvjMIjL8VMEdc/vAQoepMl44iTQ4D6nBZ7uP9Nn6Zv8tkoE
jLXeEWkVG6GLnWGx1H/hN+Jh80tuiCVYJjmBBHoU/ipYJDbhwNE6JJjgOzR+RD4e
M1NgZiNvJZQUNOYT0PbvYdQmz0h/w/a+EaBExnIffVDoJ80yv/ZSj0Y+FXiyuxsM
h/JirSy26SXfol+qm975paK/yVUAsdUiznPWB+wQNMBpC447mC6NQa0mWvXPXKva
NqwYlHJ1pcotBamaMoHP9rlLZEtsnKOteRy58eFzPcKxW4PUkRtZXpu/iNYLBbqW
VLiJkW6o9DCT5wabK6XYlcsfSWj6XipSXTWaXD6r54Yszd9NNBXDW5mTuw4WDeXw
6ocKWGa4VxFSm3dGqwBFmGwhKNbqIEUUZyfT2lBIG+uVnDEoMy9O8lqaTtGy8WZs
Bgxbb/6lo+jN8ArG63kP0tQbc/pQ2O+i8F0r6pvQe1kPt3RziBjPLExBpvaPEj34
GKf6yYPcz/7KKu0kuG7XVP28Y29QAyp6ELtH7chfjMTK1iGzvw8jWx9abm4lbBml
TuNyEu6dRVx1dsxZjJBXSWVfMH1zqRKU2AHJ+0EDWAyTtZayLuEKhqjhbfObFBRt
B0Ccqbqqz8uGHcqwjFZmbKFhtbBGmdlfmnJ5XiUXIKGH/aIZtSzAllQXkhP1n3Cr
SDj6FBFwPaYfcfMROaeZG/VZ++IcDI8j4aB/1C/CXGRzGmj+mBMQ5EMK6Zp8lJJ9
7f19YDnXzblUbfwONXRpFqXEPUbMAsPuLvlyuDHM4qN2c8gTDWNWWjpy69BngVa8
`protect END_PROTECTED
