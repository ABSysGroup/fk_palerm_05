`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6VapUCkcjk4XMnTz99tlO6WsjgIcP2h0SjNW9qKLcmJs1z/i5Vchh1pfeFbT/T06
CkMOj4Y1FEWMtnZgpppq2DoNu0nSI1/pLnypGpOz0Pa3F31UmRaDJVXwIihOm3NM
XdLejQBKiWZbW1PnCOpok3x365Hh/EQiz0RGSLwz16Ulx6PIhDiRyaeQ3fkUmsp0
OrVLc8eyWupG8D/TuXXReGsDNIIIoPW7p6hPfSgyqtD0ujTKfz5u9QulUKwq/fu7
pcNu2Nt5smSLrl800tOG5kTwLIewdB5YqP6YxZzYTOWH+tkXrH5hHNMGVsMYQ2XL
+xuAqf6PBv/BZRdTE3pOPMHs8SesMXJg3Qx35GjCYRhimA2rouvZAe+TB+Wa3/0t
LLRgaQPId9s0K02WMLDBKI2EfwvHKazVjJPDKCVX/uZQ724zI62NYwI/hm5eeSry
B4WQB3Q9r0q9Ry7pTaNB5ZjOSdXe3CNeVzBZOTI8UtUOJMBtlu9V/YillQYD9c/W
P/cFvWXi1srO18BhimTt0RZ7qqNIDXTIaZ3znqJo6x8w1A62Fnos0o76zT+EKzhb
xPhHucd4Mn0ZTQCUsoUrNa+wSGeFSCZRYrl6DcE8FbnC4GPYsAr2pR3vrKswNPtL
o7tSfLjSDJFhQBwCSij3mz4kwjkkDAT7T+zctn3igS4=
`protect END_PROTECTED
