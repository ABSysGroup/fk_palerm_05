`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IqckFwuJtb21ZlLKLEaYx7WOfc+mWh46yWrpnjXHlDHYwn7ts3hPidmWOzUPoUKo
MC3o/aEJdK5kUsFOoJi+KNQgYuyedUIWByF7UA/zeJTp1Bmka58Yr4zT0IsfqywO
8g2MDTSaa+ic2JPBvPySt1HN1TFOczOsq3Le0yCSOSXGFrn03z2X1gOYb7akux5m
nXRGQFlHTYOWZtdyzfsgivRKLe/uNnolSbOCOMVw8IK/9JYP+cEHe7tUQShm7Tyw
0+cZCNnpGLAbTvQHVRV3fL3sMaEw6Z9Y2EEAmn4Zzz8x9JnjktbMF1hgTK9JyV+d
StPWv+9Le3wLEHY4gXCBhneJfA4M5EEfpEbkt2b4zpAUcAtIOmjZ+3+CwXB/08b9
J2FxROhXtq8SUlBoBoAsifuncyNXQN89g+DcKZtVq0GHnyXRjX8HIjtM7ckhYt9M
Sbx3meYnif5uvcd8etcRf8z4K35cfyeRFaBjvMOzZEnaYcDlmqoqltedwFiV23Oi
23XBmmIS5iQ8K/BalQ2hUsMqey4+ZCHrqgOkCssmiZeJX5O3ChFpqx+4Z5juLPEV
EEW5ZroRyG9ZM+LsQzo83hIoU10pzZ5bBdAnz3IuXtMTttYiAsvAasT5Bg+ij4YM
75HnE2vgV54j6kmlQv+HORQyXFlHDCFvWsXuANsNrYNjHvqIB6vv+klRvxNZfNRE
nVZimYTQf3wnuOJhkS1daS9MRr2O3WIwaEPstZ/ZrDYGOQJe7W8Bw5HREkjcsRFX
K6DTatUOe3VbhpHY4bof3KVtlKvsC/VdU2kTuP87XuMNmgvBRVvloMI9eTBtCpPb
uc1GQafrfXjFG7bDE9FXlSosVQLCkoJ5Hbxo1xaH4lY5Wb/6iWcj/X4DNOBUO+El
c5/4Nkn3pxV+G5SYHVghM5P6KYUeSbrCzGrYIKYX9c9FEtOQdp37y7LKsLvntRm2
Q0muLnWU4yLYuPvrvkwLx4M2QCFcFs9Sz25R9JfTlz/RLvLU3xLjRbX/nASWh3ff
GbqrNixV6k08xrLIeIwaB9uyKji1cHTmtmcVz5T+dsheZkGVwaVjBPuWCvdHN2n7
mA4ZUfawBsvaOK2C4ZGRucNG0UGov3KQbzlVWFCnKPKchUWY6UZcDII1ch8aF49l
`protect END_PROTECTED
