`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tcjEExpgFpaYS+3qyMwzZiSqha3YZG0VxMDXotgt3bmpt4rJqHUeIgRc4rrz3nKr
BLHgaBtHAUrh1eGvh5xXuyBHQ4LPpWuCucBEVFF+xW+3/DIHnSj/k0lzm9uBJADJ
V0g+Z4ovOTDR64RQpwgyw6I97oDZNjCLRhvyhosIWeRhYt0pjadgo2TBmJwB/JP6
ES7yAgIVA/y84+268RA+b8Ltb8Os+0wO33+KYUUJd7432SwStoky8UovZeJfpMGS
UnMJ+zRZ9hQ/2zXnpFI8eyzQAsbGGYYFREO6Xtwb2m7+qD8/FOC1LTYYtYF55zNY
6YSusHLooIEK5ir5n+wN2zFJHrQmz7SuHtNQlqC/WTzVRB6Zs2jGuiCDOo0UbVlu
axD3AHUCUZDtHViz5Y0dgAl+uyHc8nXGu0Ai394/T0o46llhe4bbMMEUuGF7Anje
++8bPIC+/fwXQ/BpsEYZ/WfT+Nr8NcHXkUncNingSjuwdMmUmc5PtthI7fuf+6ub
kz2z5+z7h/S9Mr9KWr4Zw/b3c0GYfYOuV/9Vijs66xOHz8Trha5bTy/sAiQfIXl2
DyhpIjLGhz1v8mVKDLI6KZOstUwgqDHQ2GTBOZpO7h4ZssjAuugCyB9dJmGY9nYP
EOhWBfGk5aJ9kn1zFxdHNYWzFRDHj5N2UNvo7c5Ew1uJ9hFTAd00T/AvHrEPfR9C
9DxaSFTxqPB70cVMQ4OANlY63Aw5WiSYE39Bu/p76/3vkKl4ymj/vbVWw0UYC+Es
WnR4cLX2PF+9hGX/2LzvuVp+qc/tlhAT66cGeC6XqLVDGnU3v4Ywx8ai2CfliChF
Iz+9HkV9rp84jdl2RPV3kjbF3IUHxz1EmeIdQL3rplBiXoDT+3tUst4rHjB60yMp
2bzw4Hl0i+8iOzhn3V5CeQ==
`protect END_PROTECTED
