`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zunKY/RlQKS2dx36o/dKI7dqXe8UH55Ghw/ihIhEYF5i71HxbYaz7XiXR5lnwm3H
SlbSPtvqW6lh2j0upGKh0GkoezPyOslrIrCawCH+M4sqcYj2yRDpjBZknxKEcK54
aHPB9Vfha3iY1wP1v4GIXygcZQDmJOoFydYQWi7wxMLmOVoE9sMxTZMx+Jk+mHkl
/+AMNXlFYvvPkzPBPqsCA3hUNunKwr7yug4Zi7lflVnEB/n8XGq5EqGCqXvCZ4zk
aWbwQ/4GBKdSnRYTgCemAX3GiRei1DgKMBQuegsLWM8=
`protect END_PROTECTED
