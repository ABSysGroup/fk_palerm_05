`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1j3HNUWguBN7H2hSkOUVJhKCSUURodoHLp+luD5eA6bgQhzfPRbeobUvsWw4axM0
k63XYTBJWuJk8c6ypxD2pcRY4VdkbUMcCsynEuDYHR0XERr31v+MTWzJQZKWKrPt
kmufiYzEpweed7FFoXTYvyasqfTmHfuAkBqGadE4ZLqBTZco1vSqcLRnN7dxnYFk
VEepoPoFwCHq7T7AhdZg7u1XIj7+SaLiZMroLylEgLU1nLPMLMNREQS8fg8oAHTd
PXm6875pRn3gh+NjsyCsvmjv/pLiNP3N33est4QyaD6wtHzwKCz0eHQK1jnc2Fpc
XYgSHt1xJ8kJyxCT91rxzPyQD1QXkA3TwkHzAKoGvsmZ67xrbZq1f29ZOj7ILKsF
rrveq+TffklnuP9dijQplUm5eJyPIxKsJ0Yg3i/8tYjAmPHtLy5L0wIyGi4wf6qs
RybZuPCUpHQYoJmRxJlD13uDV8CVMOUGnN6mbEq30Jtxh4R+rpN0lXnbshk2KoSr
uoWpWB7KSErjM82/3dCYDnaFuS6CFpDo4X64pQYBAR73jTIicefo7ajxL4tvZGU+
`protect END_PROTECTED
