`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gbfJnjk9Fq+L2nia2XcvWE5+UrXT0xlCIY7oFzinkC1zBJidfHEL60tjtPjy+QtV
zLkF1O1Ud+/rQtfCizgXaOFe6KNCqCRGjOKlduLZwn6KmxFU1hk3XUVtKr/X4/st
7MyDSTx6HXoG7Gvo+VSmcxFrJuah7V39eJ02HnDlwJvhIwpBlCbauXvB+H6rxWwq
uBYnfFxtoRWZjG2HkYu7W40R269PpygkBQILDrn2h20DjNjTS6iFyqYhmwF1K9e8
jqqKV9adjAO+2acWPyBBf6R97RMAKN42XAHaW5cgVHJ1SgW8PIwsarFtBiflCekh
W3XmwwbiPDJFSIgI9SxILVs6tfJ2nic0LViMFofhZ2vL4Ux7GR3p5zr9UkCMfYIK
ZwLlOZ8OEuYmvQZCrhBAIvGhKDEElqdmu+zZSxdcOzMcytHnHUr6AhH14a7BU79V
7vsMhql7y5qD5oGWQgftjFcfJ80p30DdQtT3Vr9SLpbcY3fMLsYdTvxEUB/Xt/I3
fxhXPUcmJKk4OZicrg06Syjya5F4U+XxOieF49E8NeiNsfxdBb4PdBg0nNfaofUH
t/lWwxqqwLMlpufpbZ1FXz5ADrQ5rOUDZGt/LQ38EiaIIxZqP/ngLwT2nJuWVmrI
wfY4fPplUgRFH5WtJ52tp3wziMMwwOH9nGFKcU6Ecl4XQE3lX900mlzKfD78L3pb
gQY2rKsqBE9d5KAD3sMEKDvQQ9Ya01t+/ftWwC10oREiKQF5pLFg5u70uNKmVtEf
ZnVm4kWeTsCFY1OmFNl15IAA9njTpEdY5EzuVEvgIgExW120A3oj1E8utNhd4Cc2
dthx7O+jmBcIbOENkPlEDKPgoeDLw6dh8rKuDqj1IewKNEloDMaNi56VGqMfAZLO
OR4L5GRVKBTxDKp8yZvpP41gt4v5Uw7JsuLt3lpZkKJ+7nMp6HYPOpn5QgXb7Eok
Jd6LhPBTeV+31dvSvbMmTadPUGUY1t5l4YnFk7+lT5I=
`protect END_PROTECTED
