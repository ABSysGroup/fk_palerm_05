`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rpfdNCnKJdePvAZL9aeAL8rcoewpTUy+HI9cUYk4ZkK7F6LeCuavuKKXt7JMke/4
oRJ8BhNZwtFzP65fOKibofrtFhuXk0BrqxHkQgCbRkLFpaYBJGDYnTGUHmQZ2X13
z8T8Y5acSkk5BNN0+Tltfe0nNv3sqCDg/t9trDevCd+Li0Aa+BUdTaBhnSUztELF
/oMigO2kAmRnfCSG49rY3ArS5tbmEI5wG9MYUb9k6j+GvDL7qg1eh/JtW9NcyNpV
Ihl7w6vByqvOUuy9zOgbMBvcb6eeoDLRsxDvJTtfgBgUiWU10yv20LbRdTrtVT1p
UVnmJbjHDsTYdvRfPOjzCyvk6TWaZ9IrU8V3TWOGaHpKpmnx4VDj/KF82JTxvd81
2svUQa75jfTWaa7TYas9Wg==
`protect END_PROTECTED
