`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y+Dg3VUvqGdRIhis/SV2fq7Ty7HPLke29AC6vqzMy1d5gCmVpZ27JqiW0dZo1Jg9
6RR7bSHfLTxFYTz8uwNoHv3dB8a+XSHTOMPo72XVR17fHUhh2vLq+gubv/w2HKya
y3J31qmnZttsvxWOhjGBXfih9AJKPRkORddBnJ2DqeDPrd6wS6GqlyMzk0qiG3Ua
XG3Iq0KKF1Zzmi8HOIUyxghwJ8GMtimE0qEkJbzY5va3Rb8PQoTK5/SN4Q0bwgRc
q74AwP0KafzTMmShDniUAATl4raEaF0kWGVZjzVoa0zN+cVK6cW2JZgqJBDF9XOd
Hmko4k1u7aRdLUHBugHBayAKKTR2f63TC2T7KKR9FbS+8NwkM9zGOvFE27G6y+vc
DBIDVPMyfj8Dq9eolfzve12JZAv8MRGV+Cv4dD/o5lCMy/OMnTb4vsFi65ttFqeh
`protect END_PROTECTED
