`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8tOaVq6Rh9Vb60+2cpXXxtCxQpg8zE4JDC7xbTRo8F6sm9C92O39yRqzZwIZcv+W
9ngesI0Pz8u6mKa1b/1UTQeWXcDmzWzj3aDKbokyNky4gn7kEH46B1cTOPtnkQwU
MvyMDD6ZDYqTMqNeDp5AXYRGrrr1Av6tR3NOE1Sg8piXyBXgUAIIBK32Akmmht/c
y5vzV9rbZJ+s4OXhpzuBXvG9LLkRyi7VnLCLdb/dsIb9ZeBPLoypzBUvU1e3HNSd
Kawgk/4GAzsaoPhFrQ2piFxr+TjQmfrh2657toD036PHG0tdcs7AAqj/pYNWpJ1S
dIPQI0Q4amIC/MLj8SvPa2lwgIxZkJRbfdN2NO9JIU9wphjnzP62GPwKH62ib1ci
YZsCXgCC8L1vREmJYennAuKrcPxh+oAX/ZrJqU/S8BSKq0nCQnVDTrAeFUeeHS9N
CryiWp6+B3uujn6BugCQdg5exUjDvlskuk0LfWqVfFUJY6mM0GhDnvGffEy0wM0J
0Fun3E5dPxFGpqTLuZBnpYZHLDvg7R0eVruJ+tLxaqBVsZF9KcqjDw0gK+Q/26Q8
Poa3Hr66AUpp06PSDq0bSKO31gnL+IZQH2ZxJ4VdzHCRd1lecFO5wHK7KGXRwb1T
BTdvCglE/RZPcXal//1SXRqlQe4J2CZx8gfcTLfoNQSn3djfSobVVHrwj0e6veWt
ksSosaMLrTkbyUl9Cq7W2tkT4A1or718vGvS47AKKFhp8GhAx5xft7bHqmWLC27U
qiSva15GxL3+0ak4FqnbtMArpbGITEGaCn8+4+K7b1XSUv3ZjxZs2KITQBDFXkxK
k4BWmhaNxv03nQjlRRqE88gXmmKHu1Pd/VEuLUSF4MAiiV9cH1PaHAB4p8ituT/q
7y0WWWwGONnzCQjT3y1NzT+xQlIkh6rmZrHDt+tdHA6ta9DDcuW62ZwR9iqk0BGY
kyBApDNzUzcyxYi9NGkfb64GVzg6OdJv+/L6+BmzRQ2X/sZxKGM709WthyyWeNC1
CBZw34YJTIn3Bp+hKh7vGRZIKIYmFBG8shzA2vQlSz8kg43xSpKMVTmYVn44k+07
FW46Ks55wEC/QtmJJnfX+wNl+CtLw8Y8uzLm4D2iudz8yeipm/Bwd9fbLR2M1LDO
jMXvaHqlBJwtAHPo5xZUMa3zggHYtqIjzAQnQnXe6gG3BujOUwFgwHNpQuKL47+d
bsjECnqgq9Lnib9pjx53uh1ae6pdibeYgokObfxjDtj3drdvppid+t8QnHbRyzKB
t0dNgqXx06vSZ+qp9lZAstufBe5QCta9QQUuGoIa2H39Vn1ezVqb7jdZr+LcOBHh
/M7HmJq+j6eczrnuFa3TOcaEuNA2af96PAIwXv9Y3tR4ZYwNELTNEBB4d+uinx6X
A2CcrDdl/Lm5i7wW/bBME+HlBUOEVS9/MqQpxOJXv/MAo16w0Xra0j7z8PdiOhXM
oHp5gD19qWhYIUi2yb84RuHPmfs+4c2FSFakIqQLdv/mu2b6GKw1NWSwaMMpzOjj
4R/aIPV14Cp4QLagBxCwYuew4Gtiis/Xjn6uqrI+hNbgyh33UtB2Q3UXzUfUTmlw
y9pNsNHP1EsOz+FJqqKrcpnRinmtOYxAFwleEJ9+YlZeueD6vEjsPYwZgo/NcNej
wDja9EpXG5IZh1+IB9f2jMnkzi37gNn70XuwJHLdQKSRRmpRjd123/hHEupVaN6Q
DBoOmyzQMja1K2eL7+EkU83II54dRWUIt+SDA9E/yIIoqUMwMWkrSNAfCno6+rk8
muTCL+W6EUH5p7iRCTySf8n+cQ0N1r8zeFqUS93DQSK4ZgfR8els1Mlm2FjzGUAc
tinvHW3kjLpT5Ok8S/TcIuS2eDg5RY/TmoKEBpe8ZGBqsoCYpHQOjLUhwejkuPB/
rr4Z/u7lGaifspj+WifMt6DuyHmByENi0tfhnyrFzHUr6WLpZNQIosxsZOqXXO7M
kKiS8u1mQquXvGpKrE7iGj3kv+hecimo2SEHO4ZSwVoPO2fgroE6IKZ0j+g78yvw
KPmVDKydMNJMFewY5as4xOLKENTO8RAkYR2xxjlrd8gS4tunaEmbwEVg1fuQuAGb
oMkK35PS3tiIKSYhDtOiyUBoyALl3FJwsnh+sWlMzIwwJHf0UFNiTwqXlnBcf3kg
qL/e42P7abFEY59YAswlLjv3li3kd2D5Jdc1PzkoUnIFmrX3xNbw1USbc2ScLJn3
yzMmqpuZJkpr/hDP2PZqzNdNGumApALURSK23F7/qK+SWnFUOLT+nTh9lEXb4SoB
HWBMbFMD4pRCtGvddUtl7sDuKhp+YmhEUNY2f8b5YdgpaTmCWLVot9wpcMfHEYsw
aH7j9cGETa0NZ8AovOSsLv8NDh6TQyo4HNHjB61uVAfplR8VtDB6cNyLGu7NWrTh
JmXN+3RjTEiEIwynhNQuzcOpxSmtYf9Qxom3W2ym2w3L81/VgLJYM7ygd5GNLAIf
oq6nwzuILl+uA4wdK1/bCmB1rY+GI/jEbKGWnS3j8pBZw75l6zrSdvA8vybHBQaX
qdGBPDVqrWndk7NczLj+aqvB2+51/gmbHnvIoW4Gp8f4xlaB7j5WiOkmX1ms3sbs
DNPrXiR+PicLbOqhKKGKsZdPJ5iXzsvk9mGd+suzu5lmEFJCqD8h25AV7UHjs2dY
UmtWa5knc/G5P5oufe9ghhrso0HW2sKreAwJVlKZ2Z8HvvoOGiISpFOhwlb4UQX7
Z+Sgi9cru/ZPdIKQ/Nl4IYInqNqCGDBXMnhYOpGno3eAMuY5tiJZEEDlPfAo/xRf
UMceJ+pJ9RQcA7fI/CSYuiKhchvGPO5I0e7Wrff8EA/7OMYR/KbgVEPOkwrpok5Z
+37I8L7u0M+szA5hAYq1FWAUH03+bCcBEld1jhLgiVMzhqWybMzCWNmvEO1qNFIG
GsB9kKiAsxT28jbwD+o7Djl1jbIskbe6UJmbO93DcJZRUD3YI8DcB2n/9AXSVtEr
vtvyd6kof5zw2iIrfVdY/3qMZ0XIdDzQbJs6Dzfj41cIcYSJ2m0HwIQJwFYCgqq+
4Tm3wanF/C8YxLII5ad+sZRkflI1TDzUh4oCwh8ftCNL5GeHAHi9d9s8lOL3E8QU
KdC9L/x7YaHX11A0/s9iKwiw78qQx9hsXmfB8Kbu0wj50L6VA+N80AZGnZkA6DKO
d58lUDbtUnbiwnCXEkYsLOPQnSlbFhsphRvRtKDc0CiC3Trc04Tq9kRpYm1Pom07
5AN78LLCdSqmpugABCSGlPoJ97jWSlt6ZuHCNThK5QMYowppHraVghCVqrxY2zjt
rGPmfCDP7VTb2QiPpJASky90XAiZNjWgnmJOaH5BU2/NF9ll/51w9wKvhVWvcPNQ
QHInDiW4LreVrm3Vo3rHR5BowLqyViBctA6HqLVQiO2cojDwBLOl/AKh9MyN1yY2
aoVFqv9CaWFx7XntKqcnfBMOutKAm1Lbe2MOBgbwSwHuK4VkR2O8J95QD2lgNxgI
hfYgNlGOdbjDQ8efgFU9Rk03MAq8AKtl2k7MTwNBLC08nF0y8DGtSHFF3g7pANWS
iB/GKE2JQCjFGGhcEdM+Yk/vWsXf/KesGsnm79XK0BhdrthsY5a69Bv7CHGC5D19
g7uTBfDsvF7KYAIN5JqQqaERVZSN/Fwg7k8Bgp/NTTjE27BD9d1XHmgdnPxuaLBJ
r3qTDj+edC/cT6uEuiNAsZPaQX83QV0O/ikSt2VxDYeN+u158K4PtYJOmk+HgnDJ
kKALVGkIVg+mzBcg54r2e/K7+SMW5x0sAeI5JlombruSfK+jQeYnBahj18Amkyrb
Bv4YYVKH3eFg50ywJiZnUdaI3OVeTpN0tV274tUDIwd3hWZnglB87qbHLUuJtqqs
tkGhDsHKVZyY9cCfO8DbbzJoaQIJOeIyorHOwQSA1L4Z2CSdBYU61ZNO2IhQt+oW
WlG1ss7oPixgw0v/0al4eZk2tSD33b/2ISxt3hnUP5CI7tGK/vd5ttluIXidHpqb
DFor/zTfExTz4uPSx7WeLA7PY104c9BLGqOVPZ+fHGZ+d3i92FDw1nRIR5FI8KEs
klNcIoPJmakIQb+CqzalGVPCJF1GcYf5JvZZRBlGHf+EL7Vc+1qOK5LoZkHeKgDN
FTDGSW4ko3v0PzGed2yjWLL6B2UQrh/54okVIvMkHF4OhoK55NjR1funqlJ68X3z
f6ZlA8qHIaSpDTq45ImnHG6z7kf0+wxAmD7WFdv03Ulf5MbqcxC32zzJoOzHWM/R
eZ6gwje3aqMh3xcwLHcSY8Ta7JdvnVUBcDWORMsmNklzg50C1+zEfOARTmQLP2EV
AUd8ViZKP10Ih79v07JXQB+ZIHA81mbzEuhdn7wM0A6Mv4Z5/lgoVViHGg6k+g6/
y/yyXFE7UszgCSsxoGD+sRABz1529pRhfm8q+uEpDjPnk1PBhv6T4UndXioP4GNW
gcMgRFbIXB+9p3qslFMyrQyCL0IOTtWVLZJcKNuJqYjPAgkOX4QuIHaeKocxJYD9
5c9QB93ALrMaZtUYjdJnlKpCnfqEOsRAsOfuRVmOe4YlSavnpO9yCdy3eO3iAGzN
yHuq0tsE0ABHlf1ZuNtvmso1afrTpZ1MufmZQkZ2trao6hXX260Ri/hg6UNcFvgH
npQv7evJKHDvcVwJ9bVcUJFWjy8NaQpivfnky9sBxFq+uqcqEA7D/P5LulReTxVg
8N6/d2cpUNUvx/rimg6k13igij568C2ijZ6H07bk/9dSgAuey12PImvILkS9ANTK
ekLrsaKSKZZi8rYyWN+x+w7F9PkoQPhdQgpLCRwWLs2i5LezkXm+9LOPXKmO6c3O
THgxcRk7oXPUk5EtghuMJlIRvFLqiTpWHPqnPu9VMA6ywJ7fyQL4SYVaf56ozdmc
oGieRElw30cW0eDsVNOkGKn4lOn8kRz6s1ZheiehmJeNlHBVMnvQZ7zk5nZUDRjp
4tR3cwlFRNZP7MCKN9XHfGYOo9hWCmPRa5urXD6NtWT1L4XT7I3bnvviL215QymO
N12T0JbVogOo/YeiSAy97eJkW3mJO/rN5rgV2fL0QHeIHnjJDS/R56syl6ltoIDB
Nf/Gmi8IM+RIezue+ieAlKUKwidTRODq+Zq46kLf/TGgUjEcVb46qFHAqot/MmkG
jBDZgTi8T+BNnYfTweGKstU+s2uF1uueCkz9dx8jWky4wxuOz2Bw8JcOFNq8cWAi
ElGnPuxIjZ9dRgkGIcVqpWT6rLzzsELpV9yaHpnrOzadH4tHoPS5VPFOkfYaM7mg
rcQGj9IJ77WDw0/yhAoTme7WlBCH9yxLZWHeKdAFOA7V5jAYgMczx74/gEec01sI
UBN6DyqmsiQ9lSxfPtkC5XwZadZ1lGKzFLDB0tEiLdIvlx4B/p49iI1wSITYNYHm
qSwbpIYz4mqwfK4n7SUTDS3LF6FaGvNfQkc372KlMyPmCHUU9TKfjpNGbqsZHAdy
TsXa58yLi9pbxJ4iWAUZ046oflFCr0WnZAcfjPYGcfRBK7tdxfkOWkFYMOi4sQsD
7gouUGnAqYB4OrXuhm1So2WeilWwhek8IseYk3wB4vJVU/Rk3bHtEN7rh5DATljv
qlhXubiayqr/XUD5I9BMmuMlnxql4I97559YbEHR3GrR/QgFj/PyYdZryPFaLGow
zRWqDMKGMr4GbeZCR3qB5kqrx77dd9jTj5gmtuPKdaSyBaz0YYZxpvT8ZuxI8aYC
QwQ2hRa5ugwlqDL7Kzf/qYbi94fTokrVQtg6/74Goy69vpdzTKZ0dq6IRaZ5ZXos
s8kSfPUj6IruT6tdf1UtebK7Ue+9R3nUKlxagY1cwiouq98y9TRQIMuU83QQpuoc
9m7ZQ2uTG89a10L+n5sR6NeT1CqwXUyiVDOtP5+W8GrTls5xBh3+h+lbMRQ7Uh0F
glZeVjeXS4k2VTiD6vBpSyA89IPT1GheF10h2WvIjUU2cSFCtq3d72BidUxPyjr0
dgALdos1nXk6Fuwlj6DWfGvwPsPiVGBV5FA77gNf43vDx8Tji8aFTkbsEr1H5/70
gvq+qcEVcE8QCPwRNTwkOF8pL3b+OFbWOeM87T271u90EqDmeZx57OUIqaXGiKvs
6b5orD78pGbInvuKwNdLyM5JPABE9/01Me5USwsh0sPGQ969aC9FIX1xO0wkt4fd
3oeKjXJmpEoNq5mzLT5EYoa74n3b9D/j1KQl5jfFh4M4z/O3LiZRtHKFAmS60y8v
RjOi7DFxcaQDYktAqorkFiodpBjCnQBDiLJL/CRtStAlQGmpI0jclHWhz8Az0Q1M
APrWgpZnfWWnmpbSb0s64InbTJSnyCwGCZHxp+wh2nyHmsISIdtK6DMlIWIgpt6N
rR6DsgswSGP7vL1JdRKp/UiwZ52d8RLZEUhkZLLc8Hlg92RTZU1pMzPaf1CzHsT9
sAIiZ9NqWrJkl/ax8Mt0E78biYr1+dW7+K8fKaGaxHNeAhWCIlZwf6RJLcj7041q
UsvLEwBMgLO/SQkrUvFE8tbA4x8HJ/ScNocv9BMeR91YTDBu174ekEQFvoheSuVv
/4pFPEazbDzLH1oxqnrM9gNTwfkHiYGs3xc/KovG7BRHqaTqPxEJXu2ikyOZsJdA
CMSi/FAOHHwA2r9JU4I5kAQDOI7Fz2M1wsiVFlPtVa6CMlCzRT7nrypyU+gyI9T3
AIniK0alTlxVwdXuWZuUaPOltpD0iQZ/0oKlridLr3rh6USw2DOI4RjIvBq8vP6g
REmWslGYmKX7SnmmHsjctpFsALefuy/yeZ57ZY00c2ECIxodtKiJ3EaQcP9FoQeI
y6uMB4AuDEsNAQd6yRBKeq3psqmpOoDpQER1Jg2h4JDOhCSJm9oDIqcfVLUPcR7f
dPHscbQSKG4x+S+znNZsWK5Dhvoxz7xLR2ycu6t941M5ME027enXtK0HyvlJlQ4R
bwkB2oktJCVoynvVpIjAUo1+MHrXmkeobMrkni0RKnkHABShZWK6eO3vDtAJMyLZ
m2RjucLnRh8uN5E2g7spUVlqSGYMgru+O53ukfCukjpUujRVgvdpfmLfCB4CCELi
14ZEd5OAK/ym67i2r1KquNRFpv0rCMVQw45ybIipT0hIgNFRU0yh+FeGcEv3Vd/8
RzSZiUq5wJBAw5H6KU/FCAmTDmrRmxHeE8IsQJXDFeEM5Mj13d7lQ/kJeStTn6vD
CiUOTnc1XUcalhr9v8cjiCZ7pRFoHcZP0fCt985BAhvBpbOS4XB5es5XMMpBK5Mp
FYOtcKGz8Mt+CSv4I0f/LUTa8S1ucsCupTAEauUO7ool8upLfCo8dUG1J/mJJQIT
ttsBlMxXRvhPpNpEUnpuYXspGo8NyO+wiaPq5oRLT3H5a0CfjzxjhD1Ek8xKkyfc
nPVuNW98/Arsjbky3i6JdHt4aPjuJqYpjpImv2ajr/ZI/4Pd/n1jkCbeeUAkSYJR
/LaJQLsd6FnLr+MPYN3HIKyrIIXqIuVUg/iU+JWL5yxaPvyvHSu8Ek8UqAMPwI/m
P/axDn3yy2xoi+eMc5NtbED8kyhnpZKUAs41woA/byGRTk4cvyIrxe4J0VmECOoh
aU9FQRcbUk2NcN6TR6aI6RtagH/a8Pw14hSYm46sMYtjpChCefyhMtUnpShUkzO3
X23oQE+VkRS/W+bZzOkvOzbEwub3EH/zAO1p4XcrbEltcEbM/2+5xsWREYCI+D+2
XskUEiIIZgRaZ5IFV+PpHgJbXIRrunn8/S5XGIrj0WElVjJGqQyF+0tmHlCzw27I
+g70XqvrDgNYefbU6GiME7sKhHQqorIQR5AA/L0dtbH7M6kH0yMXJUn/X1PstELG
hLltz2MA5QQKAuKHgZs2AOAU5aPM08WARGJBYUkLUENxZCPD6GRPC/PGRpZEhFS2
/5EufZqhEcCT+TcYL44JGllJfHqy+SrVtZ7WvkK8Tu3OJWsugSdiV7Ryf/XybV6y
YRG2JJqYWvlELbBD24v0nBOSgDgpqFXAqTtahMRHb5Pxy0VBVqEH+5n6vBrvJadO
uEqZor8uKzQk0GdbaP9vRV3/yHuX3KQRT8eHZWVsBp46ccr/inMqODofMzOHvnBw
J3+QhBjIOHn1CIj3V7VDoXQiGOrw1mvrW2g865qnqMuhvkKtRzkl6vmE4wh+SYeA
KisYq/39skKMoYzu3kE5VqVs2EsSBq1LqI64VvqWj6m51U+Hsdqap13I3JzYNFiR
E3oCK6ktSUsSHKrODT8hG1xt2BOxDWbsr3pz2oGlI3u0pL4227rKv1YFKjCOKBgI
28w49YrNbPtVSw7EddVqcf/2PQxf1lOhse5H8mfEAZSZYj4b3zmLq9xT3nQIbEwT
YyVDSO/jDv0DHHiTBliObCb5JDAxPqT8py1vnWwmlZRuz29hqwpFmysOkRwOkuot
FD3TuPBxrId6u/FP0+Hca8Eyoho/2a7cla36/KfpugSVJZj6VL36kd1H3JVSDLb4
y5qADeOcK1r4a+Id1no1z7cvFMfGXaV/KKSHmz1EMVspCY42Udro5jrUfGzvPPf7
aHPbDdOnxz04wA9KGK5JNhkm2+w5VdsLwtJqZSayUG8XidAIjf7VtCOqpfD+L7J1
FBoTuaQapaE57UoiwVS+SlNwYuVQL7J4LD6UvkklJqNHwCvxeHUmmw0bhhtOEDGa
lz0wIigv/jfvdt4vChezAlZs/K8eSdbyg/JNF7uvG+j4CNqx0I64StpCTC4vmlAL
JrcBk7SKkmBziveo/UrgCDhZQVLD+ZhySie59BGBQWTsse+FtAooR3pHK3TkQYoi
SPw2VbjgyvG9MDPAG3Wavpiqnf5r+ifBd2FXbpgSqU2cryQAnUjMuwB4qfCga8Fm
paxUFYZ/xjPAA4gY+tlTsH8c4uwFkPISAxSEPsK1N3lXCjfapWx/82KqlJhNjcmV
CjIVLyts0IaqM2Jt1HUr0W5ynamwYe6BFw3mLtqDrA9rR/mppRS2ZYqnXOHBiMVF
BuehBF39UTorg6xM0nm0t1CSjit3VmHPTOqfno62hFlk2xfmC2UHJqhY+2JilI3a
ZXbCTRl9RaYlY+kWElZhoy8aUXf492wxeMvhPuG73iaL85yOMspO6GH8D/l92LtZ
9zwfPEr5qmDFWN9SFgyohmvCN/A9rBVw3kVnRUD2vjgPk/zfjxzGZfRTg+LrIpBR
mPhnSrKP+ursNM2TUGbcjWB7fMMvqqHaAfkF6WnmLcFpwiGv84oPIQfU5ci+4TfQ
i8pvl9dofaoqVXl4z3bul+n/pW7omSzKiSNxDJfxld4XK3Vv4R1eYClc8hEt9t9n
pY/mQzNkjFn0zQGKXjHUnsJQyFbxMELCDlznB9R2LNupwQXHXP2IZgIy7H3CSuk0
fNYuPkRx2PlSs0cZCG1eUZJexC9sknt4ZZwv8IbNZi0wvLlXARuxO+FCW8rJO6eo
4rGJwgJtDpVMutNfonv6SVSAbILsRuQDqXfg+0GR3obqjZw7Dxi48VmznrBzEWy4
W63hB/ffZlPZhSKq8/rZtkO9yIAYYQxCBqWiLDEz/ohY5fzMLNwVo8u7+Z/2CQhC
socpy/o1v1y74trSjRrsdjCD8dTan1bJ+crIcIgPtcySK3lOYMb4pEUB+eUW/CTt
1AWx+1/eZOPnQmFPMKISAe3lt0whG4E1H8EcEOyQPF4YzRPPOQcGqPK6L8X/gcIZ
V2akaIjtLoqGCxolMIJHcKroQ0/T3Qbb6h/guja0M19Lkbdj+k0h7cIjzJng0dA0
1YdVmxUoDZC1kWOWmdPw0AtDn7RIpeIzaBQ6zq9m4YSmiCX1hAeN08CqIRNZ29Ir
C7wvbtn5nQM4PWcgH0PtqxSyR9KP3yqDQuTsCxQGon8pxgdnTUKDBbJGGX021dqJ
jLELdd1LsQ7mVsnyTtfu8eIn1vZcd+D7VD4WjTiYRZjw7dybORFGQoKY9Oa2dAgc
fKYgINSO5Bgi070pLT8wufPXH8NoFPGGdlfDhHbddv7I53sJbx8hxNOSIX5sn7+8
ghJXhB5JkXz4xrWxdmpkYXeOoFWoJ83/qKdWHTACbt8nTbIAWRreCbZhHKs8rjhK
bkPJBdUYkRFAhiTLqy4lVcGDNlXuhFl2tErDNhSHa22HWL0w0Ki6klDbr1Qp1jlw
nkLZTICRAv6+cT0QEQ9DE6PemQ/GCa1sVO1WdLVKzfqzJmEYJBWikCu/B71ko8rz
3EX4JJs33R8ToYzRNyYAvy1eZGy7U1VeMwGhwSlnR2ApJ96Lr1U1oROQtR/Wv+2E
U2aknWhufOsrNbQqgef7o4/IYPuydO8T6b0hxwXvVM/8kBbfkxeTmqyO2xYggAAO
eJAX2mR2tVA12QDiSDdBnYyArrfZHQ4/ci8OrpY8urHc0WCLPkLA0BBoFMnRbaLY
bvXmtVV+X1ZOQ8HDo7cZ0SBMckw6QyHUkJ0plxjGQY8T1JpqFYyeVoCopgoPlb4m
IdncZ8rflBZlc7dn+UVUy/jacTrsDJlC3cMSA8ACsMSDQePxhfen8srePh2324tJ
yOE7QvNNkukyfRlvL3haCqvuBxZ+8Vpxh4vPvQuCS35kfZl3gPbOJFZWgT3SfFQN
fAnQ64nKA8+EOAanaqgPIFXwtaO1yi13NFUtb7Csu9yYlsp2N2ZBJhoflbpJ5pOQ
Aoi0yXDPdJfutxxJ5y+/A6PX0GJ1MviYFjKyx8UgZM2xJ8GHuR3ZOFCxu1xMlkWc
JLPt1nfMVCGWanDmG1bILbuXMhyQk+CBh35C1o9yHI2fd+Ir5R/7zreBluyNGJ9D
JjFWjmLYXEabAJOEIszK8X1X5hJ1Sr4GNfMxlwl7u5QnhX8UY13QSRJnwcLlvnrf
wNERnSZLB+VS+t+LkVkujIeRGO6U3T7+lxfJs8sp0M2AmTJB4BzTtyY/M8Hc+lYx
E2NyDM1C8VEuqj81oM1TwjzS5U93y5tKdNm8BmTJyuT4r/1Bs7bqFhnrr2i/IMqJ
lMG6nBsZzo3S5Ll5Hu/cHCmQNrcgpon3t55O9q1hcd8e/VCrk9pJku6klymvTesO
uU3slU7CQ1aJNMS25dqIs+fNQQ6Y+mubkXzutTL3w814uAt7hlKWwC9TrudOML0y
GtFeu5+tJzGz+IaWA/wRE+zb3kDB345LsCXwtpCNsXhRNFceoBK3BnemBTYOcwIq
m/QkgBebdRtXT6YFu7Pc2EX01aS8QOjwHEF6bwFawdeHNe0vaFSunFYAGcCnEA7w
`protect END_PROTECTED
