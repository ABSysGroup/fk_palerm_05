`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kwcvr3/OB4kfbCHWzIpbxQH9eGhSGiAn6Y/ufXnnEBR1yI0Yh9/RxZY6qWKr8iCn
f1e3t1bPXlSAWR+kE3hsRf/ohCfJSTttrHqV4zTYew5v1+ngcS029vGC6Id3f3NK
bzS6hmKESySDjE+HVV/Fr6Lp9R1teVMQo6nZRsLvDR+3rTJUXcHAQV50p24qhcXr
ns8f3rUHjwJzWOO4qQIWYq1EwncLNS6hsDmbw6+z6zjn6mgmbjP3+DQbZFqEgMho
Ii8vnWLJaDD6g17kNCbNArp5u4N7D9VcH/IAuc5QJgfZpTT11pmoA2+X5zepKXea
H2SBbAlpkd0AuOELkLUntKVcY0NIFmeRGE9VMfstX/Q=
`protect END_PROTECTED
