`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xWVpcHLBHXKA+rmZ+c09wCpluI7ex44wUmE1mkCVK89H09jYzzEkw+xNZ7rUIxJi
CVzS0Vp+DOlMbSz1JQm4VAVpmEMFTx/3LjQQq/0+O5W2XH1BDQC/f6ZHN7WW7bXR
GLvM81jsoXuv24qGLRx62EMRVwtqhzPzUnIuDFLR04zaBi5weBdJ/W5BBVVdDkID
1tMvqDUsbGqOk/Ehi+dsB7pkKaN8O2DQe7An22T88BSFSoAuQhHNzfyG0zQisX4e
hBJix5wHwSlSrP7Tn3Pamx9qq7DYL93KDO4Wh1BL60ucgwP3eadRZjWOobVBYNB7
II2Ko5cgRgjyImCpFrrbUTdppQpWvayG3Q5qFFd6vCZ7QtprBMVqEzdbAy1w7eKw
sF1tJb335w08KhdGWSdZXp28cO/IH3N2ky9SOrhDxbDRhMIqFPTD9gDax0A2ms0k
hzSjmAXO0Pp/+ghqEBPcPMpzwWpDXs7AH7TNWdzBCFRahwYv51uL5uemSFcsR2OA
Bge6ZV4nC8/c2uyCcMGDNyvYwUiqj5lBrbUqxG9Arj3xp811TTOlrib84axhdaHo
SVSwx4BnvMEFonkmR/IDjfJjGDvoe4ax2HZwJ2QVGLOlHPgKuUn2xNlXo93YxcPX
a1Ubu+zPlrmFPkU+svpdQzZnXjTylqntxGIRfIMJVMNcbRH7BXSF2fMBIvkdu3IB
belWkKyzZFAolg4ZSSv9GwdSIg75jJbWAXqfzwrbPRuruaoi72iK9WF6vCOAUkJx
egtINYg9e3QMlxERqJIpkT2Yk6qLe9Ndf7uDeJMUUf6cTKSOMMps5te2qGPqn7qa
pPo80akQDRXi42B9se28vf6uJt7+r1HuXjg6fqtpbH50Bm1DYbNhW47loRHto7Sf
eVq4fSrOJ/UiHesNDBKPck+MVS42JfMO0F86Nl3XDugJ4IqEb1R13y8+JhXoYtFF
BPkMuaaysjy/1Utj9tKl7A==
`protect END_PROTECTED
