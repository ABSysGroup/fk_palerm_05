`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UASdBoSS4VCos0TmjNGGua9xgtf1nuxfTrP9aBqR8FIPs7L25FRzNKgb81odwfpV
liQumfP51sboIWoD6Y+Fj4plbl4t/OUOsYrDS5do9qlnyQfEznZdOsH21//Adwlh
RTg/azY5ImV5B4EX6LtvRjYmBdvdVa60M00odqtqyzzOiH0eVDPXODc0/G0IgQlu
T2BwL2Mc/C/iKRASYt4MyjlQBBZgvKXy0xyUwpZPkxElFuP0rK1NofmNHpLKKQjv
PW/k+AyUlNHniGsCD2rWtFu2KCqUIQKVHBHxpxjgwubNaWmJGoOwQuD+pKSr/RQL
c0E0P9ecNNzkgHd6KWjMBQ==
`protect END_PROTECTED
