`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vHZQ65vGr3mBEQ6BhmdINbp4RAqcQvYee/kqnaZV91M6AJks9RkUgqWV+cfbGSNx
EVUvCfPWP5UOimgqr8pFcF3sovLiFBejw1/sYz1P+64Mk3d5irI76t/1PBErFB5j
rRXje/x1gqgQDC1VMaqtk5K4mma+t5JpE2LkFeOVALjsdVE5XoAkHh1URZOD9oen
gxkAm6AKaa9H1Gu42AwLOYGK5jM3WPcpSHytPyE5rfvJMu3ZvGIWkX+UEYbjL+Sc
Dw71nQUpwW+7sCxlnh9abrwTZdpPk5WrNRMBdcUchGAFIj1XaH9VwczqLVumd9/t
1yo98krluof+bOauDHCH0Q==
`protect END_PROTECTED
