`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AncvJE17EIAed/djyy+iHYIOxSd6UzVYQn6v4AWzq4AfwZuFEuk3MvUn/+RhVGY6
ovV2JFgkBvYfFu89EiOr7YpxKQniw+ZdTnsc6j+0UJcDZxkXqt2uSrCKCDUQ7g7A
yGCbdhR4d8bxZ7vR7r8iic3Tz1hFZaCCEu/hUnemL4Qtbm4qoFgrzZ+8ADf8gSci
oXyRhfH9bU4WST95BSMqJC+jQTyK1u+CAnfJAL8tw+0RYgrHZXLKQyBffarwWdIZ
QF5ANBN+C1ONGGTVx7QHgzQYjHQwxgIPZQsB6zb+W1elEEwc5tvzL+VkyTfYWZxI
Gj984ZYPOZYHsFS2aAG5EsAEfxGFEyV5BKVLaWAtoUZCrOg2yWb8O1ggeyrJYaAo
zPi2Eu0KSXXU5/d2bPTdT4ghA/JBtJFOY3AR3yfEV41TIuwD6PFsVKuNLaul35X0
MqD7//aSqBGX/9W3rhMOsRCVKKeU3116WZXXHqL+ESKV0ewyron0A++XyBZS/+jH
WCuAr0n1GjXCJKA0njFt+0EAwNYese9ZJol06VNW9Zqj9c0px1F1wST095gXfDAq
KY8/Zm81iVuSXQ9z6SKBiDyHnytNh7zWqpb9VfXooZZrmjzcob0lRRVbNsKARcxB
dy/dcgzKXAgiFfSnlpGZxfei9y1hmbdbusuHd3AfyE5LuVPqQvJiS6QiJoRJkxfQ
sZMV9Grtgc3Elb5WpG4dZw6/t98DILSQlDFoHkItS0KUH6NGDqI8E/RlKpKqyuDT
lTNQ0OsD5SEmki/EvBIS1EasKJrfwJjODsHcysJRl8kVmzwOwm5SOdw1JXvBQ7o4
3N6j6ZQvSpk2G+ykKdDp8NFDxbd/P6KtyaGteZkQgaSQ0ab7JLCMx0HXYAuFOhT6
Zj3WDYfCoT+h9636d4Rya5W95WT+0q3I4uy5IMEIByg+wcXnUOMa81D1tRqRetMU
7iUI/FWKmAXAmCHIZqzv6oWD2eYuruVeBs5Wh3VrlO6XsJTGLnYdbNmIN9xbqm/n
AP9P1RkxcK1uWXZCJ9oCFld2ryYPyUGn6VdOAS9jMkcTArfa5Xha1I0UO52ux5RO
qBgCYm2rQcvrBVo+WNgP4GjAdZpXwjF+XDYedtzIh5i1TzCQTmsyGXelFGtLVK8c
+3Ps9hRhv/FFwE22w2aiokj7IvuYWrMNCw38IQmaFgiFcLHW3OPEFgUoGdo9LcYH
z0pjCwTGcqxwBiynGfmQX82z9v3ucMWmIgrYsFErvFaXi3A5l7mtpJVklLxaYQiC
ShEEY0OMG2rdnvfXNWIKE419cyCowxqpHde1oZAX2UMFZflBGQ6GUthKhkR29IY9
iwd1g76McRPRZmzOk/PKTcdRo6ROcwQ8JPkbupaq+nyxdDzBTPtH45v/GI4OBOXs
Ir2oGkigHT2KOF3aZIhqXsLXuDnhQmWSLxpfcVVAIg8ulrXJXqb1+I6nOQpaXsbu
sR43ae+f81Ez7NzfOInHkB4Nr+UqH5nAGjSV5ThNsfOIu+wJtJxQsEflbhjBVkA5
kFGYz4NARsliMQuIW5/xqk4J6Oj2QyAvzn9+WQhSbOGbl214oF2cz3yHteXllwNl
SgWAZEmBrjfLTxtarwaJ1Aa9GGCfReLm+dcZvq5Y5rMF8oeXLefiimLUOK0CTwa+
lLaJ5c2gdDN/8PMnSXqNok2wA4F7krCBU53wPdrBgWTsrCor1Re4xsXgBY4ml7xv
vS9lUWYeG3fFRaIGPkdSh+tckwoEm36daO3+XC0eQ3y+TQ/qm/TILtKi9Bupf6aD
a0GVGyoOI0htu93OxFB1Xxc3Lkg33V2pg2Y1ZLAA3kpzx9ddA4qXKplNLkft4xKx
pUhay7Jnu2WAkjCV89i4V5OvtuzRt342HleT29LDJvp99sZlWEIDWY48rshcs3oi
RLRS1yUyarcHiOOqWbQunL2sUsXjqK3X1n0zYzLFwqH49WTOJY0FRmUCM5RpDdF3
CLClCJz16hdpugookb7LWybQFxzHEBI5ak+Lmk89bglsZYEtlWCbL+vL1MwhroaP
4eSB2OADKCitRu4FWnm+P0dkaJbAyaJF6Hs/UACXeLuegy6ISo91fwituhF7d679
KG8hyk4gzULUH7fx4Y4mq5xYF8MwJrBk6cBDyqSi90o7skjdVYEiRJcI/tmdVQYz
RKk20JX2TH+IPPrXzH8vgWw1txBK5YARS15rdGIZYaSrrJvwQQuOdYUPaLMBtAfI
imXbgnV5AevR4Ypvdjt6wh4c0w2Q0LVaD4giCPxg7Nbq+BvJcZoMH2MKXg6jaPSl
eZKl/uigJhbgiKpU1qTFg8aJMRUy5L9FPxQ2X6/QXb0yKhuQykxZVwickKSE1mhn
VKMo4gw+xT7YWJbrOOAKaNeKH5dfBaqMXs0pEVp77csdUlPKZ+cHsrYK8Ajicr/1
P8nyzvxZ5lnGLHFLWId0TrkAshSXvqdj7DwlQtSMKn4EJ249IbUKnmL+ACuACuet
L4n9+61wrY1VJT3dQC0OCecCjjqZ0m/HrcP9rl4gLRo=
`protect END_PROTECTED
