`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+VaKJtP7nFHE2FSK6la6jh37uSyxukDon2t5F7LWRaj82v+jrVyxdCV8nRQJk1er
pbQqdysOwaVSbA6FN/CPQaz/3TSQfiKoOYhlfO2YYiXq3t5J5giivwklw5ET37p/
SuoJ4zQ0G5ON4D/8F/YyReFdxlENojVONYiUozxMbwsaOcoi/5DTpgP4L4gHF6AY
rqrpC9XRpnCRETwjTETxpSRGz3GtM2QVg11vgMMJLdxSxD5JBvXFKeEXzweOux4a
vGqERlZdHPbv4cmAR3L0N5GtpV67HBm78Pa1vPOKW3oTaZR4bDZDS6htj/6Sggm3
YPLXAyTl5cE7LyUoZz1yYM/SJ6ZVVp8AlPDNoeEqk+cYpUly2trK1jELMGyPosih
dWPSprsUjBk2NKNcnh927IX67VRkgLh0i4B13Zs8qj4IPXqTtroL8Jr4zrv/7IHE
gy7IjE+qAimyRjpo7pIk1QgwYq/MHODkUKOxXRIqrnf3oUxcQYrHyk6iHdD3wxTo
8GeJVwF/vULb8IlMLXLb1E9M2oLIv99uy6uieW72p3mrcu+t98Pcw31+WPxIyw3f
izBUWJomzfSgTxtO5eO97c07ejExQEJ58r9Yc101OAgx4C/GOeRAW6kmP98FjRfJ
xJbfmvlgdnNyC1dLjDxeVkluSmEiDCzlK20o0NK1QJZ+XH2pj8UI4hyp6UDEgaKA
tnn+PdXlYKGAUGBgHo52qd+kISbW0DIC7SSmS5qXrYOJz1f5PfnNwwkV7gjpobbQ
l0eBouu7qTXrF5bGQrExMg==
`protect END_PROTECTED
