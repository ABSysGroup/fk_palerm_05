`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oghfwpa6cqWiOiogwK4OJl75d1Nl2aW+WIK2LgrOEQ+AQXIi7152qY7RXxu/BpjF
6tmpfCoFXmV32PQkTtDHNAyxM4tWHJYHJ9nuZbwsE3WkKqQxFKtGOKKZVnYBr5bW
osKYS+aOH47H1ouhBuQubxS7siS4lQcbXTz/xVPEP4zw9W97hYln1PmrjrdRporN
nMm+dZrN4HbzRAfnRBcbjFrH+wIYfHZMJEBa4S/pj4QE1NvBrSN18z8J1X2N7PKr
l7RWAP+XcxCcztf96nlpFMbuV40PfyUL7iROh/Bd3QLJNtumvACBTkaAN8nQQk3B
3GPPQHOG9hwdoyFDoYfp7w==
`protect END_PROTECTED
