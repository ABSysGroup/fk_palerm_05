`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LJrI4IMFvEhUtrSi+/4DB5ez1unxgXbzYTJl3oD6PxNRDkNtsKKXtyvS0mx+Oalf
orsuDIjAaEYCaYlllbab3rP91I2fyUqPxq4pJ5SEqWafRULnNQbgmKf4khLt9KTd
BXZlj9Xx6un7PUMokZLIUUTtUqY2PZgh9dKa1nSIoyY+9gNmtw3l/hFNmod5XDBH
m09d1HvkUk8nYoMHwlZsIQO2wUjKEKWOPPbrB1JbzvmbwAscIzXfMDMmDGOKefDN
lxEVMbvP9IeQKoj7F4dQ8yMBIuJlLYK9NUbLh/+TGeeLmn5i8NoX2bwhOg3uPWDt
sHE+l15gleYmENL+9bAOyILdt5r+poz28GS/UAmq57OI3CVeaAKS5X/57wjR5Iah
K073BGJPSHnG2fgTE/m8lk7Dqd5BWjuxWIuoThq+qBjoHA7CuQcZSPUynFpTVLsQ
qhM6ttj5b5Uw2fsLdl5uksWZl7vzRXX+i8LvPhLmH061hFy4riPvLvZKQKu4Yvok
ct46ptMidSdM8BCEyeHGkHmWGB4S6FzPZtg4ThXsruROqJKa1ZunZhJRv/NpDkWb
cwUc9GbIdmkojlCnkZZI8qPbM3K+W3uT1KPBxXJGZbkR9D2Z9KhZbC13675CTFEG
EopfD8TaZfZiidev//GxL/mYHdB22s/5nK+96O8a0+AjWW/egFM6xOwmEDnu8GrK
H+4ptuwuzlRhEAylBToBceAQ37IVuGHo+nFOsa4DLpK7xZX/Td8ZBUJ9UzgLuLbW
PoftbJt/U8yJBO5abmyXwtTAGGl2LB7uI8+0oJtEHIiJWu44Ochj+c8i7pcuEzSy
sPLhvbaKwv7Yr5j9ZXY+Prgi4bPzjce50Rc2BuQzKbbkP7fpTALjcYG7Bz9QeNMA
uShzldvO7jNyTaNLlvJmmk+n0uE8qQB8Mlmlrk6RJc15iNpeuFx4sxGsTT7Xyixo
Hbd6LaTCjhElz1b0GCv97JBe8yjWGkW9ng+2hTeTjl00K4Zdn/cMmRHIr/vCRKlQ
qcYCXXSFK3Fo0Pj2YcHFbxc+x17X7niHkJVM7YfsT4/t4/IObLbF+VZJkRrGEjLF
uM5qu621LmJMFU403yvXFXHL1W+I6gcqkVc4lkaPkxHJ77gKw/TSBaYD/oRvNlhR
IBolX4wmcAxgf3aGl4jUJCE3Xdmm5bzPz41SCA0PccbZuxFs8IYF4mHBVUGkorVO
EKyZaGk3NeCvhBrUnmQ65m69f833XddtzR8dM/mRhZ3AC63nFjyVGBt9exj7xhcB
T+cqrRDo261VKZfxiCsEFA==
`protect END_PROTECTED
