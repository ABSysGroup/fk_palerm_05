`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8NV6qELSbqdLw74DBG1cp5iDEM+3Zm2F1yJcQdFfe2IRfAdME7g9XSXh8Se2DejM
g/aF+XzOZZNFLrXlcdN9UfFc50FrDbiub54feHijJS2FiU7+kEvZ4Buz62YfX7VK
+B7eBJz6jEEc5hsg6TcuSB2sy9X3j9r3mwCr6pRK7lz6pn9E2D/bG9U12/BHF2DF
fMqXMNDY2oPpUd8+83x60vl+J2Xjyw/KbeEmCwEbDc2B21HtA6AbIbnGAYKC1eUN
l6kpPrjlDBQUYUg9ahY+VE1Hw8JNVaCbTKGUhLtiA/vN+ZyI8Xi680aae75YocLg
0zD53hl3cYLf3X6onqQIsKvOncljIP1xSWrE0xkhezAvofDE6q+n3Aas/s5VgfVw
tI30LXi5FxGBEugDu5qgLAO2PtkAzIIOaXDYqiw5rA95ZPlAkqI2nl3yo9FNC4gd
nTaE13895nypGzOsRl6ZYKND/R9vxt87a5GneXDBMp8=
`protect END_PROTECTED
