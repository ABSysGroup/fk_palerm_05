`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g100WEUs5vj+m6mcMdWMFj80G/LxuHXHDvTM1jtw3jOR9/TL0nxsy7Wix0XEpPXi
9+6JNNXohKWz9uU/Nvx2/m/SDDEaVU9I9tcFrSpIrMJTlABTtYicOxw661JvDjnB
DMA/cV1RYWdsgL0mKmZocidRKno8Th5M/hIrJ1uYRgGL/gaxQqAClc+s0obx1Z93
dHzy+5z2puWJ+ugsCz+Sy7cYdKy4GeeeVDqls1E2+JZ7dZPIjceRUccdT4Vpma+e
P1RFSCtOdQG6o0AfhOMmDRlXLg7n108/mSZMOHxXO0wtlld1mISKRe+zabdVI83Q
0uQ1uhFFBNC/XnbbaOZ6+TaZV3+37Fyp7361SUsKnhSkPycUTDMk4/CZRm5MAWnZ
zl6B/b2ATJlWFuVsu9jKDH97nCdRfwBsgORnE8TW3RMvyZ3+m7fzsDg9oJUMsx5D
djZJzDV2er9tGKt0TzZm7tF+RDn6kFt0lghidpmDA/0jEdUQUS76CriirnaHYBAK
VgbQ6QmNzvsq8EZOcPRoxYr7pQHt1UAs18qq5m8qPjGzvTMRKefcFM62LXJgSjvn
YJAXb4Kei5xJIiUOJ5ZcED8aVcWteS0NqyEC0GA2XoAQxarlhvCflr9I3P7xwXoq
B8ENIyGkeI4dLELS+vzhrCTFsfPJ7OHgWt8S3DT5HfOUSgACo/TxbhGYDV3Hh01x
N2FFqWh05STbuCu/JLbVnJvE2fbiLv7p2U1ETwOWwDI3M1H9IgI91JxBJfa2jMtL
kYPAE3yJHYeIDtFFeRXEzCPezSgJu9RDT+q7TbqzPLOpWWR0gTxT/4znT3hb/Itv
TmUFgBrSr8mZbWL8liQP5/g+toakR1t8bz60P233vN8SERaXQ8JQAB0+7K66CqLp
ap/kWg+0WPh4SuvnJiMoWNEFgER1Vj+TrgJtvortNFwxJmxeWQ1HOPVnDIkOYTP0
QJpjAnQg0sT2C2o3ExjufV7/d2B3pNKroE61tMe8tjR1GuFfHyzXSRWGuyziZNvk
P/7S7ct2qwAn1QZ+U0c4JDiSJqipxxtwbXC+wIehOBe9g2vf72TSm0CHKF+ZgVym
111XJH18R1iRby89kFINNeheQfH7XrarORScjQs4Aue6ly5WuFQW5HpBX5NTV5l5
FrjbeLNJ5wMkWCSvqKKtJI1nQxnvHYd7IbEB4McnQEXhRQU4aRdHHjr7/mldsp+G
OetHZ8SnTZa/WY7N5SUtr7A07VL0XWcDSOPP23x3Uck=
`protect END_PROTECTED
