`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sW/qfB14/76+kTQa/8v9g/9AP/yrvOA1ae1p9GyPAPm4hCNng5xA2rmZpwhJh5VF
qtAs4Vot9Tis7jwIYJn+JctB/WAcRbIbhqxV7mqiIi9n0MKAFLKpeTYWt/ccUz34
c8lATASbZJidfQTAsAUEn3RjJ7S8DNRpktjzQpGCFDtDOOrZHkeqQUwtexd1XT5P
NiYObCbxxzaZrGZB3Lms1XM0jYccaKnNZ+FNmS0cVxZNzOcx/1RACIzJkLsKFQfd
V1wavlWcspHnlHZUWPzycvmLOaM+kL03KYWo125lJkoeLcbYUGgAFW67J6tNENIn
pio2Q19HjevlLdFms1dD0zJV8A1gpIzUl409iOKA/ok3QI4d0J9yG86htCiToGDQ
ea44H+9C4FivYjFT4YBv40mFNCrCFQ38o43dk8ya1QWi78SgNnmdN9+x3r9HDcg5
6LbYWvn1gIhKnpUV5xFtfLcciJxoB8s4A8zevWQwAzDfMjIn7f+eAJ/Q/6miaOhF
1jhhkKGxhT1AqSx2zIu/vQ==
`protect END_PROTECTED
