`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DgasD8Jc+sHYd9pyxCMWTKtVQoLo9wKg7IGkj9QAQxWmD8/f6C2p2hMS/B9BYoi1
30cBGFwbgvFo1EDsh0VG1+0M0nPPOT6uCYSMPjNaRi2CPd1sWjZ+INQEh9QLfBH4
5eafGazJmb7Fhme39ajVgOd38gvMi6U01yVA/rpRA4SItg97vRoVEBO/2f2JuT8r
V+jx1f1fHSuaj/N7qEA0KZVNU8xvK1ZyM9G58ENJOHOOqSqfbwkx8XUIJURwNItd
yAEHerGoyll2LdwIS0IpUs5yaoCZsqIrjuLD8rq2dvu/2hKcrGPoI58YaHR20Bzj
7UVEGlU58jUo7VhGgyXlGlkSWwuW8suyDdua+Z7OoSTh2AQ92jkRWTRFYW+R1lqR
QttmfYvC43qJLCP8eBt8p/3CU/scVi485hR/ahKFfaft+SrBzyVAE0rpuFHDa3jD
8MC72QYRWGAPm7sWE/FwqScfjtnYJT5CduBU6t54aYuQ0yJ0GAJZkkMwXkBTWz/3
WPp5SOJBcHziE8yLFBLAChw1wWxGS7vkc3xHIpsHqb285yjzBNjn9Vb+t1ITxdRZ
mGiB8G+Xz7ORIS/k4B17rv5B1DGxK2e0iT/7Au+jaddjfdXimOvTW6BEwEHOun/I
qrB5YS5d9YQL4PI0Mg/AVV92QMGu6jwDURb/v/BXy/2ALqxPhcoOvbg7lrg4+Efs
FVtnh74Sl6gfhicCcTxFYxHajUCmzIaGlD74hFiKJehhaV1RVLdYujAGZIcfGWNn
0h2TvhWuzbM3skCmV1KQg+oddBhYgv4EeqSLW7PxzHFcDOvUiJ0TCGOnHcP6Hb+4
pm0gPcCtgsEe/Y+KOxQdgsgs+uGv/Z53VJY27vzLQL2iV3gXjwsdDglpA8qLeF6r
`protect END_PROTECTED
