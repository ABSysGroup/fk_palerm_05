`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q/FTO8Sjg6gVgLEsS5gJUhvDR0Xo/D1hp8UWCKeGXTHQ99/4zyW73na+iBfxDoYH
09wXp0wijofV5mjfiQ/p3SxZt7/CnbZOwSKYhIEw3XwZkE0oRs3UwkVDsXW6WVV9
4SIh5r7rNJj+rKOZ7Q/VL00lx0n/+bd0xWPalAzh3YQzwOrZQ5H4cuArKTuslVWr
S95mReIQK8mdCTXp4lQ48lhPrABuqudw3HMlyVdp5+3dST+JJOko5i0whjjtTfWw
NijgM7x/Z7Wcmwew7i5VjbEI9PUsibPLMkEC+1Lz4Yb6E/RdeG6CDAYOrjaPFeCw
8BYdXnr5YHyic+O4lnzXWz5tHONN1ptRVF+s13JTLXj101/X4SGYnK1bX57kZ1n0
Oz+iK14S46s+2/3lfMhS6EVKwNqskOfMNO14Vfz5E1Hef8u0ystHT6I4+TmAO1RO
nFL0dl+6PGOhZFlhX0XtkB/k/LcT4AD0Ax0SPKpiRAvGy3ZtwI7j41fpy3IGp7JR
Vq36AmMg4F84YhuCRWko4dOTO0okBR4lt7prqvneAWJGhoR5bFdLKjhE3yCjNtrm
0qCnJ6vvDqdsb1XyoclccgvPye4gaULzDz4EzHTBA9WweXQtmIBbhgm/XtUQy7E1
d2fPRF84DOZtldqnLwIiwSWwTvLSCXGGGvCzXD1P6+vQ7SIXwNE4oa3Ct4JhP855
jooaWEpkfYWvqa5X4peOLMb8BmMNgiirK7qUaPBASR91abmmCE7TiNNNAjgnDR2t
c4aPuLQLnmKYkb5cSBi5A93xjYkGwM3yVVFy+mWp1vhueLftRdme/i1k2dTiiGTJ
jwQx7BFOu8Me3Xe+wStY6+iYb4/sqkCx6oqVnsFX7YyOIZlBKiWVq++vlDxRec3x
q35HdsxmYdIcJih2XIyDlMWrooNiOC3prUokngqcg1JULXCyEifabAHZTZGQVTyl
u+0DnlaRK8Rt9a5IMSHlknsA5aXDZQOAUm0z8sNrgNH6VXBIEWRNVukwVeRsA/5b
MHWuNjXtlSEhgKONJ041e5nSsvaFwhAP2NlvLjm4M3ZxSpfutxgwhnb4yJebxyz+
AEwxjUDbxGQ2ws9g4fXAzw==
`protect END_PROTECTED
