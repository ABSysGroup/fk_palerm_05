`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GvAGmpmysIUbTQzXRlLLDVmMZ7lwy6iB4PHGX9POymXp/Ue2nNbdbzTmOYDhhzvC
P/Q8oYINncm8fESvxC91EuVKoPDFnYVQEqwUpLD2cBwjmBBC+GihAoAUGXnXf9B+
lqI2H48DzGN5+etVP47ZP4hkZbi5h5vGg6uHBH9FVvffwvmEjxfkh3KXpEO0gc99
XebZwjrt6yV+MJh/lIW0z0CScWyC5d2kNjDtDA1cYPWI0uumfYNHwIPM165DIMPf
fZV0fSn/GIBmEqAUNPyoLUuNhiG7zxb5XbN9V8GT5XkeJNkkgq3uBYwAVgOg0CK3
HeeozGF5vI7JPtUHoldJeclLOtppQSSBDhLNKetwiU+zdYDHVd0NyOtzsil8TkcE
zORWIohwohA1gBz3seVrk9uF9kztZS99XNhjecw3dy45TLKgo9mP9NB6cjoZQLfg
Ck78EGpzobn20sB9gKvJlsIU20OuqZGmOggpOSbBiIQpWnPbt5/uG83RTM9QLRFe
0kiPgf6Mqd+X3udBsMiZ41/CTTJuOP1/7zC+4PP9GUfu1Wc8IQcp2sGpJtZXOyqQ
MSQgHA2a45VSsznwNUOtWEpyW2SSCECehDA+FQUyYdNKCTDRNBjQqLKFF3wxv41P
pmcSzO6wSyftAG4H1kNJcfOFmJ1b2iL3V60RbtR4vVjrZ7tMcxvBxVTRdBYgpF/x
Y5oG9M3Fa7egrTHw5zmRPaUJ/Yr+3Oob8KYXIM5cs8OBbjo9egvFMUxoeAxiwezZ
M+MQikO4m4cNpdM/ZmkmSFjuRZLWi3pNs4cIe1mBvDyRqLm7BW/EA+OkKduQ1IQU
ydioLelwgadTFKmroNUJdrmEyhnJyfw55gXuCTv9xd072hX+3O3s6obLI7h8f6jC
DoEsPNMY4AHzSuuEaQcK9ZczW17Lwf2FsQ7kfOLvhgbuLhvz+SlDIzsydQmjZi9K
k8Lp+egniryQgGBwUk3VVJSdeIPbnRk/V5HMaE/C1LSpWUIoRYqyNnQCohtxxr6l
nsvpEbrZSjMfswQ8qjcl33SUBvHdf3kS0w1WLyJXRHcsgrT81ZqhijAjBS8Wmx0h
zT+zc0q285QqJAPVkgSzR8U/omNh5la2Rz/tYgRYgJEVnDfvShX168tDZ1SHy0Sw
RQv5PyZ4+j3qExnT96p2RHQGTk/iJI38wFL1PNQwhMxo7W3ZuYBT9QEuCl2dPEiu
EZUBDCMLdacA88VXcejewBvDSDtYgigKJXvMOdMfRYckVHSNcOG4rORrJqrlGnV3
yQ9LIFkw0O2kR1FgFp5cTXGQHNHnOd1WMeCve3OGBY1BxMj9QXANS2KRxE6N//tR
o3N0glNB3hlbKGQQDYMDm6ALGtkeq6k7o9V9HDEDWy8hUgWMOno1mVZO+gpPaEoU
EAmDi4ZXvN7PuSQeNxTnRChk0uXAH/xEankZKHpUIOP5Tv6UNEq7c0Yo1kQaBh8V
6RtgM7b0oT1MuUzpUNWmBSsmBFR8prf+riUsryvikU5rC2PtJvzazaMMuHpKnOlE
L9r2mAipWjoI/Oreuco5GXx0bV14bckGKNy8qO+hqIMreeAmlhrcYNqTrktmQEga
qy1tC4khAtdZMRuQXTlQlpmpkMhnTDuFdnhkLT2YSjR0K5SdTqDbeYd65nWsdHbJ
2Cg49YlRrYtxHxW+LlXq+MRBihWqT8UxyMjq0121NoL/eBt7/pKMEIcNAbNSQB99
c9oEDGJuuUdfZNmNRf8/08e7+cdd4GM6Cc/o25jeZU2HdV/okhh7uvTK8nUIeT6c
iFTaV/BacevB056vqBaLaZ5DqX2L1LHoYPuuB9N4FFmhFJyGeUzWQWd4b9zY0cri
`protect END_PROTECTED
