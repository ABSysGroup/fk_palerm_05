`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/mXrN4SDcIefOfOM1VKpCj/qgZjc2rKwW3/P98r2v8ZAtAj608iose/r5lfMUCxc
1FZo3+XZJoyURjahiMrMIgKXkj1n6/sEWR88AE6sfBEQdRXJt8hLYW0qJZ322Y79
gtntYjluab4gNJdXiAvSlgFjteN2qORWmWzAuGNGl1G9oydMkkdlWOJiNicd1Z29
MhzIE47wqDGPEbPzXcBkNkZhCOn6xGP9R3qHhlzL6eaHPOjF+tctcmKXVbgeIKha
B7AHhb7V4u62YmB8wQ9d7s2ce65kZxowAUgyPYsEOK4NNw1UQK91p4DjcjpQLaun
IF5iyacPXx7pLAUgl7iVMpqOGSIBkJF5fmxOltYyOe85SE9D9Wqzcx1Et0DEqm6E
WXBkG0krkqohKnZoeyWFel1B8VOSdJT1s6kmLxZ3+tb+tKolXBjXvfcgToA9R2UR
+VetWLXZGZnZu0gF7kuQp/Sztx+sGVMEUaSxEOHm6T7LEVhiJ5NdXynBKCE8m1x0
KHIRgce7y7O1E4I63TdoeVGIX01wsYENCcqE31KcvIhOG3pMk3swYsYiFn4pSRkA
cdgS6uVjd7JCBdhl7Y89KC2jKwb4V0B6mbcszhSZnfeeRMBqV4kspt/bKc8XJzid
ZmcDhUXERPAhaPXmyI4VuOWkeImNALuqXpt/GoVuoVW8VWED11oCnffmjNZMVovE
NUOK7U42Z7RRHqO+p0dvzwpjXMbrjb8kQDBTpIPO6DOtbTSrkO5qSchyOuiQ5Ywp
js1Q2XTKfkhNCtW15JTY1FS4/HxSpr3vZVDNuJF3cTOVVSFiPTYUDFfxgPT+N19g
u8e3MFplIbM0c+93x6/HZ2q30xQvBq24MusEew7dN4V03A+pCLOBaVDLhFgBqr5j
0gE83ofKvQyjeOlSvzOCKite4b1rHHiMQ2gQrx6Md4yZjOLRlVWhM5L8N/XRL59K
`protect END_PROTECTED
