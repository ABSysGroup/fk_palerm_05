`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zi6cLzrbuYJmciOKuEoxQPPKPW1dJm7GBv7NzunHyrsyr1UomDT4ZCfA4RLaRLYr
FW/0v7/xUHPKQ0DqLQ9w0WI42p1/K+tqiXU56FRNaw1OmxH8QeHI2ZXxKHdg8GIh
llAWAKa5m5TQSAD5ml+4bWvCqZXWFScPdqnbQVTRsexPYeMgQOkaasLHdLPeRCvr
2SxufDAVsauSerqMzRGv+XDOISr2G6WJEL2OrOm/Dq0cghV++WKRINylHah678O7
MaK7+Ab/oTgEPblRXrxRhRKPUJxoWTjfFzRnXSU6m49zHzKofwMCexola9+kBEPO
wTVUB8I5rgB5W5oQiTafLw==
`protect END_PROTECTED
