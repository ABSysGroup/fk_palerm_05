`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jg+NdVM/a+CvvgcU0FwCUKcNB3rQk3GzYH8TUbYYKKXIukm1n6XIthJJkXsqgQtl
xnGbIhu37seXhuMXYNehauuLdHykZ7Gh7XvLILbQCynCE6LX7D5SYvDZNdiJYFym
aEI3j3ieDF/kj9u87nqVwug7XuRP2jQfv+rNquog+Mfn4a6lrMKSWKwrGpL4f48F
Gf0jyV/IEob/YVFi+VFqauayKPy474wi+RzQ1ylYsp3N8TMp7ezO5Da0L7xkyuGv
KGJEGwEl8EWduFV41er8WooOO+i4FhANd2ssMDQSvw61JLRC6hEocKi+aBeX3BXo
+9q8t1wNXfw+5FIQiPdJXQ54pO7Q1KW7d+8UTyQXg8RhT0wvJ9QYze46GEybd4uX
qDbCBIgNby1ug7QHXsMAjpJUJ/YxGlY7HlLIIvTToFGdN30YMMRPNdoDwup6cHun
ST/htVBhiNqEgxV6DA6vJKp2VYn4eylc1OB5UOJWvku5hpGBJ0CZ1dd1b3tTyU8W
Zub1FlieJ/RSHzU/kzeg1LWw76SEYcG23hBT7Myh7njKjO1WeWB0lxwWSP5aB03j
od5RDbU5Ly1MAGM2fRvTre3LPv3Th+4ufv7VNcGhDEQv0KGjPU6KDuqP5HsbKzjM
VqeVgwv/XcaVNCLyak5yqD/GAlye7HTdSwoCJEN5jZ72gCFX+B6VYNlQaasmS2wU
sr/eNFXaB48BtdVnoQBnk4AqSKL+ifztRZOIZvkH0/8sYYTVWZ7Qu2u0GthCax46
sQHIzcLqZAlScU6+XYxxnVWcakIVxtzKTHI3A4xN+oV7ZYbPpOT8ri1MZIv9/WKS
rUJLVktZn303CHXRUY9ILuV9plaaqnpJFYndwHSElzBOPkptDy7XVPjWIwIONs+R
sQ2e9MphtwwitJmuKOpF57h1qIZEBMTI1CuksHEaz8fpq69YBQDm2PZrHAp850wr
qA6cfgBQiwtn+jjIqXevK5l0m+L31B0N1+BEuEw31kte5wvYo05s13wDKkCVCmZ9
DHZs56ZWs0JJ0BV8qZMy5vScshx7f7Ijo2ocWy/f3X+sV1C6YJ5sToV7bYonqdRL
BNpmW4ECQO7hVS1jxmlf/wi3vl6EKEpZ2dPUGuSzPOjUrwNq8l5+1EY3amUUhZlv
vbK1guUEuxVbrrGi+QOAAi6lraKfPuAduD+51hwY5q6h4qeXX6drn5Qcwet1w6nd
l4hNx4v1UZkyYuI6phUK+lOtliWNVsJN5VmZm63njj7rYgH/MNg8iI38LG2BIsJ3
7qZcHMYYLAL/FfRhzYHY1Qg0TFYe8J0IDmNuMbn31Aftaew/XCc6gBx1CumIP+uo
dJ+aVYH9GObgGVpOCtUuiIelitz7wPCaBnBsirmvtagC4RCvXgIpw6s49nbPUj06
77jXMJHWMdJekndIo8/nwUjg9EOLaZK+NowHTsACVauH5ugaKaksSgAWmVnlY/k/
KoddxCxoZwJrtnp+FLT7dkKdWHMCKKbr33QQtFiivps95RNP0A2dYO3eJxiZ4TFd
+tr25wqG/nGRvSAwrHQGGJVPrLbL8nn6RYCRIfX/b8YIZ6sILr9jtOPIUHEmCl3W
jUVtHDZjePuMACKXrWsL8Kg1r95gyqXOx8FVFq/YHYo+SIaYlnCEh9/5L1K0btK0
oikceiMxfwXSwch0WIG2vml0AHoJ3MAbI4iYfTVemOpa1QLRbhS7HM/FvH/lzY66
7VqprCUYIVLf9xAnarF9401mE8ypwUGxV/ykUUndBv6LaWxgxyEdg2CCRGJa8iNR
DIsYdr44G8XGycujHyU0DSyseLFKUIEg11WiBJlAsH0tz9w90CONBvX4uYZGsSNG
ceV7ZLRKl15CteNNFZuHgUM/8hQstYmYXCf7ujAuxy0r5WlkWfA0ICKeAcCNzJ9i
rpE2oslcZme8VxSqgKPEPKyKoTPS+NJKvgfRVK9+1+PRuquDS5vVadTpbpisyZNZ
ZgFeY9OXsvRGMycwA59HFC0Qv3kufDuaAjdGRTobWMxRzs2ginK7HXiM6Ia8Yh97
qdSTBT9KIHQB7O/DoHhcDK9u9hZw9UiED/aotn7wwkdERVhctlxvNY4VMIpQCeyW
OrFUaIzEYYuLK3WBDNsQs0XUWwqPtnMkxLhBFlOuzLHyPuAwhDocnPfqu9nsY7dF
jiBujmxN832H7fedihbgngmX4jkkkZRRJ/nJ0ChXmfiQJRtK9TOTDXehf4P3s5PP
TdmJj3aRgWbkcKzlSaRsiQlvFUBe4hKPykS+cx9wwodnJXr3SDhZaaQf4ZxU5UKe
3ZFAeXjoIB2sBfxCT1ZWNqjD7VsnY4+VMspF9Op+iyhKbCHx4srEhopNwwkVHMpq
MJppQsjslefwxuCl66yUv4WiBNGWeoqPXDz4GoncS/XrgewCjOLCVLtmuxPbKv4u
Ctwj29gnKfV0keq9ir3SBu4b5/QpwwfzL0d/JD8dzSdTjHMur55UonbdYCQbGlmp
LxVqZNlCszt4RgvFJGAwMiIT5YLLNF5PM/tU/l1ClXvkSGueqtl6thwrzcdAX7ud
3REQ11d7l8Xt8O4iRoJJW1SmWl9ekpg8SqpUw8inxVbxgBZa8HZ3parKjKqFsCUu
VfPelQPKsUjrFZsnsOKgLc0+bV7Siiap+fAdw9JGdwiUXOlxXljjLv5YZgnsOFqE
oCMy1U7zc6ggUTK9z6z9ChRkyth2jVk/F6FB4Ap4+lxe9pqcD21cwtaekJu2Mk55
9N7+ZakQdsebiWa2BSdyyukTyDZqczEhR2s67XDy34eHpLZgMzw6BQYJJlkmSn6l
f1qmOC9pYXRx6S3D8nqDHuzLBhTFQcHCGtj6n9Y4vZUAKA9L8yPDZkaJTNgDNuyQ
xk43/ntDniZPv2Y2QDTgUAEj/v98/eqjdwbSs8CWm7677BAW8HgssUj2iT53kkwy
qk7gH28X0N9hBAMmlxL0uPXcriQx2cxHY4Mgx2T89fktRZ5nw66lI8shFykFGU65
/0+UTPCXgpxWW+eBs5EfRkcu6zWtuv3874bzjao/VNWKvyM3VV1RR2QKWA0YRRa4
OT2qpaidz7vJeQjqw5EkxIJ4sHCMczQwHpEcacVHU/0i4t5IYlmlsCrI2nKoyS9E
uQ60ENcV2vENVFiwDxQP/BhlNZsdzdOdYg7TZ6pwEqRITYRAEw4LPZg8lJGIQHb9
jpA+3rkxFbJYNnsq5eYqpyWpXidCh7bIzS9AuTB47TOCNndl4mIsVU+PdewBpcYa
4RN02FMuKN46Mh7Xh4O9jTQ9haKs1pvrwiKhTA5UNN//nYnSEaMv6WytvbhnIxIo
Xp9YHDWhOaCFex8w0C0PdrS+wizfgdHOiUU1OJkY7PUGTdi/yOnB8dyCeTj7Eaek
9DWPbEjV28l+qFmzRRUgC92tQb3v0dbpkDO6LbIAks7NyzxamkEhZd2bWypWrOms
WM03okBJYSoZasoyW2EndjLpZXw4IttO7rV0z/K9Ay3frBCK6kmbvSWVY6T07NKr
aM7H6cws/9dHkPojbmkS5YLGf6/APZJLV5SxPlZ5vI577tl1x5MNGeVU1PrT5W0R
lkTPtgB/x9ujJobj0a76ugSymqQH1QtwcoQENREobU2dyKNmr6R0Wn2vLA2zl+/Q
uuGDZ6OqlKqYPkLAbXrfsvUcPhLrrXfaN3G5kXUIhhBKwfx5/jLLUHq+j4tSYyYo
6mFYdsCNStokjGyUFUTiAavMMjM13i9UNleqCuOw3HU23WzFKvmFTSfXtGmnIQjT
u8nqTpNI7ff3FVFrbIgrRurlKJ5+zqA7IuCRqgsqoSkP/Ip9n86sh4bX8m0X3BhO
cbqiUw96y1rvTvE1ld1u+kO3XLc4a86Sp0BZp2/OFBorlVWaWFlS+ttkVUCfRISN
jqxPjeIjIN+elWKQZw+tAAH6uEck92ckFfNMtTfpTMn9cdvIA46DqomjTaCjwMUs
G+0c3ZzTkqEKON9JNdLf16wml+A3riM2xNRkVUf61i201jjKI+uufJ8WQXFW8Y1C
vzGIYr5VUcEsTHunAjFNAS7/mx99vJeMvPW/TrnCnQlVs7QNcBof+C7upnakfGzA
kRCDCX5KmyTqiYZrYhc8cD3a9Y/E8jJXo/M43xTlNergdJw9YZY0kqa/9B5qVWsw
/39WOywf2UIkrp1U9qi5z2f/Tpn6xRSc28BAhXVexdTX0cqkIOxt/wAq1hRtabVI
Vr9tvbGvNdWB06jWAJKyVGg8VMWPuvLxy9BOybQZs7moQlKWuA3EIM3C8yCSyGhX
d1njS6q+nR8k4fIZ3f2VT2DARxka0l6ehMpgXk9WHGSnMvi7dBj1xupXe/PMxvrN
hDUf0/KAKQWedhMCt38UPdOmY4royYdZxgzq0GhzkWkGEXFKNRDe3d6yDcuE0ykN
igyYMEMk8VJqHRQzN4Gpdvi/tD9YO3KVxAXE2WvADEP+wgjPhQJyRsLurnshRGRv
FFs6zQcgPquJVjYuUXHixvEA4Qgj9WUImulXWFLNTQDUVUGb61bLZa6iLfZPPxQj
544fe4zMU1iqPVk7iTakdE+JPacz5Nq+K2bo8yEEeY7RY3moeP4gRq5yqJdSf0tM
7fxifD9ALwJc70Od43wJLeE3Lb4V2tqEM57jNVYQMh54EWxEQvcx5Ny1jQP5eWXp
dg0LD0Heshb5mbuzgJX8U+xku1kUyyS5tIp4XxLafIQ=
`protect END_PROTECTED
