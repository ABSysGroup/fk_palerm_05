`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fjd4BXA/xZLDaNGYCSM1vopGfHsWwO0QsqfrDqW0Z9pCJ080HeyZB5X7Ca8wOa4T
h8U+xm7NQ1Bvkin3zZIawY+B0MBxnk8Y6ueeEGLKSKvx0MWGlEpJU97Do0lIJsAO
8UchHQgbypL13ohWkv+rAJlP8QQCXu0jJz7LCgWwsf8WR0qjp2yqaL/0orjBg3RI
gIqDJUX7iafqi0JnQ08GC/gUYs6MWwrj7VteXze7GO7eRvLqILapiUOoUijIFqOV
aCgNS6+8lcBX3bQZafDl+ezOqCX6cIuCl/yLLqSSUDPiNngE9PyFewTnEVu8+wgm
XlOGIDTttJnwlCrmq2j9B3bG/q27cksM7Tcv/okAf7I4GJL4pRJcMg3nbiTIrdLG
16GW07nIuGYUD/WhHn0lX4oSQ/HQgko18LJxlf+Olh9SBwUT62+F7RwqjhOWEU/i
jPgz//xtf/RyQZHiZcMuQ0J7fI0vfQYgT/DQytR9eKGL44kcG5RA8IkGqQXHEqsn
HBUGKQgncdBto8vsyyGSy37de0f3leDlBcDaUTrQQNgc7iaCn7PRWKLhTct47vfO
unu1f2Of1lSoZkYTwGlHOMtHUyrTbd5lfNVA7T7+zM4j0T1DZaof4MLDeWdwAT4g
w6i1AeDcxb2lbrSFMfr7q5rmUss6Od2DZejDiebM1XexqgJSLezx2I/D+sF8nInR
jK4WnuZ+qrTrTexqzQUi/SDaiSnflSmkWsPL+2yDToZpxjjp6T8VeHanp0eGtkBu
cMz8DETcIVQo3wOjYRsEXL+WCaV3/mECWbK7KRhlCgOY+aLINxaoQdErns9ArLcp
59rBEmG3iDn5agtE2e8GdnctEZPrqwaLCFKI433Cr/iuRqWppNvDljl2cQnZWO5O
HrWl9xGrJQANH125iAe7fG0wNzNk/7g1Yqemtw2GvV9+QR3ppnBGJAtDxHi9z0oJ
`protect END_PROTECTED
