`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vOfmg9XZJOgegq5F0P1Bo/RW/mFQxRRiUo/PrvOZnn42BTw1LZmZTN95othSWCM5
6gqxzszxsW2SRZRAkBZZi5P9Xrhoeb5LvCb6LvREBBWaAzwDTbk9p3nB5RCON36O
ELf1KZXA8qGzeBonFRYmIJ2VIkWrBoF2FYApjC7+Wcv5v5YHTbkVC3CmGH1+7gbw
PVdJvwJq7zLM+STfA0g+mFmtkZXryeBeB5qslqo1dMNdfu0BQrUkj8CjW38fQ4+V
D1wqkl3a1Q8LqwNG7BpAQ732hvd2ZxnfEaEIsIxNX5S5vGaHkdyuad01UN8KJfgP
yuUJ2QHBJ0IeSOkSBetuabqLpItQ5l92pkmzsxK3wBbDRB2PFQ2ZKYDp2CthwchP
naZr+PPQ1315fM6mO85922F7PY0cXpJLdp+c8RVP2tkF42WfaGA3KOsuR6oeqnma
3cNkRxb7wVyY6gTZcH66EyVmtEYCncWwCVqau7LBsD6U/PHHi+UA3+JwWitl4ZoQ
UtMZRNdd2Hoq2T2dKj+NUSDZUgDGRfHLQ+ZxUZjdgRDfSvAQN2RItVSsVmcP99Ot
zQzzfufAyo0Txi4ZVi2ZbNIPQ4m5M9yNBiHhQqQpBdU=
`protect END_PROTECTED
