`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qv8yTGTfQOxqO3NjjPs/69rCfibSBYT3ZZqIDNwDbAnKuNk56AZSgkVZbthvIQCF
apEzlP7Iyy7K0igRpHnUIYQeTfHRJOeZqVQ77uARN3HVSUPyt03moy2/G8nZLm4D
CnVHjrkFpKx2828LexxOfL1Gp8b8k4S+2zWCKi0dzAHoY6NKWHnOMf7NqnFav2Zj
I9pQkIPiEUdMFfAQHGiSoFsv3Kmxkz8Hvdlz1/FvdVFzLctTfiB5y2eIrwytu0VR
qRSiiKC/SXi6Yqn/wKSp5YkiAI0vKujO6GhRw1dweg4nSXBSDfaCJIsezK32xdTt
IlZPYTFxvY41oxE3QRNoicjwmmLz84cq2zUJ70eMbUwXo4UTFkW0aOeUA63DSmhN
sADL3qG+KPcO1o5lIto1SDyI+gWJBlaHsov6tCS/vw1Tf/Cg0WpRAVqQmN3MaNZR
8EoeUdvG3ikRm5Fbj0oEUNn+AN1a0trlgZNlbESJPllOIeS164SFYAznR3MIRBvC
QnrbW4do1zQ3BPj9JPO5P37yNw2amr4M1iFVD3zaxzlZiYcAFwKc1IVayufFh0k4
aC+YIKJ2JVvs584DMsoakchoGI2TfKWPWI75FEmkNLtq/p5nDo6BOoI1t7EOO5rU
4wyREwMFOTzTRGzwU/t4gKM3XGcp9j9vkOQYHJ2pXpcJowavsJI8fd7BnXs60BTX
3OoIai+yBteT4lB2/r336hRIkmfZXJAUNnoUTL5tjzdrO3uiuXr1rnWskw6VwSYb
zsafZmDtCIffrYjBm6FwNo76opxEmskqVGqmlfY+3j8RCwg+EG/a7uvOYVyco9k3
KeyB59IwGfcJI+R9ksTBPNtE7ledGyMcQmQa+BYvci3EJBSjNX8WoTHiFmp6odZt
LWeH+ecBkACQ8ufctLaKr3OBh5Mbf6Blwulw1WY4SkKH6z2THeXI6pFk+ZXbFs6V
YvBFwT53lr0u/6RmsALy05a1Di9LV8SqwzDlXpsZlcMZTey/RtXZxNZ1gN8yeLyK
zEWN0sU59SjHQs/tjxnhgSZP7TrpE0NDbVyje69O5QErGpR8B2dro2zxQs71vLcW
LlXfp00u4BFYVyZPemvzKHeeNXxaQLsXvU2BTIvJ9iLtOb5OELintFurLsNg/rAY
sC2XhaHhQzN9snDd1dDxtDc/F0afr8+bJty7SC5TIV3sZNdcruIp4/8UUDo3yKmI
6ovZikyvYzAqM98pFRAxwwueqhKAu9rk3h/BlpLWyXq+zqZ1w3emXgqcuFZGZHci
8l22TfvLI4Tt73jmAc9sSipZBPHE8aBKaM9DRgy2pNc1t4oyHEw+ksWm7o5kjLXP
iOUkho0yoxx+PzZP285hMzHym/zUuRSjglSrxXK7uszmHK+j2zaOI+/nax/T/6Kf
Oxs//6nfNH3Q8mGzDlsc/fhMmADDHjWcO0BEWfa/yFkSovhAYZWm0zsU0GBxtfQQ
cWpz52ZjcGOIr1St6uTSXd582s453OOPB+euERk8W2//H5EBDm67zSv/lfBftEY3
AaPYbnT9BUCAIh7AxoqfTGblq6hzW+tCFK2D4hj6K4ils7kqbEPHnOdSRTK82W6T
pYaSYds8p1hSIDfHQlNQnc0/CyTzieR6pv7xNGWfDWjwxLa/QoaZasOP2Neo4lGx
rGUCyXZ6/NppBm2dhhl1RaWcwzPbfDgwN8j2/3rDfNKFpYyJ9i4gqt8J43LHaWHN
kzUgvtmvRzBfMQcxmkkCfrBbW8m7eOKMqw1VB2qCyoqlqOCjB51sdAozOopNFgdd
WKkoIXalwq+sTD9XET96dM5P6LYgo6vektIf9ZlpJQobjihdWyupkbuIFj0+lDJw
knK3eUkEMPPqOIPZBALzdQu53SaKhiU1Tr60T9C+BRGFITyqUHrJtm0852slgKwj
lvks69G8CrQcMtBA9Cr/W3HX6lWcJvJERHLH/MqQQT/MlcqemnWDw9CcSki0ab+U
`protect END_PROTECTED
