`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SNdWbjA8VYzOFCCy+5Q3weHS8j2WTLRDuTX/5k5sTBOpV6M2dYqklbT7HSk10ZrS
l5mg7eT3MnHLklEuMup4B2tkdJGqZ1E/x8ET80765mHwILdtz1Phmbj6z+EnmZJK
4bJJ6OPhNjEe07cJswXiZTtEn1XUO/yruYMNYdSON8R9aR2tWtbr7QCZqjk/POz4
0SN2CbozH1RXUYWkzhGGaaBrjV9XvD+97KvbHucy15gM4CrQWa2R1mmVYBZQ20qx
HBV7QeVEImX4K/Sq/Xc6sMtEnmM5u6VplAXeHFmv55gRRhss60uUYaqN6TO+H7em
JGF4m0TZAbpkXIMgPRUaZZyhSEoSYPwi+xZWsESh7ym2QAWS/mTxUjA2Y4uHNluU
1kFT1eGFu1P9m1SzH5Uv/nVNgfl/BMUqfqFliH8WfNOvaFLX9RXv3P927vl2ndLc
zwdeK0CNI46xVHJX09FzIn/AEXVh87r7damNjEks+A/IFH0m7xp3IX95D700U/oY
MLLBVv8VCmwHSvZyNUMi0wGOGuodAIXUneWs/9w+S+XsYWrH0CCH2vfCX+ldkCEN
Ejm/0EVDm9m2SLjyp4+FogyXaYY2kmXfrslc0tOGIuQ7oyiLYOGPw9xHUbsd4d2w
wK3lM1ks3GGRCijcy/d9tXZgdoz3ft942QBIt2Q5ULlXgsaP5U05PZP2PxOZFKTv
XeRK+cgPYCnA43osNs52tRWSo4WeHJPGTX3hQzyS6UECMAzq/P7PQH5YdC4I1LxL
IT9Ap7h8jmKtsNHoLPzsfw8lAuaFoEIX0iv3ThsMpmlG3h51HcLlF5DOpwjoEiZR
6s58XOhfnEcAddQBzjtLSVG6PbnQLlO9V2D7Fqv1+1oKX+iIcBup+0XtMx90iw/Y
O3mWNNblI6osD9LwIzsSjw==
`protect END_PROTECTED
