`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Z/D/uz99aQD5VHMRNwdmh+xR8AlmkZhGwWrg9ybo0zK/ew8mCWdRSe7tW0eL0sD
lsHY+xlYCvZJoDTk4GqyI/B88Eq0nTaorXtEsuLhYooH5n7o1nBdNlEHq2pTIE9K
YYRP2zXR4U31rFPYQ6uItkesBJc7N9emzcGUAtlXEV1kf/P5E6U6qr70Ta/X6TfC
+OmlmCPJh65jwTMQCnZuUXeUYxlhG7VORtQGZ2XzpbYbXLIqkaWeYntifABipPy0
yw3DtuoI3+iWKS5dWx9uwl44tnTlmzHYtDuNEWaAPwbvum104nHx8nxqIabpVaXp
PgnLi+scXVLFaof6cxJ/KVcdQz2HoOpu34mWJ2LsLJ6ZyTwyvXpe8D8DpTW01nG4
KZD/RYTMMnyhyhffELdcTTRylLh/pV8jaMXgEnKIBTUBTmW6cIy+VpoZdDuTDafe
Bhd0OXfFcoYOUTmqWzXl9ITOjwzc168OggFUZhpqXZSA/N4VJN0f0faFAXHTVc5Q
G5BduXFWuHMs04eLios8jbIS3x1MJvqIGjiU1Pz7DIhv69J6hWaGkfjsgmqMV9P5
6yOArKRb8i/q7NfxDHSjxQ==
`protect END_PROTECTED
