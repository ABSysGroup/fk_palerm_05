`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p75v1TgExC+dh4IZtqr1p1E8o+rr5Gs8vd3dmXCOuuxtlOECcmvL2cwlDp6tHrNV
lujYNFK0cqiq3eEpcHxIM4omVBUgXPr4IFdAFlEWecunaSnMXn69Xhq1f+KQfPeO
v3z6UrEiw4B9fF9BHSb3fwR4q+sl0r3ELhhU3GhjWcIYZq84dYJ9jaPzJioT5qej
ulqx++YmoT5H+PwIpN4qJL01BM57tDdko5McR2iyrg60LiiQvZWtbH4HsOsJQLdB
tk+TZ6iX/bq9R1TrJFvjlwX/tb/kf5hI2Gl/nykGxD/R5OHEiJjFsROJ27fBYCl3
1sZCQbqxw8Srw8TyAzD/jD5M40OSuzu+o7/dXxPiW8yWSpslV0qTzMYDChpl+sTw
ejv38+ZtgbbKzggZrN189udAT5CggFKsQ/neY+XasLP9/+BCNdKjkScQ1NVdCrFQ
a2L+xeo0Mq0F8N+8+RB0ROEVv/MwesGEuio4/RPCj/SUSpAgD9DOPF07egFhGX3B
5tfcCXctzG9scxWo9Zo9djbU3ARWKgSiS3mRib+O3ejTH8kmp9g30dMZ2IhNwSyT
UESEZiJh2a0ZoWWDW1OQtTp9Mj8BhABrGjwG6X8gTrDDZDrmJBL5wvOhY/O+ariO
rtJiyiScWrTkn2Kzaidi9CIdbWymduE+GexLYEd/Bx8URi2pln37ekNtHU2apdnt
SHQLRp0Qtn2LNHtShGhZNoK1Da/vm0Op01r3FNfMqmeku+i7Vql4W4qv2tlqKrTo
YgqkcSmxnyrg7p6h2reOUuFFsuUpc+dEPDftIQ3cleqz133tYFcBOBroNqkepvT6
BUedai/GEDtRop5X3mGBnFS/Wfrxho45VGJQs6GJ8hxfHXkBBmwNQPNcnN4ETj8I
cBLYZ2ywq6TimBvT87T+Fe0rZ+HlVhqiwMU9iSQSmGJSMMQYNqFKCG6g8oGLe8cS
6Zw2qy64cxd4EXJswX1bPyc4+60dxotx2gyex/i5LsROM+qloJdCftZcRch64quS
2yF8Cs5KvUxtbLrB3Sw8RP9Fsj+RxFJThM5R9UkVpDYKCkDtWl42VQoUXaY64MGg
4j558R3yi+aJvac5+nMnKA==
`protect END_PROTECTED
