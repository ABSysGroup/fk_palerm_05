`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wL6sU3Kla5k8YL6fJul3EndwteH3lyway/d3cHVhsDxkoMWzj3sSb/U3YuAU4NR3
Ey0ORMrrImhca2ylP5TX+6zmcTkwq/EOdW0z1I1rG+BKuPsoO4D/VzZK+xuJkrq5
Z+F8DktXoh8uRkz0YOsTA0GdaKL0Mel9vueU35cp6UTdfExVog064NXpdAEsYqNf
em2sVdmoz8aVjscdtSxo8ApBe32s92ZDlJMaX9WDqUnLp1yarL0Beask87tRV+6c
5pD5pP2SrdHAQ+vgl98apcivTXA16Rupa/FPwocwhP2AJddvaX1LLOcThOM5j4C5
g3ecSgXxaDb74lYwbSBKsv2ZQGOLefyn40i2st6AoFud02T558CPWlFrfSa7PnAw
PXcE0NyEgFb7LrTtjTv7+jtf0qFLuv1/1v/9QTiqvSt00opALs2sIp1WqVScwhyH
x/1HYFQTzSSEtMZ1/0A7SHn+tGD7epFAq3dAAyt49PyNCAe4SKmEFDwc3iJKJbwQ
p2TNvRCskII439oVLl1omSk+8NEidRm+AUHZcT0O2bT4kffqI/KiPS/ZylQRZnvE
G0qPEYAfKg00o+AdMRpSUZ+IuVLobotzTfGPnDoYBFfkY8AQBlW3GoAp1ByGfA2A
N8iRWvPIWGBFig/x/7NNGSzGm/j4utJlllcsfavAU/gjWLIYNGpB6l7YdYpf63zz
/fZqI4vHSX95LrHA1g6h7zAR1lhq7UBKFsGpW8B1fihR5d2G06ijKM90nYYEA4g/
DSLXOuyZAuY6K2B0ufE/7G7DjHqXYIRIczq2TG1VLwa/JZQxcnPTDaVHgR3ANb25
yyWpgMpGIyEHNfD+BKsT39tKILIGuTmfOH5XBHhzmAaU3HfkVlH8faVuFo1BUEyt
gLdE4/kUV1+BFcFEvNzo2tMharxj3uGaz/gcq3e+6ScPHDC+90x4nWrNG87pm2KR
M8L7XHuIzIEfJAkeP1XF43sok2c6TG1/YTsn4NPY0TYmnSimkdxcNlj6mTxIu8ek
wxbpiswVcsO4mKSCsQGl5p/lgcvYZz7Ih30Ssq1lmnoPplO/n4EZB8qi5nLLUOGY
5r6ZyFytgT5COFm8+S87LWTI27SWjwutKJsvPxgwk3y32WIuAhd/Nq4b8vJQ3kqM
hzEYRtRtgaAOD/XGSYf3O4OYcXfyflsfOsngu06m440EM4FZe3Zd1/wldTCn6tgu
c86h0+V919GKr7PNAf3rvePYBmwwDnM03rBd78WuS/JZ5kf4hmZI3nPIje0jkoSe
k/hLkuci+t23gQ6TGk36eL42VA649R26hYk+559cZc4e/jwjUZhBZUMrP6QpPo+H
EOmPyw+BPzAMcCKsX2steScRomE/9NphxguU/cBmK1ozxWcaZvecTfCtWkrCO/dK
3wFGsk5tCtuLx8ijFkmR02Nbr7T39+422D7Z+GA4hpW2znRbOgat3RIKK5b5dqHi
Y42B2XZn4G2394sBZO5Qo+C2ogZECXzVrS09M1I/clh1NC0ft78A/b00HxR1rQeo
ZHPiqaJgnk2U0MubshkMqTylBBraWzAomwG5h4q6CZFXzE1/RZYOvaO4Td5Xr1Cx
2xszoWH+votpfwXT0P9Sb150/cMFh0TsYJhAdoO2Dp0EsXfF0owyY2w4XKNRDiyW
9rbE09SY13i3p6yByYLuwfJOe0CQPcFArSiNsE7WjhxHDMCIQimQRLpplixIqlO4
OnMH4WnPeyIseo1EQhe0Xavdwtyt62ixNggmR68QWEmEU2oHJdNHn6Wky3CQ4h51
B26yJVuKHG8nGwhAFNmdd46zqcaA/999trYwl1zNC38=
`protect END_PROTECTED
