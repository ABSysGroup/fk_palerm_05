`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0i0uYyP6iqgRvj33lGpJCcLTbwSqWk685zCcDukgBsdj9xHRDp21KhL3wrlnWKti
+kUxJPFIJE5BCor602UWxm1KBjhQ5FiBhYbCd7UnZbQ1fc0XcbEeJDXrCtQHoDhO
YgtmthQJrvMsSntF4ElKCL237a0R7M634qJ90l5L739v+0s34ZSpevsWSKYmtQFa
B2IFurEb59vAz6kK5GysCdZP9YLz1WmRfgpEuqq06gCL5FdqMh15VwGJ0l27rXTj
43eMgm9pO/qapyE46AFIbjRHe5GhplDLK8q03SQKlz9jhtnTnn5y/DBq/RYAl+wW
DTuh1kh6EFbWsRSsr21S5g==
`protect END_PROTECTED
