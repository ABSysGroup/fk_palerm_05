`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uYD/UxwtTAPu+OXS2aULiWCIvYrXdeEEWarS+H66ApdS72sphWn/oFYxxr/1+5QY
v/MuBjQneIQmwiKOgFmEl//uQz620U0zFZo8tKpGAuv6qodLtRgT/gMHLdvmsWgk
FfwhB1LEKKedRBKCDDer9aF8vq46enXvF+dbLIr5wqaBSM0IuKw0zH0SW8bwwmcM
JGiAgEVYRdEYgeuunbreQ+xi3uhb1wbcUj2duNdTeN7pTwMnqwKrhcjzD1JAqjRQ
1Rp67gTdDtoidudMcm7D67zbnriPK49m9qeius//ZOyugMPLjocAhIm59XtLCaPM
FgHOXcxScNz8oogoQ4a3dUgHL8U4EOgC6VfhYy/lCmpIitHZkK/oH5VbtlK+HTOY
4e6OTcvOhJ3Nzf2vfj+FtHcb02HvYcR9rPyUswohfFeE7tOKmwX0/bh2A0K50cjp
D9LXzeK2XmFLVozMe5uvxd1u83grCkGjYJwHRg07ca6dFpXrKi9fZXhYU6ftniUY
xlxWpW79wcE3jrI2b9j291qUQI0EJca1VvMOIXCo+i5pZbzBHL8w/R+Xv+d0xx59
QAfluKCS46MD6s/mk85IV5KQyS2wwRhkDy9NWq3qV+jj5e/QHuUhZBX5bZQ1QDoD
uHV9Ah7l6GExxxmA5dNH0A==
`protect END_PROTECTED
