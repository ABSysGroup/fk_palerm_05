`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VhpGGoKlcn4xFYo1mm4CrSZE6Lq4fhooHoxmtiF0dPokeMD8ZNkOUlXAeCkjy3xL
teOFd4j/G5FWD/5w/c3Oyz0RmLBsD6c+vEbOCYoaay7hZzgGsPkqRmyI/IIs/PZv
T+aN1SVBsUZGVYRrTDywhMMiyzMOs8zGWASL/AqOYp6PxBPerG1koYIgZHScgkOe
JEnLUrs/x9Jp9rCh144BeyYrQA5VkJaIfK/hxmnW/6xSz3xGZryOL4XE3aLCcDH3
X0yMcBTVKp33RBiasHk96c55qx4CjAeHVmjRo62wG5Wo6vmDvjA5pciUiOL1J5aE
93xpjw4p6DlXwbQkNrZGOs2QNAqfdfhluvtIuU4lBZmV6RFD0KmrXjzxLtzzSbe/
2rSvSsF825DEvrooKPzZN4xbERi3QSbA7HOPhCnIYvlsis2rG1lTJpm1qhu075l2
cLnPqpmqnprMkQ3RkuMWzQRjUjgrEGiDUv0432h+ldqRHyUM+rmj6ru/kjzy7P2W
`protect END_PROTECTED
