`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
weX4pfYYGfN+z2ul/j54yBjuCJwoh0b+e6xIyFivybXZpEOmZv6Gm/NOxSMl5RFD
dpmru54kphn8B3zdVGEQ9Jm2UNJxXEkfWcfG6N1VukzoRC4pi6Mu2S+k5Gfy7A+N
urnkDBdJN89eK6gTj0paIJIK/52zJZveiu7DOJ8wHYnQKMQUDZ1qLVmpLk0fDteg
DlTBf6v9WR2Yt9FsgwqnwSfbxmVj8jmEJDMHX2KagGv4Le7fCgbwejGXzRtr2gMF
7J9HSKI5KDJWv7qO3dsguPZ3Jx40dMIXuzGDUFrZMWfXHxgygKgGCFp+NCKLZZtc
+ws0jn3/HkSS3VBxiDvoG8+sN9wjVNgjjoNebXRxwFrF5TSKcS3VMFSPhC1MzECU
L+8ghQL1SBJ+GRe9XwlXomz+wmzGOWzaDJCfc8GWnKbchsXacE/ioFY8SmxF0IUA
vi6PFyApgmEXB6RI82/PTMoXEHYEu24P8QtTNhWrKW0MP0VohcVZmL9g6LDAbp2z
PFbv4FiDaUpJh75LT/fat0sMFdVlvgKopB27NL+FzmT1TmB8pDyLGh8bZsMOlVPq
d5VYLP3Or7DHqlhW/bXup2ifNoJdGR+SOy56bwFf6lb8gZmCCL3LkgBSOj+rm1um
3xPbij9hPktEu7kM2+eFy6ocVvh9Pbtit/837Bb3nhNPGePVNEqM64TtENyVmbtA
MAV9RxwWkAY9bc8CeX0sxgIxksPCGFaWlvZwa2vd6kc3DY7nbUAvaKc4QwjIdsLQ
yxXAqEoRYs7bzNa0HV6eLKHOkRzHij4jJKHbi2aVy8eBS0Z8QAdzeVbtcIJKXEEx
QqVCUm0xonICmi4db0xMZWduQ72yC/DRUi0A8ymINY1EbAw3sAPNTkMaK09dK5y5
7c+K86PZjyX5GIWfNWz8tt339vTz5qC6kGUMqIi19z8sxB32YNBe9PEomwG8flr1
ABprx1UOBwV6uvCJDrRYGoMESj7Krrz+r/cLgCL0adFkDiQNAjIbdurDPGIPASwn
pMjHt9tDHbPR7qjhdMOQwH+lM0hWmP0NzuhEfGoOeLL3yeitVxGwDt55fmp1SCtO
iZtA6Ox4mMNSRR3mAGLZQw==
`protect END_PROTECTED
