`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m/XJ9WXzgOLXsE7jVLRhwIGMVnFeNLK2gw1RexefvNKRzJ+xbsBrsOUB0REWZi24
l5YgdLdqQtWVZxp/C58EEzCBSfNwy9XWAGdBJcJ2q2A/Ni+qy+k/xx+iOIbMQ8md
HC9ToQ4C8nteMvILy6Hr29azc9DI8luyV7u7CijuIeSwTVvtHknamgkeWwQ4whUo
8IDfvz+PLFUEZ6E0r/miHL9BXv8oz6ido5Hxu7of3lbyMWOlXr9YqnPeucH7U56r
tD7VzYH3dY2unww1c0NlBsQNaY/vYHxYvH1RKOk0z6rKhc2oIdTcmpUUG8+cslTu
3z52lOD5tRz6SEwuTX/siw==
`protect END_PROTECTED
