`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fWw2KIhhhkMVa/uYb0OSdnFKQseFpHCYrwtfDqyiyTiru38vgeOBGC8Pr5k6RJDv
ZGKSy0pdiWuuZyUCohRIqvIQGZ6P1/0ieVT05adI2+wfjwvK+r+GCjEyYEnAGPX0
h6kLmOCXv4Azy5nouRL6H5gRVmz1gnezWg8CoiN80JM30G7keiJ8GAPqV44Cm0oa
2tbLuq9ouVmJ2L0EP6XHNXOj3rXngTQRDMtxDorsii4oNSYQETIxqoURml1jc4+k
vzWXs33l7vdtxdVJiBDWfJRmH8vYuXsvVYY5K31FOvF1+KUStbLI1Kjl1Sqz01ul
xPbiaGS8RuuFZgYSO8ueSRFiSi+m4yf8Z9hCK0MKl1gJT9Nu27W88iFzTrJK3hZB
XBnqqtkBzgInkz3OQEiPREC958CP9gt3+0h1qm9YFI2HFqp32ChIsG45Zvce2shn
nA1Tii0lwWnojoJMhfYmDdR2BRts8ibFkyAw9SLKqHEr8zjd/4GzI8NvrfcLYdzV
InVe6kuhTVntZv036LGtYmiIOdVJfD7frhBTlv/YWOxo3wheXUs6ILi1ZxdY3TY2
gJj9OTUy8l2+NmhmH/QFtNj7d9Kuu7RRrXabHp8lda9LdkGm4sI1envW1bc6gggW
xQ+Rzd/ROhQHpysfU5mT9B19y8QLj/g7IzHSKz1n1kh4hgDa8hM1GpB7QonMcMGn
HPF7lj1iEDuKvCM51GUmvuwPvon9xqITpJMNbIP0diynnUaKyhvDNYFbB8sBxY5X
5ET8nTuogJWEo0ML5EcclxiedrPc/DqswvZCL/H7agjRXwIBnnJW8cwsVGyp3BTT
h3SdZI0TzFNooJOvk8I4gaYfFGCxSyOjX2+Ec50lJadOcPAohMEQ2sbGhFSYeVjT
LJ3N/PHuMCXmdO1lnSBn7kxpIbw7tyB5frsKWtqJ3tO1rTpSPviiw/532G5PUz20
Rdd53vGzH8SOrlCBLZ8YZY6ESlnU5Sot49sJgiA8bp3+dFnVmrsSnAWT2B8crdbn
P9ne3zdQPHPY5wwxn8+GR2wIYN7YJGylYDb8OQc2T5/2U8fSPVndjvbrIfdsDMcx
foXGuEoaS3cYsrmxteVhTChAcnaWGJi/KAwmvq0KCPQ1FZBz7CgEqZkAKSHmO5YZ
DYj11ZLy4IybWPWpxnKHpCz72deH4reg62pBx6pehJKYJzDxQ3J/bSoquODxQqYe
hFwoZ81B34gVYIyTExtykCzDocTMrv/hwNfm5xVkHMBhp2ivppYWscfib2YSVa8J
cih6RJso4YSqcKixE2ETeWtKOllCkyfG9z+DGCRrUJB5WNoVrI8ejN0u9NnyKGE6
EvyRBSDNiZxGSrRRIDGPialA9pH2tPmZjuSJNyhM9vw02Hul3TFOONMVaMaiTcYG
999wqgzmXhBnWOg9Ym3tkOSprSOTg6VKecRuCdGQDy1HsZS0JBVAM4TQl/MjSmqG
DE6iq+ti+n453DyYQaPLiJgThXxbeNigkqTdXLv4BC9P/s4TdYmF9Z+494A/g499
1DsKPqV/gomdotkQ+uWGhCr4qaqmuFQ7k5PjPRv2yVe4VNjbpK93QVTiZN59AQAh
7txHAc65w5RzGqXeFV4k1upfRvMfiDCBv8iei9hEvWzeeGWKUfPgpw4N0TqW4koH
OciO/l8IKOyipdIWCBz85UrjZvc3HEbMPT5tlLY2rlLcRn1bhzPgEu0BuFovfx/V
RqU//6ojIP+hK6QgXFOz9MY1UOTDDTdBNkpyD7y7PqYa4utW/MrkZz8glroVj7ly
5/u2dgAb/ImRTjGxXOGUV6x/SRl7GKONbVMCJoUgAe0XzN81KUA0/EEtLFexl6Ug
B1gJyzy9kvmRbSSitdo9+Glo7h2ifMmi5A/bSzgdhchYfCIeiQj9Q8/elJxD53Nx
TksT6SbffT1e2pczyPfSs6SIjCXHVzSK9bjz1K2+q+nlJ4E8xH/8uajLkKnwEXwx
3y3XhZ7JTlzZnLzRlS/SA6AMIqW56pRKQYXJqw6qSQcUx33iWL0aJKr7LUHorhLv
VeoIEmbAnpJSu6KHfUcjeJaIitNAwPsNVe8etNWUnL+TlUpcbUx/E4lCBjt0PLKa
ASbf97Zho7VvAeJoWmauQpmBc1zRiW/CUM08sjK9aCJlU3iUMbDJuSMZxGwJmnun
yQzqWcJjWYfScdUwG5yGQ+4dFG5RRgpA713bGnZ3197HS3t4vCxd9Lb7ljasJY5c
xfBXkGJKADJpShXrP+UekGt5wjKGaO9hqSQkWHEtXykQUA12s2hJR4y9moFK/4jv
GpK0RydAd+rTmpzjICshEIajtKyfj0gVhjVh+MT0Gu+PJFJ4MvI1yFhXyZeDYetC
3sst9/8rtOwAXKITp7steGvZ/b0IuHXPZvM/fE+4XJCaT+qcQ1pCZMmQwuVqhfOD
rDPZDI3WdYc22Vu5AAPD91Ipn3T6BiD7+Z+RsOzJ9Vn1bv0bjtBFnZJe98V+BJ8I
ZGQcalCfarrlnq63YlO9M6aMISJjSRHM7CKyhd3Dto6NRXZ6vfyDXRKCFiMR7lCa
2oYCkqNcHtbJ8YuSAmaeOxqCsr5k8hGfwLYhETmFr7luVUv+xPNwZNGrz1fw2wsF
QQmOAEVg5/ZzSydaKd2tlk6rmob/ccM8LHQ+H8ogbobPVnp80ovNUSmRUGbU7BRy
I4Mj5dWgZTPepdoVhjljneEgFnZJozCF3CMO1ahbVRuoQbx2QpuGS4EtAn4Yr3fi
K+LT8Ii29kFeElknIOtCul1cHbXb+GEp0FInw/Sy0dV1DUw0uc0jX7yl+zU3dW3v
A7zzWzjkFY5FmGoHdA0YJmnlnoSnRSYPal2KxDTa7cfeCOhuvyo9VBbAwzHt26/F
jqIb1AnTCZUHrXdkaHHtpGweuzsp/zUCKXzCxhToU1ht6WDDGBkkrMrGuHY3t6E2
IKq54U12+vvTDd9cuBGlpio8A3+JxTi/jpBRDmbu6UUzvSvHAUVWJMacd++z4Cf9
+SUHEDpYw6juKkFgMZuQTRec+TLh21gBc/Io3sSaSEsAt0KnKcS1m4T1AW7AAMKq
7VTP8FCuGhUM+cfRMpwzWFx8zuHm3uyeAH5q0084YCnjOpACTyIAk++ihuenHIsa
7iXOmy1BSikgWx3XAL7VH9YJ1j/HTLkBdcLyTFZnO7GH/9gpOUP+rIPFwYr5HleU
8Yl/dZbvKcx2AwDaNEYlI5L41hbajg0iOhO+f1kJ89ru1nccapWPmHchIHaDpfMZ
q8sCKxtv6u2d2bEcZGGqanLMaiieAKqf8sFtF8sxTGFsvOrSuN5taE9LX+kSYYt5
D/pcxIhiUeKKoYfHxtAHq+bQRGGKHEP9xHqLMv0EmgHMf1qbZyvuG/RoH0YdrnfQ
aA/5MPBKw4+Mgc3rWiboVtq0t6z84mz4vPFCuND03vVbdT6YH6ufJ3xmpPjft2ib
XYbMJXukDX18dv9r5EoZ9VS/76YtfVQhAYbsWg7SrplwpBkxJFVGQ6sTsopHYx4U
tw25Dj+mxGVqcJQrscLT6YWGD/beYAqK5hFHjPYkpUyZ5scNNfRaAq+0LHNVq9vo
mNmoKc7DKyvclBDC6sf/vfieJEvaE1OWlDlrkIUxKkxh6yjZ4gE5A5h+MyZ1bZ43
t+l87kMrTIPwODRUPXFzH57SySOn27i1p8aJc/Tw4yld/ZzrAHjTZufrm95JicrF
Ps634NQv/g4XHPeh0Rs53p4GnOV9ZDTR+3URmn3fahp+h6FXCfGaWuhMwN6PWiAq
6DAe7bAmbsvy7ORXydsKdPfpB86BxDpeeOyJ12jwtXofGwT9853ItlPbcmTpmsNt
XMFP/jLRwMf4XgM90+X6VTEESyB7DVQD9sDenNsPSQw2cWPDnqbJu+LPtIPgMWB+
EIfz8w1OgcHTu93uGlHExmlTKDmQwjSjMEFL14sJUdCoBT2+onGjt9u0KA9m3CsH
Hgf8YTzTBpenYkU++aVXzca8U1TkdsX0mvb2Qh8ofHngCtLkE1wThIp8K5GrOybC
pXK9/DvXmjxER2HDxuVYRf0a/WXz5/uze0w08AQuAEerlrdcFfU9tQLw+R6Snu+m
AthEQBfFGrPRaXzA2EOhN5smlU8V4TVr6rFjF1hUT5w9CJz+CvbH/+yUfpVB8Ziw
s0Gex8Rn8+UE4Qqvi0TRCVt9wQBimmi0fYxEROSNhTGhg/IWvCUAiH/VbWxRkQbt
S3Ci3Hfk+1+p+3hvZmqlgv+dOm9MbmgQk+KbbADAwQSqVFis+jI0NEcicuafrzVf
E35bdNS94yuaVg0rCQkkc8VSHOTP1V+G/3ikXiXvqjyZdTwMdySUG3NgZS6yiXsg
sOuqoBELPlXozTbAXVLKyebzP/hOhE77K+h18fKnpL7H6j4hpHgjzK8n6P6f2BY4
CT3015EICFzaNc8yytUDiZ+gPilezya1IbFsojONqfc6p3Yvwg9LmI6ubJ8LR+F5
FKaiwFPa/2fqfvBlBPYuEuZjAbBjlAQ2evqzYFR4XNNEM4WdLJqNu2AX+/4ZJtA8
2TrEMSvOYoO4G51EEB1SxA==
`protect END_PROTECTED
