`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/tUqmcXvmny/oxGj18Tbnu7/ZEe7QnzlFkAIJecW121fqI0HMNXz/+hrZzYufQXj
ZP2MHoT9SM2KYJgWVjz0mE6E+4UVKZU/Jy8lk2Ssa/qq5q/vNDRcheloCXgVuO6S
38kdBPGQ+w81CMwjSRXh8haXr584hcxqO8/8EL8geg2tyGfzNZiH7+R/U5LUVxiI
CT5V7rebpVtn3BvV+36NQF6+5b1uWE68smKUloseVOCnyqmXO/SEuOu4GzKc7InH
zmWDfBmemxtDBIunaXUgLPiPSvWmqBYXtyCQUZbqFvk=
`protect END_PROTECTED
