`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
No86wS2DcKgcrGFNN6vaqPN3GHdeIQiJYJbRQg9JfyPgoXmWvlEZrDFA0NOt6CsZ
iThH8e7t456xbunyZfsWc39INmhxAwRZJVmUIwRKTv6NsZ7AMdp509Y/AxVG5Aoo
3v4OFynO7n46WDF84CKQez1sk8exkQR7e0ufP1gukDVuXO0o8icfWzJzbAvNH5c7
uwoaYXDtpY1zP1pU88AfkETbvcc+8YNIbvPxdahaj6pcASbQzLIfn1rz4xp/dE/3
e5hoj3Kc0AZb9gQSKrAES1esCj+EBC9PZgQpCVVkgXmMB/wpbn675YoPXLKNNIIG
kdDXj4LNNPPH0ut1aBPoZw==
`protect END_PROTECTED
