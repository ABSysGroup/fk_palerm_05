`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WsrSXyfAxK2R+E0isWmaf16x3oLBiaHB56ybTnOOU2XiAVxHWCUcUeJash4RMpjh
jmDgDSpdMLcb9k8EGqgpdyiJ9bCsua1StHoGD5Xz/FfuBmM/ILXeWiVCcpu9TACQ
jki8GahypXqPiq2f+ISZi6Ej2Vh+wUJZA9rg5Q6yX3vUNzZcGDkaVOb1h3CZ0moh
CEXIbY8WIPhVKFDxT3TwabrAbpLWqzRrCHh07n+xy1d8pK7hoyN11faXMf6oF2aI
GmfxYnrmKt9Xd08ivHA6Inji2nu6pDkGT9mrR3Q14/XsxkB4cef0R+uY6vS6w6/w
NnJEo2FZzBPGfgLqpEaeUX3ViuNcgMFZQC3gOYQ3jeH94O2psuy9KkMNXE24FTaB
L+4rlDJEOMJFdLtMc1jhTxCIK962HbbVA43ZpZWaBKyIymmZDopM3LJ9eco27xTT
`protect END_PROTECTED
