`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ngCE2TrLe2LV0joGracUjk4euz0y9025ILpi8Um83d0vYjnuCY8wxb86VrTS6O/B
nAP/zF2BExX8C/jG6rgayw+M15ZefmFQ17BzVVwmRbbwCkrAQ+0isQsHpUO6PLbj
MZGefypPIhfEIFbt7DuSyGh3/r7wd4vJsgWYCmSP3r1MinNugm6lV1leZ7pJDGAs
hOsNA8M6ZXSZNq5L4gt0KUBnd6plxYu/1v7KKOh2UXcgnzgztHPUdH4e0R6oU6ti
Fcfl8zV+wzYU3z+NjkQBAzVAFMnYFpeGfXrbVkHUWYok5sNFi8Z8Phb0B+pFTi73
ghSUG96Pfps//HQEIuoLy8piav/PYzo49c89aRayKfxcofowtYwQiScIJOCj/qW3
d8IJwLPCaO+E2sDE+M3ai2qSIiQML3J1fAnCgYSfg0c72SbQ36NbK12S5dniA0sk
oOPRLkB2Zc+LpUQLEVeOQQ9/2UwmJTHxVG5C9CW+g7iNQ8Boo9gEQbK49H8S9Q6O
gcZvOQkITcfj5WROyBOL+RG1vahok2unj4VchQHuWabj0I9WFybf5Fi1juptPrI+
kA+VRDl34EbOGCZbLZE+/kwmTyBZ+ZUezConwFy1n8vjgbkQ0I0oo8F6o80TxpsT
KKZ1Z6xL7ehDLYMcCHvNvspMzAGhqw5oq8vE2br5az6DBvggOgvyvrnj8lplOrSA
eFdQiosCi0o2BMHiH308F61HVvFQYHFhsG7P4lJp82MjlNY44EJvzbzDrin6kbuV
IuGCexYJeYCjdX+n+5NCz0V+8gLvmRh+vOx7AorJ36sXsKlqyY7kObsOXWZzhjGN
qi7VkvLcuCeOIHMzHr2rwd1r6XlANw6J0be5Akrukj8+L+GF9SZvkw+aFFbWOt9O
Xl1J4PLBK+3k+kvXLoAsqXItyilaYlRvXBMGNEQOAhSjqfh9FupWCh+b2yyaMfWK
`protect END_PROTECTED
