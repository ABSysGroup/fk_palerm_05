`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Ifl2P3oML3Mo1cBXpcB+uRswBjUtpYFNsTQsZyf6vjLS0Pj31Khw93XveHyzYQb
D/65jk+y6Wm+877e+J7udJFqTlZy1heGa0Sr647JaVLHrxuYQTOD5p6x2KFX80nO
s6kGaQ6Kh2E28eEYm7f+Bid2QyRwOm+PaaNF4GCC8Gh3V56fFnx3szIMAyEOsYii
spkGCRd+mYxbAwzItk5RsnODcfJqH+CMPUyM86KGenyJUPPIC3nlzD4lgHO6zFc7
neVLozZgCLtC4gi+OzMf0QR7m39yApk/sq3+q9HLvJGQotNObIJa+7InXtj6rnwO
uWRBD2poGXf3cAoD851qH3+H5BNxh7bRuAaJQ4dGJS6y6WaKbxwpPETsqU0nvwnA
Y3pQefidMSIlIv3y4+WfCF3tInnSshiBZAHurZwuL0EaRdbTZbHdygLB41qgujXw
sj5UHmBCOVCja4KAayTVfteMro1+GFlenSnDo8PNIBz1RLRCF2F6srl5Yc69LqU9
pTZc41giBR5+QllYMBfwYrNFCfPv3Rvyz88odim94u+wePAoXbZ0w7Lrj84MjDL5
hw3/SsJ7A3GZHOstPq8OuduD/EGiUqIcfTDCmAPT8kyr3gL9X2HAt+bz+CJdycuJ
rRX4LX3gcnKiRDGhvu0vguT5VELXe5hT4ciEllc5IT68OdaReKgqTp0tcfmSarX1
257XEueglNkKUBWpb/l0HQg8HR83CUtC+3io0li9h6gugXEM6ZXTjHkFvg2BN2Bx
rmEB0Hac6A+yEq8PuxTorLkYVWbSTajkMTeh9XlwSOtADAZ5eg6k62nIF0Kz+Vdy
kVc24fiBkR7hoKEFAE7N22Z50XKo5jmuONSfz3XV7Q/SyHENAVijvrujUaRufzrG
D/eoG7RECJlCaXNUk767ckmjxHDg8yD9LNWayWPisMFyOJ+NpmLKQQ4gwZjHEB5z
5rTLClJ/GYz0zfs87alguNPkE2FEWGspUQbXEkr77V0zLZySgAUPlM0K0gaVua87
N4/cUiJy4AUR0LVa7HtrDbyH2jqTB0BADDj6fRoxyBTWsqWDbjqjfXXhKvsLT+Ir
EsSHB6MTKvrtDdTbZMEF0Muje70TL865iYRMwA+SrzZ/abVZ0IF+ltFKQr86Y63w
LCP6csf5FeWOFivimkHLj6BkRv3/BbetdZqqW+t8IH9lutvKCXoW+ZQfeCDI6R3/
ajoIUUkLdxeGX3pY+tbTkieLqIAjv+Xvklk4Z8K7SvsQwZ64R0RpmQppPsDKivvJ
6SjbwtzstmVI6wW3EnFk0IsJAP4CEY39tAj9Ugy4elpq0J0ZZTbpkEgjF/3ptkmE
a1lUi2am5PFveEpeDirpbPLk+85zeGRhxqMKXOd/MELTVgK5h60Hp5FjYGt5BBTd
WBACBo/Wo+f5suAZTfKHOz3aqnzy35Vju01R1d9imNG3sz4S2OvIHUmUH/0Y1Vm9
orj0JTgkVDH/l87QADScDnfI2cevD1jQzPtKL8nbEtcQbKrvehZxu2lrRvKl4lel
hxUJx2wx972/ifd98TlX4Qu6JgfnDQsVKjhh8gAa7t4OA/TpLsl+7QImFqn2MNz+
iMX2ouynhRKrcs1ZyY61vdJTfR7TugguLoUcGlS08V7bfQHtRbRlnCE8Aq+1f27i
4NintX65g0EQC3jQUrNiHIyJ43w7KP2QTnnkGEC/LYpLiHHHUWFz5H0qE/Zq5Tjs
XM/bt1qt7Wil7VWWYXPBQb9DsjVxOlO+HSR/RZ5cPpXXGArC9Jjf2mtEYPZwjMNg
YtJ7rz+FbXNbVag1gRrumbkbsKuDCfF0I5BwI0c//mRKZLLvGJ2plJrDpPwroLNE
5htpoVSuXMTH3ParQYAnyo6i7ngv6W1TwCT+oCyxhX2vhsy6CCjgr/UiMq+ySyp7
xQD9AztxDon9jqCuBOTgH4f6h9DKmSgIIfffgnkZTKQrsLF4AZNdesgrsXyiHjXR
wPRKJT381yN4k4Lr6cXYZac7+OCTzXSYL4+SL0WYfEmIk8HBRgCjZeHyJ2+1LotK
v0OqYYJrj92nxPKV6UjPnBROyJc1moCNE9ZG9nZzJoHq3hrK+GeaJN1KVdseYpjo
qbI3q4hSUvdpIPq6IoK3z4uYfDh564dURZVqsK1O8gPNkul+StpDKTZHL4TQfdDI
VcM6VkZNmxkECSNSG6mUxwQsnIEDx7ihMJ8RuKjAqtuLFdS0eEWN1oAqDB94lIy5
/QXLdfaAFBtJk++jCN32A5ELOcAyMxhSxyjskBQXWuqcAW/BqFxycii+hKElp20D
`protect END_PROTECTED
