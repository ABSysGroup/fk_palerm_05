`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mIs8oH1//ff2ZmwYdL1+TvtE/hQJVcWR1Lw3IamrHIISCBB8QfBlx0Z2U0SLR4YM
HsIN6vwo07n0RnXPi06aMQNiCZULVsNvQ5nY6FiTs1Vzyt6E9lTMp7uPKVx6+YyW
kKngQD48u83ciNOvqujzpFLfA5I/ZNy3yTEvo4IcaVGDynCzQl1XfVIf0qWEsoVn
1x02UnvCFNfh14Mboe5qfwCOcw+e7UC5p9YpRbAw32B22iIfqmnVKbTA/E/JgBlQ
g2yxpS2QJeWa4OzsukAeF0iioFTKIhaGzjljJd5TBUTB8tj5OZdWIhEqJXJGatk7
Alj/Pmc0q+CxI7zlvUKCIFGIWi2kitT+EYze4/QdZaYyStm/4EQCtz5aSLYOqsNP
J6hgLNs0+a+Sd8X2zqMpV4aJ2ggy2R9cdx2a0DV1pgV9g8XsDOIQKp1H6dEbyx7n
AdZUUUEE+6U34a3Pc66zKbYSaGvx1WpCfTS5WkcmaQ4M9vnGA0UhUx6mrhQDiGJG
Yh1G11bbUOxiHAoBwMgl7ML44Lm2NCrGBvRvWEhpxENepyPH3dhhSzt0AdNv/v8r
oskq0ULUsKIiBs0c88frK9bU9LTjqCssKEmY0Vmj9m3yz21iwk5nfduu2BW7rWT/
Lu6n47U/eQbqP6LA93kk1uB7c2lRbr5wuRlsfur91rIY2yfX/+rPTWLKBbOy8LlB
u7FwQSHGSoJeqOCKklt2QkJqPA4cOJKHFZafxp3iXPQCFhqVDlgpmvyQ3Jz/nC8S
33iSAyaeqW6zpY0x+nqR6K2IrLV/K8/gdelg0l4ul0XFXRRc33wOaXu9jY9MYMUe
tgUjmMz9uNUGqAfN9Yg1X5BVIfafAfa2wKX+5ajSBUCcwvlOEIJyRTGl6qpiOb97
1nVwYSBTr0ZDTyeztoquXqgUQnB2FMhna0myFYWojCGuxZ2e/d4PXe/Cudv8yp48
QZ/O8MssyDLJwvzYmRoYay3ccwIxe8n1JkYKJhLo7u56bJ5PFrLGC2uuqXVcV4ty
o80VWaiVSK1wYkYEr4Kya70AJB8yXLoyH0lvMpMwNyxemqqu4K+tWsleLSdLw323
d3JnxstJUy9SlOO9p4aSAmaxc1Xn81RKQ2ejJJMuk25JJ0MJInRTnDZXJWzGVLnB
ddcyE8NPcQeokb4CzTrAqbbnx/L8RrQ7ORWJ8bccKJQzpf0mov/xQbJeOy435llq
HG4tj3Nih3T37heEhnQajrtayMaK4AMtdQD1Gqg7wZtqfRbtWpzoK+MSlxrHcMTo
w/2Zc+Cd210dXhRL+UsFY0HIAm/0f9nY9KmnxLDBvDgf4TQMMBxM2U39PrrcJHH0
t29bvLJq84twajvGNVTeAwX80mKhO79E2uYHLjCcLpkfhtVnv2dACuljKuV14HrJ
pnq7OaQm45oMGsizs9AEMmIKtVrldBJz3vhoEWUpxC26sKu8bb6W3IU2bI+QEqWb
dL3SbF5whQzJu9xtVfeP1A+TDIKIwefv7yBpTJEIptV7PqK4+GUCGGIdgW9t5Prk
BU8TmN4osPt8nndORZUC/nKFB5+SgdYc5PhIGkaVkFwnrgqwIrWoH03bQrohUxgZ
WnSEyr4n16alppoPmpbAJtV4LB91s3iNmNt1565e2zgqBQNqXf+YYksqr6wGLpDj
EZ9KFt/SGuA37MVSzfkaz6aDNL8MQDyvg15XKM2ruL02UZntBdZPKCaXXiGYoDRj
XGvcvGASHZ9uUVmaHu63pAUOjCUrNJyBXkmNWFhdUkoCeeNFr/89imXBQme/Kj9y
0QThA2EWWfatTR3t8kUXX0G4QzRLn7d9K3DPp6JjBqWgMQ6PsyVavSR92Evtm4O1
9fPirxjjUe5jsTzh/cuRnruwhlbaRfUIfuk1sxbWc2vQvAw0VAmxDUbHFxFlzSDh
xYMR4U9tJg+jllusp8JlyS7My5fHO36KR7DV6jT/NN8tBnK+qGW8RzWv043EOCQD
AQLzZaABJc1Q8SixnDodprx8hdr6IwO7Kt+smHf29kcsQSwCkr8CUxsPxNZ9kkdw
wGr0OX+FGu7qO5GkK92BMHZ0r5B6Vqbv7zj/P4yVMyrr3hUGYRRCKUrr4Xs7vThV
rVixolaLcsfEXjoK0pcDmkxcJTTu7k1+z0MZbZZzhjKgLbvQuV45hi8PfTvAivRg
XDpgbYJdnojF5t6BwdjbcKmHvfuOtBAzH2DnASnuaMhV+eqlO4sX0dG1JvUDMqqe
DcaqaYItnbLoL8tn3D13+Al4af6+m3Jl3cIzgXtmbf1nhUs7UsGgOwG7UFPuGE/2
q4iTGM9kcvhbWeV8pURTna/M6PebAoPV5iJL6QPA9j3JLJN9zDhwwjjj8VemQWi5
NG5Gxq+8rzqSdOg8f+Ub7f/mbMukaCSE9jfW33BddrbdyBNr4yCgH7GPNYL5XOvM
DPW1QmeWBKUk6YgWsUA6u39AMGUufR2IqrmIxC34EDSDSCe+igfBDDAMpFcyCpo+
`protect END_PROTECTED
