`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lb/cPVngoVunI0GcYdAfWxngYZ9Rp0x2uvP8Iw2rZK6ZGYsXxhBQ9kBk/BZyDDNh
Ff1bSjLGM/5q77Gl9WTWWp8Z9Ew5JAbtZh79lQX4E2glNreTJfl9LBnN7jWh6hZs
KX8SEvB0n6nNUSitAu1gk24aWy1jF6cV3TdyC05q9v9U5+IXOosQgzxnRywCMOFp
+Fw6k2SphZtO9ZX6TqkfufMgb8s0uSWXDuvtoGPq2y6M8+E0XlhL6LBUuFKZahit
7bcYXf4GzOwYrgP9/bx+tlVbzo8cwEvPSUqAMnmjRqCcG15gb2LaPW8Wsk5zWxMC
AGB06EwknrX7Uj7yYjej5msopEE1MN5mpKkgMiwAIbBvZjE6Ku8733Za5a8R4+8S
2rvCVgJ0EsZJBMihNfUYPJ+Q22YyHKYbefRXu14PQBxj7DQE9dxeKRP/N2ATmyJp
HU3FeUUqxHhkltUkAGjCQ4qwRQllOQ47uAWXlXznAEv9BLXmHg9dbHBuWjxJNBVn
KYMRTqSupW5G1zC2zIWtxpc0iXEHZ6NogCGhOrkxlocACPTZOuIagndIyCXeTKH9
`protect END_PROTECTED
