`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CrGQ8bjB2GpdWu88fxk9ugf3Gr8KkNHb9/uJRag4LW27CebT6V4NyR6ZyUqQ2iYB
Zhr/ZkjTHwi/fqlHb+S2uYhp7/nlTZizmmDvvb5Xfk5GdC/f9Wd7rsqPnHMMXau4
Ftc5Itt9T18LL8BQbr7Ni8+zX6Qh5BrpXM3FAePnDGlYlnflAUQXj2MeSWpYMH6N
tIUbpOfANR1JBCqLw1PJegJ2O3WUdZAsbaQc9W7iDeD3WseOPJVad4s7acNavZD7
FKGrZ5EZgtp2ZbR74K7hWMU/divwCxe4F2IwfpGXwVlDNYZh7DJo7UxySeV968Bk
rdKkmpxQqUe2swXvTaiG2S1pz0RoKh5NOWcewN1kbajvT2NJEuaW6KdjvCDu0feX
D+NAQg1jAnbSry9GdC4GphmCm+ejBOuAYJRdCbC717qMFyupH3ylszDMnTxFyYkv
curwmdi0J2oawcGmt3jjlpMw+lh/GuQTFMbnABZAx3eHOGw9oOQtrykRolt6DNTM
`protect END_PROTECTED
