`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ze9kbH+veBHYH4LSz6gn8rZW0NzZJFHd1y3IhzB6Dyaq643Svs4KnYDXyd7H0Kkx
W9vFT+Vz5+qOxVB4wjSkP0ey3YBSxBigjlcOop7pUz7HWIv4cFVdwzT5UGoMnsDQ
+lkctJSV+ncKaEPyZr5apookD23cp5tRshs9AtcTnpOOcF73BgVZ9k/OiS5+ynBJ
LnIjUWnv/QKNk/GcnoFdhvgzVVbIr8drgnPd0IUtRg2D6dI7nrG4Y62bZiBv8Wky
9x8XgvTOwmdd7tYGkUyDojRHSmJ2EzPrW/iXnHirud3EXzrZa3hjO7dVnhBHi3zh
xnK8kc5z0ugbp4BMIXY7D1Wxmmz7VStnAqA6yvOr1c9g0EVviD7UUamWDm4mvL9b
8RU+o7hiA/8N3WZYIst9SA6ufx5YXQMO7yw+1YTOX4T/XQHeW2uI1wcYuv284s48
Q6IOZ9GBN3hvJzchPKOA63NtdL15i34Z1MFTbHgbQlrIvIaUTCLj+2+LlTCHEp5+
6cmL1W28UGHcq/aBZjGsmMofZIPu6e3QZtRoVsgcIXY=
`protect END_PROTECTED
