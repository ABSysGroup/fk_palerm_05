`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8/jgqw6NucRy9z2qRuzOoz3D4zlSSDbPEgEOdWoVjToUhSrmqvBR351EUaL0UCkA
oOTpPK+WC3Bdc+fC7yf/g+6/wyQtMK2rp8e9dPReISaSAEWnddHAO0Zkq2UqmiRH
7jIII16LbNBru6/ZCTDBLiPt1bHRt9SctlUGWQ3pWODnwVaUFhqdevwSK6aWqCD5
KEiM/7zzWAs9tFRKj3YpcuwavxChss/mSltHZpetplW4nEbeAlBszraX0APeCCau
tkky30hodvOlXRWaIcwTOqWwd37hWDjCDii7I2wzFv5iEzc+B0KSuxmfmarwWKKV
PUExkBrtAg6sfeZaH/+/+pB0uIPeWhbWNE/IQqSPWdXTmde/AIGHy6cKuhACkPQb
iQ8ysx/1bYszMlDo+xea+c7Arwnw8OyjGC8xtd2ZR4Sfdj4kkJHArLkiVLPkbKDT
fo2JDqB6I8fXXrhJDWtUQAAVTds1gwZIAee3RPKHT6Lsu+c27c2OiNRgI/1ewnux
XUQBMFXV56I+NIuiFn+pHBuDiuvzBEDoXz5FLEFb8S4JvUSW/pX7HBZ1LhMxPTDA
uHbpcCsdrUHruwJ4I+aLleq8Ce4MCHfTjwoIvkFHczWTbAinx5/eLHvrwL7+bsRv
ijy+5BcSPfCQ5VRV3hvT+IlQC9WYiKStYez3FoAkKQaVeoWMbgxIZJfGc93z4nvI
lHBnkqHioCEIw0CN/E8kaAjT+hjU2Qa3Nzj8enzF6EG+4GI1+O9qCT40ySC3ytHs
dAsf6WtBUdusinkH8nUyJrwbLRr0OHvvVOd0KQA8i4GRjr9fRTbRzpS4S+CTLB1O
LSV+8Hbn03qsMkDzADC0g5C7VMFiMZP/t2UIYvFW/KGIxqD2uphAzrluJ6g6NTbC
NB2MqumzgYPWD94yEuImKJ6OKOXZR+v20A1owxXp/pT0+zgSd0aTM9OWa26BR4N6
sqaz3oYxqZB2uDkkR0ihESpD5/3NGzxj5IISuKsdQWUphRqdMFmt8NFWvjpnNItX
BI9he3dF2M6s9qf6skMyVvardHxCHCPhZvSjnN8PG9xnrAJn6su/rT2CMZ+rV9Bp
tWDec6uTiSs2uVTzInikV3ZKvpZuui3KNfRcrhpnZvObiSHreGpboGvRwBUUzeR/
O4hrLP228mytUAKNWEiU+R05AaCHHjtJY9pvmoMilzJZ1SKKSIgk68O6dkobCsIX
1z9Fdsyt0S63VcAXGY2xwwf0wT5qg6s086r5ZqspyNiMG0TELkSQseWgjXEJ8V8Q
fITkKJQwk1P0xcUdxn9tquxDsfuXrSUnhXkPtxhcQivvU9YwcABoBM7jYHPwl1rl
H4pczNO6wfUArC4WvRoP/CaLZ/sHMUT+PEFWHc6shO+QH4aJfz8t3lLRQsQO0HgS
JWWMjwgOnyQPtlK9930UcNYq2jKWpOyhrPTX/+qS2U/+PuRXZjb3pg8gfUzDI+mn
JiQj73EVtFEIFN3Ee8eY9ELtZv2qpuknvXsKK158SSdXyDiKSUqTzfUObNE2qEAU
qlvDuty95b/R/xN4LldUWxZ20KLpN5dOyZzL1qXUxzAYScjbAZfW5AceclZ9nPx3
ArapN9TiAAEQOgdojtP7B5UkoekCgBDb5zKDOYSd271afGSzgVx6wScaXSszXIoz
y6HXbwbFCjj+gA5DYi7ZKFQnPEdirAeOi5GLerL9q5+2uCONHRbGySAnPaWkkr7q
PERPSUIlxf0rOxT76X3Q3Kq1L9/F9GTOKCAZDPz1ygliA5SCqMQXAqzr8pTSb0g2
q5tqd5K5BckgSe7RjYu/MnidKiuS0XqIDcw88S/avY1YoQ0eDMCYPqisSN3A5Hv5
x8aQLzEDfdV4Vpsa/hhDvJQUgIgLkx9hvFKXw/UwHzvpavXgnnKOHb7CoSEm/FKu
A30OLEtmRacgPA6+iwzmgykecw1F6Yi4qD0W/7Drb+vgdAYSgeGFwY4+oXKBSr8U
sB1dRF1jyZK6Nbfw46mNK4VmIeJuqy1CCms+ZhlI7rqCLELllqEosngcg5Dy+Jc8
HKk/jUSmJV7n3T9ODUHEhDAHrcbSdnfSXhBtm/bq54cPRDN38wqYmiTEbqsHjDEk
MAvE/Cs3VnXiV/ENdiwzytIqyYstb4nQzEzNvvJ0GkZstIwbuFvrzQx2XoEU9d3j
e1wPm6VYdNUvFuZhLM6E2QUhOikOxAMWEvGzdxiDGDo7nnww3fRWVrt9uL1bkz3r
dchJsslOgpFDXuho9gkbhilt6o1bDZTH+ixBFFr864C39bnGySAG9wn2oX/76CbC
cbcRHKWk62wvMsXv8S0VVckEk2Tw8giQikqniomUYOXzSlMveVEmCHVtsqwiBsrG
UHTP4PSH2/ohPuqUJ52R3L8HrF+pwnriuURxyKxhyeB9oX8PCwxVuXXJW3aPY5LO
yhvuby88D8F3aD1XWf2V1klKaGUA3smRVxps4GxKRDNY0hNhmg9spt2dJRd84hdV
Kh3B9SXfSrFbCkMGMA6FBMsfes53ztB6NH6bIL6N86zn4FuwbSmh+OYnkEMe3lNe
nffB2ULaql46S+j9b0W7/CiA66tDbX4st8P0qDagHi1hJlBQnG6TFxu5sKbqgjjA
M+nsJF+VDjsx0qSpZ2S+fc+q/l0RNn6+s+0YjHzbMUwpAE+8hBTiSCWXUFxQXobh
1DcLVUArZtpuvC4yV7oPM55smGKLHHgtAev/k9aTosDWi5ev3x+KgmhlPeq8OUY2
m9elPQNcBGKx1hxBCIqQcwELeYfyv+Ej+QEGkJ9gqY4Cydlyiz8h9u2bqlcizQ2N
PMGx1o/emJzcS+ngHX+ilLF/7yfBsTTyEOCuXC8hVL+gRfO8z7snzJQzMhq7gHVc
mwIqyh17n5bYhKXn5zvwKUFe+89/u9Kz1gt8sMecOKfDouE9ya6mO0tLOQVk8eSw
Z2wpaXBfvrcITrZdlavOrkka4hvM0L4WAkBgNKQQeYEFhFG5bs8PUWHuqmwi6Ggb
pd9R/saJSnTiJiKzaHqNnBTsVuqEzmEzHx6k53FD3xYp0fMyvU+0gxBbBpm2DJYZ
5pFlAQol/z6HG9qp6Vv3/RyTY3eOUM2a0eahBmj8G4cWYnHgW4ndcAn0hLhcAPiC
uifh9ji7s6FyOqrty81i0I2/kTNSwE2NNLwCRt75P1qjK86tbqiTPuMV29dF9WeY
MqVVWWHktmN+e4bznx4FZ2vOY1SJJf9KzxFMsHKTubzg7BifiGMlhPE5KqB/4eX0
/hgHYR985+Nn4LSAKdg8rPjuu4DZsau0x1329zCGVWDeZkCo1UyA9ecxtMbtpkFw
pIp0M9XDK78dVHEkLttkTUzF24inorPxucV2JgyOsUakL27Dr37PK8fYbIaYea23
LyoHZ6PK3CToJGo8r04OYpPpgJ/vjMTGmc+SJ8iudCcVknvc5KYfhvwl9Zhaoaoz
rE1hHmoRsw5nhSl3T/h8MzzdPT3MnlqNpxMABH25+Ga2E0zKiyAyas8m+Wiilf+x
cznw5WRcYZkHkU8Exdk/msIMKYQwuzyjKKR/GOjUrSJo8kmPmGRBS4j2D3dtTYa4
zcEu7euYsE8MtOFj0YUU62s34OKjVD9VPfD4Lx+Ofy9m/FeUGCS1IzdoGWZ+zos+
a1KupRxhQ9WDqayr3O2DC6ZiC0CTmksypwEGckC9AFBZ9qwvN45q9+dwWvRusE0y
k3Kpoe9I6ytIWIp1CFXPUFM+44T075eEH6kWFVgXXD/Z2GVKcc85V/CL9ybMwohI
iF67Fk6BZQM6fZ6bm3pbsmk9BvsohwfQcXoFJKjJeeVALiCknKVIPRDTZGiwyAgy
0e4ZOxtVsgQD/6fsp3dno2CIWeOEVz+xQLq1dDiZZG17jK2RP4m0vxz33Td5agjj
ZuUqz40SieXi8S96jayNSIDCRV3LF73ypsRF4YC8ozPl3/D01MFvsKguuca9xdtS
8XZjnblNlLbq/msiDxXGJDIdPjEVTVANnE1grYyRVA+XzLXNI7nEFy1cqQ1GwTbC
yfjNBzyhyRo64R8FRFSpdu4ZaGjchygLnD50esn2F+JnGlPLmNI4g9jZV7f5Zns4
zHguq6Je/3NSvr6sRr4/nGomYNRcu3sf+0FWZsFaGByJkIZDjTZpErzmA50GFoFL
sDXPxgGaSPP1T3LI2+wfUyIm0DHEx2qq2DvfAB5ZrGg27Kmo+c/aWaS24b9j/S0/
k250uyxCyyO75RcrVBrgQUt8Ed4Xg7FrcmXITkW2VnYMczenNbkil5yMroRcmAeb
Hw7/VaMdlwHEgk49Zb3OsGlCqSHOF2gu6+CjE6njx+h6UKG5nkKZNjTP16YJp0uw
X5HbkRCVcvbbh9hH5cQIQexncsfp9S/sVdQgHnLDA3dGlLOGX5OPi5OynQuUTz2L
0JLVtyx/mrucoRuhfOgmwpxVJerCz06Dnfy9UXvnHUqoBZ6HeTzShRijtW93kV8b
hdMvjIBfC/oeESBx297Brc1I9vWxOP7n91eocxbG5S8hl7z+C4sHnucwqzL+gVuB
xxVnlfHh72thpB/3Rm9jipU24vZ8O3FZDAFAe+uieNLmAVmQVNPvEXEe1V25kjFg
8crFhq9D9oQ/AKPKg/iWdc7qQ0Qq1Olrv2Zrt+FqfD7Pa0DduPB2hGvmgw69KNpG
HZ8JQL8EhYTYbSQwtCh9jg8zckppnE59kyYBNd6C6R5WZjUKDJMl/Kp/Mx5DFfv0
/ElpIC+BId3OLd0stXMy1WJBVaa15rPyoXc0xkDG8kkny2wgK8dWrxugAtnmBlsE
murt/pCpTVyzDeLHfES4UowmmFN0I1thR00LVPp8r4y3m2NUE3JdJ+0O92Y3K1kx
RG30sOfIoc1ppd0+lilv6FULGXa0RpPyNywBOqhN1H5nYSIrZ5oIik1xLn525OEy
rdiLqjhRm5xDjhOPBR7KFMxsMem2lCmugYyzWJe/9AASZYdzR9nJgbCQEIozUH5C
1dQYeseHz+OkZtfDzWMIslDMJPjcVEEkTuXIwJ3m5EVq/LfBYxU19SEgHrLaLHh/
RYhII6S9fmjDl/RCOQRChSPWsVYOeTgl5Rg1WLXX0o02kOfJ6E/mtCnOlPDq4bOt
UXTN9ZTu47GEhV1bXM0fChv817UKXr5GR0hrUVs1ZnQKeOxGLQxSe+RaUId5tr4F
2E59TDoP/YZbeI84j+bJ+UP4DoBVp7z0898XPjUhW8Ex6pmsCEHXR90VsI3VfU/q
+LoKGS1n2JO8FHgjqVw/luT4nDlL1Kv0umCiYAIG/KisP+0oac6jYFlIQ1ejIyDE
KmghYRmt58pFC+YhrECfq/r/o2yLGxSvEhhaoyslA8OBLhKxrsmOw/pXma0kZF0t
htJMgxjlCXpGwTjecQFVRmTcQ8zMP/1lAW4CWylqUhTShreUctknAmR7mtjAyC94
EmPluJazrbY54Aq34K9uiw9gF32pc6+cfeXRmrG30HYj/N3pTjz3ybxcPvMo53yL
ac6TNK41+NjI0TH26YBl9423MKCSfVvZ7fpkgqC3PgG+hPry5Y63NP8PrtQXDkTZ
cdJC3Z9RTk7Xa4tCaWSvmPjUD4ni7HVZscqZBfkeWPbNEPw5gk5EQroZn7V3uK13
f0mzxQgt2/7/nbcEOL4L/04IYfhl4oCF8bwDKQkvtHNcLelj6dVbKhCNrKPFnX2O
bLwBAUs9/yVdwPJ9UOOnr48cv0mPOS6qgH4Qob4bcyZmNDVraZurCcLyhhla6AXE
B4Zg+Gt64LMJjW/7UA3P6c3sGPn0CGn7TVp5IUrcWdnE5mC+6Weu3c2wyfat4hLz
JhQRpTa2PtAcA7zolGGrBx6qnE71NLSIJciDxz7hZ6454rvpimRIGWSbwpPIa0Eo
X0ds/RXkrAsH/sFg9tf5/jKWD9+kZ8oNR1hz0C8IrHM15F3BOodqrb+w8Eb7VTMx
Tp2EI5V/ttVdNutD0DyEHJSDwlMDj+PsyfKF2ZSA5A7tp4FzndItiolLRYMWglED
3V0vBCcn4zCmZ8UgixzfyvhkdgDcyVGo+IjrRVH6SWnvb1xXXq+NNzXacgT5Gi2S
7JNc34YT7pM9RfqD26AJSiTDa8ejK5CXjOvd9lG/VQ0ZPbK78LADskFUwyywALt5
uCOZVTXoatdSc+DqrSxbLO+zNgjdh3qzilJX1HjR+tUP6Wx3uZsfg0yNJ5FHCrUK
NnwtvtQeskc5+DoFV/HwMiFLDt4Y7Xv+MZw7cm1bpB6qxkW6aZpTKOfk3Eedk9qU
a6TYkAPjWWfyBveJKDS3Pfk62JeG+A3uNb8FqQvPaVYIbNn8FRyIMRWEgwYoSsyi
BFJnFrwCGz3Ez2jn9ypt6AtXQsFj7E7QT1uAJhBulNMSnM27bu7mDedjAUe09ttU
+7LgmqhxEAt3yfNUbx4Xga3KXmRoydAJAVrQE8+IEzVDkJbG5MkYWLoeBlN6hQ21
NDHfWgW6PF+t1OEswpkphMS23TFyBDZxyirSKx0EyRXK0be1/QEZ9cHIn6w1pNQ7
tEkMs9b0icEL/JtvB6aArVyE418XIA5ES1u3HtfFo4iE9EnpJgvSyVl9ESaF3qkh
6t3ym1YUKKlbodnHdDRTmGr9Y5yx0Z7rC3d3yqzHsPMorLOYkD4TSswedxGRA0ni
DcF3rxj9w2Kr9KGLR8yKPMPqdcxWCeWxCBy/HiFpiXwj4CqwUaTxi8hrDsw4ibSa
+GcQRSneivYABfPlKxa7IIfVchzZ7AxyPW6j1UBVpIKorCRIF78+0Y3XmYFgetr3
RsKFsgEpxJn+sVHlWTRRcqXRaWD6wC32HIqxoGl3Qb96JArf4ha6S8+ZCqUc6Oab
ryKsf7zMWpdJ0diK7P4pBkohg8kR5UOqGOapInujELmxezOtOmadkZeT/lD6mVC9
o39yXip0UCPWJ14IcbE390x2NfwnH3uCJxR6awCzwskvl6OBKSubg1QC5juWLyRT
aQMeEJ65JePceAPZS+NYHd+Od565hzrFxvuC92Ici+JHOMos2s3vzKtyZ0ZeLIWU
wutEnRTS3i+A2dghf6uq5QkkMAa4CDADWFgPoCFawa2xHKYQTOaDRK54MoEoBzpr
urPBylb8HSwCPf5i7oLNihMC4GJL89GqYgGCZg9F0dDA7PDIHkLQDGrJLntlSWM6
nvXUmQL/RKPcITEzFuCSFt3Sout4Jb/hjhLaA/7LfVVMiq+TpSbAb8uOW/WQjCdJ
kJxXIUh6mmE1xri4hRC9EX0cvdb6Ot0yWSDywRysERhA6NVE51juhA2IZ+WLyR2c
KLkuP7w6WZS+ERM920eNtJkctaVkQT1ZZLWtrV1lgd8UWlHaE3jowAlJC5D0/6BQ
F2TslLtYjs1FAtmlrJOl0FeS2hzzb0Tai4VDGfGAjFmJdF/VFaiEL68fMesu0lkE
2DSv0vZVzLsICPOqOapbjpwGVS/zGAtXmC6bVaEIK48s8un2J4V+w/TEsFNAfw20
00dP4u66g55ulmLPac5dGahy/XNg+lIZqJIbeKHvlhpQjGpo3IwJhlEQoK5ReqyQ
Yy85H8089WPsQj2uKVgYVnGEWVMGqD0nK6LE/U7SpKusuEKi3bKJoOqdfpLcoOgX
xnFZR165IvtVfA0MOsVuclWz+WptFa23ON1HdOC2TGP5P3Doq60lKiBhaIg4/i96
w/7q613tnMAmqOdKtJzJK4yQR+1w/9FzJbvK6OBOulC0QJYwvtOJkdwx4yu/xpkV
I5t7Vf6q5ak94Y2IpNSkpTIFOH6o341Rd5tmvkuTZ+2Dbzfn5/VQ/+iva9ZyaAwB
90j6499e9lqnNGFggxF6blNoBCy7CBAVggcqScRzbvcvpOJQwYZcIhYB/MnTU+EL
KF2vtIPBSNlbB2+KzRR8H6SC+qrjKfvqcUIVLygY/rT6g6h+lYeVitZlyUSl9I1A
R90WY+73TzqvKdjCesYkizXRDezdP5Hu490oauBZyPHfiUXRWp/kvohAn0pixeO0
6hkz3wvDJwuCeKVkkH5SsRb5krDyIVqrOTzn1hAP2vaRNiIXoqEJRym5DlUOYSJk
FLJnwaCceJcwl6GOHc9T6bHYOPSsh6ZUnl9jm4x1R233MtOoOU64deEVpzwmiTAA
K2NPOGlEivg3MOiTsAHtWzZ6LivjyhFGY/vAyBwZDa6uwTAQ6Pgz6VWI83P29l29
D1M8ICW33jw5fVjNya/p1EycrSIKefZRlFusBe209hYnKbMKLj3Ys0p2GUIT4Ohk
WyIMTk5luxc/XWQw0/oExnm8a9DSdJIPpUZfYiOrSc7ztGzPlg/HpeJokd0S7pRf
aGPks0PFFByhijasCZ7RDMD/uY64uipZDFG3L3XdYWTCsAhBigbQJYfnmUGhe4aW
cPSsmwVG1vK5nQx1UhT1vWZvTsTNgYuL1yTCe7J3/DoLAqenIX+9sbXbuWe4GUYl
conHBvqEbecwcueZnLeawvLzDOqMliieTuNkh/hrXCDDvevkwtT3Acyrg/sXEhN6
fplbGxHCdNBWYkrvkd5cBkpziIF4Da5CULdEXY+x4O4RE7DVJaSDdPr3Oq1Lb3Zx
3yareUixn2TJhT4fbR7Y70qvJrgWDsUFkF2CUQVzoNy5+OTLsNwlxJ5+20ov2tCA
iTQKlFtl4YNK22XW/m6cPdmQ8POXz1nmIKk5m8qSfFPHC0K1qzrQuWcv0B95C/O0
cqhYl2khKTfO1JAuLg4+HU+K0htq2D0hbLe/vLyJ7ghC1MDO38czR6RyMOTur3hK
JmsgBZusC/PAVRm1hFbncxd/3unG2YT+9oH6n2otPwze7curItTLKxQQM8H6UwvI
pDuLCaFDs+alrkDTQNDrYdNVRgeM/kas/QPtX4pBlh/1aJFW8GVFJfUNubTRi+f1
+/FmH8Pve0Khrva8kov36m5XHtsdxcPDBv7Uvi3xQey9jz1tXm5ADnCJYtRu19jD
0khcnuXFHfMc76DUTQBXDiiNaKnhlogRm8w0Wird0QeOqpAs4oaXHEXYDOZQrbRV
VnzyS5FX2btctYQGYVZd8ElHU8P6plDImqSqrc5Zvqvb3zDCFVNKTCv2hH2Hi+Qt
uVKi3C8dnwMXZ4d2gELmZnGnmAvYwynTbOPPVbENWx1rgOSEN8q03yZ9XPJNR8UG
IBUMyRM6l11gD2501eByGGo0Q1nCdqeD+rBK6crnZVbBZAqDEAng6ufFnx9gbYGU
uaYHEYKEHDnz7SmUA2mIuIAkQv2flcn/xE5UsoUzHZa0/uI2q3eDY+dVzy9tczz5
LbgAimz9i7MUvHv4B0K7w7eO7SE/mUovc/Cdhv0Z7AWAh89558NW2hb5DGgA3bKs
aGoC90YW+YUlPxrUQwnMvONdOkXMF/wrr50qxfkTwiT4w1WOw/UY5yAeSd0kho3g
y3u1k+DdJ9GwGomufasVBByOsBZU7YgmPIQR6jBNrCQw5oXN+YjSbI0YKICuFSkT
u8agNxjBQDW5L4gwUK4XvYwUnh67PaMdQam/n4LsgItU+xD1MHvIccqMhtiLOdEs
r5cyvIOIu535QmznRm5FZdIMb3dBGAVA+LfiE0SVw06Xx0RzsVxO7Ul7rpEozCGa
9SGcvwZfhnMt0gQPCfJbsnbVoiwx9d0otuMcnWRUVpd26PoGcs0A4GWzmMpR/Kv8
4AoXDSTQyoSWPwnGO0R3OWWUqTiYJBKE3/ArQNDTavOargm133vmbUKJdRC6KV47
hFNYoRCBn17FspNQzD7lcgohRO3ku8U5C9dAnv8mdyEyPHbxcB+RJlCq+++lvNS0
xjeKh6YFSgTaABfvpeXh7wGTKMCtI53F2MU/5Vxs5i2smrPB8O3kwo1+G3UtyxqI
zNXkR+Ro+XQEMan3shWaB2bbcjkxpMC/YcnGueaOwdaK+i98GoWb+INS4vadeJxR
QDxEtaUCYBGxKvuCNw2zhNMBZ+78eGIQP1IQ3eg+q+OoUKQGxo2fEnvTI9kIAqsz
/oAeCOBUEatAWjHuA1GvbnPfWuwVk0pFAX+vgvQmHrLXyt/CV68gl/SRcN3cpebE
MwNhVvUIPXgyqBFFAbpBPbTABmQ1GBa1nD2cZbbv/55hH5fqRGwwLx7C5o9zXP4v
SWzB7WMIUyLidA1Ean6f2SeJ55zuKltSr5+fDj/jopGQwM1+ri34MN/NPMIW/Knj
Ve/B22atqzwqDVDVfIetRW6ecQQmpk9BFCXg1vNkKp+e+MkOf92rKEPIxf/sJZ+A
c9pHPECHozr6HVSireP9hZ+rE/0pGwFX46POKVy9+41sgt9XMU6u/QKmARSug5qn
nNGsd65VtsEiLedi5S8lqHOqhiasHlh3xwnrJ4yTRwYXCsD2SKH18ks5GQAeu3rz
SCT5zYNi/REz/Zek+s0+V3+5a8gdT6MRw9TvYE3uoIdH/0mZctAJZniGwnPTvZ36
xJbwUp3EQa9Js5jnuPN0WYlU6eyG7lve8/j9z/wh/Z9N6fvAKQMwbcdq/kkjWJh8
xSv1Bf8b6WShIpBQpqiYnAwwdy7eaQEEZ6EtGEx8i1O2BH8aJN2tVUsZPcVAySsN
+Z3krtxOqu6yyW3NoP3dgIJnZ/Mds8CX2pSsA4bepHndFhgaOdFJYJzlN/tLpPqP
nztasKsVSu1GEZR2UIaHZLnK9kUjgJVrgrm3T7xNcvFOWQTgIlHbicgd39m6xsB1
o/9/Us/ohGVLQgizoOsRpnl0QTn77mR2B8rDG7+DfulWIPvnp9hCCl/I2nr3J7Xx
pEhuj/roysynot+raDvoHqWNDhrPyV1Y15Hya6Ox55pVK/YnhIlp+D4fn7ObHT57
LUk+qvv/kWvuQT+4kUpY9bH3sLvsRxhEDeB6haOQXAfH0I0NjSSzVIOUUIXfZVnA
OyVVDtJJmddn5gXljduuksxQBCeFKzP7pGEilIDLXjQAX7Px2dFNg2IzqWpAyzGJ
LIHPJXzEjmyx1C6Qu7z2Lv9242Mby7ZFzafyR9PPduHKOvm6AHg0PZpdAd2rm8uH
+fd01w/9YhW9hEU7+lTqojUUxszylLpXbbR3trJaVDBiprM7OczMQLMOGyARCv2P
BWVYzbMpp8nsbGIoC0k6uF+SQJQII6qPjvJLvnOZCx4EZROECJP++cJt1+qpi0+7
s5rVO2RRh02mZRcg2bNKWGy+edi4jCOzj9jTbUzwjF9EVCudytaa7Nh8knrcAbLY
6XLrvtCdUSUfwf5JCWXS4T/Iy73PY4Syy1QyVnRpgAQQbTIPC1ZF7EqkYYetvZeK
2XJN1bK5y6qyzh49NgY6bs2X9qJqfG952r9Unars0BJEyQ93R5HSZrc1Jicgb7nC
YNd8lvninvm4cpBRgCz+rSj2wtWQ/k9Sjp/Ly4qO8HY479yPJlB+fxzMU9ttTDqh
FTDEem+mqHC7nEkdEn0Ea+8HxKfiSFNz8eX12ERodK3og8iG79lowT4XNO38PBoT
qkq23+q+YldsSa+bOVoD3S5J5eBLyOn7JL88HmDEscznjOPJZfXW6+7i9yUgf/VQ
vbQoamyn+Y4n+6h3uXFg1woppznp8vOQgsLNr5v8DdB5tuHtduwkatAWdxJ09H6Y
dWcPvt9pGLBv1LlLV+Nw7UoWWP0LJ9dMOpOaD9JYGEpDvQoqmC30NRrEkvRfBHL3
+PmjVn7TLc4EvaMnEwIyDWUv5TbeTqQLZoZgmFMO1uoiXnVuQHZjco7ScGhWGiEU
HWeuWfiv4B2+OQC1bzQaQA9dsil7he8JcXZqkrosk/1OTZESjZD3X1mt5vLU3Inz
bdb55ET6te+l7aswnu96pKPQvenOm8/HfdtrIYunHdhc6jayeirRcZNgc8NCTm49
T2gPNwLAx5sfU9TXFYFDl8K7eHHJHCOJPCzyKipBkWXxndXiklodkDtt+1ayOuKx
mHgr3aoDWVagv3tpjWQP4yq0VaYZt7UQpgm6iUIO459TMoiKD37LBKfW4FvIhMDR
3j9elrGipnLqYbjBoBPIMJVdVg46QiMWtY/0FuPUsEcskI7EoGu7Ex8JlfHIvjd9
gwu5UfC03DBa3c/q2SIHjOLN7wAkl4i+0/vaI1PGAFFin+Y+CtofybTgTJrcUNPj
yOFsV+3y8RaVhFbASvC2cMWTV4G7dOUIgR3nhJSpM/pgW88+XoR1rGHKd22tfZEv
dHhixuXUpk4wxqvh4pnJBrP+xZeV2NHLp7nHLCe0/amezXOY88GRgA/cLT7AHyke
sdTBLyuoIbAIn8L6DtncHvKb2yYMa2D2JHRcmM+08oo38sJWDAyp51nu3ZBWnwwL
fqvivGX+T6lt+bLhfRVU73BzPNtNJ6zz9LvU4THRBBSIgU5ZhDAbvXSxcf/EGOBs
BZRO5gF9kl8/q+9/13HuBPlXfmZUIQURMe8l6KTtUwKpOzkcZ4NrXm9SatBRKkim
4Pmt7ucKo1biRQMYMEFn/N3TSaFbEe+6cwpE5Y/Jrb737UXLPsqTP0UvvHAz/RCI
xMs2HkG+HGz5hKNt8jXaembfvcfoD6iwwMASYgRc8C9bx6QWfKgDIQVifWoCePpV
9oai6Jt95uCN4VVk8DAFedEIh38l1iiZzH+41x2ljARcmzcwYmKzpx7teudA41n8
dZJ5N4JkqFfdPNlwmOaGleqip9jow7Rv1OyxLr5eXN0tUjG98gXBzkIT2CnlKTNn
mzbKSsH/peiwQiqgYBUfYPdmqz5bKfp2UQsNFvMCVGnjaXfK6Hdy5xRk++CSszwo
WLgrZqFPO+wvv/iq1I/ZZlQOg6RCgbjcXwonvOevkk5ZBRPEXdOCuZdU0OxCEv8c
g+oXvhY211RkanBmTuZMzwVphj43IA73qPnedtt4PT834RqMX5VaKOdpGLaUt070
xdZX5729dpGJDv3PlhGRH12FbpcrOYoJCeQXkiKykPHw6ZbRKaOvfDx9t8EmuFQy
6D3YqVZfoNwIWB8Mjs3zFzO1isYbl8aBwMDt6M38OekmD3vvspXdrrBzt5jF5siE
oRD87wSAT+PzwTk2yQaYiedSm1qhqvZ4KIOfe6ERoFNRmtu5hnqCZE8/5L28C9JY
/ggX4h4rb1cN/piNiK3/vOf6c3EgkbRAXBaJG9vH8ZeeMDpy4bSrwa3AQO9eDshe
lVTumZa0/ho2TDrV3viGi95siLFiedCKMjGUveqPsmL56rOqO2VrE/TBcvpbFcxk
YCaJ7W8Sa2g0D4yPqnOXD4NVIjM+x6AlSVXKjoBg5ECTUPSbpdYCIm7WwlXQp4vc
Fi1Yy4CecDdAv4rYB2S68+bxTtiZZUoj0O8w7MCY4e75YaQST/UzOZM8XEfxiUAi
58KN+CF11w5z9ZgFfS1Ae7Ldytx+Gp28cJmG1z7aLKVJgDixwfg2Mfn31z4BYd4/
LBCOZ70MJypcI2G3PPKAxNJxw2DBsFWO1Qz6UiM4ggSKcVZl1U7egHYPfteseYWt
4gH3aZxsIOyG7Sc9bcT35hNvPnJJ4SMELzcLegIw9ZNOw5570M+CRnsaqTqBh9AV
t3tlmafU2ZZhUDka+b8PZrepVjxaZGxQsMWyZqAgAUut5iU9hZpqT7L6CHvwcK1U
AUlSUG6VzyQCCBKCccjulr72fUozCwyIOMdqVAyyPHMaQOZOTKHUOA6Bq1dgpFs6
gkwm0Dn12tRqfOCOrIcudiOu3qei/cEXSfFSFpa4KlX9YDf8Q4IgilCp1mMPQwKb
PBngJ9nu+w24kP2LOUuJGEg9x/UiFUGAUC+GE7L7NBIbgM6igEBxz0Xugc4ICY+T
2gBtU3WNZw/s3UyS8unmpspYiMO+wTYSzu/G/uKC6ocuglsfeYmT6sYEQwqT7d4F
WYPs0gR+bxTEb7OosxfLHZVXLYS3vEu1JG540xClFBy2+mQsxm4jqSieDCHZXeOF
J7sRb4UjZ4FSHSs0veNEeYeYK9x+JL7WLG2HBJJeGxoAO/AV+o6M86z6U9xaGvbp
j2qljxQO/NQG4uSxtwAiMdV5SpO7r1W6HMrNbBgZFsXFhLt9c4GL4O+CG4tbBo/J
oBL2/+8xISvc34baElRre1QqxIplxtriV7RZSSQFDxe29dT873pAcEQvTJ9thpHi
EOesFUpxo8j5XkQP3VZzD3/GauiUaWpme6hSYlUvK8ia1AdRNgv+U+b0yIreZfYN
UMOHsJussdk4bb0NMFKXMUV6SmOSapQvrOD+pZsVp6+2udt8b7uUr4yqPBmqlrSr
FiqZ5PAUotHc3zANDKmh8EGcscAu2wqMiqPxaW6Zw1r2Hi5NZJzIPHW+G1jf1l61
T462a/Gkkb2YT2yUy0MOkbLnT/hAzTJxKef0qDXMcDdlkM9yTDudEtN3RRkD/UNP
2GhHaDzvmSvWGI8tqzYuRrq77fh8eqUL58EatkzCA6Hy1ifB9aV9dUECPl142npR
3Rjr7HIuW/6VtDivNg4kvIwlUApRa2ymBT2wPEs3ReJHtlFa/+ZYX9/ZRZnTa/M+
ViIdODDepPFGjLsqfCzcvaeVUvoTvat6YZwjoZxctKytDBZ4X91+BxnkHN8i3K9o
VNgdb2FaO5egJ5DTZZ2R12eLkSREkd5H4tXbkjHXHSmLdZfO61aNPZ0Z0AFC3Vga
qXOfkdNYM9vMW7+c5m05j+6p5/MzF9CMzca6X8/Hu9CFFtgYpZuQZ2NIsJFP9TFI
hi9WHUXf/8K9YTDAyoR8enWh+QC+efLkFJbEezw39ppb5boJy+aAB+V2r3INkHcC
flpATXSVVr0xkQyzleVTcKD1zKnw1DaYR9/8+XK9Wv+nJVs+XDY58bboJsD+lt8y
4NUersNFF+g6h00yUQ+oxTmwMJmzBmnU+whkZgBdQQto52v2tFTt6OodRpGwzJGC
oOrjC+xfj5CozCBGyqM/r0twL5FOIs5vLToozCJ2C5SVxmZLbEYyQhEO6Pv0Qn4q
1XlzzItSVRuRgxeZcgFcwPGIvnm10fPMPjeE4ScrVX2WO8+q7b1mcXA2xVrSS1U3
oAQUxlO/YXVgSIp4/e2+wohmfaA3t1bmZ/RtOvKn4wRiFrXI//dL3t5i94Jfdtn2
oAoWOhVCOu2mC1pLDgvhu8M4jxHXpmSgVk+M39zcYrNTn/AkvdD9r3O2T05huE8E
aZVIAxShftoLkBacH8rZLvuOGd8g0/voQ5APy7PqL7OH4iz9p4kNL3SQTP7s4SJM
IZgLkB+TrmKUKweh7lUw3++BI1ga9+3oiVHxcN6cnDvR+rVkpNFPClpcV4GQKtIE
Eha3fk1hWtAeiXpVaEekQM7Wp+yTtEPxmPtj6Zk/TyEs0kBB+11U/hyQOZW4lerA
CfPD3I4fi1L/6ew4GcEK4AAIVJWcvWj31QyWfEV2kNlnwNp6Ksdb53WDQmJzxViy
V34OktXv3zxMTVX6V0hQ74jpTObMduu6+b6kp8dXN6wFoOKQC+9Yl0pbA28h5Vmx
Od9iYK8fxP1Gy549Ksn96qroRvQYrO3T5FdkwfUeUSMyknAmTy7gHrlJGbiBCvL5
a2VEreZmnGqEvHouAEP0uDVs7ub9/4KwE486P+SiWeSeeApFYR80Ou79nHYxPO/i
jli86FHC4kWZkdfFW9RIy2PM2Li0M4PSYRLJcGpPmAmVVj2ibjpufKtzoTX4Pllj
mATlhZHhYt6saPHni9acfI/YRxwqCg3SngPQyjLnD90AriyDSpaD/1RIsk5JDbZd
3oPhdfe0J5onIS7nMjSc29HMMRnv5rJjA9VbgqIxck1e+BLSEnpEKm6eCDwZ681K
Lu/mv2WzbHIP+igsK0oUNcixSoePCuXeGaugGR90sijJ5AiCOpEuKGmYbT1HChkW
P+5DJmR15/H/y6pO6ve0zygGd+O4z04AMZlI4YsxIYTr4NxGxr3YLHrDP9BfDPvy
H8U++AkkyJ18ZHN8f6sm09q+yr66+HcW1+x/viJxbUeJUMg2cWu5HdK61SO2FSy+
goji3aS0sGdA1W/NLOmY/52KWiQO27go85zJHfpQGDyGBMzLDTTa3xGZOVu3ztM/
KMbFJO1v82U9Onxhczze+yYfEumVYe7a0Gz3f1Ot0JWuhA1cHqIYBnj1eiikuot7
2DGOVALxbVXb9unPXRlmTLjDVIOj9mSkqBRtbMOvfLRHMb935MCGCuPA2ySPqIT4
fy2sOKyWsDSZkr+vXx8k/mWjp9rWnIUSyQM5w/DN6oBKy/8S93GqW7SI2o/9yqze
/PHKoC8iyRneSo6O91fPZ4mWqYDOvdPgcrYYrihSSuLu7bGx2kDYlkO5vaB7ZL15
Pf/YNranm/lvThxVq93GE2RBPsUTPnPWxhcxLsKMa8NOVgQz6g/C1JwwZnGDL18d
xIzqpC1agYSgeYuvK/gVpbWUX0ALMD9c0/3vMyfxaUwwKlLsgMB0YUz3loH2vhfR
Z9CybRCJz+EixwgQFRlqSiVkU7hQENbsXr/+aed6aMzCrIxZrrS98CGC2cv1+1Py
qdQTy0+T9DCkdtFRWv0oC3hky12rHroiV0IA+kmq9VJLA1NZAg3nO+Oh83Yzi/HB
/RXRdLYCVSQPea8Y8OEtUvK9bombZi1JY+ujX5JQ/eGIp+UV8PRnH1ldldjtJq3X
6inQzMePTZAg+bBcwny5zQdlI05UbH8HOpuFvrA5WAQrcEe/oqvb/b0I1oERPlU6
UGoAv/CTBFq97pDsUoSRGd5VGbCPpNHe5QPmboCwt/r6v+Z6G92wRQw2xR7Cz7i1
`protect END_PROTECTED
