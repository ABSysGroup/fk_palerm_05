`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q51IWzMcYKjsHb3qZCqYeLLOD21F8FZ2mAGjezM+M/l3K4nWWol7mFC55ptUNK6t
dO3iXTyhusuc93DofHbsl7jH9vHxiPXWoXEHznQ2spQdJ+4U7Gu0C1EsCN6dE2o2
Mx+zAIXtFAApSO0UuEEczPRbEqBScnEvj6EhjKOJ10VoghUvIX+CY8tCeCvAICxH
iYhw1tHlGDb1FnPkvxMVJJTGiLPPzBDFHpTD7BPPbMUqEGsFmtvP19gg+vcAt4U5
wW+S91Rg/3bwsB06rKIXxDcbJn/ACkpD8RnwEW6mjm774w8Vway0kSqTPr+RQWga
81e8VfctjFUg1aehKHskkD2gs7YZ5VIM7OJsUJlvtH7z9Zuy2UlWo0A51n9Flvtc
4+rPLSBiUuBrfP/KppDXIqfWF8hWABbUF3yJK09f9dTvIRr3sYBQHl+s8eWHhdFs
Uwn882Dt0gVWUeZqXMfGfdNJJmrR1sd1g8A6HHxmaKI5Y9Pf4YSZV2v1t27kdpKY
mVJYGMAKAIg53j3GvHHFOEkYMkohedBz5oIp+nJ0vu7WrdO7od6Fja3HaanLozpw
RKR6bk4DjTW7Sd31Q0z483XHc8EoFlAipiY45IlW25eu1C5MB7UuYGAz6n9DcoUo
TQZoKhyxDXXSU//Ulw/+LSM4v9xrB/igzqVIVdWYNq/iz8voyq0XcRuc1oixkEfz
3LlZGKcCDs+R09o7NpmQgv5tcK1k9FeJzPO20noqgD45FxUYZiGI5XD1bbc2nzvq
k3dVGqu+TejXIepqUILz9mK7GJ7K5Q+q9oy5tsgCgx/Rzgkao7v4je7fCuIlWRhY
e1MVF4jcJ/SiZKpY+TFqVvEeAdLV0jcV+sPGrirXwItm3WBG1XmlcMW0iKLPOP8v
kqtBvbRaB8D2uen+bVwqMt+6O4/1wqDorFKZ4BNANJQaNqzrU3obdXi/DzXMchQx
rOA49qI46vt03h9SZ+l3Cc8Ifdbs5qAFXt2SZVAju32mpSQ5cmTJ0ZdF5TcHgHQJ
VwXXcUajwjSJPCMc1FoKk9LALYcWKkmHno+EswI4rmrSaYWdR1U2bvdDHSM/tOu/
5y9v52VQ3nsGMejeIs/5rxuJnRJMf5e7YaIhkLs0A+9o8ZLqow8Ky5yzAb8hlTAN
0oVnbX5VHRfplaxTysFwzvpcMt0HRylSbMtKO4aB12wyUH6IRcA1W/DNcHSUNcZo
lnx2OmD7Y0gLTLFSAm9SOZSTPv40mQAVw5ypmNAdkfL6Z3221UldS/FM8c5USBNx
Cft0Dh2m+ZaqDm6ZeR32m94Yrb8BycPc0DTOWBlgiZFu8eQwA285xODCu0sbp0fC
oO1DGXItXftnnbjwBdpGv3keWBywz1mA+VqrhQ3qGgU7QE9XaRpdnb4UbRQ/L7m3
dYlHaWb5WLB8HAFICNhU1FITdxAUCv8aUrhQR9YT/at2FHsceLZH7YWJ1yprvKmV
3ffG0uSQCiSHQo5jmSKIa88hUjRLbe1dGqFsVHMZSdavZqYjpVcV5S+DaYlNF89r
G0XA7W1Q0rV1pvTwip2nkAAUA5HWUMeeWknThjAx7yH67gNSsM6ZohdnArUL1NOZ
uZMvK/w/qWwiUKijsDvFXquIsng1VFk5eSXeO29mSnvERePVwSF7/gR6O5dRNkpa
1doRfpuK2Tim1CuNY9ghTHSmSGyjScQJq+g7/v81AMKExT5vpZwPjRfpK5WCApa3
s2SBthTCoHP2pr3KyX5QpYA+OvpOP27TC+uTSfZCBsvQUMAHK4Laoz0LT2fznYq+
v07f2mM+eVY57bj5lxAKizoFZKm16icwFTUnZYsq0B5BOJztPRloLVSN9KR9dNaG
YYIzHj2Y8p2UXjLhNOYmAOu6BiJOO0M5iaVODpUHpMAjIZ/axnzPhbWPbVsA6M/A
Yg2HUkutPA2mAiiijMhthcBy7FpIomGZBMRiFsBuZNdMM2tFFvShNN7F8Kvn1JHI
kwvb1+e/xOXUV+LUh209Z6lSxxJHSkUQOJTuG+6UzIqhzIeYX1OGlV/Cro06h9oM
J+HH1k7sdYHHA1vADVaL9h7KxarDP2NQrW0BLQW54sJffarRsrnW+Vp/zasWsjq4
cUXTo+dN50DUd2jpV7mYoV/XnzgWQAAe0HBxunH5FLjHe1BMOaDK91ff2Bry3rn3
B+qLfJxLpW2cQXYJzm+I4Ztfd9V9PQXgEhmIN5D5L3R2ipW7m5ctNFv2T4yRxgMG
nEfqnuzyXe7/e/RRuVM1OUy1pGonTfHww8AjHcJZM0wScHQw2VlLIsDtEs3MDnXp
RbrPiMaU3W7fc7Sm5xCVHlttgjjsKwa6Vc3HYqfI0aLc91ptFH9AburtbBuzg3Xx
KrFSRlDWPgC83r4ptvcuHjnZXxcuE8gfPcvNt7VwUkiRDb5U6GrefL4XoKUxEnhD
wftFAErtIgmm4i40F1G4pg==
`protect END_PROTECTED
