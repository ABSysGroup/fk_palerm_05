`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4x4wQwQwjlzxCOSEQwc8N0q78a0Mui7dMhhnvUPnNPhQvfB38zYy45wzW6eiJ9gz
3AoMYYBPxegF//RdBR84jIpnjKpljjeKgf2pmKKdBOD+betVIe8rZBrFwuLWvm3U
vYgQ3JFgV0fJDTEaXsXlXDt0SOdu6uMYIJKj4fioFbBZ7s8RLTiEhdB7UOUz69M0
Q4BkU5ILoFekEfeV1f+UOxg6LV/l2O2QvucTU7ICzNMTv4YJEbhVEAWJU89kjE31
b4hgl8eUkb7l1mIz6NTzB6x2jxMdRe3KU6/bO0E08CQ1eeSSFWeBCkDHqInjWQhf
yqDcCnSTgDTHK0CMkFD7hFbUc6PcpbjcroSKMTpLZMLoUVsgNmlMXqsXNqepNwGp
G+PszW2Jhmq/swsD+pXwOeOXWWj8EfYpY6E3Z05Is89fI6RDW7XpbSf/m0+rvCPH
7K0mLdB78rkVWYlIj9z/cGxTP2wMpORzzHWogyUfFF0o1PLJDlqKhIE5oLbIGFDG
rl9lhxKQ+8gqCWKumU13kgiwhI+lKh/OUfUfK9+49r3pSzijp+Xm6+OYHQ5jMktR
EHulR0lTQrU5/ZhAoJ1tCti4GGWPh8r7MvHN9Q5UuDMyWE08es2JrDHP0o2qtaYj
toN8s8wkQkbMOjjwwtHxAPaPHn3vr2OTb4gmVpxzu1Y=
`protect END_PROTECTED
