`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XzzNX05yrSw2/aDa6V1JJ0bqA0WNwcutDL8NHZCgVnBIes6GjuPCz5cGWkBA3+bJ
3MZd6Xqd69TrtsTCJoflI499rGjheFUECF9Q0qdzRjvBE6mAlqh3zi95RkYImg1x
pIucs84VdfJCmIzGCRImPwyT1uy+MvOAcNqhEUMQ6pHXXL4cT1DSPCUYQky831Uy
1n2CGmv+KXtA03FuG8mYzs6AvlmyCQ75WxUNwYjUZgPgF2FNAwun/mFFRtO5aZSj
jyw2AlUV+YOZ9/0loYdYx11uTiHxJ4S8VDdPl7V0w1AfLSkRckOzRvLg9NbDYZmC
qIt8KPMHOd2zotTFhYtkGji8RV9LQeR33rVFFL52BufFjEtFCN2vAnb61iiGcPJk
ARZxFc0UEjRvxc+4wvlq3Ui7PvOP9rAMaPOdfjRVYa5AEhJTvS+TsA7q37WTlGcA
jM7NH3NyxFzuGeZDclf9kKVfcMBqaG+sd1nK7tuAU4PSFO5RSY7eUQybT8KJncOf
AFk/ExGOFb3gx7x7213miLSMK7fVK9K01OHMhv1BWDbudTLeAaWkP7Ywhyok7oy/
OKDPTjwYG5w6Aqhc72oCeoJ61WZNdn1PboOa7y0RVg0qO87doI1xLqlAP34VI5lY
X+ffri3TligVRyBVIomLzQyh4bnugFvHVQcUheLTuLPmb5Nm2x3zO3KG0J/DlYXS
sgcveuWr3rFQ1WE4mNrZmHR6kK0zSklBzuWjeoHSnReoDuG4fZaGD4C0VsbeRh6c
XU8oXc/74jiRG2OQ9UblWIXJZJlfIJejJXi14jlCHvvyQ+DCzI7Jkr3Fwev5A6Dk
uK/h9tD8610E7cBHrkohRG33sjyb9Gkm5+m4pdsF5U3SYn6OZTr69smF0Dqu2f+A
18sGvuKotaMd20B7ub3Hu3Rm6pHNqQcY+lh5GcErD0TioRCWiZTu+zDITZB5NbUP
hvlxJ1Rxw3QH9m5FXmi2unXS1DCE1W65YQi2qNJV8Icj1p7HRjbsqoQP9sebVp+3
`protect END_PROTECTED
