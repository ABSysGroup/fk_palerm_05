`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FBn/Tz9Kpo+4Q5CG8ohufICENTUTAGRdyiGpiu+ty0IEvmXvwP1UTzOiFcEbUi2J
bVMpqO5gBlQsYqhmblI4/7Mn8afql9PjfOjifU7ek6cQC5NcJUwU7EiATxu7030I
HxP1XkmcJR032PLXBzR8fJN7Dppi0Z1ux5uHEB2hEzB9ppsF5hhgnqEMmxxXljoZ
3GGtRsZ8MV6thPEpahgjwNRd7H2crpMdDxswiPR1BVpfbVZ2sx5aF//T6GjiKZ8x
er7x3AAUHcY4j+2YfMPRO1NwEUfEyVP5Dj/Dk6wt7dfOZDLrnE/X5Bk1EBBlbIZH
CVyY9aFVKjDv4ypFwBKZ7iJjCvvKK6lMNW5qrTOiynlQnHmryaEJW44ZZy0o6Fiz
BHSROgm2G+IEjTWTJ6iCLg==
`protect END_PROTECTED
