`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BWtpMLf3+UfJfsd3PugdaAFYKMcrn1mllI9gU5dcWxEeVLtuI8B8ijR22K1Qia5I
UM5WPvBRQ7NOMI+S6nyIFsc9hf38lLd6MVSp6PWAbdYtVb7MZNdoZ5qHToeVy2GS
KZDpAd5mdo33xQG0S6MzoMuyYYUtYRCfJdMaexr+7EaxNiuszScHld9zgAaW6IvH
e4Z1KylPFf3I5EdIJRXdMrlOqKbkjDVwlxVflgZzEtxCKL+wmA7C3TFVghwwB2UD
fEKgmXzzZGE3YMfZW62eyyGz8VvubdYvbJ5QlF07UDG05OL/cVcjUonlPtFUEDoQ
kqYksgbhHOCSQtRgEk2trNcgA6wSP0V1VACkyJsaqRyq2yABGhatTLXCt+7xcLzw
GVofmYl2evSiphmfN1bH+8VklukyC9UIId/eiEG8A6Rsb+P+7wOvRQW+FQJ7bLlG
42L8ThJl/qjrBCz/gvkeHMvhlxZKf7dNtxzWea17PmdV1sPgOW3rpLQr7FiT08JC
mE9FaycXqmJuN2GnfCiedQ3rHy12RlG/9msEFXNuqsyBWV7Ybo5yz2U+LVYpRF9L
zZeQp8trtGj0MoqEjjsVglO3hGTxwEP7aAfiUUcvAl0/3xEmpZXkPFkS/rcH2+HC
MtKD76UX78ng1cNP5+ulmcMEzPi58YfXAcg9LWgAKOxobkFDbsm9tAS9U0u+yik/
CkqWP6V8TRA5NK26L5gdpIf/XJYzBGBiuIx8kxfSGONfTEAZvjfUoupw2s34q/wF
ngI/05GHIkrC93Qt8SJF3oKlqF2KjAja2/7Fk8/mb0Htblb3EdZt9/Cpc/GYzGFb
dRjeJikYwmx5fcUxl6PMvKdibHM5iu4zE3RfC4W3f/1KSpOgV8qRCKif3olrIeZq
G73X7ODvGxVtSRgjpg0HJOGbj17ecrRh119vJgIKID25Jiesf6p+CXQsVGZ7SxhA
MXP4iBy+7NmTuBo/+/ryKA==
`protect END_PROTECTED
