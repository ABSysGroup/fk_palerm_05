`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hA10HVc1RMfkALJPbTMtGcWw1mWAxxHikgdTmYJ8XJJq4qzwUJ1X92T1ADe0YmLa
vaeK8dzOtDsROmlVG/3v4/F4yeDIP0i2QOM190npq5DR0ZoE8hkoIA4RfQIVR/t/
7K73AzjX+Xs0LjJbekp7JEvVKgwnuFSPAYXv8gsvFwDyrb0hEd4cfO3XI2fbm29P
Zo+mikEtfLNEjYLdg5ftw5W2ZZumIgTzcB9D9ruPS6r2khd4BzU2EfJwkX/p4y3G
F6kIA7MgF3so7k16pEN87RUOxwtgdDzAxCZPZGeTubL8sipJmk4GkHHnPpIaYpRh
+lB890em5ZKEcQt7GxsSpM69qgvWLisqqWJwzLFmIzCxIy4Lj8dIwrBfTNmv94SJ
+BRjBphAqlsh2q+4yXhxNrR/wWG+iJaNqw9KtmaKwJM+1INLA+KFLqPgr9ni0cSi
ZdvarwCTpUOGEf9a7E7KwYyRMVb0/aaPGIi74TCwCT9chMgTG+6t+DxXCf3W/ON5
tlJOqT7JPGVuXyJpjrUt/LNrxd86InrfdPN3HHyEgwPqh6W6IM+XZ9TrSnWA7KPj
2WsRzd3vHO7xPEIXYqWD+4TZiM9fSXaUFIWONG8MIo8TrEo0gNqbjMoTLSnlNPvY
QS8DBSCaZJLl59kXhLwIuoIEdqo0iUVZmO1e8Ljb+6gUM7votjZIzaMC85ZrPyyQ
E8vJEzI9i8Tmwk9uEIw8vi0fDz5WdSMgZomWb/iuruLM7ntPwAqjICNVRoce77KU
oiIy+Aq4Ut4vdOBx9ZqaHbJOmWm+nqAuYfobW7+4kFH468wzTdgtmpNlV38UNN3Y
535AUGLavcLT7Wmti8sH9CBHT83y/WkFMXdem2237C1v/4x98BJdYjYX5GLxS8Oo
LM4ZXnG40l+xsY/0IDZBChhsj00P4hyYH7x6w9rUWsYyBsTwOKjPpb4Yu9DhNIdd
xX11gCDGBioAkerFYPLrHXPE7teYwZ71PuysERpJ4r6MSQZUx9tYZ7ELuQ9oEz+L
XLanO2Wre3qM43npJscQTe+bmcK7wp4pDgK+CwM/s1JsANEgpD+sS4RmhtGYHD1V
Ls9/Bh9v19N4hHEFtF4BrDPy/UMVh/ZF9iHy4ANTLRJQ7UAAlU7fBuhJTKhw4Y3U
m4OGYU2pWnFY3WJkx7zM8WTsc/O0VceLNO4qUPySrt+yRuZAxCHObbRJXqeg7+pq
7kSuPXHkmW1XnUN17cW4fxi0RQWKUQ+gbHLZ5nh2D2i0NXE4WmPBF/DFKhdTTnD4
qQiqeduot283wgIRbsDD84kPY/0drdZbXza0AIK3UmBJUZC0HqH7SbJ4a2zraE1h
AXNZunJBQSxb4LTJB+507skT3+McYj7FLQJFLblAwPIDODecyFQrcX5qEcwnq2CW
gnBe0JfDgJj/SUaQuYy6QBSOoWbbPDg318gGm7bAJZ8RwMUXFumpHLpCPV0877JM
mVCTbPq5f0DEmDbH2hVsyzlQmzOZ5yxmJUP5kX5WJIeQOgHx8A7wUD3IRDFZMYpT
9CjXgG+ddSLaLhvkw93aAhNtK8vltyCnzIMABH/nyTYjzpI2b6Jrl1xCFmT9FXWV
uCBuVgu2ct4eXfVx0qdNV3mmT/jOuXoyKjsavkEZBSI1Ns/GgeMU4CRJ4ZA+ZWcQ
zB/D6jTG7nQaNHb3BH/Wt+Ybtyu9ljtPjfFL7nlNDlpYuF1JA9RLDI83r7RRdlZJ
J82guze6+nGmN97ZuBUkIjEFJ1HSpKYGfgpDAl04V8obgJRoJQ5FRzyd6SfP5ltU
LaaZYx5xVGXtW5mUe3U8nmRqSCoLvV3Bfzeb4dyOT7PTiA5tP5PpZ7mi4Y0q13ow
mUkt5THgmQNXl2Dsi5bh1+EZ+qXhabdlUQESsYyfiVz/oONxc7lPWK/FtbdD9JQt
iG+sv43yumNAlGWKnyZTbQ==
`protect END_PROTECTED
