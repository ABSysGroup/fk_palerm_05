`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gsafe8ui13w8mEwz91Hdw30NagMhtLrnqWP55dW+4JsgudewXkATNFhNbZp95oqs
H69b141myGIIfwoJSBmqQyKX4b31EJD3vK2m5gu+gg6hqMDy8w36qJlrUdVBS/cv
VYCVj4IxHGI83fKvmkDwEJhGeEBugcFKVo8V36zHr0fayZj+JFenu1m2nfa6wBIo
CiPcJWyaUdM6NVv/xG3PcYlViRFIRVA8KGtNC8ANYCAON1Xo6gL6SbgPC7WYjcaG
nnWKJcc0+GSmoV9BNZDr8QdbhmLN2o2UzjzuzA6KNW0I71jpE2hOGYlE/yZLsRyu
4UJS549247Pn6AcGSzcqSnTkoiUYAS7b7Je0ZQWr4nG+vjcHGz4AvUtxJQIpSNEA
0SLS9vu1OhTTqljrlSdhODXg53bhThHAMEULJxQJcS0f3Nr2O7LoNDTDWMVCtYv9
gMNsf1FO6VCVzV1K/kxk3ss99QTm1kBUOvTT6gsf3ecWXVOqwzqpdUctFHJT87bo
FyGi1RWvh1nMu+/Sr19PBFTrgDrRr1gBzfC+rYc4952Q5nZOWYeHgVke1/P6KVB0
ioj9DEZsLJi5k1cyPmIZVztpjnuneda8phpDjV7gQ3CcbtH7C+gbZ99um/rSFTQl
UlA7Asdv+0zSJ9xZml59Ew==
`protect END_PROTECTED
