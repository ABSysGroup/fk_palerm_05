`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
thp2kEnbsZgG3LmTU6W529ftjyHcFlbv4RTM1ZgepGTHe02YedvVbnlc0TME3Y6J
iFS0hmwO84HjYdfhGSNbUI7vNO3j43cAIh1Dumlj1wcsdNikLYmTrKHsslwciCD3
GBLSJCqQAkynfXsPCEvA7cq1oTXBPtnCRGkyloQa4kjRBL/TNfKTqH8wAa7io7Ct
tzY/26mXFC858+gr0DeLX6uUfWt8FrbqOCZwhq6rpCbABfrOSLTwWs6G0P/nxXI0
TCj87HxLfkPft8PsDOGNS0OVoip4564EWWFPmw1+RyotKcqKSrqdWatJBqHiiy6P
t10by8ur5mSYKFurfxjHSuLNoT1Xsy5WOI1f1cqNtA9AeKIXhZtRD3NYJaMgxVtW
3Zmqao8CiyFgTRs3CblpGOi234zbw341TL7BgpVxIva9FEYphoSPFjHsMhrS5lhe
oerfLvrc7J7GNAcdTwe8TxuR51EVy0a3WONUnugXS1BGLE95DXcMZHd2rv3dyUTA
gpSK5q5E7aFngSL/YFEYA0ltUcsbchKUXqICFqLxgSgPFVaALQshI6PUVsqLJYMV
`protect END_PROTECTED
