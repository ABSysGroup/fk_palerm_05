`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p/Ky2UVbYLQHy8eNIeh5sbeq3Uia1k2HNc+1nT0nXNThPv8mKRfRiTlj1KnpthkE
cASNSUyfY6I8OMoyICYAslHyEiP4fGLC38tvOlkdh5ONXhYlmIO3Fsj2GYNLNPTN
jniPIE1KJAKJB7ETRCyyszPYLKOphfWFVS2Ljc2A8pTrm9YGGaLK41FGeFy9Wr5y
g2ecChr3bFyu0lAwu40olrZGWyLdjaH2exvbXuzMfUvCstQ7TsUj2CCBE4H753jM
E8vrYa7kGhtbzk6Q6fyWlpGrU7SNHzNZ7j3YKvtuV+wLiQCOb59htxmsSwwP3Equ
3s+tZTbpcFazKNF+snkLn1yrHKX4sDmi1tz3RRc/3yp7c7TgmUUI+B4om9Cgr5MI
rX2FKo0g6EIKGzU9pdeFFdKe7zo/OIco9hd2cS8Pjqe65iF1bB8vODVi5mzMdPfq
Z0IQlZdw/RgGbj7u6FLLJeSmH/YsLJ2Vwn0aF/Eu1LZe/S7ArtFGsTe3/xZ8f/r2
I9q1QowPuAvcRLke5UYsJRa36E/wwtnq+bkWKER9QUYpKweg/gbI2eVmCWy46ooH
UT+54FZkjidpq4zuCuv4izLO5WCaorDmJcwtU0Xa7zmKWBN1ml+UuB2dMTQc+MHl
HMSZLGs19DOcLhbntSt6tw==
`protect END_PROTECTED
