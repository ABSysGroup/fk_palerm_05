`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OCCr14Iru6ODme5kuzQJbwpL1VpfYQKx/MKW7z5u+UB1FJ+qbhzwm+QFALM3GPKB
UOfWRcSstmwxBFlV//4QoRH6hcXz4XCydUCyR6R0Ri4eUOYW9NkYa5ACR2rxZ/gn
hKX0lv/lBeDnFGBN9+AhuAYXfQbSHTF3ZwTTfakV6CZj3guisrUsJKs2WMHG1/SX
dE8611yB76Jhkcei6ohOF7ENRfuIov6XDNv6zzVw6bS9WtilwVWYwl+RyMSgJRxP
1KQr3+wBtxoXruxIfCftcU9DW3SwDrfMbrTmjqEDo3qwdvQUa2Be44uXdyYpsxdX
ifCUEEA00ZymsPTiB6kkxA==
`protect END_PROTECTED
