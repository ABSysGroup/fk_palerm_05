`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8E/kQNWHBSTZR9k0LpNCFs+VAgMor84s+FFc514PQdZiSV7MSHAO6vxkzCiykXm/
HQM1AkoIboBgcDkPqUAozeNlvGlwaGoKWqwvdoXvqCUijE018ueOxVOqaI0w0Ao0
h0WTEC97hTsTePYYxKbRf3OKSNHs97QQUg6CuUvME/its4PIyLMJhf07HKVn9vn4
WI9au4GiK86kz8LRa9kdmzW6UtVf/O4+GqABNjwYOCHkwwi45hegDYGcA0uA4h9Q
`protect END_PROTECTED
