`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WWwK/zs2zYuDIbm8XvBgFfMPbA7FJ1rzr7XEqwDa5NMsBvU+aUzyIIOBWzYXrlAx
KRep2y9bugKKspBSOC3ZSY5IR5bww79rHcJDL8fDB3LHofMQIX2qZIek7276ptNp
I4/hW8OHZ2xOEje9TeeIznlHk5Cokb8hG5v4YG6id2BCLC4MCEBmTY1A6hz+FBFR
RApqzdS03mykY+5NBmL/msZYdP3HSnGpDDJHTZfJEltnK2OPB4agxHImrXvjxuGj
pi+rgHF3bP4VycdlLUGNK3q5XjmZE0yeezqDK+IS+vsycvseV8iHOq1N1tOIoqfO
8xi0AAlKAsFg00fJW79865q5t8BW5X0LBA6rR8tRFtSpyZwKRcgtV29QUpKRKASZ
wFXZTpp/9llfj0SkxR2LJMG6qiBBDIqZrnVjYhVIdukXWF4LuOaTlyS7kFz7XV/a
lepBp60DohjaeWLaIZjn/l5BOBpNg6hFs9N0Md5bkvDIN3cFFDN+4xSJdiH+ZCAP
ebSzP0gbMUQEiw3oEu+4V525/TPzFW1WA4flt0hit9OuEGq5VbKhJUuNvSUU8eq2
Cutc7TPWjzjkormyeIMzWVdB3ER2jgBfJkEBHRxU5nznMEjBzE73tso4r8AMvnhf
acDdy8uuoZVlo19GJjHPAvbN4e2RavClxyivHXB55YfyrnbuSRtRI/g6mzsSmlpl
FInAxaNOGGRxuTivmMk44jWApUK7B1CiPjFbub7BacMh02VWlSb78y+/kBpJZUi+
hCbKBuVNUiLPqSySrdBQww==
`protect END_PROTECTED
