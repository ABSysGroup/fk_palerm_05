`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uITr2YmuCR5f9+o2H6yVtmJTlsRfxrC79AoGJED+xvXVC2ap85GNwS8klym6WY6X
Z58SfQbPqPTtwztgKJJRmXicwJpCzusUTh1IKKkEh/5VxJQqhUjCSeB/4VTVEh/h
fvvEzdu1TT28/MJqi+BhB4JsoScn3pZ8hi8+Xnfb2Gt1g+Y0deUD2l+P2Db/f1MG
TR3APaVyTJFe36kG8kh3voGhc/3qw4ZntkR3wuhoBrdD2WX4+Z6YuPp228iX4emm
RmKC2MYhTdHzMWOmXUHiqf0Hkt6DdlvHjkp3puRL5nqCBzh1m/CPKs+pLxptGuKh
mCtumiNsLV979iW9AItEIuupE1M8mX9yhzmx/yxk9cO8tKpbJNpCbE98IH8+hKH/
jq/zS+jIszocotOVGOQIKLCgzYegznqmcI14GjooXFZn873L3tCDvWMkYE7Xx5sn
`protect END_PROTECTED
