`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g8RSO7Ep7TkbkRaRSeyIJuJms8yDyEaukeeZ13pU5cknVlat2J5Oi+deKvrXOcF3
NANXyAT1RXZ8qZlE2CwO/zF+vJ5JWya1dvh+AbO1EQK0PQNSwFS6lnNUX14fvhYa
DXOBMYTBxqFD/zmYkLbUQI3C5oHf+ZZsfwdJsp8rUXQpJwRgEszmXKbM0gMzxjf2
irnJTEcGpdMng/w2N1mY01/f8DfVAWCq/ymiSCjfMIVpuDx6985pWI1wIYyjEWS5
jWCmVKLjQ9XTQsnupIqo4CfKG731aHi2LdWiO1QLVG1B0gcQdmnNEED05X9kaCDb
ojhaHgHKk6X+qBlXSgdHetpU3tlHuqJoKsZl2xfCZd79bbAbv8xxe9Qjgl8Rvvc4
Lzx+akNtp4AgYAivk3gW03+2UGSuTsbzzhn/XEkeIIYoia2NKdQv00MNvfBaCCy8
rpgowfDfxTk0rjLdHORsvw==
`protect END_PROTECTED
