`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nw9C7yzvZUDUHTz6k9CqHhkV1pCAj0dmu0AjJHhFo00UAtwzvdXqZKJonc/X+lcX
0uX8rIWueWp9BuWiXZe8adkn49TsOkr8OZJ09hx138/+W502p2nnl8KR+7ATvtMq
P81r7pGhD/9YpNoHKlDj+cFC47P3enIhJ0vpAkWecmISOZtW6hUYQhGFTxfWqV79
ceuTdLhlzUuzTnn1yj54sdQ59p8m9MuUcbEfD7P4G4J2sYfKdFOYbHnwDSKtokov
b0GetBuMwc01DbwS8gldBGTGPorXMdX5DmEy+Mga6s9pOZSabhG9ZQWdX+NhTNqy
ho8uFLc/Z9w24k5nokeRvLqvpcNdXHvfWV7zuvN7lGvrzLxJON+dau927q+1NGrm
yC0Y72tC0YtcfNNr1Xp0hf0+buVLy3KXDuSM9Mdn/9BP0INRbR0qmos3IenR8ozI
qjxbS8uuMbJ6jKYL/HS32szvzz2Roy61z+pHe9frAFDsaWJUKIAWsQI0rt2nhhFd
`protect END_PROTECTED
