`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZxZruvzRbjDQnN/iaFEdyVwAz/+a+yAaQkkWeatyclA/eUN9zOoBk8CN/2MQgBZw
wYDaAqpp5X53SnoxbZbs722rHZfsHpRDt4YnxGOQ90URZMJF0SP5xpjkuOUF/OsK
bPAketYxWueSCiyg3qVaEKB8XLrRYL7OsF8revDcAvJknN7VXThq6xMXQLIWfcjf
Whse6bZNlKZJhI8hcv+j68yBSoH4Gn0vn9fwFjsKqq+dkP6svg1oLrosnHlSChKo
4M37PMrhYDCIfwx+jgZIgA==
`protect END_PROTECTED
