`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5z8ibMY61erfFzJBEPxbJ1+dDbPH5d1aLio73qOEJpDA+RVvrY1wZurldnG75qci
TKVU0HmxVtNEKRJE1pqNMlhxEkfyBKvC5G5ILgqMjllc4FOes93ndH0bAN89JO5S
XAlPFoyf+piQUdAjnTTRBzLdcV0AIqpe7dBAxMJDEKxWvapJs7hmrFurQIRvG9Ml
1eJHVQp3gnf2h6OY4vAh0EeTFhuxH9sm17ADV4ZpSCFsMlfoi7UYSKduYjcpSJJl
OPqJ/2YoDsszijnItfGd4qk8osecNzjbsSTSYM132jQ8Zk2WkZAxvW87KslnexcJ
F1m92hqXZpYtQYAcPnXO1Lz3AyTG7X79KcucxX27ZSffs2JMrDixuzE0YfnygLPx
0fT8wnMZ4UUB7gX5i+wVRTvMZJAKB1r+zRvIE3AQcenQjX9olSjOic887/dnSrfG
gVPaRATgXGv91ZATjNtv+GUE7Ip5xP8S/ZU+6CBLCLeQeyR6TUe56IgvZX2Z2+NI
FU6PzO2c1B019d8/bAkMuqzan0Ue+2n4SbSEXWw670Hc8GfDhVZZlPYwiyLF/HVk
o2AwKZAgaTt7TpSsiSEQfVtlk3iIa6tamw9cjTufa/2qULZn6pqUNIPSPhiQDTLc
zRMr6pzWLSpffSAXzH++99MuJW42LMi3gS/BRX9pCBk=
`protect END_PROTECTED
