`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GOOZG6MERzb9LOSZWHjBhk1Re3pLhocc0BKeg27ZbAQpjJ3m959lio3ZUXeyIAYV
6LZmToTF1AP9OEOaYHmI/Dmk4Row+2CJ3IutZUVp+YED+nG4vRY/RPzTnl6m2HvD
oC+L6pNBEEsZRzyd9yDsNCw+J+aqent+49PIDsaP8IS77Fy+aYFXsbAF+vDKK2cO
MMmXcmXy3IMHLIAAAKm/2a/W4sTf0FcogVEIZzPE7tTWL/TCq1esIZ+/UbfzgYnQ
+2dPORsEMMi/LN52fQLRQgVexFRyrxDy7Bl9XRSImqVPWb8Ke6Bv97xKlVdSy0ej
HMTPlcZ6PpV7E6ep42SnyLEo5Eld8Kg505y5WDNdtPp+LUa2pA+6kRPrRjG7Q83o
SfAL8TmdaKokjf/UK8kpRAX/tQkU1VSXvuJKqXiG7lUvqrU6aA7gj9hbakAr/H2V
ozpdbnGnNm4XCU7LZBaozw==
`protect END_PROTECTED
