`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FvOzELAGgCEN8NntOcxKQq0ml9UOIagNWZOU3qd7ABdznwONZR4GZJ4m9VGcEUW9
HzhS+UtKNlsRByev3tnjqJx2jAApjEqMAtygQDaXXwFENdjNqoPwyeRu2ROQx3vM
B3UFWMr/i7af9Jotg8bD2S5puKyR/WQ2TWDG3U6x5c+fBzf/rqLV7jghFoMKtBm2
l5ExwfeRkDuNuBNmoDxkuqV5oEHfAaLsfXpIz4UG4f91hJlIPO2WDBmlJMRCCkak
Q05CWtfagaVnFMmJ3K6dKTuSQGnT3DJ/fDILSf131U50T3Kk4wcwTuAw+rwsS6GF
7VPYXHCQrp4POq6gF+LFBbBcb97CVT0xZVgdbYV1AkHN1wisGsrf3hprZ2Mw8b7p
apfbEYcuU7bIk3blaDXztzSYq1bJtKa8srb+fn1oSJouyLZLQyA7N7dVabLlgk4S
aKTYZ/IorKeW2ACoNZG4vmRfPZb9+z8MlGItQFmWtLWkz0RD9sp/Tmblew1InlMw
V7uZRVFPvU14OAtiZ8HbIR3BErA8pQJmBaZNzWx5xduZIVbBhE98HcMU2KWUvZFX
9H9AdLJlOqNfE5wPFySD4IfWgnnp505MPk+SqKuO2Es02Y2BIt/p5GGkWUAbNehp
MS4EOi4nQqW+Hs+/0UJuwSpLwRdgiNwYAEiJiQKCOb4DhpiBHguoOpjjh8/punzv
XS08fjCHkrzDudZd3S91hspi9q8UaZBgQ76+3smnNxiMVC6bHbdjWz/X5YVOtZNV
x4Hy1QFmK5nE2cxaEemZIYExYKy4yw5ojNraaQ7KWmHckCpypnz+jmybOh4jLHbv
grycrlPxboG1KHCiVRqp3shTvTASuKvOCpiJI/s87VQKT5UtmrkPukN2fTZll/3L
DMivu5eiukBOIpKe9PddB8wsVlQL2md19O74ibVjrlbTd3m2w+kcrMF8SDKOBDta
`protect END_PROTECTED
