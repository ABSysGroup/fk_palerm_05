`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E2JJeOcNH4t8EOFWt8pjQMk+IBQZgmawfndziRPSL/9EyDawkZmJlSzwY8PH9r5W
Ga4gp6sZU9tZrvgzpRFmeQqdKczCi5KAydGfi/mNGKa6snl8JkX6n3Ofz3qwQDRR
mqIluq3NmzMojNhKYtZmSijknHNLS76UN3SbB0oDb3WX7jemGom2pT9UAI6FWpIP
2Z7pamcfZZ4hxflSeYWYSu73Z+UAcNwBfb4I3eFvFUBpQVEOo+nJ+9HjPCUzaL3l
Su1DAi+2UHVQaK6LXPUOD7QjPsWo2/Wu96u+VueM1uV98+fRGncrXyK6b+kze539
aMArIi7flk60kBE1euKjK3MhWxiO4joG0DTpxJ7NolVqOyz2WypW7l8vI5hZZh8r
7Y1nFU0lFi0QcE8y+sy1uX2+qnSbOl2ey6TeJHlEHUYthWiFHYQwvl6SkMjj/ZTS
2hqemK7xBFub1JTFshVBJMq+3H4hG/7gJv37HUIz/xl1VCrg/GYU5ScZK7xt21Ar
IGtqV60C+XlYVJ7NZNd0cOHIbEZA+VeZK6CkZ7zJooPf6MQRZ57DoY0m/NpT+0GP
z0/h9CLzri6DduMWByshBkP92w/yiOyP8Hz77yyADdSVL5p6Y3Mjy3biSuDZHWlU
vW2NUSi4Vhu+CMeZxEJXUPbAi229XgBK7kOlU4CjRFIjOwxvGxoubUhkvatq0TWJ
2nIv5cgHB5Ii3E5dO6GE6yrgY5gF4lEzJjwiRV5mOhEd9zB+8A0Xm7BKk+zPIpSO
0WsvE6yhD/ovfZL3FsJ+p39BH39/Cs485D32o9Hv8k13bKsHD+gOC9ghDq32c/k6
FX1daDVT57fGW7dH1RWxPFE36FbaMey3pKzhbWXD3DiNvNBrVWntLcOjAutezxzk
7P0VA9ojCH0xXRv3bvYAhLREKbhIolQc7GeWWCEFtMWc/OHf/lhrMuRw19FV/wXb
bzL4ClgI2RBtcPbkVlwaB2XWNEcHlYyfubEiGNgtJIpRZpd+yNon1+mYJf5hxTL4
fAy5naygSFPWJRdhORiUftzNVZB7rVCRFcO9yHUfhFVu/tZ9isp0qEIaEYBObMWH
Ni2TXpKbrTOtTYUhEBMpqC3RcK/TRF4GOGUZxPBrdGokC3oLve3W6iPz9diRBw+x
dzMaYGzvROzncdOxH5oT+lnOqXXDkGsugeNt4Ly/Tel8Rv0fw+lUBv1kdRzVh/sa
/XGNwgyVo6pjRETLOSGa6lKarQIob0edxLKBdq8d0xdDaKW36tX4DxRM7xcvHwcc
YB1QKAZPWvwL80PoXndbv8ZmVUWgK4wzBOVjSCKGW42RSoRa6lUBs+jXjk8RiiDq
y4VfTthIkfKYK7BnnlCuErqhee7fzOAx6kyyZcuRJbw7QS1h0RYNmSW1muxTJoFV
aCQBDULFF7Im00t1PGXwwOHNoBRXQmIKxuEmAiAvrYLRvNS3xMj04kihxNHsOGUA
SZpMr1DVtt3JCY4Rf5IduT9eD0EinT6bZkl/UWw2I2IXT71QN2QB+KBw9Nr58CQI
UVK9907+MXToOCzX0vFuM7QTmET7HwU5A/qUbPHvBfHrbfUYYUwC3Wk+Das9Ao5B
dk16hvri9R0gQ/CRCTidlF8AR9k1+5luRU1OqgUqig7pFu1uaIV8nQUe5XzLPdfE
QEglfgE/LypxzwjUzGWNj14jEDo1NXAcu5sSb3CGt1eO8q8WaI0U67kZeJnXiRYi
1suo8nvG9VJHP7i5m1GQLXogKnvfqCAAUf3wqAzrpK58akr861dMGyIBU92vCfwu
LgNN1RGJwZcziu00NfxqjapHVPukCUUtChHhcRwvTuQyf+d5K1k/au9dG2eD65AA
IVfkNQZz5BTWbzX223lVBiBioneVYwTTXNcIrODlXmIoQNZvdOCeMRDEDiaO4TdN
+0ZN3ZF7ynLT36dY2KemxtZpu97b1cCk9+4xUnqB5RUU0fCyTmZW+WWsZwEQhF1x
FvIsIGdTBcs3hOPeV8q7DAB4eUJU2B9ILuRguxFuz+6Hhd9RZjorXUbOuXte9vJr
4Gc2S0wRy5WU+D6N/FU3bp6uUqcSLu2hOLMQm7Ri365Q9mwulUDoP4OKXMTrfz9E
WnB/qwrv5L/FTLBq3csTdjr2XqfU9Ppra4oO3N3VbPipXELkL5Px+23qFV0p9v91
5sNaVv9EX6Vs2dd99+cc8N3lT+HLTxHLBL21kT8sf3gh/kvEGSFCybMy3mDg4mrP
SN0uYw03tOebKEsDanNru33sYaCzoXcTCImseWRDjCQExxPNmhgutp0taN5xp1VP
pClxaa1CeHZ6gk1G6ksjNDV+8TE7nLgvU/XY2dut95b+1ebyLTHJKiU4JUBZ9nFO
yg/lVX0o1DdfjeXyynP2n2/EEWFNw5hP1ahQe0TmXjiBJu8b+JMA+dNwiyDZ3Yoh
eYIxfp64zvuZXCJfD9AweAHXdmq87LCMfher6/dM3pn7cfUZa3jc407FE2O34IqB
kwlhmdKI8tnjiTL/rQroHeeRVbqHXeymxXnhjHf+lgjI+1Rs3su90dfcR00IIeRZ
VJWRjxAUhQkabSFptkvXXxfM9mSWmgdXwTyCHU2MB4OdAYkdeTgrzcUTxryG6w87
XplZjYSVSkDfqxRm86nwbGIjpXf9BrWglznzkwjPwpczO+zZRhlQZZesOez6nuWc
p6TaN+dJ6FrhQOkKpuppJujt0kk9YOhgyvg00UDrh/iRmZFsjERsM9LS7uHvq4jM
Bu08bsTjie7MyLcT2JnLQ1Fhf7lYAGxlCYQBvpMipRsRTU+TTD3s0NryYE6S+bem
ly4XylTqkCeiHOIW9o+OAfA0/oxAqcEUPNKTG8hgDWyiC7JfbCUwgnBhAK++vik9
0PW+nIcNUGJMudbq0z7Ep4PrU7E11v0FCSmgdSnMe7nhig4Gk/1wP/fxuBwTVg6I
xr6diBt7SfhUHdcXIWQkNuBic3/hgQebEl38Xu/cbXOVNAzTcle1qtiRcebk91d1
QId0yeH1xoyqLS6Q/+hebzxZJlALtpEQ4fgM9Rh8YcCMyoR70QxPyeeUuCv+VQUa
WyjxJCg0bqawcA8TU0qweDbcAtd7j/T2QT4vk+KqaxO8u2E2OtXNQrDfEDBt2ZIY
d0zo4zb6tJz5kUZ+qKtdXo7+7dvjrg9cvTAkc0wHlpZ3+VfPZ0RSUSeiZSx1OCdZ
1FSCFDR4N+f0mc7HepPIJf5rVOnLEphWr4FJuV8GkGpDixlBQebkjfEZjkYBx8TO
Ke9Z4Coze9ErfcWk0l3sGUJ5Dw7cvjA7KR0Lzo+ubcZv4LFFJKeaSl6YWNAKVT4j
BvSRIdkDMvGcNfC09GPYBMLdxGcgBPPOcnelPZYtWC1SiQGMKYDKAjVmbrg4z1by
v7Gi05nkLiuNekLwpcE8r4AAz2pEnm2/+2EVPEHZ6fS9um4fErI0YhiCO0hvDFzU
PdUWpDEpGqPfQiJViBkgLumYczQoeSjE04UYQX3d2zClmHIMT0YBzKayH441gg4e
COkQIix6x4q+Je0iIlm1jiiXnCh5ETnmAlphqinojKJ9YX2emP4wXN0pAZmzKLgu
pevDo60gNgfhLwqIwcHwPe6+IB/0AjZTWGaYVdejygczKyBIqN3dTjaE/P1qbxoz
wKsScl92lAFz2pOXx2Llzw2M8H5VHGP3DPA+oC0D0ZLtNA9kb63Pea5f4ckteTMg
bXtl10l8Ya/nj8e9lgqXQHXToqSo1/AXyoGao9QRztScUrYaoW2gPjWs5+/0E/Wu
JaUYL9HJ3nXibKmMLK2+Ng4LOfsyfRXPoSIZZ00JWzPZodPMkfm4B/5xLByIOkbV
9/lxxkBRbtHE/KpeMn7aaWXZJB8Q+BLhWfWJDKggcmTc+XGmR1lBTaGwcglE/5XN
XCP0cZ0l6+kGLMi1Ozi1AsEoT9HdYFCJGHe9SnoqqKRLV1FoKLNa1uvaenD0g/aK
bTGPjXD91rxnUHQAeObEznnpNiD7PwAaIjf70hoB5pwgWquNF5LvrLTYpJ03G0nR
eOpg7atS/x2s+uCitxw9KIJcgveMfX/2/Qqi9bzKLwSRzPPQeCb7sh9H4lQ4D0AM
oRM1TNB1vnryvE7DSp8qbR/OBhldgr/BP29ywLU02Bq93PN3JmZXSo2KQ90Ppsjo
2I5nR4Lv7fv9I3W2tGyNJpTS/xaaHZdo1+zn1x9FgowU5DL+7FU2Mw9y9OeA9HTh
zNOxiMcMmOjCCJnyhfBNZHtzr1LZ4WxMX7Je6hCSFmXDLholNCjFd4KJiY/yZ1u1
Ik+tTFwhNnyJMtexpX/dNaY1gL/6+KSW+hfXpclh2X2Qac4U0fppQHktu5+61zRt
Y/LoNliW6LR+K2Hb5nNHwy6w3it+bWveEgTvkev89n1SJ40F5MbQfXLwcagv8uZI
NuxBgFQSaLo5Tdwdz0vUw2PI2y6gkMojBGVMNmtUboxOBMTlSYZGe+kSsPG9ZJFg
kA6hU4iaXrZV3M1rtm5xRHVSPRzTAGF56Mq7xpsl7qibEjpLjGpCE7dFKcmiJGak
+O6BlZ3wEsaPwZ7sGc/zbU/umqdWdt3++oRfLclXBJ6Csx04HodZJPZ6Hf5KyVSz
I46uNyVM8Il+8bH/wLi3gtDpdtRj2BZuWSNm1iatrqXaL555BZY4SMpzA3XdRX6Z
LF2o++Kv/VMMecCXf46L8qvu0qndWSFk/25+YRJUVt83HUcaCDeSDgjriJZs/sY7
UVGeyLog9l5Ui4FGFnSCc5RyyWzg1clnVdInu7Sctrrd6qRpisrN/NfnN2rci0Vs
iJEC3ShJWVld/QDJFh8zCLWxDS8eHbfTsFUSxW8GNvCLQ2VNve5cx0fe9ZeswzK2
nhLod89vVKOXETrtJPsEIaeISdX1Ic4hOCeIbcTlYnr/ZX+uKvIe5y8tYKJJY2KV
7xdOpvmW7bgyg43hs64+J94CjCOe0kpWSsiS/c2/VwQ3J65LX67CQJZcU0L2V2HW
g2c5J9UghFmjb9WzLiQOAfBqwYBbKTIgu/ewd7WVnc+y/WBGJJBA/Q1gNlyD7Toq
0WxeHL98Rcbc5zrUrOsiRK0C/i+HDQyA1sDZpMFEwtg4m1CoBi5/nSLfqT3xAHWl
vfr4cz/Vxn5IA+ROL5EV6HSrV2FuoXlLPWqH0PDXG5cACofHrr+x4vipB/hgR8ka
N7wJXnLHByQWhFsOvu9/2sqgN1PZaGKLOszNSeu4znVHEhWgdzmCKgbocDap1dCY
JTjPkB+C+aHWbDdRcXUtb20Io5HlYqKI6uX2DcLywzKVfBRU1N4w4xNHJMmZsGOf
Sj+qyv1ookevfCjiY7TL21r/qIAQmbgfs17o2tHugnuP4x19k5YgoYW097yFKDAh
og6X6Bsu+Y3oxtOQeW7UjtnRbb2WUr1Sjqamn64UMEqXd7oxfFhZ2mohTgyzAZIo
RinE5s+OFEJ3YOAZsba0uuMQWOY2FZX4RqpQ6bbhKIwcROglGAj4wZoVqn8/Veyf
91+9aDxGbOWxmmokn9jWZoJRi38mSKaK1lylISJ0dtnr1irqqIfTXHRtA18tBaOd
nhMHkjZORDNV+YB2WfB84IzWK/oY2N584uy36rCTQw0m3SI0BEajNFhbUAKDY/9P
4sPSY+dotWSVfmKImoDd7+uJqhFFB6k0UUhMYRZx/3uQEIMBrkv3joMTeOTru1DK
f5EHEW5QPl5ANzpX7apEiG4s2OUGH+kKbaC4gQpwLtFgZfdQDU6nINQbS1S+ORTE
ZiPF8kquFkEaANV2ryGGyTRfCJ1zI/kS3rJECwaH98RTgCNHuFNFjXIouDNB5qdv
/NeoZQu+l1/xDAKnl/inQpviu0MXW4bjBHtqGceUUTouke1F6NwA99hBzjniNtQ0
zSJKxVNMKakkmw2niooo2ZNLixuczxntNCA27nixMw6rwcBSVSJ4+PN6dYQFxFIf
dESsxrYug3AwBlVqz7MaCgxOzzaQzqZjGOPgwat1nJcVC1QgMS8zTlZJhOqLnUx8
HrE7sfPMcvoRqwOH2Dbwwti6BrV/JDBQnwKWOgTtjhmhUDYVzm2qV1yC3fWlHkyA
cADNzWxgErixHajQOjw/D041nqf7KGMm/5rHDst3s/x1nO8SZh3c0vjLI/K82Ubi
HykAJ6f+Wbi2CNhHPZxYtCdX5Q1CWpw86Yk7hE3LdOyjIkJU/Gv5Fwm0LxaTn9nT
bqY8dvKUl1oeRswgB2UYGSMXAg9UdSbIrVKZHWRU5Vi/PJNUxq1N1lzbP0uIOdsI
E2Acxntnt0vNcomZWYnOYCyf17OtBN4gGUBHfUGFfWf3kVIO+na2eNYc7MzRXdIw
rmwmu96gdSwNuh27xclbpWxqwUkT78nu9Z5NIvq1xxz5ZILmQst89grV60gHkWYN
98dWw46aCfWJLWZy4b2///fl7D1VE0AYwvSAITF53vrZYmBicua2raoKSORLx6pQ
osPC+AjH+27DvTk9REYhFEjX0F7KDPvmsbECypeRJ1lVf+eE8xHfFo0wIWlYpC1t
tTUh4PN+rVOZfBYRYT6hyYBqOH5zKkFB5CHaNfKbOxcSBxIRjvegWaz9paJWcM9W
3Qf4nAiCWcm7gVuV6qFSlKbcnPSOvB6qR1+2m4ofEc5yQHO7bQy+g2wxzZQlY//+
LgFnopQIuBz8aZCY87+5qSku7ZBMCHEopd34dFESzxDMqAYOcX1UJw/gCjvKDlgL
9T8H49239fFPOArNJj3bPriE2LyyQEslddQXrRNtqfylRsz4CekpefHwdhVXfrbr
Dn3YP7ps6uAxOtBztmGkUzOx+r/rJ6tseRNl+JeAGMreAa8SiIyvV+ckuAFBVQru
aPn0QuORj4jRRKXTNcbrzGh1z7ZlNkAwfaZk63lTKv+0m1f5WxJ/01poqjBNb2p2
AcGgkKwTXDzb2dBa98TlG0jDiwhxPfQdZxPvqSf64KYY6wu15TVvQeVs6wJig32d
FYFME/fsuU+Bele5SWU9fsPA5Cnjru3X9Kbwtosx+G1cr+kFLLD8nF8PuTz06I67
BJ06GzBQLrAzpSps9UkCUNN60HYPZrIT0e4khBLktG9ESQdoCW0MYoIKyHdI5OvU
pBzjNTtepKAdi6Nedv0L5kmBWScHoZtnCbd4jdvDxgwvxXuzAbcthxJzlINY7UTA
B+iIUvWor6YBp4EqxdxJXJegU76D48xM0Ev/kO12usCXpqyt99nQviqqMNqUygjZ
TTgzNAVwRmXuptOYDWE6+ooPhXET5JOnE0ELRNTrhb7kRsBpH0jRA8B0L4yvM0xN
sd++LQ0rRq4ZeYSkvBJVaSwv+hbI2wRVZ34LkZ/CpiZklLUK7V2Xy9yF/SEwK5r5
VkgU9TnvfnP6lSIyCD+re19ssOC8OHpGfpKuYhyMA/Fv1kzi1rUNsDr4t/lN3Omv
igLGOGpKs171iBsqIgovMhubXNlzhxg8UkP17E2xRYYPlKLBm0cAHsZJQiyqw5w5
Kam6nefAjSM2EZ8Pl1jrbK9qOREuv91P0IsFWXbgJwQin5ed9Ifm6feqNhE7evx4
SmGa6d/egKBMssw/vLQjraN1cfw1NqCRwb0uLnIlUUy6vY1BLjFU9yHSKeLoIrFA
JuR1cv1pCngpNLO2kkCvHQADCNLDhyB7zP/nJwQGNlFOj1spEl/ZjhH3VP2UYbk8
UxveXnSYo6Z4uwo6xzHiSpfDacBOIVPT4dexeYENYoPIswKYf9bX8d1IrvkoiL4u
s8/YuN595zn6U8uFfGdlDP+4uaXi06CPkWyDn0epI1U/7yyQyVwJLiv2U2H5tosy
XyU8ch78BUb4XeVnDHCinpE80K1He1MTeJsj8eGhHSmMuW/KwRufYHBH9RuXStPO
3MWoAWZm7DAA+H/6za+PKp6LfKEkE4G3nTnwO3eKtN8piVpseKswXCL/C5QkdbXa
SO76Sfgt7CYCALtl1jS3SlH8oYSzmbdaAasTvHlsCcykIl8IdwvDwMA1uBdUYPs+
xQvmw7BEuz5ydQbMmXVo8YqH9lDJ1WXiMxrtz7H8n2q7IWzTPyfVjBjd5tGB2YG/
vfTGiR8hexr5lDZR1D0yWR9Yz/YxUZCqM3g67Y1v96L0i8tElcQSsLUEqyKLy2QF
cIyvNywFAQJZ50Y8Pt2RGSxflGvWD1ikIVH4Bsb8eEzh4OVdimK4EfYJNdeoYTT8
DArwM7lzsiA9Hg6OnUDyDyePbgDvPZxLFsNwfF3sGFpbI+zejGkB0eyeA8kjJrSp
6unbTt2XeyPpJ0OIYwMLPd/pSqKC9mOCKRK8KVXHJ/f/YzfTxrBbJ7s136A4OtTn
0XubriqVKQ0Q5kIWL3FX/sU5jQWT16t9Z9k6WptjSndMqkvggW+7dHetXkxXwaOU
92OUqIbQgHOKTPRKaAwomuJPiLpoq6KmpftjGIGJOlJFGdXKOPabaEzocJ+bh6XN
cjHCxSvaXr614aeex0FOSzqH1lEiP6LRwVTce4/7IgUrYaTz9z1eQXJc5tMiPNEm
xFWuts2MALcNNasC/pyhdeD1vS67Th6DyxRDoZVjEODULCTd7iQ2n1R7+DvrhPQG
xCd9+pwyeH0GCeAWc75MricsOk8L1eBEYDmvY+acHjodvznjKq/UeGqQ/NTdhyiP
Kd/ODZwJSajX9gbdr3XIx0V9KtFGfhACAGaa+7JkJays8SiNrgN757TmffnYmpTR
lLVgrLhvkpcuCijjPocoretPNxhBe6+qbDcn2srRaYe8RHt1RPWcY1MoNfjM2keR
GWOfop0YqjETdhHRQc+2hlAOYF56hUK2EAnBQUu4cD9+aMxvc26PF2Yt9feNqGnQ
oIR1uJrjOR2jjrJLRZ2GY8yHPpenFmsFhfXlKnghzLoVOyzvXlURZTk7UXHKnQ+P
u/IZpi84t573G2viXDfjsKJBH+Y0kADN9eORM8c/okJm2x2NRMK948+QmNc2FkMm
YVbrw/b3nG998s5SSuhp7RwxV8IOMFm2teneT69EhOK2iNaQotE7mICEkdChrZob
zUjxkobMPHlHfcwTmiKSmAK9iS5hF0KpGHOg4qbyaMKsX/zZjJOUkglzKijuNIkv
NxYXbmW4ENKyDdc/bzvPV5MkhHD27jj3wi/0WwE+w71J/u2EmKZIsox51eZf6AKJ
sGqDaTfPh6OnjRX8+lH0bF2bxbMWzbYTFMGQsqfEcwZ9eJj+Abj93v1ha0xHe75i
plLf+95ThxDu970npI13ElkhUgQ5Sa9vrowooZkqXRdKI0skqapoqoKa71LR/XPc
WyVBmOMO4kz0ri/wdl1rCed/LQcHsk7wabEnWujvsfMKj5YyRDwpHAu8h63thn+u
VKf8ljk1u1gJWnob2zLH+X0qsolkx11fO8UqaJ+iaZPBXW9VdZoNE4F3eaL+fYOl
cmvXZYB2BhZb+cQF62aEU2aMIDs4g+iKEebS8+ocUKNx8dS/Qm70bb+ivKkuOL2+
B8qT3LXhe5TelPeRGAkBcvfKwqyVv4j8yfzDPCBxzJzq0TlFXB3mV6FL+C42Yn24
X0QmpIX3374P0wAaRoduwczCS0yalBv1bro78nVmWv31ZFD7GV4JLGmnfySiF/xF
cGJJOep39YlQiQpMH1r6I7TFHwGVSodUtGI54gtASPMCOHxfdYvPr48vJWgj5FRe
v4D6kbSPyiNEq4pIZENt3Kdp/bXchMqa5z9MI3BJYynkzcpoYYZpRQpITniyfrbG
AOaq5xsTxH3J8LRbAATohgohtP/If/4o+WQfrFz57i7OkDB/HEyeQ9dsyHt3uom0
xVwVS2evHXb8HPwenQWYp3PfoldC0jAYOFlgbRjWXKnpqTRqXDZOJJWy9F1bQkyV
xmvYlRfUGCFWXRu4Hq011fNaK2H91NjQGsrgwQi5Yhe31wY4dZ0PykWu5s+ey3ws
UlN3OIPKgo9mWVGs3ks2JBbK8dEy1NxHwKx3LJTZb9ohJhrR+f2Cpa3nx21UsMqv
EK91E3MGmdD9evms2y7oinIEELzTx+sK6g6NodWpOhVAIGzxHG0SiV5WUxlKSlXd
8E4bTb5XVLxWTm9hhI2yzsirYiDP2k1ugZrB4kwk1ByLDystmAplC3Ml9q2aVCUD
3nczRKk8r+EKuNArEouHf18kjvRiHNU8nURAbNIuue2dKw5CLMOYxIY8ds7WvjvL
CC41XLJmFkkyivt0jVC/ZBZHwbtHNtAyccaPAjSmdQYbPDGRx1BfYFRuuu1M24GG
4/0xzNCFMdG++c04wDNQRmthqwIxjQOZrp/OPaDxBjwe1X90zdRCuqnHs4EoeUQ/
kNSbVhp91bug67Jew19ZMhX4Ta0mswEwgzkuIerwKTYZvkFfNR1FJorpZi9poUZJ
skG+ygAd6GSE9E+VUPwh6fBTyyjUSpE9y+5p+q7IzBA2BSiM/Xoi4dECuyZ5B4xe
nYHaTSQUy5Y6izWUFPuXlCtE983UGNj7FrxJ4ddAfeLPPyvO/QwAnQzziis7UmqV
dMkp4YBpQL9l8SvCYcDCp9G02gKnTMld5TvKcJYGRwTqpuO82vW03EZMNXeE0pbs
H0Zp+k6qyIkp+2rlLvyKPj7uYK+Cj7FDM6twWVNFnMbNF7k/emmSiF3R4T6cevC4
Ap3cZYtMQbldRJ8Ug/bD/6HLk/Q417fMjPC6oDwC1kTxc+pD9Wp1aFLOueCUXaab
UBqtstpDrSmdwnv/d7FIS8p/gEvv8SRCjsKlFP6WXfW8eZi+IeyTg34Q/a3P57yZ
/HPtiJftOiKrWp7bcsHIdrpl1RfPPqvAPCL4sgpHy+yuTdhzaFEqQB8RQWUt7Agi
6SPxxXj+3fkxYE6Baw6Czg9aSSYItDnX3rfUjD4Q6ELEfV3YqeTCi2SaTKp3/fa1
OLQv8DAZuEy5EEMYtWr/2+DBnm9QiIvSdVyGEPGXKAJBoXgQBirUkjqEELm8Rruf
6rbDqCd/AO5bz2UxqlnOllyvXEgSoAbJAAJFH1g4fZ7qQIAVIuPRz5R+JGQIdkxV
vXMZyX1j9YD9u7TgocvYusEiLUudYivfKTH37d0EQ+NTiaSpmDdMZ431KQF/7ir9
/jsli/lTKYQ1D743rhLfsmPFAv6zw5pibpApZtOR/4fKB+RJspeuFGqS4zvQfbul
xX7wQATuMyX2Xqnlx0Fq8Q3snEqMArIXqqo3D4Kl97m3qO7gpGgJzEUY2uUN3WkZ
W/BJA0FfD1ExRr5ZragO43OK3tLYrDglzJYH+t5T6GVtNkABMWccjE9FprcaJq8i
xZ2q6/h4cCO26oocH71mURwbY76ZaZmDr0ROcRKHR6mgCoS3JI2jiBm5b5Spv0Wy
KF0HgJdp2nxAjePDhOzzlRMARnNXmIR/QDOP+R9WybUHPND44sZ2CulpqH+AZv1C
Fcin0I51F4kcveuosYxqGmXt+YFtggp8g4rkrauRLnyKcddUltOfSuMIPX93TTfH
x1vwN6UWhzRV7MYNv3Ga8n/a1ft2supihQvmVapetNaHcEh7o9Pcp9daokwKlj2U
Tb1OYOXaHr4BVi42lNWcsH/EoemWl6bFHUbz5lg7tjo1+3qtGwDOZl9ms3O7+O5J
yVhg3A7HSK8t0x0z5LjbDjPMDKwa3CiKPGxa4cGapOGiUUkSJY37ZSo5OeZ1kZ/d
mFv0mpo1nrHw9D4sbLFq2PJdcDFc4SJm6rHM2kh6bFKk0Me1jVrtDrHxnaDyzkbx
xld0lPyEmEcZlaf6e/UAhRtQNJYy+9IIEvJzPWIYYZzo1wjODbYORh03U69lTP+c
Wm6M70cgp3C4hjRFEBbFTiEIXGsAudJHeHk6kLcDsP+5Z33+T1jy2bo6B1FwgoBU
FglIKqMnfz9ukB6rOPImxLdcTxwiHsSZ7yviKpx5Y9X21iOvxQJk4/iPhXdpqxWy
y9fO8qLf/R1mCyBpfymCQr4tGApqg2sWDS0tHiM8JtfL6hVCjg7Pvng/l1hgNQXj
psYkfOhhCaV7q002tXwgYE7SrocGR0/NVd3sNCQ+RB8kyMPcJ0ETzRP7Z4Slri3d
MV749aaTyftpL1d1Z0GG3DAyMxbpM7pZPwisqJ26rwWRx++HoA4sLlcg8PDCaLeE
OIP2SNzzsArbPRmElXqTluAMjcoo6YHTxDBymKUnoKUFiE2blXx08gp/Ds3ErkMr
GzmUnuD4E2h8z62Pb+a7J2xteZSz/iPhxmJM0UInT1v1Mi07tYc0G3YOhlA74SYc
0dEcJ15nyUWIx75+BRLpmnAuXryTPxcx9x+ixK6Fdj71vk3VLNuSfwI3ZYGVxdoc
llo6KFegczuBItXHMRvkAvQ+5PB08jioo9Bovj5miaa4uBIkxTH6zlp5wcg30tv7
x0i6BB41HAeGUpO8t765DKQfSrZ8L4QigBCsTyjF/AwdSdiJeDUs5frn805S+9Ui
0vMdF2b5NovUNJOsCSen2a0pRguOlW2XE+liVo09r8jhiyJs6hnQJO5gqSu5CuyU
bGflDfO7KwecoFo3ojg+D8TEoB1nxOnmQP+eQLJOKdmljhjO5c27A3HSghyDVjTM
fiVivCLwuXzxd4no0wx6bzvNQOMiWmn5BmXePOMv5sZz4NIuG0O+P4dbu5DGGZC4
rEsroRWx2eaPnhW1uaNowHiGHP+j2NQmFA2SRdpj4l4W4AoriV3vl0DWISJo90Kn
WjtIrYZ8x6xAONWZl+5vMmwzztsKm0qLcAFzh1/ybYmL1qlH36HZ9S9TJX7lj+0+
lAz8w5F/DaGMQmaU4NUhKBis7HwdAoAEHnL055Y5nxrAGDKk8sS8486ksqd0ZQXH
GE/m8AE2I+nsjoP4fHOviV5CbZUeloRvxEahstIC/4ZdHLtmex37rMX/pPPtxt80
GopsT66CxlKf9kYit0gyPsY3gaweGmwokcFjGWwExpLURpkaAR6LfB7N+niZw+WS
lVjOZ2MOT2cFrIMaA1YWTYzBJZoNseUzMyLYIpEhfEVXvNvPvpqIyR7E1t30J4Ra
SYXMVg+OnMZ1770rojouyfWyJAw2XnUPvAdJs51s0sdOmu59hSmeldzVFdwFmmI3
dL4Eyneu4sQ/6xkN6ixPPiZkkvaBrTTvM02hZ7n5FpyKugyoJV/oihID/yQs5sUU
Y3XrvLDndxJ3vhMfWDtbkYtJTaxB4XJrJ9zQyCIoaQxOPMJRhDrNoja8MxfVY8ak
Vx+Bszh4na6w46GMnzNbiC2L1hRZ4pz8Hb1iDcmO/bf1z4EG+0Ai4z52msEnXHvh
Dcclf5L6p3cUJLzcwFMqhwdtrgqWGF0wfN1ILO17z9Q4XJrRvdThP5xR04/Y2PCs
LyUTyXs7MWyJG3h0dxZd9e0sjkao6DXtVU1o4pJb8H1soUXrq0y2+gQWdBCqRuHK
Sk3lDQwMmEuPLefZ0Fvl6lpAmBAdH68GfWI0lYLdEg4tvnDD4qXx+4o5+f+xFckk
8txEAjvniBJ8KhrJdREZ8fMJyMTOv5YEEejjAW1c/gUuGmO68vZlHpDpSnKZI8sR
BK5TWEr99gE3/UiP5uXYpT5bNRfnm8qE1osr8mQapIGEijH8u+3zrlmv3S3UEdJQ
AV13TQkbQxEsNjP+0fsvhjuyxFbMQcwL6hYjwmqjsZdBkeaJXJQcfgEMn3UKLRit
P21QtadjlT8jTDzmclh3bndby4HUaf5O//HkrD3jCj3Fz08JXmXlFHQjxsacEmRB
YUCxJIbDOIpCuQFwyOFXOUN37YFkffYtAqT+lTUSrYENCrIcjN7IE1fJRrrmfKa/
yKLk9TPCsyRCJ+bQC4b6VC6gecLB69fXYw86chAUT9FrxFcHJGF41D4/n4FqBWYR
Tgt9qLaNhxEVEZ1dsqsUpjyj51WPpWWpbQ9UUITJ88jkCRbF2+7xLsgtftYL8Dmd
yAQL35FKFc08rnQeI8aiF8UK1KEutHqILSdYXO+8FUdEU6JV4LZIOPqJ39GYgQZC
f5m2YBNaEQFUvqfO+GZtQTEjRSsfXZgievOGHNZCysCC9m9d2gu5ynZaw3giHx1q
l5Aj0vEVlI6JVrKGhiCLI8/GU6rSkx5eDU0ycliidbMgzuzR7W9ynGKIfDvf9bvX
BQxd9hVgdDuOc+3O8fjien5rKTOr7UndwRBOYEniWSVlAMaVEv0wiL2TzQNKm+bp
MWq8+0t7PIYmCKQk9CNHas6yxZPxn98dMj68c6vzIHcmrjKM+12Nu5pNwot7+LS7
Kv5yhFOVA85qjIz5qvBaUP2OS6A1s47X36s8KMILuVppyjY7+tjti6Nz3dqOQimU
zpYwx470hO88ZDbZ+aX16n0AYFBiIursufQa1AfKbHhQnBGNIYclGxC8P8CTafb+
R7jzVzz8sQwsU5wgQnPqs8F6DHLtFsLiddVsaPAdyy2znS1V+aCy7wROmu3yhfeX
6U3GQgsoyXq5SerMmOlXRsTj1o08dZjPB1nyOTOFmOXaca7S4UzwMlPoPgJilsWB
5rzJ0srFCM6N7IpXJLsoM8ETQhIyS8CNyiK1g83NLiM5qFyFyHujPgmsk0GbqX44
M2tZVZjVxB7HNbA8qsgHh9D2RHrftgYBQkkmByzUd/+hK0hugKK1uPxnBuoIn3/9
sGGf6VYjjalf63cYuBt/T4DLGFfqPH50Y9WT/p8LaMkRMPF/UB/fkY+DOwNcx5VV
iR/SJSjzSJVAlpXMRraM24XBL0v+dPRvmtu0rd36wPrdLVXJFjb9HjZC7o2+lNMy
81tqaH1VIAmDzyYDrqGqcsAadXeeWkuA99nuSHz2cHYwLSGCG2gmkmvi5QTWh0iW
wL95kjc9PGsHRoNzlyR4bEkOdLljqmOg+aO8lNNuXlAPwz4CJB5Ow//dfxFtqjEq
wIllmXR1ssJkJyl+797FnDjQcpE3XbrBHMoXhLyTP/SW/5Gd63yKsG9TnjMsSaN1
QVRj1B/LWtimovoj0X37kRULMsVdgE3JPOqLEXiQiiBMbifbjPHtJpkq2Ekx6t9I
frJ/N2aTSe/wsBOLcziUtZ3NrXQIbfiHMlBVUOU9W1d0kWQX/r1Wj2xGaNGayHfp
9BeSRMSr060mV39HBL/hRFPbqrWTbM/79OhkhPzIDkUflBwMMtf7rebW3EjlfNvg
dHggDhObJg8xM+JGwd+yVWjjfPnaVIYFVr2HpeUUZwWRFith2ufX+2taCzQBQpSF
FC5o7tnqccwOF1GbuhlvVSOxB68c3nZU7N522ZSKb+Tm1OYjNUcoOaFHqboR21Gk
f7MyJPae5M0q4Zp/v5UTvvYHAGGIvEoNjzW2GuUxZf9kFUUMZYl8EFo5pRrNgmpA
JQ8IXAPUTJ0QY5TS4eBIm5uIaxdU7CnmbA/tqvFqgzQEVCH6LdltbX3jVlpQdfBj
DSYBOvShVrrp7mJM29uvs49Esw4d+v6y0h2SMgn+qHoQF7xeYRpBG+ByPWeXtJxM
G5pmWvyS/GauleHKbVN90rX47q1MUybzsPh594T4JwSe/4IRlxtB82R8Udzyt1Wi
NvpFMbaS8wiNKAhJGgOYSg1HokxG4MXP6C6NBZJKhwsOMNgb681K9vSDsSQIsg96
jXs9G2QFy4/qMX8a/czAZC0zJ1lemVgetjL3J/rjUxSSNpvvv/mmkStcuVJAyn/v
VMiOijnhnnZATzG2gM5QviM3oT2Ux7lea5e06KsCoaJL4pquV9JuDyerxpYhzsi3
Hj5z4jGfAfytPFu77kJm5LbYqa1YoB/Bny87+kA+5jKW04+qNWoYVdEgiheHWBoG
6QwL0zlV9sHRxkB+ik/jRLw+JGIFaMnYO+xvR2vyyp1PG/589v6YC1WzQIB5kaD6
4R/nmEMy3WPZM6yjjLoP1ZZl0RazI8Nduzzm/Jhtk6JOZJ6BEfR/rNyUekeita1M
3l+uCguAnrGPq4Hn+Hy4rmfPZliDUGueyTFii5MFozOJhnPBdcU9SulG2Sku8D3r
RROKzdxgQnwkWLNqSS/4NkYvUMpes9gmYjgieLWh70q8lL7EvH6fyT9QPVjSbjSj
M6cWdG7CGN2gRvq77ONWjFK7XQkUwex83R5o14KwgexEPmRf9ksjdAl5alP1bJVG
hlUIB2S9rXr14+0z7+8YXgGWwiXai5IBrrNdMTqyuGKXikETOSPp1cH7ydp0/4dX
1TmQuXOvWqHfNWRZh2KzAWesgtVLbwuuJoxedTCh6XDz928Hx75ZqkuQuDvkE6CV
iiXzl74nKHzeo2+lVzjF0fus4DZobVrH3UQn5Yv8E+SwdOLAtscLpX5ATguuRSD8
Rke3Yc8Vx2frFUNyD5wJCxp2Evqm7CpmUo/WypcOjw8hS1m44VEVkzCOjA8N+kwq
jaCl+YJombhx20uvoYlPtV3kGZb2/H6kCnFXibqR23ceBS/7ryS4ER6bMQAEpz0G
vyPvE6SzSBuI3G6VgWQs7F3/v8DDX2j3mZasVQH+wAVC+r5qfchcKRlxYW1NASZw
X0jIjtSqg2Q2mihJ5b0HuWzflIVi9aEKKKz9W34P3Kx94KTqDlSIxRlG+s+f0RIN
8wEyZLUCzaQGF7Y+XbgQgukt2lrZJyH8eTTJxVSb1PNZw56oq/69tvrjGQQGpkVk
/wejg2Y2eyt+VE0RqGkQJq1nLPnjSP1u81C8gcQ6gMQu9jaRV+OGRZmpvSJLdiOD
zxvhkvfK0zXOW+6+kGNf8xu5cSXop/K8Dt6sllxc7HVlQSqa/xePwJQqZOnckxmD
NlupHHnJHsCGoDFFv6XLEGQaU2Ae3+CESnHBbpKK1f4FBanCB23MJxFfUW1ubKHA
jnkBx/8TegUdzgFMnzKs1/94voW5GW8CdrzYz5pnPaUKgmrRQ0R85fXceAFVIwm4
XxDganAy33f3fTEyT49sIBAqBlVooSlLDAdNhoWuT99JzWnlt8Cxrhw6OIAot0os
lWbrj7A/2k+yWcmiEFfr4b8rVQ3Xke42hSv3PA5cwWmRUBIXFIFjgapoL7e7oCqx
MhFHGN9Dzv8nQQ/W1tAVl+/BAYT1nsHvMa/ieYeEk4yg8LhlkXKGUi5eEql4QAds
ozHO0xVutiia+RBK9sqdeW3rJe/NO4u2Oqj42K6H9s9CE4+MmzGt3A+FNmoJpjuF
olZRTUSzGKQ0Waa/SJ3AnKFpuUcGnwDb+or5D+jIxjBo22ODUyY5yFiOWxZE/3eV
UaINgIXI0IvL4P+NLT4J56gQibIU2osTdEWEdpBz2IpTdkJ1v1u/q04xIraAmONM
K4+Y0sHa5rKi3deVAycYmxzftrZRn0gtbHFecXs4juSQODNnbF6R6HqYrQemmgJ6
VyToSw7MknsZtyrjgZFLO1QbZ0LhI1Jqs4cPX+o0FESUXXIniLMZq1W/BzXdEgFt
wIh2ThJ0FUZZKBaBfuDo1UMYh6DRKFR9+Omey48l5j+bgmTmhnYoxZPkUqG7+xYr
AywHjgtStCxkXDswu1vgl7umuM1Pc93iY2cEwSSdXL9K62/KA7lRfVreYNaD2axs
ttV3ehUd/qzaX+QijAFWde4yQKYqxLC96S7WGfJIdrtLTRYAX2rA39F/Ph5N9PKl
`protect END_PROTECTED
