`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Je7kwPHpsjq1i79cOCDWm+b18xYJ6uS4YLW8BXaL6Aculu21Qm+bxNDdmLaez9nR
2i5B62pDYUfWCTigxJJyzuhOKSR3LiKojd1uRatLD0flN7tTFLMj8DzvuWA2W/kb
kxNxBE5Vt/WRPRWB/sItpkyX2cPDG7bOL18tn/0ADu6zDn1Je4VOa/mVFbtLlxYS
5WZNrDvpDPyWWgjuINLRWsQ3mw8O0obYcffDu3MMW7tt/3LhsxA19s61zNCrT5OX
2dvOaVqEPNiW2wFndS6eP6MB1fYn/9PGXeQxMvSrSN+dSqdLP/SNppJT7JdOfZuS
yHGZup+8xeijiMSx8njUmeGXslgtEy5GWdwoDyfUBDxzGdp+drFnJQRT0WmkWjBf
qZzRE1k05NK9+TIl+NiHhgGKja8xuO+gV/EXeHLbTGZBrEp0J/kBpLhyRmbMz841
qYp+yKR+svQZSJoGIBKlAJwxMq1PkVVBffOHvNmXtnv0P3xS+8Za9UZRt2YHCNEe
SzrIU2bv/IT+/qqYg4CgnyYSszc+LcIQXWF1todqNEdoD6JBXNC4y7KG3ydJpf27
y+HXETeZrJJ1JcTrZQ/2THW0IazWfA9mFWWV3duVj7+3WMrzwycHZYbqRk6KoJoV
+5rjZZ6J5GZt9B8Hk+BL4Ao5ZgSAiFrAmkLmzIMvQaIUuS5Uw8dyEW7qqwu0tMFN
26Grde3bpu9ELGDBkVYe00Pm25QA/ddT0bDGEbP79o6eU5PmZIU8pv9dTz9q6aKB
570mMzYF7tJIxekbCGp9ZuRCE8X7Q/UYWz7PJq1vKJ4coTGT9cg25YEk+C4mCcXj
6K5fF3+9anDDbKKrKGzv0eD8dVvNhAaqBOaoXqqJ6pWvjchfhaNI9sFoFZrOhkX9
y7mgBE0060NdBCRZxrX8pflBfzXENCsJvDmitskfxQAKrY3p7L/EmSgZxZ8nBURf
`protect END_PROTECTED
