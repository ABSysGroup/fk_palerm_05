`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tlz5uTvxKzB+W0UQbhRbtkfyAL+YMh9RWvWEuSN3NMQZyqztzwKv8dmCbNuIo81f
JlnQlDEYsvegoYUwsxPCGx72wfLzR67l9Ve3YcFV5zJ9T1Dh8dvwXpqmM5uS94z+
pT+Af0hCn1LXDqHvx2WAeORokVy1+w0BLDoSTu7l7Ve2NhWeDsBTu4EiM41Uej8m
xjJyBzhlSgwOQfa4W2bpwowX6DgK8fTnatQ67vw1VQg3I9ClLW29IiIv7AGV8Yrk
`protect END_PROTECTED
