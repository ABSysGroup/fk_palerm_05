`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o+D2kTZTeLFVxfTQMeQeC7Opl5fPTvZXRrbTBF/lC71O0Jbb4VuP0RygQkQJdYTo
dc9WXHMeiA87BmvkeBfszyHkJ3SdPN19H/WhAkzMQjbYKHvrebePd3+eFpkmVx9/
/DU+gljxc4bzCr598q6xDPByaFUxWLEGoDW5c2qlbakpLwYsU75UdeNizzgbc4qP
GWyMqWeolVPKCVKmA+kPdmNIY5p9Ks/+F7NDAbqODcIHkpr2rXCWCFml52sJfr+l
BPLnrGp+hwrKsanm/W+cdvnf6nTJxhcIqgZhAT6WSI0qjTjF8pVpFFW2UJzC9OvF
WTt6fI/yvURpew/5pqPy3Q==
`protect END_PROTECTED
