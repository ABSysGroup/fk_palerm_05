`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ax5Lz2dyAcLRwlz55Ke73yZFVjRBCEnEliwt3f5XltcyG1YUm/Pi5Nnhi4klwZh+
LPPsmOQmwDTTpygRfsu73j1CxiScNWIBTcZ3Icnbx67lrCk3xkXmFzghk1Jn35cd
wUVK6wlxomGWBSj7a+O+5tyq4Afarln6c0+9ZFgZNF8/zh011VRa1IfoMhEabsGz
EOZNUgFbVLm9jgjBFhDnobkGAT9yCpPn7QyoIFOcDK6h1V2m0zO5o0ngaqxTRX2b
SJ4fcQgyHlI+nuAQGNlbmKlPKgCuKC6MmQ/qC3nJQmLvb3T7NKGwO3J0KELDAuOO
ygyPLA5vnBg1vHvU52leA44clrNyXkkcaxAFV9VUNvahVaNYKwiBwDJIWbflxf0c
VIvWxxUEPmnuC+55PggPNuN6eWCf/xWUkUbvdQsB+Ma48oivzR6xCVkkzDkUyGJv
`protect END_PROTECTED
