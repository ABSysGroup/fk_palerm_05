`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c4izL3iUJ6g3mmTgUVMRsg5be2XCI5WnkNjj9xN1ZKBG2vHDrsr0SMl9m1wW9YaR
87sKwoUV3h/214ZuUUsKFfDADuBk/Q97zA/lceKjDlyeauOQCPEN7Yrj/7Vwq4N5
3PIV4mEIc/LGVsO4NBo4cEBnvIA/ATLi3jA/PekHGJ089K7kZskrIWRsvhcJCuLy
DrWdcMt2BV3jtrLg3UyC2KTgOO6w/JwcLAbpZpmni1LPJ1X1VDucY+m3gITNVSLs
9VkmfTCkS+iwKq++QWurAA==
`protect END_PROTECTED
