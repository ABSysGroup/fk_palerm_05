`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iX7P7eoo/ym0S8S1FK6SmdgD0JTjUbGLvWTd0yu845Ojb17djy3oP2jcd3jdKp9d
pD+yGaAN/Ak8JQ2hsUyh1h4kmXA759ikiMRDS08zMUMGNK5BJgVCH3AAKT9VUwCP
SIOmqs3LsgS8bDcyg9CEvqvq4Op1APhXFthR/RRQa61Cwi0b7BrOcrPHDDyIDeI8
9eakuNbaeZlBUmKVa8KFqSE1PpL8r54wEuGVVnSWcQ+w+cVpqW7jDKTCUzKQMk5C
BoZmoqAkZJI7MKxxWeGfr0Td5qI/+X6qcl5gdTae/7AEP4g2WqJ1utKonU0ViOKK
HB5qpiBuUHrT7Ed5K/XZEVJbpCXWRHBLIu9JeMenEAVO9sxTvsm+si8tlLmdNd51
qSI5c9TKNo1XDiDs24r0jPHe4MXv3IQC7E0BI0t7tGg=
`protect END_PROTECTED
