`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OPiX64xMHPSaXAGe2/VKwxIVH8k8p6iE00KeocfughjeuQJbAZfJ27EX9SKxsBBj
5SebCZPdVGjGpoGZ+fBWHpNjHu5Tv0dZaq+M7+ri/Gc9AGV4hs0tvn7EpROqjmeD
/Kqz4EFT/bjrOAAk03S0MgjHEZZzHJvfbLDU9zpugboCVb1roMGvy6QtE4rVzfqy
5xN9+NIHEDVlfvVrWPognYImNzJIiDObn9YwwqTh9KQZj5fMczbsdUjfY2LP83Qy
UGoNB4ze/tQJE4g9pwc1tmwzUMsqdABvO7TtvDr+3b/jNu1KWB0gcW6UcVJEJ9rR
VETumL17h8RmC+GimeRMrA==
`protect END_PROTECTED
