`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iOf7RF6piY5TrJo174VlV/4vh6rz4EVLACvGTEmAQAOskd+64hAXVlM+mvCFyziQ
EdbwWKycjIVBqI6S3CG2LbixN+CwzcqLeu3nTsomrzm1zJpyC6Sx0xuraUP3Onfz
Bkm8UO6/enb9WrLbw7qR0sXjwUxJND5cch10vc0GBghdJumiJqziFeHic43WXQ9m
VwYpxfkmQeZrGDA9N6LojAxWTKSM+vBYw3PdQvIzfp6THVJESpoOS4NhqTFTIRVB
ciVfQCUkz1ay+A6QsZeUBn4kHL7rJlFUYx4/POcFy2ycVLwR5fnnhHpRnjNBLo0i
KidMlFNb5MiwtP/ZPacWN+BT/jcvAB0CCcYy6GHPvOyC88aHkhCas4xBQxS6ngsN
xHqY7/ImjDsMLmsSaFmUR/w+zKyuXxKPHY4IJyapv+y0+rAGSnUERWg5u9v/Ih6Z
iT2hEMYm4lz3r3y4nXANNd8tpwTKwNZsN+CmfVYPF+gu82etscwItZOjZRokSQhZ
t6pR6XEcgKOC0fMPWvc/CjoPYjo7YzF5Z6mydFUO/P0dkOybZZzXFAB8i4gYmFgH
0K4/c52ChtOsGO+AuyosFI9oRUDyI7c+ztV8wUqEZdfgHybbRxcEcUNLYlwAKUi7
6QJmTrhweKeq7npohyp0TvouB22jfLLAygp1sNMQhRr1FgZOCRbifQVXMoGmzb8J
qInCTDPAlAWCDWUZwOSw+X3EuPeujX7lDuisar8QvAt6nZ+oAHozIRpz4iRXNBCL
txpzo1nRYvVYLXaC3KIWqzOZ4WTILEKp4HG4H44or2jm6QKEoSJhPYwW1NcSsO6W
8h/ACnXCQtz5rjsvecn8H0GoJ9aACmLAD7AkhNdCMr7VP0LZo8XG2IRMYKEccetr
+clxx0bWpGY69GN45lUIguyE47yyBi/0GI9W37ShQaJgeKUVxck0lJGe9BYj3icm
`protect END_PROTECTED
