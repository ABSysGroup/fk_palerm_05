`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T9s9KBpKvPjuj6svepImQMtlRKR32U6zHdK8Ok9CekpnX+e9zuLWbJnhMjcBI0mf
gko6WDB0N84Pqr9btK7E0MV5Y3I+bsJ0zuEStTs6CjOqoBdx3Hx352zSIX1dEM15
fOcN48JYUSlHY+stqFW852IuDF5pparCv+AhAihbmVBZFVzuDXe8EdtPnBYDrf9d
xY/flBhzNiIL1eX6ZpVbGL79UV91Rm658o2ch5eFjExdMnOmxwIcw9AeUHMw9qS4
FgwcAsM+BgbvEBm4mXR+IK/OeeZx9RV4GAPLdTIN/54=
`protect END_PROTECTED
