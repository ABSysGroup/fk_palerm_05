`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V040Rp4hL09FroSOHAfHooSVGTgJwQWi2dQFVzEIErSP55eo5B+cesIeg3EgKE0g
fkjWoScJoqevyELvyLq+k1jNQgDtuj4cA6LnqA4GjpSnEv8Vs/Lqwm7yIvt8U5Sa
mVWeB3jTOkHVeSVNAht2pMApvcjqBdZ2tkgxICw3n7Lq8dE5SBRw1yOUfAzOC/U7
C3OIEv6D7kwnj+G2eiyF33owTodpkidA8isidoi4uyF5i7ItQL8fccSytxhuHvxN
ptJPBO6RtKKsDP+SmCtVoO0P/RhFUjMIk/62wf187Kpba7AZWVKwZR9dSOiOwBao
bvQUEXNrZZWE/HYJg9GMhzd2emQNCyy9wGkt7aFbzhragH+7qnGT8ztiqVhfoyLX
xkhMgGXY66orl4sSkEGJ6A==
`protect END_PROTECTED
