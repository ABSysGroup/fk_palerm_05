`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9urN5WLWDYbQ9eSrPgKafOBQkb41Mx5MyyFHp5Hg2w3t6ZM2ehiMkgJoGXt6O+bO
jEyKohVI6x0e6H5OQ7aEdo8YAurzJj7u2qgJZ6timC+T3LCUv7go4xSZERSoTcst
OvZqwNXk7HYhKzaya2YFHQktyR6rsulF4N7fwiz73/ae/bB1yA8wYdPAYq8wAnku
xkyK8BQsltbzd3kd490tgREctfOfrK1pbT8MWEeMXT7A7VMhs64PwRmVfwQdLh56
dcha7RXAgXMSBN2+fWuSV9KH1Lt7axopXVkeptnIYBMMSzLrx2S3YxYQpdAOSeMU
U2NebVlBWAt/TePRS6RilH+1KIPTvk5YmyKSDillZKtUU38mBDVhgLmjW484Sjva
oeDiK9sMe4JXkfS5AiFuRK+eAcAB16HHWvDMYESIdmDSgF6DXeikUAUywbl7P1iI
FmX6zV+mggrn7+nnZWIm5LjfdjOZpl8MWl1xc+6RyqLM6M3h3H2WmtQKKOyjn69t
Z4BqmdXZ1ezKYYswBfRrSQ==
`protect END_PROTECTED
