`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oGom4XqEHFOWnPHQoqpC1Y3hXMPWyw5Aqw+WRjxqp29LFGLQOZJY2AVZj9+74bwB
pSlbP2V3TvJGwndNeTygLQAFW49rLR7L4Tozq99MnYlcidbLuD3zY/HLj4BPt0da
JU9Mi2atNUmdWWkcg7WO0oecyHGeUIhIbvllA3XY+ywAC0K9MlaAI/S4mO1jNfrY
whlj1I43/zjbzIQKctbA3amZMVz+6dlSTpnFskzWT4f31sGzSMdzBbVn02kto2Kh
KMDM64FWX1IiduVqTX+0w37lwzwu4TIwf9nQPsoF/ms9/QmfBfJMdkZFtCwfZXON
1GKeofEZlzHJ1xcgvVd5tRWz0oZnizu7N4cBkTd21Rvaj2JAbFvOm4wxmIV/FQff
2WQVuET4gZgSNPWEUOEoW8XxSCl8Pl3NxMn8RuFrK5sq0i192icc21PUSJIH4JPa
Qev3bHu8+IzPpWxdkuB42KF43LFO/h28yiQEQpvlYU8D/MKjLJ39WJzxBMSJ6gTw
Z5AsULK9oYEStbREY1FsY8+ESKZR4qBFjv6qT2lP3k2BiaLZ145E7RNsKxKfkWpB
87xUimHd2qPaYYrd4HGyB6bvNY3dp4Sv1gjgDhh2yjBL0BjJFO8BYjvtUX4qIY8g
YRQFCE8mGVI8qmHRvHYr2M6S5pPsNF0RFxfa1Et6g2gyV/E4uA1P2wlo/HGTgTEG
aB3ndZyW5UhA+mrep4127N89LfZ84tF/aP/sqaN+NKS2JnpC+JMsQ8Rr6zAEMnL3
xwptNyK/wf3T8+idc0FnJNl/kcG+NcSrv35AcM1tUgn7rUobMQRTxwiJ3hpBK6Hq
Ba0l0rS71hz3wwnKZ0u3C/RWTizd1le6rN054UzFU+hwXVE9k2fLfAPU9zJvRxFU
YPwMdop3jqh5NttJ4TN1qbI0fZnZhSglz0/KoY7wap2CM/4UqBu3kbTiKkSXBAUC
e3opwwUv+WzgBOER1f6jvMt/XMJdbgTDKvgkpC33iRXxuREr+5tfWUkPEOpvYjhx
RlJVri4xkS+hft0wBgJKlHbW0lbFZxJemAncZMp3nJhv1x5JD1/Czo6jgHR3fey0
vmRqhCgfxoLSylo17A2X8Q==
`protect END_PROTECTED
