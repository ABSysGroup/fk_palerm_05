`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JJv2ZYxI4aKki9HajGANquajSk8Nsn7VMVFSjJaNa4PB3+ThgnvdTPpP/iulDRhS
MVlMH81Q8RhRYO0ue5vUwv4LG/yry0txewjYD9TJcpf7eoDqBWoR0PKaysjdqywr
yqVkSdxBN3i1RDi9Iz43kErbkJV1ZpfKo8mJF9UlwSgX3MIRmU+ZAU5lk8j3VEzG
mBq5+YFAcNnhrIQaac8/TAnPtf+U2E/BODBwoYc9Fq1qArQEu4JiZYIAUVXvfSwv
IhiGWGf2riTY/DYJGZRIwAkpdtZs0xNR5JOY8TCnU0/ORduFldcLvaEWuP4Ss6Q4
eCe4AQHePBXbNx7be49+PgpofZr7Z+wGdRaiMxA6e4zbyidPxa/wHptrZikWoyId
X91/ezY5F+LnnOsjL7KsnkKqNgc0ZUxpuFNmaoKvcmzkgj+jgcjLMSlDzGKhownD
bFWu1+CSKpFBnd9QYMXA3o6JDkaa8iT+ot3knhdLp8dbt4ys8lXQa0xefDM1lE2i
WMYvvGHO2lyjL4WV/9181TaEIrK1Bo/WmwYRxULLcfGeB4zY7LqmH28s/WjuPhi9
1urC5P3TAODuVysuvQHMuMXOYfxo5Ks+fYRSmiYa3AfFYu9oaOqedKV5PdZss1P0
OWdRfb7+2rWx8nvhsiiJHKERtLkTtogow1zyHEMtdcL/qfLU8J1vp7lsfYhGVz4h
znSLJnx1UfpHNejkmww6lESJxQ3H02Hlo02JYpCh5NM=
`protect END_PROTECTED
