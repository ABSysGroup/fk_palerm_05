`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GENs0u8xQyBH2WV6lorfglX5B/JK4dik8izpu39qQcM3ZUHjItP68onH+DmrcOxz
4XBLBv5GCJ2+2q3x9KlfAMvmh6LvEu8fRqoBqwQVgz6HBOHiw8QfDPn4QASpGQW4
1sK4O5PeLnMqnaoB9SF+gore4JRyJHji60nqrZ46pbMLpbkFjR+kYV1D30VozctI
RwbXjgllJ9uAcYNJdk3+blyweR0SeGZVQkBU4kxLKviJUP2hqFLa/azuJoXPE/hk
pkIta6YX8OUQ7yDUuvLqNd1yKCzJW1FawZ/G+bfyTkkYwHvk4dU8B1Upbv9YBF7P
aOg4/wJQ/zgSURb0cKIDWTN6gBZVe4pvBirQCGRGNJZd208cVjt5jLM/tOkLbErm
u0Mb0q3LV9Ew+M3r2TYBv9P7PAfBN9NCzZG6EukcU/Yk0QWwkdLIGB50l2auWZDW
ltFjVkiRUIXQx7HuDvvCbI0PPSBudNYDeZNyXZz6KQ8TmWdLcuAb4i6orrGdMRa3
lCw4tfc529LGKU9nbQDHi1QM/L9GFJAPbNlk1GZTD/dKgAqM2BiidcYw5XNNATvS
snp9IubF955T77buy9wQ6qKwC1DdK9l+ExmxOCR3cZJ1y19XIMJfFQvqE8QG5H0n
K7rl3S3WeAZjgaBbfhvmWG4x6MBHoQVxF50mOPK6/ZAxbSPXX9p4WkLNtdcNjF1r
uGzlZ9FQIH1Z5YNuPvAnp6D+F5UAjutdEkqPlr+ZqI7jTVLd1OiEG2WkvFvlHBEN
Kzgfcz6+10eiMbarwZHW9Q==
`protect END_PROTECTED
