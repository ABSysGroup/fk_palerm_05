`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ntJQBS1C1bnBi1yEiAz/8dk0pzDh3pJEBjZn8D0I3Wi/sspS+8SjPggEvIFLZIF2
GfFV+vCTx9BAZGC6WeCCMQUy1h3xj4KKh6QdQX2476rjvwB9TE09Duy71PZbd/Oz
VcXTkVGvKOxuzCEDlJ1JTx425FKenfQhVwgkOzg4gLx4nmBPbLHbFZSuiG0wtmwZ
UC7TanLvy4qRWTlSAl9HNZ0gLuUpyADjmJityYVuvXOpzDo7j7FAdv/BbYfpShgr
2gHj/nt+SmvVFHRYplGKcv+TB+eu3QlSP54PWYt6IJZk7u+9qccb7AUXHexq+Me7
4BW+NEUXirbiIY8rD9A/zU51SXDVBwfZ4jNfgXKpce/lwyj5NlwGZooUrU6M/UEn
yGPoX6eVseSFegcV8b3mtRZkH2oNgv4v8+MBsA2dq6q9fZ3c0Vvia/kNWAtRKOC1
6laPqCKk4EBfzEgJhCZ+VhQiepsWSQtKPjuhhGw5W3jYNdEFyNSBBmPX9EdljYWN
yTQxnXR7EVrrFzxDjd/1YgqgWuTxQtoErxID8GF50HOOyZFEAz1lBxYb0wH6s0Xr
lEULPC2ybzKd3RFcWsckAVtAMcNotCgJappCJTv127GZ/KMTBsLqOi6BUDg2rkrs
J/qNqd6ECTKsvCrXrIWyrXTVVH7u7FFAKslKt+W8s68HulfnjiXYfHizPlWX2eoW
ykssIz1tHhBVmkpcFoBOvBDR1eyV1ywikY2UTtupb5Z+U5ShSfmm9z3q3yFQBWDp
0XBHIiPXVV4imMxWkgo3wnro3OSSYhZLA+JptgNzyRA7+V3p8SX9+aXHFnO/WSma
eNpPJ8ux+yt8MswTOrTQPpTyvryiWP6ND5BjVbuPepC1Pinss0Je7ZpWJFLyFFVF
W1ntPwRWk9ezcTgHRs6vyx28sorFxLbNL4qcEz4gEhRC8/WONLliUM0Xx46zGfwI
`protect END_PROTECTED
