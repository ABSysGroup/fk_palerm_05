`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3dLJKyfD4hAVPCiFYqz70MYDVCGW2SIn6CmNIRkTFTIspD8PY4KKorLiVkADi/eR
rbCs3KfN1/uBgqSrTNhy7rgPjAlqO9tT4Sd1gbKsGAVCyVSzDFYlKYevalrmpdqQ
ZT548RzPF/tfYHMKPIDQ6bxmh3eGMylBWBMulXYz9XEam5DuV6fjSrR8yrai6rrf
bCACNJg0JRlbmSeHjjbvvlmP/Pv4Y0o/QHvFGPAzOIQm/Kw4IlOvdIrXH7JrD6kU
qFPXEwLM9qy1jcQMjEnCrSnDt029Z3k04ifmOWDykDHkE0LWPy7GNWeZ1bBBQWrp
Ara5cBaOvddUdZ+8X5U8AdFNDTWtlgYinFoaAXnctDIa7uEZ5Z+cUIHqqZVbSSR8
yIYSALKWX93FNtvm3UraDbgo18OsHd8NTR1vBOX6EiV7O+4IMQtNCKMOQwrif1kR
ffxnOoUVZV1lLGm7rgL4fPmlKKJT6wDKXmFR8ZutFgYwUVrdYXyEqQweAQLjkZgF
/k7LNeufDL0qjXvugw9bk2LGqrgziEew43z6+D4lveFbIt7lIR/DznpD605bUrMQ
omh/dsA89TxUUAK1VjqlwA==
`protect END_PROTECTED
