`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qmMHVtM5x1Rw58eHAHITsgE495Qa/6xKSUMKPRQYhWD2GRbs0jcBQf8AleSuUzll
nWajP79ZizZbfj7L2dV6Wpbk9M8MuP0AMbrkB6g1JbAKkLlWYEUkrwj30i+VUnY4
uM7q8/tzR42U9BroXTDRq6EOUsMbooZ4vx7IiWPddJ9C6V3NkYVjFQoh/2lJ9wbk
O1ThAsiHQs2PscnA48Ly/fUqp6RQ3UUt0QxjE5yhJU48OL1XwrSBJtgNw2xjEwAr
cUkPni09dOTiHQqPZ7PN1quT9xUzR9aAaZhmXfWnTa9/Ymn7eySnfT9+TIhXAbov
Io2cCPL2pm8iXCH7+JIVoWj94rPmwPOBWiyQNo+XnjHysmKwLP63qnc8uO/PiJv2
kF9LtPFRqgRYSwKrJWZ35a7ZLkUevHvYCgyO28+lBjQgIyQnC1QMYD+KHpHZnMgV
S1MOAeNg6iQr/pZ+S12sn8rpB4UNJmj8KB+oAqFE0Vc9rzy9kNqrf0MU8IlvimM3
2VrE8tOim5BbPo6Fyc5HYuhmceJyRT0LAlveOM7uTbnwNUq9MP0w/ErYIoLXcSEW
pEFAxcxgzKjr88HEFF+WdLnwLasOknVx2VKFwrUj2XKQsDXi3d9nR/zcsEb59Bxq
qx2vTHE0dO31bLAyFEwYbVNXumEx2gutkZhXX4BA+qOWNpbWld3PyRKcWqeZNIqY
zIirBziaOLn1/oD97pDDlA==
`protect END_PROTECTED
