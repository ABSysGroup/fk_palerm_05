`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SLMAOZgxTjmYPcXHaXwqQFM1aIl1WCqpMPR9nF44TSfdpri9eoy39XtEJezD7r7D
UQhFxfdO/MBdSwFenCHT3aYWfjiG4U0gGMEpa/ciUpQlfkATWij6bMEyDVciPW6V
GSminEEb+iir5HaGl6kyrUB+78PfO8t3ChHupFdfjPLE+Ryfu/iSTwXCN9BxkFRX
Vue+zLOySPbRl1fEdpG39bzv1jbacirt848iEMUipx3zaCjYBM5sd3JAw79KSH09
L+P5+DLkY+5od6ORAwYMlI/NSYcZJhrENwp/nTF4n4tpJaXfADiSE9dNen+D+StG
z7gH4jB12nMEeHsCh7l+2imsMQZz6+440i04BpQcmwRaHYIzcLOxMjrUepOeNm7l
bx3mgodsSTEBwhbY7t/h11aJi1BhdVxyXVjgnMBd6zPHxUiOTQcs6cSZeCmJYG9+
nuir81J602JUw9eLHLkxRt+5gQwKGkvqLo9nmUgYnEo=
`protect END_PROTECTED
