`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sTNVOer0pyQSoKWgfu8hf+WVGadHZX66bU8tc77rdXRCi6HAt2+TcV2Xzt8ydU7O
V/7qNINW0oX7QzeauG9bE0VrljfnHypXQxieetSuP5/T9waa6FhlIggMHq8tDBIk
gHdN2jgeVD0FWw1GgRJK2RAVD0fZtFjClpGcmf9OactUFHXqjSawi+y0V3Q3XMxp
CbjGd4a1/SUbfDq25XW+KNvLsALsH6r2BybfpsYCjmDweBNMQVjTccx9AKR0FAUw
byBBBPtMmwv7h4iz8SYJsIA+5R+cxgC5GB9rm8fiiJkP/P/GVklgFWhldFLfsAvH
RaR/qyEjg5w54ieIPUnXso1nuBhw9Qf+4vYgY1hDk+aDxiV8jke74wIW+Nv02Sdo
KxOA0CmmyXzoa2PyAoah6reyv8OTlUk60gcxejDiloEQV3sbcNEI5mRT6glY2cTR
HiYMVHEW3Inp9I1Q95VYTvfkEEh2DfvPAC0BeGVssAUcuQtE7Gq9nKdqdymx+Gro
kWjRnG9CgeMLFJvo0R2Jw0bVAmuoPzxtYjfbOLxFTwFT+VGbUjoyVhuUsNy/C403
YUwCC8EjDs08gV/AZ7YQSaOGSXERMmSFJzrPHz1r68h5SJ/TmbF6OcmGfXX76moI
9Y+0lb6UIbVRwRJJeF9rArVV+ocXvsEqokED4GIBqw0=
`protect END_PROTECTED
