`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QwMNnRWqXgflLOaR5i2TzjL0sydnJms5VmIodpA2iRCwj0jVSluZsCfeXYABibJG
fz1t/w9WhWR0tBcxICNymOYheZnqp7nbJpn0i0sK24eqCM8fmLUUmepWrYNr1M1K
iK8X+GzOeYTAuGgY0W0MUg48Ap09mAz3FXLrPHcusMBS1TLE+JApjd2sWWNlS25I
5iITOChIzc2n536mzGDm4VRojKL9m3eYEsBYS65GveO2YlRC+xVM9oe6rE2eTpP8
ESkLnqnZ4nM6ylMxjuVzItIJbu+sy7SjrXwaQz1MozM5KC1aEfVuwj3oBIogv18f
qs7Sq9R2cw9cLBhTcb9TchEIVqVOhOX+mTGc5TWdWiFGaO3x/VHGWOCTFjUedm6b
MMujyFJsgG0ywoFRL9CdCtWP8RNJkzaMvsqlFC1DbduxVAOnYKlG9/XnTpS72tGi
Z2gSU4UMqYbPVm6GVCKrKf3npMMjkovBDsgH+H41ziHz5K6BykWk44VlnnptBKa6
6s/naFCKSJMq1cOIAhZpV0fAzimPrXxO5AUJ+qPfOkQMGdn38psXytn2nNCOzddD
+DrBkQ0gnOAzBZpbE3nTGvpYfUUhzSUXqE4lXky4dPF1XGwrJT6apCKZKHcY7ZA0
0j2MFYg3l8hoRcNTRL+S8g==
`protect END_PROTECTED
