`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QZZNHosKd10XgYLyq8ZikM2QPxjps6Bw/azPm6S8HAwNM9Iphg5qunyfeD/tr0WS
NvTFpi0f+DlNqhYqH/I1gZE05ofbpt8PPXLBfaOb9fWxtCW+rPCEuhHaJgXfsqMx
B9DQVnOMRBB4U2kqLtTq8LvcFiOGkEFK1FtAWlEENBDROiqJ21KavaKhoWkT2Fil
qt2+nKK5Snwp4Hy5YvF/PKSf73Mo+U6ZvIgP5J3k1qwyMRapA8JKLNIKRYXpqEjB
DrUeIisvs4LGR0roF4hIV+iaDGkp4p+8jhCDIcAjYfP84Twr22XWrfOtgdBFRRXF
UkyisUf6drR1zmg60k8E6LLOVItQXscN+SlUVMNpR7G7nXvtdHMR6m8fxXOnZ7Rk
30YvSQy8cLRAVK+z6cAJJ0RKp3Gkg5cpQrcqo/tgEa2xl+SfV6ldw5bLx04w0gKR
xu5vxCio2tqxR8BU2Ww1+vsiZfQbmjEQJ21V7wqM6fX5vXWK+UfkWIDTggdHaDq9
mPnfv/NpAkCiUufcmmg00nGmWVHo7AzAKtxDxG/LH3+9AUbUgH9B2twprDSRfRCe
+iCtlmWswtWf84NuyXFsm0rR6UQCgPRYo6nklweOdo37b6upVvjs7WnEfeUV3pxZ
1jvUm+m/n3rMaYEnHNjJQreVtCJsSlF8VtuB2HFMyd3NULeRbmmbHOhqVhJ5Jz1C
GMoceT9MfjZnUHSucON/sQlk51qLM2cc1WkCTLxEuoa4HzRoYUttxSJFtzdN/M5j
KKE5XSqyvEbmH3rin7fREndLwo1ho4iPb0Yvnm6pmjXC0emPiN+z3IZIX+7vucwz
bEPOBQ4ziJH3vFsB7Gy4kWHnHtw1F5WAjB6qrceCwPbGi4sZ/jHrqYdhKIOPKuUP
/zzGyYezZAOcTb3uyPX6u6SyuovQAW8/eJ12E1H9K9o0DUJBPu6L04AIXX/PUnAB
gUSmksrebXIksYDD8YNaCBpYrrFLMhMh3/wlttNRR3NAU4P6tkcKwOFQMSiz/jO8
LUScsfzMHwp693on2KFLEZoH3VXCbMjh6VsozLq0jCymOsN+bQuaBvGXJflNH3Q4
12AdFY4ejN1LxL6HGSQelkq9WEEkkmeQJTrZENhpMX3CZfWzl2NmElM81ZcSIsso
qPSQUaTfYdE5vV/YfoT29PVpCg9Z+wlrjnB+/euOUKIP34BdUcRC2/tE6yAnArsL
gEGf63rK6VvBLzvv1dUv47iEirvKIdUjAqqwXN7+nWi1xTDRD3r+ehnlVd8qWXJj
HdmpT0gIaxG4Tey9aRjDX229wgTtS/oAVZidjFM6tirVjezwzOFHq6DQoDfeuf9g
eYs7Xf2ZMvBaq+859eln9idIreaV54T3HlNcC55R85BXrIIaU/ImtkF0rU2PSvlm
dKeDzVLRKdbs8yXdDaCNYJo/GwJ79/f/WS+KFUB59eSd2Y8pS1b8XrHfjjmne4zm
56JFsEhmuXpjocFKxLoG0F081mujjXb4RBPqvxzQwlivXDnkNf8iSmxQWo+im6yn
Ea7Ia55/iSYTh92HB0WyTsPs9TAQn/bJZit1C1tG7N1Oc2rtzL0SNuzSjTjAT6Rt
Z4auTfMYiHd3LUqI5NJcdyrQ7mlPndBGuye+9qXWcyyC/lu4lu7dJWYIM3gdTyIE
zMFbg6jNh9EvFFp5+b4Ej/EBJL/NDwqfVTcYI+oY8139bAnJiZUfKPeByJJo/A+H
ytLFQ07r1bzB3i+SWm8ExwQJOPVlyOk5Id8V5yYgOyOtsCaN22GCF96I6oaSTeaA
eyQeG+Gk01/xCyXqznN+Sl+4Ohq3YjYv4P8MHEHlwjavHBKU8iAjKzlLBmu7LFC1
gjzU8vmqz55AJa7nasftn1nqynWMGi4+t8375qDhcNE0hBxMqQXhZH1AXwVvnfHa
yiacyeAYD9ySvVrSEqE4K+sf76bSf/BgUQVblmfSUAPpsrEw+e938pmvponjHddB
tOrNjFj48S8jO53qaN3E3sxkPlDS5hRMW86GjpY8XWe3yLYxp4ldnFIa8p8QXubw
rT/tdDRbDbQXO2jlaJ9wIwK4Hdg11jXelHEihK1Vcp0x9LrLlBoMHJ+6PisVeMUb
Zj9ZYitWACcC7zLSFIP3J0E8TRPnUUvUWCixML5vH0hZehjgH8Abd43YOtS9lMNB
93cWm4027gI6DzI7dS1a3S80Z7a+1P6qolXY2SxajnD6JXGZgXPwtC7mAxG+8iFS
ncTaTa9USK0dlwrczww1+HDRLEC1iaNX8iCjMUFEESQrfS4EtxycbPvliFPZ+5+I
n721rXbJ+H2/8cYlMB85LOgD2dktt9thD5dHREAzRhWj2otIGeq9pLOX3fLVSF4S
JyWX1ZZclXbfVZNvF1O7QpETs9HbnjiSH7Fd4g/CmSfXtHFuA7xCVgV+UTRTmWH3
X4Q9XE5Jx+YrUPGZSqlnLoVuMyrSwcJ/GU3PbIb/aXP9kF9mDcvFJsy6oKihdoPy
vmwJsnxxSATkN5gN17VYJbvpgahyK6euUIt++QAhUnFa8Wc0RTLmpu8IvpRfrg6Q
LGZjKRV6ZofqQr+BoL+GkgdKGzvYe3GfYuaXNDnbaTJ5IocoGvP7iGHycRy/1OUo
gBuE04UJ0m3YYFF2bt6TaBdN73yzU5wLIGHpMwn4t6A4W3YpeGt2vsAd2XW451jO
S6F1vJwkqRkw76mSUGXMlqToI1LemGyiB8sQLsvBxCneban7yYdBGANim7wdMPgJ
C3eLnUOzl2KDcaIUTRtueDwapMVXjl4X0ZepXkpRts7U5ptrQNcVErKT+nF/2cT2
vrZ/lV65r/47vuHTRrZzHPH6TrkyIX65Sy/sJGXew/TWQjLUaeWVDb0SRHi7uBZq
CqBqkB7LNwUuMNU0dYVMuyasB67B43yU4daSxscoIoLeOt4hMjQJu3jxjvLoAMui
W/sASl73HbzLcbZyPrXfEyhXThK6+RWKTY54PAkWp53yJar3Rf+Ic0VZ2gHGCoBl
f2dcEXfgljs5aLVCHcUZzitnSYilv0EqaM8t60XAC6aOwk2pv5qjGImCu7rKk3og
gHc9cL/+a/C19mWssczhbSaT67yDQJyj80TqfspeZTHCxF7+BZoUP8EMGuq4EueY
fXOsS1m+WPjOtgLwVDGuz5JrWsRtS/ZysqzKFXWn/oQAHAqegHGNAROw3P+5hwpS
cdd9cbqKysH/rAEhaEzyCGS3FJe1Jryq6AiE46OG9ITSuIozeU8/i4+W59hCj7gk
Z3zal5HgUDHYouYyyTFNdsS5YXCyuK2gGwd6WU7FNmHfsR3C5Okqj5PHmwUgkX61
5KwoLS0xUaZVoSUGH4vq78CtZvqvRdb1XotykzqJG+fIy3tcQKWBd60tFa+kgErl
2Az6qt5H/MT7gmXAznUcQSyqQfhTpDh7TndiHQP2kl0iE2qpurlDaCqEjy3GjDqe
S37ymy11wa6r0xAtvybzrAxAxKHsCPs2vx1g3r5eEsz8aUFIW6OD//GJAVB5R0sN
IPrge1FL8PeJeqJmCddQTbo46l3bpbNOghb85b98FILFNPjT/lTLRz17CspVXWDO
PATl5Uwmy7lSk6xjUPHd+CskNk/jjb2QTFtdVf4jt6US9AIblh3/DWviiXLDu/lk
7Xwzb43Hm7hRsADnySVZpc0zZqqU+3bEp8UU7Axw903gi6CQc3zpvnB5JAndG1z6
hojh+Krwcy9ML1NJ57JdOkqmYBtTfyHYwVxOiIOvOFV7GNStSc9bLroxM9iUTf9X
Z61EzF9eYTGPUCrEDukGj4O/fWXHUPLdMUYjM1EsVKePGMSoywyx8+hIzbifhF4Q
jNpB3pCnLpBKmOvZT2uzisY1V62iYi4ZXO4rcCO7vfebVVDUet2142ETIojd496L
DDUfBq/miV+1QYwO2agaY7WHXRypgtEF/Aq+8q3oGxDCXg50E5HQMBhlJADv1fnU
WHg9K7ayv8cxSeek4U4lGQz70jV+t2mW0dXqxxXRwRRZDFm+0jQW8BM5liimZ1qR
K+DOYRWiNE2TjT7hR+0xx02Q2EB2tg11RzQ/WlRxujvORyXyLhl7ydpx5sc8HwF5
c88lvrziUjWo3lNu+wAqE/+AKSA+4tpBfCGRcvb1BstfEU2PpguijQGZfXdPBKIS
rt2Q5pCsa6rkReptJ01Fs7wWsBiFVUN+9gzHJpQtXENIGNENg4TcQ6YY4mM4NyeK
5HGrlPZKDOA0pSoTGnLbbMIATtFWEHM7/bZsG4KgVKhknktYOxIghQPwrKMsOQIF
LqbefOgPsynhNVk6IcpnU2Nx6AX59VBUUiuASAitIoiSeBMQTKuXikWwCmlfZUFN
mPK9wrvkQu/qchf1qFx0epDsic+N57QIcNEhX1GtEsyzT/qbdn+wow2Adpu3f9Ed
i0mTXoj6xuRSxiAdpecNvJZmcQvPwOI64HL1nJ8SYNo5bzTkdN435o4S7Vf9N2jP
ewLUPAbLqk8YgB8q+70GLVfmghZPf8FQhedXm92iNMW1egD2o4ZoOUDTF8vZWXZ9
IsEqN0RvCthJzG7rq4rRUV9bIoWp69l+wsvqJacL21FGP5dw6eeeWCH7yUhrmBxX
vkqXH+hmv33Xhkosx1BSiqrlyJvK8An9NWdreqD8maIcPZzQES6E58YiY2o0dvqM
tQ/1QMyJpLJqiPlDHuqHdHw9j59elQIew+9+CKBZucd8tXC02CwuPCSAJsusLLGb
Zg3jfu7eFCK2wl0XEWzG7aPKAwZhP/gyDXH2VXeB7YiU/WIi1hWXLX3cEB5bTjwr
H/zEEg+JBr4jBTWSf12oL7Ze+DPa79ujAWM3TGeHwXW+mPw0LNvkN0/IDKx9CwCM
pzG7lRLlMWvy2CTUEbLRnkSm0wycYNhe+3xCLeQU48WOMFNX+1I+Ie5H2NRd+RFG
FQIbIKZXb9Kri6UaWoNEDo3boWFH4fgmbDTUGsjfg4WsQwyz0q0WksibnLBrGcdg
ivFOxelSN8Fq+dRWexXK2lzZSpTf679kw9CVRY4e7WaQckEaOQxjT1DxQscjeR5x
zAcI9cNeUEGoyxqGUwneH/d0T/ikfRGUp7MIvROycNl8v/hpYsY7eOTpWSma6eL1
+dbmw0KaPfaBEexnITsn8OX3DCMrI2lL+S0Dp89DqOpqT2uKTbCI7q1sOPTaGGPw
h+b17TJ34ZugYSFamj7gTq8IzdX9vJZPVc2EsTFXnnWMnb6WBdEPlS+oAb47gw2B
po/VGGrnrN1tgB2/FjqSG02S0WsU0nvTiWaXDZowxcNJzc/uXKBKBpQDVRlpVhT2
8XngRQvNUUqw0cwkxlVg4HSf+aatpPiyNm+IzJfI8o2TwGSj29dJI1h7q0VAFvcC
m4FpIudSi0V9AvuKWnlqafl6XbC5ORZSd5/3BdQ/KEEqFtYFqFjcigaLWCogDFWc
7M8RYO/jiIKpP7j1d6zd/B5EjAOFgsNtmjpmegF5G4FSxtvLf3/CZB72DJyDur4I
Fe6GBI4zGsdWFOqsrW5Vau2HQJzAwc6RZHlYslg/Kw8Gw1QhTjfv73EYAsBn3vcu
JMi6Pa1o2SHBQjKZKdkEm70DHF7yLksn4DJP2JVFb/qnhZ6pICnD0LN+H/jfFIiX
9D8gcaciqwxzCe73MU9IpSDPFi3KrURK3paueFWvKeQK7nkvLvCPwwI6lNblg4rS
V6AGJu40Zmi/L2CEMDYPRXZu25MNOPeVXBC2HRcZwtIPJMwQJWSchnPbZrDBnWWq
RfsZPVySv//aP25KirQ9Al2yAc1wfmlXlZXkVBLtdT9K2Blhzn2lWupIGSVo9LIz
6gL27b1OybfCwAPxvqp1L7VsBKlIL+eKXWQMcY91ibuZerln76kxgzA/TwUVz4Pp
HSScOTWJ9PCbCsDE3xSxXZRe23ZEygcyN9sNQIueLqBYvSqcSIB3lsZLxjTpQ0yf
z2pI231RP2N9noEYI2V5JOYn3Ae4cvjgZ1H5g4Ar9qnFHE2HLIGlKq9dXsiDM/OQ
wkvWpul/pq1MbTmb78DPmSiCQlU8eDLz6R1oaN6uAzJpuzgC3i1niB/1IlldF+Np
30kFQ5OKPwpyPE0IxZ7CeJS1A7mdzzDbGYo22j2GXc2dQcCi/Itklk1EyZuzGQA1
BvcWr1Alx7FQePX1nICLDJCp7GhoFZBJkklxrvHv8HVQ3zmJi2RKY0NJnfXLAUW+
Be3BTKGA4KZf3i/u6t66jFhDx5EBOWjnBsz2MMT86M8xEJhvdKLfzgT7n1dA7Aan
nlFRcd1EG2/X5c6v6D08i6rtbEBE0uD9Uq8E2yQ6FfBz8AJQwtKCevE/psUYwc8z
zOb23aRjo/ZpEB7qy8ZgDaNYTIzgIbxoYgs0WH04as4jgJDtCbeLouq830r/ns+X
L4HPtw3FQ7zIF5S7XGbUsi0cyWfyDy5f9M19+nU5lYUXPx7bop14Ndn1+aag+l6x
OEGNwQJ/9UzewMhSr1LTHMv2SsKSbovmUaqlkWLGyvPCDSM48cAQnVBslZiWtfw7
iKxWjXLhWiilBXZ18juPHy7TfrYOIyQPhLTrkcPEqVSu9l4evS8ks+1Moa1befyY
yAYAFBW9kMhQ8fwZ4HgNFnf+hz2Fy2Q3aY4kyk2kRhRT18/r5L4p+ar9XNbmktee
Cshr66TWu8GahZDPd5rXmohR+pauh0fkB1Z0KnOr08Bp1gTtbBISf40/CDUPcuxq
mzIjKAo7ncNeyiDouf2PDwjzwWlExu6oKIh9q16kyiUkDg8Ee2ahEsZg0OkZZoyF
yd0f54dmyxZMe9Rb3yPij7wvF/I/Hjq1G5VY8ngXhxlendNfyYfKkJEWIjKRczC0
KnKTkkH2yoml7oKeHBBSdXmZmiCu8OxlltgXL41LhqpBYp4Gb2hGpz2ICQfZ+SpI
/F9cFpuX0M9Y6PQgMxL86XT9oiRl0G5mv51LxEzOybFhSOad26rE/nlnTSiL3ntQ
QgAHikPNv9RM3JnqJvLAB0pnmikMckf82h+0gL/RfnELOah+ijXU7Knfu2UqjcW9
a7Po5V05DaGMlIFxhxhbRdc+doE4h1o2zRpG0Bco4YWqN5YTyLODJZ6t7mgMm7IP
nFkleCdLaFMH15AOOlcvBeWZp30eNJ88qgMV/PH9/ks80dy+qMnjYFXRp2hC9bUl
/moenXvd+7lz23FJuXcp75eJUJNEqISHl51Ac9MzftgMTORlp26SdROmI7Af6BMn
/U9e+MPU6PW1610khDwe99tJoqZzl2CZssdHldPAoMegIoMb2gU5IruExHo5Jae/
CqeBO+emtnFq1pTuNNPc5B5p7DPMEIVGXrJz2b4b2z0pjhFZ6wunx73g28Maoar8
H7dbZepYl/+lH5Cd2s9TEK9i+BiQb1rKQDBngCq2+zJy0HxIaKJUDh6zDnhPStk0
/UH9jjQs9YqVPtTlisY7O7CA0zUw0yyBGI8G4KkJG2rxpURQGnFyCiekiu6rZxDm
VHZ5QGUEqCLCH8RmX2FnibN7a42Pcbr8jGE0+lQYrcGn4byLUu7MqRqTELyvueZw
fbSwbfK4xTo7kCzz06vJRz9/wOES+zReORmMMauwECM8aO8NTu/XnkzQwdIr4lKS
DTxH6SdNY2MkpSUJLPaiGDJtrNZ7ZvqqYdP9rNRQVH33zra/BCcsWqoTLURgHMgx
87RBPPNkMmqxxj7sH4NmIbAUccNMZF1rEtStMqx4M9QpObbeMi8Sg2AV1GjfkXSI
kJFTSpfPzdgzV1MLFyiM0d/+8bLriiobficQN6N7S9zJthvXBBNJe+NJwBtlAOYt
BR4XQdggz2Hjd6ia7q7fJDdLrsmG/q0cSey7TLkR2DokhN0ThsZW+RLDsamMA0n0
Gg7us7MmcDqS0VE6UDoUJ4DuCQaYbcQijJ9oZI0PPmIfa3afLkq8vEzXEGmhkAtQ
VXSP+jDvDMgwi2Da6MtCmfCeDgJHhYxPFQQyK7UfKjwM+CTQUG1EUUmc6g0W50mZ
7WA7CkViX93QrAYYS8FQy+jK67YXLSoeD4zhYZLiM+sOO9MAKFXlcc2NB8Ciqpwx
SI0NafdwJyAp9U6jW44+OWhANry9xmSDQQuqQPV48VSW9Eis2kz6zNQ5+04k66rP
cr0QGfyhJ1flVTiD+U64YxxQwMmSqmXsy82NZy5V/OurauzNJlnnis5QgmHYeDAO
wiHh3H8lrADLC+cYLvCIvbaf72+9o9tIoEx38sVqmKJlm2YCt0mK5ukZcxQ7RhNQ
dTPnk1TjWVB9wyt4hyy7i/hGAoBlJRgcPf75Lxh8grK2hhshGh2obeWgkvNPa1rI
8qhaHH8ZrSG8StogMqbagISyn99RjSlYGZmbSn0t71tzyQ4Qu3OU3Vk0OGSDRzC6
Qf3jltSWTKGYTnGuuWfMaPvxoOA6/I/ghYBAQzVL02JakeU2ipOSuZ3YQhWrbhSO
k+ysVhEG/w+sX5FuXAaZy28EmZMdAZK0Xvxci2dsfKP4UO7ezZB7+au1SU0WlUhq
tT6wCXA/M3t29r9eeh/i3lSmOUJ/MhubDCtz7Ia+F/NzFcVEKJWLY3/xsTSeeb5M
A2vf0tmgUR2nHzFw35VlTjPklGySWApw3jQ4lbk0zvJqcIzVwkpy2cfiTp1MUe8k
D9l3ba5f3BSC0OTrycEXcWPsBD7KoW1/WuDclCdEqYM+rn3oPL/zOZUUSZha6yC+
s0WMgBZFoPqekPhkVJ5DJ4YwRk6SCEqvv+ofCLOtS7mHHq0SFhZYxLFNu1xAfNyB
EttaQmR8/rUM+TmR4/mKIk/FYXIDLL/Qw/zxrzMFIAPhWQfx8QfmF9HysFd4UfHo
HW9LcPyOPC+s+2mJSJfAP4EHBges8krBuJ7JGoojJpPgNAGN/hglAY6uptgmgvHd
7CkbTBZwf84HzUv0pzVx1OshOnet5r/sdXyqOomcvjNos+gEm4PGBMT+LAfJQo6y
unbhsPi2WQwK4+Wk/YlECpDYEin2kN76+rFIVTN9FHXMtXaS4miDiC/DQr+UYflR
1BLrXZjoUA8Pl34zBGTb777dstBWNWXZaSZBknof7f3kIg39yx6xvJEV7kAUkBIq
FOTNTguor2wyMf3k79J1QcGYlEgrVf0kiiHp8diR/H2vg0lwKdsx7jmXBDoW8wpm
twtGaxn/jsSrZHaPKqkGIImT81iEjx5LNJiawBUZFbqHMPfVpO4DnyvsS1Fgtsnp
DnyZXDb5bz49E7wBCdrt7LdqPBFQ3bKWxhAVpxF3T8OO1rydFPfnzUEErQO1/+yf
5/1qr8ZU/a9TwIS67IslcPQMt0DF25/WxgXeL/HcishGnSRlb8dHo9VzlhZQX7af
47FSjrF6mzCSnwrDwD97UZ+5lVWtjzp6C9l5Crjvspxg+E70tfQJ2IJdzercfoMa
R1+19X/pj304nHsw6DzcZLoEScFi6nNMnDICS02aBb0V7pUd3BH7mYlwnSZhggNg
pCy1g16InuYsLJdZ/oq7rLHI94bae26z2XpwGzblDwGkq0BG45B9u+K0c6QWhyTk
YoLtiDVtTAtl5U5Wdd9pwX+Tfhz2W/mq4+qRMDxvcvWugq03cSV6lJj6p9yukuuD
6inG6NLd3MI7wZnKrz+rqk0mJLFX/Y6EORH8q/4vmAUt0+fWTHE6BMd/tj0N2w8/
1uMC8BS3FERoV5x4TPDmMmVu7v8J5b5L5iuFkzTu5oXSupktNv8M9F/UnUcuwzhK
180TrrPRsrKznTpUnVp7opfTpV+MmW/Q57UhT9x0PbY1X9HiRgF1wiG2W0boDYb2
KCunP4fTb8jpDa6U+wRjigyi0gn//qUbKRYYDpn2adjwJ3Ol1RJy3k9OffAhJxru
cLnaSu9XXRYAY+Bz/FDIP3hIfH+7LI1i+TxkNBKE4u/mPPghwgKi9HWQ3Fc8SA35
5Wv0prxYP2easd2wJDiUgp6Ae1IDl9L5DUCemNxUR07dH5XbcILm3LCPwiAXz0PD
obip9bnV2E+tbP6klfwxif7rqoUaCNp/ZZ5DkZfglMD+yaKWydJjCB52BF+FmY8T
951tR4r6QscKbf1w70sx0Rw1iT1PY0vOHgyd9TMSTBQItJ/tUkOb7KfVQqkrkPrH
jCZYZY+je6i5kinewVf0sUWhzgSDCStUVm+Fdy9nqD75WMt3qdsTlWJOfPTGSD2C
1fCpnFYHaoA9VH74HtzBg4IywvL6jt1N3iicU1p/y6/ym9bnhQoKbXTWMR51dDqE
oKwm0daGiciIyDzeYGB15sOh/zvnKZ9HrmT26LAPxCy1ZQ0sRqUoQP0swaoRiRgY
i0QweShmpuyXfogKNZ2ch1QlWO4aQMmGFT/XOMe2SDjPdKDZGYzTcaVZFlQ7lwWq
rowjzJhwPP7amPBHSI8EPeMvXcw3VVtbu/t/5tVb85ue0/uCvGvTFyjpkQ7xqfY1
5+u3NOb0PHEM/eG7XdLcr00VeOPzZvvXqp1Ufg1+mdM44/9po+9Dfjv38UOYXECF
WzIRp1X8ieuwPQKR9HLDQ4B3D5IThuaU/lKSdNv/UejusNBwrcrVF3rQxxj7xfYN
528P66HPflzsjMt6D0SiuUywFDogQi4tyYrjiYsMnh5mVhG4ieeaS1qrS9bdsV4h
wSLYnPQ4rgrAivNvMH5ZSvLCQSr1YgFlUgIqSrxbqkez0QRbDj789V40zbVxJlvx
AkMuE4dPYAwTAeEp9Z0J8MVgwCF/gnwUowqs2fuSCnIcj8c4e0QpHkmf/E6JOnDQ
ZAhfwUW28uVgv9GM1Tfu7Uk3m/DKOGLUa6VuvQlNJrsctRVxUtfsk7j7wsxXS6Mx
HBJlFjmOVcqvodxwGXdhPqreo10w65zo5prRdX0VxG4oFzXIUlgBBkQ9WuLYlVAb
2FhjoMRDgRYhIQIPWZ8zM2Wh2LyyaGH7VMI4e3jlOpZ8kCKcQjW0sNt7mymulU+g
kKiowL63PkfoouZ1BwZcy50cBlln1dC7Cp6ERiBZ0D9OTXHF4GXqhEAsca0siE/m
BLmUOlJqXaEgKizbqUFwTU3XAAqoRdtrrjlhHs0Ml/xny+FuvuO5hHMvlunP1X/f
ocWNYlW2obc4Hps5z8dx4Rpb4JiJt9hiVtJLl8JIBJ3MwopS4h8rask4X3LSub24
zigMairjnH0WGhQiSOho32vrFXwP6tEOYlpmEOTYFv3579vsvaz+hkjJ6iFQUAQo
HyYfRWCdCLe/yuwzDGH5GFEx4GvQOj1S6GNmOqQ0N44sYAi50+wMXae7u4IIKGK5
uYCGaSMZPtP0QoOrW8doUlPqfJgxUmSRjpxmj8+x7cLl+yFjiQE9rK1bFiafsrET
BUhorlc5Ou+hhcrHlPgoET0uy39hb8h3o08FKuJtUVEOJVULsV6olY16/E2euPOX
fwkRixJJ+8XTGiukGo+drq7sLxJHEW76huXZUZu4lXwLPxxkNGSw6NC5GHvnbWqP
vXiCmU1Lead1ARY3QPP4tyRg3rX3QD7KsIFOeUjsZv85isFvYZY++hqK9D3f4T9u
7eNQ5uCqazOB9IA5B0t0+tAl3raBlCSok4P4nkvChS3Ad8sogKwGU1vKEgfXnfeo
hbak0D31RlMyUqTb3quIbnkYIqxHxzVnDLArT3HYSLDnfWEVpgz8guqI66ejYVSP
wLS62aPPEyuuw7Adc9Tg4TCilv0im3npgqpyjqFRPiM/YhjiU6ccoBAI0BOKwbRM
YuYNwOkgtZZ2zP6a0BTdImkheITEN8kJn1sustXLb0SJddoICmd3K274NgL4Mxse
CqACNhoLCb+H+9jG20jXMnZc52fjDtvxPSxfyjJjhk9vD17w1cYlG5ghz+M1j72L
UQvbKOQrV4ui5ppiJOYZxMbM1++27pMrEBfshIsJ5lDyctXWI5N1vjektZQNxfeo
XqRpvWmGdspJ47s1Rl7bhDnKERFo7YLify5VDZVNeqc8M4t6slUf5yL7iYV+6f6Y
4cYdLzz1vplkfYJaRcNM1PyMLknrCeYodi4iqaIH7tk4c5QIpu4L//4zHu0Rc1rD
z4NnYXwaLTjDU7iH7U+fQ1VmXGdqc+FuFnxBheqcOyqnyqFJQAwCMEoTJjjQtsBy
x4twDm/17EvfMMvusH6fKIi8W4j1pmCvJdaqQsvC8PIDo85GBUM6OS0+daPT/OEG
MmwsgCFURW+o0XQV42ZpQWnUG0avKenPjwE40oWPvENZSv5ggkQVcEYfu2PIroDg
U2L9Jev6Xg7pu+TsHAH/y6Hqpe045PT1J0xVGt41VICGVSXgt8U2B3nQo10Uek+H
MM/cTlZnbXvHvgtqhX5ZvxB+y3nxPKLt/QxNcu3Igbfia505CqrfHBNR7y2BYXLe
LBtQkrLF9Dc90DFLnKSznPrKx4Wy+Kc99SOvstpMPnhwkUBLh2nxWrHHm7xTQo4V
9qgk5z6DIysbQtJGlpkihZ7rjuiyltRNLccy7wJH2Ad7TK3BSRJI3V3N0+CI7yNN
YgGDvEN8y/wTeVccSTTjdj+UokSv7t9cdI44RVZAA0DqeANFS1pecghwoAtSts7P
gEIoEvNHG4MnKLJZO9Y7znSuQ1+OiKDy66T4z2hYyuffsBTMaTdCBgBvZnj6tkqj
V6B69NtQ/0yRfHzNV/PTjslmOWZuTO6Zi6rmyKHt6l/6zieTWS6KSMOxJajuU5Ig
dQ8DyuW+Hk+1im60BdZEGqGwuCF9TK3ffnLETYuaCCJJWhmmcy06YPutbYnwhqtR
4N+nog204cqZpzvc6cR88LUY58d/a8NKTNB8ZZKrsDTgEpB2b9ORrgZv/ZJaSVj0
cB0/O7t7AZVKtN/PwFMRmOYrXkMV4lFfAoImegEjkrdiygjBeH4vxdyPLDGry9PU
jBPA87xllcDEYmW1dwJr/kGewsbgT2kY3yc/8EI5Bw2Rg6BvQmFwYMJ1souXmxSl
QS5PlS1Wqz2gVojpRyehLczLFHcoFRYKJaE5gjvaXOAg1p6k7pFRBAKZZ0NwJZL8
42oPHmUG72xqqgs6P/5/n5iMuBl8+DT4cnqbNhqrw08Zw47tDMpmbPyD+XRqf2a8
iXCnVs1N5hn5PLf0RkixPnaryE+L6bClqBgoJ5MSma3dqZs8E0Y+sUNp8hbmB741
wlW2YW3vrGDOQqIoI1FKNLEdKi0gywYx+57VBDwHk5gMKpuxdIdGMkT8ArDWs8xo
Imiut2QfsNhDCaQVuZLw/Qkpeg/SZ778NjfHNFNAAWRgHoEOgCXJw6Lm/Awyiy6y
7XkMK7jhOYqGynmh1fX5RrDYj47bL/1S1xoAUxTIxL8vVVjWIavgOF2EJBI+/FbV
rffgolzBVnJFi0YocZlOJRssT8EcIDNwlCWn5zMnGqjpW8mg0/IUdFLpikZqcn8+
5TyaEVxEp4FHotkcn+bn6OCjfyt9zQyWBiIbSQTWzMUFIPSns4cYWtQsN8XbnolI
9XC+D4Ie+zImda2+XSV4aixEgseH7zO8YVLGpu5TnA5kf3ijW6jwWkLv+IIHhZ5T
cXJHy7gRK1ytuHazU1UeDsspKZZ6ITw6dz+5F4StdNHS2qH0v7phmBCK3TbvYy5h
5l9JOExEzmk+AxzB5cYAM4sS6DvnTFO7WVvJx8MlCbNC5J2r7mSdcoHpyBjlsj1z
s1XHSNaQ77ODlRLB9ikWIv6xri6SJmcLA5UbCs7f5wZ13kpmSk8JCZzTlWFT0r3m
bTHCgU5GvXPUu55tDWpkxzCNEY577ZvzMJ9KBcZt7ETq3ofoA7JyL3wxGPjfGYnu
LR9Z/G+ZhEXWaSFBqaQ4c+QCt+7A6c4pZq8bQVG5vYwkFtEBKtuwNMBtgjI1+pVx
eJTuf34yH0OFay2b0RHF2sRSrJrgwJFqgkeO/rw3u068IsRQzl/CuSVG5pMkQ59S
SmVWc18fq/v62Qx7YmZe91ybtSngw4EcqC6/y+sYHHQwvA6mRppG39y8lJr2Xn8t
tbiXL0bsZN2iqFouL3taM/hldTxblgFAInZH5xGhVjY7hxsUTwCrouamuhdBtFjJ
6WgaOyBISO5ahrD+NKVm0kWrAxwXFnQJi6S9ofL7f55YQ+Gw420uP5QXdf1VfZ6x
uL3N5C8iQm0YGSjUtrN8KNhsKlDcL9j69Mp8utuKDgmWS3yGoAQRqEFzO96BJ5G7
PnbqT8GfyE66MOd1W8ddO7gmvbVu04kzJOSJLjLSAZvSV/KaaCCsGDbM1wVqDMFf
m4zD4Ue048K/AD0WJMDTU/0618TwxmpKshOvLX++7olvuUvNiR6G2Ju3dYzmP+Ba
8WplPr5eSZUKZi6XRJq5Dg/EkvlcFxtKWh268tobmLzYtdlnWzIid527zdgUvO4d
UDGfmxWtuZOPm/o4lRT+eNFddHaWO4sEojKxoHqJt71TP8i3LQIxtkRlxqtIIsmG
b6UiINNpGUZq8KEnot2zvhh9VDB+wI5pOFOrAxmK35hRczF5+csFuwv/W0i9Kfg+
bXoEcnBCrxTMCRz7IJowHVliTWFBCBq97tBGtC+tuWwFrdM676f3szzzqQ1aAZ++
t06SHcVJJttTckgqx3ZVvP5Ct66UiZyOuupz9oUMplOeR6px2Ejre2i/yaP5UJCY
SW5N9FmLqfISYdqZZqYGorWvqhHdCeSqHnVJe42s8gvnwd2uZ2hJ4wQFtxR2GpTu
5KnNaH+v2dIuB90vuPXC/st3NMSkqKCdvEN0UZzntVlZmzmaqgGVe2igg/Nv7hq6
+7DBJmvAtqNWQixbEqzk2Dz59ZfCdpVS1ohRZqO01OjXGSiUlKEGUW/uJyZfh0KT
UkXttcN4M5uoZsNuH0TIVKtKmVPqjO2zZsa85HZlx0085ZrTKy4CqnOF7+WjQ111
bCMwp4B0dJuIlWv/1v0xxbn2nqFj+bq2xJptnzFI0Jcf4jRIoWITpcGmrjK+RWyi
6AuZOpmsoh5yUfg9qdogZfARO3QgWxntSvuZFa5iDgPffkeySVHtHHA/O7298mwR
AdTX5R6G9ZQH7LFjUNIIPQiP0c+iWloiwG4mgxX2wD25EIWgo/7fDueialHwNi0U
kWXPCUzcLpe8nSyEArXC0sjuvwfzS28C+QOn07z9WJRlST/5K1w3OrTtUx5ybvOA
ecJkKNYql+7K/eyXu1HdnzfVdGNGxIvsh7dsAhJvmmOTP9trupJmsFt8FAKs9z8V
c9/0EV66zT+DBPgEySQMiodCK1u9vcrJDp+ff/6Bk3xhQqfputdeeExeHFCZ90/e
mU+Nzif4WEtrbc1X3Jc1lQiKXu6nECkRxAuYa0DrYW8J5xzC/HB0KTK87KggFGM2
CWgbMAyRSJ2r6Yh1eK8lIb+jTmdvD1BokK27KD8jE6mfXEQxPHf/LL3e3uPCOTYU
YSgKWVPejr0d3K3ZQw8Hu6jgCTvJu3tpR711YDXEGB4zxoHPWnSSHopHPoUD0sF5
XLa5zQqlMT9dS+hy6cWL6niFwvQHUuM/DEJT9grBWLNsiGykPezw3pxEJneb5T+P
E2P0dw7aB3vrwoZ8K9SzjwZF/Tx8/ZHewQJctsUOHQh1lI+K33kcyQFBM01uRzHf
NAYOCnOLnx3LXAn1mrJ1OprRnFfcWZCrJ6/k8SKiYEzcJ0j4W2fVSan0OJ5d/GhX
7d2thnlgTDP7wVYJkb57GCuEYqa2iOd+Bk8pzzEAVyP0bB8VsVkibipRIu9L0lA1
iJ+TdsYpEF9x8XxwlMcqADwjnfPv23M2lhmHKUDQe+Q9XIT0H2JTQ1qlwVmk3Tcc
HUv13JrMMRBxAKmX7UuNRrDab6OBcGrhe89I1Ls6/rf4zvmICmfT7WibVHR/de57
HQ7jJNl//pU4RvqxGUh4EEW83m3c3BDHBIP3i67wFrbWhzMc79wdrPIy13GXKg5a
L1K65hiDmILfF+jH2Pfh/HPTI3Wsuf+oqUZbbz1nYqJTrv6GtjBD3cd7kgXqMMqQ
woAuYi4RoFcW2jLDihcRSREfSrbp8Nc8TrGEtMAP/urND9ib6xuUjRPy9OVrTZ7l
edgLO8EdSP9raSIJmneA/97T+oNr2w7IPHhCW5x0HiboDBUfdC0ZSUaI//ooVtpk
bS0uHTfDvErVNnOXxGbit4BDv4Hmq0NpdsFWw0StMuu7otMDhn3P/0dpuaFA9nwX
Suc3LJdPfeOYRpbee2ny8qCNjWCENf7P2SWMiuxT7hIa+us/APYZCenKiCKByedB
iZOK0NqDX0v3AMSB68yA4/0u+NeV77lNqr+02LrZlPgPWKYzI1vkq+8uN+Dejnm1
wx5OXam7i08Au8K+aqtOS8ZwIdmM5CcEMirdXes04dcP+RWc3cBBySs179Qe/Xvz
zbe7H5k3quxO+rKLzxYO3svdi32Z95KkfdFgBpqqDC0dNeKiZX+XOMN2DVeg96+a
nGPUXBwuNSDoJmLsd4i4lb4Pkpw8J2aC0cajpxZs2y1BUNtpH6N5dB8bH5FDl7kv
XULXHGUmaoncHC6rBJJQ74sYsJEfE37fcaGx7XdyO6iJJDOHFLHipGxDDV4UC0CS
MAtxvFWBsNZ4bgpPkKP2J3iDYsBcQwD3l2GeePEnNTdTbJ3uuIcohrKhR03sy1Ue
XjKLKBWkk/N1thmNhjQIzWgatWbVtvz1WvaO1lwEujTbyftiWaCck2eSBtz5711s
dfT3tHjF6O1ZkVH1WFi43U4ygzrAPwhxdteO1PoqMbNBXOhPwtfoNPq9MuDNF7c0
WUITCfvZqvBRe/UP1tHgBsrHuy04NZNsrX0keA5fty9vo1r5iOvw6GgemhfU+FjE
p2v/vDA/YqUAzHjosx4d+CorS7q1XiXEQxDuoOIHYPx88eWoHuS1TviNtAX31GWy
CKwUXdGeOXTiSuA+vmxH6qcNTozbN3MI2bIJ+beaob9NjpvPBI/7a+BCyjPsTGxF
aMAdo8zVGU38LQ/VR7yTm4tR26D5UFPwggUuU3NB/r/dsl7K6Y6JMj7cQdiwO2aj
MX2Uxy1m1koQxFjBRcYO39sccy/kDotWip0sXTWXdsDJBQxbl8DU/n5vVGP3p97Z
2AKNijSU3Fh9xLl00tW+DEolKW8DqyfaNMYx4TEBOwXVo/e57Y9IWLt4YTaFDiNr
yqwWzO5qf+BnKm/FS3FJmYB159+UE/V536YTzNuIBzByaDtbMbkMxsBXmm6pGPia
CREirFnw/a67yfVn9NarDpkeogItbOlKAfl/aVfOeYyWOkItOW+YG9koQm0kMNFs
Tg+acivu0OO+SXHwYmcgbzDeH/wYF8cXCP5r0bD8TkfntSHoC5h7vCKBy9NkBDH8
MQLh8zngEqdDh263hUs4g0/VCYPcuCXbJSsCXPTO1n2hMRVpSrwr1RNhyKkmax/9
OB21vQch6trfSk5dnVRN4ON1teqeryZOCaWPxbNE8Vzzb/EBdciTggMnSrVpOyof
jj8OjLDsakHbc1c2mnUSJDhF7ooucX39mTHp1o3CwHuP2tohHKZ6fqicI/juxCWw
s7LlFXr6zUIk1uddmEeAUb8rd3E9zheM5wf54CQ09T/IjVPRZq6LvA7jHkxOT9If
0d/D7kAchAecITwndMjMG0hjCUpywflItMlJBr2rgA3iO6DEbq57lr5Ozf2ZW5WG
4scSlmkgrNsQcC3TLr7m4S60s5D0ZY1XAiC3BtdhJPCRBtGqJyNVbV92v0Pb0QBx
JKhfHUYwE3HF7wKs3191W3nD95SDLALZct/zhd8EZCa3qnaTZCFLwdoTT2CadpUj
Dh6m/jUmGJor6vPGwF85D5yMVL74cEIayxtjHm4rnxmj9AOfeRJrq8UGeBzLJhxX
Nn/56sm/Qjb2/K2O1zsf0D60khXrYkjY2ZjNnoLvsoMhC4W3/xqyTVzhu2z7yGlZ
YpvAAk/RLKoO55ZNTZtLWlRscR5QpR/sYxeXOKL2yJ5DKUptUeX8RZr7PDdtbKzU
giQoKniSGEdU+U9N8lVe4YDueUi/ut8Ss2w7+ZctSNbpSxB2Um6kZVvSIEVtY7Pl
IhyTRkuhF9Q5/yCSqIZzdCyzJEiXDhvFdP6H1uX5PtR2Rt6EFCLGFB6GkXuW4yyk
hnaE1IaUtdctfh91jbW0XU/RMoAwfi06Wn/Pk9tgwGi1YavSLZ3cbL0HMdfL5g5b
cnazOfZBMxSzZN+0hoDU5nl7X+hRJJRFrKY+Q8erTiNrhucOcD/Z5BouuOQTk9VR
GB7/RFJ6wMmmTWOASICadrilBxY+sxUPZCNZmm7kqtyAKGBrcnlqIRecfdQs815l
OnlGMMsQ0VropwECKO4fAAEPI4Uhc5mujcaas8Lnh+laosJ99SdyHxNu4PJIWhe3
imRZy+k4FeAUjepEDpUyYo/Ao0GGzJEBLuoAsy10Kx7eQpYzawmaaBR0AKKAps/h
6aUo1bnth71AbtPPwcorrK0aZnxxMigymP7YBhvdrIZL8E8rMmoo4eZ0mimQ6CJT
w1P4L1Ir/Ile7Jqni1KltigvYv7Jg/CyOf2uJ5VZa6Eqhm432Yv0kEwXbhKYLt/o
CLYb6LTjfeYveTJpMsI51CfFjQWzM5jFikaixEOC3YSIwKYQbGOVkri/VQT4OVph
swnAv2Uw1TcEy59/8NQNdfQYc6ppqFHnRvJtKAazrctfNW3kJXCO3TCXw7TvKVy5
fGzK9b8Y0DyxcbC7f/TlOCribzlIgKjQxXpFUA39XOktHkBcTm1MqVbMur7IQjKy
JVysqBxjbXcHG4fq8jG2ZWJQlhRxxddazfoVTr/B3Y95RmDqd06MwcmqSv33Fdvy
Nk/ogS4v+7A0EsLvQcmPGNujookjDItRgoq3u8NEXUuq+95nEacscJc/DRZJevJ+
cVnuv+6qsBJ1Ppe5sdDruwmKoKL7WpxiQiJY5W/ErGg4w7U3weLmDZ0CGZa46y+8
VZ2+WD/ycu/iw3Rnz7lhHaRS+s1CWOAUARNTrjayIhQaY2FE27dGGibFnbI8mEGU
ds55IyEZpQrQSGxVsp9nX8/WNLCdfi2lM/aNAg6sUw2v23fkcM7lUD55BRsIwHjK
EH0iSE+/a9Ap0nT1DPWxHiFilaiBUiGgRFiAPVvxX6W8+Bee7h+T/gEdwyzdAMUF
TlI6TqHqAsIUE2bSpojbwFmXZyjqplqPK6c1B/tMvw92EY7X7lIBFaZt7kkkw+vm
p6BKjV5WAjXToMkTX2bJ/9cg8WRTXvdZrTLc7r4Qd7IWJhXuH8IEZcgm+7t8EA5k
UBylB0v0wL5F6YEQCVGJigFAbvzWc/usRQaFLVLSJ+xv4pSvVG7Ns81v6A2ARIyF
oEt68xJu0ZOuWtT9pH0LEsLNWY40dKpHREKW6iJEgjLYkwTOsGLMIG3hSBETlQlP
4wfz0PqaMTPN8UDMIyLIFYVqB+AOD/AaBzQuru6tBaHxrQICDh7Migsds+PWNkFi
Pjd29YIlN5lHIVuO1qDcEwIY55ty7yk1x32XtSfm3YH9DmFETqQTGBnJeQtGxT0q
aI3jek7DyIakMK1gWxrMswe+x5tGgZ9M0oqZ9Nc8l6jbhBjn/vHR+vjS9C3a3A77
/ENwpakya5eOsbT3RcP7K7L0/VPkH1tNWe7KiI+A09iQZ+OaacaihOnnA1/xVX5d
h8UyRl4JmLHV+DZ+q+nnzbbyKBPJHLtwW5yVVwgHMqPjmNxkwuwaCup8ayOuK8Ug
rFhIQwLrUe4nE7p+UQfugX6tqOOKM5stIro0ObZ8yqb+8r8a1oJKpzC1F32WABKa
EI9EMLOVGx72R+05TDhsiP9f838hXOILEnmJapL4p7GQX648QqPBK0whtLfNbRes
jndhxrJzdYhQrCapEsywed15KA8KFEaD27B69oz4Dh86rChpiH6/PWGSRdBYsnPf
5woTvry3UWBOSh8Hx9NJx0OwX5Bu3n+S9TNREoBzbKp3FLMt8o8HSWK8kiiKvNla
V1hL+ZwuODSRNk8W2z8c6dDDxqdYcQcYXMEMRNNut0o01uUstG5T9Qq2kd1BvLjb
5QQoJEwNOvLkoFSAB02fT+hMp3W9RP7nustjAeHEhdqvGvsBxLkB+bphwVV/K68B
RTcXkw1PdOFPW8dPAJkFI4K0587A6mRJi1hubxPUYNNnv4OL8dcAjEQSozrmbamx
r4Brfi34KLKwcYJWOLUr0Gqj7kWdqb0kDMYkckf/4T8KEE4xP18T/wu/JJevw2yt
P1DNFMPtlo1YIvDreDtLjsp7sJwzf4Po9rRhVZs3PABhuBaPrlT8dHOq9G8BaKT/
sWFdpMIOPPs8xIGujvSKcIZAht44uRJqmWPGgm7CBHccVylvAmB/RKoElWnjElwb
EwioyHE3QmCvJeZV4C9Xl98nbHNHj79kv+XJ42AvbPi40r0GW1aynOK0fwXNl9m9
VmEefOajsLLo/S9reavVUTidduqwQBi03KFzMQzwcPrFagz5NdXWpwNCzY+3wk2s
xbO9csGgooLa3OEc6DLwbuBOW72a4IOcvW91V1NVJuRND9s6myglvab/tk+RPnCT
W1hNKZstCNNg8otYzoOMrGk3lqAhiZ779FKZtCXjTp8JMexpJvMs0SgVTk46FNQw
CpI/bnzlQxpCAw689jH3GnLuY8Kg76d+rTZkDG92sSUqXbTOmCci1i+VcDoJ2JGB
HUUoCzawy5LK19t1voWge97p5IYngj5Ow8Pe036J/Ce8pK/IPCr73XjqMYbjAaPL
y62e+NNmSSUUwgWnYcHk/7vakl8OU5l4RT97L/Zkg8ooVDf5ftRMVZ7WDd5HR0zZ
+eApkgQzYYbaKlp3XlVY73Or557+jb1hoxg9RIu4lQ9vdJu53LMdncLehewrCbKf
nyhaJzl/VNv1OB0QkxURpSPl/ZDPQwuBsxMTL40a146rqoVptn0zrqNHnLdJeYPb
DmNKpI5FAiZLzVQwbx9qFltzCTO7nYIPjyU9wo0LcbtjMzLSKiwcO3iLL8iU5ujY
l84hnXP5Mlb5NGuN6lklKVbKbsma5nOYua9BEbo5ZiAKIGhLelLwbhJravdhSBip
X/f9e5HR5dm4+JU8EwtGyh6jDhfXqduAiKNDOzIZHuf14M2xmiH40QKpbMxKvRlw
nD8KTQNZ7NPkVKkKT92XBrGxsnA3LBnwkkqgoZPJ+nMkbyoxHPM4gK+zdWzypC+1
tS/4H+aENkxogViepIenINbyRyGQ3uC/gLVax+IH61+XV949v/q4VNL250rarA/F
uHI3SUEA10nj3vaoE1JkxTTAszSPXeIesh4S6WUNdoP0IOJJ/xLokzDKHUabDafV
fWJA34Ags3BA3n2rzn3HSb1jaesF8LdOHT3HgfsaT9Udqep/2YecK0PW+8SqoxOm
t7YCMIlqPC0SWlHnYSq/ZFrZTrV6hhWq+db0/I0e2SNUnBrkZcOYoFiUUZq8QN45
FdXwukCG52BhcMYQjHcaSbxcJeuELTbcwIY/IDS6Xjs7AY8IVFVj5P9FBk7jj1cV
w5kqV3dtK5T/NdOuRo8Z6lLcXCptK49FjF7JhB/XDwhMjq0cl4cpXPrIOP6n8Tvd
rYvIDiI4y99J79gOXV9wYlmmFW98q6VwFYu6Bo13u00enyOn/xKpF5ptH+mLbZ2O
Xng8y9Jer6BSbWMU9MMOibrOfyQSikd6T2E5k2A6Y4oIbKdt55p6F23rS7P1JpNH
zFNsO+QTcB5xwurKY/2j5DbgFDPLS8g6s9HZIhkl/yLXmkVYkTLDyRzkcztq8qZ6
mO6CmBO1cqRlW+TaHqO/W32gd4LQSbgF0VCIjI8OHniHvyy432MRpt2JLdvaB55m
09Z0uH2ggCFb/2lO1A5h5aTTub6aupXVoFcr4AsvwbFsWwTB2PdfVusmqJJhUpZt
0PQYt2B40ZTlwzjCq/4kQ7eKtRUAEE4mMKWIC6SEs84EEohmwnSDDBvo4gJsQ/xS
Y92zYJuXfgejkHGp4HUqodNo4Nshn060ZPHAxfXEPkxFjZO9QHMEafLjayA1XCZ0
EAyG+5gvk/z5N0LV/PAGMsNqoeJUDbRNXUAl1hth4nxw5Qam/H+KFXMS2FwqyLdq
huZrHykl9iMt6YMUtsvFftbWwMxCNBBovaqgpdmnDbkNpTPRmMPH2PP0jNyJqtoH
UkS0l2BfftBgzEk8iMcdwUC82Oa1l2WtVYEUyb4WaPguev0jVO3CIEz2RpgtO8pX
R808ilthF2OlT5E+Ycwyc9YGzyLlq9UzQ4zcwVIB/A/BiJu2G4NQTnDjaqABkI1w
ypYPfzJmUE95nFnNoHRSQ6DVSGk0Uv8ESzwTF3mcXhGpYqXktNLjx29xRtNvfEYJ
ybXL6aBsEqXeio88a8nlokdyUH1PTuSMNvwq7cLOyZLtyk7b5sVdr2ZTpNIkaBbP
PPR2Hbf3JWwO0tHsnj8vFAkWeGTfqA7+Cl426PY7til/hHcNKb/m7lhYihxkYSVa
oFGI+rOPc6tBBwoA5zdyklVT2reQcQebJGYLAIYH/nipzrtQFKIjpzNYr9jOHU6M
8wT/5rBVDbCFLhT83GtwAV5JBbD5gVxtP6yvzBa1gfEk4et45rhv57n0DZOyNXXJ
zoeNWBQE1D7EMIOUiQnkxWz26chV5c12mBXX5Hp/KSWWShgybBQuCkY76D3bvRnB
UvIdj2/r2n/q2ydEa4jY/GoIh5ZzbeqMucn+/O2CaDKK914L4bniK4xjenuYoIlF
6eKC6UbQ62eVFX0dyIFx5IumJy6XGVlI/ghuvZGoxvyNQijN1Og6B1QhrOHZcmxA
kk5GYZMxjVEK1hpTZi4Vex8+kdH6Dg60P3YPhL4F0PLF/hjoy0NV8aoXWov2Sv+k
rvSFIGoCclyhDfz2xR00xVw/cxvE0IZnEhaL/Q3hrsutysige4nTVQjgIyr1sgNZ
6egOf2h6KGxnu/VE4ioKYWZ17Y3GIEP6uRWu4BFJYwvoTh5gCKuvNQ1wQ4HNeL7g
UGDU0Fgrf0VcKv7SSvyTp7cPnGZNonF/LfHU1Ai2UJINdHCge5w4NIKLtjlaUdu9
ZswFy6DawNVrqDO7LbouIjy1Sr7H5i1NLHghNdExLl5TORlEWJYInmbFNnbyEu2i
Tt5C9f0GGLR+I/oAG+3X6jZVm71UR0M5gRryIRVrnZA37p5OpxwpmthWYZL780Hc
cO2ijmSrCSftlJcq+6TqaWRzRnnP0Je5xfYDAEJvtigxoeDpezktDNGbCINjwzLC
zm980iyqvDRX908xm6eRxK++Ry1OVpZiNfOKQ75ThlXXhaH04AHD/A7vYDcQ87fE
wIkhAW+Ff1n+GUklPKC8g9X17ddkE9taYH21lpIyoMWnqr2gPZUD3UGwgWU6axrh
A8mB6Ukg8ZhlTc6SjOP+P0F4s5WCYt2dPbQLzOBvNI2D9uVsrRzH0Unv2SakupCB
9fQGnS78jCmOyF1x0MjvwUDFoAEL7VCzN/rc6U8dEHpQjzV6LTzeoW5FnEPh+YjB
5Zp6Ck+Zq42xGTaRDH+E6bOFIi5oTI6py4NN7QY7IUKNUyV4gwAm+9XNpsHJiKB2
BkppyZqU4OfWQ2ecM8VELMZsyog44Lhg34wMWXjuZLuB8/ljwhfmLq56wuYReh9K
rJAMsttISAk8qqymTcPgLwzJ0cupV7XFug+KDKGX+cPhnc1lPO1yb5Kpd/mI/GLW
kzgp4JrEW9wD8cN7sS8yA5xfRDCV0LvvElD1rX2o8V5PwPMvdwl8GuHtr+cbKVVm
QOk5+MG3Atd0FishoscglzohkBrMr91EdVoe+c4xn9S6qaFTgkNPJAb43HELNZdT
WBTg93zzzo5EYBPkgo3AxyZI/7QeFPHdUqbwquzMmfhH9nvu2HORliHe/gffpJ1W
yeIanKc5NgNxNWH5byVtw8vXisjDWAQX6pcTGCq97fvp8AAAaHdguUWzj+evdG8h
kujSr7n0bVyRFH2SEl/tG2JC5GeBi2+DlpGThz6oyQ24uJZ7qYw/tr1vDjAZ4c+G
yVxFijTOVh9W356GVHkJW876FtDmqLwvqghnxpqZ8KWbPf+33iU6AaFvtpYWeJxd
WqDCnDu/qBtD0Epxh3bkZrTHKsqkKiUK2gF0IE8vr5coTGkf9dqrqpveNOVsvsgt
QFX6o7tnEifQaucp9a9bDZCjEpx7P8Mwr5JhA/yvmCuGHCSsB2DM6RBQJYTUm28T
KwRgfGkHu0Wvcolo80veo5Uh6ahQNR7FElfydTr86aKLl8f8WhDduSf0NpUFd0hD
n4AxEZNMmt31ksoQIGFOMlx5eAxP2vB5OOcpRsTNQD1ehdA/c63f/+JmLguaxoOi
6hjkmJwhL4L0fpcn4LxgkRbL3uY0htFSSRfcjn2FJBaIemZRRXkd8wysEqnPl0Nn
EaHOcr6vUxZIOaI6LkqRUs+HWosNfezZch8dNVZTmWQP1dRXy2KnBnArB1Wy52gi
PKm8b8O0gAlPsFXU1MSkPJ9KcYFWnQd6AaZY+XcRKs4d+SXGk2iU5CERnAELrwCY
MnF55mFaG0s39llqOoVB09bq99kov4CWVcy1jZUPACpoUR5OxjOvQtj0CbeOKBtS
mWS5yPiNnxYrZfFHtlbVCZmEv73qIDnJLBkLd65V1wTKQfMmZ+BghMNzsnnOViYV
JIuLMgcl9a1w4tMn+75wFlbGxCeSyjalVYMQXcvZuKi02uN3O8AIRupBcTAW5ZDJ
fndbCGcalCQq8KnRhLuhUChgzi3xqBzmFkcoASHMq17dHbMFfNzl5HjJR6oKr7fh
V8/Fn950WGhmvhdBBi+0AoQ1a8v44wG3mtx1Zci4BJUP/AHe3c2CiP/J+Lg1882t
RZKN+xZTWQOPD53unxkOPyie1bs/135hmderJWO2cDEJFX9QCW+1dHx6l+suYSkO
B11AzLAx/ePc+4paKdKOZFsqzqjSR5XgtCeKUF1DG+nEApA16OQvaYiNz1rvEJDr
U3KlyewWa/UGOeHC5B18BRrxBBgESxY4muEUAifSKVgOHBjsj6Wkouv3uDvNODnx
SQhPXIWxXK6rRZFkXpHchkydws4b8JPLJL2UypUZnyArnPZgiVLMK7nRR9vaD3S+
8FeYElT2jkSOLBJO8aRJut0m2awGuCDlEkupBKHK4CAtwJVBljbxBt0FMLFUpj/Z
1U/m0FBBg0dSLFKf7X7WzhtrbPGIuYsnJTCcKW0zcbuRJR9hE5ZzLpeOsXCbLhEg
DfgwKgNUooe3Pq9MyJMY2yhf9NJEeSb3pl8r6Ng5lc6NNJpKykctogOleU62rd/9
kKaFG/EzeBcDT1EGldjozGHdPOmD9EBXRUJiV9Llmd/7OzihQY79uWBI1mE8/BtI
6Igbi8e6TS+aqvdud7qBVaKiiBjw1c7wtyUJ3jYKwPq6yoJznFZrk9+Nbxth3Hzn
8djvdAN1BDACb7fIgrujaHQ/00uM/lr43JaLGuh5kp4xYsyHxBI7AjBi/JL7R4RF
C0VgU286XOrX0I/QOiys3KFUKUrAlrn2dIfNF0zXZF7ctuQTxGYopplQ6mpJHNgJ
/L1Ew42Ej628yNNQWqTA/qNZKgcqzx1v7JuxCmD3EnWgjmx8nlW/gcZuaPqTqdnh
CZp5g/CEcPA+hUlFmwMQ8caQ5cXYo67aT59B0pPNSB6T6U0HlSreEal+xQ/Nkutr
yeH56YY7p+XN0YY9DSrY6OXW4vHUPCk77l9uuP8HMtLIEGiAvl6+UBgLl+cPJCUI
AQ+LDvo7nK4tSZcIXOO8GW3UkjdhPmVZT5g79rn0foODc+i1qlgCZoe+QJ8Z9Gmv
zD7EFpeH984pF7Cesv+KIGcuYallli1sq63KbuKZ5Y0qJU9QqElUaUADYXV+jJE1
Aaq8NeZ+RAYLQYDe0PvhFHjQp6JBlijJ8YBJsJi3TxmEwOgAVrxl+45RG4APV8us
1lva77CIJkk9asZZu5SRW3IqKQl8oO5N49+2wA2BewKcIWq6QJ7vqrHkATnjRJzL
QGxzL4xrrVyPhnamlMN1Pk4xBYK1Du6fjQBBKiImPdMXyuWQn09MmLCLkneoup+N
yIPz5lLDlnA5j7BDdk/lZYKFalVkoe7dW17Sq64eGFtocu8TW6AGtJBWr6DnO/dj
zTgdjveR8wvIRoQvOPWz3sisILaxZFygCIIlQdhoytLTleMDcLHamLI+YRXQRY3q
/N1gPj31s7jFfPsacP6gvbzBQWhE9W9I8SS0wHU32qW3oXbe+IEn69fPXilImuXR
PP2ksQBj1da7HJsgS9UYJiS10cofVWYg+hEi1/a/kR/k4XPRsDa3kXyktwPKuodc
1QLnscTfwV6Z+Ve4xWwjQX73m+1fABZizq64s50XnBuIhS0PmQziuAiD/vfNo5jC
vArAplYNiLFRXUiewMAIbMyThT1c+20ubglr9Rf77jMu25ek8izJXQQ13z2vnX1r
9Eacpc9Or860kda9C8RlciKAzbvDxrPipgD4SsnzvN9LYrDGY9zOeOxXOmmrPzFF
Ri9H7i7T+CqXga7S7CBLRQdU1yWVrxTf8VFN/ffo3idqccXMX73YvCd4lwse1VcC
7OeVjZbmdSFBPDosQhLYRwQaMLoVBmy5/4WD/5+U1B5VNlyVTqerVzM3Pdnd5JGz
KsA48Sgi+gz2qDLM5DmOyd3PSlPLelBaiGYVlCVzTuAMdgrK7q+ajG6XL9Vmv6ID
DgT79p3N9pXrEgbYPo4ZXw0kZRVrA7NjiffRSUdFjwczq6xrnYPMmiJmd77zw007
19q0YEG6MXfI4wp6G3eC8lo68ahz4Mh/hMe2QVdR7n08Kx86y0dv4U9T7pAkD2gM
N8w+zGWRTm8H4NULcCJ4RN0es+LxLvW/Bykcxp36gRpbO1Ijps2OgxMLHA9BkleA
OfXcujj///TSjU+fJoEB7W0FUe5Zkr5y8X6R42LWQORixvL7UDuoz1xqEM51gc3c
4OTvlR5rigVHJ/kaFp0YVOJtXY1UzczhqaUGABLBugZyAbRY/dooXyF4pqB8tWpy
lR9+e6SXdQyJb2jf8p8N5c2FU2Y5ssE2KviiSD/yQbKQx0/YKPkiHMFoq+dEKVkB
54pv2ZPvRGxIFPL0QK4qcyviSAX4u9379a+9mENnRA9889kQwyQf924w7HtLXxcp
O/rookXuuwQXTyfD2czGKCHEf2MeXSVlv/bAq2YdkgWqcHtMFfjnertczgQMxgPH
KsSa9Gx0+cXOhyws/L4xOKnlAeOPKEDmFT72IX3Ik63M76yEHT9iApLZVXdTAqrx
X4VRltTv9pcNUdkmq14gFqktEOLfuBXnt7XysAgzZ5Mk6/2oMyDn8QC7wQ1GsNA2
uBKFDpqQ7zYJ8gVK3YqYpNFUwkOg3+MW/B6E6oKLSX9OS9BL4wCy5x1l5G8mq1Cf
XK7humSvyzCtoblzqzKN9tusgm6ZYcvWb2KtxW5S0rUQfLZIl90Jhv8cOisdyFro
wSiRjf7OgGfyXeutwSNBjUQIGImHJqN2k4Ja0+5hhLeS+eN5l/xrUa1tI66dYTQ3
z53jXtNYjcr2g3nv7kMGsfD0tvj+Uf5khfZVZCTIISnchelnBVqSWreeaWPPfdvN
tAFpLJ2kwwo4okRZB5Yw0VpPM07lLMG/xUuYh/ojO0z3+kFRuifUschT3uGB3Vqp
Ww0/tlt9KDN5UrpGOQiLmR9pLXgXafA2FdTEYjQgN/7JyH92Okv8uteNVK2sXKUT
usZ/VgQ98Z5r/mLW6ylSYg+iwWwsmeOWzfaTUdb5YouPUdow2XvMbUMqbtadPKp3
zZyhveYUdYY3ibJV8jAM4F0qBnLcZDv8i+vbstBVbJoiGrQIPMKHO1BxHvutb6qc
j27SahTCyetdu98aeNGEe0uDbI1jiYjgjfXFGW1+ZlR6BWLhQ8hcoT11wgEybrpP
LzIVP0ok1T8pauIERGLQjk9q8bF+aDNgf4fi4BT+9BR49iGzr/ypYkDQ01FxR89o
rcmFYTaB3pFozWdVxNvSZUOZ8FlW6mHXIF+/TT7Yd8U5g5v9HputRkOtEgrCYxR7
eiFwnBspUNu+dTOE7VX8nxK6qOasK4paRQ/896ypbkJRPe7k61y43UfTJBU0Qywu
VxTK0cjMOB2JmVrqamsBLyoELPL/PGd/YV7XUoVaIKEYZJs4nmCOCqaDOBbpXAjo
jaeShcYKmNXl15MF1AfO12ZdJOx5WpowP8flZyXRURIPrwQfCH7gbd61nH2D5i0v
YyDfnxbjlFQl7CsKPCVKlmLp0BZ/tR+kWpiPagXdw1dt9FfAQmROn/aoA+df2Ola
29SxtXqNz7SNpAnKXbtD9ISzrBx5dL4bZHbv6T8ImcqkTk1tAPZZgpLSH7kGBTLn
wX9dF3vSKFbrLmPqmiG/mO0nq9RLGA0jVXI6N1s1OK5Mh6/tb+AywuijUwOli9mF
ufzM3IBlxYd66UXHlBkaPYnHo5WHSDeCYF1L8MGLS86kD7Et+OArdhDltJTF2quv
nV06HL/U74JFjVZlN5m26GFKW70YTCj2FNrliCnh8EA3bWO6MP9+SjgmgYcQKpJP
44ye4IxcfWepFrWEJ5zxb2atCQTJmLOHqbuvJ12NyQ8A9vEuCKleVVb9W7rtibqm
Z9xZP+cbGYd1mkfLHsu2FKVKRldiukO6pxideo0AA821XslU14jECRh+WSONR2o/
HqgpIbmcMjJJ8shReSZ7pBvAC6GeV6HF9ma+mgMkO+K03gqGwVoPX9iv0Tcr9JY9
7XejztRZ9AHrsQ/ZaR/m9AYq3H70K/NuRTNnBN1zTps1JbcmmCwyHpoG8ameB+Hv
uIaF9qArXljK1N/xi9zuJJJYkh6Mi4H5ZKm+XnULU9RMQxgH67aT2YtG/ppbxbFJ
rz3rJenpPoLu2AmSSF6yg4rXh1tMGlbe8WocP7OPwuwBxnHvuCrJ7oDuWbEfEnc+
ca8gc+4Zf5Gw8GV5pfqQrugfC76URIYxHPqmj9bs0pX+XyD7ui4CRJ7Mf05FdDo3
loy/fx5llNuBhkaX+3fsXMI45KHubvqCQcggA1Vu/STt2lQI7HrmCZZCuPtioWSS
fErIHQr8rR3sTZ07RA8e3bXJadwwD+segbnvAh1mWOck6ZyCqSYVQDpg6tqdiCsG
9dX38aqmvw03P9k10z685kjshFVr+kuO6LUTT5IMTwngQN1U70z7DJMHUSU6R6nh
Dtb0yKodTWRExOH/QZf087JUU86qnSKAX4OV8cxqHDEf+ByE9qC77avKrMPPT+6S
9KWWPxR/5PNqorueibQ+kwSLqOC5cio7i/tgzvlgXofOKohpXbFDCUfXVgkCK8Z6
QsdQBSQCi4tpEmTS1GAO0zSp/dhbVof7ROWxmdDm8UD9xC2VD1NNf456isqQ0VEH
5/Q98xJM3ZIX1g2jIErFWGzbHM6QZ4VZlIiD3TFfkXtvWG7zDwKfL71rCqV6NHIb
e4w6HmvXpTnFNoUiZ2cI2rEemRc4dDigWDgn9Jvg7Ve94s81ccpQ4XjnbklOO1k0
fFmEse+Sl6rjEnK8O8kAyNmkivXTyozra6D/vjml4fpCXbFJQ9scr8v1zVgEZzRQ
7JCmN+9PdrPZ9XqZ+fa6rGn+DOkwEnARwus88kAK3onfcyHO5NOJZKGJ3TdUYtSP
RmGDWLcvw3h5eh1Ji7csRLFgr/gMVIv2x5j7UlpUKCe7I0dODQUYt8uI/02kJDnk
AIuXIyjajyWKPMTeVhRmL33M6IIli5UDI+vLVPUD4m91mOUTtyi+2CsgKgBf84iG
mXbdIEDeZzi/m8wBTfNQo89qbfKVKwCPRMc/1pGt4B7Y9AKhn0Qdn3Is8uosGL2e
gL7QmGruZcxH5MM44VTmDh0VTVqCb7EQvXny1PBcxgvpGINwAUFveUOsIvRO+5V/
8i/MLbWjb+RsWjl3GwIpWYUaiD0Pdx/9XgReY4l6/Oic0G6RRgrg9RsWw2N8BACm
CJ8LPIwBoptqvc4uMCdQSO4CwrqY/Lf0ylqpIA3DV1uN+Mkc5C/UlKddKDkFQO87
smgp6MQWzMxpE45qcGC74pJaQNu+53UU8ueLDNvbPI//Z7BEXKNsrnVzcbciMTIK
A07dusIqpq+WLtdAZ3dXzSXRqSEg6JLbtn7EANYfc2XC4wQDMptkxi5sXzhU4Gyq
klKNSiGJeekPgXrlaYOdRP33uFMTbkpdK9HwtMuqqQJViwnM/liJKlPiEemLe8Fi
j+G7bLx7R80ZeF65jdJwCDG1MYlbOIIUSvsKUW2ZIfQ+RR0g/eyVkF6iFJbPGBg4
F3Q5AgG9gRvBofOINxmsuhYfK5f5xV2xlev/ahDyZ5/LgFVxaCIFRqnDwNBqJFcD
HWZl+TpLcAINgzHht0xYZnua47JNzVU7XkCCpqoQ5e2omqcAzi2fwmGq1/+TOuLa
/7+1VGSW5FeXwneM77Q2R4t0HKOMsG7fefcVDynxhF2EcAIP/67GWLxqbRJCC5J0
QMPMzsfTEucXMlS8rbzwMYoCs3bGqHVurxfVkEGU9tdUfSVPp+woSq9nApmPku/5
C6A7ETA8MlFnmtIvAEquvQ6N/AWzw3pRevwAMfpNbKbbZrpPJfQYcApEzNM9VuQs
yjqQyY/7SymMqLXX5tKXAnzMz6QSH/bLU41YEBb2BFbJY+nmOgFg/VIXoaOXFl93
VredMEdhvFCkbELbcEadYdJ5gm1Yj6lVcenuBU74D8/ZBhmxut2L+E1uuGMqXnOn
tBa8HuGXl4WwEv1Qys1VfGduOPf3ES26yitZ+GR6qt4V0GHudtJ+tijfWjYJGepN
X+bMasWIdcaAE0lyx8DlclDchPvXScpHINpqvhXklATdUp+bN5HGnH/u3aLanFTn
abY5+GdXsd59999GfrLEf0Ey+vUYE5HaaO5wTIv9RBTyaHyoLzer6oPIvLIEu8Em
HZXHUvK8Zwkt8rZlYWWFNKDAl1X6Ltr3C6lXsjttsAGI8IiaW2mCzBgconbRc08F
Ci02XgrGIKJAPWFHZGLchcpRf2I8xlkt+UqCSxebvbDCbg0iPGIK7JpUcndunVRI
8P6Qin/IwvTQYG8kux9gBBcv1q9M37VhDb5O4M1hwDZxWcIS3MY8pjRIqIhY8FZK
d09qEYV5Vj74QowT+PQcHct/ZtZzwYuUlizQcCIcaDYIZ4N7eRMrVh5wkPxLlGNb
QFZR4e2xU7McG+i2tgZwz2S+yzVZDrpxvxaoL4rtNePf1VGOUlDraBcKer7R8CTf
Qff52UqARx7CKsrAizMQbvm0KL0Ao0rxCJWDmjAGukohS0cN8E4pwnlUIhAaJcLO
TdbckXhcUY+Szdkar7COdzus82aDnieYpKXFXicwHg9EqYlyvTdJMHZZFFfQt8i0
OpAtg/mSBMQTkc+9xWgXLxM4Qnry+oqq0h4Dq4eShl11nLqIrqIrzNKpP1v2P31t
A5RPpoHQKedPoWoFlrKpwSygX+FFny5zilGMnZya+CWyCtFbgluxnP/vMOcb41yK
d0oHbg0G/JpXArLgYr3GKej65OfyZkKzKA7OswtaTuPZeU0JF+Hi8/PXYK8oLZH2
z7w4cDKzewsQoPX5LIYBSRORYafP8Z+vw0eaTt/HH0PM5dvmXjJipnmqYtwRySrY
0lq00eHGbMBNesQKz6gN6VNelKKAjCNnyRjfj6p0I7Twu5VNuIe/bo0CB7b3GDxR
najZy15CE9boFLGUhrWKmnK7LeA5Wet/9AcWoX/qNquDpXrb7nMVK4tpJWfbune9
xpuUIllLGbcG/lfmTPEAjleAvaZlDavYEmROmJWIgam5biDL+O2X8Ehne1YAD0zq
b6xXPC0VbNzkyIdLiUpl934hoEWzGndlhVOUsgmiUX59w8yJVuFdTGYfJErkTUT/
9iL0DiFLI0cUIgHjxu4bk6u/pyrD0vbZJIdnujO69Gpefi2ThDtq4YmD789R4PsN
THzthIq6RukY2bzX+6a1/HdvUuIKpLK1V6gpiImSZWDEroSRbpIKDqlwaQcIzlpz
xpM+T65gcI6SqWmelETH2iJSN7OZTmRHvJjpcpg1ngHFz2Y152lCLU2vGrIvQPE+
ea2SCljj4T2/J8X0ExRBat9rUfLuslpLi8YkbW1eK/vxP4blQzUCsiBxLXmfJCmk
cCoM2KHMszahQqWT5PF5jkid8b4ga/0EvHJioSVMEsZ8+uzja5MNaFasd6SJwLjf
IY/GqOpQYwDN++icMz4fPFmdKpFmvNZapPnR15Tlf7UkZddlCY3OGcfIc+ouHkkG
8vsTwzZGvliCUt9AqwAZo5MQ/xtAdJuRXSln9dWmrFes2n6G/ML5pr1NezhYi3GU
uRdNzfbVdZizBuxl81Cs+SBKicxsKMYY4OZJp7aj/GBrygtPp3bY1Hrm6ij7CHAl
ZPbThbju3iQzwImoTniUVZ44doktmJ2SVE3Vn7VsEBNPNEOkbtItxoO0RuV+Mfoe
cabm/vU37uFvR47ZHu8JXjqn5WSYvyuBz1dHyRv36UDuSsC4CCQ2njuCBbHlxjos
aCzrCB/Xsv/G8GCE6lf3dx6F/qQ2SQSMDqHoMn8K05SMzo5A/zAmh88UWlUHUz6C
/z8g1cwOjdLp3frNv34clA67OBNCR6qzrV+bg7KCxyGOOhpz7QRSkZecYYn9nDOF
KFH/obYS18inI89cHDYwEWkJVwgTI2CmvXHIZPs5FPhtCE0rJt81Z9tuRpQgwG7o
QD5ILvYG1N+ndm/oGry3tY6hLzZO//ufE3DiVVKFCfOyBiw+JMnKFBDq1TMyhNk1
6me+eNxWkuWyMsOxPc52paBB/124XrriFBxUz6AjkYuIMV4QnCiUC7GqNFI6NkWC
NXsAddnoeP48Ra2vab7Z1UlDx8MVKrlAKbLnWHK2i5V9+Lf1Xck3QFDfWYNUx9+W
MqwNOhnPcvC4xpffi+bUBCwvlsFt/NzG7hssqUXJJ32mN7HIrvWnVt/ArxDOf/jD
wIDrd42F9gONcGeLWUw2J0Wu552swtx4Vcfg6NhG+tTz4v019H9a53DRPn+tJtn9
qesE4deY/ZLFwBiezrswGNfifonM25kULt3VE13oKbGYIOdP3vZ4YDKtuJMV3iF9
VR8gi1INMIRtY+5coqzrVRWs7xrivpSFK41gd8QCy3LNXtOyOz3wPFRv6IvZGo+C
mNvJZDkM7XZkVmsqwlvqgp8mOVUiapdcyT7QsWMq72HIGhY1cAsUnK0uHjUrLagK
U1mKOc2FBBS9fDspXRe4G8LD/7lAHc3L8OXFQoOpQnDX+I7ChWn+fvDyGJF5ew1q
PXQfQoYLufBWCk1/iBGhnY+1BRDCfnEzTxTO4iDZFkPDpG5vW0k9UdC6JIMedlpx
flrwCKEtDEN25lNvRB6sTEBuWZtRaDWi6NUMvv/NlzPqssbWZXBJ8UJ+Uo4uSs2I
eIeaAwXhtZVjqUDp59Xx58E1dR6UpMQpTuJFrqgu9Hhg8fY7MraAukMsXPRwj/AR
QXhIMJxkbqWuEC6586o8QHRoEU6WteqSyUc9vUCtRnfTS30CCuJDg71LsnQ7EIcv
cLlvv4dPT1vHfciw0QoUKXyypbOoet+rR77tJrwie4cCoFfX5b9ZoNUYAe0mIPC0
f3NQftkh0esc6QiramL718lVMfZWfmEdJnq3kI0ZE8mXA78nSKGg16jvaC5JWODO
GCPFfnCBGnUKlv4AvhiL0puvrnTsFMfl43GFpYrZWPTcvMi7SvgrbVR6uLGjHzSa
ljssc6PPsaLmf8NhItKT4hvf8SdzatWvUIndG5cVgKrw+WVuHU9J0/Dp07+/7PKM
2K57VJqLoh0AcHTV2hoDWrMvdOUgvlSEXDb2yxBtFqEsTlE25CiheDbUNINYnVhk
Lw/AS0eXJNPrDQEKaUDBx4vfUC8A/cmqOzX/8NQuZPv+MqwNJ7mIbl7SXMyLa1f4
QJRRSH6jI/Dm74Pgg4yDVumm806dOpYGlLkwFSIHdwqT+X1p4ShOIPXE77Jhuxjl
LMyy/AFOuja/cYrJwjeSq813lFYyYHAZjzd/FCWjKvDF6hzdJrDkmz7D30SsBc/H
maty0KdJSfSiiCEnUaXMI26EC/GxRDXAYEJ326X30E2Ye4h8/WPuhjkLucrUNObT
DXmqJlsrw9o7RzxbFTSXCENwMTd8TskvbfWYDvJIFdYu95xffGKKvWlRePDkmFcp
+rSqAnfWjcsmP86R4Ko+WAOF1MomZDbw5G16KhUwUOWtJoEj8t0uiYMYHdTHbeFv
zOnBv7dt6c2uMHoCgYtgYdA42MHJ5ZAtekqg/3ZbL9BhCjKLkpeP1BeJgqvH+xN8
7F0UFqYSUANv+zOT3If1Q7ovLgFg15pwz3OOkgCi60hlftx9DbENu7IUX2FvhstO
G4DpGcPIRbKOjAoy2UxEIZvbv3s8981Qf7vzd6AUeL1EKhHt1DJ3bx7zux4eL+XB
Io7SaYtvlQEZaGUOgQ8PL7dkoaWSQpPZsRsXLyKh+PAxw/a751R6c7+FX7+uHcuz
AOirlqBBNEnNHCXTUzWAP+SjSiCwfpOEIazwus8sLCgr0mNtg7m+hdgnAMkE0OPt
08ainDYwfa1fO7P1TXGX5bx+KjgQnTAGtKC0w8wMpFYVWTed8LRgXeLZhjtq04hC
liFDihOjj6uI+yJzgjAwSs4+ShlczP+8OEzfvC+PjqQEKbwtexPdIeVIvV/tFn+E
uwzQIla1vyygckTfBdS0cCWky4MxiFCgZT4eZhLJFXdsvAUqZNKpzxgvf8cT3TN7
vgId8jehnqkh6zEd7ugSKKgyRjJXrAIYf4Y1yUf7wa4wv1z5UjBnbmZcaeqZY2cQ
9FLR2RvGn//Ia4ty7JfLJtaqJhqvDFQlcGnSQy1MNNgFtoZWlSpCO7IoEUBo6PV4
fCeVpwD3356rhnYtHS2icNlI8853f+jQ39FrVzhIoeJo32MTWc2MG9Ka1JsvmB+N
yDd2zAvgBoSHJQmNLGcTkc2Vp2ATndnLj9Ju67HRMPC7wJItNhejgHzMXKObfsbG
pYCZ8erLeG3njL1tQ7kPUeeguKW6NLOp8p3S6wM2wtCiDcVjmonOV93+Bj3wb8NU
fVcKL8/MJw9DM6AMJHcNU6BKxbwTVKGT7uCFb1gzwF3iHjpJUuZemJH9NQA+qZXf
NQbTKbqFiPSK6isn/vbM6W/fp2UJZ1rYg33ozfkYHAp6vvEf2/fuG3kkCPX3dk6s
sTwVshQYYuRRANVo6M1EpabO2/DXUa50WLxdWgJbp6Mjs5IgEGJ+9PQGPmVZnWv0
uXTMUWUzcarhw3C2fpJy1gvwqo4FDA1xHWj2MtgKFwK5rHUPUOXbq7qHaEe+eU79
doxG2truFNe0vUrVQfiqAQ+4R4EpOzDOxD4i6kcxZCRIBltbIghQnK2Rgr1pgSms
JyW8fYWRLmNLmrkHPAmzXXbyOCBxyezxdmds8/PU4Cuy6Ys9hH4DM9rjfBkQZe4u
yXsj6oJdHW9cxq183CA7fOdJdlCSZNoTCcMl0KcHhlTwZsZaP8/7cFBUjgJFW2ry
+rr85QrgSc/ntYiOM+z/Xu+4Y0HafexT1KfvRa2ruR+lraosdK6LV2Brs3oiW16I
AAsUlm56+tGOKy2EZqKSYURKoUhftdz1bCw4fMr5k8wZuv4J6vbnzBpsm3IIg5Vu
yx7Z3TVay4uE1zHHJ4YdMmWYyxknLWSrBw08btexXy/KnEi2eOmJ2XL8vGRWHS9A
/ThgYQ3eRQpc/Fem8Cd1x1rqPJKFiKMVqG/A3tlYzfh5E9FUqr16j1SAKxgQ04Wg
Jx5MaH4J5lXQ4jKJ3owjAXn3HZxILx4WzfRuRmZIzSdqTiu/f8YSRlENzN0OcTRl
2jsfUVqOMUnY2rY4jVOUcwL9DSYisaAQG1+jHigqsWy7yNrRwlCFhXGk2woRK0vW
qNSGQDMK62LG1xXqdpbyWPUUffEIyAh1u9jexYSFxH/obCkuRLTYmC502QZTOMf9
g8XGD2AcIVLsLS/6ZNElX1cWnZnB5Hn8dBRAqVJhH40C2EGNtq6j6VIFoVdGHwXy
N66QnEIorDNXWZa4/Nd3w9wrpwy/aDPNNERtv+s5CkFfy1T69KFmWmgnl6U36NuZ
QhcALEEgBhuAmyvZLaCtZmaVqGFFeKR8KXwQQV4ZHf0HOevMcUYzZa6mvPq0cVLn
FGbUD9mcEhPFP/M4oxK9eUJ6mzWYm1vKN5C5W3dnyGcyNMNJ7u5zcYEGAdWSxVLm
6iV3HNEEsXzIimRngXY1ruqDXZQ12rqcBGF0BqBtWpiOZcd8gKMMxaWwf2c8Wx3A
0vrf0Q5pma0jwKV7Gs12wNxD6w9Vjh3WLDl5sBwGE2T0cQlLwls89C//UuOjgbVo
K1PWL/eHndCoQiKdlVql86BpKT7xvFsmQOI+EIVi+a2oxlhpaqNTSQpftxCaZYrm
AuRw33D0OhpOkF38bMvz+1m1GxWLvazEQJdlid+fEs3CPbbx8U2dq1OriQN8hOkx
jSuKNwDmrKCKaex/lU/ExpLATRrlPiJ5gZ6giYO2XchwBTjCyEpFEHaxfGvfbSC/
6ug9C9qiolkpCjMrWIQdBos+8jbRZgm+2m/WWKR7/D1LH17L6pTKr611589IyKVn
vLMSfibmbKBuaEzjjur/5IDTYLujg9DZF0K7HqiQSbNuzrKcb+FlGsKr1xtG4uCx
3Sq/+s64l9eDHoEt8o9A9mmHFDF59wgajNU0PtDkhN98zDuS63lNWmyg8hNJLti7
hj8BxXdLBKyjcotYmN1N7svctmrXp2XGDyw5nmu+yuhOe5pO2WDCGQh6aCDBbdKX
hus/YdgYNDrkQxLdDI8oXUShIqyXZFLfSplH/WCTOy3BTo3K1ki6ube+gBdRIqel
lCOyWULTyyZLZu5FyCauq+2VuSCJmIcVbnkXOdyqdb/UFNCfovcCd+zjxoHPjQXZ
5qrxOfhl703IxPLsW0s/aAtIoq2xgIr+hjL8nbO2X5zagz23xU+FGv1RnjgJfbey
+FjwJkqbqLjbkr2L+r7P9zSr9mtAAPoep39mgGyiBQzJoKrxZXyxh3pLnC7g3dbQ
xCSthHAswIihn569s2iwsZBZynYPttRBUb9OZldgKYEQFeuqmupKsqlqO1C2Jvy/
4bdL1W6InWsrGGO7jE5L5UPxlLNkAy3pIJgT8eEJTcJWOserDxIUhD43dioA55Q7
1zuDA48GagxUfPxnpAOqiQrac8gLYXuI7YIHSy+0Jt5oUdj/rfL/tSeutwpTMEHE
mAw8OteU/0TYozk+6lrc7F0xQ5zbaxMWTN9Mceb50tJUUSXqAeyFPJEfvqihKjV8
N+rKqVMGa0W+E8BUj5G/h8Ierp8FJmPbwPDAq6loipOdS84XP+AV7co4JKx4lwcL
G6CjP68qI2MdQJR1vb997sY03hb+ZQYYVJz3OggQUA/TOxQiQs6dlBIx6b+XtgmK
thydYDbPr/5kdJkCgFtOx0kGsbfwu6y/leoLqN8c+IgkY9EoAPlMj4PEpk1eBcWD
v9TxE9Z6VDrRu8zLVD68iSUo8USktYZMDzT3nBoHvTO8rWMAHVb8gB4IeSGLBg7H
TfoeIQJ+sBZEFV2XqZdVWIFkbHRWQaOwWrZfKPBz3BvLmC8a85BPfVpdgBK33nqV
rFclFWrNEgwtKZXo8ksMH19hZH2r84uChjG/KBQuZoxT8YJVL2yVPFSLAbngH2fg
60hfTP26B90xIvpo+2uQN5Fn00/wwJfp0PaiDnEPk+lWl02S19TKZxfxDYYP2E9M
zK92aLB4EdbC+qoZ63549oo8S66cXZoTIAtzoKmj+jq3AKHhISF3EhYEPOjsQQ0U
fUqpCCFy6eCZtbm4XSiKa6ktoJoBp4QbOn+6s/IRN5dy5SI1thVgHxXRro2fOLo7
4nQZIthto0maM2mslvc/niJdBD16UJawxAcUqVzoZnh8mW1b43wUMRiTaa/hin9A
kOxPrcYg64rBRtWe4LVvk7Sj3VGO5QIMwarapXAZYNbk0dXsvFw/UvaXdJV5Pn1M
sDSeAyXZVDb49KEQM8melJnR1i2M/ti8NRDOP31cU8/n3TtUrGJNqOt7QKDmFvDZ
ySRB5tt44T8kK+PoGczKGbs3776apmKV9saeEyS5ZLio+uC2WnT1LwhAyn01k3ls
v6JqlwO0QGkjj5WWeSNQX32TpvLNf3z9FEOCI1JtSa7XaiW9kRkkYOddhUaRiZUc
Tgvxe1Vws4WOYcBa8DPx/RRo95KN7qxxDnYssen24tdcYK1Zrc1qrTmnCgTo/mb+
bZu4+Ow4Rw+a37mefKeOGFd0N3ykPdD7f/tzFRiR/Ny1WT+dkfIc9SljEI1puuNJ
1I5sCUO7cDR4p3ephzA0/5EgZT6HsdSgEMjgdk/2IfgW7+0A5n54a5pAmLsocFHc
AAZk2LGEafqepqTrmXfKZ7eB4Fs+qTqoP8BqSstcLgD7yohi06xWM3HzCSEg6yPZ
FAJ6PBrp7sTFd/ETCrV1lHs+uLZ+J5xNwoWZbkM5qPCGCtCju9hnDN+cA3fVFSTI
3OHM4s8G4rhBAOd4Es8Wad/PnJz7UueAjXJdY+v7jZ2qFl+ALNVDGw9+SnOAB4TX
e/Qf+ceUz4IGMM3vh/yu9wsR35LAgXAAvPeXotlzK0H34bfEyAaDdjMCWVuxqrGB
4Arl0DclOYVOJINHMHN5Qjx7VG52vyFHcmOKEWp1gJn7Stg7Gu/mrYgOesLoN0qX
XF81pu1PD0xoUyiK0NWssN7MGfrufJ6WTcq/qHR5YhQ398kbWzuotM6Ect6YYsWf
jP9yc0BEdjv3chOkdjZcLa9iLpm+U2F/YpZhTTbVrzMnlJiSF1v1tMOtd2njePzJ
eDY77d+DrrM4UVo3NnluG+anEFRhV8xfOG9MzuqktpDMBJNsZEef6z6xBBnwsPup
qa6YtJFfW3w1Moi5QfZ0x05QHi+XnbzZ4Z5cW1d+lmgi8tGuhYuSTDPbKfQfyKy5
eRRh/o9TKp6+gtuT3HB41F64ch172cOesnoOWf757KQ8gV/YA1+mNM0PQCBCCjGU
MTCNAYdaDd6+/FyyBsdGtR8x3sn4tKoXk4EwlX12zLih//sBSIMl0Qdrv0HQ8cSp
4tR8V7x4SRk7NPL5GpBabdZ7D+2MFpenjQqHJfiQ3umLSdmwmNTKun68ZzM3LyvX
KymQXVLYfyd2CLM691QCTi9mhK9FZKX0b3iBnycoBm181n+QZy2ykdfuTVxxPWza
jV6KtVhmAIzsxrIMp+WdsLH3nCzQ0FsaiTuyQUfJT6ri07HTos/dVyd70a2Jwv1q
QTsoEkwgL86jKxgxo1y7H9FssUE/wVpBQw5qRz2agBnbRUzcTDNi9N7qCivANcyT
2BLQyGOGvMYdLQagcT3O9ihrKzHTj5GZE0HUtjdtDyCcOpBZo9la4gSMci6ZFQxY
LSuUnRUz6HXamS+a0xsgOcWKa14zRBKssV5kG6YnK0i1MMpDvv3AIvN0ihPzxAi2
2tPcP2ljCPw7jqxq6kFEpngveRkk7PEnS6K/cJ6PIgBWeTIzr6RAI/2V7tWorWHc
eOp27i+9KKzXuPUjw6nKoQLxdqiQb6x6kBzQN15MjU1F/Ah1BbkpChiJ9+KGle40
rG6Pi5UmJO71372Qkr4+V0vhR7IYMKYsgeWozUc3p/77QjiksTZ2k6M+PpUvM39v
rok4Wdr1wmV8wrZv3yy+c3VsXpxpZSsBRv0vaMKxmkhgKCcPfJVh1rYUUumNhFbf
3x6/WLV+czu4z7Yb4qEHEqTRxdzldiHnG954inZ4/BAIdTtIO9kSo3QyPD+MSeux
R5FiZPYO5jdn6dJXixJ7Ex/5dSh3GZ0aY7vnzhXO5CjKC31qRBQIscHje59+87x6
W9vq9r0tw7AfYvoJEltUqvLyYShDbShqzscQzwrc8+YPmiH+SrLa4pxww5xdwDju
9mppQdxtm1BTp8S9K4I8EMZdfczLZvfNfQet1p2pUYzC4Nmzp5wqNO0eENVyXuqE
0RLVv6xH1tBMit/lKNIFJ/774rdo8Bxb9GtIRbUgS04di79LHCUwxw+zJsBkDe/c
cMBmDLX2UVTCBnsJFSuu5jTObloCck3EwQwzvRJuMUHoneJCbLKudPEgBLQV0PGX
arJP5Q+wzjwg4URLiYrzLRQNniLsdrCIT0frCM9P/IN4SQKpQHuT+VnJ0GjtvYOe
5/J2ob2ADd58JatV0LHKmiMQ61FAs/7BnQYbVAQketbBY9hAfb/2Lff5O59/gti5
79uwuMkJidr+xcf7TGPXlvD/hSHDZsezmUTklS3yUL82F7yUQSq7YCeYfQszS4zB
Q7Sw4pF2uKFOgLVUxmktdn+xjvUCRQMV/+Gx5+kCSq9L7Uam4rgQeWQZlTQIzR0J
OU3X91LVOtI8jqH9EOj+vedmbpnALfHPZCWrNtMgNmm59PQXQRIljw1HYZK78/01
T3PC+vCikECP3JF9B4XJxRm4GCF/xO2icFztdpCAOJOU6k6prlKh+L+u+HFLAxL0
ioqbXdXJMMLnCY7E+RL/+98g5pdXKBzPmBwRDWPSVtw8OeThxosQEsn+JBStf2IY
NHCP63ok4PhfyEq7DzyXv3CwFzkHsd8Rv+ZDJkr7rzcNupTgrlEBURf9veeEaEWm
d4mekbXQZfCGhxjHiyQ0L61+Rrb4rGL6X+ux4vb1cqbiZS9YBsvUtPUlShWYkCHx
1NzS5muCM7kUuEF6UJerLeySkAFjHOluXAZa4x714T4dHZT+sY7Ub0N0yHtoCjRZ
/tW3Q2Rb+A2E3lFNKWx82LiHpHXezSY8BRC1fekN+5ZDR6XzX2gUtZNHJWVxA9ii
VySTa7Y5VfDsrQtBkBmQDxOj0tlBrg3E4f1kOeX10WB4qphqIGwCoojWuqhcoFD1
I74x1HIAHAjbAC+g8o6EOTdW+t36tCbjsqPXpVRYGsBXqYuaWoafCGJEWUXHFKRU
u4lmqXlDfoyrfmceKm8recQFD91scg5p5A7jb+I9A18DxowbMTmJ2NffW4DlsNsI
Nm8SenoOrA+zN3zgaPBnWvft4T7e9d6Lh8sGsb782BLpOuRXvkSFf2DuC453ZuSs
2k88bOwkwe/YyIkB6cw2A7NoFmDrlOc9gDJtVEcGcNogtAa7/ZHnuA35VxrdpCh5
/BWNp0MrGtONe5R8OhXokNewRf1MNREat7Iea9L3VAecadWYSqZa3Ouah4ByQJTd
9KhZUVFoYpLxpvjkvVOSRM58Hs0o7ft5u2tKKnJmEXtqMGyrjcMlr+N+NDvQ5dFB
DE7PjxTR2GeyFBMLTyOyosAekmMxJ6fi9vgXA0eaOotM6YBfR53eNn3lcRis05nb
XGcM+RCdNcWuRN4ZF1fKhkKopwcaPKJmP1wipgXeJptyCbuszNsiV02CJIx5ezCC
RSUiKr6cnFK3TQFuPsNX28WKaGbdLAmGvixUBiFbU3y09Y8Iq6lS3doEhlbobFTg
xyezuk7YRXwUJYYR1ImR+Np509q4gUe9fgmxo2oRyPLWj8Ri9NtEh8xZX/HP7kTZ
t92Or5qallp2dS18UCOH0aDasAawcX+ahePYcIXqqVE=
`protect END_PROTECTED
