`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uBPTQUXTUj2xgntxKTAUoc328yVjU9TRyxyTkVZt8683Ba9Jk83aw6XIOzPysBXi
xn1F5wNBVXNtcXCctoI3T7mTsAcYLg7fP/FrO8mqpq9ZenQaXjds9PQCtNuqV7yp
2kNBffUXhLQ3dzefeyp7ALCkjzYOINqVSvgzk80AYGqzzkj6ALIM7lr2YhxsBq1l
GCfoQjXusPI+aakK/4AW0hXHTZr4hH/RCEC1KCO6SMW7yi595UO0s4R81w8WURZx
G3rYnWbpPSwmKik3hG/Vkf2WwxYltsq5yZjaK4Yk6D19Kw+V45dsuaeo337OHIRG
uJSNlzngbsXJ5FsFlrPhFg==
`protect END_PROTECTED
