`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nsShittvW5/jWs6XFvn1YdCWuQb4mjzeWn/XEbDZe0L+yDbC23Kavoj0LQW/TP9m
arCBzz+Hw8jBXZ5G6xEGelafp0iDzZYMWup5/CiJ/tWehHsPGSXZ9mXE07UeQrzg
gUdThGLLJ41Eqvho5LDW+FmIJTAIB3h2ndQnRv/MRZF04SP38e/VigEhrFdBKikC
/gRlPhqRMSTe6rf1syuhAhZYU1lLxaXSi/UqZRgjZh36Euxgm5b0quCtknVkQQsJ
yzqQ0ruk9VvVBRh+hgu98TQHPf9rZ/YYcaDkTQP7kiKrR/4h+uf90b03yPFYO5tT
0XGFPNv/qvIm/5iGJbD8PsYGCKH3vTXprRTjjXjuNiL77h4HbGuccxtdcOjo47Au
VrOVIQKJp3E0JYsfWoXrVAXpuyBCdajIX/L26qX4fRhKv4JxwoOOUXJMiq2Mw+9U
RfI1EAvRKDfanEkyU73fU8Bdx0D0XRmOiLTjl6PF66aQ7jUJKSCGimZYrx/cyvli
hc0tfy8RuEyVqATO7BEjLAYsCJeJrku8TabErADGo0tL4zkeTeTDnzf9/vo8SET/
E4rWFn3+IQ67iwsE+hUyil19e78jF9iDZF7X8d/S9EEHJHZRdwLLxqsd75llNw2J
dqNPGKKBK146YaB5jQaWvm+AqFbHh5Cg4NrAdrJf4btJwaE4BZ/o/v/5zh/OUB7Z
BME+fLMaHMWxsFC1PO32mtYHNtPUIYqe2f7a+9LKGW3ogqTC0CBSLHykgl6GMljB
E7W85P0j0acVwJ5pCRNkNl+b4gR9PC5la2KIIbZbV8+cCtrCv9Cau/9juUoyTM8b
CLsR4Mz4N+8UXObxhbKwQt6ttmw9Gv402aQ38Ix5JR04JBG2RsH5+ONy/78Xiofu
QiBEiPCfM6gwb+XaBPRFuENWSEK9XUXwqM/JrX+NEl6XhegwTXdyibG2qwQ5HIdB
XQ6GxQhMZDFekuyfSDUquBj7kAbE1ZZn9zTSekF0huMEUXVSMW7993SCk7OH+GDz
zIxDE+ec3a0TYtaKbbF59UOZjgrHzxnzbUCRSWnKmcBUrCHwJ0gPCu7/uNxycOpt
X4JRJpQxL2JjzfMI+joJrYPcIlsIV1OO7uF8Gldpds3UYgOZaPK2YXHZdBqG4Hqs
FUkSInNV5LbbD7CKYJ4k/3ZozXbzT4rVMXYuk7Q+mjnEZa58uH2ejh+5oUe80PJ4
ETnIysLFxV/IwRcp2iIs5sadN14hy2IzUZ8WPS2wdEyK5zJoGd5V/tnvqJhkUvcf
8B6weDURdoYRyZfzpIwHjvj9SEZfmQzP2UpSdGUVLri4ovxqgbSKBzaxqaDkQjDz
AYBggj0vb9GXIPhHG65uKN6Uo+wX19UoFzAP+0GpCvMrXrkZGZLVv4D/8c0LFQGr
7K/dwHm5L5y44ohvoGXPqmKzMMlAsrlDcX9jLYORE032x9V8SecoeBf7S/I6T8Yv
vCQrQRTIyCj2ju0VtdU6B4TAu8BXt4tNdqhY1I8KT/mr3Eja5b3CnfEcVnr3yyDa
qJSxTgNBN62mvWox66NddDCX6r6RvbRkfQ/TjJGxu4Gxj1fG1PWuRMNdYqQq7Lpt
4M8T2C7GiiEOUoK7xkKkw+urKi433hnZJ0UZ90DSN3YjQL2trqYdxkJtXxo+IR14
g4P9TxEXCJ9Co7VzjRKc8Vdbu2YybgZG0OGBPre+q/5wO8/5tAB8kik8RViyCfdW
QwMLc0lDIW22q+ntsrfXSvG1egjdQVgIKx+gDD2BUZdH+qAs5hJPOlbAKx5IO+sj
PIlPjQW5FbW2B1aJTZ1yM8SyqWQZjblKlPWuKoOABksaUYEQ5+3X0Dcmv51hMNQ3
81ZxnDFkwRpX+D9Ev41ckgVwQytkxcaKMa/UzuGdMHfRWbbh8iD6EJFdPhFlTvWx
HsAqMn5wtL0p0nqAeyky+u07Li3ujaL2+yfqDTEOQSeFR0OPIJoxC5sd8nlBZMWe
3LkhA7uEFQdn4Tqjg21wcSx8/lkXE8SLLRwa8f7RD3xWdCXRCbjTxOAKgov8OI7s
RWD8eZfeAohU/kAkQAYsC7cMVCdQY5zBjD6Y96LE/jg=
`protect END_PROTECTED
