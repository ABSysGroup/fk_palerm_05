`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dKcB5QbaV6TJnkdrS4zwinZBP1KTYTk0NTKPwbNu2cGG9OpQ60o1UhrYxLR8h1fw
AG7lEzHXVah+JjF+WipmOI/8VwlDYrwJvLZT1hy2/8fsYqcnRzsNaDCtTBV/a0Ic
NH95r8N74FKTwnt0DbuLYAQg2i0FyzwFbQX8M1XpgCRtXl+y66cn+5eScc9zc3b5
k42inrRi86uWsqqRVoAUYxsvfeOIhFVk6GfgzeY3Gqfpr1Seo6UE6bFvBaT21sDR
PrCXaiHYAf+GSYYdWSfoSoS2TiXCT3wSdlv/jBqYvnN4vfUFyKbCWZunxi/uiZcC
prL6Q09s4skPYiDgSpi3IjivwN3HQF+9qXepwOLhHoWKpyNIklEbjO8QlRDRkmpH
tdIpCdh7pL1YSntd1DWLirGX8FYxbZWvPfIQVW3RMHhGbbnoSporlBEzLSOKtYxR
kPiz3OpMSg8mWINsE+qXXIWJe9qstABnHDdjEMH6FiRSC5W2mhHcCWbbK7PNNKqL
FDM7R3wZGrjWAEucGv4nHBuya0iOs4OBWpxcLAJlQBJeR3gXj6cBzdz1vAOvmpnC
PrKiHHBC7b65nPQoV1kInM9zVcKBtSk33yrUj3ellU567zda7g5RsfSqCUiilgbh
sYBRfESZ5TPn5YR3jrverkxkdK2CZyzW6brOndOvLyEkpoBc2qITTSiKyReEZdX5
/7Xy6OQjm7v1PJzrcFpoaHeh33/jg+QYz7DN4tinGZXDHSWX7hELJqdsXFr5e3jz
IH2JiPxiVG83Bm59k0hRU2wTuBc3Wef7DFw3JNUSGuyqoVhN1Wvi5sDhFLzYZzBc
hVNRNMS66QYZt6YTO53fJFakm9pSkk056cdjtuDPLsazmrdfcB2tK3MSqlXRCB3U
/DGRrUoh+VLb2OJ44NqCd681xbZvd9IvXsJseyWcY3hb8+9+M9j9KeLhZMZpYE9x
GgaJwbI3f4yhJyh2F7YWlnBbhivXDWtOv28vrcvRxufgICj+js2iiyHe5ZC3ViGy
EfYIpG8SsPffSumSkAdhtdzbv3dKiBlib1aPpMYyoOEyGsmDB+7YWXaiSSJwZSUr
Ugr+fyBFQDvX+l/tyMDgjn2uBASTz++gAjQuheppNoB3OVBx6/W/FoAFpePazVVC
/tyJQJ0S9nNwUWk2mdE5I/33SEIjL34hEUzdWuw0a0yGxr7upSRmzvJcqRTx26u8
RCJj0Yopzv6Revbz2buLmlVtqzo6x6M0FBLaNV25rtAQUGp1nEewlF9eQFLFwCoT
K19yGb/4oFPHRLphRO/l6YAUDjqz4ObcySt1eDibJJuV1ahESXIRk6s0FrUNt+xq
oiR0ERI1GsdI7LZHFpMv+yyRWKutd7fk/OhgCF1kQ+b1Tb8YRnXuhebhpm/qlC39
Sc/+SVidH2vECtfo61HI58Qkce2BYCm33jzI05Obp97f+g88i7rQFj/O14+HeW+c
dK1pl3PxyEr5uqQAuuuJ65sK6m4QsPaoCcHByVLB3q62Zi/2cU/mqrwgo3gYTUNs
vu8JsRWkD1w4ZwFyAB5/2NDAdB93KfWKMuX9llV9tzrkmrhckW8UU2Q9F+wbEswC
TFruKkX3P6FHWJ2TTtDrsKAIkRH0YK+wAUlOTCPUj5fR0TBcD5otX7YGVaTmrMT8
Sr0TNr7MBiRk7Fb8bUZaLWgSB4jHKsLSzzvjqCJ9TTEf6GQWNAB/DFqRN13mP8Zb
4fjTxbyX+SF2z6vK/qiHBKrjE3F9cHKV4An9VVm5i+cziGWotz4Ot2+FXgrM+4Vc
wyqaWmum6Q0SIvru0q/EpCl2VXvNCsyHvqBFcMpU2Z5NdtCn6twh3kjYfIVl0A/S
erJRkLZQEegkdmnzbKpmxeI/1pd/N9zdHbNHmbvue7y7ZHrX2Krfn+wCoHN5JDkS
6MXEN4kIpA4dhgCQnjHg6JolUZ9PI/MHPU0seVyCzjf2N9+xcfImThQeOXeGcxPS
K1StnicHoeoW3QlMDAyW7e5QBJHj5rO95doud0Ihu2VNL/4esCRK1xA6NlkJNhA1
1TylnbSoPZd/0/HGfJ8thYSXBhqjfhdnKUgdcIp5Jiw=
`protect END_PROTECTED
