`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5K3IPLE7zbHx1KzoCUgVcrcq1h8JTjYZtBY5mrwDUYQPvJCnM0Dbp1DrJvpNxVV4
qLf1mg6yNtZJ8L40YqOgQyfqQUFcegu6398jPJ8pmFkMXK89TEAxSYCZC24LWuan
Z/TH8sCNqO+qFMlALluIrVqCP21NQWOxNrszp0+jrX/GbPe2wT1BYw49BB8l2nSx
f6NcojmnpSTri5sVqSLrYKk5m9cFuQUhTK7aNZpnxSdJelQRUuLEhdKx3WeN29q+
aO1f5d6erO75ouiiaTtkZ9rJHQSE93kTdvFZ5dJv3F/vUGwPfxdUQTTiLuFLicqq
keLwjGYjxpgP2FKfVm3R0Iimb3MQveSNh9wNObIsllywvGv5r+7ieSQxY2GjNOGe
`protect END_PROTECTED
