`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yl9ruevE6pNccknuRI6x9RDKglSSsdAHn0rVwwaIdMpmdIqltflY4R4/QEndqqba
nuLTabgawsTykDK5cOapLtQVoJPsKMamCZIpltJxF7wtTi84rd6Jj8WoaOoeGHiN
QrKJVdE6E+moI68QaPPfwih+CoeHMu2j0FSVBnn5ef7LXPsRFLB6QSKCXVGVltJI
OSQP1ze8rdDd8max67f5o17wjHhSvRkiD94B/lbnWCaqW3724QuttC+/BuBkXb5a
2yUSHZi79lOtxWw4OgG34dvGs/LMyBCYD4q35gu3kvPGlGugVv3cXliCFgXMMP24
6CeQOsi3pA0LKLLT9NByUgtK11J3YL+jeV4sJ8VABKMJXJ9nfRfgM3xrMBsrAzbo
RbA601fezMovHRiZY8wc1l9g7Qo69It9YzgWVh8nvMlvP6QzxTtLWmCBKJ+onmDX
RzVrvLxh9rEIDIo5vmNtt5lbs5z0ia2AyvJWQsNv1hTfmlVF+QWcMjOcA1ukFVPE
r4qZMQa9YTWI67B81aqQ8iQcmoHGMkjOSVCS/LbxRYleiTNyrSY7vKXf6aMNjnOx
joSdwbbblbDiMWcxxahxlA==
`protect END_PROTECTED
