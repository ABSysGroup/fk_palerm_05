`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jNMWvJceAxcGV+j3+NxzT308h+YH7Qt8QjXmwn8rGvkaJ1VkVgyJOpp5lj+/iIKd
ln65wCqHPxEOeWRfyCuyyLe9qPtLa2mv4a3PvgnIdew7V4ZAS1mjHIdKQs99/jmV
4ZpRS2i7skaGRGjlAFWiseasbJzhDzy71WrxF16RvOP+quNhQIGmS3zY7VFe5K3m
Cjq4dzpytvmjIMmt/0+TH63z6uC423DMGXXT4DtSbvCiLWsTjcYIRPF/Cn9vImYh
Gu8E0Z3AFgKtHp+soR/rGU60plzbmt2So6s72IUThx/6GtSKfUMNCNjo2O6yMJdN
C/IGLqULypRWAkBIOn+sCFcUPxmlc5FPns4prsK33ysqArQR3fqD5N7EEExCuLeL
mbid25tr3hg4zSqwbTiRJdelHyiDfR5x1Sx2mDCjcE2mnQTrZ/ZeCX0cRPvan9Va
DBjJ/TEFZDxog/TiLig9uyP4B6JuZjp58iUsVdEZT3bh5BmETuvn3LJrlr1gCnNq
GC3wKMiPc85rto8b0Fhd6TtpWqLX1Hc+e+A6f9h9Jmz1kpjQWfWe6lE1gEer5Isd
F4XoTl2XxfkdavM9LeX+nKrfKGUg5pQZ6Eq9WHZUfYMKr0RdLa49EgXiKNHasgJQ
VXS4GGF7oSCAiPvSaCZ2FQ==
`protect END_PROTECTED
