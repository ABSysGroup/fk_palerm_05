`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LlG0dnQPNwDR6kknN7cmXVpIn62AHFp53xPLpFeC5DDLMt1PL/Ph+Z2ptWd/hY5g
C+7UZ0y1SFT6IJIa3Kp+jPumPt/2UdgKGaYthRPFEz7gmkW/78/Z0VPg3zn2Uj5Z
P6ZZWjD38kbhSPsq5bOGWq1zerxf6Jxf8RStHRaR2FL7JbO5Pjo48Bkci5e4qIYp
Cr2a+BNcokWRK1JF8TAaGmVAxc95MFpYPz1VcNooEvWtTKdSjm29qOYooC+Dr0Ox
xSCSp+6r03H13B2i3Y3V8nycLH1T2EWLC8giXGKFqPJ7aOqFAEC9UlLgu+6y2p/s
lT20yiL+StuuAsAzM8anp8DSrQBFCuOYR8YcOm3nMuvbwIuf3+/NO7IdSGHenYeh
72Xsv+1o4qzP2iCuqPpF8LrbWNBAzag37qtcSTMlRGWfU9iPL6/BO57DQyy7k/dl
j4fkFz/9hISzFSWJ43m5uBce7FI2zS7yU4kyMeOxKSiaRFpbjkYVeXN7cGIhY8tb
otcYloTBs0ImnbK0kcjF6bmuBb6HWdfsvEhs6vK97SY2RoQXs40M/dpVm8Gz4ULF
LVZbtRZjWS70dU7DmB3GecFk1eaeGf9I2HBxX2QacuFfOmgipnQC2XCZ3GIPBu3a
GUVixesRVmdSB4spKopT9nRyKhsVxzCXpfBXyRcp5m394wduA4iNzLjcWAKA/igq
`protect END_PROTECTED
