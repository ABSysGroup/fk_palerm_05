`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W++evJwOQynqqnmvJxqJ2E5aksDbzRUgnDmbQFi+MIRBlEMLeimrAeFtdZIn7+EF
oiLrxPYusTIyWsIQMKAerO6gRN6X5XCAmnjk6L8ofFf0xgn4TZm43XmP6tHDiaw+
tNntJzODS73bGzL8e9C8cLL+q4vAv2o2IBQG/iib7thF69/IoxQvRgiORxN89s/A
Yq50dAKuP0nrj8iNvVnLZh5Mfv4SLgh2S/z7MnKxXEEH/pNpeFaOpPFLUqMrM3n2
PlrifUhxQcXuajrdFfsYLU8bWyOnAbzd2F+5g6VPtTBptZSceDQCZWn368c7ZTJv
gOG9qxsO1Dp6QQHgF1SwFp4SuiAxxesSd5L53EKvlerafL9V2MMm0QRMt0nHcmr5
F6rPI9H1y3Hk6iwfTPhRAjJTvCxpIdsMWN323NgRja7zOIuq7CDQ/74DZREd0wJR
`protect END_PROTECTED
