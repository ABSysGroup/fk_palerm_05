`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DkpDqS2g9btXmLJ6hY57eKYySOBWOdBYoHfcEsTbBz3cBqD82KflecZFdpKWOKUO
kM64IaE62CNXthVMCCC6EJ+bH4CU5ikp64yGPXLTNftB/vMecL/kR4HmxLidpIUf
eH3SWCZ689Q5R9BX85MknrhkijLod/6GNgOia5rIwBB//2mToIy9BzGZnApFzArD
Pr3ITtYAnU/VIla0mYOgKMHFJf8XS17jRLQg12gS1K8rN5teaMDBKjgMKA5oLVS7
LBljUvY8pgcG38/BQlV73Q+V5rcJm7jmPgpFRJ7H3nzuPOsi39nK+FqmyxmZLsfd
w0XWyUbuwI28EElqF8Uthw==
`protect END_PROTECTED
