`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D71v+qJjWEPqDCLl6mvKcX7fdxI3A4i3lRqktocWcDDDlFyIHsTTwt8exeF/vQep
1iyoivyZPW3oCU8OeoIjnA81ogtxwz15to83eFBeiy8PjndyR38U1jFnCD+l/hUM
sDsbjiWtQIWUUHuTq3woe/BtPSxh/+dTw9oHFpqlZSasnkfXPa1qgHT3UnBksleQ
zzUt33RWSTt8aUrLDi9KYUK4SVRae+H0NrmrIC+x5hVDjSEttO7DjeufelKNfAar
R5USiPdNIiLm0WTgAn5eOJfoGDfhhW4KJLIB0/oNvuu3efynWrGPu503HKP4y2z6
PLZO3JYcBRcUrS/wffDb0kJm47OdUtiwA7Eouy1yA6vkbZLopNl+eSkf+8gbLSZW
eZDy/6ttLOWrzyDywPzjTDwbRRhD8R2Yi+hs7MOujNGhfu8/VZyjzDgkrUjBo+lX
C9+RqMoI+1X/jHlIa2gSdzJs03H9P5TiF1t3c0F5X1EPwY5Dt2LnfEs1pL4UoZg2
CZ+eEyWly1HnrjTVdlu4MTmMkScvmvQ7eanRrW1CXR+Lli/mAYhDUYMddvh4S6jm
fCh4Iw7xUIDahQ/3RXdyBLlesY7vRQH0uBlYoEZ4VrC3+D115bcLRwAnyWzft+sR
1bpU49+ZaxnbIg6tKJEhIcm9i40RII/5m0XdedRfGfDcoWadItsE4UNjzqHpF0Qj
BxWMhJSuXVfTV5xOKRnNfj8iNisW6WkgJUs6/qYl1gX0dqazV1cns3jqYAynHUKZ
fAguqk6I8RFJ/paRpL6ZZkEsxuUl0wX81xMyz91qkgf5k2nSE5EA7JzJX/xhafKQ
xDu1B7Mf2M+SWDCUgFrmFPiJtjA/HFIjonZ6jSxT9k7DeKgvJWrCsGC345Lvixyx
PelM6yReRrFYbA2VUuC/SBGu1fPxppNdadGDmyYu+TbuD+paDZAtrBCE/h9A49tP
wu9vfeJqOpIVwhC/reDgZnLakkQ151n2fCNDHTFlwTUKAt2UwLL/KlcKLPZtHGMg
jtZv710xvLILBKAcHZph2zrfr4boa0Kah2AFcbUD+WICQAqb9YXEAu+JBRCbFnoF
F0hIVQQhgp82eH3Q8YpP5qMNfY9kkLHQ7wrhH7dc0SSGw8ohxKU6Oo9PGxSgTxRa
o6UkyKnSRQ61mkWehLFYttBh/Ag3baKd1EmkVyxIGz9UUdB59PRf8FKu3FpyaUuG
V5iIRhMAmRVSjeDiVCpAvDwb9zPQb8Eg0QiVdgAYTOCqxxpFRgdrIt070drMxZqI
QEsDd3Ut/5mHrw6Jib0xooSk8rdNhQAMECnm09pjWXvdobDJTWC6cXwnOMy/fyu7
27+8qJhe1h51rYWO3eLQ2YUFIsaJsYeqYOZw645V3eAb6Pj8HxQ8qIYxAU4/H8r5
B61KtTLjjfRdCf8pGVOyMqqFNs/WHspVV0y3fG1sRiPWOMi38DOkn+DqG6quEKBS
Vl9Or4TZGA/vCvs2AbWA1hJojdsfkQEbfznc5lo057OyWS8rd5iyNzcE6jH/hWrk
uRRASgxnXyDbO2tNuyp2HGVGZ8zR+8BqdlMOvxIYtpI+CYavaZrChyKQ1XGE0DhK
tz1Cmt9KFiTE9kqG2fCbClji5qdtzso5TFYC5DcZaQUXELQNwI/JiKgUXQFkZcZD
OSMMTJPN35AUYc/l8E63vQZzPSO8uB8gqY5xMwy07+DVr05PyOvBz/am4FcxXKlu
4/nARzN9CvZt6qBx0iMs5G2Zj9OXDqjeP1ISu/CTxjfF37lyYry+p4xO8Gu7+MSS
0nKbxf+v5+hmC8SVNqH1p5AD3hse6i600graLhDF9az7sy8syVV3K83Xe0Ut5XiY
QiMU+/iExKU+vr5mOr7/2TGYMfiBgF++NGDCab+EIlQ=
`protect END_PROTECTED
