`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s42MC/Y/CW3Dls3kfh03Sx+7SfMMWwZO9KGqKNBjYiUzLzL09YTsbD0hmXfrJDwh
jy3k0os/AQL2jYQB4DJfYk/UW/YNUR0YkJwdOfc2VTAWcNvw2p+2kH+AageWGkuK
T5WOBirf/CQhcC/Vlrpk7tlgaHWJml6x5LmxWUEf926EJeYL9JBR9LC7W/ILsu0A
IX0eI7O8ZhZHF0tlIFhgyPYxdUwhcwSF7CQ1lEdb3IEIDLcxvIq1x1MWvZBtbtf+
8CJMCX3MjnP9WBvwQYb9ats69v3kERV+nwuJtkWAe1tCK10ErefLxx8nkfUUTXCH
tYhepnpkJv8snWi588hAGt8BboERRTxPLLyJACzIuXNJWSRBh/Smb+rxrqE4QG/A
g/Y0egJoJ8vzPnw43xI/FPQK28JwTy7xZ72zUHwmxU1ZY5WxPLjEXrQe4P36tsNH
rGwmnHGbpMnPbIogRbH57bTsn62s+HDjTAh7ybQWtenl/y6PH8sJtWsqLMSDgSvB
LKkyv5FLF7XwhtTUUrGBfg/aIYNlMyMBxfRU++m77xhF/KxqJj45MS9zew6gpfmg
sMqK/AaWDsZ01i7aTp2zAnBb33m8s4Tagkao7y60tE4jc7/Q8OUA5k0Nn5EF4tx1
/ynq+f3CSka17xwpJ9+iPFTp0c47NuVDK5OhcKnfKSQbJXpRoMwe3/wgVGh6nhf5
KJoGHw0bd7/i4xCh3mk3+UgPLdeGyeWa5tugOx8+CcttJlGnweqXDiC6jMIMHyPu
BdWxAhi6RH2aMFXkSiZNtYp0kxwLOB9zNcHu20aTAbZxSubYC7A43O+mcej8WouV
PSW+SbBKatq3xkCZL9XAE9y4QMKr9dU5WyLKacCdwN28pwxzSXQTBjfk3dT5Pysj
N98fwhgsSLQ8rvqEjAfSa1khudp+envRSWOtxBsyCwOPCKiBOBPJSOXDXAizoCZf
1CxtdyqapnfSIlhJaStwZXEhjG7zvz7BD4LAs5V64yxx+BzE45sgW5sJvNk3aJ6/
jVoKkDIIbAd1+gSHLEq+5y20h6Fx9PIP4xY2fuc/ufJIXs1/qFPPCVC2KGuUZQ6H
h3oE2OhEmhtw1dxHPSqdR6Pg3ARGbWb1h2oP/5apkx997878Pg6LcDCQEvwca0bL
eBjJ/VxEtY43ESE1L4v5r3HT/Pd0frvFAFKHAixShIEnKyElxFfz0rpMm2Clm19t
lGgeEVVE91Dq+Afslg7gu095N6L75c8HnnypTVU4DXgMbu1XyuBhCI6caXg7nvgQ
4+eXNm4jaozOBmNpDY3qYkGp+m4TKd2BHnppqYoCIrN1XSHaxg+ISUfUnRrKB5YE
INerqOAZvtDA7CKIqJFrjbjV6+oGXa9A3D7XW7qyAO7kkH4cyECoc6emP/H5d/WI
ou73Mxn3nnIyfLgODlTgg/R/vYp3+iQFaYaGGcPEW8gJTtwVcvI/ue2XTibHrXhn
N8Ri/NMctuhovUYqaJ9MI9uZAfc4iRZX8dSC7PgL9NF7dzzXij1SUxxnuuOzL8+W
p8oYoc3FBEeeNWtoPD7VkHyQxH9Q77hRHy9OyYLL4UUht+4uXh+8dW6CE4gH7DJE
7p5/8uTdNIjnZNxewCgLH32vpZdGDOnbEIZ5FkNlp/8SKcx6oW1lykApYFb8xz2e
vQLZPIWgWc5q84p02IMvgNOTumabJkJtX4Azrm46fSnUrTsrEGPLwr31kcRcpzm5
qaMmVDl/UDqeQ3H3mixbe7jxMDH34ZB11OC41HSDPPIQiuhwHNiWTPLdr6nCeUi4
`protect END_PROTECTED
