`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5yT/sRchSzSQ9D+EkC33rFCX9a7k2oPIdDrvbxdRBXZ9FlaniN6+GX7ou/Uqs/I1
/+ienAHDR7WKN57X3Uj82fhR3/vt1u1iNDN1AI2lgtdS6jMHj8aPE1e1KhNRY68a
cWBeieiRluzqLVE1qiZdD49CWi1ykS9VaF9rokSwlkTZUXXz8SaROWtL5BBi7fi3
FKvRe3luYqgK4DPDsFR9af+nSPX674bwiT5obfqwTgfQalouCepeqXuA6Aiwh3hU
q/SQ20j9OUp8EjKtnJjda/oLMvH5h7cmwYm36zWmpspxqY7QpCnJXjbVMfo2NpkR
7vTOJUocGCM2JnzOAMr2M/sB2udEKRMm84UOXs6I5yEpzccARCAh0J/FLoN+RM93
Yo8VBjdJd7qS8WIkVvFRJp4yNaXdq1ItHpzjSRil1egefPRgD4JF902cHQvz+Qrh
AE9sjAZW45uAcAvhmH9/vWIMfOnrsGK8/sTZdE+gH6FnyodNW9KGQXsdTH/XZKaY
EWff/7sN9iL1UesbrA+FvL4+4ZLvY6M+byxrIdcQadxZ2+t9qmYBj2m6FltmIrsf
6Ltb3J79gmypV2fZaoBgll3EFmNLikmHIOJwpT1PWC3AK3Wz5ByPDUwUZH5RSfSR
PB5IacKfTf2+stwFold053dcj2pW0b3GRpBIpjsi7Rnflnq2yN7fqNRWazp5XRba
ZUap3jvl4A8Tfz+rWQ35AiqY+41DFfwcsYmeXpkPRdYpGFv84vfPnmKZufPAgD3z
rUb+AUofpTqxcvb49DZwpX+3tB7acpTDFwN+12Kz2s7OknfdpNUi1kkk+PAdecqn
2i7MnSyeaQnWeSkN/333Ag+BXFY4y5QHHri1JhlrTrdN7kfwh2PJGnjpOhekqSUp
m/1mDtD8u+VwTJXvmK/igjBdNAEPAI/yRdwglP7OVpvnKuKws6upugMmtkUWpMNY
`protect END_PROTECTED
