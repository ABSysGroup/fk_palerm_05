`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yA/MStniy3ccxhWGqQzvWacSo7X2LSJTd8YPuYE1lMcMcjbotAN6/ZBwoJQAX5zN
KLpCx77S6KSuLKjM8r3iD80t4ExOoYrXLe9jpEIb5NCAUhwOhTFc/4U+dsVMgaND
pfbeAebUQBz5hvhy0UZJWurmyQMgXKlwXZdSTJQzl/aQwUhOl41WFOJIkwBdcLoK
KDEQLNzCWxCgtOsNEmFMHzm3b8UEUr/VnMkd+IiTzCLJlvzfxg4TztWSuUVR1MSj
8Y2XBQda7K2HLkU5cuctag==
`protect END_PROTECTED
