`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CG25eQxOg1Vd/0lcr/uWuuZ6HgzR+vLh8jjL9hKnDZxnxGrQwDsP0rl+V1kXoECN
DJp2PCw+uGh9Io6pHRCx53heW3TI2c77LD0+NMDhlpX6lZvZ3JR3uLgSabG9YSrM
DKiqBSBMtqe/tdKBIYy3y5n0HkyPg1jhSzpI/BZr/FKInGQt36IcJpRY5OoBHWay
oETcPW/kgAUBuxcga3KrXvzRTmLkdYd7TAN1T06AnxP6x2/j+cpHt/hahjm5s7jZ
y0DnJiwoIaVxJ6nrs8Qz3oTkD1y3896xZGx6FRdzhds4uFmhhnKOiNZZjfuLuZ1l
gm+LUZhWAfG3IT9wRKd5elZBVPA2CMmuTXMQIRGD5pYrHFFWCw55QOROV9M/Gw6b
QtN9Um9koPUGS1WxhKGJFO9sOxVq7U1qW7DEF+vMf11EOTw+rAg0ZJamb0gwLx1c
a5pwG1P2Ss46VmELb6rRlQ==
`protect END_PROTECTED
