`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A89qVyx0NaAvx3ztAIG/wkDPv725OUR8K1b2N7nE5UXW3SpBZbx48xXLckp26qSe
ro6snxfumdosfC2BodBBY/6nseVaBdoovGsD2czKWFXY6YYlJSzqYIG3KnQhzSQx
0IVxcjTMYf7/sBu9PPwxrsdQj2Kpj1vqBGwCLOItsbjlk6pBobf2gNOIQX0MoRrM
of7oUen7DqOKs0Qn4gZYtg==
`protect END_PROTECTED
