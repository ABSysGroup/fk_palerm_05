`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KecY/1y9qpgtJe+bi7emeC0mdDfE7PT+3PrUAtSNOXPSfjNhhrknrN7kf2LY1bxN
ssUN2uQXeoH5GmI4+wSIkKLmLPGfTHvWSsQuUqRrjGYun5fC0r41l1UX6KLhsx1P
bgV1cIusBeNJdnCQMt9koUOY8WQ+IJqfoiI1AXyAC9b8tdarmUBvokwtNS47qSiy
xVuDcULBGSylRSTVlya4Uvl1YAEHTjC5xzfdUbq29s6IbQ9Y0jKntNwsdXnuJ9X6
95rEka6NDOV/w29IWVyqS3CvkNdc+2VP85u+iWrwiegz5lu6I57z9puF3Dzrb+NY
CUVEOrshHXS/BKYDojNDryzbYitJQ3lyHx64rtgzJMlSCX7yUHE7nZj87+N5Yhnb
SOELzXyteGJPGNf/QatnJQa24Qj5vhLUNo3uewBEiQCl2SlcWtuiEonwy47ljyU2
QjmRk/MUDGb0Q6KjNrnJ+HmXNntcL6zYnR4GP9W9Pu3tm9oDq7xo3NrjKIplT/rS
BP0ATYgO9b1wTICnSZG/GxKswHPIWawMbGY6ZmE4Rl7e75STcThBtAo4hqcunyTK
NxcjSr1wfIxlOLG+W9WncVyGGjNuDGFktrYtP+QGptnt+XPIrWVw4ai5hi7nI7Oh
`protect END_PROTECTED
