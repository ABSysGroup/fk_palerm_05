`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3komYzGdLrWr95YYmzJisnlvPZjR8Mbyb1YT2x17wue28FS8C2Za+aXXxuoD5rBC
BLSr82FXjzUbaV3rIjyIZ6qlT/LfiUjAo7C9y9opN/9YnO4fvRsZh0c7FCy02dxc
liLDGETWiqyKl2EHrjh6wZ3RblHeP/tw2g4uplBI722kJcVfL8qLwh5qirIIStql
yqcI1uCHF3vsQT/LlubppBLwI5ymU/wM1ghYh8CSuDmQvPO6qaLURNzCmtESaIIL
Iwg/miSQaAvQH01N4pZxymy8eg2aUiNdaFSzsyzPpd0KoY9E//cVr+QmChWlEEsN
41wESce29hTwF1FljWqSWLbnPQR22U4Zf1tRL8QaApqCv98UZbK8jU8SR3oZiw3J
jTxS7ZzdFJz65e+lYk1vSDdHJE0RvpQFoEsmiJJcgaZz91I5ZkkcCX8Li0aMcU7K
dTyp2o/fEuwlA7O2rK7x7PVFgRhmdAoXSDUuoiwJRZ3XOglPTfEWgfhMG0nPYqf6
0G9yArUnlOLLtocAoopFHY9OMRQSB/gvh6m/VrFtfVawaeOG3wmse3v5WpejU71k
5AQi/AdLro6CnnTM546UqLzvwtx1H9wglo+ElfgkFZ9bUp//at5f0spsz5VJ6eOl
gSKnkFbD5mbkZhK/U9kduw==
`protect END_PROTECTED
