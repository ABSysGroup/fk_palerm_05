`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nb7ziYJQZY24m6xdETUeaa1MNwSEjXQ5OdVdICjV7zkESMdPWyFX7iY5mTp1QWNV
IkuD7/FVXwP/HVvvlfK4ad9OEWGKJaEfHAY8B6UAwTavhyhGbD4cIoFNh0nH5Arq
T+GELAOrRGNO6iaUXJo6U7cQ0Bc20OtoN5TwXkv+l/UASIYudTrDfwF4lEaQt1yg
v5A4TWO9r6inABYogN+TqtRmCXqwRpNv4pXo2Gru5KxtC+pbNM52vHf+siS+YFVQ
TKPKx/PChDsD+HolgXW51eRqiZhWvTE4dDk16LrMFJHz2aNUqNcJiCsL1UNniRbA
yQtKwQNvrnKI63AF/vCRXfnyW3CRysXuZw0Qbi1jy3tO9oj6HoZfO/RG3Xzz5mtD
L7JNiGyU0to+99QyZtlEOfWrBstS1Y6te5kvceyVsXnft5XgaWOwq7zmNAhkb6GQ
svJ6ZuUXI3GBcMO18PlLATOwGIUGk8+pme4YnovtJfeuYhkYulWabxWakPy2scPz
6BPvgWvLXIMN5/QfpGh1vovOfC9nuydxN56UzoU4X9nWrwK6cI7j+DRtap92Ybhu
BZVwkBbd5iED64aOOYgUQlWOKYKN7hN+SFoJ1g6V6TU2kVo/cSuehjgoyQbE+jkb
QX+mTT217e+0KifDjW17yHP/JrCrMqwbipKnzjR3hxzNu0nqfdrvZist9UJ0YoaJ
7AHZqxGW/shvhEdO54B1m1SmEsspfs20uBNOMHK62EZ5LW9qlPXJucoY/0IVxpKM
uO+htC6vwC4ngGYVFJ2ZAQ==
`protect END_PROTECTED
