`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iB10GnqVI5t9NQMUKmgDA6uKR/YeU6jRhpWyaapec2vcC9r77KbFA0rbDJm1UyeP
JNN2MZkxHzh3uvaIktG0il8knGRHhVfYYuUBRFuc48/FcN/e8P2uLXo4dwdWYOv8
+7aGIxd5J6arN3QScp3+uzzpJe+0FYS+rifTkWvX/2N6lPRYWz05RzBNguwlZBRO
s8nEN/oKcqNEQzbBo2XvZKFlq+BEYy3Vnq3RMzBkLWMG9F8q3cF52ynXn8tf7f7D
aauN9kIgCmduz2MMG7Af4SEFS6V6TmoYKtHLKvFFjRgNtuh4AK3txg80awA86JYD
RIAD7ckSoVR7hTXro1EA6IiHUFMSMNK/tW6c5pbwfXzQfEJnQ7RXeJcS8KgZCTOt
wPjI7E7y/A1bm6L3Zl8PMsmyZ1JAUwOmnpLbpkBkZhmD2poiXM6mnTRKXd5uO07N
bP/CYgp8G6/33iORcZeAUjcyQOvyJLrg0jx/8zn1kSVfNlmw9rfaGBiy4SKv+t/z
sWYyaY3Wr4DoEnnN2tyO7y8FJMfp/Q4KPQA0yvcMAwLtvuHD9NQKkKQ38+LPv8/e
eKBe+sDLS6l/ViRHV3///pG5N1lmFRZ6KJmR6L1qiF0EnNT03lS0zX32oo+F446L
kp8ZVinCzWMmRn2MwTr2t47FRHMsMMv9w1jFE+8uvL/4JQ5nLUSocPufuC+Xwov9
gRHNMwWbo8rcITlRGkX9syq+uU2GeEWiqRrVZ23v1wmCKUlDtiVwXgGwDDSLZa1e
UEZNOv3p70HnF66L64QwM9KhJbSWXaozYxW43dT/lrkTvbELVBRUO9kkiKn14ldy
+9t1pAX0rYBIC/29Qn4SHVSL6MbANMPAWdqQaf3RJKg5JbbPfx90+Zs2LpEjq/Ng
y9EttJU2EkReOOsy8Wap+bgdpmJu+cRHb4ZrqZlJLWQCeGERZB+5OLYvpMqQ0W+R
z0FQfgbgUCXBuc1YzYUgW0hxob7hdLjDWbs3mt8xQOdr+rqYTFaVTRgYbCVGvc0/
B200bgZWeVembudtzpb9hBg5EIDN7VjNAjBqFKFsCyXnaWyM2H5INEpfdc6b2lc9
pODpcxYurU+FXfKE8IUza8nSa3KIpjdsKCCTXWcNUJyfEmcuCzknqlDjW+zZGvbZ
Q+SQLtX3YB6Vb1gfT35aM7LE/YtIljxEBcMJt2vRUQrj7dyX6K5TOKGtJr5VuN+f
EWOlZlLuoevr1jFsQU1rHF9DhPDP3/6lKrlqTyqqaY6VCLs/qcZBxVLqh2Kr7Gx+
8+5MY9nURaHu6dn+OC4OD7cWdrXhMzKEPmM1HX1W/LQdiqnyqiICQ2mGCaYwz74t
AID2nqCg7kGDqc3NLtImR18W9symlUiHjzq+aKv7UauRvddJU05HbK+1AmWAnFfk
4y+V3Th6CnwmYvlqnF7UfsL8ePEkNP3IKX2x2vpnpyL/HR1bYZd86QRnkJSsiJRs
S5PbzcXWMSw98fG9cgDTxpsAWTLOqS+Chjw6QH2phlYcByAHtlZ1UlQOe/FPfFd7
s44MAQtHBCjzug/DR+07Wpa5dVtZb4ysWKWXSGoA9/110Ioa2oT/RGKD0ZFTAhjS
J87AyUj0K6xFRrbHWA2i/ULHZQvUn7/djzhaM2bh1RXKtF32lhsz4Mm5gphEkm3b
K8Sr16Ds9vYHmHG7bZWMyxKhFpKIJJDEffJ2na53bg/0v69h+USp/u1LqTxHyGeQ
TYk63pY+s3IUhC0sODxfGzs5h1RH9vOpzYujOqOFL5dKWN8NBCqrlGDqgnhqDmAc
6YNPm8LWo7ajjzi5YLURU+iTIyJuG4/Xev/bhKCR4BQqjNQSTI08JJK9H0kzWira
eYkuWZLJifSt7QiXFsphxutFXcnoLCIrAnwHqdjMRTTPE9MHCwYDjWo7aJ9Ig6jh
PGVgfjEdzxEOEKiJ6Er8KBe96VkrzrvjjCq0uKfYpELnvobGJbbPoqMZk1VMUNFA
cevJr2dAXIjo8FtU5EaYZnV3sMZGZnT9FlmwA0+kgQyZissfrXnBccK7uel0JnCx
gN/dcYqqAHosGWN+Ve/oVc00Q2NW8cGnXdK/+c9Re3z8rsOda0d/bJjf5w5JK1J2
KHV65BO+rXcbZM635INCFBIcCkb7xZPWwwRy81kUsT/sv7Z5yRioGhnBXSxf6gvQ
PHJJ6cTusrLuax/WwrX2VrvQWF0XVhqnVuUHH24o/QNy2Fq1hJELeqkRtPq+Agqz
QrP2bYQr7cR/uPVRr+5q5U/ksjYE9eBGrYX9WrItjIK+36qslbdNu/z2ynOCgkck
LbXbRxe+JhxejczzzkrCFYVmNabBn2ejLLrkoc4xCshfPFq1at+YJQZEAPpUFVBH
EzeLV+jOSPQPvEpqoPYwC2UTkkHgwhq6JiC7KyFqVIP/kIGhw0/dbXxJf3C+DZ1x
1WyzXsXO3MOs5FbLSa4lD2Nvx0IpBTxkEPTLBXRk8wnHpJkGYxLlsr7hDm/qjr4q
aqdD/Q9wP5BNNpZZAVuHJuQWmGhcL6IjJ6CiBre8agHYtxSh/TUNxVaQxaoA4jN8
Cvsqk0rvBRXhIM2UJ0UudITJbzN0AoBGItO9em8vq+ViKjxFxIorJc8p0DgXs1zs
I/a7zx4nVBvskXiECWefG0ha6sCHSTCjAtbjlkMwuzE+FIEVIdavMyOxGH9i7LNF
7cQFjWujfHsohmhcyf1SeqI2yf2w+P4UNJMcJnvchqohok1GqS4qfMADm1KuCEnp
6WsWief4YCRjcWaYhqNcH+yXQ1kLQbFuomTqQ366Wj8XJyy3M6OuN8VUk1Kk2dMp
zgc/QVe1zzS09970naJlyXfv0/V6MfoATrGywn88iaEVMAf0huvb1Uhn2S8mybJ+
4a3M0kc2XTQ/fVMahFuBVncNVN+P8OMOlgRq19f0lKYDLYr0oBzYJWJ/psA889ut
3M9JBIRL5Ia4HZW1fgawktmIhqVLQg2FrUozJtLP26yItKBHfd/5VKsSug15+Pzk
nwYmAKWnMmIF9h66DfaxB/mBHzKahx9THW4MWFQQw0Hvyf9vmfJZuSp+3I7lIj6+
U9O4uJNRKi6x1888giFOQcbFzAz1yde22VtV+hSpexiYwCovYXjaNdG4Uxlg//w7
BnROQTpDjAffQOHOuNbpRPNqYhTIAzV5LZJdgWPkOTr/4zxVuzgXg0Gi+6RU9lgr
qZX70gkn2b/hp+WAzakdnEsTfgSg06T0UxJB1czT3rbgue5mPzntiRlcgPuj2yOj
eWXJg8k6th8429yHyPWcQdzLktPDBM253euHeItkZqH9LpOwpLM+HsFJ+HOrm/ib
GY6POdOsB2maf26lmNCM3CZ5pVI6hAo3HetzROhoW68An+dFQ5gLerpdVk3jO2u9
0SC+L+dH7mZ3LZkBo86tL+vcjucISflT8TDfVs/4jjsC3N5N3/6d1t/VHfl+3OLN
t227kFjQrTd4L5lbk+etbCDJv1LnENG8Y+J8e8Y1LIV3/6EiIy8ZVX8S9tSbYraS
/P5+4kQzH6FAK5w0HmVmkN7vojAdEVwyp45gDYP14WWCl7ky+VIcdCFHdu2cjC0H
AvhlsvB5jBk7GVe/U6Wuu3+MxnTDUgR6WBVTRhs+ekIwLBkMMh4KSB4sbDevZPtv
RSldwe2/+IJ4k/G2opy8/LbRVmHWW/Blt7m8R8oSHSn1ID7G2zY6ueujRSVVO4RW
u7NHitwaiqLYbxW8+C3JcgD2RHCVSPApVWKuTj/MT6nAUcgqPtB4UlL7wiAhkk1l
HhKaXil1JivCBQXu3zDcJOTKYWi+cRnNkKh5g2yvWbZD2VXSRf3pu/TF1wwjV6iO
7VZxlsPba1LFT4zmfqMXKHyfsa4ya75l37Irn1HoAAiWyP0nAXjOsARMppQv+sMZ
nBv8l223PVSUcYLZI/vpFqq3eeN8PoyyCm2iBk+QhxF61hRmDV8kwW61Qvy7tyae
+8y2MjHVHitenCgdlsT8W+onDIFY2VEKZ13f6E0hXKRwH+Lmyv92g7T0Gr7O8uxS
8+KXldHsvsf3/h+WIZfWfBBgTUmYroVhPO1bIf1qCZIAtQmr3/vMCLmGnbpOySYf
rc9KwJJ8FCP59SgHEiQ/9ed7SrXDn5OvEMjwU59p0VM=
`protect END_PROTECTED
