`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nucKwwUMqPdkikE55x6IfulF3q8Vu/PvLZ+xChkjRXEbjp5q9F7z58OyCI0mdOT0
NEs5sJg13Rliu6o/AU+UdkNEEg6ViLR2wLIjbUJfuaIBqzlhdbDF6rJzOfkjFRkn
SWaCHOYf6ONsbDQ43DUn9mEqnxxhgwYBBqUjnZnZIhzYeXdsuDbmAdCNEQINcF89
eIZCoDW7CFcxil/L5MPRb3JItwlCWpaCRNg3F0IzxxJ1I6QFH3iTejwh6ccgT3LW
lNc3xewWhxmgVl/6n3ZJlKSIZHG40bxxwBtkJAsbCb8V31NietU6pFVVhNIan5HI
q+xjn0o1yrIcWqpplgSWkB/OECnx2Fd/ZgVDpzIXQkEGUAQQD51D0wW6wpHH9zc/
5XPWoWJ2wFSp6s3rkSE6YfHfJvEG1p5fcYBGJqfQzyJMdPn9DJpX0FuYRSL4LgzI
9sagxEfob5xszWkIf+ZfoeG2ydq+vbsv7+pqbAX5/9gStAllh4pEeI7IrYe1koXV
VopxKdA+hicI283gw5Owj1AZMqabXUrXGmfEVr0Rz7yKXOgCJStJn8E55hFrK25N
MXu8GnTNvuSoSfWBPem9t3LN5l0alfzUbe0/DxmXflaPQ45U4NwBU8QsMYlg7+f8
AK34N/a7h1V0GAlE8gWnK7/McGwFFPHIgblPNpBuP0W00pQHtQBvr8u5RKJNDja1
GL/+UJCuEZo3flplvx8gJindw4xhlVficWVKz+DR2A91naWZib3elknYSrANw+X0
qbzqPPK1J2qIwDVhyRZRRdDLGA+3/cikhmrfvVaCW18gD8w3xVU3z9vA3rEJ7Lrj
Th0AjL0ZC64XrviBb3N1xWrN1yn7PFL4lIUD8Wds+IgszHyKOsPTs2NfLgKqfjXX
cWRdME2AUwVRzfJ/d21c4I37LiBeg6ggIgONBJ/yD968VBv3AYC7/GQXQuNHa391
`protect END_PROTECTED
