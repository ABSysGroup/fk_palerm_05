`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mkZicD8z4TJ9//bJJIpQ9es0vF5DoUsIA/PlldIMYb4I2Y7GOHIRJPNnsEP0TkF2
XmARQQKW4sSRBrj1OtIa3dswNeCqu3qjlKwoQRgX52TcQsDPKSfERixjolBNcE/8
Gxv+6tJ1tVFRwVWvA8bTzvan9Y67PNUoJrOV9j7Lr/A89BamFFGxCD1ND7paEwf0
2OCN9myDuHT36sHe9uwipkIsOZQ9uYJNrcjGfYl9xiM3MV5AzaKQx3Z6JjPVkvQz
jyTlTkjfthhZwK3BZC0DNfSCxYYyYt9I73oNK602wGgk/TtWoYjQGT4AniID8gRd
xnXcDnHjfoXVoPy3Mxhaa+mhEBNGlkonr+SAZkMvoEvOPy8juYIzGYl4I/wI4CR2
K1pkBqr9m1Qf0H35WJpVmOEQaKVRVkBvEArDOxG+fIU23GG50uM5c3240zKLU7l1
kwE6463Bw14knb0SIob+52tlGdeviuv1LGYTvmnd5Wggv4EQVSRB0YTZZ6yyEwUG
IWQhifGbryRmX/wIomMtfLhei5CYsAUz+47U6PO1KKz+Wp6AaOp3S8R7u7R0kBq6
aktJYJ/3dyRrfzzna/h0acqG1rBOn+HIAr5hYJLDkcUkbwJzr0uMYsg++eozFH0o
XsEzi+f3dio52R9TWK1qKaYogAV5RTaW37fr6k0mMS0=
`protect END_PROTECTED
