`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Roqljw87RtCmEtBAb0mnvXxHgjZ5tJWedR0E1lHxsLWBSrqYPuH8MtQvOfsHAUIl
uCvTqfEvfZp2cJTvzE/9BdsG+H4/ZrEoXgx+8RgXaQYziIfkR3b2xKf6pLM6/j/x
bxzPSwLp9UdNjkoJz3DzQta7ha4T2RwzJk8ZSFTg6A6HolXZs1+0V7zw0zej0rS8
VqJByxllOQ1OItKC9IQrVxsgjk7xq3zrn8SkGauulm/vWK6V7bP3BH2wipAJdg1M
6jCuFkoARFBn3DxbJ/a4iwME6PIDrlSZJ/8gsVN6+qBbAqEaSyDArWrsUiwBmDR/
6pgMUIXutnHT7iTaCwGb9qfvjXQmBp+fxV7lW+R9M7tbSK6Jfpst90ixbgauRS97
T+RD/cCtHg5oFWb8B2cNb9g12A27GueLLOZJbjsZBrQppBrW9BsF1RQttesI+5yj
CKyb73Ijyx0H7ZlIaHmNScxiUNCU3H9goJmDHHX3wnBfUVyi0tC2JFacVw3xTAcX
4CCZSakro7FpvnZ+Eu2EzZJnpxizDagVPpfUv4pexC5dtJ8juNSpBzlmy6w561SK
nf1dpzyzB5m1ahThWMzOvVL4xNNNIFnJJuiXzfHZHMTpzzdyj+74p44shD+Pn0LU
uS16v/49LgaJr4VTTBd9d5evrnVyzbDn+JKEH7jrIJa5SnWswtp2KH7EF7pzeybC
T+cPxitiRNzYVYYt2A3PCP9QcXPRk6/TWpsBNsZ+PfG7TXHnvsdFTbkOQnqFxOb0
7uXGKmZNFxY4G1tbLgjtBMrRi7agB56o+ULfz4OzOkRVOQ6Ai/l6WfYrCdBa2o9k
lynynZIYmDLkBFoAI9djEjH1thflkVX6BSieU574cljhUTgkied0upr39ky9sooa
cEdrxneII9f5BZNZQ9v0HorFk+ZvfYAZ+im2tv9JyX4KGaSod1Z3Zlb+A0z8zgqz
s0Q8WtJqvv3Z/i5GODxoSUrTDAdWvQtT119wclE5oMHugkhYmMW5Gg8QCkEEyarv
fFqxly5uF1983T+0lDYZVdIQYhZwcH3kUq2SRlSTzKUMPSFQ2ZieXgGlCNpcG7ez
FaaD9E40xJYRM2Hw5m57dvZF+8zN1CFJGnRxdSPQr4Ufy4KDDLyWPqmy8pCyCyPw
dSkT42VOxziYPPRz8+BH/jUoY+ZsJP4g2A59sidSUJ0sbN98qlI14XqB7v2UrLTs
9BSTkjOSu//JBkSwA1HnS6HP2m+o4oGnU4yH2p0q+Gzbs1l1WUfrSh3NrXNqV6ZN
/opmxEk268mFbeqxyzeiTsnlLASdCPqs3yg1Jo6SAhBpV8IhIEHt/4AJAwGNU7O/
Z67MgwzB+RNYrTTmfM7VMCrGNnruS5A3qhwFoi5xuaM=
`protect END_PROTECTED
