`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3uMYagA9F+wwRC5nW+IDnAUcPOrJuVU+e7g1S9CD6zapULuq4ux/mjE32CM8vyq/
TAojMmIdytZ5rgd48tRwhM6cr9M0n6ArVL4+OldMBXhVUUWoN30fQN1es50KrCWP
5NrTmXkrVg+uzhn0ENiRvKci/oZP6jTjpPqwXjVv38rZBIz4hOJO3bXP+OZwGryw
lZ1Jsb/IwBKVVfAoQiBaqSexnUuSqFCHZ++pc/HlvP5qU4jGkP+4npyZZoVY9pIW
FfIbmZnsYDNGGo5wm+GM9qmpTjRWctKB/8CHTYzB5c30oV048Y9zCjBYNcPfpw4l
I1IVW/M26VjFFYsADdqLxHG2MSTNI1KEDSSzmQP2gGIdqGZpOMi0EqEuJKb98RFU
DknlppQfeapD34IY17waqPW8RFlvpO5ubtBQqQjXQ/+LCEqd6r5ylZQHaW8d9gtU
1pkg97XP0d4XgSZnVnV04ObiLpCfuyH8JJtRGpbmsrOldi3hmhVib8VUhJYvTLab
ycMfXLqbyouMKxfTByCJOqfmiLb/hYaQ+OXrpGroQQCbDMxZfkgZ9vJ4xUpkhCji
egBYi6yT0aOzeXQvUX373B/HmvNsf81Cx8qLkoAGolszTT5fB+bltzB+lGZH4McU
5HbCH/JQkh3KfzYsPtIDGVe4kUxZUI0YA6ni/+QO8V87jfWaxiY6bSHwkXm25Gvc
ia2wNC2BGRtEmNnOhmB7DO1TsDuCDR4Q2ZlYv2UWlX0qgFqU81aHliTejXiaaouV
Ii1DyRP/OTH+Wbt038y2fni0vjuFrpIe+67kSBKa0yeT0A7cA/8agDfNeQMphNAH
RS8yViuLoH3YLHfHQzIm5q+MHQs5/LQ6LIcg2/TOSPilKVjzpEq3cGwMJzmOvi3k
zW2J+XSXbH9q65csmp6iTN6nKfZih0ydtONNQdMFz71W2dbYpvkSFSnuJ42299K/
Ejova4fnc9aRsT1fwVf6no6lv9SSHlnYvy8GXCFHMYP6MJO9dMf6uf338+5tm5eP
1lQ3GAJU83yn1luMrBn6YMu/wmBr5QGADwwFWkZefaaN+rrouSC985qBQo9ToW+a
uAnJ9cgO07WuFFchCXVEc4AnhVZgGhRgv50a3xZHYt15NNtPf5ThJqPDiOxi+JQx
lo+5QqOw7xcU7ym5ZVzTH0zBXu1opDVSwXtpLf32nirVm4JPf8oJVP2JdFYtsK4k
YEb23VUENK9oTPFLNt1calzxNFqvrB7nGzpqbCELdokHuy9htBQawknqiwaZr+YO
r376aCCDZD0qH37K5wbo8yFBFVpxIZsio8GR9ZzYnAcdSAqRG03xPfF5GO9hRVE3
issZeOHR5EdkWzVuxZ20S43+d6ux6hR7KyY9FMq53Tt4cDemuFqADtwac4zBWp8q
QXXuyQswLirlV/BYaiLcjwTuLSYYzRyb5mAGHS65GLVX/g43S6/4wvrVcV0Og4Iz
nIGSCbthbIkKrfAAiQaG3FgHIwuSM0l7iqNFME41gKz6Lnfp8TnTuUFQ1hoJes3J
qfoT6iM/rtqg56FgAxkJaBfjINPuH3TMiJ6bnAva5rSCN4gXhcdwlIk8Uu8bCM8R
LbbnK4Roq1Ei77oMW731q/1m81x2V9VfXhaWobKGJr19Vz2HdNsYohFMyEr1GGis
KujTsHkfrFEoj3kNwr+l10lZKTe7TjAR+l2gIZaTZrQNuS7cs0T8GIh1SnQOp+XU
530VfWxNtzzgeoZEZBoQgYJAUi9QqBp/mxVxBXcM28OzbtINJslVh2EOqf3wZu7E
QMdVml+Rm6XbSiCY6O1Csv4dQy+E5v9VNLfzSHgBu00ST9W10krfuzonxpTlxYOs
AWAJu4zRSQnXtmo4WPuMIGPv6gUqxHfWKLGftn0BGpjvpLOIOdgTR7U6treDT7An
Wqvex27G/ljKfrjz11d9HaLiLS4JAX3purOFvX2a3xhALq89s3W6nOm7G2ykLUW7
QItxyKjgLLeWbBzrTGgayVJ33YTH7sdCcdcLvxgz3zceHnS3gkjLS/6TNT7a3W3z
Nqv9+KbYiyweBJnCo0PbNCQvfKT+R2xXAllVTkvo5hsG7KME5A6IBqTCGpaLvxDW
KDH0UPc2NXUCWtb0Ko9n81MWQE5YIRcuyE3td0GNCu1j1W0tHV5JOqjkQqhgZ2Xe
AotjZQuAMEfFttv17FhPiAA3oBz6UJ5ewv2DWS4506qhx+k4gwRptQkXkUQ5ecBl
KsfX065PezTsmx6lblkhrxUxz0CF/G8oBNxvm1drmSMuWep2oAlmWUpbOgo1pv4M
nVhRX6R3VCKgLZ7oHgXpjW62LYAZfrI13Ys+5QisP8kzyU8f9j4QYkSorlvue7xM
x2pJsZvVJNjWR/J9I8/zdmU4PAObuEY773Wnt1/V578vuoHMrCsfZ8dBnsNDJMSG
89nuD1XnlHyzPBlfOXr3MGexRXl8GZV9ZiqQG62JqxVoBbagvKo5IMikijRGwq8p
SRsPmY8IjgYgVnbwJb07t1Gph7nYh2tTTVkpQTvFrsGzjOd/btAVFnTwFAyZoiDM
U9LrXqf+AG4RMP9WhpXNTaW6JwVpyKhfmgBPEtHEjF0uyQxujwpHZas2zrH7IWWC
g0t6PU07eVkDe2n5jk8x8q1u0Z7SsaTY6d5eLLTxIl+YFCJ+xq41v6XUa4miJ/eb
jSH/TII2cm11KxtQc0ey+0KOAelpBa/as2l/sNtuIDH9sgKtQA3o8QBhe6J0uIP2
BVVo8AIX5x3Oa86lgiWWaLUAiQ71Z3IAA6nx5Hk3/X+EHwU8GtuRh6uNdyvsFunP
DXUUYxvgYU2wrckuYVJ+65lVj5HZWN7bjYp8t/uakJYsCgHCXBbs4LpBzg7IunFR
B3bF3eeKJxgcELupFRkhLRabP7ixq07DK94jPr2MQOu32IQ5Y1apAnkq+T+Qr2Ju
5SPLV0YlZkmHDCVJ7/27+/uRfCV+gMvwM0buAKnU87lmolQbRx4bYzeWvzGRD3Pt
M6eHsAgEGiY3kagsyHj10Km0zhWIy/zIc1atGwIBP2gt4TcKB1kAdil7CMIGeRrZ
DXs2wyv9OgfggSlJfbR7/5mlP65I7u0Faxz9oaI9eEnpaCm/NM5ai+/UaBiSsNel
kl2nO8LCpNXw4PiYim/mmxuFmjWnlmSnLo1REwPQaVPF5hJIdRQLAhOI5Om4ElEz
1GylGBY20K6HK4CTieoVrVZKo5bUPZ4UE8OzSqlS2GBb/j66UaXx5jzR9WUiKSmz
Cmw7hUIkieGM9D44vExw75O3sV21NNMbweZ5dbK2hvKfLYqyqbQosJKfMJjn5hr4
mO4NZpcSrz89SImMOE4eR7+fHkguKyxsZS1cWrDmapgWocbolFSIkHc24Fnnprno
sEd0n46efroSJTkVKtBycVZDZ4fMZBy68fBkDlFDdhRg1oyKv+PnKyYVAHfkCK3s
PsY7Qll+7DiHSpmSnPk8wTxpF5KoIjst2InK6mgH38XA7vGsa1cWTMMU2JThLuSj
sQrHS/cRvMvKpTCtNb4cDDOmiLPZMDymSXesay+dSMgwxV6u4F6uPD/+PVJgYqMl
MVNYPa6PX1SQC2R919AnEESl7jgCch7kAxX0eXF3j1QbbLRdIT5Ri8nDELh17/ds
U1LnEiiJztxNzYKnWvaAZhIPEPypQZ4J80nPwHkad88fgAkjFCx4QAawyYhOocCC
pW/HKaz/dpm7iYklfY3c23E9VRtBiUV26Ccdk/fAmZC6kZ9Wc3BUeIPMQG6ua1jn
MgBrjeNW4FibJlz77c6X9JvWUn29Qr7wIFDO2wZTVax58xRFhqtT6t290E36G1YY
vYiQhC57plB5Z/ScKHOl1V6AQNbsDQouqgbhH0J9KRQMU4NPzKg5PvNmLkWgH4lk
RdpjkJLh5m5aIM7cDtXFb8IPSAdn29EPUdlzzMx1+dEaUbvqL5b21vS5ib/MDFzI
WjQBLkjXYeXZDlHrO4bSbrLrRMGhYzvHElrgVANrYAec47yB/xCOp73mpTDIoEl0
pWJOlL548asVaXy/tuP1vzWkRKCEssZf56ENnImYLDlt4s6bg3HhDBTaqU4cv5t/
kN8uygWxY/9mwa17tcMUBn2YEsbMG6Aou2CH4uwsp57BwOJjzEu2Ad73+E7EeQCg
kEvBjOAigZrcgLp87jvOM3SFHZ9bG08oqOCm4Ynx7YuASitPeKx617fk1tMUQwge
JoApWgh/1ehYSEbQZnzsRHk7dtWTMt7Up3AXZMwnOhGXE26whniSosXJOKGQcVOd
w0a0IyGwAiXnSse4S/LMBrnr1dcfIm33LHvU302eNHbFgMWkxgUuUc5HfMJSmFtI
IlwkE9L3P7TNltNb/mFfrUdIYrZXMmEvlE5LKWkPqkI0k2+Zw1wiK4eOViYk1G5y
iphC/h/8TTvvcQoobu8GiJrT8suMnuWOfUAxoMAJnteupuzw9HPunu1HtR+i+6sa
6494PHd5yhFRuc6OmZKmrTdyh95/LEcy0j9f/+GH1oKV28B430e1MohZOynGM6tx
8SYSkpu681er1ZQcgo64arQzHvQ3gHaCmjfhp5burrFwI7t5mf8uyHzBJgibLhah
ZNV77wG5jQb0F8jOrmYPhNTIr/FHIXJCTnEJwZITqs/o1FCu3jkD9D6I+K1rKt2E
g+Or4YDXFOzAQAcrMxF7CFc+M9wH3wCAvZdkKZihkZyJGn/dxrejyPWr4EqV69U0
zo7mjF2wM9fA3+LIMfmEcvXhvjzhZUL+pHg3tobVrH5e4fmdrtiC4YrOB8AxD1qy
KxzgRzUlzrlTNPxTRCFpyAu32QccZXTeZwEOKZFcjvkVkX8vUqaDRE0xpu3gEPgS
LdleNLgIxdBqabcAY1XMOibTUzTHiuUp765Qqv00oc7vVXzAlpyBLb8WD1WqeT8S
zCRCzYk2MoFabYVAojPevlKChB7uiN6Vym4dFooO9Qa6jeeV/JjlC5z5PsuvjBo+
jn6LpRgPnZmyWS/xDAN5SvFxKwnwOJDJ9perkpqDq+zVjrkiel8RCLGSPreVmxRu
3MyoiZcEw2LCezvY4hIxQxjtB8dJRAODfb+qqT+Y7od+4sTU6ixwbe9HrUxdKzwL
poTaAf9/v0wA5SFD/6eIHyvFo+tM/ulcI3c4zxnYxv/qVK3MRvbTR/dzbmqv+U3r
3AY7DdmtBaGlU48fRp3fQKrZJuMMLH5Hu28JcSFyS9ft0v30LrU314a/e8Ke3KE2
BnhzTPHDSITrG+v0N8wvZUXNJcf0RLIZgNWbtuwc7XXouRJ7p45ukPpIE5OoxDeK
+mhxzTPSRJu15dHkpTDVD8CyOUQWelg2fHAQO5Pi7gq1nY7hUNcU64rmpN1CT2pg
F3ZIxv0F+VvRSvG2kkogmvWfEEqIxP89EOKFrQzmpTgGFKR8t39ou0Rbxw2kYros
kQb63wb3PTEu1ReEzyfeM+kXpk4z9Hw4C90l9zQxRP3cRmrnxSBAsuzNThNkXbgq
5OBv91Y3vJb1OS8VfdQgGgq1YLKrQodYX2vL14h4cNXPpIorRlrSM9Jk2DNGp72B
EKl/xzmQW+FjPDT6zpPf0w==
`protect END_PROTECTED
