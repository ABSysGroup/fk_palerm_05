`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5vf3WE7DVOo1GyNTaBohdbWetn7ih9gpU6kaXatgEXvkxDgXHLD+iwYrLFWAVjEL
5u23vFZXu+xti2DkGxE4z5VfBB8XWEIeWzVdp/1zDyFH5azdlZAl9aPYjaBisLvk
hGT8XBmMHZFroPQ7o/NrpP0Kx3N02aQ00j96AB7FyYwQnGa5a5/sGcIfRkbfocFP
zlQkH2ZuR2a/HtNJibj6q39XRJ2mzWaqBL/Vf8kQsoA0mipTsVbSh6rwG3MmWhe2
A62A+Gicihx/Z1fLkAk0XVUMo2ylLgGC0r7YP1AeOx6WEf/332Dey3OEoS3dRrF+
xkC9o/uCjtQutMU09RrDyzZHy1nGsWh7rulA4eT6jepj3MCR+Pwk2UFpymmm4vyS
XJTSu7rFf9R7+xyNfURtuzXR39FqBFwjWf17KKUUOPXpsXZTkHoeO8ZHbDXxc4ja
Wp5eoepNLjC0kIkkzpBYCDyxqtdmrWZIChkPqQeuyvU=
`protect END_PROTECTED
