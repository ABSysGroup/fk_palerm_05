`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MTnsWHYyKuH+E1tnGVjaLqGgFRj3jgqsFSmRI7GPMx5muq75lImkRkL3ZsIL0r/O
EauwUzyKe8feLuIO2thdZC2ftCc3ja4R+UHvJtQloL6xn0diKvtj3sl7XliSkzlN
/ZTQFqbXshhJrPoNv7BSse0I5uERien9tTsnuyy0K8AxoYWwszJ6Rir9KmMjeE+g
t81fsZjhndjjk5sQpx/wPA3AOOmu71TYpdNRXJjPZHjEjn4cG4Kr8MmQhBQ6pwrt
V6A9HCRtWhSU0lFalZ+CpXRlCKR2+duELuXE/0GTXf6EnDq7rF29P2BOSaVYyS+8
/zMgUuJzxgZUNz0EWI22pUZLVe7B1LTaLjnv7lxPkbO6zQ58olqxLtPOuKd+2QY4
UNnKecIgiEeLZw7PLG12KP9JJ5rJh9Ym8dvPUkfNVZqniWZ/RBwJYwqIjVGYh9eL
bgwgoO2RRVCQQxXPXwRbZc/Z8Tc82lKnOaVZDyfLVYJKs0QhxVJg84NdRKOytZz7
8hUAjYH/l1KtcrViuS1PUwvs85ItwS4IPDpnRo3IDhsQ0u2UC/U9RGNcHUp41Ty5
hrs3hHw6+DyIdB0P44UrsH0lSjkpuBjZc5O7KpxrSNRyTuGci1zA31UYZTQhHtNy
DZOtSp9l+6tCh5GMtVci3/VjHkrMhdKeZ4sQgjU6zxhIgnd3k5Nugvxxh84RdHk7
WgvZX7c4Yvjjw4imUL8iyjRXWnRPzd3sQV7Q/X7yXWW3Nbb5rMBoBV4V6oycUCq9
8B5B1tFtEe9iOEujP+lSG4y8sFaqc8jjqcBVH6qkOzhmEQgXbke0qk3EorvQ2HCP
aybfkji9AbjlkKaDpJUS1BvTQI3qiS9iFcmO57VwFHshuXK6unXsvHVY6eBhnF1V
FvAt3YWOS8vpjFhVI1iK+cOdlM1EdbFEs3WeeIgcscgzSwaEIDpGsycUoM0JMiXd
8SXBdmkpVhrUzgvXlX62oSERkdjW81YH/Ozng7aqVZUcHEf1JINrOF7CLCTjzIYa
ks52tiWfJMf3LQxX1CP5sRDLwkVhGd3erHS1r1OjVjSoCSWquXwGMvDM/r0r2yEr
JUC+7hZ96SF3E5WW0WaU1+JyyN5uoWh3sSjd2shbdjhTOZkgCufbgkFnE1zUuoH3
73tBMas99MwkebnXdDT2NeCuTWoM29e+9cXH4RaSlXt2TBdAcGwNN8KFGnV3yAGv
2CRdg2tpbK5/uSfqMJ4zc1zh3u4sfNq5egFPn7BFGTSToupswhvQEYo/NTz1KlZE
0CxABFAvL9CHhTLFeN9+9WU55Xv3WcAUKw6le1yJWyAx6uZ8YTICCQJ1rKTWigZt
PUa8JMgXOchyPOELZ0CRMlVH0WyUjTNlSRVd8bYac7RL0wTzCv+0lgBPMb9/ts0+
EBpAhehy3cJPrjvqKcfamb+JviYEcJPChDzaiC0YkBpP7WqJO5SGtpQnTjRqaQwO
885l93Tz/muf1MuVccNSkLwwKdf2ALH4l7FEoNRTX1xJgP8j9HLfQOXUQ/WMn+yw
Ul+vUrV7WpJYoSk5D+llc2787HkXqg/qcUjg+JfOPRlWifhUTaLYKXXrWgTRmnhA
lX6U11Zfq0YaranAS6Y2IaHco6C7aTv++PdLvkEYJI0pL/KFTCQA5DyMG48M1eBr
BYC/4UH8u32MqD3lkTcScKpsP3gwC5pS7qp2EDkkNG9REXD3Fe8XfhjdsiVwmp0T
QkuguDJ50xGh59RLcD9fISrPBOBEVIuGWF/ThE3NUCTUUl1tIliZxcVn62uEpZa4
XtwZS4+H4AKBPqzxF4dtT/WVPgkBLhi7I6PSnUg6gnzf/s3d07a147cTpCJ92kgo
l4XKmuXw90nvHBJ6r4hgqSRpM0bkHY1605VybINkX/RlIsnggQPpJAWsgM3N8St+
wj2eAkbzTSP1WO8UzPBBQuekSnZ9OAr/ZTLvLUq0TacdkepsD/Cr0HBygj9mLeET
AYICG1po6hQnPzZjoIfFJbAZwnaw/BAtJdpaHoDQ/Fte7cGt64kkzPdUeoOOGnDp
hnv4/w2Uj6mWWdDRb9Fa6pAYzhxNBX+aRqJqMNyv2bfttx/y10JjixtjXsY/qugC
XA96dvWGrzWcPgq+d6Q/GUpr3tfaiOvckmscetgl0DyDxMWSj3GUv27VSIFoV9fQ
65sALFYmjkwjaJRmBt7pfXobENSexmie4dtPyrHKP6qckeI/WlmQW7sOQuhu/eOV
WnKjwTf/9ArLIx0EYIPts05/I3m+ndf1Pk0Nr/DGRQJr6ijDkpXwxYg1ZSJW9Bof
5MsaXuPBkRQngr694ZJL9c1BsBE1DrIz8/B7ZUjpKjgB7I1muqhoM0Y5V3liGH0/
ckovljGJWfTdumFct7V+q3Idfrvmu+Jw/6pos7p2ixMsBDefdi+LGj/2xa7J1SMB
`protect END_PROTECTED
