`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dwBgsVC0sARC5hR6TGl1YB5Bzop16yM5wS0U6nG+tXAj+usxo+9XG9r4B2Mzue+i
ZWE2w2XxJPTjjhztViOHKP2mKndL7SKSGzcHh5K+xICVJDQ+eOyEYW1BYVHrKJDg
qTtZiyQ3FCj2fuLE4x/i+a2QL/rljcMxlkQXgz99l9oMLiNJmKT80Y+GEtzjdxH+
9VbZFBeJzDQxlANcq4kBfMZBiSGDHkQ18h9bcDMhQwBbBXQxWX75/PZy4giAaAo+
5qmO9lh7booyB8vTunS99zMxrVJZbbjBVbzfOm2D1SNyaL5uThdzykJMCtQyXngH
G34gdt2/FRJbt/aIDDwjFusNIKiU0lZGkmhAttNflzJffq1pb7RLBhIxAqj4jSol
z40zwcQ1/wUtqJQ3f4/ud8QXksEqMOu8D34DoYnBYSkUnlOl6w/iRLrfWiqTj/MP
3M2XHI6J8cgIKaVluCjuOk2g6RyPcANrjVieJK9lv1o=
`protect END_PROTECTED
