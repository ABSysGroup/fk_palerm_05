`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
upJlVNfhP151XtGIOOwoVF+myWtAaYu7MyVN4Aotr0Sh9mAQVPtqHVmcRBrvRbGc
bk+/AQZUsoNLoZC+tCA4gSMLgSDV1yAagmxXRFVhzq+7XSdcebe4YpImM008EnI/
fApW5hZNVwlrqcjpiyFvQFMFkwhuwiKMhhuLHKlnvBKqLoH8cmlZsgrV34maVXeq
Pu5daQOFNkxPmeWKish2jlzdS9yQm/P0LxFJObaFcNp1PPNn007EJfHqYQ2gYZ60
mdAiqtFCFqIbsM2YLW3npXNCTd6Ip7/rkAZvfl6anZbWiN1BEc1yr963yfJ8okYA
mpQgxbFP+xneKuiuLI/l0YQyEMbv7FsdEPAgwv4og/BlPiyMiSqS2ies1WAnCeMc
qyCpBcQmVtP0aJb3BQ2Luy+9s/EV1BVbNtjU4NSH6iCn9iWgP5z5YsX06AG7Afty
AK2LyyV/tpGhKUe2gVAcqVP1hW3tH3ymNoiF6z/HTMSzttJFwb9biwLO7TX2CXVL
n5alM+084GEDw8ydP4Z+Wr7IBEJ2Z9UHOAGbTnUL6EZVEXe/2hlTm40VgfuTikd4
Az4+PzIXSVwsHJKPNmKt0WLWJX8eVZuLgrjkcqKjI8kehFbnax2ag2PlALiHoUrD
I/xzTi0Tuy18Ha5fhl6Sok9UbkDc1BM39otDNiByMzQVhu3eFsRoTVsE8balS14Q
s/D+xm3pDTuEwXDKSamXE/nlkI/YstHlDbceNrSLkPWcZbw6O/8+PS1oy5p5Mxf7
F/ziIvAmDNNOcjAjsc/qnqq4DLPPEvgSnov/A312VTSoywEMHy9r0a9W3KOuHW9m
IVMEMbaJL4vuttursmt1YcXqtnhhmjUo+2kcYg+LGbIp7v5MEZljYmrdDOmDuJe6
S6g62F6YwaLtXNrHLicZQ+emr3+501Dyxd1eKDJtzhVNEYz5JtXIY3TOFlHgKJIB
VeZck+NVuArOcFQ4kX6pcI2OVQdLRFUPHR3QwOUn2Ev14Kinw8gZ6xou0I4ziKsW
`protect END_PROTECTED
