`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GwjT6JbAZi98zoGWf4PUFLbrbfI8WfsSpMotRS0TwX31xSl3oxM28JMBlcOlZXWL
EKFQaP+Zupn5keZKc+XLvH1BNG3lWp3ZQZRAfrFpTdmLPJu6/MAPNdynMy7XW74H
MD0w5sh9z2A1SNdRvFlb6f6vWF1t8DaMplSpD+hnCrq22/B2MagRjhhra5xhPtWl
+YmgBX+XzTLrUoWPV2R4i1Xy7/AnwfFR1aAlTvw5QXpVJXYMUPdM0PeUQBB6SOYE
igl9ZZojDgauhIBrgUbkGEyBShpxmPJIUduukTSqDf5FtNP+s3ZnivFjfqtkKwPD
iPYEYx5YzNKGkJ1CatUZP6hoXko0tFdonyKLUuJVGO7vTCtWyRi23qAwpVdKfWoi
ufWBn+x4ADxY5h4+aRgg5WvG+uA+8b0UG+LQGV66KbEkCL0JNiyrZS9uS/9MzST/
`protect END_PROTECTED
