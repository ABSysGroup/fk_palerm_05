`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S0+uWTmx/NzBhRUVxYzp/U2p1jfWtv29Cyw0Z7n28oqD3JV7YIbY0StW72e1dzL2
A5GWhl4QzpX+RFTOGqwiVik4FjQmTLmgoodyvpyrTAO49CTSU2VyQbwtH9pPEaEI
jG/RH2WX/uOSi+B8Ku3OL5LDqWqImGcWfZpGIoKVsvoHX+986MmmtFoiNAlVa/yK
BhgOx+n0uW+pL5opVgZFTv1wo3dVByftale772IC1a8hUsTfALhM+7Uf4u/osSh0
vw4Czg9gUKnHob8QoxB6TJIvnUFEnaNMw0hztGZZ+sUITKZYfYPKxROprJXxxaiR
9RAhenUr2bvenwP1NlWIl0KHfVZg+YXuVddwsFyd8gq/YOIO7p/i/IDir5DcqIXo
+JvVIrzGUNgrwB7RqjsdbQL2iBJoOD6HUKGjUZCEuygOoUWJmu4FgzMPKNPLwZwT
eKyUG6eEFckH5mUh5J/9ONj4406qqqezNRo+K2fwxiX8MPOZbO8Fdm0VcJnOxRiR
KFYCj/ya8h1/d1WT/rz3HIliDOy6bQ1158x7tIsOFz6RFlZKD3Kaai6ZMUio551j
hYv8nHaK6dAMg+xF+l5yCLz1u+pFhuSoGY1CRUgT+P7ZX4eHj1N+SOjyL15BpHjs
UFHMIwGMqUocPcx3B5/YkI3TXZTeVjLtk8GPK64RYIWxX+znBrPL8L4guyIx2lQg
gMQTz5ZEkoO7JsIJ9v/bhBbaOEMF60RSCK1bBZ3N2elKQS4XEHkofUb/ahUTOJxI
bCZqKQihOG2lBI/RhTk3Nvi7jEBaKM0u/RVCkBZMF5EZ54HEjTu+GBfLcR5hupOE
NYMMGbVynRMhAyIxeYBeLUcPkbnc/KOA/0epGgNXMMhFk8QxsqxU/bw3nRpf7WDT
jTsQ7bCOg3fbMWv2pZyFewq6k2uEpY7gkJ52N8u98BUcsqHrZTaA3KwDfJ0PXmUJ
C6Iq7aXEal7YmsyXSJni3w==
`protect END_PROTECTED
