`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J1jhRFsQ2l6aw46q//DoScoTIePYsI/IVF99x/WpSBUXhXJDTq/oXdZBk/jMFR/1
54C3s/+F1qYpLjKWgZQdttr0PFQV0KPItb9YgLnsshNVMaUjiUifwhJlMoSCBbrc
hELKB/FW1Uq+f/mTVOYow1fTQ8gDqZxDHr/j13g42639stzFwlw8T/kghFfnX8yS
BvhjJNNDQ1XiHkQIWCn6x18Q16RLbC3t5BrEtGViQSUEWL2rF7olxWwsjua9kUAr
rbIu4GU9CYTxppygeDG0mw==
`protect END_PROTECTED
