`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nc857IdLmt9gxG49s9kjc5h69MaYuibC+DsKZ+ecLsNHoCXmrcY2mQBY1XGpIJMX
sDWr8e3RqsN1TZSBSxUO+bA1mOUZHsO5/H3E434z/62hRqlyDZ6tNl5a3eqiydQJ
weDWx65/yjKbthDQEo6GJjlkJb0GtVyw1zsJj3TVuDvEGbwGUQcWfDdCSllnt7eA
Kyr+TxvpjvZlpRG+VVH81RAzNddDSBvtgCX6+Yk6GzP9H+ScKMyFehC6IKrQPpse
zk2Z+e/74zM+YoqhXE6AqTVptCFK4uecZQft3AjTVnV1U/2ZwPEh0fHaK0FuF+Q1
iAWM3GsErNrHQz7t+KczLnqGq8UrnBZ9RfKGei43BN7NaFbYZ2dQiuXYJ4SrXX2j
lVHciTOrEKwIr3gs6z5SuKm5SeqhXq4xsDu06MEkKyO0wG6IspLb51Xtmfo1hGOZ
xs/A13/wVuY1PYe9vq2FN7Z+HjzGXR7v89XE3mJ9z76CFerXr+n3vke2gmexlVID
LCgChkeTyv3LnSvBGpU44tJA3slcG2l/GMxxLPK9p5b4Ygy84NY7oOoRlNSOQXyF
fHD6WxiUXGqgxox/IRrxTtDbcdLvggUxqid5iU8FMlc=
`protect END_PROTECTED
