`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CB8wFxYEbAKLgz/Ciz++p/iy1T9HoqAjkGMCWu5daof6b59u6sOoFOsZTQeeG8vo
Hbys0XRdUpM/vQhSjQ3P6wJ2kcapaZNB+eitXSN6bZi/fq1LnIY9On7sSVcgFMzs
TuxX2lMaD/FXEXcIX+4ZtnS0bF+bVbyvVFhhgqKuW6gfC/iFdwL5P/s81vEiU7X6
wPg8i8lyKEKosI7hrlc+U2QwYjWx7kNMRKc95KlUqIq6ODkKHuHpKtzrET1mjs0k
esTJvLYCoJLd5C4Ga+UJ6OzbVz/TdXDH+cfIc33K46Fs7+UDtv8i7oBD8A1SU62m
iwzYBgUCdymivos2p0+1I7nlm2KdzoWL6ZfxD0hw5abcyIV/t9BDmbPNjO6qCwMP
OPGqpq/mpPCrwwX+rNmmtJL3/ksE+zQBgrgvDK1vGPtSlmPhVhh/Vkgo5UMrmC0p
4UyPtu8IS1TLT0l03Yi5tGoxUUisGAaIXacrCxp5jqLohizLt+mJGOl+e+2odjMY
XZBE6YMO8cbnI/Fjv95I/wp2PsBiN+GUPPo/T6gRvLNY+XGjvH26rCOrpqAmDl5D
LwWt9n8/m4UY/3M7QLGZuXeBexLurLWdbXNIrziJ/gOX3K8S7viQK+iZ6NkV6b7G
NHHJdnOLtSsRIAeS5dOhkgFNp2Tt8dIViFM3sp63kBFXBaU9cDJyJCzhZ/PmrLVJ
U8ZVPvQxAyJsg42lcCVsNkiuTG9Cb7zuqSED1WKEgAt+QZNjTgLPdXroeAGo1oF7
SdHlzOQ06CHNyDuqHsUApjLtvUamS9FNkNjwHtcvt0gzhKbgzKvufCfeoxDLO6cY
188T6/a3qPQwYwkyBhYcvzAowOPw5Cjms+hV5LO/OhdV+aKyPVOBjqSJNt4WPHgd
YKN2WcCv4Yx7R9qvD7Qx6ipTfcJJ7UOi7j2xlVowW+VTrT/1A+jyRPAo2DMp55AQ
LQs9q3LFFqPj3V3MBs7ElTUxWTF4Qt78idHhnVUPLM2UfNmvtl9GDHrVaBnFJI1w
JsygAsLUUloLoCrWzQWWbSYPTX70rjIDQod4A3806jXRiCNFRfIgCgNRSL4+2f6T
NzpHPzP9c497hWFk8ki6g8KVRylqB0tz4pnhBXGEkKdm5KBn8Ll4vCsxkVf3Hzgz
7jiHW+Vpm1IGbOrvFSYS5iJFxHj+DkM6L2YyZQ2J2XkEBtJbi+C4S1a5lpRI2myT
RWSO8epOE4s3FASDQXWaCz8SrRL4tR0HBxNwTetS1ff0Fq3lmjO9lLfm7IdR7GBI
sVeTyYrgkFdhuTCDe/90VmJT6E4n17H/M+M0VZunr8GFAjRguzCpWu8dlPu2JZra
1691tJyxBQ4pW83+3vv5FM6tlb7TIP948vswQeLprkAikU3K5huZgPm7qJSF4P+Y
JTyBceNqk9Vzq5H120l3akVvcqPCeSXPmdPHKIOTH/DOAz0qzJjad0DpSch2bC6j
rmmjyeEX2aCOPB9LsHCjsFTZEKT0ueLwB57N3eXW0S0ZgvhcXZYJ6hKWC446nmxf
sMrnledBP7B8Q3/RHwoFI5+jrCqg4alQMyZPqlQYOPL16nz0DHhaeEHdPNflfFpU
FrfhXr1xefF27u4kkIqVKMJuAAysLXOjdVNQ2GJmfwxOZFvdTlsloIHIBnX17pPl
`protect END_PROTECTED
