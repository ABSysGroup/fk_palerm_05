`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h5F1FQi2kbWLM3sjPttYFzN0sLFb6WIijLzBBL+AbcvGmS25R9BgxqiQncaiBnz5
dugkUQAEOe6IVwigbpIT4Gk3XYpHKqHMbPod7uczfYBsH52NQGSz00aNCabFheot
b4T62bRFSnVC/9FmD8cNc8O2zelXtPI3vUoPtZhqhO95VH7RLILBhb46vfqWGCFz
1josGxf0UrjEnN1d6x4/z73Pge6aCwDT3bUPvoypO3VOYhNusGEE7WQ346y+gR/l
G4V+a/pw/swHtMSinuQBR3HSFYq0YvsnOPcULWAe9UqAssIrUejdryquqHORlDm7
Q4IO6TayWK/WCEEfTpvmJTJIDiyWNZhB/zRPAVStzhnP7sC5KjSwlZr61/4I+56+
5MKEsYPP/fBg1ehM3sL87sSecqgOH9KCMZBXRlHdG2hMxGMPmorbKRtJlDNJAmlu
YhzxekcQfDJNEoDYBJyB1WBtgIgiGVsxCG95r+pYmogrIRvA45bXsa9uG8ZVki/9
`protect END_PROTECTED
