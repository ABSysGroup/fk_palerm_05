`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gybdvfgI1cNNFmyyPNG+LR8H0IcrzfXWfutVNJmzilQ5omT4vn2Eo1xYCeiOnEwu
mzyukrtlSydiqU+/RDb3XAtKiAFFK3Y6Dj2qLfNJ6ftkoXvWqgehc+m4frb+6qxA
9sO0TS0lq7UXkXwQIxMw3xcM+SP1PyvzoKViTRogfglBPvktWjLGpmnMmANKCvsc
bLylurhS7/4MFgJt+ss8TDNJU/0eueV8Gc/Wbbwe7aR97vPTYnj+ZTwib4m6AWpU
erJDUJSu/GmDvHrFLY3fn/H1r87HZdkW7WI02+a9nYtjTisb4NyEEPUy5MFyqJGm
I0kmzJNx7um6qPe7FOhE4czpHJy3stFDuzY3k558m9J27HZsKavOY+Ij02zwEolz
/UAk5FD3eqdzuHnaKk2elua5GW2hWPDdXUJjs9495ItCDC+KHSPTetyydofMpxni
RqUPhWQrWX1nYeSckc68dg6AUq9CrSZTVCCCp+IcXMm7Q9YQb0daYYVDwkg2FZEX
4BoFmLS3defzOjVJ3kaD4VCtTkwea0ECUAynBoXTJacV1M+IVBJawLBz2BNgQsnf
irvV9nU84jimOACGCzLiqwASDIkIxgM41CDTF8tIE8w7lHnwOfhUHet8ISXHgZpx
9sRJHOPe8uCFd5c4BYBnekTVGcwF6Ju080nVHzPuWX16MLmFzuWjl1UVvFmP3u1p
08GvQVKa1BivfSskcEfBqiSsjA4S4qlEdsofNQkIMm1spVPfZNKnmOKLoiKTkpc0
IDhVj5hyaxSYCFW7Fz6yyz6Qli5r8pDubCkfcuuwGhLcUdI0InUGhQI+cciu4ZxI
yuBTOAKrc13kQ4gFGAEMUrgLJSk2XYJIdswlE6rNiavGf18Thv9BDbwM3c26CACS
r9F9KuU0WpozhsRYF7XzlnAW/me2E4aIfjCz60HjimQEThbghqPFjfthjPXd+wNy
w9llzzJeM1hFKcvXNFOJ1QRN7G5WQqeRWNX6p7aVF1Gc2NORuKCZcHCngu4cbfvh
3PGfnwqk4rUlCuaKyM0/6ukKoa8+djvDCPYO68bulm5/YoDkrl8vPhdX9/quByWo
8S2YlK3zNCZR61/hN13ji5sERoNuGuJeN3bLLhf+PV5fQ29gJQ/mnHmWxV8jWMl3
jJQWsLSpVVgfhhx4onHmIazG6LNHxwGKd/hKAz8jE+b4p1zTZ2KEyXEXIVLjzUaj
WZteOqpYCV1jKygHg28Zj6H4Fi3eQNUjRHJA0WLuqxDKMRP6DU4RBb+eBgHGFiRn
K+i5obn3ffGfpoSE/YY6fzZm9VtqKZIgQdSf2ne4+T5j8mjSqMxqHza0JF9ORVro
4wHy2EmeTz4YxkWc+3E2J0a2BdonOqISy0GfWTtImO7WigHSVmuMRaOIo0ilcND0
aovBIN/EJ7SHMY2GARkwdQ==
`protect END_PROTECTED
