`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hwSW692IlZZQdQ6iwYMcQ5wrBF+rkbqZGS5PUOYFdpmdvSjxlvyKWcCTimoAdIAP
n5kLygOCj3HvrH073GSgFB+Ii6+bH9gX0cZg40idfi+aWTZQuCsBJW5+1LLWESvf
DgYkzxk/KiIbRLvh+xE4+UmeFs8TlIUwnFydNX2bcWToZnrJsaYcapWhbSNWxNRX
xyGrrAQ3g7Cfn9iWN4qECPHVvQtnror/hUYBCz30hYpeNB94e2dmo89Lurz0Kdra
izXVf65wSojdrKJLbVrPYi0bIOlLamsI10+650DNmG+DwCsmZIh7pA4qNHpXCaqd
0+Xfod/IatOpqCkRxyCVF4YbCokHbBzMlWNWiHLX9mA2dIBGOKemwZ80J1Dhi/nC
ekPtIOy3lhYypfsbCsaM2HoMZQoUE3xr7g2RupehTh8=
`protect END_PROTECTED
