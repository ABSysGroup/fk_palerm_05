`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vB5gxeT6VCXaYikckO+LTRKloLyengKmfwh8x5rcQukC7oTyW+DHmDfnooXEgm6v
Upr357wXT4ncUrAKmbQSGAr/Ub8sn1g3CL0aSLy8An5gfP9KIzr0A0GAYqX/TkkA
U052fxkOM6xt7ZzdLBdlTGLibHZE6V8w8dx44rePxtQsAxUMNy2twhwN4VE2Y+qm
O7paNILiyXc1FTCq61uXfh8NbsZTONr3/sLPAJqVGSS27rDvudlgnQYITaW9sK6L
ufbim2PSP9V6SETF77cBuEQxnvNKDLXiv2sJnUkE6LjPslR8r3qNs211H72YBuyT
GYElV9Aa/qe+drYfjzcQeH+YBPiNaEopibgIP46vOmCLNI+SmJGkU/erWh2eCuKi
wgx8ZGIPa4+XdOydFPRSGn8wlvROMtWWDINWTAYaZLAx6/mGyjp6YOTaT+kPFrXa
F3OlyMrvogqQR1KTA6iMIJyiNDI9s/yAw9+kkgEjkLc=
`protect END_PROTECTED
