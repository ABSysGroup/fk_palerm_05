`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
za+aMijHHnOTN3g8IC4HWgsDpFTCl0QcrigZdCx2rzewbrJs0fWtlDG21X8AVN9t
Ja8fkUyUSdMB30H2cDQH6rqoz9O3fHWDmOYiGC+Un8wn1jhmAfX/YAmOo6G7cgIb
iADhPOtiwwRKHON187+N9+skbmh/0Z2A34XxvCEr266iF+mHLEpowS66dXSZBjme
ynKqqSeMF+sd4KyAHU0jDwE8xVnd6HQFLXAKHc72KofYFBglit6q1waf5+yrQeIg
UvkxIi0IcQry5oo1EmxmQhXB1+6lE09l6YXRSifoqcX6sNPhR+HvFhQoJcZjTkZg
FX2TygpsSL+fOfvswdCStuAfjy1wkn/PnsJPUZ/CxGPg7Kwbktx1Wf1KXWc/zoYZ
e8vndX6rJY1+Z4z/3yU5T6H1YNq89Zet8/6wmnLdKQ+sT9rOdhY2KJBGvn5apZbQ
giWyLv77hOep3bCaFyXFaXoSqu4Rbmm4ncI3FD0vDR9Y1TTQE31cBiQ62Jx2OhyS
8vIu3uSODG89hykQgksdThr+F9MZ/S4tEUOeuxs0BZOey1nwr4eZxjoFlr0naJPY
/i8H3k9QCbD+ST+g4jfJ1m23ifYqFucvhaeup90bJB4VmTz9zpTVys4qbcdAiLxW
zM4dURSt+7vgiH1rxRI5UgiC6zF/9b4dqtL3XCuCQ8scigbNAVqsJ38ki6+j31VK
cTPhLshPYZZgV8qpFTcBwRAhFss/qaDh4IPiupuqbcvrHUx0xeeJXXlqqQ/jfmgo
E9f0Q25zwqEPvz7do3ssAOkY4PfzgThaomuS5DW2TbTW/HI3ik9sR0rjmYWpYaBK
N9DVFcEq1EvzPEXs4Q+9mb6tAhar2hba3X0fV3IyFn6UXQ61yNkaopSmjhOsdUf6
0HFpHy3XYvynPLICcYfH07poFxbI9+kEEnfbjD7cQVPbi3qe1F3l4dLRSuh99WeY
anuh78QgWTRHAslxhBuji2AIzN1zlbqnEQk+MxC2JL6JqrG+iu3o9kQ3YrzYVUOd
C7d19IRmPJaGMLjfle7xUxLyDRah8ODb6wC54uzSu0AhANiS7yLf9LDssWtgAhV9
I+4ETUE+WKJM26/1Xe8nk2ITZ5VGynQwI4RX3uV9TsVCgtFCjW1xDBgMPYtWOYom
ozsWcIebWRfcYq2XkmBE4gq9BRtL/YzXvzG84heB208vBcGj0FyQeAzjqgZWDX1h
j5yxBYuM10s2d9YCnSJwKGE2ClAbbC1fMM4GRJDaoTezTr7ppCd7ySHkRp7Bpvcw
JSjRsc4Iv839knHwkcn6yTGdAw/Sx4pZNzyXYEPL5gedn8ds2C0lLACpBO8OWrhV
soS9TW2syqnM8TDOMDLuAueXHYlZvFeVDlOpZ40FH03mgn2/72gx+yVZvWxWK9PN
GEU3W4erhCIPfm8CuVwEURyqsO1xYV0/Q4B3VBQIxQD5ymQX6f+InpJtNlfQowS5
al4flTUt0SJb9uuJ+dOsHaLiuhpKQvnvpeCuTmwEfyrqmMfcNq0tsu+Rdz9breSn
dIhc4Y3xEIBuvcUp0uqSGWWa4qhBCqESncPPMe6wHkflKEx8/DQKfERbR7gCkRgl
oRiDcbktrQR+b+/lZJR+LWb/TKzSFkF/eB1IPzbAolKpT5P3S8lO3LufW4u12SwD
5ckobl73OjEsuuMBm1+LudO41gjNDLwBPCtC2LPZB29QRftQxV93QgjrhKTVhYjo
IYD83bkqvbvmYvOPRYYEGHAMIXg74mrnOBsByqtERbSLrrA+UwFhquVlZWJgse19
q3js7qBGuOIlrYY1FdP7e150HaV7Mcbja6HnOLfP7ood0scLop8/RMmiyBLCmIVU
IAYRThhLiY4LUjLxGh7asCYgNL3BRbCIInxVTMHR7EN7G4Xs7mCkwMssrm0SkQxS
ZkYerzxCVm9DPhPLQzX56xw0/5uFXBKiD8AmcPymKdTkEanqb0Jo3R31i+UfMbA3
HaqJMf55sTLA5KarhfSRaeKic+kfta/e5lTMU2Vn5iRjMRyzxmKzUqpGWclqi3bu
ZHIc+2PrpdgOKVikWtZVJ9VlQv/SKWAhXMO75ATUkgEfUnTenO+KWs35jdLNiKul
c+9K+UDwx0d+VH0SlPLYAQ6k47fSPx3cO18FGWOxFXeD4wsv7X2NOOL0b+Cz8bjS
rrs0DNFxptYi4ShcujFfK/yRbF+TIUOp2Kt5LFr9IZIpncmsAooqchu5EJSE2wxJ
0CD1MbOwcgP6EA1z7J8qHwneXgbt3ouSD8YxSQ+iPkg=
`protect END_PROTECTED
