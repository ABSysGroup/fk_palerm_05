`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AD5L07x2XnSK8Ri0s/cGUIPiQHc0JEG+QS6l+Pm7uswSOkg1CMJDWu8oo35khAqj
FF9yZ+ulQ08RmzYHppecP7HduWTRj4pY/AHKCFKnIYYviB70Xd1GJ6xWf2m3HSh4
8SGiecWfXzgTdOyZBeFuNr3TJawqhHHW6BpmpvM0r9FpztS7KsQ3NEUnQiwu0VH+
At0i5z4WhRgX7qMmkoY+02EFrNmVMcYPXx8j/uGklrk1PrdukXK5xR7thG904ymz
/6kXcWlvdVqBvo2u0KUN71Z9Eoei/NXg98hcccO7t7C2GCF0lf1sCVPmPjCPfMiM
BYirjAXqrNEv1M7MvhiAPGYHO9N+uD1miz0GnP8eWTMltg3JENBK5iI4qDgNfHPP
k+NW8neJei2jg4n2qNZ1O0wG1wKPjde3TL31/buWAiQXb9rTPUptncpHfn7Up7wp
BMeZDxIBp1mo0fGDWFcggYYJ4WTqLVLCtZWtZDw834XimWdqShhdEOh/jkLlHPTU
PrRM85EABVUddLuhnRJQb0+ZDHFfFv2MgPrpymOJ/xlVq6i96t5EkvCvx1JeEBDe
BM/Mu0SzEPlCFJ3YHjYL6t2vE45CGgLlUHmyPC0SbvydNEM+bcsrUYPJpDft/XJH
`protect END_PROTECTED
