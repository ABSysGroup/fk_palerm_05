`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LJRiSzbwNBClUv4Gei9CLCHaIDJ9Zdw89O5LDoAJeezQsQPTh2lt5x98rtipXdsw
ARvCedQX5/Bks714d3PBwO2PC/P0k+Fgn0qHoSuAE+lGAE8zL//epiJ8QGSoFS2p
D9JASUy/UvSkL/XwkfPL5X8NAU/IBbSoVckQ/zaBXrTVG6dkJbiCRz+lanyXTwxU
E2FOHmreVjWzjTVg5YaAbW7EWzrnclfn+gMKZna93bHkW/IDj+//vn9l7KrQf1eg
t843hs1JrPWJvoKNg9WCk6G/G52WHF8a+ZCIFiU2BkfpHm8SufLEm2hQ734ldArU
BzOKD5sP3GM99TJ3CxpSYQmOy+vfHJh2Gz/bdoSZHLo+LWrBnDc44QvuHaj31hiE
PBLAIzXbNOHaZx+e48d+lMYwZ36UcvzeiJt/xgIN8S78j1Kb1FiAU520vFnfrwZM
qKzLsP5O+PmDkHdlyHB4B++DZm6U7a/XmooRcDCcLlX8fNIln6q8SQj9BtN9m2SQ
3xJKjwKSkS+wAOczJtnNcUEggSqq+ce5rQpGrSDLbjhEcoVOLPc3NMs18V5/OXbu
tBZ+tlGUuShlUVAYAamyogWI5Ik5FGy9l4BDs5h9/eXQ5qMbuzlQ0dA0RBJVJaQj
MoFVgsg6dVmLnDcfNoz/9RcXTcG0ve8XOe0z2y0GsiQrTglHggajZZIyD/Y9juVZ
`protect END_PROTECTED
