`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DTe8BVganiTFNKJJGVXQSruVOVHMzHxyIf169Bm3BZef3OLfWJlnAotTJZAX7Q5i
eqbY8AuAKtA385uVH+TtodNZkYF2zo8lqYTOgKn2kwYp7F0TJV3jPGtVzmwm0BJY
087fjxNFtxzp/Fu9I1Kjj4wMondp0QeUY/UouvaFo7uiA0bEHIe+fU3kXjmKaLch
CEFFdvOB5bwFZ+86UrSbruvAW1NNSWnH/M2WZpW2nzsIpXarTp+zI+BTYmt43Gz7
/85qMU6g1CaRKprxHciRjQ==
`protect END_PROTECTED
