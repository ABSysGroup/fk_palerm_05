`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NCU6R1Muf0UwyAvHOQ6hDSWEcymbZDqhJJ6IkwnO37PPAkEkPo8t61SkFinn2FlV
YYL5uVbYVZwQhWr5XjqwPCWVTru+oqxCrQK1HFd6xy4PDb7qOm1Pd2CILVeL4Cyk
a/xE0qi9k75VAoVyI2Ytuqq6pQsOxQA3wdLwv0RlbBmsBC6g9Vj6fWNs9IPkkUCw
5YpIZwgli+q6idLQ6nAybAa9F0JATiXSoL6suYa4IwsouL2yO94dW/GmL+J9LvIM
qPkJXUCUL9VCdYesD1NfxDkhgmyzFis0ENOlH8nXNrV6u45HEEbN7OnD/A7kS6Dy
kKFysU5hmrBIvffxkUBRhGNsJW64aq+tnmzqIAogdgcfFt2HWOhUwFsmS8pyfzdE
ORZylMeK7TnbAYl3oVJIF05zHV/4EfaSZPOjBfxmVCZg7O69854xjHsQbcyAxznn
6RIHn+pyhjW/bfgIzlWc9gkZ80caxvtKIZCIcH1bVbKYIGF9ehlqVSbGYf4U2Z9H
8CEPOg9OtzhlNF2P3LujV0GxhEcxkrVHf+aFEbUEoaWJi92/DkHaoobIKN3BIvkM
HrrbQHnnUt8naU53uKmXSwsc4P2nMp0kXahNVrrYs0HaaDOI3mUK3vvyJhLc0QL0
iihFGuCJFXH27VBp1b6hvq8aeU6eyqmoartWCpprOnagvhP/tzqMzVb9UnQKnCkG
xrXedTo+JUseaNTIEV0qODICKDcpNQzT00nE20D4diyVtS9YZasf6bRD82ioj4cB
2v9uLuvelZY2OmYmQeyG3w==
`protect END_PROTECTED
