`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iitebjKunHdBBXLABQWVMhPTkMzcRRAiIFWAJieUVOYpXZscWdApJVORh+pQW5oz
1bRdsafa4DsmRHPYPtb5ptO/gxk1k5xpKJsLBhtTlqRCGhAN5Q3BT8I+Hg8BAW0X
LzdB37bYMmpIs61uGSsYD0U8T6lDC26RCIXchBpsPtJRPU79dSiwfdb0K/KL6k4V
/2jr2bb9wXZO5p3Ococs3iY/d/Xiv+xRnc3Rbr900D7T5B2P0UacQ9Off4twjieg
R+8yEtS8DEEnc+BlFg2LrUzaDTJITGsX79fylYRp1IE4+ff2WgHp0r1hm9+N28wl
q3wrA+gqCS+7k5vrMYdXxsr3JkaApao7ACipsl9K298/XK7LBpKlZ6NrgOMR6bmP
0U4lmOOshiWDQtRTZtWErnehmleQwiC1E+GrW0gqoOITPL5lNtvJRphxmxir5p8m
DLmqIqXqXe+1PGD8adQBMqoqcXe5Utb0xxlMynpUnBIZVibPHEA2YmP4v34Nh/gO
jJwzSBuZQa33mUKBgaQqt5ud0TC5ouj30y8dd7NvRsYlwNMFpb4hltgG23wsvaxp
KIa4lnHgwhILjuwRaqMcmJEkO+mxyCMT5qE9uE1wTEaFCfTqAhYPwGmB9rjK/tJS
fGuUsVTXEkIib/GfcAGFKUBeVsHmwJXWhvkCBHxZnTsuRKDoEh+IIgyKcbotPXDU
HboFQL7SfITP2JBUdjEjEUNYHfi76dfROa+xjfF8VKT+4LiLqYJKEp7nqwLTVIgk
Cf7wG8H5FSXfVgRCn6EDGgLgzPSjUESTQ7NnlNO7ptO2dXOaAzboby11L9Ev7BXv
kO6ori0wzW7QNM1AaX2fxm1sIlNppuKF3D2umEM9YD2A8tC60a044LPvrHLH0Jvg
sSfXNyiPa1Jg2YtmLu8JNuELsp5uGtOmWeWAfC+5PkIgx/oaQPsmYQiCfZyDZTAt
8tWGF+td9DR9HCrsu+p8evq1R1Qy99uNTwyCO1ersmm3+/OL619f4kDK488PzaFm
YfEwAipAObG8T9CLzWUknkw7lGkE0ZylIxiBYATfF6hk9sAuzyYwbCE0hWGV3+cY
WVcZHA+gGuSQOkB4iUFjdWyUYGarzkB8MsVZ5m7WXwXnbRJSEKC9dLR5Rn0vBgR5
SAHhKu7XEBa2LnwXf5+CbpJvKvKaorlf1JNNyHInn+79S/gSqrvAZw+NPv5LLPs1
P9d23XW8ahlfpswGqSmRYjR7ZWPExoLUITycOGF8BQy6s6NjsFkGvOvcpIIqFU/F
mXh/RpM7DZYpd1yuYj1PuwBikcBoFdj2dAklVLdS8oHaWeqOp6fFT5E7oxpxJWFG
iJ9vQ4hW2F5Anet4ZzMIdFPz1eBJJ7B52Hq2DWGL82XpFzMBQF59YDUglmLi1P31
hkcbQQxA3M7RPO6Hck414zuctrakiQcdglDpWQ7En7DNnt7JWhDkVfDTflFlogLm
It9e4xZNH8g1ds7+RQoBq7F9LUHpKLf5z9niv/3i9dOqCenT/pi+E0KYXlbBloaJ
C1cMeCxpu3xHro2OaQen9+iAx/LvlZHGYqWPuwCeMAiWkvKGl0JfMbznaMeQWRNJ
RJk4rQeDXJZk6URw4EF/UZpvRaFLKemJ/lajlEQpZmveM+306G5H1AUoF2nRGfXh
HOWXxz4IPzhkajr11PDlp+c6PGwY5wfWYx8QTsuY4CRSMxGLzeMNSKgqn4LWDymM
F30emL5qzbyCa5/stlOdjhh/jou60HfpASywAKdeIdl9Ru1rZR4k352sGDeNX61+
EIJMAhCj7rPYBKxHKCKvaI8fR0hAViuAPeXhEzEHCy6OcOz52eYw+rDULqrM6Dgn
5dvtAlP8OT3jF9DFYNrWNwc0fEj1v257q2j2UJ4nWkM/W2up7djUjxidq41UfCNX
GCIInvLOmcxYw6NCkjBYjtjdUNUHDh79MNfFGhCyU/OkpLPrgojJNPqO3zfwyLR+
lQl0f17ZFVkxKxbBXkcEsSblc96p5BJwaM0JhsiN2ZfRR7xsei0Jc6al/Ftc1A8J
QMxWaXRzuku+FEgJCCmD78ipk6Fnop13Bt+jTF7FQ/AJe7I8SWzBsG+9Hl0ov/dw
8vFkTE3rLx7f/pHL9nZ97tzqlB4nAT1bLDOFCf0xy/etcK00nBKlb9apiE8bIOHI
4h5YBzfxsuzIUwbvYxyrtBuS5bH4BQn5X80rUbTgUr9+bpif2JFZ4wRW66lWcLkG
DnZIhvcj0pVvsAnPTkNgcW2uhlLEM5VKno/fA6oaAmOybZavh8hDqHQm9VAJP7Yk
HCZxjnVR215T+NPl2zvGvUKSoC6lqQJFERE7hYYIsB0v2E2yPa83cJLzOqFHUIob
l7C+7Xz7OEaW/cK2P4yQNioMcvt7xX5aJPoywptdvyo7mbpSEE3QhgoZPlAHE8ru
OCuW1qbfQsOB9vlVqOZLDaOQGzRNBvQ1mtRAsa2nFx91fVKsGZvegYG94zi8bxC7
EPkeRH9DsPmMJcGcRmIH3lHcckcg9K0xU7YFNgGAaZvFQrnP244Ma7dKw6uXhQqx
uw7avsWRyC0yjV87oI0KvVFz3JapDeZbjHRCLBWgzIKO+vTHG++p+KAhO65LTR4C
t1OX3x6uHb8nc5tdfSAhA8DcPQWQJ6hoAq1VTqD/vM0y8mD8TXA8zlD8hqyegDwP
Fg/hxSYIRjwAKVMnzFaUvqhTVYRFJf34DXJLLP9lXKSc8geDsIZLTvnrGYBVtwiu
W2avP3tOJ2witYaiEEN3jYYN1NkPOJJkVAfDR5S5afxfTlYzrop6niGb3wf1i0AX
m7q8FMfppeNdHO4aO6lmRBW6ktYc5IEzs2LiFV3ud3nstGSqZjbQ9rex8IF4QWhp
34/n4qYqkg4+SizeiELQM/vzUdOXyVdHhs7e/HNS43FoVhbEKT4zzP7rWPAXJA9D
TYFOK+u13m75gnmoJJSaS1Ec3IVOvfMxD6KgkctdddTcbR40cl1sMY0T2iRVuEmK
l4zOwPC4zXfNexvJjH1ocvSLtqVysdXsEE8IraoNWPWg6qaMuDHBvafYsUiltZ1s
wvGnInFSqf85yLKLCEdctL0Ubm+4DRFBT2eZzmYSbtzqSVYv7Xg/6A3vyn9XVcYG
ceTU1g7pQkHHnGzQC6CSZgDP/m5bm5TdY4ro/J/2FR85eGYZPGFIkCaIgaUeRm01
OyqVrXU6VO2gCXLVRebL3Ilt+sZIqQMQ+UzHlLI5/CRiKyo/bOCVpmsgC+tAANvR
O/MMcoTnn5ET831ZxLOKqaiYefZtelDvF71MWtcDJ/LGa0id5+cPSfV3k/iXvNBr
fY6rRjJBuU7mojrYxa6gzaeB51qWhFH0H45TUahJTrk/ElswY++Hzzb2qCLyB17N
ra9krXjsIXEZfb/RoFRTFs9vGg0+6UaAcpjo1oJj2a5JFCOq4l7fACfeBVgvPh5C
qgK+R34InxhTa7WHD+ybiR3JWZDU2tGonZ8xyjpXccA0wUB8UFQ/ep3W6B88DxEw
GB7RucqrUCj8LOE+i6Fi/hMtYIgMGZiaY8v8pgYgYS5HdF3PzDPqKQcufydW9+8u
Vg0vUehcXOn3FhSvhoNIRt4hejY5OkckOlsmeUPBmZ50J2HfHtaxfqeqVI7jvK5h
rxZ/Cv4+UYDg/5TDzTDjEkTqQ9AHQmYdaacnFpIlOOrrTFlQlUGicbmC5s1AOw1S
R0c/M/06N/VImQ15B+I0cwFphEiQtHS4ZQtu52lHiwN8ixm/T0iOxFhVT+xTWwxN
1EkKqDK/dYeNWvs2Y4ReD7tWPP5IfvteJNe1GB5xIzFgeXOFZWbuETofQ2lcEEoO
DA9mm4P7slSGRJWMpkkJ1EDflL+033jo/uEIoRFg8ksI8nHOZAy8hYO2PWsJZJLF
MOh72ZPlzm/sVc70YHWA8Sy+GSyvhZd8yMix435FBQ44PY0wIiMo2H81vuNm/t9R
y4c6hFh4aV+aZ4J1zkoVVMVUxSeKO135+GBCtd2+1g4/kTxjkvFFLwZ6yhl95VUf
o1plEVnn1Krx2+b1DDnjbvW/hVBrqNKIS4tVaNzEegak2J21MRKDuduCjuulInwE
fA+tuTjRLuntNcd/BuB/eJLeummcQFXy3EPq+o8A7vbuVKrXCP2N96ZK/asSLs6a
oJajrb7TQPRbCQCjrdn7woiKsfq5NDBX/5avwBZrU9c521i1vIoCXgxkH/lQK7nc
Ucctc4JJiRV9UfkBVCzBzjFDx89knD18Cej0E1MMoNW4kgAhMncaO4daNAski63W
E6/XNqhgHKfB0ypHClIi40R7VL63DKcgWWC1WSYRiLAmbrMsiVb6nigTLkFmdfMe
bkknG54NO5ZESbLARIXziEXTAPpDaU7HivmqbgRzyi47kXmRiY5GE3zSikj/W2XV
0JpDQmoQ4bhHOB9XS4FrDvvr90RBxTEXBnQClzsgGcdl4HdR3zs2gJITFK2+ffs6
7MA/edMTYYDEDPVF85aGcwYspIWo26ibXSJZfQ3USajOIh/Ke8LvfJB/VOcudVvu
yzOMC6zpthnnO/6eKcoOxze8NSxBgdr5abzwlAdAHq3mzHZJl98jsgKuIIalNn1t
5D3DCS2g73vUzrt+9H/RbxP8OESNHWoy1yyudqiJrvgXx/uhJ5hDYGa5YsC1Ox8W
Rlae825BIn84jfdTPPLx/xHRN3nsVn/bpt+/AGf3TiF4/lVwNnx91EBA9UY4UtOV
PLWmyQYlXPKLo4ejIXzXskgP36l82BDMGQW5J3FzlgWEry7zreE9cXeEg0HZYGHJ
nZOzvn4z5KgyUbVnE9JQFcTEmyR7HWRSUjkJLdqjMnKd3uNvYa2fHiz8hYHz2c9V
pDyt2D2LHK5BH4U2qMKqfi5aAeK2i5u2r85kPVa5EuCng8HP/QphnytYK5km9YLj
W4N2lhi5wNYsXuSHB//0UFgwTRruOXiTI4+xhM75wT1m6hbqDd2PMgY+69Sk+vIX
qpnuxKROcmDd/DndELO564LUQnlfw0z8N8+F37ONXjTOHlhd7qkwu+c2WNe/0v38
JA+aRWmMhSkBuY0gIYe2cyFh/B/VX+hZnS4LYzPxB9I3+9PGkjRMCYa6mZgt/Dwc
Pf2O3yjLEfRfXyoS/zpAW42b0sF9FrqOETvFtX9rDRIPHRBy+PELLDIxcvSlAR37
jvkZPelSarvUo0T9PkQPt/Qkc6zkw+RVXU166etlAplrcq0EqXz8d7O55xQr8bOy
8cP9Y8hJTuZkW5fjdiubjTQLYBMJQUImNdIotQCi2yLPQPGSGZYinJ44KnMSkhnv
FeiSkaVnqz3qxFm4EVTAQzGUyw4YXhQSx3gfZ+6Lis8AvNbY4T5hsqZT+IKVZ2i0
lzVGy4RyoCPcKp85tVorK3hHKDhXpmoPmNWembB/SlfJiXejhWYXwY5+q10ARCII
yX0V4kDauJzjIp1NuS0j7GyS+hbBU3yPGWF09DEaVkeMfNxUb38N392j4EAN+4k+
T7qYhZM4mWR4irrgPbEhzK0qIRLvoPJtNHzFjVrMuroDDfP1dDG8pulf/roHxl6i
aaAEuA+gnCB8Y4C4m4SdRQUVZ1CSkPanxAnsy0GbB3cWNU2xAy5yRyDAXaIr4O/m
QeSM9o5mp1SFyqNKi5DAqhAWFalY+zhCo+NvpqA2ssF4VZhYi4z53enafcIQX2Q7
SkqorQAj05yi5Cm+6p/pCCC7z4jrBgS28DQ0DI7HdfgPvivvib6NQ4z3y+zLF6mC
LYVd1BiOXey9Y7s1pYWUVCQXao8dW13RFT28gZzD7EgP8GeUfcq0GZ+lWgnVSB/a
wHEWjOATDKwIJQ6ztl4IsorJEJfBMRK0K/Z/TZfkdzLLdRkaAnd0LC+zdt0ASzp2
1rQCRoybqq7S5VtnTrSz1U4Fsf0PTsqTxEDFCOxspSp5WFbrFEkLVkYhjYMFxNaM
5CCjKNky7WPiDu5bvjabbiLADG9ywVrnPJLx7iUcI+S+lFBDaHQ0s3YAemise9Z9
Rm3bNBw/We/rxsfY/I2DnHCpmgSkKgtmjjyQIXRHjcMRqGX6bELbW6bH3YcieBZ2
Gg2w0f/ceoVtG1hldBEggJa2FQEBDuqwOYkWdfgvqUI0cNmUYfNP2Suz5XjptqYE
UJqwQl0TgPdlxLVCrYLXU+ng5yFMCk4//UaZesOQQyYuxdICuufEOP844fAJxRx4
/bhWtcYq3LuNHc8hNQ3vYIhNRw5vriKPwamSr7znf1nUg9NknSbRjSy8c3nCCB27
XJJNpicpo9tNWVg/GH7vQMDtLAuFD45nKJn1zlZdrlLRnyC8xHnn4z76d2INXWxR
hnhL7/WPqCcspHCcMxGBdFbO5pDPUknvXHop8HmcpuIQyjzsCwYptim1UCaR2uP/
h78e2iY/wDhZ6Xf1CNYeoK1NnkTmsTK+4AD82k3ZCaeF6CA7Z+ccEtIi6SaKwi/o
EnzRNnckC2G2eDGTczkpyMpCNdFHizoCqFRhyPpkBjcFyma47tYqpHDY1jlmFrsC
wJznndhtTys5h+/bWXFYSb4Lx+3n9e+nkKvI+hXTy2zfq7GfeVTChxzZJ4SBpoxV
lUN9oUWVljfi/x8SY1n9d4QebnXrnhh6jzjlCAiMKUajzOGgFKH8fwekHWPW3b88
jHCxFOwijr51/D+DrGP0s63MCP1kBc3fMCYHW+PWFr6cOLC0rbiobWNbAWgkGC60
NmITN3lG9ZMvqRFDKV6NaYyM68yLO+FNnvdOy53dGSay7cfFZ9q41WjHz8mjKii2
ExibsFa8vUk4qptrTwMIx3iThSA25HltRYS1VCywUHWT+i7LKtzGAGWc+16uAgLs
xBMfjru+fEYozSizflzKGYnc8gH+DAqpGnflGWZz7GfOI2V4EDTQF72a61aqnTS7
VnjwUF1QYYKeagOZ2ilLkrJhtwAcJJsc3+jJsmaIJOP00SpcKzwPD6+7yj85Yh7o
J74Y9SeQv1aQVEQwson/+WkfXZx+Ex1lt0b+9OVUDN8I+b7/qr/VhLZmajPU6z7g
8ZUU1q82bN6hJLNDzq2Emf4XtA4dwqqGUn0AEYpeQ4TmEapQBVksHZzdqPJw4baa
FU0u68Si4IahvC7ryBOXqhf3ZZ0hveUNhYK/foCA48yaMtEdN73mMMc0QyFqhgM+
zpyXtTLg/KBEX4zJ082axi7jc7wU94PEE0yRJWRGVrl+D41Ej2zfCU2T7K8AbRwQ
PpnAQHEfGVHNsJnzQHEB2ksxwhSGYBXB4SlQbh8FH7xQTt2PYK7GKbTpATy4b0ML
RUanocpxOgPCM1eVi14fkz9EnUw8ktbBq46V/vHZrqq6r5mktfmlLd6wyYq/kgji
ATwDha6wO/Cqye7bM8B83an8JQex/u39dn+iX/sNu6UB1PK9JMxu7SOH8gUhESZk
OtfmHzI174gE3Qj63P0/m28rnHaQx38Qw64gqRZLdNg8S607N6fwAnPrBNbmtIGb
o4VyqYqdtWMSxVFNT8iPyY81qumkb8YFldTyxhr3vdQ7cenLqHdJvM0uhUTcfOQF
r0Z3kK4hDPUL4h4eDx86LZaUlxGM70gfyfM+jw2S9mZgOJsRjWh2k5TYtnTW72rs
jlcabC6RlVpLQs4rXuhO4M2EBgB7elldR5d9MJPxqdXbAVYPMSFuUMYvWEHdGLgH
JYHSr7EraEU1m+DndH9H/SZRdyrpdJ2RyXtunGgxfhg5zc1fFW82DpMO9UPcSc2m
Jo9pq2EputINbHxkTpZdRz77gWIQoPm6KMHXpd3y1iqNY6/1k/NvtPy4W9ee81D3
1QGk9pwbwC/kr3sspszwNyDOzPUsMwWmrVDrl30OvwP0ec2ojhcIWzAsSzOROUsf
HBtatRUej4sL9rWCY1tVZNIjbDs7VksD57EpBltplIQZWXGlVppz26rQWuKOfgnA
tzM5r4Ysmv1k0QzG+dzp22vizGWlqo4GM+u/ekntMIVFEXBRh12L2ZAHS0e5udBk
uAIzOblQEBgA6K1nL5My2haBP2eGQYBVBQ1hFKBjl5XjF88N1hZ5LfvQrUDzLCC1
bvlnGZ947XcxvzVMMqL4qxufKkqfdeBh5avnsckgsroOYESoMPDj+Ez6i0J1nsho
NhODOTxGU4sd+XbMoc1/44XK9Ml3rAlsB451PgrC5kJ+D7lEP/uUhky4TE1Xs4U/
2njdue6Ble3zZ8EaqKlAroc1j4WgwmB+4itJvQH0Tn0YCOMMSGn+XwtviVympb+y
m7/klJBrH+6/pYU56IPR9BNWAkWcWCAU0ckoK8ibHtDkz35I8VbtfFP1gg5UaVdl
RCIyFxeplUnRyAYvJzWO1bhhCE2AASddiOnYe80kLMPMS8ewiCfGtlLiLlt+y+aF
ApGQTTdtuqsxbuAgrHel55luJP4OBL5vIBvhZQ/aL0L43rDHOok9bOHfyqnxiPUC
TJ0ZXNp8sMPKfCmkO2UfxHCIEs3IB9Jq+pqs8sXkjKeeejFOM3kT2a3Dr2d0LOnT
bkfQrIQQQxDKQ92OfCz/du6W23CLIE5bK0V3J2W6LgU+WfYvdynOkeSffTxTx4iT
GZ4lQkveMLZgl03IYcqYhFlyfBhMXyFpO+XoZcnpp6LpX+eapJp1PvRldlbBHWwk
Aq2qbCJxrT2GZvT7PRikeSESykwgrxjhQWqPX7fkD+sNLLJbE0XnkUcaHoe0Nl0T
EUr3s3YLpFThPDPBlLruc65d/Xc2SxLo5bbzHvBQVPlFq9m5J4zoJhhoE8NmpOs5
ayOMX/x5rzK5F4v1eKBH6z1bNyDKe8yY+3rRVLFLVagv92fNgPtMYmmZZD6XwjE5
2UUslgbaf/+9Y6UBudjkQ5c2iOpZgdtJkSbPTQ5N78BtYE40vYBUkjH4iYSHbx8w
bcYJSJ0oDlawXniVe/1WRoXho36efRX2PrsLj1yj793FL6iAqdPKVjnUEHg96FOK
eyDMFJqmgZEUe0dFhoEeeHpnovAZrvyCBsmaacSNSHOJlxZn4Fl9fskDS1Pz1eQk
G7dCtfLkRZM4KOQXXzja3UxTu2c2qU8vFDBO4uO6T8KI1r2gvy+/y8mrO/xA5EH8
g15lv4wIcI+j2MVH+taiVZZvyZ5wWRRZpQYY/My66Lblwhen4edX4pFd53ZgeVB7
j6utJfmt+yQ3Bfrg9rMjRlstDPvFeVKgagfeVlfTEIJ1i8ImWAhWxjMSohWa4Gad
IK3+yoRSCGBHerQ/+KQDfnpYW0Y5U+Gt8JlVgopbuuAKdDzBHUuyqXKF6fnagwpc
4UaL5+5l/sXKigDfLJWfs4tRycGgdq4oOmef7WrNc+jgoUYI3SXy40FDgGBY+6Dy
n7oA6oOZafBnF6utTol+0IgpBzyP2dMDMj3xqe/lumTvRerm0YuwOZdnEcuJSV2Y
bmZHJLIXaR2V6E9o2hnZU4iNkLnWZQ5TT8H8RJQsie23OzPqeW48DJA1M/LKO0mY
WezVC46L+95RADNSvECxy4kPBeCzWjvBdz1nn/1obZ4+J6RqPT+h7dPxpv1qrN2N
ln92All0N9KY6e1c2S7iQ52gUTb+CdQnoqkyQKxMfjZqBOOTqODQzaP3TAnzql9R
ZvdB2khkl9Av39mDnl1RET0ZnbkZHiQ75BjmKl5WnbwK457ANTeQxRvHDdKQnqNR
lGxrz4ZHEg/EZIXFe1p60CYaYSjy7MaACMVX9TCT+hHZ1R8i0/NqkSDafyCnDCUf
GSFn/xVbLuKngYNF8sVcpoboCalm6H0/8kPmYOg7FnpLUc9niAauDZYrtDeuUFi9
2y0zV01EbEBwLAPod8id6zCF6rf/egGw6Qp1ZQ6alzMOWsSAPkC+96tfKjgkn0Po
KrDfN556FebzF7Qy5JcFUelpN+DK4Ga/YztP2YT2+yg5tC3jUayeYJnUArSCOp3L
jiLNOWJLt0l2fU8LWb1OB78NgFLrShfJ5XQTBIxJqO4LnqX/c/U5P7Dlxt1nhDiF
DNlNC+XHW3njfF5XsR9kK4POf51GVb15eVNT2MrJEMn5S8fh6JtSQh156sFwRXkq
t2R/JOzFnvWQK+Cz7JvDb94Fmb4fUu9I46kEdJF1yTzNmzN5Mee2g7nQ6chY94mi
I7LSglCfjSS+ioNlOJKAANx0yleFk6tqzoiAz2I9U8owsUusWSYK4hg+nnD20rtu
Nn/KjbsNk6N/JWkGrmhghdyVbwM/7IFaYSRSjBWvufzU9qmeD4XQ2ZXnM2WF8b3t
imYKskfBBLEqJJYv5IH/HCEJkEcWYAIuTlN9lgUB78QWvtxZgvZPosvB1CvYzbZd
kjT8tb/RgvELPRFkkHDclOZvfq9c4hatDq7xd5Vyrm2FQBkt1S5N81kUWoBmJLFO
WJk1/8Yxqzdp+rda4yc6Tm5p7q2kWWQUho+jMMi9X3/jmAmRaDA17R31iibGd94G
vCAzS/rTEup4EzLCaaBeYUEKFrJ3vKl2EB3R+kgs7v9srof21b/li3TlhVXN8ohn
iwS2Y/L+yMT5rUeDs1mNxxFERE4meBXXX7/26qbmGFPV4qqu9cqduu3OLfGn+4Qw
OWAbfTdv/Snwwiit0wxG9yi9o2j8J8iPZH0OY2IxQ281IICPDeqRsccicSzOvBhk
4JRsNxr6JGJ5Q67A+sYmekqaPdj+/whR9yQhgj/5wyphcuhrv/DkNZBUwhhb1WNN
EGRPcE4yIIRpGT3/inmLsXeq1Dg8gkD3UI9uyN/n3h5hBmqM6Xt23+G60eQ6bxXb
tcw/MfpBlWvbfIMtVJhWjsRMY/Ryk/P94FJz33qpVHIteoJeo9j/vjeoKZsWhXSx
NTkGHyX/0iurhFTY0clgjYKvxY6XJJadCJMlIWgkE3Fqe/xJKo/XegLWcIeCt4mi
mOmthX2t1ZsbtlqXQKeJuqEqpLv9m8r6cn90R6XbRgZDacnhukGCi6QjgGkfCQsI
xh9yA+3cbN8X1ztKnEfUXw405ALKssT3rEsJER274DZeOTxxT6sDy2OoWXF4H7Gm
08l6hkxO7ULZ739I5naygxGb1+CGfK2usW+xhux4Tf02Yef+B9UEpe1fKMKpc1cr
GKBFGOs9JL8BZA7hY31g9pCgQTA6wNhXusBYR5KTOjwbjZnIz/Z2dI1TEjbbkdYH
I70BAVMsK/s3RhV/vWDjToy7tbHqSyrJs82qlY7mXnuR0X1+gNqRtoEvs17kmJ74
+nKLAFf2FbAxy8JDPJoDe5QhYUZ5yiV85q4ven10TNio6TGLF02114nb3RmGqM2u
VDEQQepAtMKt/Mben/B7MY22HERiydxps90st8D2KvGQsxNPie4hh4KB1AXHYyIh
S9RpwlYny/KxtZZW0i7TqdPqx5UZaoBsSRPL8Wq41UAeuofFGqskzODr/I233c79
GUyY1zFjpNoL+Xw0EBHIJIf5xviZpdstCRkFPRea+cARS/HnKg4h1w/MzMDhm3FE
9niAyFM8YUzMAV0SlIZLmKiSFKEWmN7D17UsBVfxFi5RXS+FlqfSmJa84TLSK/UY
UtbR3ti7YV8oGOxZQ4rDb7FX6tZhw7m6P4WABXDnHb5tugjieUL0lfkOLjmo0V0n
4JS2oYGftov5Jko+68EvJU9P4eIEY22AHPSNjtJSLdhV2Ztb/5+T9Kg4zXaH3oah
heDmhBmaRa6FAjPR2HmlDcwU67BrzJc5xqjbI8aMB/RxlNH/AG/xuOLxbvZ9B0Ee
oF3chUpnI8qHr9M3E5HoOPFGO1CLw1+YZYeXCtZrdqxNbuRRPsimD+bVmz2CdTcL
c9csg8f2I+odY3AcHdgotWE8RLi6Whez4obeLtmKpy/TcZwS9EaXqGkW/gyudM0Y
xZEmTmq4l3IV8DpRfq9/FSBGt4TRfCPBRxJMoAcyOFy5gyEvfdGSxVKdPnioKGin
vl+pxqmCgstqDNHPOyo2y2c36odPn+LE02l0W8p9RnDVx4ob5yBcyvNZfZzsoxC8
GY57Bbp0iLzIKbhQ5N6GKXlxc0uupx4oolyP9reigpORsQFYOwL7YoaAcVjUpvT5
muYkLjLeQeUJvjMCATnzH33z1vrTgY/Sqsn4wOKEQLZ8g5OmkRDrtt6Jb9kPgolj
o+t8Tju9hd6sp6rOvbdgjDnbQZkzdJ2A/hzMPbt2jGCKAN1xHa47pe8R04q65xIA
ZxmYukHujY/J6aSbQHaRVk3ug8rLLSUuOCnRJlMiQN5ITePHXc3l7DZpyslLt3LT
HrX0NRQx67KhGrJSo1V7ejWsRRqRb4yThLm3Svp2uMo/2Yeyo1nNecXGOTi2od7S
87fQ1pj0WvpcYKOTDuf4FjRPNFqsZzjMkexSL4RDqMSUlKDI30NvWISF6Y0kgDNt
YVoSmExk6hj4g8BxwjOiQw==
`protect END_PROTECTED
