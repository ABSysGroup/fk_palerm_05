`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bo2QjzRMDRsLQlL8JvUKUj6CONvDUcZwlfJn+DRr60inqVZHOTgPJl0i5ypUc49h
qhz24fyKeLHxd6xNTqDWoB/c6jguSOYlcrMoaxyTcBnUL3EfatU44MRqy5Ao+H3G
t4r3eElLCWci+4FH0Klo0b0TAZnXw/uNFD9UPgEFtKk19WAnoNve5Y9js3+KLwt0
baxd5Vu9tZ4k8MgWVvwMbWEdpUG+t38up/AqTqYgT0o8gZdcPK+5fJQcZHZjV6UT
Vq1kuiR24CEJALHRH0B2m3jmxhaNqkYesLGQXIyfnDxdNdiqCaiJcgnHc+76MIK2
08IuNdRQ59ZYcpYK4bYAoCeJ4/cYbYWFmu84kSct/8LM2Kq7EWvPLGq+L0n3YzLU
OOeoOKOs4G3mhduay2HoCjx2v5C406wuG8cZq1Vm9cpNrrOVcv3X7+Qc/v3mpEUh
HHMmrpctVub9OFVQUZCppehdx0fCUDGzppS/3NJsMNgXvs6txvD9Ucnga+0hwYRs
CZm8SFDQBLRJZ0LVuB7hohtwc0OAM8tlVn/4O9jW2/w2vbvAbY6eeey5ZNYU8dYS
2xo47NfJwFAySw8zhuRFwULcZZ1DbJOHOvmmgjxPiCdtgFtc8/sI/3YTYBkoxRhR
DBH5oR5WIE4ZbHOMONMGIYzLRSdnYmAn4e1v23Uwrpwd+o+hfuAodJfxaIsh9P8L
dn664mO71QcS0OHfd3WvbXRWVrB5eTo6fh2uHmFLIPRFULbt7bxyYtZKuQxK6/tP
AULJS3IGaLI0fySwJbfpNz8dZZ/IAQPl1UnXtup9X9oTDv4X3LTnqONt88sew6KM
59UTj240k4FAVpgZP6u+ufaxrYd5XjMOS0HdVZzWxw4AYs2U55jSf6BRz/lL1DPe
DT0Ki+JyS0QtqTwQQV8gMpbWvcZ/gdc6cqgffL0jrvnoweyE1OikK92BXuLy7+CJ
nuiBFPCqShIzrdQJ0ULVCfjWZT95DNdWlGjG2Jz/9hluHRS9HWArMJSu83heUJU4
eD0gU3rl4kLz7gr9BtHWEl41eDfbTLktkd3Cj4vR+grWLzmwBFe+/E9uSswbCpOR
7Vm+RomT708MrJtij0OR1WWHBYJ9a5WXpeNuVaTHDv11DhBdJ5K+dE7jDXm/jXyT
V8SmciYdjGTffHZfp2zY1ZUXhC7LnoJGusUkfPsvYMSjQr6RG9nFkXwFkNPlsvzn
dD6t93mrPMEVg24eUQOr+ynVLyaM9ha5M4CHyohGLutpYGGpQaVrJMKUqY5Z+aQn
VRzUXRhIY7q4K8rS8O9HUs2nJDw+XYnTPUQCIbvVswh7ecVnfhBNSaRM2B2u+weh
UuBiqQOZQ7nmlOs/rR7NDwsMI//AU/HCy3WaYDiXmlk4yWP8clqJJ+CietYwuds1
40UIk1drpRDTpiM0FzaL+psRa4M5xgARQrOvfiwOjPodhiJ7pB8m7vul4DkmpNvi
CsHHsslL5gKwASVbfY3vbPsw5H2ML1on4bj2K8QlRRqMx/a2JFQ/Q7beSKCw7KsM
Z4t5XG3FxtpUMtjhMqKCJlkPjbE0YnxrSy2Wq3M68EhdJ+I3yBhip1WzuWSEVawB
2L/AsdZovftT3jRQe16F2fBTv0JxvORCZMV63BeFmoIsAb4Qye5JoaVXKoQzMVF+
T0Sny/IcCGSjPgz8iXNLXHTqj8W7WnGCy1Ao6RhQ62HLuulwU9inJQL4rykq17Jw
T4FHcqOql2UlW2padbk5xFg1/C6CaTcB+C0f+U1jD/9Nwf6u0EJlsuGalrtB01N6
AgmI6h1Vv2sDKIiSfUgukLMrQYtF3LXx9VRIzQNaBZt2RF8uYI7sZerk2fTypiCg
uX0I1KbrXjec0eXVDq6dP0gsMFnSCsBs+OEijsoY2JxAXLOv8KI2frZa7Zx3wJpa
A+H+AbJb57/vVAJXPB24R39FAf4TNKcH7N76oM0rSGkpbVJpjTT+D+oPP2HDe2bi
ZhMu7WtjelRuoKxiS/ANLw+ERXoHyWhCRymoJwqGUc6oXkZK6XwofOM6mNZNUn2H
TZlCJvbpLDMelnnEpFL4APeUJZpKHtwyCJQEkC0KrLfjNrzzejnZAe3TSVgUSABy
9U23BJ0yMql8s9wRImatL9G9YLkGjFYfhhe47GJUBTXSWnxehxun7q9ufK9YVjB2
we7McyDAs7l8WhWaKhgOK/0TD/fYs9XtGgU87mqiRKTfOWCXTsWXtSm3LR2XCfLE
fCjztKK8KdqcUgjYFikIMJG/K9sZwzQ2hlY1hqnZ39IwaYfAGS4hzDTeljrEeezh
sSYOh5WrZpPwLitfBctSN3bwBD78RZNSEE/ubmrBR7wEZPIYj9yv6MQpp9+3RLVr
vWJIrvjjV2kKlonQ/zoD5obYBFedV3bBenMjBrZvMnMOOKV4TsygIHIGQM9VPgKH
XNwUCS3TKm5aaLfrgjbrefi/monIdTPlXb6kf8Lf6tR4wNW/kNx8YRQcXpdn0c9c
STfXxZGpet5BAc9ofuRjQ+uYXBYngKcsrEYrPNx4e8AzPIVvxz7wto+PkUA8fVm0
9c94CQYxT6KEJDlnN5/LC9MDBpfeTSNfc5Vv4l8C2W9Z0k9kxkUFanYmH0y+3oII
n3AjZ6yrTpGnLdoUEaTeD2eweGKBuwMAg03qVWot+v7ymzq09Ex5KoZmW7C0hsHd
zs7sMeEINmiUN0OSvEIKQuBomdob+F3F6YRCVKt0qeOFvLvG5LI3R6JwKulIfv3C
6vmJManLZntvQniLRPEwYTiZfY/kW9enfl5WvmJMXFCKE7kX6e3bHxxFZwxtiNUA
R9IK7GjXZUaRY+/6p7oEDn8N6FrO2mk6+kVFILXs8xfAwLLGDbkeLOb+WQ3DBIcg
WvBTvoGrsGV5c/e9LD0KQFcSRO4mieJrdcsttenmvpWu/m72+pOc/wsqorrf9HzT
mQYFB2a125q2QOcyagQYFguO76GHs3Xx1WPHlAh2V+V3AcxOzqifyeY9+0kfyKRa
9TGqr+d0Bi4r7t9O15GaBq1DS45IZJiaEbhfwzFOdM6cv5eoqf0gimUlUaSQrL7z
vah+gC0AVr/yN1UofCwtJK5KqxJiwwu1TYmu2l5h+plSllANjZS8W74DvqrYU/rn
7km3WZWYxIKNv7odcvAa4/6+MbJ3xZI3b98Rtg19LTsZl39hH/d+8BM0Quw/37S9
T8l3Rb+46MWZcq9lsn7eeQ5533klonUcxbGL614alppw5olLWUM6rlgsn4vT/hrX
JkGucv1CSxpz7LZD+Bb8E0kNRhRZUH9lWcc4zlMAAEjvtff2npDOzoMJ5sorBTjU
f24ycx3r8e2ldAN9ySrUu/00BJomdFGtrODhY1rK8wNkTYYHBcjpH0J5kJEhqrmD
vrnuZXc8fF1LLr3tB0TiD20IaROi7BHG8wzFgxuVCH7maamlsAmcJNs2BmgDMgVl
3cm6nMoX9eP9d7mfJahHNle/AqJYyoRd83NklNt+ag2cJCoYc/1Rww9r+rQTVwa+
9kYLk0/T0id+L5+JWC+5JnRO1u3xsUd8A4PPw7h2a3G6SfUCoIwp9WBPtCIZ3B8C
Al0OSeIfC7Chckjkt1rejlCWaCf9e9k5Vbj14YS0atX/3HT3s4YdOW+10+5isLNU
DOOdmHgWb0gNuN/r7VBhl8VOtfublSeCASqulGJNiHoxvanwcMxYpO9kwamdiFl8
4gb2yRRtwtNdO6mQ2E+R+HJS8EUeXlOhs4JT1OvKUBRpwSSybDc+VR9IVA8rA/tE
R7bMNRZqgvmpyKUHfYBKkuDVdXGFpc5I2pxkBuoXUIHCP9HDuQL2rPQ/cL+CH04o
i5271zcwuf22o+nms8oi+FNS4DzTy6Df9045/M6hVQ8fwFu3/lYVm1HkzuU+nRaT
myLOwsLrhd1HSbOsjI0Z48oUqySz+C6o+07q0cxHSY8MWOCdR1S0AfA+ZXBZK8L/
EW69BP+QUDxaE3cc1zYqe/6Clef5v/I0J7RbizI2FPJ/wQkULbJw2NWVMLL2VxoU
LcJI7gKkO+4NwS8By2SEm11IsiC8VP5lR0AHg6+UtCaJUDsmMOaG6xtLvMRGBGA/
Om8dVlj3MwYOgsEtbxH/pfDIJBag+btJXJ+iLfYERiYs6lqF0xPwSdo+akkzqHSG
K5VHFd4dyFAwm73YzazFNar4joj78/LCHeMcB3mrsCu9CMZBHM0VcgFQtpUDOic1
6j1FQOc4cVtBuqj4ogSCDq6pRNhv+pgbE/niWshn3/N3istkXT6TFLu0N+htsMYT
2MyVE7f1mP4ouLNUM1q2gaM91W7Inhf6Fxr+9LLN+yXUYNZfXKTeAEhm9GkZgT8e
vmxHlzODFprR1Tgx7epUcYt1wWiRpnF/W64xh5yVMBoVUHGvdEGmkvuSOJlSxc6V
6wrGnj+gozb/O3afzCyitBL7k2NcllSM4DokBrZcmSQ2M9RyjZu27upbHTnTZGY0
NZjMRvlTEqr63b6KieWH2ph0jy6mVVutgsICMdKPKGHbrdP4Xe8XwgEgANX+67N5
cw6knB+9sd1cp6ajMw5fOF2FNwlf0mT/LYTtVfG/yMG7VZRr+5WcHOk/XPTk97Ni
vBJ4/WlgLsZAk0rosodT00Zdt0l8uTeV6jtrOU0bfQfKi5kI/NWPIeSqDQPwMCsc
l55Hcep5+xz2HUotYBb61etN7awHiPpbeEdfVXB4AormELGcyZyhmu+xZyT9NGUB
240RjSkDhEOxUSgvzteVhO+vNw9aezdKcLDn9c4YTDftkb/MzDowsqhl4EyQfPI1
a4d6nDGRZGQqYHUGj0hpHAAqjYecWTt/wBa3VD2YbpL8efg7pRiLoED/J1zsI+DH
cji0m6b7h+1O3U8KI0R/IfKxFPh3IzhTR9lSMWhjNmQpHazolPzssGwWfwW01ZZy
O+4Z6HiAjAkwqTr5Kn6ssofgXsQYw1sbBCEV6e6ZC8PmSl5leK0vwTLC8OgFkfbZ
6Tz16z69YH9WqD7vRgCBj3OqhsYmvUYc+6K7RGON0sYHUd2UgUF0y90iVN4xc5cq
LlpplFtip7rBSJxvtvKiLaNwzLkvUIcuC2Y3pOKbIzmnD5jtV7iuw5J7+T03yfVK
OBRZzYziQnirVp8jYOypCvoRCOKVnXEKtwKfJW8eUAfgQNUoEdkZkDMzVjy3I/PE
ZzjzN8XqriDn6OMqi/RkWVbsF5xe1SyKB6sZlHIq7d8pQTXSqya7JVoQ7AdOpUK4
whDwLFCJPmuomI/TjuOx5MULgw6SpGUGjYdmm8avqThAm/NSbUcNPTdYOWjl/Gam
m7xDknE3v8WzyvbuMZgjan7CJISbPoMxV6ZxnDPMYdfp7z+bMm3EG21Mmp5DXD6D
UDP2T4Nccs30VswoKOHOhT93RZjDSeAHDctv+wdhJ4mhNGiL/bnPdBA3RDZiTLYY
rFDBfcKx//LDpGVSAfwNYKpG/T+vu2USulFH6ZotmHbXc4mMGX9mI6m9KTsZNWS0
jYaHzS8Eu6nC9IbOUW1cFrwMmLMc4n78ih493OKhpwOQtjgbGnx8b3hp8sk7Nk3r
u+PkQfEN8CVO8l9JgWrvU06Nf2R+GgwMokyUP4faPIkqMM5zhKpEPAUHJt4qr2tm
WsHJ21clcvLlG5Jr4NQHaA==
`protect END_PROTECTED
