`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bKcb3RsqMDpip+UMRdmGeH4Hnf8KVEywGvLZMrJnuSJJjYCRJe0spwo8ct5YOJw5
YeL5x0uqKm8aDG4Kaqbvco/CfW+oUOEH0qFDqGAPg9hb8QxAyjzo47mKeAB7WGvC
In5ugLAKjEWplfcvjzvMlfFPEnCSz9SnH7KJxKDkKyedAEvyj/1Sprhkvbqt48Zn
FbIrZyIerjMAqkBOJ2Gntg5VND542eP+ZKrkVq6e7gnMKyMtD6xy3ewCWo+QWgow
aKfzeoKGlZboFk0gZzgSJUb2VAIxKnbQsqADAyrnFzkvqWOfJ2CLTV3hLbUHN1os
ZnhHvPyxQOb8u2an/Y3oXl4Q4fdrUDo+TweGuhKKEfcgVfCki+vERnuwG7nRl1x4
PWcRIbArfSRO9QKfAAJx40NJ4ZGSpaML26aJXszwHr+dkvvz2VEcJOFRTaHfBsGe
To6y2tHjolhvzgqw16Ixhn166Uvw68qEJOhDHonkzp6xzt3NLh3XHXNTUCKfilY7
hykWvooSj5hHM5HXPoR48bVns1v0fNr+5qGoMsU1KOAho+wYeSBdE+5pkFcJDfJh
VrvMAKoh9Qs/wiVtLZV68WmjGJ036RXoqKKT0t9MFVpWr6OL7IO1LPZKMIqimK78
qmBoVIQUPwON2yR93wdZlFQBNRSkzZncNngFIrf50T0VOL0xgkh3yefXruVhmRu4
kAGqF7STayEdxbx6v7tvPg==
`protect END_PROTECTED
