`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZJI+xe6sWKv36uspApB0xATItM/Q9W9Ousing9MDu+vQ9FenbKPhxAvKm64vARW1
egLAqdRcmnxiAiwOgiU9EsdOjCrwYmfWp5k6OcvMZPGPX7w9UuYcA6+o5qy3m/en
EVBcH5w69cdRVwnOL52L2t1YOFR0u1IR6bgmTPegr5dN5wTAdSGwZj/Qw6VBAeiR
h6fPRTy8j9sqD26s6LIOxm62OSI5Ntr8BK546TrgaQDW74K8ESXatbvrFH/jyoIJ
bgc4flCSgACR1JUTyzJgZDvsCxz/U8RcynSFVFzXizYfnOUUvjmK4lkz06BstHcQ
rX+BanNDW1b81W2nRFMQGF6Lh2sA92WDAqtLjLHvTa2m4d0POplOcpJ7j9x1vMxj
IIpAU1VVOPoG2ItfA3abUXYJitThbNhOLo+FMNRzzwVn1VgpDZC/67D3y/FwQ60n
wy2MQddvQRm/p8/r5T4A2l2TbqmMiCBI9FnTiXHLSTQiRgYKDhSOmWIAXCcM1hLf
Bt+5ACD67t7P5q3MiwNG7jwdxVeyQKPegiS0dXw//G1mYoa7Tf7PbEClY9MChn6K
fltyraxnX8osJSVMwmKX0DWyLXGtwcegjzL0CuJDfMY2eaoW9D4S60C25N7h8WH0
K0LS1vHkM1l+7TyQw8oi0tU/Lj+CaXFfn4OJOnC2sLAf1O5yMNdNA2woUAI8KY1Y
rLalVY6Wkg/5pEfOZEaOi5+Ew5qq7n6LHHJfBMMZ99N47+C/ASYWROhjfcIG51xi
BtAJ2sIRvdiWCzWzZtNHcw==
`protect END_PROTECTED
