`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u/siDb86F4aHWP8EHNp5O0UTpI3/sWnisoLwY26dq2uIIrzZW2ndo7My1GR4rIQE
BPbSzDGXkggSXuwwFOF8dzukthUzh0cxpzECckHukmVK4E0VQwDyT/v311d8XJ7G
VBikFk9DmHcKlQAmDp3fMCoWPbUK4YhkkzKJBG7M5T3N+LhgcNlY76hUtwNRajas
pTDHQ6X8E+jN+sz3K/JCWuAya5UPMWyeqKr034ItZi4hjhr+R6R8l09kKg5ItMKd
rqpgmwPpAyi6Sk5F5RhWGb/azd/w37K/nc+D5YdCKB3bsn0Ly958HCiLLPDZo8kG
Z8mxI1eFJjfAvHuojhDyvBrRlXwdn4wAb7spQT3XN1Yd/2OvTP2M5XXldzFH92UK
w8zJQPUcca7uEq8h++SrRil3NXE7gBk5qwBV+eI0iUs=
`protect END_PROTECTED
