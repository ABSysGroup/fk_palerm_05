`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c/kN2OAfA0kIZGVG9WrT6lJIbfGX0qmPwK5HyvI3jVsjYLcf7kQOiVVXOQ3yw+0Z
yQS9MF3YpcM4ZT81uOePchvkvg1We7uAmqxD8whvGyPEoYMyunOujiY+IGiOnRBZ
RwECKMo5Ab9vNb7MOrxdbPmBmuquKRYSstYSIRWHOksV15FItl73LKUXkxfmYBCX
AflUuSZhgYAGARrF+O8eixoV8VRcMM+Fm6KTiNFBGYe7N9NWwQKMv9ekpaCuWy+u
IroZahCWfR71WoAzoECYAetU2rqttgZdrbbSSf95MtmD3Lh8od+5M3gdYiaOlORh
sB5Zdi8Uo8y5qRmsawb7xg==
`protect END_PROTECTED
