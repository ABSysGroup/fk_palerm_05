`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aEdpyUXBhXm3blJAK0kG3Nw0wo/EfkNEhKi1DWjibcxu/vEL+Q2AeIcEHO8pKzDa
P4i1g+1WnJvg65dqHHQOtK+fV1OEFA3wStfpuJOVsIttX1CBb6RTEJm+CRMyPShY
wgZOLsmtn+czSAPXLvunAoIkTfaiZAFJsR6iF2SQEKMCNYXheyNMtpTHasC6AJF/
VcVsRRMZhAkLomjUiqRA2BTWGGXlJ4evmc+mfY0p6dNB85OH1H3lQVMBiwPrusWO
jZlV9RL5/X2dhQF3M+IrgKCr9E2s0epaNJme+WMfaxvIkWakRqxGTgWV89PeTB25
GVdnFwjRJCenKduqjgRH/Q==
`protect END_PROTECTED
