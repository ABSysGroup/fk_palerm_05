`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZweSPtGdeReRzkTl5N6ge6iOYuvmSXWgrzn1pEc2XBNB7hD7v1th4PawzAmYZuUn
PQXrJ54R+HaYut7gvU7kZrrxWOwwLJW2+C+764fnk8cw4OE5fZmrA08I/CmgvHK5
LPewEZ7abrmCMmHkfJ22qlRJ/rlc6xNGPkCtF/mTOg8XBr5jmq/10yRceC6XPqqy
x0qox7myIZ9N5So2e23nmqFXMdMq7YlWbp9/BrymRjNc+jRqsYshT+ZZN5ABOG3v
9jW5DKVDhnRrBQpjIgvlyIJvoTyjrDYdcYpqpgQa3Z3r+4kF8UjuWZMcOOGbEITh
yhoK3XcOWex4k3b4sceeltcB/+s0Xhj+ElSZ2ZWFIc2zbQHJkXkGwPeo+7KxzBoI
bxEMgJAcaCUCm5OYce/DBDICVFiZzVT6e4tjaIBtKm57JHeY+16yTnT0e0+EhhGm
VblITqf8vdKT2oK87zSzFaeCI9jgoYz/gXk15BJi+rnIvPckAHq2pT0bbTi1N1WL
2dbr23SvQFxs5wFV1ycuO5YCzZ0v35SgEGDkrv585BHm+RuILh/vrmOi+duguRgE
Mem3dbVnRELn1XbsWPN+lmLWPGNkiOkGhVSiwfqV9d4C0HcPxulJx2N9jkscPeYW
ZDVrZHj8J/vaLxURYp4s7urmbvTtqDiYA2MLsxY45js=
`protect END_PROTECTED
