`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qSHsWM75Z7jmKsRTfya0WqXsP/bCN4OaM11cOtQKHWlZDlVhAYlImf+wwLLiDR3l
oQO4vk4eSALg26GuJRl6NLeloFyX8ighgNaLMUxojapyKAtvLsdiwKFevO8FRDfu
6Im9z/KP+XnOjr1O4ojHPtABzxNxqpTRJNXx7x+d9X9jXzQ4Cii6xNQmP0lz4NMx
69VRnDaP/q2w9SX7BYPszAEGvqMYu2paXuNsJeqXaqM51i+sqezcsCk8IEOIDSNH
HQD4m86aopoaV/0iALKHw+vepfBvBmC8+PiPvgQgqyx7+F7g56WNCwN71GLhFejB
/Wk6ztk5PboL2IdXJbshwMmoG7lGG+30shQNJr+B/Xy0gatkFQH8F0I6tFYIkMfT
/MWZ2Jq5j6sFN8T6P90h/0VBpKhOOLNRz797S4TNxez3Ix5hk8+OJqQhcU0IPxfz
7HH7KG6IUkQBt/AhmzDxjHpzz+tyUmgfcPo1GI8FpqD7hg4VqafSqzYhGxqSH6OJ
HxAt34OyyFT1aFhyljvkvzUNgFYoalnzJDA5N0fayMJ1lZBX4DOiYlGlpSl5F/Vk
ozlyEYsIKHLj2+3W3libeoNe1aYNHVTB7OqAQgI88mE=
`protect END_PROTECTED
