`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CwioLHMnZvfBDVtozUzxA4oHp5JWb5gF0GvJh9KjcuzMkDuoM2WeV2JjLCBZu9nN
spt5py7/NVJDx8U6sWXCotzmNrzezcwra++0qbHbiIEoTRpmDrVXO7s7sHMJ6MUa
d10hO0xdrG/8ng1rqE9KoYAcM3cykUF0f6RTgzS4Bktvdv+5UT1n2pkJRxvRLZPx
gcfduWnXvPNQFK5grLOCfpwsOCwtl0eKFMemuGx0qEevXEQPGZgEYzwm6fGhzDJx
YPZN58whVvJhLDMP4G1V4RPR51g6II74jEKJOmN5vkv9VVhyco+AXkNnrAeyGhGc
gDev06vz0mXPruNgZszFDmdktlVZ1PIzcnTZcUkKGMo=
`protect END_PROTECTED
