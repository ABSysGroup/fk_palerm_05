`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uNxxNyX/Smnh5rSbN8U/Mo3zS6FZJ5X6uCeyD8FnYst007Bv7TV96xOWTCiO7u78
mAmyTBP+UwSSA9wylOtpMtd9DXhmONjOPePymjGtYQfjwqlOeraxLzuu9MK1ciPb
H0pcCTKH5Ipb6u6xtAGfIR6bh+QZsS2bAM5K/+8ZXKPTklT/BuXi6I6IYcqI1i2b
ZIBswZ3DrKt9Au0jAEBwWAd7O0FoRG8qPjVeBkDR6Q63HgJVygANzoahlSJ/lnHB
oDOWgQxgpD3dfRmS2RmyEmJJDEWlY+/kdI1Px5XA6iM1EXh4aWskVuCX355B8g9G
KQldgbEQ21csjP0gBI4RvusBrl/OLWa6l3O6BM4YFNSoumkTkkCgEm8kPuViyS5D
7RDMoui05l7DH4lZc/q/8si4HcNbbz2KSayCgXQJVpcixnZgQ0E81F9g06LeYHHA
XHYGFfjr7cRBQAwNmLrZZ5R8rupmv6noJKwiwI+jFfgyMWIM53bPhuoV6RZZaJbk
e3fUofh1Unk5g4XaxzR74Zwt2IJFLEYQ0TiCiNVLAdHidwwiTZOPavcViRFOP/ns
INwhTOOQS75wusZ855OcvZC1GAbkM11Qa6je9aTHQWzyPO5whTeu2nWlacqxTFuh
nfIpSmUJBPWAUib0Vx5RZSbo+hGS1ok0IHGsn8Oxmdxf7eExS9XOQCnR85c3SrCI
rlnSTEHbaF9KcKdH967kUHR9Idk+7m8QYhxF3LKERDWakYB60+n0FnNVprz0o3sh
//MlWtqA4azSOGjH7wJof+yxTCuZ76QjEIvSgCfOzHKoq6ofWQxqu9GhXtzoJjjn
PFabc0C8jkvwg6krZHxL+awfjUpUTlxuqRgCxqvBHji3sqDX/YXHawEXlrvjgCVQ
pP85x/w9IW/3UyEVyphIffkVYkS1B+rCxJEqBnlEVeldC7CwyN4Y1dwU3DU1d6DR
`protect END_PROTECTED
