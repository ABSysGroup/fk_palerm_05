`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X3Wtyn7W+CptkMXySEZh+zOec4wPS43xttiiwcykYzgB/1k2khyzyfio5JSBuJoE
3iQZ4QhlBk+Ozeeyi9O0L0HAOORqQQo+NSkBGTwaMbyTCZYNneLhsUtCF7seSDxO
6zVx9vFngdPBLGgJ2aQGHSQWYOcQbeBwpql5o88L9rzEIx7auLT2Tb7zCAZYdD8f
rSorpxWcgAnx+/1HEW9C20go/gdwwXslcYlR4tyUFbefc/sXG6u6x7i+Ozdjj9/r
Y228JGo0o6EasTPdlYYpE5GxY1NHpUAVo+vSqHEqm5a0CFQndOEM3rm0uz/GYkOJ
xL86umMbscXFlqfah98/4cpu74Jz9WfgxcpsJIhAEYawq4G+Ys5+LFQR3T7rg0ds
k2rqEWqMSkprUF0A+dwaltHmuEcAK6Gb4AM2aOP/kxMWwuF8sW21xt3uvzNyGn3L
1Y6dmagAWMcXRa+geiMuyA7i0BYlMaI0va0aXPUyz3X5j2hy2VEizeV322N8Ud8x
XsgpQBLkNl6wqU6twCDEO6qjZIRyCyjYhL+aWaBGYpCjXACUJL8329B6J+Qz1/4m
tK62eDLyAgrMGQ5FsL8KjU5Tm6obqx/EMykyXQnu4TbueNl0KZ8zv8zJqHKzbxjN
MDD7/EDhQZjTkToRn985HuDe3R49fdB6UPJvR6ViHRpNgZC9WtkeJGXuutBVBJpM
vdbZOIJDFs8Aaas9eoQ1v6KaVSSclSb+eRYUvNtjMmcisbeMwHL7WgJlDG9AJYke
rt6XJcKHhpSnzT61YcQfI3fdIe0RNP8RTUVM3eXycA8BefKBHDHLT7yVTozkxDsV
FzDRGEc9VrMN3uTJcaTgMNlGng8rq/8qY6/fPOHKAhHB+TQ3zWvC2XVkhunjTsXK
Wm5L1XYp+jibhMKIyN5KmJ8UXRQ4AT81FJsd3T1auF4dpl9CfHw48Xs4RZEBz3aQ
`protect END_PROTECTED
