`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R8cZ1SYh/C2oxEIY7wqLfbIRnCL03DHAwUsv2afqYyvrDlVvdXq7bhpM2vE/h4n5
9+7rg4hA8VldpDgnNS83qxzFJUOJgT3jwXMKRZRxJ9FAK//sL13JKjmA7V5OJGsp
9GuYG9okb1r+7T2U2SWbnt1gfFVTsqEpxtrUHEJzIjyhuMT/Q23htB7WN1XW75NW
iiG2UdkpMRUq2P8obmpExr/Z51gRyuRvvi9HDFtBNtGIMAo+RBe6x+AQY2nOSROW
LrbzOLN7rxVKIUrCKyuruID7PkgUI+5VeBgHsxfDFdTkqPkRasnFffzwft/btOyE
brOFP0/j2IJkmT++PFe7Gg==
`protect END_PROTECTED
