`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OhjWVgS6dew2p8SgA9C89EeaAZAUQGOtjvtis18E6X1M69qNtaqazlC5nixnesaE
7bcIJaw03LA6w08MbSAfLVgg1TBdtQXJATfCkBxiwmohAKnosX7n/6qHlxbWMHq8
b+cMK0Nl6J8XhZhhEw/xBiX5i5hQqyfL7PJfkKZhdDslXNOZZ/jj+3en3QZUhZc3
MEoGcv7XYy56BJjlufoaHqkpJ2ilBdC26NUqUgOrO9njXFrHuPq9mvtSoV15jriC
tq4i5rcBK7/T8ES6IKjTzxhlH4nT/jbKD8t3TAbnMZdFhPlrD98D4s1V77+qjA36
uxGsw1fx4GMgH0TMmdutR4sr64j4H+3VxN/eXblRWgHROBNV5rZnIb1icDH4pWgO
5EzP2m1rj2K9UvXPYhrhCO7nKblVIR7lCzIxBxwADoUEVdT1qb5wVYuJxWnpHj2X
hE0amknxLpcpJ6JaUYn4YxGb6iryk+W8tcoXzPMFxSBu5ghkRbeUdwvjQ5WGKRYv
`protect END_PROTECTED
