`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2mZIHAakvCNosDHOSdYoJRlorVJ8koPOEyLYBC0l2HJBwJlZYGmeFnAh30zPy3xl
wUJZRus+wwrkriTynSJdrjheg0scz/eFk9nMq1TbYJcGCiBsZdxdxHMDdgI9X8Si
rgXhYZqzKxd6qb1y+EVsen7BtsK6WZ+Ntkr1lRhZP7RbgKCDY5R4wukbe4WelKH8
NmH9Efpee+QWJXn6WSc7F8VjWR74PsE+c0XRr34qf5wCER+u4p3KsHM52Whuy42Q
LRYVWC2Pspte6Skftp22Mfp90cljGSbiQ1N0MUPZc491Qe3O435MlXzrEF5mEgXU
q3s8aShSyVpFxjkuKiIjcbOEDY3+0AxJgZk7qtF9F9z9rqd4FnpubEQyRNxdwxVV
bv3Itwostuur99COfJL5cGXNto4AV4JdO6D/Va+W1l6kiAEa60BmjtHn5FzKoDwu
av1Tb1Cy3YZ0Emm6uIWqoy/nSJUQrZqDL93V9bm2JHYR+j11DVGcsweZDJzuP7m+
znggciKzzyiqh+gQlGRRL/ACP9EQ75AZk4uK5rNN7LqBfnbJe7v2n8RAiEUEet5Z
9kpvndAGJ6BtoSCZtGn8cneOqJk14nABwOMWV9FgaKuL1pmPkI/bL1Imoy9IiB6J
V4BVPwZYLxos38PTmV59St81amBOg0H6j3b4w5MbwzDAReOzOF1e0mvP5XPxt1xa
HuyEAjJy5VCUvIBu/sGriZbwjzmhKLl9gqsiKX6pLO3dzEkgqEaLbco4Q0nFBytb
0IDmuDqbXBDgFe6gS10EvO6DqKNKwIRrKOCw+jxGKaQ1+scjzWKDbG1do9GtbFFm
1metnUxyGnTA/s2nuAkglg+/wA/P2S815DAfNB3/7ua31BWLNor4ny/b6A8XgVHY
i+Yqrgso4VLwGMfNb44LgTPy5jvsLf33JDfegpNd6pwOng+gGbmcao5HLhfiyw4/
qawjmes+I0Y/4vjtITU2GzjfM8kO/0GoG04JhHu+9xFTDml71SrFxLWfJesPKKqv
wqqD49Xc6NId+uhdoD8krbSW7q8h97HgAIXGS6ri3OO0D471Qnu72NDAgSWCANFr
MAEHyY3pJtgW6BLsuYghIPXXDBxV24uKZk2WO03DuqGnD6j8uJR34ayZnjQ46Ym5
PpZxUhXP5lcGX6mFt1W+XmucR6ZQw7GeV6NlkREejIroDpSMI9iOYuZjxBuVqZ3T
Ts8mSnGGbXkXs4HDm+TaHATeEliamBrOgi/y82wFTF3nRldcGd87aBdtg8Cps+g6
c/IoTsOq32ZJ0thyawbL3TNcrAiW5vDkxx7++k/xVE+sIhwKjdHpq+mxsw7DA/vl
9kbKs/iK23zZNd0zccNfSp5oatzUzD3CfqS0YK9T4YMlAkRNgWfXib0mEnQ1Ktgp
XtLbW7AYF2dZunK8/Bxv0CMR/FJqgJo6rRVEqi7q1vSpmVpaaH8M/vZRZHgth/ZH
7ZOBlJquptrjhF7MymOIJpT1MdfGMTnncaEa498uQX5fWDdu7+Ij5obuYyUCBj6h
A5Ag+D7vOWB6T3ZjMXZq7vt1xt8ChEhmx0dn3I/KKffyz4suvhr/SXqD0Ji8F9Dw
qOOGXgkpkK+AjcewPOSZPoFXpB7+DzeYmUbT5aaa1VA00DfiZ+rN6yhvqARa+BWa
nmrMrlPzmxiphdVEkRPkhTSQrfTvgnU9mtZLzh31EtEpnuGvK1UEX2EadEEDk675
un7/dEoT2n5oYoGaar4T9LI+V0OfVkYj7AvEPlxm4FDjpQF90qHZDLqeS2vFEwJ6
BANNDWkL4RcQrhMcoih9sKgMHIpF0vcC57cjBczsWScRQ1p1Jbek8TXa1JCYIcpT
r7LzJ97PH/lVW77bhJIZwjSm+soUUMqv9FfKbuHubnc73X1Uw4E+lVJDY4CiXeOI
ZxkMh7e71WRc4VEhhi0zRF4fJentPoRhTmbGVQGfqjidOxjrvopUUYtwYzTxN/y9
TIEtQh2023C8Z1QUZrlR4jdAMaOxq623yQX+8mwu+1oWRPoA3w2j3dHqboIX0kTC
22SYMFTFLyV9IOBv765PJ6XzHbKr7hWs3cmeSCobz9GkvHKMWUw3A8yK9y8AndAF
ehSdI110/CbYIEQBZYLpfuBEQK2SHmQfyX6WNZ9DYSZMlYfIoGLxVX2d86KoaRr/
TviHc7D10wavYhEHz7a4QAajS3u5H4q0oKl8o81d/UCqWzXSftrH7DiWl3YOMs66
sQZQe1rBw5Jg/YTksuIIBvgJLdb5bXVtLMUINK0xrorHeQVz6temhy88UNlv/Emk
va/Oa57lfk31idnkgJSTDC3jUYmniXg5u333oAmLpqRDMONhXnxQWx6or9J8syGK
gYMybWv/N2kOQWYzMIUem9/b0nYBqamPu2He7Q8OMrIBhykyZKvpeCl+JhVXpAeN
sktFMX1wKJFBAC0qAHlDj5hMNrv9FesRUmkLqsjn0oNJJ/BL2ae/ecjI664lV2Dc
rzizl3g82UvlBK7rM2DsD+e2MtSdXZ94yRaBRd/0aH6i7JZB4cyY9grNFVc2nCQr
nZe48k64YxE0RYVQIC3QYymqZu2epPQn1lRvbcBitJ7jrCKllEmppkR5vcbfrlQs
D10m5lXTN9mkrSMLzEYzNLXVHqlM3msu/IyW0chblwfWv6y9rTQPl20wMm+wVrF1
1ASOCo1lynq8YQJeKOtjhNhCLE8Cd+V2zVOeEnmQX+9c9GGZJ8Ddn1Vl91+QKNsG
K9BQLKOyEt5XrQlKL0vAuVxAhVBuEDlxRbrgR+ZPQb4Z87RPmFnTeHeDDJdbYEl+
vyqf1OGI6o+xq52clrZKCmTZQTkrdKWNiSj4+4iDSE1zbHHlLrl9pJPd2Bga0rUz
BAuGvPLgB+ODpm2IaDRXUtigMSiZ7inBLNHubSYYnseHVOQ7HwqDq7iM3Qsc282c
z3GQMVaOW1YdNwB9x3rjJbqFUjNN3VOKgJ2HIpJys2honvDKUPJC0N9Nz2DRnNVk
TukSqPeL1HRb0bOm4SGWfVcc+St/M8KfKUG+Bu1aZo2vr0CfjkwCpi2R446l+uIV
nKQXn2XFjs62ejNBOknRfdvRwFC4vQvYP/LuUi/X2buCw1i21g+ntzd9M8L13S+S
ryQl8Sp+tNdaDoMb7lsAiYQIe5aNv8ZAY/N83AQc9x4fCnBizl50IqzV40nC0oqf
jJq/GtC3gpYnp3hOcyEafCBcvDLXqL8UMLGBZHIiCT6lGUXGD70v9Hp0d0ArJCHC
aGWXOyGkZMGcGjuLyw2bFly5gwI2AMVIgN5iRH9f4J6b/Qet4D3XViOt97Ho8ZRF
/9e1Jf2ZHQfE7PJEx72rcanRnGV3w5K6RV5X9e2mLGvPdJswhBXblG9li/90avQD
VRw+4Cz7q129Qq6PitbUu909/f8+DuX4Gtp22YutBD/CW9VzZ4q+7045tEvUnnD/
0TSZVSKOasneGR5nDCOI9BXE54vddiWLAjB3+3eXdIzsIixweeXUawM21rLAf5S6
RCiAao6na3FWIpZA3uQmm6jV6dTzaZ5wU/H0ZtU72Im5QlI9sSCzGS52o8z1I9VK
E33o0NuK4TsYFwDzDtyAxyOHRATrh6+s4N1GxtnDjL0I0CIyS/8uhVLJLQ+hkxxW
zAuJ4e43n3kQertslUSqefdpqJ5Cys2STNg89MBsK2IxPXWdm3mfukUTi2TwjSn8
a2lsDh87VrKSgJHzq5mLwLtvwJqFuJ5kC16AlifVLAJpZYe8PInkh/93yBOKEbx7
MaC1XPthorqjJkIaamdi9qvLS3i2GmjGMPrOhv4DfC6hWYld3TJts6jas1BiQJKu
oETplcUihAoVEu4uOhh5NnxxdLtmpjMsSP8pHGp6NfvabUdIzgGW6qWUuxd/Ue6d
kPYk3Po9jWrxgXrJNg4JxJamMsKRAro6nnFxzp14f5FJh5bk8bdeOyw/QxoVYjOQ
NW99qULxmV+biIaCPk5B1O3m09TNOZ5hUl/R7s2YDtwRJJlrgzgz/Am6d0B7EP5m
JWPVCkzg/yzAnDSsTiLzGW+sHofcOnM5zXGj0nGvoa48bdDKoYDNRLMqKdOBaVS9
bx2/wKx4IrsAGm6wW5ZrJHUx03hhvlVMR3SkISRgAjM1mufntdxtYB0D8vtOEf4w
tS6CKcy1ranBrRi67qswSqJCraVNijSTIpWuuaYEeOwweu+Hwn70W3T8MPJZXacG
FDz/hHim/BpFP3k3uBk5+9OHYHbCI1M7o/Pl5R9funSK3/UfSHLB95yAdXM2CkKh
DcsPk6aS0dYmmmn1Hf4ABX7cBQvUlOb8kQwCnHKyGw5eU5Y9T9JaAlR7zUZyQt7d
+ApwyS5EfvZwd0SerHfAh8xLcuCNfUg4OUMvj1l5kT8Lc8DLlzw39Yb1BgsTCIs5
B39mxrzUWZJqvMU3EFzVA+vBcgDV8itJrEHdRlmcZLcOqRCvdZcUOV9J+e9V6DO/
ZE2t/Gg93FjeJ1uAp5lv3IcroPRrwPPQs95y9NXtis0bCCanYDaYPDJGBn8cpoWS
uJwSdDvAOyhuD3EAiCYdM0Z/n+GwcILR2jL4yTw1IpRyWyyRmnY/2E/FGaOk9ydf
O4DShqfA09J/oPfkiOtMIdgRXfLT0jGspNjvIXr8CpoCQBtaa9ci8sHomoupMnTm
TSUUtQVJr6/c5ig/v93WUtKFJjKAEzNC/uW2fpaAb/TrS4Jtc/+2unj47Sm5h5N9
uHQ4A76C0GsvbaXL0KIUNbU9qg8baa5y9Ycp+3A5xQAsbXnBRdtJVmJkV1+DZRF1
+iIlFEBm+Im2YhD5y87kyoIUPKhk4bpADka1Y1u9wWPusiGBb6w1IP3Nb6ZtCmHB
RlIYp1gqEjRR4DruLruPoLTEP8YyHgplSh8d9kqACVcUNyxQn0Wcp3MEy+ozLeS3
1nqFeRB2WG7Jdhds9r9LtnKJZu7hMq8nw36DfWWgGD/2Q6gx8+4QgdLHSUUF/1uO
8lFKjJKMCADUROnpYGRqRIH6XZk3vcNT4ql66plllvMdaymU5FgoY/20IQ+4vMZe
gZu3FkobU97jhgpF3g/Lfe9ReFrJaICRbH++MXPTA7AMhvmTpGoKP0/T/8dxHVqD
TJzT/X2DLKM0pN2Y6EIc7ad03wrZegwdheOaE2QzqiQaFkkHfRln+7kUeZONx4br
pXi+03MdYS3dFoFyWQS80eN/feg8vwarkzVORDo8K0grnwYSFtbYUQd9V08gyuMu
/Ltwr11ES2hOzRowDK70bnZZq7W4LKSL+2Ho+a/VxncxumVu3plAW9ieypsO1yN7
YPXZp8qHNH9RcwlEViBVvokqNiy0Jzjr0QTbsVscXDAK/ops534hYSIkM52EuY+G
3W0cHKra5AprmxobHyDtrQ==
`protect END_PROTECTED
