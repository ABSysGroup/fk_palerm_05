`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zr68/2olcZiHBuYFVa6T1jb4dzf2kfFL+789d8ut9JnyJLexmpgwdhHTOx9EIjuS
hk6bW0418kto0Vp90gL/Xlq19sCNvsK0GUIb02Rwno8TF8xzSbgX+TbVnFsrHUha
PQvt1EMJHZ5SSyyzL6bmKRFs/ocKpyPepGwK0Y4NpGkrcSPBd4rZQ7rHMm4H2xcy
kZ6QBN7ACdlY/lYnEpbxVKkvlxevtJb/v0Z5K0iLZiKIO389Xapr1DGoXA3oCaH3
lBnn+N+NCq5jTjlqWAqkEPE+ymaNxyq+i/JXWKy8egzWB4PpYBMgkaaXQU/OmX2I
eDv0lXjbiHXQ4lyApuekvTorGyvKqqH14Y30qtwEHAs90D+9KU0QbURUkJprWrO1
H8nMurfDnD5UlvNl1bwAndepN6AqNfQetY9Wak513tO+LjT1pcAP1Fqw3Uj6OrqE
/9aZNGDgNwYuptWVfj1ZLcOC/rNNAyzZzucuQ/y71LC34ueoodEuTfaR3nkuVruV
zzUcrll0IFgwV1vAkcuaL/82FVwzg/epuCaB/P+QhWTp7Y158kTlAs43n3vbcFgR
zsYy3Ysd8zdRaVCCroH8iPSj0dC1Aa754Kp24AvlFpKqrfkXxLRVYTQHOgYG/xMq
zyeDaudY3kmxIZhZ0/0xgHPaJyRuz7j3jlPHQzzJu6db0MA8biPbQQvtb2jBzsCC
WeMKYtKdontZRn0zlxuhw+xvxUTHXpeo8LqE9LQjamBudavROhIeNtFTL9166mdI
MISPKDTVPq09Vq9D43dN/RsgjpDt8RegYe3mv0DBjqOXvMxZoYxhXAVCmo6+5YoZ
SM6SQFXDzImbFVOGu4u1SNB1OMgH66ncLNSDwlfsJNhFSTSkrt+sc8iOmr8r3jVy
kr5mgNg++ehMXZyCpPOENnII9v/wCN1ttOiw9DJW+qDmPXQUaJXBqTHRoY5e4iqS
`protect END_PROTECTED
