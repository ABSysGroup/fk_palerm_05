`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4eVLwgwZJxWZTnQu5ZttVnytSwRp71hq4DHBHEDDImMIFbDIZnnutmChof+sRlbi
AtLOVIAqieYcCzK1FQGU+tjoM54KpraI2NB29ZRmQuz/wkVnMNJog8OE0pTq6/kz
YfuO5Vy7yX6TSdUsBI3twibur88RF0b9XKxnIBje8c9yx3JEQyboVh0E1JpjWKGT
E6Ih+mZ/2jRg+KzwbcLKjoovFCO6U7pNdRsPoRJ8YvQn/2A9iqUGqgpuEGjJDxsA
7vDjrOJxFntdB9pWihSku384mGtl8po9gAOkMLBeBVfMJn3ZrDYEU/TtYKl0lfJE
cBG5zguYHzaKDkvmCsg/tmE7Y3wpR6t1fbTVyAtGt4iPnoYyAyB2IuSXFQymjhjc
7wCgYd78SnAuIR+ADySg1ngNb6pS4NdCddQaqgQv7o4hGfDoU9y31h5UCquRnbmc
3ZtWx9ZxSn+FTcXk/idLIxV29SgA38yOF7iQN/9ezg4U91NFVae32srVc3dWIMYx
R1DQuq1ypPKo18oLgVBhiFjmLg7z5Kvktl7M8lqJRdzEFk1vGRgYECNBAwSVLbZ4
ReX8PlDj43HGIWbaq4zU1GQy7jLDw2PpSW+E/uX4N5kmnz2QNAVnv+5QQOJUFEIs
6K2aWQDMZBuKFpAvscI5BswAgmLg9auYObVN5mscWDVweV1yqwcleE0W1uZ12R/A
NA2dqUY/OQ5+nqA6NPnI7smFaEkW/hwY+sxUMSj3ORsPcH+BceWCZf9Hwq3C6gPQ
jxdSQYD4FOMo5QND14GmzPspK5fu7WIOFS7cTOe0KSWsm71iImdfCDwmWqRLZQeF
ipZYlWdugOLrauverV1rTjjyAJKn4bb7HLzp3/ZUvhLMcbSupZ5HDZPnwHjD7xdS
5gTKHsHgLxgv+As7ZPoWqI19+AjfpvtGwPa1NIoFxGIPdi4PQ9zFL2Z47eabcKJP
7FgE3LT2GbFeLDZz2Ow52Ep+uee3tRJpKByAq/yfLP5Hs0KX3iW4HHpU46XZTIWI
t525ZPtOQVkAgEpobAD/uUNGuPALA9r5K2xm/P0d08ryRWg+AkIdnb7FsF0/LaBw
+ZjUmPBL8/bFPW9Py0OLu0WNLO+BONXTZNJNMCVkZ94Wl4kvGKAkDgZRyo2DUdBa
2oLXcWDp632wHl2uCMgbzAVZ2eYyUSj1RGXSSnbW1nbStqsd9xVLgjCDNClB6i1f
EqWSYwMLlS4gaY5b+E8/iGhi8YqD07wxkogdtUO50cOBL1aHT9mGCHe0wNxmux1t
uOIh6ysmbhRQPYWqEsMsH0i0V68s2qeggvJBmL0kdhOcDU2rHe23DCBNGVd+2dyY
8DiaENbsHsuHyZYPTVJUw1Oo9Ns4CuAA6TgDQ6+4KFc=
`protect END_PROTECTED
