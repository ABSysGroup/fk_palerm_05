`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9kYD0RbF3T9kt/6bepJmQCBqygFwC5+Eflc2LLegLehdcOERYjWAc9DAc7Tn25sc
6kWg7f5EoG6DNccyMD85Z6vus1pi/6Ai+Ud7LY535oZzKTjIsRlWaxSlmWt+RxLQ
98k/V0wkvizXaQWfQ9/H3EHhF9zPNz6fZ7VyJ8KiPrK2t7gDHtGGxcONGdBO+7HD
f8Ktw9+3ZSOK4lCsYfxljVLEoUoI1Yp3noVnvOLPrTI0C/B+R2jm0mMNtOOo2V0r
yyawU4kPd5mo8Ec+PoVvMOHeixaLoeDigHAsyWrTNGNKKJrJWLTuHTta39tcT00e
fD8DAuMFJu+blKg+GUimKrWddOAi6UEYb9D3iMjYRdejx15uNU1l7YaYOsMd2syQ
1gHP+eSa45ZXyWs2M5yYLfI0vEm/fcZWzN3bHeF485ozivzHszGUM75x7MVQjUbn
hQmwXT4tGd+vPlOS86ijg9uv42sQ1Uc1OLQqH7a8psX3yzhgBGk4ahrsg6xGgB4o
LvBRjZ/66Mgy+sn5jDdToXZOyKfSho2mlkTL2H7H18Yw7tdgDxVCbMKpXwYez76m
uZKyueCPMzPBsr2DnT/8SsYlV5PFy8uLOS5m9qM6C8M6Lpa2UTvwRma078s9DxMZ
nvwshNOWszRff6jSnzadfDeW5guR5w2XSTqjwME0Ji6RpE4/Z4EXVkgMeG0gPrE+
/Ny5CgG38MtQnJVPVBEgqJCfaQJJcorGo+Eavd0CunDfJK1i4Zth3AzorqXr9iq7
xtXrdM0n//cBr5HiPJE5xkf5xmVbiZizgIu7AMxvKXmbyHl/w/cT1IUIuRhbbIYv
rWt1Hd/lKBbh82YzP+1maKMrP3RJ+UCcYnML8bp15hREtrn7nE3Zekvj+YmcJCoH
YE2b1CWjX8SG9Mn/VfyA7f5NYILLvJTjSGbcgFlb4wg5rkQBB2bKw5v8qP43ddz2
TLLFiGjXEs3L5LkdCG3IlImdW2i5m1aOVP0cG9BFZq24LW7TWkKTgP0lWurmC/wj
0EIJ1UmFd9IZgCfySZKgJAcWfqXJFCcvIFuU7ZSeg61JBq3Q6Yft7v1aVuNUmd6+
YFltuNsMtvLyRGiuvWUUMrmKiqk2iqEoqi0891aUcaSkofdemMGXjFs6ENJLF2et
o1rx6IEEQDqphVwgsagZsAP63aBOVm+yWOMpz+/i9iwvXV52RgeVJLo4BNDuhdNX
lEOVf6XZwI9ch0lktlUsKUj424f0EgJuvs4KqT8XxsuNm9b41luDNse7xwIM2G/v
rsMs2ootYhLKcavB4/TwqxMiJCIenYL2qU7X1WTkwLDrC3j9Saqp4kNiJUN8rgCr
iGTMO+wQANzroYfskFJMLcOeKycNxjC9m6NsrpccwAr5Gs1dc39/XhBJrVDkK3Y5
du1GTFg5wCzODQVJ71CTsU2y9HDJITPNOC63vkiF2h5U5P2mAxsWymaic4+A30t+
9RIxWirbL7hPw1XugHay+BnXDu2259bxlQxNsiXpZL0tYE0TRBJngseoMsu69DcG
aYoBlJEwx9FRsqOYaVENXf6xvWey0PGJcoYV4xiMg9172opNOgt40C3mEj1KEXmx
FigxvU3/oCTd5xI6frlc2Ee2UhpXNRIqYoBFCUcOBGtZZVuhwSTIREGDILncX45E
ERwoAngpffFj3CM9nlXnY8OPq2+Skc/8Byx3xQzZSN51fLT0C/FkYJiLiKnOh2jB
rKabNUWdYf/UyKQ3GpDb86F2WYBWc8cOOgYWdaXe2my/TLItUMJCIXritDE5EITl
pGnNEEP9ndkHwK0qAgkIvb8TEG2ZDVt2wolghZpWWgZ5mq1OnLEdGT2uDl4qRbrW
uaC4NdxUJ1GrAIJ9nTLkbeJoVhS5X5f0KhToUvxjW75Y2FCBJY3+sQrVozHEEX8D
JGn8bnhgjuWSh8AIrZqe/oWcmwFassHiiM/RGR2q/qb1jq4c3NoUYbca+ux0veH1
XogOXoywNkj8Cv76utb12FVbMMkYLiYkgp8nQhPBJKeen/9p8y/p6UxR/CYs5moJ
`protect END_PROTECTED
