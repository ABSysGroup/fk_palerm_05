`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F4WEzppol9D3l6EPkzSmvwr4Lo9OmiLgUjogzj3vYPH1mmkO346smKecV5YI0PPM
6Jw21pQZZEOPTGMbzRa8RE9xzNn5nWtnZsGogGkC7lvGrKrVl3snAz9RFi2yQ4Bs
E2Ew08dtLcuPJhftsDRMfdMpXdCAeAeji/H9hPUAUCdSJW/0tyJq7BVDWQQJMeQX
FQvIUjtS5uhA+MisnSKD+Kg85jogaBwCZvKYmaoUSbpL5aRl0LvjBBej7JWox9JS
aRyjln+XIE1WOv79I6kH2TEicq7sGWRh5RSwT4lTBxZkmP0y7f8DgLT4C921ASOM
bYNBBnewDdoHlNngPXpqgueEBDHwuvq5+OebpNFrMd1C8qKD2YIV1A1gV1I0RZBN
zBffaeImNKy7iEMFx/iQvsIjnNCYNVmnNSpJwj9S2dzKwLLmYf0eKTcWemcO1jRn
TczdUpXTL9tcRcvc5SoroKfEblHDx6ZiG2cm08KL8plVEnmITeLV0wMil8e37y7I
hace4G1YZr5Dpo1geTlOieZ0/mHRykygozKbRvgxBVR1XbGQUDWaxzMJVxcB9CDB
03fY47YeqNxvFaAJOIxOXzDmWpQIZx9sv+awmeZ+UbQYsvl2Y+zC0YUZ0SnJCUew
tpxxAjZpRJKtrlndF+OS7A6RK7jdtTjiQuVU4MW1IgyU/eGOseEoPzJpmoUoAwtD
g0T1Pk63LBdV4KHLM4OKNYIgn3W0FtVi8hP8LuLjPBGRGNRvAo9Ekivf35A7SRCg
p+ruu4cMuNScJgXNT/ZBbWqfhiXbKBBt8aEe1xrFCwoznw0W1IyUiCgz6LxtZfnV
7SDtEiVa/rhPhKZTRcvdgPNWvIq/7IXSuqN6or2qzL1BwVpRN1UbwYv1Qg6ibkgb
HR0PITWF3e+PAOMQevqnwkT3ERFWSwDoCWtSgXbxpESK+4YWBb+Coz6BfmAhQxGr
nbkGirS7nDREUWvrFrciyLOJuizhc4RBhajBWhPxdw3rMS7dOvM7wyNb3hR4HDeL
tcDBAKTzEsVAYFWMI9hx8TKspj8aRs7zWneu869UH9jmUMhD2m5q0XsbJ8dGo/Bi
7XMfaRaU4ZKZ7Zoo4T5oRT7e7/WnpZDS+w37yT+/xGBymLPjZ4kzaUWWNXfs4RhG
WRnqsccpR6WG4Z3E1tqZ0uqhq+tCZX4eqJ11RSri0K7y6I5zF/aT9GzxvZ2zwmrY
iJBBw1iowSGAyEhDr/XTImqUFYugvTdpQj+cVntqye0Xy4baeZBxodZbLHBHVTcH
Oerw/AtOOMILQxdobS1/OIkjHlNBVJqGG71PL3dGc31w8K7VscDnS1RybxLoiY5J
SB6TfU35TA0Jxv/+V+CCeCARPc+QbGS1YgThCzAV3Nyh9Mh4e7e/FBLqrkFq54tf
NWqcfIdZ9dDGbeeWW1hG5UUU+g0mpai7slhdJw70iZP86hI3ujkLJ5HI6NeWSPQN
M+pUj4tPqF87qYXonw5sfGHAsVOUu+Zbt1UTIKMQhZAZ/SD/sD9xsbI5cS7zlG/r
1wr4YiFyGLPBd6i7nKTf2pAXkWoTB9mYJf/piAoTC+PB6/d3BigvSkqo6y1X1DSn
bQsiLo0QeUbzR1GRLxktiGNA4dXnUvScL+B7F1WdKR//wKzYhgZpB66C3xKSCdOB
AVzrMlvZLKcWnXeitzahU0kEDQU+CvlzXsSm1R0wB8qYJZtRCoXv4jIy3eI1cju6
50FEV2lzrWBy7uTjoRlAYkaPJXWTBnO50sCiFKipDOV4Sa5Cf/IozxNvqjUeRwYB
+nMA4Y/CLm8PGD+jrW2u6YBdMqydrExq3HRcG7UICz9lvm8S4o2Se2ILyI2Afx/y
CHPn9Rimp9U8ckZDj1WJVqcaXaiPx13+XXHLuYouiGT20YFbxCKqWt5vGkzo60wp
RIRD8L9wHsmkoyQM8I/StP206BN31utotUszVbLBqhEMbGjcP7jcEMe3IeoB288G
kpIfb5OcqrCWe9dx0FvKjpAQqzwxuGDvTNtbMctkmijQkWAAebEBXHCsiw3j4MFw
hFDvoJc8D2irFmYXM11kUScNKBKrlmgarzwo1/11TMHkIo+T12fgz10qDVXeAEyy
+zvhHkFxTICxOPi/MN744ZPTDdmRRMCKVGuyxr7Ps7LtsjpNXd+boN6py8cn3cZ+
PSXy7Q5JCHTNCNRDxqLF0+wZl/ZMpionjVqiv0v60tRiU85mnmtYxZtcu7syf8CW
s0drTVWpF4LzXtof+KsaPikz3wOLjviLT5hfmXZGfpeeLc6K4ii7aZ7HDcc2ki9Y
qRyJQ9IH2MiwBiqp5nkm+GDCrG3tvooqn5ncH4ofF1YqoGtPrW0/8LDEWTnErAQM
tMcQNzxFCM0CkznNtS74yJlN/aBJ0AQrDCKGjPL1VdoiXA9qVJDYaOcfVzZVm2G8
HGoSiPoOK9YvK4yAUOr3dXklHJYw4JUn6l437KTznota7OwyDk5KiAYU6e3+jENl
CloZotztwaL9SkaS7YjT1ZJwR9A4BX+/QSb4li4Lw7wZ6E3qXXuXlw2B33aE9us0
mqF2dzg3UN4XRNiXyqeSVFLqdVUuhEbspNWRe7RK6dGmE/lIdsTxiz0J7iVySxpf
Z0hzxC/gxw9Cur6nk8zi055kYkFC8jMAz5fXEXiydwsAJZoueBKHzbTiuHnGSXM2
vTmkoqgdPJkPoGXGZ9I+f0F+Z0EagxeXtjjSFXS5o/CqCRZy31DmHDkod2dFlJdb
aw00eJg8VnYlJYvd0uyO+NMok2dKkTfXZy4cw0Uiq+xIbpRvMUhUeDXY62wHMpI0
KAmdIxmLJVIZZhrmYncEhH/YF1RG1/57VcpC+agVzF+N3sRD7Tnkra8hwZrYXDFg
ArC5q9MgdR9cmsvA3mWICK1xSvcD9p8qDhtAnJMoXBIuKszpadLhoO827P//UBTg
M43toR6lJaemw8EGSsKx31DsFltqFvJ9XyljykT3gIBeh/UHWFHl9B1OIHdGbEdK
ENuNTtqcTqzwK1znp1Js92EbguRcGU/y41G/SHT9N3yON/D+80SCitR6QMMPphWi
EDtj2VkGESXHLpxWbRz8DPRPyXVChvuD6p5H3hQ7R//h49TMRREKpJarcf9NaOsV
dvjhTkGyj3Q5UncK5TKAAoVxXJDl+8wIXkny3notxmlUrSFcgiq1nQcQrt2shk8E
yrUIebNPYGaSy4ozmoLlhgKdXh3gnzaMIDurrPYzDatvmzugKB4JuEM9G6P3+a8/
3027fOHoI5IzA3ZxTf3IbfNdzvgBdw8NIAJSvQ0YBYoN0AJTIh7Mu1P4JdtDHqe3
7WDzME/XNWig17sq7Y952TlmM+Cz/A2IDSnJJwjmG9yjeCsKL2y59tQuD5JSRZcU
4Y11h5+ceVlpAZtvieV1b90M2pmaKbrkYX52Gf8GxHh0YplKytulEQRbwcdLhwmU
cvWfWIR8rvTN3VeUMUJuFatmB4iT9mbflY0fFnqBY4kl2EXN1Ro/fmgSUbQAKhqo
JcFw5lHtYNdzYbRrYqZhpsygL3CfV1iRfmKB9OUxWl5rd8j2o2fVY8y1q106btzT
DZ9U6df/Wg2jNJRpGjrJPuFUw48aQdE9oXl0N989UpYtWBMTGA626au1r3TDdEEf
ROt/vLV6/kHytrJrohb0PoBhfO3QKxyUYSZVsOoFuaqVhLw7mPiq77cGZ2okGZgU
8ERuhvFH738YcYhvR40fDmM3AxSymqG6JMw2n+jofDN4tkmtfg8FuSnD5fvXq/pS
ut8vgQA3A9iEU5eucXaxvNk24wulxSGnSY1JQPwuEWyNu96lubAPXHzYcZlWwaek
wcUDwEwsTF7qtLdcD5SnrbREAGNpBfjGq+op1nH+n5oRCeOYXSODiyOhQicJsVpL
B40ipLvuHDYC2RT7W7qJXaUkcxFFbfvVMh0sgcUpCswZsvvJjuidtgq0NrmpUyF6
4ThAm8jveoLjN3Pcm/OmDPmjis9n/1VjPVJNXEGlBzlW1a6D1faztwhmCvNaXqiP
6T7sU7nIu2ydaA4yPxjolSosA48zLdJpnJoUhKA2tPCSXlTK50jw5XK1OptJvFKW
8766d6XwULtNsCYAJBRppBzNwGhwTNVTpH6OwjsjP0Bdtqz8qUk9ARMzLkdLyFH6
8/EEJLvG5DBJOeh+ixGrnTedK65+q40zzqrUP8IvPzEqjBFCDSwgLWqEFmDxwO01
42cuRgTP0D93Y++lfumUcnYtncUvkAcEVMTzesSKa7FyfPGw/iJwsMTep2KFwE3c
XORkKaPGO1A9eIghRVnSC+ieXdox7yjnuXSOEAfhVubkCmqBIzuiDJ0TGhooQTyH
WYN8adkS567v33BM0LBNytiNzjIdPcEn17saLgxIMAAjk42dF/03MyCKu6NQCdVY
6Fw43dVsAAIUEC2UYEMYJpaIdUmpJFgBXSoeWHFI7+ysRgHoIYt3sJgPN+Rxe/CZ
IR7qC9ivbseTFypXEpK2mctK3tQrsW/2Pp07MxosozYaWh45xIQTyW2OXmxFlHnf
lxhk8K/2kIHKdl9SCT5U1wbU6Xzl6ySIxyCTAuHrXX8Qga1kqQCKi2CXynkQjycz
OPsZM1EVQCyPNzUEDpsdnAQRD45fJG8U5VkHJ8gY7aH+qyuY99BnLYkwJcEiT8J2
ZdDo5e3EHBWGKKmjLNHQpPJuHlMCWM3YTKDKZVjx/8w=
`protect END_PROTECTED
