`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sDrmomHThmaXvMDhSC4EDFSu6k2OplhMy5rDRhurNEZoNaYt1X0gctlavkfLesWt
TpFZnmimOD8yCHfbXWNZ9LKQTzCknulN3SYWYCbmwshg2aeEPuHl+joORGWshn0v
UQLFUCxt4n28yhZ2PnL/enRInt3dkSRCyJeckpjqQFPjIbRbBFhdiMFYHArvboaN
NTNZsxoCRfaWpwH0ZHMQX7MP7hmTBuY6AYALEHpMVgpuFnlfb1JBH+dEg+xFL2hU
NnV181MOTw7dfL17N5ZJMs8rZUky1G68FD5SxL+k3LBGVRs9efJzP394f1Zy+uCr
VU2Qz09ZvVo5S7A0T5CmmgMHp/u2jgDM/gant0YOOj4iQVhRCgwUqR7T5iupb5q8
4NikGmqE1pEfsmZ2r4asbA==
`protect END_PROTECTED
