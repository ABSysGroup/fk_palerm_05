`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
869Yd9s7M5+UVyaQ2Z1l51W7mmK2edHxZAhvpTXQwP7QwqrzH2Xnv/1omLk5qlBx
5AoQgVWvZ7bA4jqBPUgWn5NUFGPmnETtlSiA8c4OQ/2yJh4+7Y/NDoTR4cmY/01J
qd2HEPGkKKV2Y4D8HqGcrpaXzYi99Oz0Vh0RyCM++wdq8VKAjueLW8uPp45zT2ht
AY0g0umyE66bqu0ychNZCL+Z6hZ3vEbZ/huk0GK8LZI+QmX2/XnQUhRbJUOdtQne
KHXJx2yANEJ2jrwokanve0GOVwuk4EAK+I9Y4c4bsCyw1IygDYAG3SQTmxSZXgXX
f67O13El0tNySBfAf4wbFtG2QkpUvcOTIj2eqqvibU/m8Vq6wbb10e61uUG4JLlz
yPm9x5+vzM1ztYef42qXpHeerlaF3CAe/1EWHj/f1Tg+yQFMVqzaX7KdbLBg0IDW
Ob/HUZXEFsCly9G10Yix2Q==
`protect END_PROTECTED
