`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AleBfcPp6cPFpzGQ2WRv+REModxvfgKKbTO3FmE6AFZWmTxdZabcNDTk3kgcuJem
zsdgFMX07ogKvjTCdJVpjJWIW2+cFM4VFftcUM133C78A9CBvCsXfA5hM8x9zRym
3lIHs8cHICv2rhtGZf4jocidGmIjMjZLUyBlWF0L5WDFBFF4fGXzghd/g5Tykv4o
L4uXWklteJ1HI3tQADbKzrXqsrHFm8Uq0Bsw1vyeINIduFNyPCAD64dOrZoloOHh
q82pXfr6ILWs7ane6nMuSPmSF/WF6zmqK5w4yi1Vs68vXLHieKxo3tJU7XJXFDfy
lnPxJ2J9KOMs8bHkwrEKy3HE3GvA86+60FZlO9Rupr6DhvgeziVfxXhWrjGMRvgw
2RZrcfy4RbOxls2/iB3XatkIQvBzh4S9q4NamvsUYOSKTjjBy7YeuEaNu4I47rAJ
dDbW5Pg3pV5D2+ba56RigKGHT5DRGhKVRHigFlyW0lSAL6kaIOkkKPiERRm2ObBK
`protect END_PROTECTED
