`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sCehYI2Bxf9nB0QwhHiSHJue3gFNMiwQsGBAI4mZiZRD+V/twc6Giv9NT3h1stO0
5Iq0CkAJcKswohZAvkPpHFPGfKZ3+aD1mEJO7mjQBos5RlOQMjPyVd5soK3Dwzat
lVcUdRIACVfS4thDapFY15epR0GZyTOZ6a+8z7hk76bPYdBwPYQEaNrZU3Q/WAoe
5IYInulMpdv/HXbXKr/EtUHH4RMbVeoBGLi6QNDAiN4hm0nVkbRSW2jYu5qOEfPk
n91FcjXaeboWgkq2zJNqhROwZtI+TPbmkq9ls1HoLV6SDwRW6Ab57U33TmAHXt3q
kEwXEE/tpv9eaa1diG/8lzvbOw52rM01+kOK8N0r9sPxOC6abWi4aOCYuPrZdQRQ
yBXyPLGOOc5ncgPzfcPWBnWd8XFFiE12GPHegUIHLHq4N/MRGW0CCoK1mzwXsUU2
VCgYqZ58HHkE9CeXMFRZH9BNvPN0gGJnozQJRa8vUQkpSugrhrbCOYdxD/f3vijG
ustlIVVq/K/YZBqN6CtgEcv7STvJqlNkYHWU1o4pBOPFo0vXs59GJlLuhT4/eorE
TB09XoBgUTR9mp11Lr4O9GrlT69mv0xPOirkfyFCe9xFtAbyHiFM9rtKvU0U5tP0
9OKUVOKt450WyCtiOvSE1nWGCIqmOphEUtTMNCEq6kUqwUahqxmNOAwSiVSJeaJc
cm0yr/7W8cDjZtrqz4Q1XTVle6oI5g1sUp0mzedF1GtHl26Z/N/hqzY+3E0g9wtH
dNhd+AKhNPaggXk6mZkHefg1+3qIveotv/6LHQMw5u7ApzPS52SOYjEQOQDmjxP2
c21Fw0Jvkqw9fj3iCH/KA9nPnyse0GhU2J30hh2oIbGmOS5huuqvsVK6fF2MzOTX
lz0mWxzfFLuAlOIBxCQ3LalFF234H5MnnPWunqiLS/CYWBIDrq31d78FGdPHbIMK
OxxzNY+Uu76nZaCKDQ9BWDUll2unLgAjEKwg1uztUeWBShktGlwNdqLz2K+FXchV
kH/I2Pd0ogdgjaQo7AebiMTEIt8KZigMVIW5tHjPUu5e9rkq5IDjJDtHAkT5UoBP
4UVO5lfWJRtCcYbH7pUv+i3xftiV/n8oiaU1463HqUY452yRwxkA9Gpt5NKWuHux
tl0WeRk/4y5di2wywxMIbuCt/EYBHgzlSF5WXn9rs0fr6wod+ohEbY3V1XKtrw01
J4hQ/8scrCoiaeDObk3gLd3TRmkBL5YqDrgk0KqowHwgc586D4gD99ZwiEzr0JVo
pz5o6dGDyHssIsD0YTly3gtu2oPagwrX2ySYKRFoSRmDfWQxVulkwsUx5l8oV4dE
CmmG/g6/5XG9ZJnjuXpJo7487a7l+ImISaRsOM0FEpEbNUAQnykSH8ZeV2tNgkeM
jOv1WMPm7PFElMiHqUYwGcTfAlW7AobuOTkBGkhITWGBJdASYNrx8QSR4qtiO8ki
0BVhgvXf7NcUaSKE55T6qa6Aq/nbe3yBg8Rdq9rrmwhzzUcInRPypAqJlbZxMuUp
jwYEtpjiD9yYrNPSfA6SyL620SnURqLcG1ga6l4POtuFSAS97BmmX28O9w7MyE6z
0BcdCszaW8+lAMUy9XHRH0KGOz4+rMXZwFc9ZXpEfqybQe4CyFLVGPi/la5JRkw1
ICNvM5yxVwOMB6mS8TzucMf6/E/R5EDODcg4wTuOOAuMBOZv55x2zrnJ3NgGrtOW
xoFkmLN4KcqvHhsm+/vDpRiIJ7lIo4cB/Xoy3VG2OmttsRn2gi2OmexTpzUmts7j
oepnYiaqotAmjlGnKk0qeIHK1isC/8+OChYu2wzJj/ZHGmf9ZAEyXESuBpVu6bMU
XyJqZAwzqbJbH1co0QezoX8vr7lpmuJwDkEQEtLHKMTZqUA2LjkAPln4bYktPdhl
JR+lGxGrW3JPyT16zxBIDU4qKZnYIbpRDOflHFDvKrz1K/A+L5rbLCWbZhw/YNOb
rjQsoXG4aneJ6ACI7CyBvHYQNspmk1CqnyeXH2pptg95V/UX7HRXIawfsTs8Z8KO
t4uF265KilOYTB+ZQMlxtL5FRK9cI42LpWlgSfVoQiVCMm7k6sit9kPL8DK2mCUQ
YNSHJkDGonN6P2Wmwo19esBM8h6p0huIRBUu0fw8JHdh4MTnkhYLyCJ+S4BzLYUd
m2V41R4eSz/o0amleEPQBwt9v4CxrzJKPbigXfxHHTV0g3i1aceHzuZ891kgZH3g
SMpt1yeMOz9kwqQpC/B2ZqIhp4DvxFEPwa+OpZ7UpP1x7cVwxEkme8ClkvhlrYhO
RFblECV5LNLfzXmdT2j/QlVdM3O4mNK+BbDUKRXlUnJLkjtTmuUQLn1Z2gxWYnBw
3V1vjcbYUKvoIh8XhrbAtnh/1ypRWcMqfyWqYPAD2263Gd0LaLWWML2CmD3c6sEI
3w3AXEpyfyknC0yFWzvx2/sqkpVCz7rSdoCsKMHvQu+e4UuDUQWxgyQ4iXu8Cn0Y
h+3091kBB24wkaLKmvIfS6ToTlrCgQUbGGur4+ZQEITcn2IZEAstUbTqfQJqSzx9
hL/o8PFXLmDiLPP6vhxV1mz4oUJrYQVMz0HtVE8GzxIGpWojHHgS9tR+R2Q2vuTT
BusLX+lvEHdkv9qTGy+qmJoLpiMkpV5mzvG818BqyuiMeKh1FfA8yF7gp6lC2vZG
+PExl5CR+ElB7s9DzBcVITjhpmQao7KKT5IwV+C23tmNTfVjUoB+x/8gnFGfvbQg
vJbnV6wqu4n//5QG2FWuHZMhfe9pN+oY8jJTEUhBNDH97oLIfQ3u7EQV+aNm2JXK
t2NDl8HhRsIN86fPQQ+mjG3c9gG7734c+vJ/88jdR4p2Q4J8HUsfjljaA0D0CWPY
fLLxrI9pFZVOi91kupUwIxFKPNZ58lIRzy9KGJvdJfP+CN3P8IiepjIL8uelPSHY
Uc/sLgcLjcN3KLe/bOp9nn4zISGgktvYlxU3Ldz4iF7zs1StGoKLHjyor1WhpN+n
JIhk4qGh8sJ66FqSijB7d00DpPzjSPMJOZE3qIdJFJlKdl1lctqYx1LM7FkUZewl
MQgXW5ZhcXmLE4qn1+tbLzMZAz6H7JVi/IvslsxcKTnS6WH01/X8HOk9TTseyx0H
+NHS1F3CWTxHFD+8L+gJs/nMPfA0IH3VShgb5B9eqaERUUu7S96CvvZ9eSrJ3Pka
1U48B0bPdfm7uKyJ7n92Yg4tnf6L32hNg0NQpO1YaRUHVllhIgMKOGHjzDOTrDO8
fTHxR1tEsCc0j1aE2wXkupnalL27E8F2jwZXaKBDzBHqQj4XDLxapq8+yHi5ZT3B
U0COvXQC7MwWOBNFDFKZapEPmK4n6cNa2+likbNGthn1Z6ScsjRagRHvQVN3yiEz
tCigNDeXGFQhwdaeSaL/idn9J+/dCXEHs6KuiBJeEekqEGjPSpzL8Utt7yTvei4Z
7caQfLXtUgvyZVARQ86Wj0hgZxhw4YFrQxJ59dv/rO+xgt50mjdCtt1+j+HkGmH0
hzG6QOo04KkarvAk6ZurqKWvX88hV0aSytAIYWrK9bK/LWDn1T3k0XdFzWwc+5Y8
KcgMhErswcNhHXAitZPdWF+q2STYhdUflUxxGR7QQO+tIDwprlBN9Gp3BBlXXFug
AliRLzeO4bVPtWC9TNiPWlTmgwA9vhG24V/98uVrx52JFoSmtGlrhhZBQEiLrr+3
uyKValgEaqfxxug5Mg/vBWKJYKd7xsGhEhiBpCxwGqn4ex2LSSrbe48xKIKJR1OK
OYvxkXIQ+zVn9TBBNIAG4Sh3nVm62xrP0ewxodhtoDE+BwEHw3pqOlTX9DziEimp
d+5l0gDIra9CUYupQkZeNw6HbXlyef6X8h8A0UQ7Qzpqxn5+2JSOJLmC1dWqMNkz
8dLOJacRfb7LnwWNMqhUilNPz24TD8DBIkkT3XseeugIipfdq4gVmeGjp1OKaCl9
lNtmiQLXq1qTY51HIzYaHU7yjOVkcWEqX0+pvhjubk6uiNYF6ZKtGsMSthWCMdSV
PYcX3dfLgrMAqZqvqKTsnStQN16Qw4k5eoyY/UO9xYnMXPqyQzCeD3Yk9TSnpIqw
e0Gu/5CqTFCuRUJGdxOu/q+5b//WxUFXPlhdTjLu/g7/Oomn1SBASrPz1WBiJHT2
rMtQ1FyzLc9D+wxkxKaCVgIVao9YAiwU7llGTrz2bnyO0+I9NCOwXFmp1YoIuDGO
x9IrF5h2+xAKPp4V8eafr98eL2UZqgAdo95xBCYza7vi8JSDGs/hbsaJ9yXRei8d
AQUlA9sqG+wd445Kz9Hw/SWegjq/Whc44kvUMe9RZAdR+sHLjqx82Q2+CC0AnwO9
jTcOBP8GyNArwTjU5myEaQNgvtbDNg0K5aDfdIFZwqlJb7LR/MhggDxSXzA02zAO
c9HI7jip6E02bXKIykxTf7QaGvEr72AybZ38WefhSv8ZGoqpJnwIyvC36HCmmKnf
lxXldObJmAGItpcMMqz+s+D7YUV+ovEp2iwWHesqqyk=
`protect END_PROTECTED
