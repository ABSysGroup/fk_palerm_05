`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sxlo0UB+Wos4OidW1fsq0E35WCku4VszHyhVBmS+2p4sOLG2UYgSHJb2b81+5t3E
lzsSEvP6/NR4k0+f7ZQhXlX+DffM/a2Ohpe2qzuLmDBHHPXW34L3hxW4+HvekWhH
mOGFvwydm2d8QwEOxSXhqOtzAGtU08+G2oySc97lSYqbuKcY7oN+D5fLLVmBK0c/
qRXw0EtzlrIv3AZgFyPN/gZ/RRcXaCRmAr3IrJcVGM8+3ywCzJJcizcP01WrncGP
3w/UabebIz35tD6UIPWBclxA9hBl9bXZC4Fwu2cbJ/a8+lLzwEh4iv9q0ahKD3vA
QOZtDFDpqmz6CBI1i+5mOg==
`protect END_PROTECTED
