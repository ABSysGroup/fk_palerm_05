`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dv3etZtYAGx+OkEljcdqlPTUAttpKP/EZSj3kyP3SV8rhg7s53pGSPREBJc9CpOX
WNpAcqJlsw8Cg+vZJd4bMbuSXmJfX659M0vnEZqkjhCCnC91Upgv50kmWSS/P+nn
j/5nK5NeMnD9mv1xiY2ETeQwXjWox0yA5EYHgJnW6aMCZ7JlvMJJuDVvb1v7J8sP
BBny1AXgaq6IziD5u6wl83I2mtbGFJH5kF7xUfeaqw5T2/C9oH2qtxYQa8SLxu2k
gtjltt3ce6fwSQcprAqAuzCAl/6ZacFF12/N6qLqlVqqUsijrtE9kttyRxTJv1Ov
9q0SzFIajUlWFqJC6yX47oIp6PRyVVjr7lOYQF6X/ENKW/Okom04YVKnn5UJlGTI
lkRV6//DcVxXb/adI4sbguCS/FCxT1NioFgDyK0VjCOoBXfoDw0pfX2QzHBbU1Bg
jk9Sc2RRxPDPK9SD49jZku+w6Qy8zMNY2LlIM0u6ylcCtu/UROzUKQh6FdMltL0F
SeQcUl4JuqwrO8uA7q3h2Zjx3b2oWa8UtJiOhUfGirxKW2NXBt4uuDfNrZOTlLGg
kstcB6eS26Sy9rLRnnpLOaQ2gJu1cps2vh+MomomAcEYasQX33sZW0hVJIA+zPRx
3MJsiuxOdTDZrem6NWfraFamtiOUnnPJPaIe+gJBoI99zUNLdcr+VLViaHeAxiBb
XA+ZHuE32UQOwDDzG/KYhtq4QznTrAb14oPVq7dmRE+kqzyjdk9+hcsg2W9i5wsC
RZbNbWlyVZXe5yEygTgI4e0HRPSQFzLxdyGXATlXx0Ev+jFw7ghSw+NjJ9KL3wss
01WAhGpDW3oGPXGmEJ0QyA==
`protect END_PROTECTED
