`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TAZscr/e5K/ZMYfXNsf+2wnlqFHoRz9r8LWky8gy8eUA6QV/BAjN9OEDt6KJN8V1
8bLm6/ko23Qwi2WIr32lKCC/GVrh3DEajbGvtY2iZ4DAvRwK2u+ydBsY3sYKD84G
jUTz6M2iFBtd357Ig/SKtsBoG3/aUFef6793O/WZMYkj5CiBpgnK0hjcjzRxNW/i
GT9JE+sDqT9WkNvcVGH4vDX0UiBfQv9kQdn2NOBoO09oqawR9mB6N0mbakoTw01H
iKAGhx8iugslVXlXNIIk5qXbWBldm40NbefmrsxF0zjpKOortrLsyiGkfS5A0JXX
p7YJOvxsRuE2oL+vevnQenXw3YPmuWUAqLRo1LF06wz+HHaqL0wSuBMltWZ/pCpS
8ZiA5E9DATRUpaHzPsNdocgl8LyHr+TwObPEXTan+DiskVSyM9Fh2u40cvxBVNyQ
BYrj98LbtH7eU7Ip6RUJWNaqFE5XIzxSR44ZzKJ6i91WvjWfHNcuW61Y8wv2zTN5
Kg4v0FjzZtGp9cHr9hQEx8o64mwM9pIbj3dK3iuARZFyeHbGmZ+YFIruMeYngIlD
CLF8kAgtD++6mCJ1Aye3wb30p1mBDHaOzRQ3BUuibPGAL4XJlwXMKsbhyRaSw394
Sn3oomS2Cn+tG3q1h5adQZbtf85ICwj3jLf3ONTDOa4RrvcNTC1TA2fIAERVqJLi
MyrWXqJEZ2KdCbgIZIHXFp+RXuCEpVlfDLmWnD96vu5xsNDawwenahdVGIHQoORd
8HlbPvUlDxlrkdqZ8j+5U9G0LouOfzYT+KzL3Z0VJVKEyKp9wecEj0NiGjeH1J2C
DzkUopiCKjcHqEXsNGOE8ZsqoKZHOWbBttRk3Wax6WGszqwXzD3VEdFhs9sKaDue
`protect END_PROTECTED
