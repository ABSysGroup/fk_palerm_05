`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6HDyfBz/ksxVlapmvkLkXN0D4G9zfyLAHLyiAIJKSQUQ/HPMMRKnqTnDB2sh555A
BTxgl1t4ryVnpIGxRSfqnyY2nKNFHYki/26yxnOOBpf2PrHjP6iqFrCoGY9fQAJS
LSuzYiQlp+FxACrH9oHl9e1/32qp2xnDgp/XTqbdlzp/8dmQRSd/bWgVJhZmDC3L
oAnPxKtKtkpThZ5NZEfKpqPSUL+SbK/+AuVnRbSDyhfiJpoF+2NOuP4nNRXEBJT4
UXkRN+acMo1RBYtuwhJNGAaGleWfLlkInpWqdr4cOjuX0TCFN0U+3bBZVB3RkHVa
x1WuVA87wYHKgWi4iXkRJBb/9s0tiJflsAn/4bYMUxfesOpoJxRCYq6dwMaZOwCe
gh/f5tEzk1f5sNOm78HjT7yZzeUa1+Fsonljf2KFFadCa3A+g39graSz6giT2IRn
bBGdbXjPVzvkEUCHT5tIP3gFsC9Opld1GkKED3wacwUaeDa1IdgHZ4beaelwvSwa
WCxfH4hjI7r+RVPfjze+NXH/xUtfxVscXWpC5wcZqsS8h0RIidmLBLDcjurkyCcN
zCU2KZ4PC10fZWxayKrUtuFq3Q+qbHxj2t+UTa1N9ykHes+Ept6zqDTWVv9JUzWb
GonczDVsWUgzTnnD1XXKfOwIQibf/we68wsWMR9cWs/hlbqWEWjxjiiSeMkMZxvd
p2WpPx9szBmVvCSJZYMMbDaXWe13RiDK+eMWoqL2zszcFlRqCnwZ8Kid3vpojdDR
v/i/MauFTDz5mkR2bd315AuPzIE68TlX0RYHl6CDhQJc/1CkEcx6H9Oih+guqxic
nuF94+7r8as7kSWAwERnyaB8jUznttWRkdZuvi7uWsPYDqWpDIj4nB9Cd2PY4qDL
gJ7Es5U/wSY5me1XD/2hp0FFwCiE5VA8E1UcoJOiphElLEJOCyrhtVyyuffU/sn8
enybf5QfOKaQJxB3cdT4IFFFcdcbQavj4D40OPFk3qhhsqbsWjs0mTdhGjQdflCo
b9YEeuC6rE2BXAuWpesWAClg/093+XRoVqMguaGlB0lnIr5gAjzs5MIwUBNGD1oj
dQWj2i4RfZ29Aw9GPf7mZAovDVhvrbnB8cjDqFHExGFnqAqYQpxA0wBa+6LksX31
fVAp0ebQomEmiHVX8WcSXrUsdk12igxTjGEDeeKZiyf6XHBV9GkzKTfnpvapWPQr
gmvzUMr/dv9dzh3Q23GrCgkxD1K6Y5G5pyP7du/xcgVAy3s3WH12Rcq5IDtbiQ8H
c3YSZ4uzQRdvuvS4unbJIsa3mkIb3UzLk2MrjHL1TqKbQDIHDuyHLBayLhJzBxYv
xITUQjC87T3/BNidIh5wr86kW5w69o+jlAvFPNwiK7yhWth+5mxrS6xVtJGj8ozb
t8bG5mPjR76gMP3mrDjqvXvkadNcmePqRKV5JPyB+jchnEaWUcMczL/48unS/2T2
B9EwYqblCU7aI5aVuueMhfKCQwD4poxuVv1tUK+dBIv+1jmesCA43ZMMCMt0kuRa
jBaCo9msTP/U+YBRXsRJ7VVQPKVAhjGNxW4yUkJequ65AQ7lOSznxbHHsaczxnr9
FoFTAmEfrNCxcRutGiA93B7KGWJdzQAKA3x9oznyGqANcA+hIiHzCJ/dsZon8RDs
FePcxzdLWA1g8Y8k07k3Jn9mai6mB2cpOlJ1Vp6QR+uEGwNPl387Ryp5GL4YJpnW
C1IsAcgjLXrwJ2gsxYWEiXAowHmg5tCr+4IvQHuCfvN2LMguY2KOgBmGWEc5NRKK
HF4nf13pnvj9q18NPq6C0cpkL3q4d2v/suC0R/xkXRhK7g917DvKKLDk4XpjN0YD
PT8k+O+t+1jxU8xNadZvLAkkxuVMCOmseadUZy7b0JO4FC7oUNTeCO09o13xhleo
n7pddJI/Vs018qciPQ7YYurcQTFWQs2nKPv3L3I4fcpRZcGGlZSJTTSO5L40gtUf
/elDcL/WpoHMPNrGlTFjYbgAePICI5q4LSwuJhKtrQHzR+NoQuH8lAcp+KcWjSjB
BRvqzfCwc6A4rffmXFNKyw0iHadbV4advqJ+mH1vBlE+W9FuJLt7i5MRrHcfDU+d
ht3QRhrN7cvcWZE+HgKtRrAl4sRGFIkzkrq1FEti+Z55EZkrw8zh01p8tYXiVPdu
KN8+dr5u8WL3hioGowON8q1O/E4VqFGRkGDWGADkc2Pc3Mi8i5alipq8oqUk7kMJ
hrZBl9kZPRDcXL4s6WX6v7alTPopaWV1O6nwJ5UM8iDwttD93ZJZ4Colla4rd2y4
s1fcam28x2FX8Fpq/wVZDqoJaFCoOttipqHKQg415mhiYXD9MnsxcfzOL2DncxrA
zjRzLzVY4c9B3VRN0CCgJMb2EaV4e/mhuX+++kkVj3zKY9ovVH9rOvLDdiWYk/fK
0Rx4X8+zWkCPSkhGVO9PAWL60j4IpCe2Vn0e/aceaFsSqL/VVJmw4T0HkjmdjfWz
bThMB+h7uOsBiSYOOhuKmELg9G8tffbOjhRz4HzCAbpIKjyB2lYyWE8P2udAR+pm
qFdvnaMVmzqa5AzR/qQLhnloY+rYtO+wuFHY1ToYXmZs0uEFZ+pBprNk4qibrYGy
YyrmWWFUgUfUVQGpukcN14e1PE/TtN8KuVBY8xftO6sJZAhUbRfOtodbcQAkH+aC
FnVZoStfnbeEbtlixbAX+0780MglObLdYFiuUJhMmJDEMAL991HRAbjAB0j1XD7p
P94R4wFb0f9UamHQRS8lrXRcsALgJaREsB7bft+vezVv8fj5gdU81dVR6bU3wEW0
yuswZ/NAkwPOMU/AnkqUsg==
`protect END_PROTECTED
