`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2oOIzGk2JW05WbknizhqXRVL/AyErbH1SPZA11Vb6rt3iff08q09x0P726k0J24X
ORn1Ks2D+qxQ3TSTj/EwHNrIDvLOy91mC+ZNp+qzWSBo9cDv0WNvu2dAIoJTDjgm
Xs98qYCHNHiEhYkjKMEyyAIPAyDsuGSEHWQUavRBPLamfhBB/11yS9UVD0t5TDPR
i47nqFVXkbCTOJSaoQuAeQXjcPOhUTMQRgeTN/AazvK7IikgjJSu8bOJYKJn+5fR
TUmSxNJEqo4WK5RqspyyvRkTcytQJEmHrZhoONHxSk0KG0k5G9CsBbVdtApg1vLY
UpH4XyEmkAcwpCsIIv2J1JYJLA+5IXklJnB49Fxb92YTGTq17AEnlfONOovtp2Pq
hGNsiaDBbEemKqbXNiG7eSE5wySZNCLcJ79XCJmKNcIJJFZXYLHHwMNIeAXUytrV
aykY/3jZ0+4CcBP2HaiSGrWtsVv3JpQ6LLTYSbhMAUT2fKWNdCSAJv0KfGeIMu5R
oUjWrc9TizSO0w4CeYlKcjOj8cFjKUYpjNCuLCE5N6wljn++HHON/A+tH42sFc3d
L+uQw41xpPrIVAjUTSRbRau2mh8SEwX7OvezSQ1K8bo=
`protect END_PROTECTED
