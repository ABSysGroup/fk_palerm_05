`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dM3vFPxZyc16nLW6DVa7OvBvb7xNwdPtFyImubH0u/7JfCF0MlvZL6dZdWv31YTE
W3JZPnvUGeOi1BHBRSRydTIexudlUtsN9HISuaaPvmG8xS19SkOG0CH91v3N7Tkn
axtO4oyYFel58rqFqpzfHHVNQSbxJrIMRNLHfoakw9w4P1QH3PKQj+6CGGbU0szl
PIyrJbq1OGA/ugJEh/a0+KKYLjI7+7o4HT+5WAUltPS9+tYWeLdhC7fIKCL7IFoa
AefH4dkJw/1RqKrfEGAW8Uu/8NvrutLTighQrJL0Mt0TIzcuUHSUagucODuKAk1k
rM5BrtB4WE7OTl96q2BmbUEYeQq9fGm5qYQpciJYJrN1CeIttB6HL6/0XzZW4Bci
hTUkkxR8Wy8dpY2dIlFYv0+r8iyD6JnG1SYGkMuZyiw2+zSXS8iMEtqSMFrNSfOr
+dIzii0jbATEOkQtHw55fvJmv6wI3V/sG15vGuRdhmvmFpdGNVrsplWsrtyxG7RN
CygQ1vxNfLhmB+aS4sXTkagD3fDv3NTKLbKPlErbQxGTdHo7fxeLVUxgPyp2VZZE
`protect END_PROTECTED
