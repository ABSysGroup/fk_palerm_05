`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
beaROUPsoIiGRQoSlWXw873JU/8GxdicAhIXS4rxjPVPMo4vUABgov/EkLfeq+pB
epr/iV9/PJPwps+IxNSxEzickF6pn7Or+Uz/pa/TUUBP0treIU2w8aRUqK7ZGYxv
lO32qG0QIgMbpXUl5PnrB2aOUjBM7BxgGhgnDzK4pCUSt6IZ4x/aODvNRUt1bEP1
Z5RHO/rWnMgXWID1MPWhKGQmxSG4pJo27TBKh1gf6B34oopSEnUVwbnZicRyZJzw
4V8WsSxsLe4It7EyrOOpBzpBGB1HC5sP8ud1O0rCt9nkoSpk7vyMogKiAjDhVxCn
mTgZ0hepVhpijFNZ+Z/0v6qUKmifrx2gsTulfujg8OIxDVDVAZM2orgl+4F4H1q8
`protect END_PROTECTED
