`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eW0z61takepNJrAd/cHrTdB4CECHXkULHJkV3rILTTfhWbjlGZpEgGxw1wfjRRa5
70ZpxcJe4Q7H6omee4e13fuQwhy/lSE7cK8jAwVbvdqDYF3M85I5HotQPW4xXrDx
xQEdqkEDxs0t+uSuGhoyAyjhyZGP88w59wjSTJyuPcbBTPxZIE5bia4Ryr0lUYlb
VeBij6JrXKsSEc75MEbp20sft8mCAC/+21DYGaNDl2BAMvmhBjFvafXFOejUEhnX
VK427wGOYo4LmkIG4k4ISyNqtiZOlLAqBWL+kb4FRdBU0cZel+FuFZtb5y0z+iZO
sq5tsapJpAB5FfLKPXnXvqLxUtr+52g0nUzXW6zOfUwFosJpvolkGmhhY8khwXDV
kLzW3AAeYy90xpNySfMjXoTsTDRNXl5bneIwQERHQT7xqG5m/+ThsRPX1W5QwDJE
+4fhgN8wEEWwFn9ZzYf3V6yQWHUNdhV8IiT0kLCeIAmylTKRF3HI0TG+kUDn8EgN
sPWwVSQB8VThdsLAHs3KWyINim3d5OCMYwLqPCwgrzmTstRvdy9WfBW3XsFn8EnY
5MblYbltnWkHqstvWoFesc8ZbMfPpY7gqxzOpEIHcUjSy+2j0cLzf3B895+IrUOB
wy+X4BOA/ERZOXk41pjFMp9uoQWubGGWPNqJakyscZmP5YVzY8+zvnfSElU8suSb
5Ev0dM1dlqu7906SV8+kdwdqaDZfNRvj7HtHduJuDpmULvjq4Tp0QH0u62W3Wf+d
X/N8N7hklGoqnlUR/OGSRHHtu+rxL4Y1krC8L1TCY0vtmcT4XBlXlOcgsrpXsdum
8/BU0l89sPv6PTkcsogCRArkjr0rC+0NJbZi5s38ZRE=
`protect END_PROTECTED
