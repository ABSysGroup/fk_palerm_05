`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YbAGEyeSacWaXwcGg5Ap6hj7XiHlo24gfbvVfndtD3dlqzshxpq83O+nIynazKFB
WlX1Vc2bwr0RsYdSY2ckLrTEjsb15vw7+mNQAgru3UjiZ24gzUXEPZKhiRyx4YVc
eEtXPH9rezX6KU5AMphdFautPtuNsDfJ/0+lRluqDV3HrWqyhE0rvBfmTjRGrk8n
zBHzMBxUqWasuoqmcuHKO6D04Q1znq36TYCPUQFOrBZWhMOfTxy9r3p09wR3xb4q
vrCQUO5AzW3dGxbTofl1IgMsfxze8z6LG0tLplVl6FG5Nikl5Vlb3/DZr4PIvzR3
Yy8mSwbwSDRdbxp4nTa7M9qRdbdxmYrosjQAW7RugZuosY5OGD/XvJc9Z2hm6Kpg
woGi4u7ki0RLoxnNh7XHY3G87ZtvIeTMoRFyJOz4ofk6XdH/ev2+p2Eb3cpO6+61
OjH+rUy/aDfJfnF/QDG3MITLHQyyxE+r87ewR5mFfmDPqn6s4QLoIuv39rDVvy1t
`protect END_PROTECTED
