`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7HQiQlLMSyNFqFqsHGyRUm/Dy97wrNp0UMBrpH334Hg5iinubqe7MaHjNjB2kU9u
wjqFsPni2ehIAuVBmRvPbaJIwYOsjJMO2OEbgN9nko4IH5wgzHunrdWxzs8LWAXu
uEGVXj6A9lIPVlLwqla0YjOftW79Nts1wWVl6iH9TUugn5i8Exll1gmfkX50go/T
+JYZhn6ojOKGGkKQ8Phov+Jk900lRpPKZlOLhXnIv1XAe/WlPSqNk1OQjuCSRYB5
AKX+ffk5GAO4SI0zw5/7qbSw3r1nSIk8jUxPeZ/len91viK9P3nn7xUlV0/OR+oj
4xMpzHhPAz3XcjBJWLILoMwna/s6ocz4xXnsGCQ+S7H9kPq6sFGOAziIFmJ187Oe
cf/iZpGgDgPAlRUw3j60Xwtnk77PwMsL++BzsJtorJwxagiNWOXC06IvC6wIHsFR
ToRkDQxgMTb3o8S+/HjHyujvE2phX9YE+MJDm0kDaEyMDjDym8wKPt6U6/KY5E5x
kyk/CwcumkA+R5IvHzOOcJyzYEAqpksldRIWosdPgvTw6MhsPcerBLzRNFcYBcPI
5GAWSDl+Fgz1dmubz2Ux4oGmnCdvth7qR8IXVA+jEw6PmGvnoaqMIIGOhTyW9ZQH
brYrRpACVqyF7P1pv8sWrBAl4zN4Mqec9KeaBzFWjUT9l9wR3dJe1iZq7yMgEiYY
nPHVC217HBRwONsk8tYBehHCAmuLeOHPBkp85goWc8zzImbqwBybf/vRo8XW5c+j
+AFk7nmVEzX2lZFWZk6EbfsV7aXaxnuWYMsq+azChPt0fAnytyb9Urzz5MMfdzbu
it+WAZA2nMqESdlleffGKmbsd3xIxuZvQ5lC/0SUIRDKqmmcqiMdGAz+MO9AY1F5
1DC/MIsra3e1+12k6JG/JBWjEP8Gpw7Z0XnMcQChTD6elOqWdz80yMF+4f4fS0hi
CM/vLPf+m+uZGxw/oGa/rp8VHSGlT4tqv97vKlEtz6PWMbGell1wagAjiBI60t0q
+jl+ikK/7Z4LqNVxRYtgx2OLaG8WN7LV/xU9KvylUSO5ChuIwvoQWEhoUyi0bMli
CVVJdk3xmKY9Qg4iwvQPhAej0/2rsg6lc6X4sLMoA5TNY/qqNaEtt1U9o3bC3STL
2rSDSuCdZE4tmhBqPu1m8yvrk65KBh2rD947prQUM6qoZCU512kCo5Aojw7rO7Fs
bgjd6NEK+y95oae9V0jbARR3oXq1zpWiLPY524SePk/QyKiDxf+QOrpYgWXS5+cL
3sCLlhhzTc8ezW5ySv+y+/vFFFsmnwwpnXAgDSHJPl+ikBGPB2W6YLs9d6XhOh6D
BAU0cxghiTGoGd0Vd2SHvgDekLr6Lu5J+huVNqB9JT7teBd58Xc/TWcFyl+1ymV7
jecI834jufE+ZSErjidoEP2BtnXSbVIbYF745jTQYIW1rLiXDsFRE04xj5cwkFuT
AC2Jl1XOChr/6395fIohpg0Etw/itGkVg3tS7qDXPJTk5kDa/HbCl6/u6ddqj0FN
f7qB3S/8L7/bUl1ay0w3uVDSrKNoB0V6dkrdwGZsHg0l79Dkhc+lk4lUPtJx34wX
8I/ZB4+KlQVHE6+cOVRdy6KC0KVPQnN6wxdQLODIRLEYL6+uKxVu0CbInxc6r0A6
Ue70OLpkPYPWDe8VB1ZeFUnA5zTniepH/zO8Xyx3cs09MJP6TsiwowS2MKvbv95Z
MR0uwE9Rgq6Iub0ORMdxR0FNWd5p+gl4BN5PUH6Vj7FAPyyAMd/eXKntuRIHZ596
jNyLT38h1YHtB3NOIMU7FsudYCi3BwrTqin4BehWa5U62QkkFTw4ogjDrsUvtwN/
XVoh6SZTMxs3shlIX9KUIl4L7ZgyQmPEsyhYtLlcq5H143riCvFOOf5TszjDzrn8
WMMBXN5f6lPA76aN/w0VbNegTqXf+r+i/9CoxMhe3TMwx8ZtbTRsZ6TL8x9L79bu
xYZ6xM1C88UrrSiyDwJSYrvRaOlI1T7afcBHDr563FKHVfPhxyk1PF6K14wdOzm2
OSXI8t5p9MAWPiXwLc9e2upgfHSJIaSxqXRdbN+rILtSAaG9RpiSU+U7g98GhLML
ossnqkTh7bnzACnsjfdpAEAUfOqOtPt203eiQM32otdupjPComGzRjykkguWT9b9
UVxgos9IJokODbf2m/oQYBGtAn9fnBvGDnewfVLXz4jcfjHaFi+49OlKmtcyLLlI
bKe909EjKL5jYzOxaY9WJww+7l6mQXjU23mhRivE4gHc3ePQl2dvw2iCwk8JnqMf
1D53h7Fcrdg64f6KpQ8GwVuoud7VAWquD9nlVadQSk1qMHAjwlZyLVMBBRIdc+hA
wyrutHiHL0WEX1Jx2yi84IV2ZBkdW4zFM/qG2GtsIGwhjwVvl76E7boK2MSM34Xr
fDZtIqUO97rGjLpbFXMM7Y23CBv53E6AGUvJAvJBbQBcGFkR2qLWuB4Wa1LtCpeJ
Qx3lFZHOpwedl+kp93SPRGHU5yEzZwzSzRHDf+cYhNF6uO24g9pqnTOU8lisD9At
qmkIHn7bIEe8RN//ZcPrxCMc9thb+MjK6HKkRPY5hZ2U1WRFLsgUpepc4K2OgoYq
clQzHagihvkDMXSv4TMDQJ12nwqTLBM2K7HMpO4oEyA6ZLKSXoTGy1pEmHwV6Cpm
nlg/E7ACHwb6bbISeTWR9a4ujULfpALP9MNksF/swBxmLv38RSx/kizS8TsmYfI8
FPIbx/3PCxk+NXigQzJgI48MjSCrZ4CViqUOT20h+F7UdLHs86mL0sEo1eJeQfjJ
`protect END_PROTECTED
