`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zQrxhSCpvGVOrD6yhL43Qg5v88EHWd/UmBfos/qASg3AzFJPmowzOh5ZEDFHhN+c
zZrACPY6Cc1MyNGs5EYQmQZnqaM1MPdu7Y3TZoFl3ku/0a+GmwZUoEcCWV4kg111
1VezNOJ30Z0mZwqr9vPJ+guhSW7K78lmTm73aOizudAWaLImJ9TyAn9sNTl5Sk1o
MUY+Ub4ygOTx8eFAUco/3lvy9KmE08MEQgspOIatnpNnCpb9ZdRA5sBooU/33tGY
Z25PC+UL0pCDvJyLJJprumJiOV9MRfzQHhWdk3pOFQVcNWEkCTEf53cM6IFrKiUx
peoHLTonpEG7EDcvsNEJByFDplPAUFWqf/zVYIBqAUvPzPV1hqJ3w/YW1TApWVkm
IRF0TJgPN8QW51DVIbm4R8pMtcFzgaQDh5RxND25xhjoOx8xfA1tv8NxkE8zRBCp
H5YmUXAX+MDye5pMAhAcl1VLn/LzTSKBrdnTTULdNE+dlnHdvG7LGn4YQ9lx3e5p
EWOSIhobHrUGPpTv1j5J/KrtGZec95fFTsTMGPPGOmahU6zSMkWmORSrV6cC2Lfx
f4yJsPM6coKM1ecNWrAd7YBvTyULlZP0ofMEgdMB0KEpiq5QPN44wyvqU+x2+dEV
RX5P/SH+QZILh/LlD+BznGt0OSNTVsNxOpu4JtFqBSmojDWrqZsIbAg9gfHpm9kj
ymsHyatdEX5fMEAy7PBH7k/U1zBRbuIWMx+BXUJtIXILOFXNLOBar4hEFE3dUE7L
BHMctWGyIR1qtbb8TGLGPw==
`protect END_PROTECTED
