`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A47w6FLFioNRafCKSUKseXdy+uDvrCQZG88PUcv318bti3F5tNVsw5uw45RxnYh+
kdiTTKs/SW6LKbXTGDplFo4w3FavsjPhtJS9aCSKJKDc2pIIvQvy+wqC7kAtIG1W
1ynOO/ejITs6iemALq0qNFrwXbzYcW22swGUH+S9lSEKxbSNPDvoSUyyHkpkSXN4
5PNBu0lQkInqBY3f+sDCISvhijbSKEiUlMpGn21tXuHZ0vWBNMjiYWhY4s0Dzpht
zZyltv/yYfJJ3DoUAsybfUoFkCN66ZJ289986WfIUjnWw9sCrSbnOqHHPwkgxz6l
KC6UWJLzTgVf+zr5b+NTQpr9j9MK7JGE6JE34/0Pis84nDN2+ecZM4K5wqALmQjc
k0+ryihSLbLTRMQ0c0J3lLnaFvfRQKCvqtXGbalvA21Ac3fnKLF6VCLwZeYAY53J
n2h3ogHfSHD87NldSI9a6L9f4AtjjSi9FEPPqAkUChc/mbG5qiolON6iwlk+wf6M
t6AlqBHvYJWOgi4hJGjvtfWgo3lCYy3hKCKUS6V5zIKeWQ5zfFxpLYVMC+eCL/SF
w1vW5oG6X94TnwmFAgrBSgnFa3in9g2kTMbIM25a6BEmlLQbhEmT4upxDtea5THU
gnRT3ZDC8BAtSs93K/6U/ZW86mexKs2XeZvLtAoakZc=
`protect END_PROTECTED
