`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zs0hyLMJoV8xM8p5D2fS4wqTt6EO+en6ZEmAhWM7ky4i6vDz0LriT9dI8xsM/B9t
Y8+AyM8lrlJ785xeCCVQ/DFwCxjQ+A9m4BJ1HTZ8ibuAcyqHnYwJcpG3F6NhFWxv
vIlG3xwH5atsOptQfB5qwUpk2xdS9M2RWvEcwmyEcoe5apsaimwNFIha3DJqSLN1
f3QYEbxc9IGDmwpP5fbynCFuX6xZzzXjD25/QG678PYrTG1TlxGdhWycn9pVjjoQ
g9U5YQn3yPRsg2+LqUrAqmj0Ag8ksy59mQd0sOisXthv9iyrBVxL7P0TPRChpmnn
AGwPwTPVsTe4dYyBw028PRXu8zdp4GX1TRzyWm19SdHkh9lL+e/won0x1EgjuvYo
mF0sDfbYniMsZpdE8G553gBGXOcOHVZg6iH8xsOn1nedk22pMvl7iYD8kczSTb1s
MaHU7C2IHsEE1CJmPnKdb1BSusca9XxXlxATwkU3IseZh27ReOqI/Mlt/y6hRalq
rwkGTheD7NxGDptvfOmw6NoaJT/ulMqpLT1/n0xcwCyukdNgXVk7hPxLvF7nl/U/
tgkdt8D+e+flH9DMUQhwHsVpyhGgbT90yX97kzk2+uLWzEpZX0EOuudHWLOX6AKA
XQBwxBhpdwNAG9VdoU2v1A==
`protect END_PROTECTED
