`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lTFulNvXVPMWFdqCuuLqijeHMXk9SetRdAa5aEdXHFmdTuPFAxzScUr8ZXYyc+En
q9phSZQ47+iy4fF8w3h8XoNs9yZJ8aqseNGOyxCVcO2ibE3yncNlBU+s4c30bLsw
/i8+HKb4nXPbISMm6SACFdLKrNSDjS4UCMs2GiKRZmtwFOQy9EoeGCweS7hk+bko
nU03AqC6gRHih3hjJOerz77FygzT55X05PC5I+Abgi2ES2w6wJMD6w5Gwv1iznIL
IQsV7CXkPU4SIQbZlP0/NK1LekCwcUWlwHzS/2yT7FVrwqHbMQqjKKEIqbZmhstn
PzUfpvzgrj2JLJTKYBqzvILhtYaLpys7PYMoQBCAPpp45EKoOj4jwUSU8XC/2RDy
XX3oZBCAvrH/akIe8g/azL2RgZzM38HWu0ioQxFQkHo=
`protect END_PROTECTED
