`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H+FJRWfaUwvOT6L4nGa/xd7LBa74det7J7VikrDHPkr9F2d+7mVPhGA1XkKstyeX
YpNyjcjA82cvjAmtTj+zXsqy9ZYoF+KhbMKHmyevoc/2QGQ55edvRvKgIw0uFssk
Mw8qSVlhhe+BZmrtbg8VmueTXrr9fVfis+jfaX3Z7R74aKvrJsJvGGVbL9YBZBGH
4XHhKawFWZctR4Nf/My1F2Jl7pid3oE1GWRj+BQMSMeyRFni6Jj9oBJgVMZEM3BK
N5SwPMuJaS6FljQ372UBLJZhKSwa7YUFwFCfPaOaXPUghKUUOAz4CMT+8lmRV3eb
b4P1GEH8R0yzsv+V+YCynuyccj/KPuoX9UR0NNhtZmgK+4+idV+QfgHph0YWOvO8
ybIbTnr4HuRDfQkLiuaxZsIKl5uu4uGXKbPN1wJtZAoGWv6TJ2anuKLFogFHT0WX
RiRVarbdar+I7h7pfIp/rZL9/YDFIexf3njEpyZTVsrg7iplodoaRoRsEPVZwxk9
WqsqkRPRzz3TeDFSg0AdZv52LPps4zfIN/5JKdeNjDO14Hl+1I+z7DbQR541sjk+
eWq/z20e/fWanW8jmrRt1gFQjmpJgajYZTCjorRei/8vs4522EYifSp/06C8ZcB1
dU9GdaDxMwiNdiVTE2zgFxNPqo+0zTiXzYyYtqJybzk=
`protect END_PROTECTED
