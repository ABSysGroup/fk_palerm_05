`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IRHndld+T2z7o8OzxqWKD2aryj/pPkL/4VAzf5tNtsHuDufjXbZCxww7Ol6cEY+8
4Oe6YYNQpD2PFW08pFjKuMA9XDc4a4p2omJXQ5+cRlSoBIpMpZNnDKri1Iz6SDpL
aZdcM9667o25NRhPuw0UsHSx+fZ/3eJdVkxZltPnt2bcjJSURFWZTkf5pfWq3TJ6
hsXstV61LhLSK2pz6G1kUOUXiem+WdrlZQTKXXOFM2CbtXFVcIJklw3Iy97qaxW+
lP8cI6TunikvWkTePV5U6vnE2FHNeDgUxY/ItyroNOIY483pisVSVXuLUYCIzOR8
Z3bfmeZ3WUsM6twrJ6jh2Weaz8cXQ5p6kXBh0uYinzkKWgs05HNTd1AoGIqtl3vk
E0NSrWkoDkLPTQBkMEwwP197ROp6yUxfYsRxFAjievw=
`protect END_PROTECTED
