`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NfuI7C8qaojBebyke/lgYI7wPfxMU7+tPNdFDVAvEUvyG3pcpHxgtJ40NrHxwNBy
6HGFBCmY/RK5HI8Mzjh3VS0ETsASCdzSkdxBFcoMsMX0xdlaeqRBSNGMOr3Jp0rl
ws5o6IDYzhKLQgCicnU4JKv+6B7JU6WnFZ8o57olP8KU56kbbTqTpFlAiT3WvtZ5
CD1P5mWWT5idwOhv0ROTnB29XxYEXaATAql4yKkoqzNHNjQW8T9ZY2tY9BRoFldG
7K2J0/buIDsb8ExzbPwGvo4CBFYfg1M4720u0ixvvS0pQQuRZT4bARazBSKpEZb4
pBJbNqZ/34A7oupTbfuchy09Pj9yJ384LaCqsT3mDqtGAFeKbo5SLPhYop0PHekh
7T51L3hUCvGwaBZQ9VyQBrF0tfnLyJV9tJ828q6DnU8j+x/HxJTb2LX+RvcycN6s
QxriRTMZsYKh6HN57igm/qQKFdn1vOSHvx6uQaB+jjlxX6+FSIUNVl1Fyhs6WhXZ
D9kk9p4mvAALtNKUqERWQZ1tZObXPnZ+AL5Rgiql/hv4ofPLv2Q4lSUotCwHcM8Q
RpAwLDUxpAihul0v8gNoZIEXaw+KfGovSBUl0OJWXENwd4uAstZUYVPljxXXv1wq
aHJbDskBl90UfAJrJwBhbw==
`protect END_PROTECTED
