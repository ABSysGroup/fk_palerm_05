`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z3pTiKrUpRaHhddrzxYgoEGDvL7svCcE1hBJR68fE0xu3gKoeCScH2WyzOQv1U8e
9YpW2NcAGQUUFwKKfgDUm+AmEmr8NJ18rZmsC/00PPx0PkCKWBH6gKD2xAegVecv
qjhFVc4bMm3OpOPaKku6p7dKyNkD3/0QqDvye3+f2Kfu3tLrXSK2XJigoQar44r9
8of57JnaA/Znei8lapHaCqXnpBdyGezfJJ3bMhZXJ0sj4PhdrWJHwJYqWdo70c+W
Q8/PL0cYxX0iamaKTHDYc9OUGHXjUqPoORAuRlOCivfjExwlAT78PJ3rz+3XRBm3
pUiM03c3y6JZ++cojKdLrw==
`protect END_PROTECTED
