`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
drNwQb9XyfxxgvLre4W+48byyPOTXv7E2KAUBTkK8dU4eJ8z1EpmdaBhUC0PGKo/
068oX6qFjoL/XklclFqArIHleSoksYgf+KbZvxJj1QYllXCYGUq2SEWiV4QV+8Ro
EtZe0DTEbysRYksH5/jmf+eKWCycMPs2hEboJgj0BRkiiVST4oTbO843/H1RMaa0
Fkl5KADhw7sCGYQ4UMs5waA4NPrYZ9g/xwLNJPb+Wy5t0w0TmCoHUi6XawdktdFX
LoLCrOiFAzMTrTJGoSvxjYkw5k1XmE/dHDonDu3OyT0tBz5H5Q/4bI73PmwCnVhw
LrYIMVGEZ0B0R+i8kMEM3/ijvu4JRplUjUYoqvZTAZozw7KikHHRfaO50x3ALUKm
PD3BSv/szxEJ0kWQpzlWEeqfyLudaAicVIxXtCzxQDqTDV1zd/XRxwiZUXoFx7CR
hKMg1dVzSKxeimvGP7oCvMKkkA5TlSQ93i7WOQxRRqS+GBdKgqR6Ipq/37rU7cBG
TnuwVTTHzXQGCpaoYBIMs+V7Eqf9OrQm2yrImVU5wixKknngwoexSEtQxtZVBsj5
v5XD9YnCwBFMj9QEV0K2YPin3uovWAseYgwsnAtKYOZX8t4aPqEYzTwHIsXzE91K
ydbt1ja61Otauk6fjwt6gB6vioPng21eCN4wskf3nLJD6ghQufzmptAzopPhpWYw
56m0hjpwu6xClVOY1RrYH56uwnC7Rk/+GNDjVmwNaBtsuH0pjpvz58x03Dt16ww7
xQtUDGhei9jzf4oAHlDlJFTxoRKGTHlrJxNzIZIqmbrT6KOG7GrEHXmv8UaVNGjE
Va0fALR9rGmZzH3Nmpjj7lsyAd6okW35L4ophId2V1t46UnIunf2yrOb8rh5gVDn
qev0p2G4IjkyJxx84TSK9wrfp4rnLCtInWQ+vLjdbunxfb3vy2NKiA6EO0Yklg7R
/zsAg8tc71PRm1uOx5j01D2ABSNK19NIWaoeS7uh03taCJHzP/DwOQPabWNkeWj2
Mf/7vX2SDiVVAzWMIuHMMhzF/IJrVqwzMZih2qxHZlaa+gNf/kieBwb50dnjePqM
UDkEt0mDe2BWNwdMhENDGgXpSMkIyLZ23mK6RXp8x2hszWFriBQCeyUm1/0NW/A5
0Fu06kyn2yRKO9VJ8wV4IvkInqnBG3xDp5WcPFfPDKBT8RBPLjjg5u3hu3wvZbg9
+M5lPw2G5AW3RUiQ7jiByA==
`protect END_PROTECTED
