`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
24lTbw+Mm9dF+19sp4kM9s1itxD8EzRWDUHoHDuQlHkBkIIYJezNspQ9n1tPbT+F
s5D+bErfAsdPz+jHpJ9xBuieMfbruvLJSPptvRdfROYHFUJEg4nR7VOSffSU1+Ab
qVQtwr1F4y3rw7C4Uj0mP43g2J+hEhsgN4oOX1uSNBnpL+rMMR1s0AXcvKWsNXWE
rmDIS3qvRRqrCfmOQzZeTLHyvXF9pSRFsMz8BXk/owLBxo6FkLgWJd+H9sYMDxI4
zEK/72Tdk3sASOiJ9v9jnk/2ZkSn1m9Vo608x65ZSfu5zY9K81SeSaNAQEJaioct
gNqLdL8XOaVGlSJaIo18eVSzN+EY7skk5pTjPifLN0j8NSs2cTFuK3VcqamBy0jR
XUn8AWMe/Ea2gjDoWnMTP40ow79rRkYAUexj1za5KAJfeQAS+QOBo9Kn6uY3+8BV
hFHe/HimkXiSSFU88NXVdw==
`protect END_PROTECTED
