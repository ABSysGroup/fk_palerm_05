`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mikM9mMrB8Zsmuv3LvysYymxwRYRqKOMK5PJPsiKnAxHQDpvtstpw4qAr10ZRrR1
b3HBs+5Y2Akwlr/v/hmrHkQwZIGcCvPdSnirMequZ0GjoFX0ybtWV4pKGTaiBRcS
JWT49hZm3vBi3i3Y7uITMFBzh1xC6fqSj2KILaGiRbGEjzdGVDKXDXSpq4q1Sc3b
x3XMe2dh9EzvUcESsv9AvgInJK+Erv4w43lv2s1r9GcsH6BKb7veqQpYsNH+cv08
Sqk8sJf07m0aW8H/Bjkh3vXL0/Mp0UZAYsVXl25xx+6hVU19m3HBkXEH6m3ONF/6
DmTkijtv9PH9M+GLkirvLO5XxC8XUEL8vne3TIEhpC6WASQBwZ1pOKK3RjkUhUu7
loD0pYV4j4lMM/i9zsj4EuwCd1xpvE/gfxzXLVVNX2wzHPyIgZ6YBzITWVrHWFYk
v7eaIEjFrBM6dyKCyxSGWl+eJt7ksjIivvno0hDLF1g=
`protect END_PROTECTED
