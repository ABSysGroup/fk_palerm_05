`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tAr+1TIbYkPNDn32Vf9Chladf11eksEyap2DQKXpnhqgdY50rCLQjUXSxaTNDYRP
DDmbSYeJ6hszYh7p9DM0mLaaUayfgJbF9L+kaDgMEqV+KYof8z75+KpKfrzWvTrU
PCkD8OcZHjdmIm/qMrt9w+XigmbzfRd5pw6rJvkCvAd8Bxy5yYpqLHu2GPdT0kLH
nEW4zYRUuNdS9xcYOjJd5/FrL1bYHkpog7BJBaw/gd6Q2MeJT1eoc5GkaKJW7LPX
FLAEoka3Tyjv91E8MueTDoulrc8TMa4xkMdj8LYjYqi7egkxNomyJjFtOkUrCci8
CR2ZUfwm78wYF5pjm/f3ZDZrdhqKi4EJjfyiB2Iz+yQ=
`protect END_PROTECTED
