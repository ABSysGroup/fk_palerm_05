`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ym6+mU+DLToD799qEBXO9tR0GJeATaEYIa407sXcFFT3giHufZbSxM3VYfPFeH3/
HgUs1idh7TI7ok75RnKRvJB2dLbzt4kZLmbEH4T//xQv3utjKiXEjRVqy9Bzp0QJ
S89VPuhnqfTJAwB3CIKTIaFjCrq23iHzy3EUO2Okn49ZitKOd04WI/D3otd//Dy5
t+HUxYQIuL+nhfI0QIt4F/1GXb5XBPhSRkIqrJCM5JAH+Qo+htuogmRitlOBA4Rj
8315BRSV4/6GbxUoUe3Yc2YdLuPHbukeDkyx7QlFGf1AuqYtk6xJqxFrDqehftPv
/hpsIs+HX9Qo03BLpLuIJYl37OsOO1+V76maVk2CSUO+kdnGhl2zQxyR2ABn/E8P
xWL+RCUtjoo05sxMMo6zCKODP5CoKYuPPV6LL7laV4zFjWAU6VxwkWFTNDZRkOe9
UWOmRtUixJFqnAVYna9hzfBNM+27ef8P+QsTVVRWZljdDRSPSd6n/Eabrf6d+P4u
IgZUEMoVhOWL6YZi+FWuj6Pq13EaZ4x3od91QbZZcgo6+UMvKXTdD8zxDe1qER/g
`protect END_PROTECTED
