`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rHa+x5S+0Cj0UlsafDrmMCuGdBus8vWfKi1EJttTV3tDU9uEMh5J6PISdY2OAnuk
QnlDSKScLpaDwueWQ7b2aGP4KI0HZQiF+pCedTdNJfb53yph6SCSq05fdaJYbHPx
zDAw4UylS8ELwmQUc//6CFwRni0q006iEaKqYVVHknvsJarU1Rj1jx1SaSs5ICcl
CFQSL+XlXDOhU6nqKEEkLI6k7BirBEb+SvNsaG4iReoeEoHvFcVi9llDB1yfqfyR
rcKHVqN00eYzcuavrBBeZ/tWcAj6dpXtIRS1apkgeGltLqJGH/RAZzFs3x3D3Sm3
3Slf3ce0EzJJDc7v9kHhLo3AZQuBHYG51i8BXgjsX6nsyD0TxxPR5YKG9h8jdpRs
1t28YWGvNaGSQyldvmPsRjXExIDTXNFjDvWmWTL+zKRo+6nZiOOdrSd7nzdZENQB
Ab0Zk0+rbE8QVuPlinTgj/MKmT/h5o0010f0LIHZFBjru1RAbWLfUhwF0B29mUf/
9VFl+9xj5rhwK2QashhwlnVI8lHt0TXN5sz5iBNj3qjj3b8YGwnzUy4VPDC9TebG
vyawqRY4wiRHHVR/cWVHf2THbBZaba8wtgnpodD7RsVLZ69TBn2d1YTG8t0tym2G
U7HJjvcHPt7cxqy19A6uvGuXK3Z/pXe/IvTUOBWmpcg=
`protect END_PROTECTED
