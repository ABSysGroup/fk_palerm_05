`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/6C6vTsjXWvLFlcXhdu0HkzfUpGubctV/5PwcSo9F339rf3mVkOTYtn0IiM++ZFU
KaTjYENfE14mMxzcGy/QHBGTqUCJqKE4c04+evG6DDO0XUxZOsSISdFQ0QHzdGGf
/03kq4STkoeRgpQfJbDAocbxmeOMjaXELIxcPsm+zz/FaQBqWRYGZmcESfsgZNi8
bu1AYq7coz449Mv3t2mTnSxk3xsG2jU4bi67tbuOSajIrR4W++F+kLE30JQhbupx
AklvUSNXm0a9tSWRM+5umyELwyBQlZjIssNVsnx+zq5BejEE9qdoCO6o+Nlw10Nt
tJsHHkk9lzVmJHqFcwbL9Q==
`protect END_PROTECTED
