`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N3qRjU7fMReCrJKWfyzz0nWsctJHfaRqU+HNFFfspNaZuttWiqlpufMTxKL6SKRw
XYqdcbCtoVuCy5oT2Lk0Y+aaX2rKDAjTUMUZd4pV/85q05UJiF+SlRI2sny1fUyL
X66pSHExudhhDaT/L7VFWYpHFlVPrtWmwb45k/8921Ip6yQ9rPwQx+NtZ/bwfqUN
1IsOTzLQcOqXgXCASEWA3/OQJj92PUpirJNabQ8wKI8Rgp4JmnxiHdPz34HLUHdZ
xFjRhtMqh55e2oyvceFvbrJ9SSQWDY1oe3OhgvgOWChSs49U8r5bAuxc98hzS4EE
tr8OBxTO+rjAkwnnORYDBQ==
`protect END_PROTECTED
