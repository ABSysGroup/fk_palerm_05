`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d0H/BTlMQXvnYr4qF+Xer6/0sytfr6WyUtMviQsxASa4feeJA/QnARLupt8Nlo/7
FK6IsFtrwQgcBhmhFHxA8IvjDurAjWC00kJQ6ht7B5iCUt9RvrOk+xPyY7TWTZNJ
D5lqxZRxNyyu5+We6DRrY+cCGqm7hMB04WWUfQgThehkcMhrNjIKp7mLk1LcIp1u
Mlo8/6BSmxM8jv2SgP4eX7lhOIpyJFSsBeLHLsp4wbmTGo/AyNItJhq5zZoNnrh2
JQjc7F/ZI4qWoGt8I3xXL4R82p8vZnGnKt6jYCqkO2+RPRfpQj5K+raB9WP1RdUn
CNyXuDLnyeVR5MXxHJdaRU69PSg/XUt4Jw90YRu++Vq32hgGYghXYwYhuYd9ee8q
A5EOJWpVwUjPy+E9fBDQ8SSUEFc1hAAXLDPHyPRLsBuLzoenNBl93FSDLjuV6w4A
op12W5vErUra8tPKhM5aFhod7ielcfKNA9R6cx0UxcTwqVp9dnIbmo9E/b9jCW7q
q9fk/gU5efFHHOtb3IDNJKSdP1aS76FhvruvlBdNU0QkL+ovWelfvkA8ZiBIRi/v
5XSLX8oc11/0iDc4ixH4RHOOpvgvgf+VJLb3ZivSHGI3T5PNTtxholNjeHOmjw3Z
t7C2496etJwXWaKf4k+VIgJQCqlQ1plbaWXzBv/fzszhSTUp+2U/RlysKuKvtRpZ
AebOHkTzttqmNvWaiPxrAFkCjzAu6n7ui6nZ8h0T5V9Y987drLiCwhBXQu8ut/Qb
0n03UANilClatBHnfnfdENFAUSntn+PJiVxRZe5jeX+Tjkj8xrXhr17PFR9yqx9/
0ZAFEPf00p6PLZlRpberlEDSHh+JOosEACLw5SS0hSmMUMh3oVd9x0OkxbngPm6Q
fRAbgIu97+9qWRSXTAMRaoTqyjxMrUSYzGfaivgPt9+U39ZZLJEGdgDghCohG2Pk
vhQTfXTv3j1WB6ixmuUQvVlMWy11RNhagBumCC32+9848XNDDX/HwyCo6T2oywJT
3DUn7qMbcTtS/mHN/nqSAq7L7bRGjTa21fVHTjNCAydxHXqcgWU1VMPov6T9wlWW
8V+KAkbBvoPsJQNfdSu7k613shSYmYbtVScxYIrA5IpCTM1zXfNKcOju/Vi/CLu3
+2Z/gsQAtVx/qQ/xmNo3bsR2ei6ZkmbZvfDzvHxX8v8ZQ9GQ89O9JLaIlZtDbCkn
Ygs8fjtdHRtWt4duN9wuTuu/WCPiIKj25IScubsYy0Vnr45745sJH31VClZJQ5yI
NAItfVPO9kq5zh8XGMfSSG+PfXhUYQ9Ew1LyWx5S8db7NrLu7OVvOSj1QdAlGkcC
8w+BDx8eVzIvdbORs+NbcaarngfQwSER4LcvEcPyfyESTSvxcC/KrwOtxFMdFMOU
nodAmG8sKwM27TFuvq/6KW5HrwTMaTVTCMmDuo9usJtxaVrQY9Jn8cniBUd6TECI
o8h6B2gNv9B9Cr97Hvz2nJ12rqXJaP8UHGcx6lcR3r3lLRkaB1jxAcx5tyYvBhSU
OxQO7bYYaIca72DtbGV/QjwxTkx4D08+5ItvRXrHlCQKlQnmleWFSUK5OVhpE7Eu
Rho3w7oKyURfN9aDu9OrI/AAsI958QFI6wZUwnHBq4M3AD82bU55JleWUu+esZvD
GZJqxM+tXQuLuhY8HqLcoYjajB80/sIdfEflcxiQq6wafySNyYcVw/1L1DeLMUzP
VxY87GVvFonFw02aWbKN1D7/jBG192v0VsQG+ZxdTT8lJ+J+j37CbdOPGvC37wlv
LHmTpA0aZs1b/RzuKMpgsLzDN4yjtaYagUFjCreBCpX3CPvV5sEiZLTT6T8oLkUg
GUAHsONKYyIy7CuI8eU34HT6W/URozrjBINNSgcPBMxJiZPpNuUmoMJAsaUEPKr6
96sx8qov0Ll5R+5HCJ15kM//zXwqDCgWD+kPv6ui7UQgQmrsuwGmEdz+EVkT1XWI
UkGN1LC+rY0TkDy/9Dp1sNitMh/xf2zmRiWKBrEgw9bDBuHKax6eW+OXxpcG6/UD
lZz4jzyRFUyi68FJddxEdVEwNaF1tJJVUY9BWgK27CWc6BbJOWnGRM5SFv7GrkbN
WwOWhidSMSFDM8/qMhCeitiP3XIsnm8cdPjekN8daGMqd2Fgmp/ZGuPNwY/usaZj
6uKuKCXEZXuMmRBS6d0WqCDdUQhU1IEqWpSMcXxyiCpRZCY63lujtcgyST36q0/F
+OIFTLSIIifh6j+6PyCW0+TxB+0Uw85MgHPELV6C7xdT7Jh/ffoe9QzgLQ1Dk9jp
lYGhNGZvL+8junWJR6wWJ45JOgCGIrDF7bPRSHrWOrfZx825xP5beodYKONw5wnf
BtdVR6zOjyH5R8abNrZeCTYmNwbrPQHglBnZNyGzslzhkpAVN7gGL76prk6nl1lr
gJEPZOt1VB2MbXQ+SR5cZOZr+MWiIfoDB7sHh8YUi9JhX9HczIv3LgZI7En0OWCB
rqoa5/IO4S0k1bqkvVYF79oye+j1nvtlptny7ZB0y8zZbhFMeoo2Q16cjxXXwIEY
1CuEgG91KslRQgSJMC3mKKeLYYYmYEiowH/l1BpszwsV+qCVRszmA4tseUtimAr5
nIHcMYVp/zNmoRjSIdXWmdR6nDQGb+0F5OTRoEd19emQgaPhv1wvdQg7Ep7Q2ycR
CcZtAUKZc8ZDHhFF1yeDxp38ZUfgCA90/p9cpJbU3HI/KAYlkK5yKvNLVGg0T3rL
pGUuICFvEYQuqn5IacT/Fzmnu41WTjKgBkJFUAanedk=
`protect END_PROTECTED
