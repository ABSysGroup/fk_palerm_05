`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yHARAiPq+/Jm/6Bdoj6Gj/YvZtSKCANNTRCLJsiCygNJv0wf2kBfEFq35VLl+8md
8jeiaCfMvl2fu3VC5doQbPE88bi9HNODtHb6IpWIuMoFEb3aH9J4UvApHYjnOesS
SGE0ylU7nXTdykLsnwAN+KnH89J+dQR5gjG9yu6hEhhbkP54SdrGSnSjQ6f4X5b3
30JLyBGtD7/+yp9viOIhjMpG9zftxWrzqH+WR4irXHEXMr5Sd56OawAPnlzXjfcB
B02NCqPTe7C6EeXnwQBmBY9Ax1m/ZIMCQc2zPGwAPRvRk3644cJMG40+MDxHmGTI
rU0nzc3D4ZV2f4vfhKumrZrBSFRAfBFUUUW85fD4sYf+1qRNUjDMf2okiAdjI3P+
QFf7X8D0RMRU1dRTTX4uKeXtL0cVB7uMTf4daMr0Fz/A2g4AMDOA+ka2Zx050Q8l
xIgxzS+iXhO0Ue1ls/BTUocJwIIz8MmuCUpscsl/WAC+QeFWOCHmEtzjd9DpHRnx
2fzoHeizOoEJf8RlZOW7z1Qw6oPZhgC7NbRXh3zjuoR927svkASgYCa8sGDCme2I
Q64u5/yxQVaB3izqHWrEDFAB0E2HdBMW+BJ0QJ0AI96m+OhEK8LDrAYH+RjOybCP
8SeL+K1lbGHgyi5pFkcDp74z8Q+sxXaPbJx0YoH3fLzLUP84MErfYdpu7pEiE9Cx
mOCrAFHVdjOT9PgE9HDLtPgSNNpx+91xyP79igZLy+R3tHW/mRaLVbTgXXWMwcDU
ccVazpWbe0UVVeYZmeMJorgaH2tRMhuq+2TRJgZ5DDs+J/HRczUrhLjyro0GTup9
LUeZgUNaVNu3sTrbNevGBaLMaMi4lNr2K2OuQl+U63GqF/CFphkzU2B+t5MG+ptk
5wXAXyUVigZv7dWigNbW/4ZT+atFFs4uIc7BDvYiCjULlbDCZE+DCEdbKhMB5z8m
U+nQ+EQvUPgQ0mLjTYfjvE6JC3Kij5SKsEfTAaChG49G/6jYy52nkX3paKyDH+kj
+m020XJvFqHkiG4FzG9YK+Poza1Xxl2cm74P5vqYknFYylQmxNQ8r9a6Wk29fUyb
Wv8nZJB0uFpvV9BykPKg55iCqnERE1dD6NGuL9KwbSInX+UcTHEPu3Jkq19eOr0l
XBORBBVFKdTOx2WtimnVLOokkBxE0vHt79FTGHcw7qqOw1Rqr3f2OfhzR12T1KC2
MWVGWUCQIhHZymmqwwhTZcjIWMIT8IylpmQ6a1+/cakVlzndM7CgFst1Cf5GsnPa
jn9F/nM7/SIa6dg6oeVK8U2RQVAzEIiCx8J0JbegtV7ihG92a3Uw6HzMN2aT8Ibt
lhleMi8Ye8fY8Bagqn1JWdI/WjFdEOzz1AUSnA10HZtPFM8iKaWVdfBn38fOtzeV
6HVLiooVSy8Ikles1yctWyE/Aqu5x6U3zBJLmCXdlf8189ajNOBtB0OKza4r9xjR
vUQz8rGBiEGroU7zCHEy9tPWo/8xl5DZFelmsukdTokY+gTGSuJl5fK+rNIVEmUF
PcCxyMpnML6xICToJCOoF1rWwGZobqYANkfSAozzot6Mii16f/oZXOEqpKTshhgg
TGUVT2aMR0/qCPgSUaulmv0STgYKRGN6Ltgtxtp2EF5M3251+9CFDpbE5XJZQ1CD
ffrOPM4X2+3P6o2nl5HseTtOBcNRFWObv/WhZn2Xfnk1YA1Vgo7y5Gl48gkonHcg
OKI7Gxh7FNS9JYhZsLrN830I1jH1oXEOD97FrmaMfnQYYL3uhDjQpOm5e9FSeFfS
2UoR7jro16qdQUnxlyEavZLWNypoPe3/iMEy7czt4zcct7hViEfXFNs6pkici6AG
Ue0B/qtlydH2HVUeoY+rvHS61ZUPEwsjoOAmvaKvA9cCdYFhuRwk7/J6la683f8T
S9QbFbqZVKYzX3gW8CQi8KPTysLPHAH5fOx8b2eTusq8wQC7gW4IsPNAShQo7eKs
F8cQswTUTr4Tw84nC7zP6zU1Lh8bxnjpYWwUIl2IC2HbtXrdWpQAqo1XE1izPuoH
J0k4LgjVP/LxyrTXXtIxLLkOuDMf14dWXbZJqwdIf28qBporT2UmqSC8zk9aheLV
FeneRIvfrCpGeHSurm3RLtOlYE8gQa4/tXRFkaiGxKys8dQ+UAMUlrKTV/3mE+nn
9HjoZpCRKnZuzYx3drFFsMMGECmxR4oyAhhY4TqD38b0y2fCb2U8SuTmu/0Vj6uF
9XP5sTazlCSgwp6qQBjnckoZyWaQB6ItLKoBDr8ljtoIl11sjKjC8u80BzEjKX4S
hs9Z8lSfYnDSTgKq1ItezsZo8FpG36aBOYncNBoQO0FC+XtfBedKpyTjuIFfaW3c
nojQqHhDALxLsHrF7iNJgHVWxaGB+nDQBDrs4QjkUmbEPos5pXqvC3z7XEuNLibo
Vzg4A3Wc9iOU0+vf1mye1o0J/Vtj82pBepSrtG2c02rO/NK9j9CwTJ+O+Wt5fCJR
T8Vh7HZzbFLnU9zF1865Sr+OgOKwNscPBkqaUtHqXFagLjJh0b420H6IdEWVJ19X
5zqco4iG+VgV2aVJyoDU/HDTpWaIvJw+Pj5a9qGxC0P7DWmTGPspdMDb4pg2tjR2
tEq4NGCQ62vO2O80CtjkuXvKuAddA9smfFWmLW1KY0k5Jlz7usVnpDWoqDlka3u1
3vXdy4Uhw4fgGMOcvhvnijYEBiOA7FnJ8oAnorLhjHI7wZHaO3N146Ww1q/tDdIl
y+LxOzZTN5s9qCTGSodht0Ldpo4B0TnV1yzIypdTCXgek8vRs10Qwr306yYBBtTK
QHMXDyiNqpE8xyt0mB1aXEC+aVkYZCuM6BX8oompWkXwPk24QcDVHKPADSmvaJUN
+/ghAf/P9VVPNeujpqWlEgezcmGlOw8iIrlofg3LAh33fvw6sXwlSuR7sGtgp+Jl
B8swLjGb5yIaWX24OWF7lVZuC5WlWt4O5DdvCF03E59eoR1ATJQAHoLPHi5j1R2+
x94gNnOkTBP6WgT2x32Myav1taacfbRugkNUIhyCy6PgkjsHS82OE/18btgqrRRC
IcEMP9kCb4slCxQQSqmLyMcX9S71SuDrG3dg5zxnhArfJVey8xYs7ZDfqK39J6zQ
2tt1D/+ASVpjoVViZyiHUzjKzbETAfrO7FjiCGlsNMwU8AwGM5hTe861JrHk2eh/
b6eF1OjU4M7L6DR30VO9kExCgrBhrir34PepLr1TlMorqniQeL0WIj5NkL8RwF0d
fZd7xVky4bGB5Tc6KkiDXq3OpnIYUCuXVkWJ86PXzi1SC//m+6b5KwFJufDi/cr5
yoAscE3EpdqdlsbyGxU0p1kFsaLq84MA5w5ofpPtHxJxBrOpOMhFcfq0Vp5erKH2
L0dRR669MCONB9jqG9li02qxyPXhAggVqS4W8okKiiMDMAmUnhKMuiMCn+nFywrq
WlHQ78XPx5G4g62x8KQLbNPg5wQRSbGws3TdGT/NFv7nKpqksAIFskKt/XSiqwAB
CsZ8AMv0nz7StD573jskKELtblOtL/1DUAG46rf7/Ck=
`protect END_PROTECTED
