`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kxu8ubtm20aavJTVP1RkTWs1l/EaMSjbOXLq63koRV0GKA1R78Q+jNPhrIPEFfVB
5yCvs1RDUpaT4nYQIV1UajOEgESDZBcvBjQjF0yCZls2UXr1xxumeI9i3b4m38fd
bygDcuW3Ol87JMnfEUq4Uq5rgYnN6rP8tfwzp8m2de0GDf9ZQLr2Z8o9dgldNEwH
5vrppR++awZt6a9GrXozbyUkKdRZJO7tt00O9kKB9PwuOrss4CZ5D5zyNSMUcPTg
zxOKq4BXc9XCB9bXDkIuUCEX2F9+8ZSCXUg97MQu76Lc0K0ENy95W1SNO5V8ilpF
WShjn2HGUKKwmZ+e9KdWdzR7mu5UePmFZtg2NY9O2p48lo0V1ugLIu1AKEuX+DxU
L4W6yAu+5vP5+LJkTMk+mqzu1gwoc+EtB1W+PHQqSgkWrfkU8ugcE6ito+QJJz9I
wjKw8okgLY6RcAScorcIXNiECoD5jn1NrwrRsrUFO8sYzeEGEfPZII6tAHelqbPx
NeGBkbILGLTv9F4jovvlHg==
`protect END_PROTECTED
