`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XyW/D4MQbAQZciO6PymlBeTpNqNjhQKdPDYUv9ESy/Ck4Iha5+nfKVcok6kNTU86
0KI/m1U9d1kOHQQ6Mxw+I63X11t41wK4vYGmC7u7ZKigLVQK725mWxRNqsXKDzqc
/VG1Eh6fiSIkrNy366neFhRUDQ2xjWFzCh3r3bNARxLCezdJFEBBaqallX3uGgTY
GMcGpsksE4OSQCCt2oedff1hODq82B48S8RXdDktdQJz0tN+Og9BFEjGYrjilJAq
XffET+45xaiPGbF643xyqw==
`protect END_PROTECTED
