`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jtQ7n9tW7pBicmLfrG/Y60x0yCUDtGAVqM5WQitKlM5bwiV68aN5inSz+0dLZOxp
y0mhPn1IcjZ1h5JfRF/VT300dafxciyP+0LjvRUzFVHcCJp5T0A0PS+W6nIZUCMO
wwC8I4VaOmZbLG/0c8tp/ihWzfTIGNTu+juJtl78vrd9DmmtImwzwei5opl0i433
7OkQ4w1+1+nDuvVZIiKKJy1erGHLXwdmqWz6qh0IO39hKlDiIT2ON7ZorzlwPuqy
qcV2X1UDDp+1x++U3fmPtWD9Y1eWe8YnPco1x7Fif3+5wsqtRLYBgdUHgf4BUgbU
Z+Tu5TA30NeDXNV/5R94N+9IIgFvbQ7fOdAWNzIqF9298dVUffLlyv2ZEHo8ynOq
0gGIO3LMZa/ANp9qV8gw9uGNdYHNqZlxBs8pBgpeQq8n+F+KEDlvqs5g/QDqWA0j
lyv+oXV4tKVfpRYB7krH0VB8M8fB+ctehUS699DZ16pW7tNvcvkyKwyGdIdz1CaH
Z5EU3Lwizm89SHsVyU+/+BF7+FtgMiUvHjkIdWTd1uKj2hajCUMejsUCJE57cLuP
rMwPh7KE07+MONePxscJul2W/3b2zLmqPf3znJzTwh43iO0Y9i7mx0HHTm53kbz/
slYMGf8qGNsL3vnDInk+mQ==
`protect END_PROTECTED
