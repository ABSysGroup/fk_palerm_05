`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lTqB+YxxhTelaMxQS5TJn9mt485/DS2xnlYTeAk73IYXIUt4qe2xYBea0AQ7TMUS
zAiMTcz0oUhXCFUbXnCe4CrDj4jFtiu+z5oa5gsk7w9xECUncylzhdgLelXKf6gx
G6uxZ8cFSwXJniiXS4xhyV6Znvfry3lr3FcPbZPDBG5XEYjsJlrBZfHFklKfqtqe
4wxSIwOhe1G3rwR4eYWoEyACt7Irn5/+WjPhdJsAa6/B4kIGnDZTMAJ1Q9CS1rsv
z6DYn2GqBNhwvW2M0NEml2+lnmQY8VlvyQdgEe/nC2q4z0TSfrH24vtpYNSy+20z
hJqrUGHj3A7KNmhMUrTX6Y0knbqqiTGA+O9zx0I9fmZU2G7bHd5ZYvxxFOVuidbb
08I5J1jShR1x3r/fGAfO51XSvz73n43AhVaJN26RzRPuwNgwaouWuX9WfELGCHmo
oL00tmgFiA9VolEzMGvnHmq2PK/iYxMkZGZub2MnlzQ/jP7cj+AoasyYWNFiLsV7
HLQrstW0BNBeRLMAK6n4Gc2l0NmUDySszWuTX3PzzEwnk6ds1T5Ka2OeLY8IHQmj
EDSA/T1MCIVGr08iiHMzKuyiAjbqaFYHFibVzKLXd9/IjJEkegA/3BdCKAkH6KuR
QPe5dG5QL6K7Wu494dcUu5Wo3sjjurUWtofnqfBtDYncTxcNc2ePDVkq6p5eTfpr
JUQpjSLRiGfLOmfBUV91BlcKT2GmHSt9ysCKob2on9TCnoBoxZ5r7inoxmCpF98H
xdgq7rj+kN1ZyVOD7jXoch2o9VvBIzdJE24gYq5eBQ7BEsZPrTtYO35ipu1e5Fxe
jPj5doJp6yhLKzHUnnIs+sNaqPWujb650oLroeyT9lBLXJ1QmjSD9YOtjmE7W53a
J90moMBpKbAG3qEcwR/zYwosKLGfRKP+YQLZXaOkomKhWwbFYAmWo52y9jb0dm6A
w8NeM4V4tixUezmWfy6iGrIdwa4eexvB+W1Hg/w/bvurwtzEmGET12kshNyS8CKA
wrVgcvyl2JBMLFchRLQIjKvQkPXbARpXSNOK3WIq+pGS2cWwgKL7qNaenjcmX71p
Cj2u9+G6hqi3Gc8Yh3KfMntXqJ1iVedVoG6oJEUDG34U/Jy/qQyEcmVFUC4lJzBe
Yj3pkXXq3LNVBz5LbZJvgZuiwIHIhKVcgwMMcrMzvXabAy2IxbUdUw/EwQfl9JL6
S+dR7y3e7RQpBTA4CRh4CQY7Bv72mSla317mTOplMdyU3LwztiXUfvpo7eyKClo1
Pn76vCyqV8Ie6VQzMdxRn6Q2+xokB9u91ts61Jd1CqLJyoQfnlXONWPm5g0MTS1Q
273dDfkRn2gBzygvhQARlnTgugfNfat36WyRYWyCzBWya6zVg+QfcD2oHlaW0Vox
j5S2GEQ0UBLWGYw9aVwRREWMsLJDF0bGGlYJSx0K2vCzoMDpVVctyRvECA+PqbyX
S9YUY6/E8A421gpsDvX0mQfHdI8CC4K6X8bshUq4TGknLLCBL0I9aGDpbxTZC/kS
RoqtVoCfEHh7gTYR8h5H/3GpWtpYdy6bbdzDdB97CDzzpky1E8ByHQ9QnS8KwhZt
69AYKTqU9p4TPL17iOXJzz9DI6A+8UWMtIjGZuJO3OF+L5ff16Auv5kQ7FxXPcx3
zR/a5NLof8n/cwQSmRNLb0X6Dmj/NB2Qjky97EGiONQYPEYrlKNCKVL2TE386oF6
VX/OUG2b/q9mQw5COuDAOXeZl5rSBstjdQP9qDfocxdUeoviQ9fw5AMkVKqe5JtR
84r5JTD7n1hk44ViSeKGouDEkwmqTjNkav3LoCRwGW2mM0Tt+ERdcnUYNKSeQ4rZ
q/DdmBV51PLO6ncKlZbesjAL/iKlfW5jfD8IARahOCBRCfgRtwm9zInG5eIIqlN7
mJsSPA8P9winJRxMDfhRU2kkTMhGiYZq/YZzEm4mbQa3E83spG5BBSEST+WYOOoC
3SsJurx1siinLeUrA3OdOFAPULk/CzWoeUflMfjeCr8PGCkUG2nRksuQtLlHCKDJ
uaTyA2nHtuJujsgV9CgMAuK6JUImS4ear4xQcUrMEnQ=
`protect END_PROTECTED
