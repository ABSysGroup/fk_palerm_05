`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TWWzhZHQMPb8acoC2tbslgdM42dbgiDZ6JocSwQZkKfcAvFIVU7OgHZbe4tDTJPC
IoSkiVMb2IdRJHJmnUXQOj2pWbeZobrgMO0ImzMHXKN+HPq19TbJZzdCz+5jxGMV
IDXM1tjoZXAk2YIIUi76V0ZaAlvXhM6gD7bVqN8TyK93JhD1gtyU/Ut9rNwdQTni
4nVbgSmjrb/4dH80j4ZhrXc9p/Gk4cjkZEuQfGW3gXTN+8F0sxfBDNi04N4dKKu7
U0fiQljTTMe52jYt5aT3f3YLDtXxaG2gWgT8LdKWGGUf+Vz2yriOF6tQIkgJ/hU+
knS05lSJYDw4GXk9p5y+yhr/OqrSOGxW+lfL7PtWMT5PWlRWF+LmcgxjSqg9brfG
mLN/XsxJj6wiobN8id0PDMM7H3/nnqvhVacvvK+5gtIgZ98jfD2fcsmMQvdxBXhM
ZsZX0SUA4qNqxSk1Oz+X3X/e1G2b2BHZ3XRPo7FNhk06x6eUIWXszr2XH5Yo0/je
YtNdiW3IM7nENq79ASe3Ckbtb1NE9+r9t9SoryrhneLi9aZrMIKeMTrfOm2uxeBg
81pbJ7hFY0XhEw3hpRfPioFbhmBI76M8g/B5bGCw04/PkHV+A8im0IyEUovlAewj
JqNT7N4shLlENXN9+8W/ugjjIRaLz1X8roqQcWyXRlI0p7tLpyjgJ8zFxhqeENSo
he8vQb86xbRdoxqHuDUP38ZaFxFJJ8Gj+DLoA5dm5sR2smriPLOuXBXt5dweZVjP
4YGW+iPcPkTogsGcQgs1jgle+ARYmbaEtDd+P2ysjOiOYxmAbm1ktkBk+YEHSpB+
bcNZJmXmjW2U9aNbAfsX5420KTckKqJofy6pUBK2GI68PbqZHuOfxGhUadmIT9X8
Th2n4MllA7AYWGhBtfETxL6PZUZh0l7uXUCUCrJQV/g=
`protect END_PROTECTED
