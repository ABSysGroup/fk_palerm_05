`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h/Ziyf+E1EU1txPmFNKMREJnZIRJ1OZ8ooaWS4OVgQOmqTJmPrl3WQJrOuElDOPi
0NVi3pnyRthkkySWk2or0LZHa2P6UYs7TI/9EN2NhzKRCJQHnR4y6CNMM4TeRqz4
w9CaBuTgvA6qx6RQlMV9cK6vpF3Lna5B2REBZ3nCCaB+7Uhdl5WX6R+t+MKzcPGH
jL/CkDro+UwMd5UHmXhqYM8gGrtwGYNWgDFW+YFC+HU5CFu7uKBgW4qMxApCO5vy
dH2GpO/8cTYfpGxyzrCHkEQ2XDMyXC14w1aSQqw0IElL5FKhAizxfrbJQEQH5gcL
Ks2CIh0Q7dbEh/GHV6VkXcyk3LyheVz9r5UaDXvfb2lk2//6uYp4YRLZyYoT8Ik2
sivbktOj7/EZfVYm8cRHlz1PnqSChxz1cznTzNmdLzmnUPUh3w24f0R2IU22Vsja
0b5jUDOxdpefttSSjohAgxxAwNUvlU4D7pMj+dzGPhv104lEtW+s6Jy8PHAO2Q5W
JyESahRvEMC6i6Ph+OGtoywwsbTwQTsZcz4/Sap69SfqTHWImFFxb/x6LEOjBEs5
YiMXXH1AYXt5IDEiIBTSlYAvbS7VhQq3zPMOZFtnPQBcS2KQohL2ddKcJTI8Efd8
irmf7vyWGfGSqMlKqP18b79/YEyTntP5FKtwNUd59lU=
`protect END_PROTECTED
