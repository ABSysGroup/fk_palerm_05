`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FNpiAJhl0vNWHBclOwj0jwo/1qJnfS8AApS7ckNDyOsH+wLuZK8rtFskv04tP252
9uCNv1CH+kLzl1Dnd97RqqNMv7lAFfsWa58DCuW3Z0QQ5t0tP8oSLk9js8j8MjAo
7wh15bn8DNaR50v61jR55ilabljY4tKti9hTyRRT1VOLmGSGmVFy6EKVjRNUdZql
6ntq1pIls6j53qH0kb6Q4KtfaIJgSRE1LPKnW6KKf756GOqwA+6TT3MESM2jl8ED
P2uhHcsW0tNYp2FVqWbU1by34GTb0imqKGmlLorTM/rtf7l0htN1HU0prDuNy2GU
gy9DqH8Ism5ZoC5c581bCFWE5/wSHhr/hgTHSMph0d6kKcwr8sy9d50uendVzRHf
zQuQyRVgGqAn0CqLEiE5rs9IqJBZ+AFnerXzgPsFv9CJVqhD9VrtBgNCD1Q8GbS0
nzvv9M1/1rnIePWai0yLbhnyj5z5U4wJZEIuFA4yY/M=
`protect END_PROTECTED
