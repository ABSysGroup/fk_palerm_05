`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fcZgbGp9/ru4F8bynZqTJylSnIpPIYMiT/xQWSXygYKh9QkbzcXUj9TpLTRTSl1E
294VgooK57bemeDKfD1BUMpPvsj6Bpvg84pkwTnzVpg9vMRScFhaIDffuBzKtiri
pvdC9aaJiQXnizNDGVPRa1NWAu+AHXhsstxhJ4M6a5iXx/VjJb4bLjFBML1kMbG1
oU8WkM5eP1h3R3YDfFDwsmQkdtHPW7ZPzQDFFQJf1BwknXcMuatLS3XUcy6jPQDi
/OFOXNEXGmLHk2HmlTtBGzu4cKQ8RvKbvVZz5I8Cd7uHvDXxi/S6njAV/ax9q1H6
rHhK8jwrSQy2egSv/2yV1JU3fiJwKJ6l6MZbmpo1Lt3b6viO6yFAWh4ltNFZhvb9
`protect END_PROTECTED
