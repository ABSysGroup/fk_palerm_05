`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7QQtzOg2rARTj9EY5urMscwv3ReqOd1SlOkAosz4b7c/FHNwHc5iaEMRsLS5pOxb
kBfyxuck7JsxdK9tFaIfozK/jJY8zyOk+L4plxtvo+eSx3u86Rxo5IL7n+enDLob
ZoiqkSn90makU3oe/QgIXgqGOEZrDfJCbLeRxMU2BjjnTFwpF9qN9vbGIE6BK/ki
WOuVKPYNT9SBZl0kTbqyFwCSRTg0vZMlp+vc2BgNlNuui0wwDOnJzoAuNfkBGG0p
lMcjLmE8x/wUCl5lPDEW37uIhaXh3lQKA8q+VgXvgFdl4sk7kCM9t+GxLZiGKU8K
h7Tc5GiZGNQQ3MT5MZr24zBANOpurb6cl0MxnPvuKrgaehewO6IOoBwzCSRIEmrQ
JMl9BXl/N50WPsiHjHodjy4Da1tyc1cRPLY8wrI58M9O8B+pvXpu+305DY3k9P9i
LCfSwU0wOAS1aEr3L6GbROwx8vJgrt/FNsz4fNk+0V7ln58II0brPWVqkrK22XuW
5ODz/UNcu1iRqdbefBcJUA==
`protect END_PROTECTED
