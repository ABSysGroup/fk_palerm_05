`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hdmp1WwnLX+67IL3YXvtHfPZNdOc6SPmymCzDHA0bwEWt///M0ErdY+LynOOGPEi
gwk7QUuoSzbd2W6Sh5hkFiXFPySqovuo9ySwCd/TfS/5H9LBKQTMUuIyXgzoCoOK
p5NQJEBaXCqXSHDGMjY37WAwF6hAqg4HzRkvH473gTdIdamiDEm0YfT/cPA8zxtT
UZry/w1Vu/v2A4kxD6ECaYZHvi+adHGnS7I3L7o2ImTUBDfjDM5r35C+JnlneCG6
mgSZf0bdh7PP+/DAob7GjYonZNi9C7HBnGe6SX79jUtsXcdb0nPqhRJOcvCtrYJV
bsqG19YF8EgiRLxSxh9itBHLDxMeYpVbHLEDAALVfzhzIkJ89SBopDFrVl3788Sd
JNaE0JKSNKLswltAwN4kBRFnSCxml4PF4OmWYEa+X1ZutXF9xR/oFQlx9KXUmqJ/
Ia9EQWmGc2ypbbVzj9Rw/POqgwGNzOTAl1jivfFKE7k=
`protect END_PROTECTED
