`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xfeg3ctlANGMjFst7zhbM87b4nFeVs4ES1hf4Vg5cDYt1f2h3IhBZeD4DgkAVtb2
kNCHoNHfqhkopgQ5gIpr72NBRQqJ7VLQFE/dgjyj7UVxPyykSKIkZi58LZRau4Zm
wTaa1Nwm8FdoxJrEvmgdwTu/rSuPCfPgK3KlONVgSSQfmhjMeIx1gUKtn93/7R4Z
g7cUrb2OTVb1iwbwQFWw5hmanB/t/OX1NDjtXE2i7wjfEOWsQJPWYAScG2Bkyii5
hd5KAUWGq4j5qu1Nr3bfgg/SpAwdR99YK7Ba/2rmbnU0S+K+XwV/BqmubO4MHqqX
YvdNi2JtMm9wx7RFR/P1NPD0K1ySF09B1+nCz/SmCGlko8IWFnPqC1/wPAzA+O+v
XAdW8vnq53vy5CAN2XUWVpHxVpR8pe5i+lUOK0bOz4KGuDsR+dbwj9jL/k784/YA
UtAilMWdGPuG9aPPnXJHKykbQ3uOPRbap0ZWNb+oMrrH6KEWwnbiGrM/6K0jlpVq
wJLJqMWBUs2iWF4tJwbb9GvV879oXy/lZiDjQgZwbfb0Cvth9XsnYq0t3Q8Pl924
5qfNpHzLgIVwkwXEREgTJbQ8oiBZAohdTur098mORA6maDThpZsaHTX/2tTjHpAq
VphTCK9IziePJrW9L9XGzPHqh9T8lJAdCVEpR85XDngseAaUItd8lsV7Aqh4dhiB
Rw7KkNtT8yEdUk+LC/3o5X+sYDc7DRP6A/dTc0ktV7+5cIf1YmsvlRsOHaxJZeZ9
pQx5+qV7/MitkX0+WtnrVeCEwgoSpquwIsf6ce0NCH/hZbBz1zNehcda8uCiwMSN
Uca/c+pZcWDJMd8ZsaWPDsiQ5Dok4rU1eicDTg0dOrKURbeH9Ag1nx+eiD+AKkYg
+d3UaiHAAXaSNCYtrR6IyKkADDVsRt/Xa95PKg/piam7ScnnZBrJfaVfxFGbB6tk
di2QlfrOh9VQ1nSJM4x7W6ovc7Y/BOI96PurQXZC0EVH/Tv1Va1s/r6iqz89PNuE
4egLiHPn/AcInRRruAtwiyXjpGLEIWNoL0CjvYAYuMUpVgWHpnOJwcCuR4Bqf5c4
Ka+Vk3GJfkq67xbI0HuafZ1/mxd8d+fEanVqxzFWoki9RSeFUwRk2b76xQW9Y74a
D4LFz+K7Z1HEXZ7SD4hE4SEou7G38yHIplBWyp+4JoHXbgqWMMFdC//rgy/rTfy+
bvaQJrsoNRICE+dF/1KE4Cx+EF1JpYoBQurRp0I9afh22WiMoYFYrw3hyBFP3dmg
Fw97D05t4ygpvMIDAYFgm+u71DXPviAdlcjDOT0yBY+pWQYZDYirYnaxpzpOQKup
OP+Lx5O0fAZWTNu7BSybCkLnftT7fba01Ia9gKEXTEAyJTSFUjPsxvepHjduCldn
0Y0fWmhbSTK7N3DNhVBvCIUu32z8mv0WZCxiyn+y+3eVBNFOMPgziIzJNlhU5Z8X
J7b+sgto8o7N3IQBBXGv+zBB9pujoplHmVXwOUBOCFX6ofRQdmgZ20Y3PYo+7Doo
eTp3jqVBAPfKubwcAUCc0w3eazCihtgOEfoShSmLDxF7/HBOm5BbgV9i0n+Kyexj
TEUnJteVNmH1edYRZEqLaRn0FgXadpsz4GT4ncIANUyndugy61B6cn9foOAIRLQI
mfaNyvC06YoA7nUMXc7zDIw5ipMx3ha1MSgOEPfLaqlDPq8cg5jD63oL5VxGwcY5
Vz8mr/MQsBPrS/YVbE2eXx0n3l6tk7vcVXYFCdT06eTEzXF6fkSg5I534m2f/Dob
dOVRj/WOzwyj1WOpbVFshMkCKJq2yMskEnajQ8cLotoYXLbxkr31nnrklu1RO1mm
cexl7sxLWHiokhKkXdLl7ii0iGtaxvnTQZlDVhLPPdL0wGrJ/p3KrU87KNFGtKu5
W7OJyGES0jtYZ8uv+S1TsOjUkZIm7Q85JrctRq/AOP1wsP6+5yrq1kWOnJRgNM6+
1SZuXDl+IF7HEObqiwjupX7PNbnNjjCnBj2Nc0j+vV9SCTw8TowkjBXy+ABmRCP1
jKb8Ijf+ZsFlOMpEH8L+BOzPeXkOYckbUe5m/vbpjf+yt0mNVhuRnlhC6s90lzAx
hIMI14u76VbI6IwYi5StTe90UdgfSGm/8JB3NwDQviKwjsPobcKum+OCx75DUZ/V
aF0EF1r8j7kmx/XvvvRaNw0rHKlisiMqknkTP1m5EmnEJvnCzxUrBAZwBXgXX3V7
TcOCufB2NWuU3VE822A59CxckAuSLdGVM7PMQ6N2lph9ctiTtwu5+KW+TVq1ipNF
7RcM5BT5w+0kqM6NzVu2TnG8/gMbt4wL68WdvoK5uxrEF5QHEN14W16Co/Mrokqe
EX2J3Boo+ekrujNNqbWQFh8lLyLKjhR4UMkfCxy0LIEjAy3RYvW63iQ4iuCJ/hIX
DRelkB0NBQUkERgWLJidl+tzDx8u8MsDnXBa7zALDSof91+ZguJR26TsWlJ2SqWE
Cld8z0UvQjxpzXJmuz9qtUmtS6O9h8pq4RsJFpGqt8tKSVK7wMl1iiYaeZaH1CXe
7PENN0iyJfPtkYjTHmEOXfvcCKdz25OKuj/1in81nL+3gw5x+rUyjLP6THytwuIU
GwCdLobJ0FXGBWNxkzqcg/52NwERQrYT7fRNsCzMdmm2VlxScwnAS7YJYsXKIMG4
`protect END_PROTECTED
