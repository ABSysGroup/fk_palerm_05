`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ccRxCbVPCHMu31oJWU6TBwXD9Ast+fgDyJAUHKYMdZlJwD9w4idwTqw/YDVKozY
Bb8ps4pm8QEqPEl/C1iHK5QD2likKfewwd4aafefK5No4B10oPVMm/TawAzx1gxx
sjOoic9P4UErXXL7qvoTnTHAU2K9e//+M7tulALvt/y7pB9Wkk56/TtREVGEHcor
RQblOvk4lTK64UxnOTRxXS5OkQhvAwUC7FM7tpcHNPKwbsoskeZmdSlFVQpl+bhx
VJi0r9Vy+7YGvGIg4ui6ARjefIzURHuFwsiryaDwRcSsuw5Kg6qoZ3A/c38JDcZD
OChfdoD5FqwysyorS1sWrswyPAaqAsNFWpviEo5aNdK0M6iN3NMRkNln/W2F+HE7
2P7NUJ+o92q/EYZ4Ko/IMVXDatsiL5pTFB/1JqEfd/0FTJgNkTkJFKLcGE1Asoad
umIeY9EEr/65ySJWiUNrBriqb2k5eQyJClyxTnpVNS8=
`protect END_PROTECTED
