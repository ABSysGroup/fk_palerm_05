`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
87KjI4DjjUIJLd7SHW4pHv0b8BkvwtLCYF7NUx+ZFnhMRMqDO++IM/cBe8zQYe2M
Hi+Wmnl2RRTe4hHSdLk3zfz/mPdUAK3H+h93X0RBgEh5JToNbljqFEKBqisXseYl
pTpavEyIsbuCZ+iXipaN4gqjpOm3uBj8mW6hrqqoyju0+ku/lhH9Au4+wlOhzQtu
4ywbbj0uLyvBoA6W4taMt5izvxKgML4zBzdYIYBi+NiEsBB06kMG42GTVDO0lLqH
8lhKikdt2dzuf9b/d1XoGbYxxBocjiWQBqAM8ASc4DpStQ3MxUBfaWu5m9Bo9AsO
Bm8p4i9dYb5ql4lhaOl15WlL9OHLRvgLHKWXwO10ARB0eG8aNrWATSL7sXj48o8T
VG16unqVRn6bknimW5Ph0nLbI4dZAgO1uvgzhAiLJujq5h7N9mR49upQtMFjQp9L
IbSIXVdfWnSwe8bTKcqCpoaAM9ReVvArbdU2a0LPwTqVMPIi1HlG1R2Jys2l/ezk
YX0jXoH6MhZCex+w5YvngWDi6Uy962bXntGC/QOGEMySkjDxOKIwpMqGcNrMam08
WDx7p854ttrKZEbrX/KtSsY8dzxFtZrhx0rmbQFnCVhQQ6YMKOHxvzWdkhZrkIOM
TPee1qgfP4QyWCp8ez+qFkPtk/2VOjilScPFZt8ot2acHljJS9rlmjkjYfrZdP+i
Z1bYKv5k55jbbYz7MqDfv0JNJ3osh0CY7bdBRJ4bRu1RAvb0Zwkv/Xplss4+O/jV
vc4i/ma6tpR1Bb/yg7lUPXaexo3Chv2nQ0vpcHrUjCkZJ3MaSSLRsygGL6NNS011
jvziEvt6Nl/mcmj3PCfbrXllxicfRwEhJ9OUuF5vDBJXLfcNV9nW8hD0e05J5/Tm
q6Sikwv3elvfX/FrrnXLJUWvPIUwOHme7lI5U9EyqupLGjkdYR6ni/LnSZodxxwY
j1vanJ6I3cFAGNEqRAsnVVLTjT+ushzMFm/Jq2HGrnqDjcFZH5mIdOsyjSPYGnbG
GcH88GMtRVHwoJpox3sdsKP52ed2Z6ZyFc2j4MIfjPaG0BktQ/W8tSJoYpBwSw94
6Ly6tNf8mD68stDphKD4Z/GSgthse4bZvw3lPp3uoJSz0FjUa1Nw9BWDk5Qf37Vi
NEJBbdy4K8XqKq57uuTL5F9kdf5qo+xxs8m/v6akQWOlg7GigNW77gWhF6NrknCt
rWIo8iF0p7J+ifvP8iVSz7BZ1s+XIe6ZX8lpuHJNd3mL/21OT5FLn2wMBde4F5Rf
OHNkhgougzD4GIu7tkgQw5v9a67rVl5LTmJIS6LiOgi3F3pArENsIly9Nfd3Vf/c
wS3u4/wj2c7oVaDOa1ud8eMUHHiW/PpjpVEfYQ0cjLv/fIDo/pOSyhWK3idXbPbX
0xTQCzxafmLlFbVy9NV9Kdv++quEKOWQ1NPoPXTpj3lP61PZNXfsHnjWwNOQU1Qd
t8iYi+6bmD4AihwRlkcCi2ZPZJa8lRPGgvAt/lOy635rQpoMm9sUNVevT9/mM5Rc
BK3muv4/vseQZnOX2k0xlRNBtRt8mt2JEYrNEe+kFUTwG2+r/kppL1q5nxypilPP
KqI49EMJisIzvwSZM4OYJHHm3N88xWvs5/lXaJbS5u+AXlm4771PB4ymt8NFARRv
nqLy0ANQP9SXDd2QV+qXLPMvMtIFmk65OzsiUfqi9K34IVBrzusq1j/keZ29+Dco
LrVmwvvv+AA87zKtGAbGWuButuDw6WA4Vm9x9kY021bIiZEVCS0iEDypWELUmD94
S3NoTSGttHmie9zVjgaNKz3i3Ef1+6PgrG9MGQck8ooEGCkgubf8trkg2p51QV8Y
XZBA2Te6jRFOSt7UNarWPlOZY+hyOVFKhXXl8NSY6MhpfiKYKs8q79lOhdzwAObi
lWP6oqEdlVClDNIgh+yisSGbOCp7W/vBrbJP6CD2EvPr06HfAfD5LOePQJXslSrz
Y9ezDVbE2VSwuPMAs0wtDY/9x4+S0ub5hZm+Nwj1JSUgqqa0x/FfQbGfs0M/pfpx
njboykX94UNsKKBf+GkdHDGOYq28ZXOxfNYSxXhcHULSCkqoBoM3GDTiYJ3Vz3i6
nv1ETlKug45pzk9w26srS9PQVU28j8KwKU127n/2oms8EdYv8QJJYnZDlK86dpkw
h73QYSnNqFnaWv8K1p5o1FPT/j8p9lyBr1QkjGoljM68Oi7Co4qHgHqlznOPAxIO
BpT0+Z56Wi26Dt8ex0p6cvD+9RqNVhb1vafnlVSCKFSxQZ5M1Y1wMLq1/TzrID2E
LRMhyEjZrT8NSSzbJyv+/lA+APAm8s+jMJXa8LJR7RMdEsIAVv2wHRx33E7j1vXb
wvhdf9e9cGZ8k9p9hV96sTZACdMOsbO9o5WC2yAFtWYxX8GGZvwEUJU/k/2yVaxU
oqPUb0U88RIQEw6Pu2NXlCOsvctqn262cj/9dsTQJdAwCtUcA61TayVMTu9xlaIX
gsnO78YCJpXXzYhh0F7pll1AflI2OGt/vu5zXbXYnfDRSTL8MhDJmKVKdMqLbDUa
6y9uzZaeIwTD58T3bQm6iWW/QhK49rb4c5gVxuDzGGC0ZT/H+k1sY2agN9HnNyY8
aOto9t9YEb4a2wFBYiqBAqk99lXdSeg4qUeuds/LhLgaSU5l+f8+Wdh9vX4a8cvq
ia+IvE6c1AwT5i+hNHZG7QK1dyTgn3o375HN0mYhVRTwEBdIC93k6O+q13bRIel8
Qy1tDnQGAEB7tR+ID51zhYJXbeCvzZtANeDJ8svFUGQvI8oueaQhJLwL0WTyH6Nu
lm2ocLJTP/b+lNA6whWA3j2xXvDzzQR0tl05o7AMOqJwyz7zPTE1O0w1lVjVxxdT
Zg3GU00drGXP4j1utJP4gpSkPoeVLUPyHmpc5Rf3nQqUZ6Lz8BprA9ktlNPVaysE
3j0dtIzBkirfpDTOTQrh9CSZpkNRccAwRAJAkyzaAoEtrYMiGrHGwa17Y2wuwbL1
jqH9DJSGPRQV7K63bq47m0CkGFGgRFIPuS6b4UA5wP0GA5MrzgQqCvujr4WVdy86
Fo+fbF2M5hRyOGZHfdNbo1Z35bcOeOe+5H3OcaraBzoBqhjQZvS4oj+IFjAQbQ0F
0RO5OK6+8+zB1SuEXaCAMg==
`protect END_PROTECTED
