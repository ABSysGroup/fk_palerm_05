`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jWPcqFq3kYBRBT28Jpjh8Xh6GTfTdUjGuNhky0+D5eZveHBbcVqnDbofui/3/IoA
UQawA2BBGYA6JTjef8pnfJKcNAOigqLbqdZPWjzMSV3cJblkYEdnTNjcdqZ747NZ
ucbM4GQeSDgbDZCmQg7yDOa5r87g5UStKa/L4QmMRxjcLBQQ2x3VgJ73RymB87Ld
ioN8RXuhdhRfQqN+1GhlPcsW69CiVM755wirxtYyP73xjHgW9kHw++PLDjVfn+H5
fzXen/8ITjuEEUQfZYH9QXwDBj2fk6GCHjTk5XYLnWsCnVY7AmmGE1sZLDFMRH4u
lrFPC+tKbPMn8UIHJteIhg4kvOCflKTO7Zn5GIP6FaZiPJRHd4ghtOtcSw01YEAT
Xp/ndCBZPuNG+cxrpeUraQ8vAD5TtDLr4Ip6147bFVABOsj69rxl07I6ng6j25IA
ycC78VvRPypnJKLzvDVAKWloG1uB4nbi6LvlnN4+2oESEKJs8Jwa667mJ4+WeVKw
XaY5LxnDcl1pfuWP4JSBqHx5C95VL7UXCdCljypq8UNY+VzDhRlW1spkicaRf4nO
HvWfbGM79FDJEW4QUwXQT/0cpGPPzVUkcWHz6Ca8oarfyVXLGboOnRgITzGp7wCG
tIPQss4V73i8tLV0/LqUTGKSm39IP4WVYH85SzJETM4+Fa1F52mTxcE52Wyt4D43
/WOFT4nE4gxeb6E4miEzjiEhl7sstdzI7dCuAun5rTT27dKpmctNltJjORWGOnq8
8n8yCqzJq6SrfxBYljNY3nIODOpwMenvppOxBD+lFxvccRcg9spwZjH+nRwCKlL+
e3DHd99KzHXlTftxRPEztStr4IziDeQuqjWxAsfiuhueOzBYkW1M9XDKz7d2ZZvT
6fuEyLjHuh/WYnjkY9aKfRvpVwceVSKd8C5i629V/Aj3SidEPEPR8fvIGJ20ZSCQ
YishfXNShHsFZtwCvYjAmAAOFFkrhZJFuZ2P64mdiGexjxrv+NngRiercI1jJuY0
k5BBvuJJUFSM0umN6eNuamT6VSNuz86JbM/V+SIFr6U2obzlXbTirmoUiSC5YDnI
Y8ovzXlAaLgLwkC6pbnCkxM3PLa78ftW8l+jitDwGTv+j+Kmb0SEF+62q6Md8dos
I6l7pUgqf85thM4RaRf53Gjw8JWjkcTrdwSCeADDlPz7FB9O4BUXZyj4R0damNHI
LPAPgwf4L/JRy5/9kFWWjS85f6qajok/DwDtvH9ZuBzVmIUS1UXHIRFV4Gd6bmvn
k7JY5ZKDoSkst8uzjYfpMA3wv/P7JzfEGBleLWWRYvsnlAq/9J5tAwqBaFB9POMK
Oh8FH7xw8c44wIz63NR9RpLIltyCox6ysm2h5ykMrZWTwXKA7/77jlVk9yUhUuvE
7i5Ip+f24anydHK1A0BRRbiLBPfOb57rY5ZxGzScmzh8OkKbH8Rbxg4TsLvNtOJ3
HMZvPkxQkwiiH3irEn9b0jMO/+v7npoIrWvk98QfYAabAgaqA81hOcPEatQluiq4
VT5U3AlnUF0ZWKCwphYspr8uoGOyNn6/Z83WQ1hL7ivOrFXU+yPX/1r2OoGaHQ8k
4X4oRdZBsUemGhSe5XA7DrcVyRHTbJmU0H7hhxXgy4KQ0jWeG2aLpgtCtOxGWP4B
+gIDUObDnsUXIE47F5/t5J76zFOCAxNgwS379w7BJ4EweWEE5skSDjvHIXBVogo6
hT7hgP6ZAI59WdBfLg4Uu7bWTnIHwt2R1CDkNF1eBuo8DRjol41WYSI+Yz+fUuvf
4xwImxTF4SIhxf3EAEWsvbIGu38No3Gb0AewdcJiIOhOKAMVu4JMBRBwK8zu46IW
G6kcmTLQnHcxetKxPCMHtEFCCpR13N0HKdsptzc4Vc/iWj9jCqZyjOZyJoqg7eSM
onBjgWg6Sm3pb6vjs7rh4n0Pj2IAXp0xAzYfuQ2MDA7DQSAx7dMIeSo042Ibe5O2
VIbecAJwBw21rU0Fs7fpVC9DqYacPjuAc9mp3XNxkCcgr0oxTiaPqTWlpAU2zKqO
quGXy+nmK3KCks9viKHHeZC7nZtxnxaTS0b3dnE/6NG1zI5XzHI1XxLxvrTkRqCP
trCG6R/v4cddR/wHBNnHO3ayt7l1uHphsKW9QYG6gF0T4mXyr0WDo5yVaDqbGRUy
Fn6JLSV+1PAvAT/ZoAyBIlFnsZv8GrqOakJ1viZT/gjminioCIh2iNxB5oIybui8
a10vb8pojfJM3gJe4JkAwSUTJDIz/HBjNYoSOuIRZIPWwfalQqytwEiroINqP7rK
khVBO80a2detgfB8aLqwlXvk1nCoJBMjBDXXSwNvyE1tD6dWFc0f/vReWNvNymj5
HTa5A2qfbX6HkFArdWCAn/pPIWHBAEjbcpxUjkyUGhrK/Bnd4BeyY9cNcBj+MKuU
W7quflva19U4dfAGiGgrYWJqA/nxlkt0+2z+CwOqgj/q49M632XeVXM6hdLIpOmv
y2NLQubJSSh0Y+X+qjK+SfZsxDDtvfYrYkOdQtzaJ2BH4PEISe2KUdApXdn4Go78
v5ZC1PNmD31WZOUY1Jgirmzkje4OmyLfdMBxeSWaKKpiLzaRKhH/LxoJ9lImFOsn
ubA0e+ixuqVT403mh2VG/LWX3T4AT5YNclnYEhHHWpDbRPTQ603kyj/vFRAI/UAu
6tx215ESr3TWfptI/Ivt86Pvgm4aDSqki9I3/NlUpEHeMVOVvpONC5tRepnZbly4
5fop/tIv9xC6h0Bsv8s4sh/mc9QPgr4OMFGZTILAHdIdpKgqLRwPW4pIyyXcK1vi
OJ/3/b/jr1Q7U+3z5p6SOePO7gonze4wHaX0lymutHn3kq+Yf0dYRRULXNCI/oF5
bxX2ujgRpRQAl4p932yZxviFhos1M3rOMqpTNffayEGj56xIe2dBwPITNW9QKN/Q
bIes5a0BLoYu09G65W+eVCCn6H3aVARkG1pldxQTzrLk+S1g5NuCftq6OfHaM54C
+021Ivb8DmSQ39tQ7vJ0HVZJbMBZjkaHRlMRr0+rO2vRx/4u7IXh2QWKnNpSBRUv
l4VLs4TlszddXEJ4giHCPX1PgDYYiklPAVZihnzpPcfbhN5TRi8B3c/oyFquPgpH
UOX/KxxphNDOLJs2fqb6AvfmcODu1Ca/E4frU3JHeZRPdGitR4SsC4Z1T1HYAASB
AZNHTRbwJdAJDz2Ai1DZdamfFigOCyXOQxo4bbZvcIl6meuaS4NFB5Ior/Sj/ltq
fz1ZQO/uaZucIrB5O1/SVAQbzNWn1DW8YxXz30uu+OdM0N1ecaWL0yi+zUcgpeN3
mj6swRgKywrQ8Go7IeEIZfEHIT1qs+ImWpAHadmLvnyurgqrMrWT1pMQMX6w6Xs8
xGah5aJiYCRlvrGDRapb9JQYzieduwpMz+YqzCKlFHMgi+J1ghrQVzriM23PaOTq
ocb08jBNNnIdv28WDieqhEK/r+dOZ0wdU0a6gZnwYDdnQOw5gc+vEdb9N3oMgm9J
Ai9FQZPR6PzWDaHkNf9UX4h5LkXuuoj9I01IePmE9aqHhd1121E8AykuTSmVNE7N
fu/MOlfStNxTpdLowEkB91P6UpLzRcG562m2nV6BvExKDY0gFTawUL8RTxLg0wNq
+Ahr9R99DKZKj0OiEvJizjIVCjsw8IVl/7i9O6TcecIgVrp+dZ9NaEgAWWFZtW/T
c4oJHKngsYiz6DcXCQkzJRkWD7gfX7XbYm1oNb/ld6fU9EC7Y605TfPHBIxjKwt3
6uWZFn1ryZ6iHjCnr+MTyY3lNlu5/0tnQHPNHZccwGdvZpZvLZn/hRqvRt2KBssr
7/h4GokDwm+tLu8rGo/viKQcafTMHmzkztd2KIjjqqC0IUa3vmTInbeoss5Np0RA
Xj3A9A+kBJ48//2/FwGIBAgADKWlqmz0i8tYrKVnHwlwHB/auzSxC+5ZwemEpCWf
Z2QALVz3/HJXPlfXkVuX2/SdWq4m9NBFuFMajLLJTq7iW33UrDbd9rb6y2rOtFNe
XWGjjKjeDgzdzbCI/Geu20HdBmZhxdn/2cwaWBbXGbL7gUGR2ej7ilKBrLbQs9ZT
kj5j6ptGhStQbr9cunZvEhwrIWj9jy511Su462GLCTAXqxpBpMhV2FeAlpuvKtKk
DTaKe4LHoO6TVSI8do320MYjTgMg3xGX8cJGPy9ntmtW85bSpE/VyABmGkMQL66t
8PYOT3fQdmxQ9E5GLiSU82PIwbtRUZ8Vu8gPiVHGwD78Jz0BxUPgsZAYKp9wGQmp
bcMyV0KMVm8yaNBNP2gLlIW4iRfiBtSP/vnlr5N+qnTFTk6FQwZ4VtRghwoaHvUA
NQekllDOBKlmDjXpoSDQk8MjLuz4/NMuO11Jw2s3jtxiK8pbb3hYev7dNySnjALw
jh82SIPX7LCxG80QubbVTEaWecYaBqIWJics4KmB5YBHCxtCDMI0JzcQ/1k2hi5h
3d1JfqG0F2x4CEQSOdCdY1LcO9/1Mo+WH4Isx6ESkyuVdNATe+faCorTgTWZS+O7
FbqTYW7/Cpt7jJ+V+s0+V08fUsxwe26mOsaxtli3h5fIpRZUgs0LHGzYopPXV4b9
N7oeU6XQaVtnG7m8cyWjxJGrgTptY281459nF2IqDQz4M95gbCrF8ul2uukn8G2V
h3v9A7W5+e3rBK4y50tZ3+cneYe3g+eIVSgK3Q+9405CMR8i4h9HbOpM50HT6P4n
kBBRbic2PIaNWtiPErBDYqWm08vvA9UzVCm8BuEHY3CURvjLvIgxlQFaj39Pxyr9
ZCAh68v1Mob9d12jK794FJ3JFynz2G+Bd4ZV+Ar8+Q5X/NyqOH8lpt69AZPH+x1h
Pkh3mBz9dWV/9uMCd2u1fBsQPnpslKU5FFhDz6Oq6ZvQmNyhC6Ow7o5Awz2qvoLF
33hyIE3y6KHhPjXo2EYQ+/rCRgmQbbxTXbbtp5V6l4fUWhQ6L5WGF399ojZAloOK
PjbRpVfB2ihUlRhHiaRu87lZ5WXfux/MXCEDrZjQHMn0ylonrJIl/TislZiv5ily
G3QDIcg2wjm+pWL5xhOPm5WJJWV3hF1LEjbtcu6yPs1Sv2JKTH/N1Np+mJyYIes4
tiGH+LyMhtQyf2bcqiMVPkXN5SAntuzqv7c/ML/HwB8YCYKVf8oxhjat0HXaLNLR
XjIy0KbJUSf6qsevyWBkaC+deBYIX/754ztLYphdHj4W1ziIt4FyurUuOnkYA2ur
QmQWcOupU83Wn6abg3arzH5BRC8DdnXHKdFSoXZ1z4aaN0AIvErC45af0R2z+aEN
xOlzzJ986q5jEUhQ4rMJ4ukI1lQQSQowmvBS2bvZpFzZbZ7JlM58zWHm52k7b+7f
a0wgT5ebOSMamRpIflRMXOxMdwH8lG1ygq1QAOADB+G0B8gNBAr4OgFyCTvLYslK
zMxOIywZp3qpLZhqfq9jmkRSQ7AUHsVdRWa5sC+nkm7+42usPX1mJbsiGAMUggoI
onWJ5f+GLEvy9iojHbXiwAYO5tQQgd7mGDQSpIkWfy42thk76eqJiA5lwvCPSw56
zl3CB3SC4EPNqDDKr734fqh1kqJ+hvlIIAo6FumUnyi8ERMs09/1BB6CYvANod3+
EjQv5x+ZdRSKNZoQ7gLX9i6mMso8OnnrxaMC+rtcm9QyI/4mMbIQG2VY3C8NV6pa
xpcR4DkUSw+BIYzlA5xpKfcjVJQ8EkBQAkx8SyRw3COzO3WWyRiAfFOoueWVrr5U
rVCmBbbjFqTEJMlkwyDDd5r6kgSE+6ISuRV5sbCpEjVMa3tr9ewxeeXyzCrKZrSp
rkLOj9/9YplchuvL/PLC8ntR1ayZQE3WDsVqm2Br81edpY685jH4ulSkZu6dIp5D
zaGqy7x4dffURwgI+Sj03aU69iFtmquUwuoruSV0GGpNNU5WQwSzD72vzMMLNn4+
YnOfJA5tEkBYjmhdnMoNt7rJKZg7edWZIVWWfp/SA//ZERmTSdtYkGEvHmsqSJrM
WeUgH5i+aY7icy5NPDiCUNGGhgnAUJvyGnnJxvX/li1rqjVMiY25amp22dZDs0Yd
qimqyjhCbthomLbQ0dg+OR0hmkS/oN+yMZ4gy0GQF1hZWU7Pb4qix/y0kISHCGAR
qBYbjMzqTxy2thP1JRFkIuM1AY+v87tcPKsQODQqmYVmARp/2z6RBrPS9Yd8f1Wu
GzMIiNttgZiyCezw5+MQ79DTXykNjHU60yB+eDzmUxjwdkXTSSJVMe5h7z32RyGG
K+eUg7cmRfNBWJDVhZIimr27d22DqzEkNit+AhCIGZ0=
`protect END_PROTECTED
