`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oeOJ5gFP8LE+otMJr0+oUA5wamYHv8LX8ySaiJvxCujc83WSyYtTO2bEkfHaI9Qu
wf80wA12zETjjoSRHg/esOjdFZavdEjg27PeQgqI8P6EW0jBL9fcAwllIBqrmHHT
o9ISkLkF1PGlkfmA5iEEIzbz5ZQrG43l4+PigzIcgo3j8TLtnM3AHgup4chi7wTl
JXnHsqoe3+elQjvvUcQUA/BgwDMPYaZQ3jEyTqu/gOyn4dlKwYZezG1jsLDhisaE
Houx1hXUMBlbRYLTDd/GR+VjpiSsb/iYBS2BcbZVRJ9Ec3QO78Gy7Jf8ML7gt+uj
jT0/Jr1XZ0+/5twwSNvTpMm6Lxvon/2Cw/BtdrSoxvnLsj2X0DFgPlfk+oICJECX
Jr9gyp17+yXgh4p+QVXachXOum/b9JELV6N3/HQx6Iu4gBeJ9e/GjP/KZFQAeKyo
XcQY+IAWWAPfp9R+3i1S6zvr+1dEaFvFL4EoUdH495xGOZ1iHvlwKPoN1NkMPjZ9
1yJ0ZCaDhAehESXBgcX8kWQdl33GlVDH7IpNaBahvgi8iw/In6XWTaZcCowRPZwW
NCddTkqJTnZ9Hvc1FgVDx8+905FzHryeJzVrOGoqfc4=
`protect END_PROTECTED
