`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NLSHUOG/WZ9jc2nhVPb/36srpVwKyutU6A1Xo/HFxOPDj+pK1enlM8tCRVlpEmbR
7G4hh6ikdtmB7HMW7fkijWmnbdf+6GNDprC8S3mRJVgBzq18M+3Dv/oB8OnlXdhR
yVe3NfnIbMt1LQxX2wvdYOoEPouAj4gJMjo5prnine+ZEXhiu5610K9Ex/iubc+H
bx6to8vzG1RzkLNSJmktQj/PUzyJOVMUH5R+VJQheCkZgV1dhfvyCRrmDh847XU6
uuIyfj3pKX6pzKE6tVL63X8wi/CUAswlT7m4A3qd8d6qjle5MjDEcwLDeLX7tnq/
PC8qbULWb4H8bReA1M5sLys2bdSlWyv1QAZGmdTfkJrR3gNs/UUGiY9YOykInvIB
6JFzprdjKFNtKK529d1N344S64MVS8NAiICtdDwojI0ievgWqFxvDuukFPT2FDyh
ywtv3MufSU1dD6P/T6wRUTedO9GaT+BE7c6meI4+j5zJ/sV3DWxBOVhlf8encmNP
qQmEy8Ta/L+rlYPvWFr0PMA5i2+HIvlgI64DnjPYhzKgKe6qVcz+UET5NVqsDHan
E6+iWdoLI/kQ6k+cjwsEFOBWU03HQQslocrqo8ickXZSdXk4TJezjQJwT7NRH1Ey
vDTesNA7Y4m9rL2q1nHmYD0wr4RDKi+o+FLdbxDL3OcU2amrCFp9ntJuyidH9fOj
VlIZyIyeZz/YDbaWsZ7IBzrE20yb+ruFXOqHG3Z5b++lN0m7H8w9964/RJoIqpFt
MVUA4hIJc3SjUepKPCSkKweIi5pDtx7vNv7jkf+hro4xp/sH/cFFraNVoFGC34Yu
X1LryCHJoNBq6MzPL+Nvo1xlQM8vXzjY8jb0JG9h/RkaZW/pR6vVXJjlo/hFlpXz
Blcr6N1CsEYt4jHc59OGHGbDT6vFJj/60uA/cQjuLhok4pE1Pm3w6KKY2SCzUZY7
HJnTC+7FStFActRQAZL3Xwutvv67A8tDzNXUayJ8KqW+D09l1MiljJ5XZ/SAdm3t
+jiW96O2Y4XRuck/comfokP7WLk9D+HokUOGm7Asg8dEmoJQRXoYvyd7sm9wTCgV
y57DBe/sujcxmx5dQZjNkce5srpvRY8QF5q6/LicZYxRpkRgl9pyvxXLXoAn6e67
uFGRSOQ4UzCFsWmt5/grHAa0t3kUSJYybC1ILUxGy/TQrWBPpq85WRO85iwriPEA
y30Zhvn2CF7kLNQhQU56QtAr6m9GXObq5ZEASzfB67iF7uOpsz1JgpCwSx+SH9//
1KZ8JLtinhT4egDilMMVACXtT7Reo3jj76P0gQUB9BHPtxjkMimJpuJni2lJgpca
ksTN9tDbnVNJHLhrZ09kVmtJypIiipwUa9lNBT2Y8p/EKWRzcDV1oe3rCO6lgS3X
YMSLGEKbHNo5Rmqx+rLp5xYf/XyQ4CaOgsZUta1I4vn74J7WxnRqKJeho1HwkgWW
arYYZUqzOhQXXcEXNrXZTHOHXdl3RpD4J3XHU7UxrzmpjA+RD0SBF+Q1BJmkjpVS
M/Wq8Ucg7xrHKq+xjQwEHM3xisHjUMDKx0thkw6MtLNxYRP8x+mL08my9x3g+O+t
QH16IN2Rs3ErzJvGEqdNPd921Cw0rskHW/VuuejRFM27oL6obQIxI7mz8BxmyLJy
e0+WotIMj/DvHBoaSCAXjfk2BWED3Sy+O3sXekywif/iFaLzbH7nFHksbpFJimCK
CEJN4SzODRwK8TtYvIb8fKDLCUpfrUnA225zmqIgwetcQ2+QIA0/nSTZGhhqurL6
OMnq3mRhnIj61giTHq0VEY3jGxiOECYBGwfark6OzxAIkf60eOSQvRaEpDHNf2Lb
74Iw+P7wtiRf1n7hzKaIiTKiYxhfzXn/gNuoRV5FVjZxj24Mamww3GCtM5Q6u4dC
00QKEwvmNNGrCKuQiWPN3w==
`protect END_PROTECTED
