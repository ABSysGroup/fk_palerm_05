`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8cyKm/SuV2rAbotVT3/j/lfF/HizA7PF0PMtOuGDoEJaz5p8Ojk7qfhMPSybcXdV
wUuNXyVpUw4bHZjad0xsWkWFF3HkwwMCL1eDo1TfotJ7/pEoHNcauyQF5Kd1YRQ3
/8soZ+M+Iu8jOMChqKTfF4RICe3E2iTp3Jot+LaxspiHXJTR0rl+Th6U3XweIAEw
jjzr/b/LqpLjgZwPrpi0QekN3PfweuUAfu2C+oGt86z8Nnygoc3o5gjERIFdpIon
RuVR/Z6FeW5cIAEhSpgEKfUw9r4LeIlU5C2PRN0IxUU=
`protect END_PROTECTED
