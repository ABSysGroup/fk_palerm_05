`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ulqBaHSDMy1/02pBoiZsYNm7buQQcAlVMh2ImvvZPfH6ko7zEL6vCEevHRTtUYW8
NFYYq/ZH5MhqFwFX2eRKF5kyWesThbCTHI1HrKZNNyB0VDWIUbEN8CptGSx2gZ9T
B9/7dunzDO1L3r5wups1cfaohtXf2Rs165fQ7bzfw/mJsDIzkCAq7nZXumBsdEKd
twU6tH+nWooLM8LyIm83nW5f2hx98qytpHSNVzT00Zknpvq2QLdk0VdOeh6V8WRn
wz7QJfsk1O7kLbqaIlpjD5RwDpquTD5uPw2FgC7s2pYq5Xm+/nCG4/1W77ZyorbK
v1E/2cf1AX1uadaRGwUInnB9NEFPHpEwsGXQ64P4VpOWgcP6BSLBzLyAnaR2LSOC
O3PtWA4n+KuuLwlxi+qShkpzHRzAs1sXothoXarB7nF7Gy4XSQwh89WW9OrPcKXt
O4pCoSuxbAnmEyDO+Xv/WHtTHGn0pbKab9r3mWE4+35et7AU/ndcbU8V/CDAfZr7
JxQYg57N7le1BgAIzFcVqN32h22YwCbd2FBovqc02KZWhZeaphEfJXGB2QlCMRBU
+2oxR0QNo9Z7vO5hHuuB9x82C9kTXOA7t+ZHGnza54LmOx9qml760xCJuwo51McD
RciLn/3V1ziR6FfO8xaN5zZv7wwlWKm1PtZj0k6PbHY=
`protect END_PROTECTED
