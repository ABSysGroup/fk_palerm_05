`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y28e+Nv15z3WuUXzM1ztOgSgIowoPL39wP5zy71Obu+UkRVPO2WjYw7hgbB8PdwL
ao6IXT6n57MpO6R0WdGKUK/6K35wfsXz+JEgX9EtpABfcSfiLR+E5O2pfDaT/AlO
Bq14G87ajUaqrtxzNZCLMN4kEvDZ5KsST+QVI6KfSF70S/SzZxQmACjxCpdxjrzp
RWEyBYEt+l9srQFtm4rx1oTqBbYDSW80xYUlHq9zfQzvcUT3ptEDhb9zj3Eg8zC8
ZaqphiKNvxGyPSxIQd/wwM8urJo5euf6L7yy4OqgbSHt4C5hJBbSFwCxc5TTjaZn
hZjtk7ncZqiqS68JOpvfakpnQ57ozUJkanRLejHb/oW0fYQ1KZALm9Qh/T/YohSq
1RCwRiUxArgBxBxQRIwWEZRovcUpoDhss5nXt+Q2qhjdeUJ3yTUJwKJsbvIbiy+J
vK/orE88QBYJQKxtlBuEW7vToymMGGiXYeGTNd4sQRL2ymuljOHJ0qWkfXAH/ycl
9VL/iKT+Fk2z64LVGGFiZdI1UtVlEcSF3tSa2ILBtpP40v48RElJnqtVIZcCkwuy
/7+lJ+3pe1ZrnfKSb4Brj5QWqQvEbtD2+gdSUIqnPXgDzfxsRjJBidOzdh3LZ9mo
ZPuu3J9o5aGnnvk9eXgw2uBBRKVw6HFY4uWL8Fi+qt74hzpvqc7xob/pLndsUZGa
lEDm62GDnbJvN20YJkYpn8uVjoa702PLjvNNCd2JpzmXJrA+/H2x1ALRN8PZ4yoO
PHYxiSC3ekt83HtUmfEaZ7JZpqbiQn+ySV8Cbny1tZfERltrOmPgQ6cBaYFm4K/P
TLaK8wefkQVraAtpGSGNZHPddw0voZrizz7pHgpmVMUkGG8k/9xbrbVxOwFgVm6d
9ggMAoDboW/16dzDq1jMPLRXQGQMmS0CW51gkAI6vC5RbMCMVq2YbLEtQXOVLTpQ
SSIgJjATt03AbZQOiv3LP8yNgvuMZY5WS+I89Bq0xRg=
`protect END_PROTECTED
