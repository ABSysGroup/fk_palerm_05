`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DlQcqxS1chf7Wkj8dLDxsePpF1b0x8p5OMGmHH0lp0EHeEIEy75RxcK8bhNfoK9c
FMt9GK52lsJRNx9wMX3mWB1GGaehQPay2Z5rOJMiAdRhh26wSZl0RxF4P90VPmnX
Siyd3tvxPLnW5Qqp6/P5Qar74ptEkmpzpHLiCAVmCzvzKn8J/gZXs0998zYm5WD5
Vfm9Wv/1VTk4szyyACaC8HXYokn7p7tdzZB/E6vYAkqw1c7PUEr/WjNTELZSoiB/
0CQatKDYzznTUKA+j5B4ju71qJC0SeZaGuxBzl9invgj2EnDcTUFgLaDpvtbIqOv
pWfLbUXV0/ZjH9pHsg9tAlVG0Ih9TccFehINve5bmOh9JsfExr1vjpXVQAliaWPZ
tcMsQ8j4SQ3neSGq9IAky+1OFR+V1EP6SlPsj7QEJsuMNr2ii/CLLj3MNOEkea+m
X+4MRSnTudJtSekZ52jVOCqiyVgAeslQofmmIAm4pVkeFYf0BD04k+iY2nSITshX
S19UXil7nat7Rz7Z5wFs9zeas0lm4/z5FOaV/X7vzAlpPKa6emBWKJYAlt/nAaRR
uGnDUT/RP+zLbj+dopq/EU/KNtty6k4JGIRonT+cRgF+hid4+yTWxYhqRIQSl31/
NySVuYXTyVkd0/pssvhSgC3EZmgxjn8cPqXrEPlnBZpSgL22pue0/S2PoVsYq9gs
S+T4zVyCw7SDEB5Da5JkNvWAT3aAESX0gA2ITZxCkMviJRBZXwsNJ4YCR5iE2Pic
`protect END_PROTECTED
