`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U7kklA6AVTqbF1UjL0xGihqGOYTbEFt5GjgML4BbGD+nfAO7mcy+eYL2nLE01Ma5
/zLlKY5eSrmvFSjLT+0kOMDWD/nnfskj9Tuchjlj4aXVFqbm32XcXsDfRjf+AFZu
GSCdi69GIu15YgIU3Ui9XPPxbfG8/4QpNufDxW+x8btTDvWQBqdYp6ECpMYZxb35
Fvcs5XI2NathBSe8LjRf3nFoj2p784wVS8dHv/nakwjHp7YMLG8CaMKVz8UBUfTp
`protect END_PROTECTED
