`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E38m9ztj6sMrR/ers/5i+OV48oru+1s7pIxtARvRsJG9WL65NGefjgAM5V6t3DWu
Ll2uxm6MWdD1yVBFeCg9efkik01mNRe+EX1Wxex+w4po5Kv2nHG9K25xOS6TigRl
yQOC0t7v3ILi6391DGuMK6QkVxTGr+0u8hE4myfnOynJfiPeQfFKmWCMRZNcIV5G
/J2zfGSf0Kie8CMDMMa6ztjzVy6OE5IFxRoc4s4tFPmNvx/H1NDwthJ7m/ietHcd
VHPQ1pYTS+3+qdLAsT4fkCSHQrupKsw+xhKQF5RfATAZuCTF5wjFrIultnReG5pP
yQ2jZobfBQcdB6kufDEbWviTq3Hfte20wUV1JaDqhnu6u7Tr0Qmu7N6knVB5uAcg
w4DksRmufsF5xA8qS+0LEsMrePsCOIs/hvzKhXqCI+a0dYRrgfOgbRRSkMmpXg4+
zo4HkJ+ofciXWDz1PYpYgIzMmbMp+t59PWKJl2XXvBnp2QBsHGtzXj7wXh1C+H5Y
u9uvhD+XF/kQ44WIGdudM++YYkEBqq8dGjUDJA/aiibU8JYf0E+MS7NbzThDBKlZ
Al4FGdvN+dg8MRYbejLDTMyu6i2mtJ3EHFuqrpel/zUqjVXUDywUrHcmGTzrpbUk
Q6ZzzrEsLrpepZ+dw5OCs4BSHhutTu+xEC46NN5rmdM1/FfHjdm2wmSYOlUETb5a
4F4DJx1RQPmb/qWjjCRGPYro6eEwrxfaLSdNtT+j6d1vO8svLUix05MtzmoBq28A
/BGa/WYEqoUrMklTR+1TGyRlOfq5wuIXgscanMFHCkQwP0Q/mUf1GwZvzRUzmU1C
ovM/tgJjdwatYC8lGPDGY3CFEUSwQjU3QSpFgDZGVS6nKNSmeul5IYYKHmn2Pcne
XrTr6o2dC0Lan8zvpwqGWw11xIpiHf9huaJK8Qic1GED4qsfnCMwTa19Wdm1E9GM
r0ukCeUk/eCaES7mBeu5P6K0B19IF+cO8NNu+9jIVHSYkuzNGDVpQCpPHjRLZzot
yAEowKTnobbylHKqq5zlXJJUVta6rqrX145iOrXO38BO3ESbrHASoX9Pc8hONOoq
D5ObYqXvZvISl0j4gNfFNh7xfIKg0P0F8VkOlGrvDj5YKX4n0C2tcivTFnt39M6+
+SlZzkCbbasoh03+Uq/xZ6YJLdrmpVEXao1D+L3yEwP9xQ5VCaGF4zTZMFxHzVWb
PJ9a61FQ3WgkT984lDKFi4MK3JQbhH+xzGsb5//r4vcrEdRiOuu6ruVGVom48VzC
0t6QdEb5iy1+4oBLZLH5tbOC15+kfuiSdFdLru4OjfqITzlozU3kDWOtkeObnRYH
KUQY3ui9UKiacsf6OyxLKU090FaHYbn2P76vKSTyxNhHLXNkfEEFq1lXIH5AkVzE
Cnpg+VJqrxpRWBGkslxAn0yj7l0EH/yjNkn9fFI6HwOCUwu5vjiq1ETkGrw5zAY3
/T/1tgBQpI+B45dtuIJHF+MmSm6MYkylzjYRZQFS2TSgB+rr3+tZp3z92Tv3k4mB
N/WvcaCUmf3ptb2CCwf2qMSkZw52ls12rog53dYKELVJfzMf67HgFLhhjw8xKsxe
lxDlcrzUkh30ExNKXRhhD+QdQXdSmiCH25gGaIQAt3fobre/ZIISYwyz804wZVxH
`protect END_PROTECTED
