`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oBLXWWw8QGeXoVexjs+9waMWyKXK2Kz9hH4TPx3Uulny3YNP0K+4GzinZFZUH6k7
CjoERE3lXXwLgLlTwOtmgjGS/2TkgD9bJKaJ0hFWM9dB0pTDfAKq/6ZG68LUR/QS
AxhV56f9SZ3qyOWvUYSp1CxGjWFShCaVXyWvZ2ccSo3mJVahD7G/mgi4bf6uCyCq
SGN+HJE548UW3tNOKRKLHYj4jzsy3qfwbZosb0li0oynh9zIqWVsGdaUdgT9n66o
MS6yYtvvsHZgnNLWdfsqNlJToMEt0IPWco42YFVhEqkl3Z/ME/3yNjMuOKh/WLxC
jtAdoNM2BMs+GHtZMD1htbCQP348RnZeONMGb6oyUEuQAZrYY+xew/6q3EyUO9t9
hkDrQ7SQJL5CGfGpqJUq5OQLQzHr9NERj8cs4zvLFWH7w0sTmQC3mODeDNIilmEK
`protect END_PROTECTED
