`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PJGpN2staF5GsqTvJV81D7xaI3B0AU0vzadpWMmYu09ajmQFrSZlaqdxkzKzukDc
cEOSUioJ+gx7I0cnhcQH8xkZSrQaZvUzPO53LMk9hqekhcINGQ2Kg66LU8sPfNVB
YCdGNhv4XKlkD7NeOh+t7sUUTlKoXMZrqoKZPtpkQHOOt3QkGViVWwsYYPo8VOQX
+WV+oFBtVeRLOWyg+O9qAh+dhVv9ubK5EpsA8ilzIJLbWL/oEAxzdanTVn0dnwic
y9arDgW5A6FTX5klG1O2lSUf+494sY0eTRpPTaOjtepep22f1bgN1RJhTbjD8tJT
fZts+9On0J6bN0BpgxBHewXrwrWyuGEgmjfD7uQ2OH4zkqqCeR2yZa6ukB7xJgpn
quvYgsbUzgTTgZd9Bvulst7O/8A7z7bJ+xJuY3WBO74dp7RCHNx9Vrsqo2I1Madh
maVwZBCzyjtaodl1ySq4faxRunU5/4Oqp7EtuIlUlQPEEC/LoTuSOgRtqX8qlAFf
MQQOWPPTUnKpi9FqVLnc72OR4m5TKYutLDo7UuWcFK/WiLfwh5jdsvsdZz/Z6va9
1JhpCDKlLgdBB8OeCHX0BvZdus+ZFqQodAVRPm4x7flUXv6al6cQS7Sayib8CwKh
jKC29y40naxZTXdQrMpWqfnXoka8zSropH2r+V031+NcCSWj5YDXcaHo2r/0KCaC
TXHmq6O4S/kp9bnmYqHWhDWDt9TDmtoTcw/P6f0fXBM8M8taF/bmv/fWIb38xzSu
VL4l1hARMkFBiFrUBibGwjSmFfTpkF5oUsVuM9YTBWvichrz60CuvJPEmhiD89qy
VDDGYLMv4MX9qMXA3GMKL9OJpbNBotCMQitGlFroC4hkequxU806fhh4pue1XkmW
6ZSSN2/wgnb0rGr0sPQtaH7SbI6/a/slc2IjE4IZ+Tojk2mCrse+W66qsnfM4ftA
FEE8GgWh+K811JL09/nN282IibKrAbEWwrQPNUAxlo+7kBfZYuse/+9W78rA80zy
fH7b8YpDqdygsMrE2oCzsBbuHLSUf480g0lppsBgYqUXf7NpmUkg52isjJdiMZKY
jqruv2zIWW5zRYMIClEsXNnLnhaCkUGjuXZduOenFQSw3UIhc00/pZcRcCdzr7lU
DtInbBgFW8lKfBCw1O+U0z4o0fNpQK0FkGvR1Qm+qQSNYTtwcWEQoFcYxULV6QUf
65lCi2lT/FRhPQMrjoW0A3RIkuSh6BWi8WufKYqfrsHNFTszzIem1Em7EjXXme+x
DOzpF+yWx95BjV1a6PCvK1bqEI0lLGrHWmzGqekF8H8Y0pnxAAurkPow5Egu4/hh
rcGZ9Y/Gb5m1ycGb/DeB1R8WQXGPc84Kk5dDJyFJ5c71lGQMaknDXDvaX5GgLOOK
qjydTLdw6Iorg26sivMso6sxE5KY1W1N6fD9xu9FYed36sJH83gGeZmCa0PnODJD
MRBTx9ULyhYWw7Mg+/qfvH3PW5ADIHjDTBtbwFipjsk8mhmfYZDqC8eTNFHuMQuy
GMjCkGmUqgYfMC5kt3N3yQcbS4YqDkg0aa+amsfIhiJa1FseBbR0tRYkLGs+VL4a
v+kJcTaU+css3fKiyx8vabQ/GyfBxeYIpYFWCi6DQnlkp/6ZfCrH5kT9wxevM1VI
7UlSuk0zg1z8TGsHVoEmFEpFGTeGZwlNtpNNowjqfugyVwiCtoTloJt+XJd/FHfY
1D7bbz7Rve70j/52VemjJ1DL1vmvxXqpV9fTv3Lp385EZSj9AL1wP4rm9ZPiq7iR
Ip+ri6GVu2Wynvc1S3JO94VEWRA6uNmviMXPeDuj7FAGtr4ptnxYmEWkZWR7Aj5L
ZZ0QYVFyf/3SzGWWpNNcNAD+xf02CD1zH8pFQfcds07fugVZ2NJkq02U26CrAYHx
gvEemzAbUtXU7mEGbHS4XelHi0ow/3O2c4fKeKlqAB8FDJ6cKk/6Tyhg34zd838n
ByROG7lH5dQEUWJNz5O6FfSBIwU9xQOJC3LnonLgAdcmChKT8yPsEQ1DaZ42npgo
7z95OZe1jfGgCoT8yKHqlvUi39C7bKPqAm2TkgnxqYch+oxy0cY1160eP/aeIpQz
hB7u810+nBn9MFZy//JtNdZY3ES6dXf/Q4Bxr7As6GozE/8SPy23UqW5s1IYN7JJ
DRCOaw8LXbkfgtEVg8tfs/kdh+mpcj4xfb2JUnm3I0jpdwVK36/JOk+AtKp/2bml
aEMNm6OhmrFxUWKp8znwZa5R/ZoEPk43jMvh+IlnJcofa7avA2u8vets9zPxrK/A
65iP9Fuxo1KK+1nBFNPj4GpWsdzOkjY1NZc+ORz4PqDLdLP+EL6NPocZZw5jDw36
jaOnua05vfn0JATl2k0Vyzx7oi7K9LRYin5WkiBUtSpBIWFeCXXZlZFZArsVxgE+
Msd9csH+KnbV5KOGXBmYqnpzEh1gfsF4/a/+zElAiZrEqTuOvkIJ2VjDZaDrLHkp
fzvzt1510AJ0hMEopOuLnoerECeBoumOd+0Gr+WrC8Lp3ln47QgRQQN6GNQ3R9zw
i6WPWVNvtxb5/njA4yRAWhzYS7bwDlKh3bm37i0QIh83AL9nV7UwYgk1jRlQwv9Q
I8pxBFCgAPWvlUqFNfduOMpDDjRL8fjuRdbIEwbvZpaKPzwHA03h9yEyZTAMvIc+
9QkmSoaGfa9y97a1RcS9sGwsnetP7xvLFMdWdQVU/Wh+iFrett+tfblyMuUDTFiP
iTJ3CRe1WMbmtA0UAmfXOdtQ705/5Dj+ic5+tmXvv4INFhFcQZiz7fbqwTu22CRr
OfRVqq8/OLnmX6MXFCFXNKid8rWB/yyBWNnmDkYqW6DdXQM7cmKabhGRgaFL5tTR
BEuoWlncnwqYKy1W8Yve5spqJY7gnlk0vukvDFZNdOjsEYPkXX0P0VPvM1nWK9gS
kXVbFpB4Jcfe/8a1K6VIjIJKjORnGR9kcMXaw7DUghgr16oKRHEgvcahS1wdxMEY
eLZ8q2CDI5XewJydebaehk2atUvx3nql4phDgO56r24RGS0kKdx4SC6Q/ioKx/Qb
F6yrqTdHEBHP20ffBZDCm70KJdJIpaE6zmO6tTLHE4+ji5F3vF3HicBOZEHJNH1r
Ppk/Rbu80EY76T7U0OwN/kV63mi71PSDtUZ5HCryTg2RftowWbTIe8D3gWLj4not
7X8cvrHctF80bYdlu0eVNB4pUrxHvuMdWrRouMh7SN/wL+d06lTt6IYwBZlJHl0i
bEH5zKy/qB0uLlNpELhz7t0SiQ0PWVN0WGuCxUlVBVzP30upYM0dMLIue3HjYZay
1qdc2A37RduLt8it7cCoCA==
`protect END_PROTECTED
