`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BjKAnYtk/krlUQFcFl6BNl/D2fQakpq3gYYC1EAPBtItKMNa2OLVN0JXKQfo0vfy
lu2Rp7s28RjD91lQDgjJtET01OO5TUwwR2oVLFuXoKQ9daDRibAY85zgVMNwG6dD
QJStje9geQn961eM46HtxXH6kWXDOYRubnpx0CWvhWVcuLl+77TvUDFSVrsZyCoV
risTRSJZLu7m+cTnGGLpPULAjksE3GVeyQYMh4E1YyztEdlbVQetX4W2f2/b9In4
Rma09lz63027KCGwRAS+Ig==
`protect END_PROTECTED
