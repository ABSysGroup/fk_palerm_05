`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5GwKnUR4elAMb2FSFf44fKkTgAyZhIXQcDKDqnGJ75TpyC0XInsitqNH8ZVq+n6L
A91xLrRfIEQXspylQr2x37NC2MwrlfEWqpLSbszlK8jyTvW87vxeoldC6zLC1UsS
ROORm1x6pP7r7zRzrbhD1MK7wtyek8uaf9Iyc/oypzb9FTbsH9kBKb4ap2tqn3sc
mE5tMipxkzHA5Qlq3sTKwvupWt4LIgjmuCZe8jDPKiMyQMBJ3UctjjOrH+nea81Q
Y4wD5qZ6w4Vww614O0yoTI10hMYFP059JCnvCMSlGES8CW988P/gVzboQJeVMJHs
nIo7UJSpYCyJ+FuLyywgx25hXdTvlX34vHFe1lUBITwiA0PJq8O6Ued8CSC1FFUu
mMzdA3pxJ/Mkekkxdq6VbjNWw1TzMOF5hPOtRCNK7PXTTMTD8LIUq7QMMAnK1BDM
+dQOLvgavNHcGVQKah2ueMEamCsAih6lQ88FX0r5aLBgP2OdzYxNnqsrN1XWxj+3
D4s81sm05/HiRx11yyS7lhguqWWArpgn5HqhSVJm+qnPzLL1StiD8e0X3XG3Io7/
/8wnGGv4pN0uifgZLtzF+8Xgh947MNWYs5vVy3Hz4TMbgBi4m5p/1YxviOcjFmoU
YGFw2r7Ujo39EaU3lw08v7UxaZ488oxE/+u9I7LpYpT2YUKLbGyebVIbE4OVJP5o
`protect END_PROTECTED
