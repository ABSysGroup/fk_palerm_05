`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
09k+O8nKoz116MH8sOQmZV48aW7wF5dwF8gmJjRJZyhTqvPS8n67FF87la9bnuGe
FY0rJsXY1eMgeZu+lgY6R1t/AoaSkmisG7BcmTdRmnnnJdtO1t6p6eLKB+7XxdXi
OfM3Tt6cRAQ8QpbXVRwPBdyMV48sXIYaVpI3I/IknvkHz3y8RuJZ4plNGYwYWqNI
jCG6DEbAEaWkeBprDOVwNDei7xjTMA0+9Eaw41/SjlWYRxET8eBmzCU5n2jJg3Wg
Jehpn5QrTJm3o2wBuKPSV0JX2i5OjjWt6CpAWIk72Dq2ywaD7QYVEyRKzw4u8wNC
mcfIPCAQGzpKAgHSPFZ2FG1S26XE1h8EeZ+k8TIWYVKv/IlOMcBARzaaKAuGJFEu
k136uMM38gMKgGs0J6TFdjiOXiwrfzZvtgx+x75WSgcb2VndrCxUm+eHUoJ0fSr6
K27SB5HDe0tpcpqYPb/VtWeaXAJziYTJbH/JSliBIYpditGMpVVxUHlrB/8S/XW1
RBB+IuSiO42klhFN+EkPnKybXU6zTilLOmQ6xA48dDvdsqEqQVkIdV+I95LPWFxN
7K48mH2zMVO6aJeJW92hH9oJq9fgYuUaSq0BiheBN0vmkfffUIrHVv9D5pZkjR0J
QwK+Bfk/3cPoRz4olFFQMYIfGzvlc9IOCdU8DjdYPWraEE5NOHP7SjcwyVBRmObS
SpU2wT2hoa/gUTfLzspUuEH8DKzth9d73UUCLqVL1RjMOkv6C7/p3XnfOUzdkYtb
tEUCBvfQvEkl0Od5t9QrijTWGZ32y1P3hOiEiYnQsDSdlvS7E+B6Lq7T9wNEic1z
gT1sydx1M/bw4kSkO2o/py6oJX2sHnON/NxBS7EemkSYbRpiIJqagvGJiCaxOtRP
oEOD88jFAVBTbEeW4gqgtA==
`protect END_PROTECTED
