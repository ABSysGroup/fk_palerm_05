`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rxl0QxsYrUoKIzmkYLFqrAL2jkWDNE8hYgFFcrc6LVzXuoIfcRp4XweLw4tMvFkU
j6y7TJtC18PS+YSqwitfaRJQPvXIE63p5nQjAQTMVEv1R8gTZxkc8KFRGWgLjy37
TvxK6RjUsLSfXFKkhYGSoaFuVjTcHq0ZhC+qvVTNc//Kj/woKjaQK84rJSORI+/u
LTQgezwRayHLz4/+GE5kdUQIj+olLhTK4XfHJy9cjChk23esv08L5+R0W4zP12xn
6m3sEzUYv0BgHX9m5D1LwFOHkylzRptvCngfejtf2e2OKa/Qnsy0ZY5dIwriVPiQ
cCcrD10r7ErLqkx72i8hGvK3qv/LnMGzcv/CTTyZL/ODztQ87jnQXCWB4n3FGXCG
yjdbTF7m37/zyx4k4J4TynkoFT0gtekqI31ywb15V/KNjBwwI6abgnKYRYx2xnO2
elnvV8AnnDGtgWyfINJyzFcJneotB371keXd7GC8Q3G6ZUiRdQr2rF417zeX34ZX
4OwyHuFwvipAmrConIhBMsPWCqJ1uSEiVD2pEs/tFMnDA/e3aqtZkOeiTiT2m7Xx
Ew4F8DEkVli28MmWQjAMKQ==
`protect END_PROTECTED
