`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iyYisxgvuHfGIye2O26EObXYt3Z91Sya5JGsxprlYNTYVfNjIFrxE+QkKu7KYzZ9
nnoIehzOd2uwgnNOdHgMiXbrhDoTcZ1ohDJSOvKHkVzATFrQrq5x2vvX7Ls80/Vx
tEXaWIm6ZTaumQovftbctKYuAY9bl9Af7skasn4by7E+j3gHzKI8fIWTP6l9BerM
2a5yi44J+OTVPOOa2KyiuhT8MvBB9EHOHWV8hX1nJ3stFe843BeIydJ+BCpIz+Du
ML5FfUkSn08jJZR2snY8kZE3gF633VBULb5cKNnZaLV6zPCUYZysOJoLo/2LMHVD
R+JzcVPKmfCl4a7Wa2C4lZFbaMz6FT6OHl/qL2rZJzlW4PO2QVgtdOfgn3sKmr8O
9ZEOfdOwvmAT/Thgv/cYURPyiVQ0JS8bB/xypPRN9eiYL3q8f1giGu1c10m+Ton7
LzR6mUFD32Th+BWDectzgZhqkqNvfiuT4bKstnpL2a3Mg/Anc5DbxLb7fxYG2esQ
jj3o8C2GOhhZUdmcfZIRlaBmQSoXF42xTItkaahPDzW7RU6Fzs2ItDGIJU0A9mDs
Xznet9Z3gljDVqySPsi5BpBuKRnkgpaAxCE6cxiB8KrkV2xCvzIPjebRW7rBwO1i
4mTSlfYNx6Pa4rsu+Mk6Cob/7ke6+7Y0VA6E8AmQaMQ=
`protect END_PROTECTED
