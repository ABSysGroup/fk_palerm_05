`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dHaLVOcNGByjM12hx5kbuz+WxAz4k8lzt6BXFeplzE1W8VilBh8mv2ALsE3ZOqNZ
kDIzDq52ZseWFNVHTB8WmClVHqZeGrvcqJbIlndxQF9Yzn5DjqWxqbhQ7wQjVBJY
18bq+ydKtaIKaMNIU0rqutu6TbFeTNi2mNGF0JL7PWCEgSzZJRAMtxR8p8mQlmWm
q2d8rYCwU6jQ2HyHMMSuB/ZSRrXodsNLuZAWCNwIIuzldntZP1dIYBfzWtUt8Pq5
Ws78dIEQ22Fg5/LMjWfffqW8+Z2HuoyVOuPxhKTSVPCPNW5jcbs+cHmfSJELLHfN
3Huaqv5RxH0APWZcm/imKE2U6GIJ5Cb0GF3WCwTEdlIKqQqzIlwnDCUrxTi5Q+a8
TCqSaVPpQyP39EHTc+aHYTxvQ7g6yBrw+m0xS0CuIvmGDkDLQjPDOPVD7MUKUMLu
iZLnZMjVc6h9aDH10SxDmdGTDNAB2zEkPNvc009SRopBFeHO6/6ngoKM80Ip39F8
JlIKfTxmRHNDhogCWVvJ60kJwlt6ZjyTtqarP+lc1+gBshebj60ixi44BlC+s/8N
RFLZH4hgMiuG8VieRW4pEDzQwcMmxzgRyXUNmfGDP4su+fF2F/L+A1nNQQGoioi5
0WrqAc2KdNbM0KFgyGu2gtI2D6XyAjnjlD+f96PJYolkm7cLaloaJhK5ayeakoX1
l3CB1eMn+OBDHO9Z/K4ULHdo8JWRSyu0OsTuHZ/8uAR8Ysq2S/nvHRefttDoKC+D
glo5LjFU7sUPApkhocm5mRH6QFkqPlQV4U5wIHWqpBEB+6Lhoa664PrKS6JwoBnz
mf78oHX45VRRSFqgNg4ShxhW4k33rntD6r/kOH0Xnp9wk+j/ms2Nb0IqOcmeF9f7
pWfMFyEfktzxdHudiVoJzfcCBS1NmGkXnjHVrlDWpOJ2DSIBFQ7JnGP/LAnqjnud
mnOlGQrgqya+r0qw8oxxPZ9LcxdBcB/1Z8C4XwXgBGO3RigWll4CR0aF/f6njbj+
cBxKgtNWd91uVpWUZD4mKnT0AA+08YJeXuRMRehoz6jAqWEI9x/F8SuWKnrPvCKE
4dUFD6PHt6Uy53/rKq7MmIi3aiJXo6fCKm777IBGDtqnYxwR+inx5wKHfvCp3rr2
+FUTvUAg5mGd81QhJln+rsLpjLU2E16LxYRumPSmmPyAtPjQmhkPlYd6u09XVJZL
h6sVAqjijaA1gy4YdbHBLBgCGHV6nthuYKoRtQ52alU=
`protect END_PROTECTED
