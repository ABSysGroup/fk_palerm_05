`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5LaOjJgGKrIlmgqSG03Kz1RRYdb5XsI+yMp/DoDGE/YFlK+AnwE15umgeQE0Z4Re
WVL71Q6/CYc9eJ3D6l6yRUs5RNmnbdF514B6VvvzG9ZunOGqwhA+1ZZiS765rXtL
pHsr5iHukYG9zWM13x5fWIetgwvWMr0Uck+TSblZWzbVCp5+f0yg6dZT17uf5ZPA
+CW062bq+E9j1pwCy5HTOuzwo/Oxilgxy1BwhWio/CTFm0XvL6rYsO06x/i4GFB1
OlbmY7xfgx/rgaOUDYwnMQ==
`protect END_PROTECTED
