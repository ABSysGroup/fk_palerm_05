`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1DS/N/+20LquvsmwgyJtIg2YQJCY3gC1DYvJgfm2XoQXmPhMsV/3vvJ6B0Oo/J0M
Wio7356UFp1nSBXIHAaQVyxUIEoPaYPAuHcbmYiksoNSOIpTc8TLEX54BNmaMP7b
PQkFcV9WpUyPuaPKOjTY2nIJtqEy9Lb1CH+NBH6eJAaXM+wi5DjuW2vfHtwafmuS
pcZAIjWOn12+ilpIzAE0LD+ZglC/TFsNReFEkkX1j51DSxIWNfdCyMtJrAa2zMqn
mggIpOEBKp+FJrHrY4qjRg==
`protect END_PROTECTED
