`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
feewE89pF0dMnOio/12eVSypypf1DSMUS4G054mJMEJuDzq97oNzlOf77YsfbL/G
5A/JzjWnbObRcmEMMYVP6nUOSrlpNbf57sTumOQUBvg3IzYN8OYl1Atqd3geRCTQ
wyr1CaHLhILA8T6IgoQfGZjst99cbpIcxajH0Fn2g+PSba44rk9lV8e47ah8u4XY
sF5war2k8KhbAtuLBg2ghS0WMNkBLIIYjns4PNyajyLVgHmh+ZkAqi3EyN4sNfDE
lPXRfQIo/IDpPM3GHGNgCwu5IiuivmoY/mmykWra9YuO09jgDtJ3NA8z7qhXgo10
Mgnn+7vc2xni5eiuIAfcFGcljIhk3yxL9e7tgagsf9zP1Zy0MtyuK3qBTlLeW4Ft
CBR7UIlF/8NrsP4IWMasG1gbWgM3gsy3XqJV0YwBbd6layNZPkueSD4MxWjvpe0g
dZTbvD3kBDc9ubQvCF4YSvQ+LZydvF0E+Pnu9Nrub7f1/TCAy2lPpjCIi0OTlfY9
ji0nyhFzOtCANXLcf4N1AgzO3c3g/IEc9E2lEm31uU24FNb8sTpQ7mhFmnTow9QC
tFOnLllzRHytllh4ORXgp38wDfcBK4IRSD9QqFekbn2Q7NEiLo2ODjHLlLcxJ86a
7Nr5OqifKJ4NmIYplLaXymT1Qyjc4+LLdbYEwF22J4f60nCwvXEvHxHrAcxzi0DS
AAiQjdcJh46pP36iOKNbfXUAgizkmQOc520Xs1NI3PevDkVEMieJZhbRtEoguSfo
TBXsyz8kPkGWRRQJhjAHFTiIbsnDg/rs45UbJUAYZF3tg3tfKFm86bGdJVd4Igm/
aHeMhNsC+euogxxo5QTiB2zYxZackiOuojDDiCQuscYlIxUUOQqIz2q4EBPU1Wf1
MZfxMnsX42PnzCkrzqaO1h9giNEO1G50BXVKVcIbosj9l5x+nBuAnVK57cxjkkLI
5REQPeOObyJ77i0bz0pabYdPXQm6N3uAn2OT9YgGcV+9nQ+6qkMyfGIN/YghBciZ
HY0Y1QUwPEq3cD8R/7MW57eJB5VpSF7DYNigeDGziqCjR9+Ks/l8NT1Ms4bk8+sA
8zxGNsIQN8GC5veup2DGpImEzkuRSTTwxyrc2q40Q/hP+FieqwQNIbwusnJg4Mzu
4ngo4b/K/1ybSv3SRMe+1WN1lmTpQhS3W2TirA2ZSlYbYVKNOm3caOksxYM4saPM
FyE0uINRs9C8UD8tK2DmUJB5W2f1u4PJgCkWu7Ih0ybOBs7XdKESJ9LRlcyOHxgF
GG7c0AiAtpVgGodJ6sCSANH73i7VEGFgXWZ+cQRcKxk98oXV8Zfc9FXlrlqpIl6n
EH4M7oYpy/to0WLsQKYWFru12PuP8T0kmeijEFKGA7IcTh3ozrq1IIhe72zOpdok
tq9sxNw9QLYEJaxG5+SnU0A6Pvpfxs72K+OxVMszbQwnhoVpSEuuBaKo54PV6lnT
RKp6KF+yCap1SLhM8Kev91VpOvWsS9cRb9TtjC8ebQN18/8oYQBFY7yxi1hXX6AE
Up0VexuTGOHB3iIeQ5NIIFUA/rLCGn7EqqX2v5TZeZNlNtuKqPx01WOd7hjklXCa
wf/pzamend8j4Owgr3igjKKN+8sSe1XVgw2k8M7UzCZc/UOfo9CdM3PZFf3ZvAX9
lSqF7TgRmcqeapc5wK/bG74oc8FUPZ3ZbdRftf+NCtcgzlrPxycxauxVzy3ou1fi
K50J8O+oywZHo1HigkU8sFaVw+aqFGOigcQrThxV0bzbI+hihBe3LCKMrecH/fKe
ByMeudns6sPxc0vlqPbmNkKy3SNVUQKwezToYG9r7PI0sZoMPGCT2/Ww85JWIr41
xSGlMY3sLKBsOXLCs8JQEHCRz5lydI+VpUF/VeDgxKhDNLizRF9sTBXnUq1rLMJI
Q3cSXrBV6BcM4daQZBZVLWYIlD9iRR83oirdMO7RsJ3/Rrhkvd3FAXMGXP4emKIG
Y0CAtBbFXZr/SYsOTfxm9wvVcZj7mNaROPvqin1WpwntqujBq4WWbn7hBZCOp0sl
GD83ry4FW3JSzChtZrrdGw==
`protect END_PROTECTED
