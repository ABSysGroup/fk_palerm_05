`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nymnjq8UkNwQjwUAUGE0iKk9e5D5n1FyHC7y1qLTRAOpzdll5j4Sx8GKvg4B/SLb
nfCsVWXdyGnbwuJktRnnHE7FI2B81IH9TBXCpWEpXcDeGKydeau1my+okIk1Hda9
fp3HMFxgHSC9ghfhRQ/fONQunKwQoXXiPBHYxyUMdyP3mqLBgV1GVEmxbj38ija3
jGNo1WzGyjg+UL/duehHFx4g5QMyyb/FY/Nvjkrn3+6J4RRlH0Z2uc6wC2T9lEG4
sPo/iprGdqiSJ4bRwIu6Tl6oCwP1RIKe73dboYX94evsNcKMCip32PuL+MSTVmJU
dQ5/0cyOxv337DJgtdx1ew==
`protect END_PROTECTED
