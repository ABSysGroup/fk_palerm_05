`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dFb6uCjkP6nUuKlv3tZkvJMC5geUsQAoTAjVQi2NNmkTGsNGr+SsxVf/SJ1u4CLT
ztiRZuPSUHwnIU5vSY57aoDzS9eTjkTHB/ESK//fE8l8HDqXdr85yxp+0MJk8JSx
YFBTyBKI3cuv7gNpdOc37eNx5exFav9oXjwCKFzrRfm8yjtFCQ3Qh9Hbsi97t8Ei
jjQS2y596RInsYWECHPjHneV/iP0dYpsNRLfnozG3lfJVBcO0Ggoi8dWfzavQPjF
es7Yp7lkccE+KdJ+nYNoiDnW3raPrH+5TuO4CocFYjRCMTAAd95Afzim4DOpxIJF
xD02oO1rM1yxnGQFuMTM8TVU/PG96v+5p6fBY+cCkJmIq+DCeQLMViz6LVnxXm43
rOYvUeC+juBqz41oDyFrhCP1/62hVx4E+bXQG/eRRkvSmWid1K9SY4Ju2hs4+/jY
qsTq5Oezn3dejbFXK9u35FN/UbEqqEIQ0FYATSqdiUWsK9L8g8UI6/RPfPZ1v8HU
itd5UoUpqOK1xOaA1xQc9ugQIxxYzQe5rEaIztEuLSz0RZKvr41BIEvByjHOGAZA
aSNRfa8/np7nZkmGPgxRzmsLt1UDTP+vO2Ech1hs83TUTh8Ue7g76OETWbwKHLwK
+5SSU/0ogRiq7oqUN+37tbMqmSzXmaZ38P+IkJPts7U=
`protect END_PROTECTED
