`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mrAvP55eDfWiWSeO2LjZtSe9Zj98F+Jyh7Ry+s6TmZaKJwaF1nmFHyG7T38Ddj+7
m+EYB388AGsLDpV4wTsVh0lD+GjiwfuK7sWqUA4FBBIa7hI3rBn+QlXtq+/fuFKN
qynFAUjNJLsg8ds9yVTLksGd9gZxtbpAPvMzajbS3CUaAFW/NlJuQpuCF5IIazum
aVxRw866uwPOt8p2amVUHMpwvg1YBoH0m+1hKc+B3wWhmi/23+ER6FL1F5/XPMQK
/ktEU0s6IBJcXN8sAT9IOLWhVsqmPo+6mD/Dg/w3YIYvhHgjcTUNQjgSCdoQZPJv
H16bwsVcYEhPSARMubBpvn643Y/+Or1F7W+37dF7Usq1Rapv4JqcvoNPm3Q7zA/q
gh+KKeIwnJCQTyH1TzD0aEsJtXVMOPo6Eekle4XataD683YISSnGzuIUjnVaxJ8y
2CQ+Ji0+R67/bNDQ8Km8ANtGYnNc3k6ooDLQDjkL9h3XFcAtk1f57ofuRCh0kWdb
gqs5eefT62s93YECmJ5mMpqBCdoZOJZFXescFddPcsS8opOh+umr1p4Lu/krVp/1
a79dvHlzucCM6gUqE0snYV9TyhbNb0zYMGCZzYsk6nglCpz/WGSD6uD+ooPVr0SU
YhvPaRnOdBWX5m8Q0Vlnx6j2r2h30Gqykg6dlvCx2YxPxSSvjJeMiwPjl4vxKpkH
zstjcmBQj7tO8p/CUVAgCEFAc5BBvWns8/nY6gHs0cG29CX+UDKjErHp6H3V+Z/c
OX6jVMOrOxfQjrzmdD95fNscL5w+EU/HeAo3IXCRpqkSPVAMb6pLjUWPsxilbI10
8z/VzMwO1mtJPIShKYOzYiSqms/veouzFf9ubHVzrgBJLXt85esc6hXy/FhLJ6WS
a7I1vZ49pIIGBKq7keKhr2rjxT8+44AqhhXIM7GB72E/Eh38w4MaQH9C694Pg5wo
`protect END_PROTECTED
