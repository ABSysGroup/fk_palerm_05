`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H/0766UmiPPJXrKKYjn6VsIUeRdNxWFFnsvLW839fd48t7pSIFeMvEMPyrN8DGrP
Bd17ECaAQbifZE6fJqyHkwf/xxcYZjkP4GJ0G8/zfM8NR0lBR4YtW/hH4h52mof/
mVIT22HNqDBabqPnMHJrHRdnM2nLqqTfGPqBGzwquikKF4KGoAvmY8kEhNbjiF6H
F2qoHZdnl5IL497Nrr9WVSauk2DnQA9tHhckYAXZ+R+zyJ2kCq1BVCYnqwBcRUlj
`protect END_PROTECTED
