`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f4VPfhfRNGZ/bSd3BK8tpQnVfEw/v+GwS12/kVRCK53FPEPpkf3MCw31uA/lfdJr
pnV07Xx4KoTNZpgtMXydUEh5NhmGkdBG8eefuS+WfGj3mxAhhSLkIy8NeNF3Zt1i
hKNk+F6GdyWTza4M3bR0BC9vXS0KkkN2y3RdXTs52KSiGY+6LN2moHZGWa/CE37K
PkMREAG+w/fy/y0SDcDX5dnv6G3fWHorVHYFSPBQms2bJf4Q34U57UIo+jwOpzMp
K9zuP58VW7JlJPQy2VRbGw==
`protect END_PROTECTED
