`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JyoE/2YT3l0BRYMrVnOOcobocgVhTO7QismmEmgYXnH+H0HCWcRPRCxGwvRFyFHT
CNtjPnMrhoQ4Wcy403h+4lMqKBpLmpcaNnFKLwyT5kWkTFB21mMuBv2WAeACHVUa
/B27RTI49R4LxgYYXRZIYBr3mX8h/3HWHhiQi0MDwrwDtNxR/Zgv+GZThgI9/Q7H
0vge6pT2nIVMW9zhNQlnCyXD1OGgFcz7pwAcnkXpJy9Sp+ZFLyO7m81xdI5Qr61r
bx+BnT6IaEKxgpkBdr7rDpOXVa8xhK3YalxKqzxM9Ne+8a/tAFbeaKeANdGclA8D
Qo0rPLwnSIX6cOGo9f8lhZnQJEvgBaP9NgCqpAFFMwEUyUzSHJp1MtGWR4WPpxip
l/W7fRyDkP0Nv6DH8yauFJf46Dyps4jx4Zws8A54nMGzwj9xeCDZpRA4COWFTWjo
`protect END_PROTECTED
