`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ZGsBclNdAeZbYxwf5FIzGdw/GyyZmpTYhDs2vKa2/4fItnpbOEnCtN+I90wkb0p
RD4WPmnTwPUlW2GFJMobTZV2x8SQ+CqTur73abc6E35vTwO1bVMyWhwrw6fOeUTd
CGHExN7wTfUsvVNua1u7SAmyVmHafxOpffogD3jEK+PKtvHq7ADsduBMl91DXLqq
X9Kdy7v9lrRowECgwRQMm8u0opCTMV43Ryg6PPJTxpmB5SG800L12nKYnXrkZUTW
suv9xENe/VO4MMtI39AdgnI+zvROFq9XJxvkyljFEFDC8U7j8DXHfmmsYTF9axNQ
GplY1UC67AW6pfA4cCqkKC+8g5Mk8WAQr4ignurjQVrzr5UhltR+W0Bp9FS/qeXM
jsz61R4GakWVcdxOjJh/KjhC5sua3jC4+AOcfoOX35ncRH33aTx0HKqefvagK0Yk
F3/9T6rcmdA2LtVjf9idtgRPx072P+Es4THI/eY9gGT8cyM+BORPP1jGyPXuPQaw
luFoDlyzsBx/FnDqouNtRou9ihuIzr+22k7RySMYEUjaj7wWG7uFibz3uGbaG+zV
RUon5btGjVPdoXH/ZH21R+4jUqRGyB6nlmW55u4kd3xZ2Zfq2Ifr0PefgccYhFuA
FsIof/S6E+lig880m5B6fAzfB0ZEA4ihoW9VR9VrdcadDC3mH9SrIeo9DtyCCMnI
AtUxSxmxWCzOzJJ0GK6UhePp+6Ti8RBUVmRWrq1FE2zNdyWaiVtlpbRjCFXaBgF5
yEhHVCz70QCV4raGgVo20g1NZA7Q+X7FFiyx2QgVf5hApotEI4GCQQfuD+ks8gPX
5NJH9IfkEdpE2zDJcKzX+WMlVP7Y7imRRjRWR1y50QPuTX3Vz9XMV/TZHQkgPF5M
ogr8EnqYhTr0zBVUPKJ2eQLiQCjIyCIYLTCTEIOhIDQMjCP2F+xbEd6PNRxiA7jK
ACDl7eF4RJBLIL2O/XLghmcMh05xx/3qhFjqfj0bbzI2W7M/53cRL44HuGgRnfl+
SxHhW3PxStIJXWex+6GfbhQ6qW/zPrywQtPa7Cq8MhB0AQctaWwruJKQ0YyeYeAA
QgGqEy9q0TXz6J5UEMKbcxXLG366JTYwG5LlB5aYjCaCcljlnIqLA4M3ZDePxsX+
DOBFLZchRzHQtdpcwlKIXuw8PjCrHlBHGrDcpYEjsc3zdStoChR5zu/4kwQ6++Fu
r1cfLZzl0NuZ8sKsZAbckmjjVRLVGz6MUwWBoTVAL79bQJijob4LcYfUuvA3dlr/
jOgpA7p2MCMSvumxEYx8sMIIUjrQrnZ68r7gJSz/OdKoFUuTpN4opAqTWqbFuXfV
SbIreAFEoW25thRxjq9/ClLYZTBsLNkyhGScjdUHGXbBcfSfevFbci9PpQC2elqQ
ziHLwcQctWLPvpvRLmsylSuDwHctaXXdfPjw/WWxfqj3xVPdWTs+smgH0dp3NTW8
RMtN+1X9xkn08ziS4Etet/4lMZrsY1zeQsBZKmxgFiK9Hh39vlJwwIh6+4qdF9Gr
7OTrHQe3HcHYgLl5QHfz9dLCuj3iihhGpp+C7hjr17sSC6X14Yu8cbacHhNoLyu5
+ZvHdSMjoR8UKJgigmgORw8bZaE426NRR6By2zVBuiguS5hKm+9BABxIf0Vk0Lna
97hogfBVBURiPLD050Jl7iIxcU/XfMnzFJBqhxMgY+TEB23SL1YVOVuIdi/iRPuX
RPOu0ASDhJdt6exmum4LDiGd8d54uJFxB3Syl+EPlV0qX16v3351yXuBI9kCaTrj
++i7bHmBXUeI8XM7q786FHibU7TKEAWYdcTqu5Ov7IGHJpKXoyFsH9OiWiFfYVvu
sJb046SfJrFkc/OVcoC2E1KfjTkcqj5QcBgNnOlOdH7gmcnuT6bfEpqZ4qaTInNh
Ld91ZVolbJVsLD585b29Q6XnvgQBZBq/XxOsuhfZzCAFblG6HwYH6q6K400XqS3x
e4e4j9U6FvtU/5lXclplPylG0JHoLb7ST1s1NffexW/zKtx9fOTYfyS2oW8srU9K
+3vkypPoYwzE0Wo+ELPC+zAqcggc2yy1myFLMrHArx+oJgVRy7/L/1jzlQxbfcuL
44dqIJ5fz15OmZMp7ES0CjNAEdTWMp/rLoQH8TzCBvwfQyzLVVrOIfhc/QdgeEgt
xslyxzW/AdxhhNrySrWJ8pXNDP9u5uR+X10m1pXwQxPQQjY8vcnQOaHykCZtCOT4
DQE39KWSIl99L3F9KEMQZXyu781p4lI137IlDqK4Lp+xAIzeHzN5ATSchedmB7Md
M+FrGtlf//X8zEfNYI0l50yWdQ4guuv4qaiqi+G6CEYNT/pLp0V9EdgoD43KvtCy
R6JQV1FKCqcsT48zSCOxnXTcRrZaHEgK69NtnLlEUufzAOmqWH7SPh0iPLxRyMaF
UHnxNzUHBW979U9uLslPVnEN/To5cmZBowrHM0uMBj1NAlufTftL7KL9adlZeuoO
JbiHWx82WDnLBSBYbQP4pORnKjXp3UMZMhBfFeLRSGibS9yns0HtUT67cZiyGh7+
YSW+MHWqoWmXwrQs+nNY+1NdRKwxvIrGWt4R9mC+yV8eIodumnefD0B4GZBce1Sd
SXVdFr5AGPG7YcCvpbk3+g11cOz/nuxfCFoWjy86RI6AbehpsKDIN0cB47TbRhly
30Jnzhky7Wlwy7phcVqYoFLVlYjURiNUgJY9XWkgqlfM7MtwtD/J2RfV8ZhZ7ZlX
FhKZjjNCnH1PP+7lfzTEe7Y97FRcYgdysxmFJe82rVxj2yzbrD4g6MHXNaW/e1Cw
B1ziM22TMf7PfCzziGa0ce9lp9KFcfo9chZSc5dTVCbkKdggUSHMCwr9nAAGctVp
MV9fEqpHsdYAUwMOQyFMh+fceG+iOuoaL69Lx2sGhFvRBOKgxl6TwJrNy5+D1kxn
o2IS78KgH6xaiDt6NF3UY4lllniMQ9V4oPHCI7ozVdUVfCoXWDHFlOaA6SIH3C2G
Beav+k72IkJdk6L57Ez+uyBl5Ru2wCNtTqrCIY8oyd5Lh0sm/9TZMjhnkYZ6mfAd
m58SocVa9x2wYiauiMEPyMlypBLAqfEqm3Vp1Edg6MqV3Bb8LL78F154Uuwy2DN2
9VZGE7U8eov3T08MhrIIZuW5VjEmROjJic/A4hkcVvRpbBSsNiGweO9qrr+QQqnK
RmoPIMTvZ4jPQRhNE6CvN36DPaUzvsrfqbu/rxgf56617cxF3sirZ+xa5Vrr627l
Apu8RI9q4uTsCGA1UZ5fngvN4HHafbAidFOB717WJ4zfWOo875eQv00Bpoq3+r6q
xpKXpEdjy5A5iV1MaIFu915Esdcx/qjtMZdP5XqSCjpNLgoNej3ayLvRfKO8uwzO
IRMsY3u18G+IksT46ky5IqTpPL8rr/BnvKbTo333MyVFhCVnJd5uk18TgOs/DYbM
iKqKfwey9Yz+0inlb2N16IH4s/t18tkv+bw1uCinXkc+DXzgAUowdy3Gb0HrLUM8
PrBUVEtfARhLKypamZ1M/8XqP4saC73qt3iXyydystHaYUgyTnCI5EIFJiApj4PC
FU/4q6dvnhireomHiuc96qjm+VgranzwLGgPnemFbghqZtN2qp2ljmLXcInYtnT3
nohEvGyNcogtWwdoJNCkJ2w0m3QwUJthehl7HbJvECWgTSu4QfzredB7oLP0kSlg
wClBnVWhVaoJSReO7ocSx89+kpU8eSNBeXpZdzfVM3YTGNwp4WnL8W3JAdinJIPD
R+rulfhlnq0CGpTduDmabqe4rEMuBMByeTkzcUvi+8sf0SpE91rjpQzlCcpdW4vd
aR8ocqvnzxVePwhgRe/zJitaiAUMXcJwETU/VOtzbFupN0hq6nt4uBcUNPp0jfG8
CevJf8Jgr7wmG0pbmrjEAttSVMMxL6biKz2IRk5z4Uwmy/7EevRN9Ri8V/hS47gA
G5dDzQuXojENi0Dd+EfRqrJUftxoqGIJQNMYwNMPcrTH7JjOkRdNbJh7K0gMvnmW
kj0a/ZowxXHZqRf/N1Fq2BiLnyzacZD0gNd9UnniSw+vqeb8rdbQ597C/SzhgsH5
InlD6AaLz/X1ihhocPAbkSgo6O0qB/Jnbh6RG+aCnHiSuZxhvPfhIvD2uz1bZ2pG
tLgNoVlqJTl4w0oeOdPHIzl86WVoKDsN4uX54XZogDAK/5rNNwRBf6V3qpCVwrxF
r7onCOu+2yFOiT7/HzgSXEcuI68ch3DjkIejPhKV2mjhMH1oIVAGkk4QKQZ2SeI+
hx2NlYgB51vAjSyyg7l69Xo4Acdt44pIhJ94X1exsyensfyjYtCZWJQP+SKMriGa
oj0sIGrwmHER09k/aZ7C8HrTnpLEeQwxFi62KWtyqfOUDMfn3Z5CplEuDA384ota
qzzcQjA8kIIk5lBKTYPTHUS7IkX/9vMWjqULygjDVsd3Y1KS7xA2+sKulymsPGxI
o1MhuXardJaubi+oSk2nd2IbbVUtuf0oSOWtiFkB3s0fEK6uN1zV3ycuHKCiwEIa
PXOClSXF3/Q24myC10bG9SKDdtD4LK8BwgAj8znekM8GRCuGseBEjOcB/xLcHdoe
NkwgujjHqIodO8mdGGSOVkwqpGIHi5zi6uhbXTmneoZWCkggGgct5tLRktz0E37M
m60We8DxD0MrVCIhsRfiJtN4AdYyK8vS/8EbTXrV2Hzdq6K4dcajq6lxhJMXERkt
riyDU0xTCqiFnQU0IMRyPAM3me164KLXzTIs8/mj2gfG8NykreqW7UmgbN8GGoU9
LlVZNjNEqCySc99gYUgUMw1BgX5vJKBHIoOEJvxF/FFRxKybwSzPfDxJcJcppcyB
FD4y421C/vz7clfe0YMx9Vw9rawLJJYVw05jHiSQ8Os/GH7GsR8zaOO/aLfdQj8H
m3ClcRIMbSnVpPb6lWO4wroaiyVF+phgjw7OGoLHOyleGa3NPFFx+n1yEsUajalB
fUdPetoCyGnZE3bd36edf01aUfEA4d6XNc3heRckz78zYPfUxfKCTbBOCMqsoF/m
4hTbY+qtkVzyFVa/NcyeKajN9sV6fhWskXd4qS72rJJsy5YuwuDwnn3KU7WFymXJ
hHbMFXGrypWO/tu6YV+JqfZBrJkYjQ9nFOHMyi4VcGV/FKpkS1iWuLVXRlBA5y77
s7uZhmxu1hF9yZMN8+ImX9txClEj1gX++HwaQrXDyJH4u1oopBnWyKnOsRp2KdzW
eNQwDfz+0lv2fUccEYwppH0SVpa1caHfWRqDE5Zyb1wthANrB7hhv1TikI5A/dD2
IjnIdA0CMbBi+nt+essbRBfHmhhrF1SuuoKxUbuppCrvGB58L8d+n5MKGK8xr/OP
9cgqrzaAXjbEQE5hXziSNCrCCsC7Gf/xgXkSAdHdKBo4gbK8YDmP5YIDQdhKjLzx
uL8ZP5Gx1OcFbJUEqSlnA/TcTftnXZPNhbcks7cKzM06LxvPel10f7v6mrGCKRwU
Tl7N19S5lbHOeKmJfgueW1bmqvJLUUfVI1x3p/9g5ylKpglZICty6Z6JJ3xryQTU
27O+gZ/Gt81lZwJzpAE0JKu6utbEGeeYuBT86okgFGvwMWLgwL1eQ9GNjkR+byma
LTDx2oY2wlgWFZFOnjqqX3Hd6v2LpsHputt91f6LF7fVTZ4FEbHakSp2s2/wI7Ku
tBFYKIx8qeHrSQfkMLS4R9D3VLJFeZIXtfs5wdCjxM81MEKelIkzuyXvc+Cofdde
+naXRJi8TGEt/gbax0X6/Coq7j0PfxWW4VpoACNYwDTwSObsy6Cok9F629p/eBSq
CqgW6muZSdGumeYXH8/iS606wlqPh99CtwKew05MPQmr7xihsPtSQBE7WMeXiV/8
7V38gR14CX64vKL8lqbjDPYfkaFfwUIdKVaN+X+UX7ASXN/5roRdSP+22zVjkZHq
rpb4kfdAzj2fw8w7LJHalNxL9tWcfwPZgrg93n2doCRFZT+InpFR/UqhYDpvYgbM
ECPP3ue4ic/gIl3oxUwIoeGu8rOfju1aZlxuHMiG/jNfv26zEGeA8VK3PDFCBXOm
NE1a+sEZCEj4VLHN3O07i10VKC7SyvrhANU9lLF45pPPKIu43ZGkU8B0M+OKScn2
XLU6kx27ne83qhnqyK9RKxy0G8IMUYsnB86M1LMHmMbHpo/YanNJV42DG9+JY5ly
oKbRt1iXN8p/S5fABKXhydKb6erGjC9ML7o8slLNaHg+eB3UsbnfbxV9VUrxja32
zHaMwSVfmyvmnvQNJOOcLBqjoswULcpDkLElvj57FhbBJmluz3vWQmqZcE1VUvP9
ujBYNtbR9GjR3yxbw/bfanFMxRnIOI12249LLatS6IsB/SU5P3+fKxj6iiGft1S4
p2ZyUqTx5LqOHJrR0lXF+EOBrgZ2X98blazFI9IqTIEhPuVMYEdllvvqu52gEAZQ
kFNellFpjYZSsqiWIjh0pEFugHUDfQw+mVFH7e1kaS2NSKMvWDSHsfbbSzS0WLtz
/qAoyDmcDFdD4h66erA7qDdupCY6Xpk9rYJcifcDrqBNlEeWS1V5rer7us6tGDAC
7RYiMAb7awAVfDIxay5rMpOkmg1v9ktbzNMpX+NVPAEkk6Sw9PSuNX+KvFFXG+92
5tGRn69IkNckbQsdEO8hRay3lu+pBwzHQaxfI21ohCZl8oSfNn+GxqkDqu0Cw4o5
BIcRvNf0bHz9jnW9UaO5qtPVqNtY4/FcoIbBZiqpbHIl8gevMMVQTPNRCqOlADvo
swCKbucBlt8oUQoH7OM1UBi50O4tg3TWra/GsYXnoK4ky/6fzK5tp+5YvEx8gmqt
IUtKA+Jpcehdzpql+zf0+0Niaw6KGpYjSCqkwBMyMz1+cWTOuuXvc0G3gf6peLyZ
TtG6nTgjteoWZeBg2ZOVxQPbCltlGCQ7rn0ex/6m2PbdZzNuis7vbHaFYo9h2EwQ
OfyaBvr5DM/yN6rH8MBNNvqcK44fdGWUrWhxV0cxitaeQ1qG0+On+9SQkm9R6HRI
TZWD9Cng96Hb4IXB1bs8wrUQgxLJJ96sWI1rOJ3sp/XrwQyZkQyG0RTGEdCLfaiL
tPs+AglCp7rUakzXyN2xiufakaQbnlUOfFfB8okYRbkmxUXmpusAdUh3+x6x/Sur
1zhZVkg9WJWHNsCPGwFt4GpnfB703cAPL7rmnGvr+UFGsMLAyFrJjqLCwQ+Vg4qZ
9w6HrPfFTRXaGaU9U/IVpqabLozSS0Yp8n+WUOKpVASQix+hAFkpRj87F4G5ork5
u7aWcfBjgv8yKzYjB+TUndTiyv7sBW+GgOUWtn8LqAHSZfCkm16WhIyrCEjZkaya
ASK0w7SjajzSRpjLoDewZttFZEbD8fDjQM6+B2HZh4yD9X3Xjt25qYnx3W0tydIa
4SSRG+zmOlXDybis3goKiKgW9kXRD/KqpaEsWFqsPwSL9FtcDit20lW5gvBrYybs
0FBTudkj+XLMYZ+zw4e+cqbY1vi88iaZ+NjwrZP7rsXNKuS8bECyTWPVr1q4cD6G
1V7e9cwfh4rAoaqOetbkVzjUiW+n1VKvWe7r/IKezwj2i3ipxllK0w62VL21dUjC
YK71RYaNauVPdtwEh6b2M43nlMn2++ZaULXr3ToalakBI09ODCMkeZUOEPxYCCkF
V5wMUL4hlmx3eYUZC3WDTmbMLxI7S/lHtQHlC6ekwTkuq5ZlAmu/T5bQr7n+NgTS
hyyJ+XgdBlDP4n8zlYCFK7BddwUJv2wkVYnuHUW4W3G3smFdKL5oFIvpxoV7RQF3
wlTxm9vdVn5jOomc00KsAlkWmLikgI5NE1WpVVhgUA4LIc9ABwYBqON+SPg/toQW
/EaeYzaqSxUvYgnAXrVpKDn6O54KRzmhIzdgWc9aMHMl1Gg89U+Zu6PFA9FZiZk5
/kZCj9ZCaMmx/Da87BrsKpsbmBnwtkJE0ITZ+YKdQDDb/GkuTqbVwAHT6+UiZqU6
j8+XDbIF8QUoUek6FOOIfz2W3he41PzPRlyVIduYGQA87sR17Bfosy3gpm2/AjDC
R+/7URrJMn9Nqhq413lxS8Or9KrRW6ftn2vp0c14u4xKR1dcHASm8g33P5p+W0Wo
pciwXcA+OC7Q6381w3YAIBrDBMhyZtRm8GXSzmAuX+4gCphVmzbChDJ972lnwq+1
PIgku2tVIrO/KJq5RZFJFy2UxZKh7XvKeuURfZ9nEvwlb4fjdOYNIoVmAnyU/Tlw
D31BpJ6s3Pno7vG6bTtCGooKULMhBlLVBzd0NC93FkrObNo4mOUEogoFYJsUct62
g+lufO+0UIj2w6mhKA2GVMJQtWdV0vzUwbHOPoRhAo71JRcPx8L3XrLg893DV//z
obYuktpnCznx2IrvLVxUEgUU8ryUf6Q3khd4WexmmBSW23E7Tkx0lFhIUMisqNz1
dM3MRjWiqF/Y16rajER3E8RjPR9BTAXuBCqes203xTP0Uj5/FcwLDsUjmwG3MtBI
HTE9LZJUCeKi6gHXvu/ANqTuApg8s2RUtqWyGbXQDwHWle1iqk6O9Yes5grD+6EI
0b9fwY00eb1ojwcIgsqVwctXHNODjAk3zsGZ+HaJzd8X3dYqkJjcwd1fQYqB/BlY
ChhY4ifr4uiXIcX49POaKuqAKqp1nTcj2+eMSLEu+15kZL2fu2L0US2yrsbcm4R4
4niCfKSOflJxPXv/KP0YziECaAE76y8owv8AUP6EZRo9UyMriptnyKpt6AgAkqE4
F3laKqykmhfIWBhofiLHhGcgFwfkAxHWE5rV2QGh2eST2VojrQXt3sSTTfn8Cbfm
4SpIYXx4OYHW9I592fDaAWOqjsLuzWYronCbvMnerHuKZQd1tpS60uZpOQUWd/Iv
ydzbhXndgRUd9OMcZIJb9dUtENa4k4WTic/B+wbZzYPmP6KD7rRPQedXlSzbg2o2
6XjPrQTxKqZDAu/1JIMkcHU2bKs7ThHQWCeUstlLH7qr717GF8g7GkJ7XCwEdBMO
D4vuLL6kIOJcSBbhxjXhadPZFoxqSnowrhthWs7lBcFQOCTF0hWKZvT3yPoo4F/z
UKNHG718H7XupMgD8gBUmdBONEm4oH118q0GAH1dleqP6ROiMZ+DGXLQvagV/IDY
Nd77n+HsE/Lx0mqYdKiL2QeHaY8ylYsK2v1Q1pkvOAFaODF/K2BgVurYMiyIt0NR
ga2sU+fu8JnxTgNRzNLy2YndrvZtznJIabj1oTghe0o3jah+bcvFGuIto5pmoDHb
7uYlXYdbwjryyXap40ODlOxN145zfvTIUFnl/F5yRliDvu8HKiCJn2D3F7Sgh9fI
aaDr985nlzNMPzyjrooMxxJWH3RxqoA+HW6fowy+qobGwD6Nu8GfI3mfxXNUQGxI
wBQ38vJjejaf2v/B/WFOc8MzPaRJCr8bhU80BsZnf8Ukj4uYa6S+zqUu9keNGLJQ
mP0eWZWl5ysx8D9qTc7fD4nCyDIoxK5Mc9tQ0tDgurGHauaBWASJwKZ3pzWhVIpx
tSYCjvnoqX84G0uqkU/CzRBdO4efqB/XFBPazt2LebgTXi+Ra0gPXemNFxixtypr
OmYdLSjIjCKtrWdiquG7CJPABGxuuk7TAMcXdRtF/q2sqoCwbh3neboDGyz6lXhA
pQgogrLNO/d2oq66k2t7glq2Ov4xExsdeJXLCybzePli+wbornrt7lRBHG0OdPJj
9RlHHiieYEPAfpeG1y7wqYKc2TwxVUiV2cIw+9G4aeLVKpNH1Jp9QuHlR3kJtaxX
/bgEUaY+UP5hu76jn2aI/IPBWg+GZrKHnyxusEkeuYLEcVdyHCE2KXjFQWDYBUXT
m6bW/nFEAK1C+mwoKjnHBTPKQrPYE8IaNreHrjTOMVrGq2UcGi3NrSQNT1D8Qgvi
51f/OO6YnkvxgnBsUj7eQ4nwgY1B6zfWjPrYu0mEjAg7oetVuQDvTbWWKSjh0TEq
WiAn6MCQ0IDHhjs/lfQDwj4BGraF3m7inMrK9U6yKI82WXY4JF/nwS3z8EsViLVk
kjRFEob7WQveYJOwGt+qQEnzx8jvUuzlwyvn85jMFXmmR6KTIv7zMzNeweIViewF
DtJdR4Q5oSrWelcG5vKVlkAgYtafwSBQoyzi8ia/OphwTcGtn6TCIW9icJUp6sg/
L9RAqobqCXkF1tcfhUJU8OlZaCiFXk2yC3Nkfb8K2ne8Fwwfec4Lr/4NGxYUZbgA
AfPLCYzLnOLGOHpRdDAU6s4M2CcB+oKHnqkoXdFffcJUVeMlT6WBcS8vKln/z/RH
GIWz30U58UQLwkfyGc3VfNInr7L+Q6DafO/kn5gftffsHtku2PLOMJE419J2GKCM
fJaDB4VMzDD4/dmNu/E1LjRdqsFzRW+YAxHYSOH1LWO5Js7dMao+U7mZFDs50k5G
mz3c3NE+hMm92xUjjr6OtQC7MiFn8iYbq5zNmiUCnr7haXUH0uLHas13tYLlPTVR
JTxoufZx+X3uqhqgZHa9U1V1zIpvydpyD2b4obRg+pV5D6G4GwMauTN7WsKjFRVb
go3ZPrX3N5+mk6/eM8juqNWwVzws437VhDEh4Zox2Q1U1JqbQQA5PBcR4zfy8WM1
hUxXz7wCnK+Rytx6nOKQnqQI+PruDre3h1mLzFW4wkSMnVw6SJQLW7YNaUiY2nW3
1ygy+GFXJNP12hB4dNGxRCYxdSndqYsGZRmBXaaWJX7Wv38I92mm44BumE0FvQMx
f2UwPLuUjgxj6elMfjcaP2kHEjaTOCgYqV9pvV0Jc21S3wbUGD3BoYizfyS5MwXM
TQQFqT3JRAvaNe6P6xZzgD4NyTDq8aWVZQlhtSeP3s6E0UnhsjkMs5/Ha6sQKdcT
iXT+8xiQ43mI3ESguZZW6z7VihoOB8m6KjA9Bk5Ytt+IRyLrtp0TZXMwS6VdDiY4
J1mCMn2NqtGKAzIUMepC7ju0OFH1F7CM7QATWxmgCZWu19rUfM3oHJ4DDO/Ig4zb
4lXfDMKFFaavlXw0xGDEHab4ueKUOkqhIkQJX5UkifZksva8t8cWzjYZrcJpKTeB
rJhZRmVlgH5ICtbVBhPpm4xhdqkNvO0uRW6TYMntf4eWzIHe/dwgKu8EZeslk1rS
QWQPvFPEU7i5WDJy5fiDSoRA0P8kYQPCvF3jtZvBclgwOB2jcKQJP0p8F/O7R+ug
fAcieey/Oy7QsYSuCT8pEh5gF4cttV6m13zC1zKadXxNcP+PRdAgOwfhrZS/pU+v
FE/liUcbJeZoUTOousI1ao/iDx3Wys6DE5maOWhaXtgKtHa/3utE3wlUqVbe/B2M
/YP/csIsb1PNyrsFfaWGXHOeKgOCKX8jtbgPfMqEry4M9YLvViCkYGTrvp2bV0sH
YK+Rys1UWIEpbiiWgPEKB27QrM6IwOVzxqQj+GktMgm1fdYQ6UURX3pFicR0sc/n
hNlsKHeUKOhHh3y351x0Hk4lgtpY+/fpzJPXmyOeeP3hRXbl9er7QhH4LCSPjNu8
bmtm0ZObqswXp2lLQIVHjdzCoStwt8UAjKG9teNf+NqeFzXEnvqL6eYhdCydENH1
FzifqsDun47YqKhRSB7vzNZqYWpyKvuOBQwBllO2v8XrEHE5Vwv0wlrPqOhe5eZG
fIBvP29GNuZr4QM15bZxJ28/rruzz3hbtRJi3cDqv+Z7df3zMhECOv6280anoqt1
waDcd/Wu4guroU9mpweHf8AFgEhFnVtxbOauPnQVzHmZmbkBg75fxsFV7dyIQH1q
iI2GpemW/ZfVYSDAOKKHIz22p18UEh1DEsDdAxdOYFoFL7mxyAQ5R7+bRmS0KmNw
TKCMkBjKqHTTHZ7xle/KGC97Q8okCDiThHUhESDaZHynl2Mef1cPBgcsrghjn9PT
TmIk6X1dYBrA64+7sXOyckUav14pqhNQ/2oaNgRy8rO/JCB+W1+YAHVMPT80knjq
Nr78D/ZYa7DMgn1aqtBtWz3db330H2NIRODwmkH8uNHaMQqVhqUApvuyt6WEXGN7
jGwhJhY74MhkNRJsqtQhv5NaMtfJxDhmCWfPDoccSJv2DHFQfvrHV43/x0+0EFWC
HHHfYH4vHbq6aeHazLuk/KenQAkgvuj2phVeSursdKCRnmqiOwNgRW2rAESOl5n1
ZunYewONUtoNdOh4xmX7FGzTd5jlU6SJToqQd+4U2prAuiUJ1Sq+gFi6SsrIWtAI
YHPwNXQMgCOh9PHmbx0S1nn7AdY0HPJqJ8WgGjvCHQ5a4Brko1xv1MPIxcOs6qmI
h6+YLAx7LJs61SS/rkOiDiH5w4cKlh26QUyeK8uoE+Jo0hGoxFJmgrTtL+ihpm3K
yuroxQK4OVxR3TtOGbPOt9mWhfLOgTRY9P+HsxQpSWtrcME2mIAWaavaKXzMfgti
O+dgLD3AQcfyT6KTZHoDvbpga1rs55WJ4xawATDHSO9919v9FZPxTBft730SYV8N
iAa2RweMy7oqtO9QA+etp9/Tuk2baadotF+6yiUYPik+58N4F4QrMGmrNSb0evx8
DrB5GLfvS6MC/sqNIBRBQC9WgBEi4vAtXgz3vMuJ/e4HDDd+nOYzE0SLeihSd+Fk
61NZmslAI6aCrMYQaKcOMGfNq0y5dUV0MGM31XLwWU3D/nzWS3+ePz8baGMY+BlG
YGWaGSWB2lZkuoOQcBAY3e5tiGyso/2aMrUjb3dXCw1tDZfz/rvxtNsfzLkiM8J5
u7NnPU6FkebqB5IWazpn+nzUXlmQMtKw3RQbxjUZ5yh5hB3Nwua0iKexSa2+uS68
8q5OF54NYTUgUPSj5S5ezvXhoSFCvdPgLXEDf3Aluol9EjDCMXNgAlbGxUOEgYip
U08t10WhnGaqIOWb4S1pJ1mrP+/r4DfSVHfbydjeLZYEUoAc0ZnOFPLi9h6xmpEJ
OHGUgHKs3b+sJ/2FA52+Uo/nIVbsQhFXAObkV0VJnIXJCHRkZnYTMTeqsQFIArtO
pXqRPsyPpz0+yYtradWKEfH19neap8oBcs3LSrJxnTukKKuNfb5cBM+BqEMHnUy+
+ZQzLrV1b4PnupHmmKXxv8P4TR9b/mylHe0mU5km8xxzmLst7NFFLhtVNbho0qAn
fNmsCNLWe0WZEIw54oWdcdXKJcEkMbkFvyxj7RiJlds5+qIckf0NMG3/1jRoz2zD
83OSm+FSlSvDflqV7fqkHVU3VFwalL7o56i/Jj6Y189M8lPyr/Z6AVJHb4GpqPZU
RwoAvEVO9YDQ3BTZvyLC3ysevM8e+QcLfBo/CrndGnM1EwlMmP8B05xVKTDS+52F
+ntJZH1y4E/rv1IBAtbf+tqcc7/nSWXx+fTHvxQrOzM4E8CTriumU6vgDhpT2+Jr
JNv1x+BCU1W0kIrGS2maDVhOdLILhWtotEFrWo6fbqN0bXztSe3A9ph+nY8Un0+o
/rX6Wvafy3KAnPmoY4zCWyuy0AE0IlC+1e9ec168lmsuRxsVm4gFnC9uz3S5BzFm
uz0PFGIZ+BVC+1xwUZCeEyl7KJYL8q8G6mR0xDhs1x7d61zVD9aD5DLzshTiO0zQ
A1QYRAIyTDeS7l9KwpP/Q4qNZdCvzIWP0jVVlw0McLMNv/xvTweCsKRjHvYVtw4q
ovVJtG+kyLrpsT0iubBxPWVwqvbxu5bOiFegqKtxwfy7CzygaAGu74YWpgsWv7iV
KOPMcdPiVi+hOUhsC23oHx8tdm9HuxtO1evKA43PO1fmIY9iXTg27W3epeiy4BIG
K4su5eMcRGO/rkOS9Y6OVs7GGGq8D4mXsHnG29ZlAwS82YuBYk73MgDmx+vwkqJB
Ae5ynrWIRSN7yWdiOBEkN4FFbOfEGxGMvk+5e5HOwWmIDvSUh9TeHhE0qghM9yvN
fLTWWivE/LFkZXNyHiUXuyYl172gpS4HNNe0IeRMLrkGc1AzvveTahIV6LtIaZf1
V6kMzJQydTHfgmYg0DnQxW4i8AfuuK4JleOK+Zbg49Je+CuvHkqC7vpBuRLb6NNN
dyli9czVWWCdhaW3dv6IEK/sWpburdFb/Kti0G5T71X43ccypbHJ7UknC0XRuYdU
boPHBFODczXToGwRuRmGbvUAnFY8rBhdWgO+9dmVHtJNcseo0h36JLWbyeVADAh0
2gCGjYCdw4FmW7h8bySpZS5lJy/t37W1KIf8Fhnuf6WIWrLjPYewQIbHTDOuqn0V
VGnh0yQUnKNJ17Rw0jQwnrsbQD7KPqjv3WXGsS4R6FPva9neQWPuDO0DerevzZv9
5UE61ZlZqnJOWV6/7u6m8ees5ibJmFiH0E0M/06QRwhWAPupsgcrY0KbMyeBAeTo
QaNwjXD8AXE6gfi6LcTMSGxhweokr6ygd4PB9eNic5ZXtgSmR4uMXJN8TnaQg40w
QZC63xKao10Hzw7tLdyBKgmsqTxQ3pI7cjj0/LiSZv3XeSTC2yAn4c/zVovw1x1j
w4XuRcLfJGWLOth7gljf1Qf0IaEKmdKfnX9ytzLhC0vkP0LDGZ5ydK22PoH/fqpf
U705Q59FkfKA5rXetttHF22sGbozG0rtWfAJl//sWk2U/nwVbrMx5mzmT3A5xNQM
8TgSO0WucIA6ehkpfQiYO3gm044gBvyn3mmWC1uJU1vf/Ki1Dgzo3wmFw/4W8NNG
xp4cnA7AZVLBuMumorfsZQ5hIrMq9FkVfHwb6kL3Os+gnkmVM2+qHe75Molxtdx1
nKVPBi3VWGpA1A8ScX7rYvBMJ6yOM9urCz1RYMPjwK/pXNb4P8xTgkXkNUrO0ktU
0pUu1fItEh8LtB+K7OK9DlrHG24V2QECptblBaXAf77vGgE+DSh6I4lrB5N+e9AC
3c3YLFfmjv5ZsdJIeKO6ZlVRTYsECS1iYV0YNtLpivEHxiezg31QGb4YcROQzv98
jjZoXr8683mxlsk7f9Q+N/s54DJZ+7PAvFnfqgMrRDhwx6uTScVUNe4QjLbkv+DA
T46soccMTOTaFnuBVZYsr4tR9ssnkEXsyRTCXL2cP7MEGx+QtzMPUAkj2jF5KRYE
Q1xMfZ+oMMB9M2lz27R/dcRt0gGR4TFwm6dL4a+4xYhUwZJOnbxLcFssaJVnBLAI
AyAEBUiZJgY+CkogmwXHzpgMsYBu1gf5vHg8MDHU+KFI3zfPbg53MM2rAHqxq8Sl
yRYLZHw3uqtMiLxA9wHOjDndQc5mAIBAn8lzg0qDrPAh27+Bmink3HFl9MVJQLbO
jRdg9oYo428kwGr5ey40132jrmZK6S+/tni2nYmkY0cUHN9V3nhK/tlpWxuPh5cI
BSehkPp/2tjyCMhiJcIyGIx++bFAAeFVXrFZA++HuSzVZrFkHCGPOTDU89UbJNMN
kw4KQCUpfDRtqBsGBzjHGpCsgYaeYF9P0I3roT1InCbIWVGc44G0q8iYGF5dJkQ8
2ruJ+PgW0K69jTbGgetOzv8rpcQDREBzeLIehANMn23GrtKzT6Cz2OoQpI0zNty2
XWFduf35voOXwMSUeWMfyLl4NZgkVXCn8Ht/lYeTFTlykm2QjqE7xkRErDEivC/h
0uQM5a3Q+5Yqcj+lPhdjej36+3wzEL0+F0YQTfqzoMTMT6U7vLj7xHRqLJ4qTp99
T2aTHrOhszJE6E/UsXLiQtALOjHZ9ikgKIqL5MdeOxA4Fx5WIlM+c839whAU8xWl
Hq1txHwnLtxK52Du9Tcx+e2ek2y2Af6cPbraatLnX3rkbc4np6QZp4ImcA2f1sUt
/+NhJUKiwK1gyFvdJ4lodvMXy5BYZSKS9wThTd8E2mUu7wARAlzYuT5N4sM7I4HR
0j2AwM2Ob/ysNQbS2hZFu/Rky1m3nN5zbun+C2eSxMMMZyVDG1kXYTZ9zfxdShUV
WnqB9x3NW9iGmAkUJ8LUO220ktBh6HuglrJG3ZLLPv9+Xqfqz9Q2qX51/FsRHRRI
a4g/31yYtCAmOWMw7H8RszyuG2Tciu5xSGmySbc15/vr7komT2vFTLtYGh7gbBPW
XGDPzIGuvFRuxIRchIUxqgwuShYYbN2HvV9iXgQRVWVsS3Nuom8fJWvKMtJO+iwP
CRDie2Tl1K0ARI1eF+TBfmaXeh7y5AHZPbpxF/Suw74/J+7Xy8ISHbrlI8qHfHn8
ZlGvJLjBp9OiIubMzhJbW3ql4hilIZ7nlgOU0/XrOIUbuDEc7MCy9Epig93GplPK
wg0xO5fgYz2qlDCI74vrFvN620U3KUkHmgSCsarUZnuRlX2zmfOpREJvZQU4DcDZ
clNwicoAzJCq+YwWWOy07MGk4Cp0J1Igk/AiUu60jyzO8CgvZ1Fn0kwLLS8bU+z2
/Ks2Z24CrY1706Z5Ob9JPauZITLtMzeMYNUEEwXIW1OhbwRs7cFKpE/BFcc0j0ZG
Qf5k74ouCQ3/UgS0C3I6CIQoeOaeFb4SbW6Z1s80ui6Um1slR0/+NygKIZgar/G2
7+ylfEzqaOXasxoUOPXSVxRz21K0aLI8wWoBoZU/z2EtczGGW185zyxUCXDPjSgK
klzwEwxjysOjPtYAhzoS98wb9HcizPu3TBxh/+4PCMoiaO5bsFDQQ3UzdtpoQSI0
pV1/DwtfaXxTHVotTTQX23uAqXDtz5vd/7MlKnQQnZySdvFngNYf1wDYkePrDuXV
e581ccQhzFx8v9B/QTSmN3yfV6aAJG2zPYDryHQQeG/zf5MmSE1SZL4vIYyHWld7
uSoIVS1ifhm9ygvYKWXbo52h3LYqZ999hcLdrLofZVafmECGix7GtX8aIa6wd1b1
fLh0nbGUT4DKDPl8JZpZGIcnB8pqmgGgVVkwA+8SpowaFOwy/tQwHe3o3A5MJi5G
Zjfk3971Nu2HQnsJFg0hMNZqGW4bTh5ymAKZHy1yhAHkO7VFaJJ0/B7XgHJHCujv
fsLV8p8ycqGAi1aKTnenUbbqJEMhzb+4HZHwGduAoDqZXyDYG2uhplHYC0EFjFMl
YNhumZYbWHXtzBVCC427HRAco6hX8uoLvuDhmR1zfpJn/cASxbH6EwmDS/TtKa4j
0MLVTf6iA26785I2d62pGKyQVhcL3ecmggzOiS18cA7dmPe1Ywn7YeKxVS8zM1g5
8PaKWkqDRIYEm50cIzEJIrZMDGZZlzp94zNLsPsE/1vjQFT5pNvkFtywPyKHGcvs
oNmiZ7aWC73Bh+oyDd9aL/4wNSmRQ391pbHTQEvYFqPxPO4JE66zVMk6HuY6BzmV
bdS7aPN1UPDYqt7fnsRlQWxi9ao/pQ6OTglcBSmOJ43FRbknlhENbw1SA+/YFJVs
PGKo+Kdb/v8hFZlgmWIlUlf/h/+EChNjSgDvcJ7u0T1bgm02e7XQUccG8zw7Uwo1
nnRRdT7Oq/CUqdgl7dkvg/OHkH4YvCNTzgHYs1+1DoPUz2yrfurpLhAXaWMe2BtA
h2yZTHV9YhEQXr31Ph2YYeIhnnex+lppF7/qc4ilLLqu4ZZdMuKxHVAavS9/G+V3
GZor0LRNNiGMQWq7Xtr+Lort1aBz/6Blu9jRGiGCdQ1VlU3JvdGE8zXrapuCIasG
Rwb2hRPvXJFcJzKT0+NHFd/T2qN+r2e5VOH5HHeItp5eaC8VMA991N+XEfQXSXGG
5kK1LfgjrapJt3fz2BPhfVXJnOPQYqGkTjhUV7/69kgmZTBLMSry0+xRwKb5JffV
Fc5o/PMLISXnGWe0D317DQFMk9NaHsM7l6Jqi0J3xGI+pqmnS04jF1mhEmnzaR1J
wTbui6dPYaG9BXaHqAb1EzjnTNqn7fCo1HnGgXzYL4hcjs8BxxgxSwvCxuEoHbsQ
Dd1Kb0KgAX+EqjvllsLZFQFjku49ZCXhtIE9JHM7/tfv7XyOe5LVF/t6qns4RAVC
5pAKkOZh717KCwAFasAhX4MQHD80ql/jjhyJFJ5sr/UPRvq3VDbB4T0MoOpxVif7
rFQF6Dt+PdpX+xoobLevkm0MdE7fgncLt6P14k21/EB0Ho8KwkF6PoirKuHea2pz
i1HfdypKNGh3ish2tt31/so5/1iEtYhuE090EM8inO/alQQdGpD6uxTPSloyOUPo
0sFx5pP1pmHV5yMzKMIIIU9BMwl3eJkHZ3p27/a0WP+igFL3uDEx+qGleIIZ7bIU
RBwMtRXxS+frq/7WtZ+Nr7HfgiU+wSr8fWqddZs+JGXkiyoznUgs/dPDnB2smbo1
hBFMtHwuSVcgy98AXkKbJ6rCx/5ug1Oucp+pUITrZ1TBMZne6duokO4mUWH9ItYC
PUzBjaWlIKsBv5jv4nt1iVIGJVQqFN7xJre+ZfAwjfzIyyKTOyypwSZABwW+UPAS
Tyj90NcSS5sC/i+/m/0y5I8RoYmZsLpRyMobx0M3v1liwbBz5V4i3WheWgAW+ckj
qsi1Vr3ok7oJqyTRzoBmowcfjOIjzKt60sORqOuaNfkFB+8Ts+wR5TetZ4pNGuF3
mDY+yZ77qaafDuTpsHcI2WHnr1+2YE7iZ8USpK/U/GdUjIrwYGb8IFzw1NXIlena
BMlWmdYLJM/6q+SgqUWnV7VDDSUtL9ftOk13aJuI3PdLUchba7NGBHJkwGLXoefX
XjMV9+zwAQO7e5QWj3ZA2JUMfvtIUQKGz2eUIKA87cuopJNzRs3VdI4Y216q8EAj
lsP+Y+Dn54kAGCK5NvoVck5iLSLNd+yXv0BmcevD2gyubDJRjmpGGbulAN1yk0Ml
QlGynb1h/yV9066zuNW1G8Q72RpgtU+wLh3m8/NHBq1mgEZJJXq2Fo+sf8p67v4n
Jkn7x9DJp2kaenFQliM3zteU5o74GG/nRjQg4x+7WY2uOGAXuja69nvPClH/LBAt
s/EteBJFe6BKwJnJuol0vBe6rYyfEBF8gkNChVL7Vxvdhb/KWATBDHm1s1pz67cB
aZ2UxqsCDIoBYxhWyElu8lWHFkotRNIvH9urxc1V2Qi/+DsLOl+Bv/Is442vhlOd
3PeaZGcl71FHRxi+grujIiW1joSSadKqbu36cp0pvzrtkJgeiC/5WIE9XYuvdfTh
UaMoUqw9B8JHvO9VCcIdF54kHjJ4mMTFHSgigP9GM2AHoWVZ6PcFxqwZ8rjJfadG
+b/sNiTKLjJYR4GXHaKptPkj3tzfdccb4K0mF4D83dCnvqQmMjniJWZpXYud4xFz
ljJnjwHQn2gQ2HHncIX+7y40abgM9/THwsoYuHF1ImRPIYY30n4f9nqL8fvZA7JL
Uzo5RvNJofiUnTJ4B8IWQAZdpW40aahtwseKTmNcNpcR003J/Y705X8T7JewM+dM
WXMDx0toCDZB11Hbqhp1H5p9GlUiiZFZXyGEulu3JTEUTbNXZ5MCrqryqIzMEiMU
GwJkl1FcZVUrP3RxrUGLYci4PTwof3nVbA94+CZk7DiktrC2XqSlmNoy6NAkPisU
MKSOp3LKjZ0Ji4fYgrmNqqygudxLpL/WSjw9bwfv9OyLX03fp1MTBopGLkTHpTGi
TJvVuXe31qC/tpU1zcncz6N+P3V730hV2AhuQnhNLOOI04pZPce8NwWRa8VMipdo
jE388Fa5fR8Wxm5p0Djq4HBimBJO6sMBvGCzoHxP3A5MrGuTVeq7JiP+S1BazH5Z
uMcjA6dm2gOendsKpVsCG/5a+eCXI/tP5l+m3R5BCpb9IXQWHsaslmH6+Hs+n6LE
d5im27sxuvZgpZs9q/aSYNWRPMMbVMA55sbCNExXfXhZ/iCGmL4NaGL24Lgpv9oj
XyJ0ruvL+kYIWP6mr+6Vc7ooqnxhtUM4rjGjilClCBI/j0F4FPR2eUgwvKgbEzh6
yp3KdNSbson3HQuKvB6/GKDS4KkddrkvZ1WGJUgJ+yAfoZaCo3wotLSBffKQ+ITX
A3QAjbjGSr+iMee0SvYAZfqdh/E5fXfD5AJx9PyWkmeAgFCpv2Axl9fjP5G4M4j4
dNqdDU8VxKtVANd8CmAq11hprZbQpssGsxm4M/pfhmcrlgG5zkosGY7nHFWpPLsF
ffsBOHflSrOsCx+fQfT1yplP7AAfFWc7C7BEV0EiMcOXJYofW+HA2SRbs4TGHzCd
imFOoEm5TQUmSXb5mW287XRmMRV+KuFUSpplUitUf9hcCKRznz7pcMPVTtT8J1Fw
UCsRgJe2Ix9iK7F4bzcq4gmLGQq6SWTPQqiPYcO/f6h4M4U8xmVb3TtpwWYVRaKc
kJCVWPF4GAjwKJ6CQph7g2p7SPRCgZ3zxJ8nymLBlIMrUZjiOxyefa/IszmI4JBd
4X6epJ7czGmEXQFo22m7A5VXWK9gDmC0WmYzzGFuk5d8zLBaGdPX32/8Wz/PnnbB
ieuTwCmyyp6SJ+Wqi6pQcjim27vUkpUbP57KfV4bDMmh1Dkn/ieM2c4t1IClrElx
jdQQ2hNTOPvg3PPlRWZPPmvL8MFz1/znj2aAZyQkx8bhZ04fc9lhwHdtgLI9WE72
ltvbVUhgFIwqeLQxmpd7HxcTenPjthuY2HQcvnI5FbZqKygmGfG853A9ohRAcqgy
awfsRp6E0+83fzuvUeT2VkPKV26QOyMr4z91tF1hRPjGjO0Zl/Z5o68LV5+0SMXg
rtBZix7kaMTF+QoVADxoCqPyCUPwJb/SP6adSF1AbvnLAY/hJ84oO7lCiIDQYx61
RoyZP2s4j+Fo7xZwHNaBkmYZDM3+ANKpcdQAYDKTXDjvcl4+ed5chXEIz4OFSMqb
8Pk+TzdEthrDcX0WSK/1VFlignXpkdMFjPdWrGbyYcLnPw4ZbM+vwAwtDeQaKrwe
RrF679EG5V/GlWHLAMvFoaXl1tZWBP6DC1SAgYP0f0TYrktyplPcWtM8UzKI4vJM
QCNO2WWpJp1uecTkpwAAPwlg9ovLBkxATBBZB5LR2EJK8F0v5uFgPzEt5yp3Qle4
SLz7RvesrOs47Ih+N5iHszUVlezC7VSZhoseS3c8zpUV7W0jpCTNuCWXFDe3j9px
bT+mbpkzy2fbIPyoHk7opLxCD/qrFcrI+E8m1ndUi8j4KIFtf4kC5st1ai213jbn
SDuQmjb9wNbsb4r0oqxxf3D7oyGqRnvV+0xhsKVX+ed8v46iyDW1wUqVGsLGZKYd
p6lISULFBUrm91WkoZyIMu7H4UHGuxabEQVVSWbsQ3WVqW4tv6mlQ2R1+j472V1f
PBI31I80Jq0m0AtIu+oWccSGB1SGGSohUVYb1OqcEEWnBFQ9GXMTiueWEw8O0x+8
YN7JRRlWt8pJ86YBOtIoekLhd6rZ8tTWJ/1sTlWOZv01MlW4jJ0yge+yyo3ASDRs
vBXSwIQpWgoh9r5DO49tsmT4FdacZp9VTYZhub1KsY6JZBJRmNzOcld+95GvjxVl
FBqKX1lf8s6U77LqwDM0BYhmTXCZMMzOk58tTIe2ePTJEi6sMmEHndHZpOb5Ml3e
s/NbOv0u7gkw1w9xPTpZGse5wEridZMplxiRP2eMn9Ngg1fEmU4xVgg8BgVl5QXF
dvO0XNFtu2RL7YyFGd5SjLh4MirrJFTa0SXJz6yNHsaVRP6f/YqwBDYyUYZ/0e9J
l5no6s4auZV285vIdgHWU9ru+/TJ7ENXaHACL3DLCcKuc0qCKVFgp7EyaNdzD5Mj
AeWcYUEQWTUNnsxmKhnfwusAqdgfPusYwh4J+uFh06hJKPwqeXkSYUehEQEixSzw
jEsqsKqH1fXortBelFsJjKS5IhGKlJ1Rdb8WOMIiXoHt5tgEXJClO/Zhi7s18X+c
dL+ioIdqg+yViqCRw+URjSDnjgyDyPm5GwGCopY43uE8SXbhZBdlwFYVpIWyJ0qu
Mg1/DpRDWtgEjEF1SPdJfQFd1y/koXPsvsMUckgD13aANnUCg5AYn7BKzvBtE/yG
cPGSy9+GotmaS4joF34FQX0e0r/fookfd9LCl2srXJGKzwkO4YtuzS3FhFbpioKl
l9CUTzjjw/9bBNOhFovUD30Ty13wmvLq3RV5HrJ5gAeKivHCVHfCOKea3zfDPKd6
zpLYsHx6jh/i7AQH+eQ9IouFRoGBYQG8le7YZmMZAuEU4pm54mfsgnPaDfEnGfx4
SGXuHTzcoCUVEPgfRNo4sQfSNJkUUHLVNZ/jcpw2pod0c/INU1djGmY4GHF0aKZu
IBDFYChZ/oZgrCBc2uJn5WfJyLmnChjscceZHE1Frqq31JSAejh1rLra7r52b9uB
3o68/7L2//MwsSF+SsReRWoDtoHGzzqGM2JHQzQ9kpDdsmbkzMEP2LQUgDEnVJnP
G6Mn+RmbFFWeUEXVktP7z9K/sxyHfiOysu4gZ08URCoFe+FovKvPTptRaiD9XDcA
t1fBYanFWhq0xEm8tUWWODxUJtETZqwkbLJpsTAsPHeSM8qhzxQYJzMt6pr50x/A
lIMVXz4531PRAbQ/711lWNXqyMuiA2vvo20kcVlTNUoPROd/nLtOY8XrE9LHGeKt
Pc6qpnT4MtolQzW7ZpgXkmamegkgJYAE8wnUogieGjsxO7rZtbWpp8IjJPcpVJEK
I4QvPPXpOxlnTi9/KG9a34oRALmfSr0mqwuO3VAGv/9g3i1SeK6z5Fks5u94rWVL
pZ4VhhRkttid/J7gGkScFqoCGypDJz+djMHgk/+QO2Adi7sV9gzV6QIROzbQ97es
lnMTh4c8UpZ2T0zbo9MCyZBIU9q99Oqcp2y5fY7t214O1lCR4B8/Qh1GF2s6xmIM
9TFjkSKrXt3Ku3zvtEmNhHT1VZxJ+UzSjKc8I4Ii4i4uQXTl0KJpf2UCNQwLGL80
pGijqs4GqiSxTkeb0DXfhc9Zn+zXKu79fQbQVlqcaE6SGVvxndXt1BAvrLDRbDyf
rc8Gi2xrW4eUAS02F8Pm4YzR4szdWQWKBHYfgBQIsRlYcikmwR7I96PO60g8RrVK
IAhKAKY+t//NNUMQOccnMIgawo6Qs2qLIGXvgQYfXpKy9BNG2h+z9YwVmBRQxdBN
GXg8JsoQHpN+sO/Wz6VBJfJ2MUd4jce2yLC4oEwLyDO2clbAWppRfka8izH0GDcP
jan0SwOleKCxMS04Qa7NrZAV0NSNd/hTIxsyxFY1lh+2S/loQfyD5dTNyJ1EvaCr
3VlV11JnlZ3pr2Pp6D6ncaGt9C54YId6/q4KsC3NK5NWmXP64X7m/u1CShl8VWxw
nAdRcFDQnV7YoZ0VCZ08DFBq/flJjXWep+Svs1xqdnP0WCwq8D1He2xr/+3xBox0
3bWEwRVdaoKWCAAoY1mP4xwhpdgF4pajiv+5apcItBV62/B6eBaopzRD3+MDwHap
YwpG1o5xDtXQM68yI2sWEDXWXLC0qtkSaPwlE1y7E7IEk0sZd+lipEUX+KPZ47+I
S5YrbMqCJSSF1o3kLIbW7HXq5gfW21prJAxTAZiK+gyytLC7GUfAoi3jLbKYm9R0
uLYi5KEkW3jYL32XFe5PEzF7EP+XaOqDCZoevYajeuh1EFeDPgmUDnCjPjDNHo1q
SHyBzHrbVLH5txel4mXBhYzqWxFnI1fHLEqnqpkH152nzQbYASldtnUSNItM0ldm
jkd/a6PVCJqZD30i1doBTKqhDZB8sMz01Cw2DB0HlYu3ftEBYxSfp+EUiEBE1K6N
k9iUvFOICy4vw956/HGKpfLyNg6/MnblLF0uEcGAuzlJ9i+h+Uk0+iaOw6Dwbcrs
ixp6gOF/fC+VEZSi9KfPBOHk3A8qswuGaeEIT7LegWQtZDFPX7xjVWDrl1/flxn0
b+BzaymX4peVT3akMc4BJrRJtSCmRub78/yrIeoDJBu6MpEm98OV0/3PmXpLLy57
N0VY5rQhgcloJet19+o2TEAUiKwdxgMvROKzX9IpYV3TAFmXU1koyvRDCvvYWV0Z
TBu3JkYheuEyOE5FAJN7j60dTQrKzPrOkN0fhoc97jfknLedh2DIyqbX2nC58pXi
4964h4yid69WemvJ6mig9bf6Zek2Fet6/isFvjto2IAPE/clB4hhfRqsPVoosnR7
nczZCCpLekYyMLtwpQJAgxjVtnHPcaINgj9lNOJBZhjwYIYmZM2RN7krB4Evv7s7
8ncSkHerFKvzn4lp3/kQJWP1t4Cw56PQUVeg/6NZm5psH646wP+V6ROMDuPZbLE4
jC3quxaJHTCk/O8tURjoxD0QDDVOTRMEKGoiJNb9UwhtMoYvCqQO9WEeTeGNj7XY
+Rx1Gbd14oYLneVOEoJNzyrNeZ3R1FzZWr65RuuD5zXjF8nJuIInTgd0TEZZCbZB
oxACMU5aLcEGJ+//oAbXShwg6Kj6nPsyAhnNhJsOAzsI9HLGg1IoB2CPyMI9vbTE
JM+JEPq4wia336LqITnB/1ko8lUbLsf3jgwB+3/wTyBEGG1AfyCTtnIcmRJ52Jnv
mvUEOGC+m5DvkNdd8h+47m4DVQlo95tP3LN2zMtxoX9L0zI1Kt04Zq4otohY3lMe
Z57Qm723XBnxkN98veDLHlyYetIHNOgLPhbiSkGz7pKQFSEAjpn7C87PRH30wBxq
WTHqoMy2FfsDc15C9p/XUk4LsrSTBRqPCqev5p74dKCNT8OZGVVj661w8FXbR+Vl
OyIZ1mwR5hO+utDE6Jzrkkzu9ScrghyEoA7cRENh4tOw7UcNQJWBhwFsDDdoNyZV
LFPzbGeLGwpiSnmM7A5pRiei/9uHfdHaMwlDM0DO3YMeAOZdB2v3hx6QpToOTsPk
70a2cNAAx9sgFp0T1sXOvBzVrfCq5DE69GJ0aQoYrF6YNjmAL5QsGBTXnlFKMNQJ
9UCilLrAGRPzzKzcxdSuIXhvacsZVfc4GRe9QLJs7gSwBH+3TJeaC3IuH6vAFaXl
n7f3E2ONh5oE2+unxujgA61c5tLuZ4bsUxbukoilfc+bNpgwHG4/hiWuE0WpsZ/6
L60yNU75S2cwlJdJarwLT+dRM49kOqAWVCKVN0TkgM/qwX+SBY6mFQddZZTgS0ur
hAwbVuH0ziEETy1OL0CiEqfay4i35AcDRcDENEh48tLGEw2yi3tjNG1b/K9hJ2rg
eEF/8SCQmGXt3z5Hxyr9avb3PFeUyJQBD1QCMRkZJA0600+riVsO69N6JsdtpRTK
pIPuBF4Y1uaRGPiErl/7ekEjW4DEBllWUb9Al+6sy7ld+GtFRyYr6cXYGxhWFg5F
pbefL+1zunV4fwphXgtbMpLirNZd2p5t2fxcMh2T0cuC2bywRvz9gaPMyZ3TaEBL
dU/jbqRvk8ZB8Cjel7UWPhFXzihoJzNOlsdUG15Qqkv+mG6jw2aqVWhnrt9nbSU/
kJbk0j86RRHm6vLUta5Bdei/jl/WOVfxmYRK5xS0CXIU0f68ncouXh8VV9mIcvij
SxVGcb1cCSLoMkunKyMXrprUGRuvT9vCEXoxIbolnHsStCcnsbEX1PvcnkO03ais
sV9x5aKbE1xu1aoky/EJjmps6FoVW6LI0/lN+ogXeVViS7msm5hK6pw/B6I1a6PM
N49169VpGmoqonVwLreplFXFJFCw75nLYCvq1psIDTLhLkoscAGNekvUBUdqhf8Z
d/+C3YyOAqhKq3VTPjE60XLunR0xcWd4VlZZHP46hv2niwaLFXCDF96DXBvoBgF4
xVfZkpVx5CDEdX5yC4ueIfPtuQYo37Lj3/aoTMbT7txc3SdRIdxvvzH4AKk4wmLB
bXdhvpkwLJxDHlfZNI6foq0oEF+xyFK0QcVZ1h1FwU3t1Z34uunZ7BEi4GmsfgHA
oYRx6Lsa5oFRGdMIHJEtbjT/mUTE6mandUotcoJjYROWYhIJDEBVhoLJjgU387ZB
qkFVa9IfLLLDEatcy+LM3WW24H0WRVaSQ1CA9yGa2e8oBdvt//Elg2tw6g3x/BET
IBm33+9AAnPbr4c4mPkzlINYbs8PKfZA6VVUHZ7RvAUZlcsexjlW5OgGNJnzk49k
JTTEM9K4IPrzoHUeD6kp2fnCNeF/32feIFlo/Pig4Mc53rfTA9NL93LFf27UVjZ/
+NKjDPobC07xULZLxSRyWWqq6NemV82uTPeXQpK6bLNL8jO+Bq3IckEpDa72ShLA
j64lfVQnDzE17vDRG+FkKSf9ctmTQt8WLtN24aJnUXiYV7qfBW6XI9cMM41bbeYu
3AON1OtjRYg91C/pwKKTia3MYAmetouJE/wvilmsU2oZNAjwtoyB3ZNSXVcFp9lq
3HCZvkV2c5WunesAyQGmuq4RpwMktl2Um2y7e1ooN2jhco4kQhD88JvfcCr6Twrx
nm0RhFaY9LFFUTRd673xwhgizmQfMCx8ra7Q1i5sn5r+IAFZuXNt/7t2VqnbY+Jj
JIVAiPYbieUeKeetiGVUA9BPxIZcKcy/SlznUBSFV7I5LhiDDpZ4JIkta5q4EE32
qssSCNexuRhpGud54a4kk+T9DzOcwN9TRQ32zcVPl+tdvKPFmLdIWqvFFKTMIIYP
27mCFkHlgXm5gPEz9HN/PsdXWvFpE5QKkKR8D+EhhSJMCiyuTDon+GHLUC8CzUNF
AAn6I8Ywc/cJhrYYDpi6rptV1uZZhuqtSfHKeRe5tfQRBm13YCtxhN977Uv7MDxc
AXpU6pCTUcCSrQC2XbvR3eJyvqBKp0YWOxD5vPRkW4eIOe/P1PDuDVVkhV76Hffs
ttmk00LeJd3Bao6/iBkapGocvbo3xlK5QYIi/4dBPGGm75ReJy4W9I9d8MH3NYOy
Hx1UOonZU1JXgUDG3vgT3hzkM457yBb5A2l0KTq23P/M94W0lQmEMGwMWBQ/B/vn
c6A6vgBzj/n8t87ZHZnw1995/YO/iM06QQRJbiKu4005s8gHW+dYptFQQkTtmkbT
hFBPL/T8DUjrzTUQNCUo6w34Nssc5jaLZhmEBVbfVVKwd4smhx/AG83HyZZE1ce/
nN93P9KLdDh80R14xvR/MZHyg6zOPwkCfpHZAmQx37Jd66LiROL2X1njHJw/SyeP
w3lVAgtRvMMNq+lbxUOenjSmxjpVn6OxkYAFeD4dLvUxBEXdetkbLSrEkOtCPzzN
1E0h8a/yEFCIVt4Oc7FKJURg5Cyh6i8i21IaWMvGa3Gq5UYIKo5ICAMk7DixLO0x
rhG0fENw1/LNpF7ZQ/Sd3UafZ5gx7NsgQy1VLVGGd+2VEN10StI9t+y3GwLPgm9x
XqORzVQTRJrr2r9Ilaa6biMZ+gCT47SgHFEtgg9rAK2Cs+juSypGNiF/DrmE+3BQ
NSq2JiKlPQPlLykz2oKnpi94Dj9tmRRatFMME33RMLGtYLJQIqndu1DNL1/OdkHD
6bYN8LpcZc1qaiazYDMe2PfaXP0Mmv07cnugFU6G8KO8sW0f3KKxTJ1ISn7myr2m
X3ewVBeLNQ6UaQ/Rga7DQOSjn/yotfQipg8iI9TEx2wCXDRL/QClGd7wX7rzAdZB
ba1cEC7l5+NBzLWzaU1BCCYTQMjUBwq0kodZWuqYZMmGv79ULIAwDavuzQAwP3b4
XaywDz+jtGz9jJflr+yCHKiWJ1tBtKW6GvxaU85O4FpcpW62R472QWNHuStUwCg4
pT6jZTlHoIzcP7cWmeOMAV+ZTVL/zPhwi8pIbOuVLH/SnmLjmzczddyxTWUJOCJ1
wcT5s/8NtSlIrIVIUW3l4CGspRqmiTG/ceXXq81g5VHUUUFrgexN2kTO+N9mZX9V
rBIiVSIMVNyuiDO0oNtWPkjF8XcZWtkE8G9Byz7VlmGQgQX7zOMfsCiKgAgQ8fvV
ZddBHdUxCKcuZn5Y2m/jLCn5h169v7EtWyBviOK7I5HXR+JgLY9E5n1QIZwAvzmR
pBjOj6kGjhbK5fFa3nG4fxNFRXA1WzMUMMzqB87T/Bu6ETIM+wV2jgCvwwb0CBDg
/dgs1cCNdgkT4iiwpI//U/bOsFlRQ4TqdzfqTp1A8nf0/mVltJK+eily5W/3MHjA
wcBRBUaQEeZb5SjLaPSmJAXKlsWOA+7qKmulax0ymBnC3dVHA7RH1KGBubRpZO0x
nlefEFay+LQyYXOjFLyUNhEZp1a9GbXRsK0Npxg3QyEf+g9zj2h6E3aOzKYMs0tI
klGQMQxB47wyspagm5dT1tucpvwX0lB8sJPiDCsyEG2KqNaiSgQdm7moz1OY1g69
/t6r/GpUv2tJwRKc33mz+YzIT3f3v5yBjZ9TRv8wdkTrrLe/s+1MX0LsOM/8ZECB
YDFBdvq9AUWCOfrEkSSbfKSvRcN33cAthh7a/JpDTRTyJmT82CiuUiYz8XkhUVue
ee4zjD05TvUBBVg7VtHw0iFS35tblfMDW2eViqsdNbo8wHQnLJX5oy60BXJumUfr
ex4xorrQAI8sW1n36srCMCFNaBfquynizLnD0Y4D1xk8GmMl5Ck/tfznfPRoU/q+
o4IvIxI2bz11yMIdpiydFcXEviiF9IAtKjnZ4RqteD6R/n1GPKxxq2QUHt17yzVd
U3guKgbPnBBNXFQ+6508SRiDy/Lg+UxqN+AM5vAVw2he95ItPGlRlOBE6Z/CUVQ1
wUlPgZT3EliClgS80JGOqrkWaqhW/oDESIe8ilXUAWwLueRqfnUq3na94Ot2FshV
lx3kZIqqiPa9r54KZxEr9u9ZUXrmSYXLmTNYotvr3v6BWz/D/XL5He+ZtiP4Kn2w
rTRx4XPlp7TFJV56avIH5J6rUh12CDUjP/V8nlIb/jY2IgySWBe+EaRf1nOC7cYT
x/sg07WCrflnefpKXj9ovpT5Q7jiTi9M7oUMRr0u9SLMekF4IwFuqO5veuNlbUTl
H5RyJYKZB08PprBcxXKzccYgEdcMTu8OBULAylrGxn5ni98xVT8merEKmZgz0/hL
m0Uqem4oudtcl258+w+jFVKABkFoPFjzaDQQCJgAFEYQ9zb3kDm3+AjNnTp3t7VK
+VUzdvWkG3f0JgnY+B5GaoqQzsh3QYjLP+7TCgDMXiq0hI/aFz2Vq5HhqGvc7UWy
o8V7Q7wM5ePnHERcELaCCqHNLlTnB6O6EdfLfHjmORRVWfpexZra/lZn8posQcqa
/F8bGZlHetN/AYnshYVZ7J6UZVhrSVcpGkkNcOCV09QDHI91nk238AZU13q5T+CC
FxOY5mKQuanH9e11TwLFUphDIlgSrOX8ZHeT+FlDJdeUPQfs3AapGHMsXcpAi8w4
mPZA3r5TAgrnr7c2LYbX3YJOitkDjJrD8SEQuxOTEP2ke5qwg8gejOjmKfq6ngDO
j7ezleplUUwRDyurWmXYBMKqEdwjGNHOqtiOV75QqoJgw1L5x1pK6GZjHS5boWNh
bslDPNG8BEJDMfICpl5QwJeYOpcV73B+rUaLTKc1kmyN0MJbULoXc8VFq0mKQW/w
oTLnyC+28tF4S4I1hLFTffzG9gRHzmD5uIRSLz3ZJlyD3HyH9vSC+1WMS4/JPXkw
g9ezamcLYPkSU8NiIMJKxsfnkef5l8mJwkO6aTjikQatlhFwEqYvS5ru96jr+uGB
4n825aBO5+qy42ihqAOEFwlFvpQVlaewqtlN73oxBtkjUe5qj5984CN4ZRuw43iN
yKYpAhP3y/OvWw2PEbJYQnMWukbkANjOQqN1S3No/6QL55KwIU4vHUE/85huzLfM
6T50m1q6iKyoD25WByyTmnGWNhDyxqC/fZZ1kLxmK8rT+uTRFOG5P6+7hKmPXeWA
eQ3Llvadu6bnT99Qp+Jo+Bux/ygFUEZN2i0vFREnftVHU4c/2BDHQyupT3Oh/mWw
PTAiiaZlkxE1zlk+z1sRxLtNjVpad5J1LN0mEPbZvSfmMXKvWXzjQ199VJOw0RUQ
tAljmtNKS9e3Hfn5vvDk6+S7SgZYw4Gcbn2niGhJ3Bi+tYebYWXxvyzuJ4gKEcbT
g8wEzEWYBCdbhQCAN9FIiysJiMg9rawx+ufWfFgtDSh5rSkgtCXr4iDhOE5J4WrH
MI6sG8oSNeWCLCe84zJo0TjPjfTj+3KhfB3cpzST1C92jd48QUjUScClI1RW+rXE
LgkywDr1xLXGfarZI+o845NKh3yct65xP5v3UTkOztpT/2LpAEBXK6r1uYe4/C2m
oqBWT8ka/rDJztq1bnaTYnu373zKNMA+3a1Ch8F5VHVEYtSjC3wA8NCGLr3P/Tbr
ssdZjfpOfUluUbRtIjAmFzxlNIvW4dL0F+4El6UdnAlQMKcRv2qdLCgERVyvVpR7
iYYlmcuAUxvxnoUlCA6Az2/SAVP+V1vIFw+LoQazcpXuiAVM7oAvQ8xUcEc6dcYB
0HbuQsEjhoyJ9CvcFWsyPdTX5dKcZWSpMiLEor6qOD0mMGOcr3WsP5wdGgON1V5s
JBt3iJiKFF1AuFWoSfTXI8guWrEqmSFIvLK9xP3cSz1yVliSvZ1OGWhg8z+QI0n3
Vq8yNa8hOAP5XlXRLheE3JrhxN7ganys2H0mCuR9uk1S4w2ewnRJGj4Je84TLBi4
0d3T114LszIV7NwvZazFcWQvhPNKS33Br6jODnmAi0GezAPL4Ru+rNKJXFJ80tYy
2LO6DRAtBUbAl41qR5syepbHACSvyi713lXZeTHO4xOfJJRQpTHDTU754kI7P4U8
36RkNVLA3VxSB0fIyndgRiqXG7SAyIPwQphnzkSPm4qQDTVQMxYCcuIInXh4yln1
yXzwGnA/S/4ZTFc5GuRqFyZLcWs0pWyiVYNbHEGbwQvD5bK6Fp85mToNO+PIOsyh
+cNI3E/QDEIeuTV9a8l5giM5nqyY20SmJGTNzVTciVC0fRtFJtnNtHhW2jjbzKeH
EqqYZRccUrTQsLuynDxA7wRPhBN8eYLmKjJEWrefPsHYolJZEBVLFVWXhrs9plmk
3SiTXYqXd45Cm1GpffzkfODAk4XxjBwA9iaLjBGWzb1LSi2LXxTzQ/ZTxfREZ+Rr
S+3ltcnvsI9qbbblXWWMKe7a7sQH8f1JWIUzf8nsel9kXHFzE8iLnpmAHA06285m
hIYtRfqKI+JDYodbe7zzQwr+gDMsAJ1nJw0x4P/qLkqZReuiC/En3Kwj6TyCYLB7
XKFNDbGJbtk15BhLef+3VLLIT2zokOujXbbSPZOQyxN5ArVB09r1dlIHV6KMl/cr
YOi41AwYTH6Q1s4tv1ipyTy2Fq8b6t1QkBmR1r/wLxju1muwmMdbt+7m5j4F/FY9
FOqHz47hNRuuStedOtSDk/1lBKTJUw+cjFGwYbsSpWj3STPS+hlV+3a3YsRaVhFW
krbYbmMwsmmQqGQtGtEGmucmnMVVT6PbuswZRIjJ3XQgu/oV1V7AFrPqcY7ZJ5J/
ijT4bIJCSYrp0BRO6UcgJ0tGCObjh11WtRnuwHLc0UdFqAbKghkIYAUXZVlxlDzc
BZcGPc4oc3fwI08EmF9vXhWFy04iT6+owpvkd4AoybJsWZMxCviDgzVCiBEglRNX
GWy0/dB/mokGhWYOhwVtOwnbUpkMR/RdBg2V+kYqSk3dhC7yfEaSpCvwfywYbeZi
poy/w9mIsyUKq24rxHTDguA+aLgfCtZwc1uDW4EWEjopWA7CRu0COG+jTTSM0YUg
7ftlksI19p/L2XOmvhoTzNJZl0XpXBt9fK06LslkomYJ9LEUDMO90YcLJsNsN+zJ
tAwVNInLxelCQZRgWIjtFy8kxlV5CZnFj4owMjESdtVXo+6VYXG6NWz+0HvDGFVY
hT91r9kiT78IWCf6/LPfmfTQwkHOAc61Y4t2htQsW4SOC5Mk/j+uDnygr9yPDq+9
37vUMjcgaAylrMDZ4X6Hxx2uYcLm/VqJIe2o/LIJHh9xbyOpyQgVzrnKS3yvj7EU
vLaZ+76fMjlEBsGjx8JgnVqcjuih0KBRXyNRSQhDYB//pLCfSkN523YgLfPGm36L
OkOAXrIOKJ6L5hGF8TBXNyHgZ2ah0iw+Lcz+2b3y4uzUYqGBTlExdDaBAAvSJIt5
JXxKAvuW86laTx++FWj+TMuJCsdmOyr3ApdLwS1jIGjqxz+znAK8Yh3G9RS7iHR0
30ZvR8+MHJB+6aPUHw5bViMbiJFsNwJ+kspy9OaIot5e3iBG1yp7MkzC3IJRp5FQ
XKy7amiu3M1O3LEriywfu2eGqGIop6LB/lRXKEmCyO+jtpIy41MPOXbbFIn3w11f
Z2Fo2digizbhOQCQEEHrrszWqp+GzRnMU0+vaFzyaqNv8+rsGI1acBcX0p/DLzXz
hZET/Cv5ALfJ0smQai8Hz4EV/IQZp5L1KdUH1TOqrw3UaMW/0oFzDqcfq4obv7pw
ebC4aytkrLKqBzY/01TDkRrZ2wLE0YRMVAM/MhoVX2vAlT8El4sRDO1cfJ5DZ0Rz
5D/k/ZiF84ubZHA1nTh4Ba/8Y9mKT5zJQQIZ7FTvgMn5c7okhhQxqlb5GVT7uplP
pNC5T5HhMfilW/9cCO9G/PX7RNOnuNCLKqpkDUSOYnVGCn4kq5w/yMmxmj7+nDZ3
/q32uE30KKyivQ6iLtaduI7FceQIlboxggpUaJ1TF3Z6t6bfXh1VlvScBMGibPZ3
gtvkApF54NSHVb2u72+KRoMFpFVpPu78DFPBiVSiEyEnzv9iTYx8Ry59rdHcd4Md
TeyFkOzSI5oGwh+1GMN9lTBeNY1KuBGV0ztm9HPKa1Oa1AvL/rIFjFuOEBBtNCX7
7nftwkVpTcDZmMyG4Q7oRGeViXrOlWvup69WWGUyKizY23/MZLvrK2M1AWq1VOxR
ioy9QDxDmsYb5s8dMxujkXR7/jvRScVBPhyUQrdIqd/OLsmSehjAtozk+WvXkBgL
Q2EwbGfw/FdbZWdW+uNaQ/eoYXCwT2zImR07fi/njTgfbNXiwUXja0FyqPYhwcN+
JiAVdUm2hYQaNpboZYukwQlWtC3vh+nMmVyGGJsXP2hKZHotYuSGURYUqKpLeCVk
NcZp5Jizr0UjIg7Keu2vR5aEz4Ry6yFTpsxJqT0G08wTjbKF/zQwA1tIX9PimExa
7itBZf0dTMOJCcCtvrgMoAbthbA8swjzUUZlA7b/ZwVVRbWu1dcEOJbIqDCVkRK6
KTaMKm0OfJbfmZ4EH9xEfrimcpuVDGmB9IVbUHrk/Cq0rGXScBa15wUUx8BxoHp5
NLLZ3qNuFqHmDMFuvOasfAJiBjheeRxgRctUy8TRxJ7mnqU/OHDCO4oQSW3b1Ugt
aFaGwrfEaXmRLSlDeYc1ixiSqTDJcXBgNwUVcqdbZHcwHLdHVPc7/jfG5DZ/FLsu
QS99x6yeQIg+wlZ5wp55ztN59mjrq6bZR8xzr4tuWzkbzr08DwNd6h7Vwi3OoV1X
uA7VqgLnw48WZR3Z3mw8WzeqrsCUj1OUYuq6wF94mqdv10hSfdk0+sBF9u0+Ga+Z
LMt39kY6kA+uhA26UORZlRMCJlC7MkeMskhMfMOxBXsIhdggxoV97ikECfHS4ENK
a++JLTPAZeQzwKx7serk+GK4Tx5m2FYtphZQ8WV/KPoyxy+SwzWoZw/cCy9AVplU
vQGUl9nCcp3Kax1XCYHHEudXIgc+UQB27zSi2PoHCR9UDsyWUCSAsDez8FGF+sna
SZVbXkgvavdEPt+5FV0nHAnd13sc+XXrUYfqkiXk03FsUzrmvurENFqRQfRH+6qg
1NE10gSo1Krt3p7V/3BScFXalvGYFd8HchQyKYa3lrhbT9Uwu79O8ivolTD/wmiw
fAcmlPQR0byjN4XEam9N82308NnWqZdrSrDnjZMXa+nNMVJblwCMCs0vCo9O7dfc
gVMhs+aAV3DGOmUYq/tHZ9r5u0hE4FYTM/syaPJULyQubAb8GelalK8aN29pf4MI
cW799E9LiUOq47yh4CKAP46+sc9ZP8dH0aV3Y9WSZU4xuyF6rtNTPvkNE4inGKSR
JQ7x4Aty1/3gxVgwsosltZOqPm1uhWtdNgz1uABHGHWXjvh8JIoWB3RPbB3REFEN
z4KZU8lxP6V1EbjjT+o3dPI5Y1jGlEUMBD09Hl70OUBbz5Cssf1NOMlW5zPayhBN
SWQ9oiDRA29jL19g4Ut1w2212muHr1lMB6F6CrUNnlBTPUjeACFYdFxlTL8JH2wE
Lp6ysOvslJCg2Q1tMQ/h0WKaU9U4ToH+n4lBUwdC0jAPAtDavSd0gX3gfqewbtWT
oARYfvEzQpsK8fLG13qknFpZWQPFbLyXHj8PQhuk7eMbfyCQpTNGfACLG6jns2w4
9fAONz9658OYMHPgtJYNThYWBr3oGYoB6uSarA2srhlnDrFmFN+k07JokEJpMeoo
mC13XqqIxSE2NzyLwO4hb5hlHQ4P3EcZNhsvBbCsaxi/0sV9g95t4XnRFX3+fajR
qzCmlCXM58RqL8hQARfhJoxT+abDXzk8mABIRMuphScMbG/hoGTkrA/9CRvD3YDM
k6p77TTfKCVb4zf0XwE3RlONJiFurUjtJfk6bB1t4eAuOA9nduatGC2DkpGHAJs2
SdP5x8JEGnZlmmsUsfc+VWlG4Uh8ehEq7RVuvMIjUYe4N8xPQt0KGBWPLpxieHLu
xTOZKnOND5INR+lJSi3TWS+shrsppLg/G5TNgZAPL2I2ecyfkXynse/Z5gnt7Se7
Q/FEVpASYupUfSQM5dl8W6OIwlkWvkJdLOLWZiyeztEgImxeVHu4mQ1FrVz+/qzq
g+VW7rIn44Sj6gAGvC36Z42DHB1yztFVv0LOFwvgc4rtNk/FMfDq+VsYzunntbE4
A6ltHaBLOEevG3g7LVmyHXUsfzc127YZ60nnLBn8TcSnx3TyP3Aj23u036miGEMm
sZkzbBOTiUtxSAvCNTgsnvVNdraKmOonCqixV91s0ax/BVTkyWqAolW1cIvGrkJR
y5uXBE8gc80DtZtkeZgzWIPFaC054DgGAHzcY3BLccTWKJn7ilBx+KyOET/Gc0Qu
3zYDViKl8hWDk0zCL2jVX92my2RRWZfuD99E6P8Be3I2bJMI/NJM573ZJHXuec78
Q0R4gBRrIcVj9/wBW2ewJ5ijGPq5/QyGfM+z1d7C7uiKSatvbifOwLRw5jwXnFBO
hVoCiNvUKmX4b0oG53vO6GMphPg046ijehAT3UWwlqjxnsmJiMltL7b7nFhCp8mT
wX3etO0o+w6Xwb+SxZwVy63d7sWY5ndA3oca8hC6qDRRyA/PMtiV3/nC/VehsEmh
gS/3I8UI5lqOjIAO9M6Kc6j6VMJ7BxoEZOpqKxrTvzMkEENr0L7BnlAhIHjphIAd
3oVFr+dwqE9RHGhj+D2n5qq6sUtFy8NoVJWVyf29MSko3N5J7S1AVSPcDxJLdSxk
+1EfUlUjJCy8AKoRiuy3lMJMbcicgm3oONeZ9XhjjXKR/urVCfwKLoTczIE2Vlru
lyNlIYgP8O9wUk/ngrZeSazzpw4AuDUxaFcmmvE6Ccc8C7za0cG+LGZSSkkbhfY2
fr1MKeKYNpqelvVjP+zyKpSF+K06J4JMduCW3qwcjB+5AtUp2njipowqjX6cHMmS
cSvz9guwwR/zwpKQGnlJqJBbOWsSgSHKbiQlVStVRP82BBM4DvQVodNME7CacEve
YSIaeMSDWDmZuCDfvmyObcodpPUosqOp4dstvtiEg8zMmB7wBrEiVfle4wF4fhRt
UUrMCJzlcUi0zLfczjBzfxeaKGIC1ayAP5/wWlfCAb1NGhV7BP8M/NpdI5bTBedQ
Ry30lGRRpZ7ZBneV0wHN6YFvw7nWLcTEsln1NqZTga9BL73C3f5fv/bZ2Lu8WiwR
i6NvVMbTakr1aEbPC5OYm1SQ82QqVaL4J4XBRVKbCnUpSP5ymPiamc+RKD8s8jA6
VCd9+hKZshKDsopP3N5EoLq+cq7Pc9hyM27p/fdO4cHnyE2rlrehqdeWWYIS/wbr
DqvBzwoMgDeIe8CO1rkP7NYZKiMsM+3tOlVpjqwmLhypsZedoDWbzr4+qvsUnrTX
GCZkvaiKZ2MTw2SHeE2buGaiYwItSl5rMiGrMwEqkV2FoDNEza2ivVQrQaoshxgi
yNCzffI6LqauwqJNvzhg3DIvkfbY2ggb8bdJ5YrV7XzSZWmfzPKCLS6VNIhYdgVH
db1D7dHXSKUK1Eh+2H3YmGFEupG6AyUT/Bfg4ze++9V68THKPwaEpjJ/viAkBVzg
/Xh4sIyNmvuFS03F52zYfhOXmXkC1hnm/KVPdhOURdFNOV3GXz4almMPsK9F6vIp
OC2ahCRt0r3SUcBfUwMDgLWjdEiiG28655NwdBzFcL+yzJKx1BNivCX9dPRlp7zK
2cE6MfVzkuz8xaR14dBa+Kl02Yuzs1M9FEMOnRu/btJTVEWMa+qgNSTFicylblXw
ev+wjRxLVjJ2999x78hVnhuFqxKvXk7XEpnnkSpZBakZBKLTFwYn0zGEck2XEYCE
lPpNZTEWgyCkzkDWAo7oa7Ri66r5AhEEs+SwTmY7m5Wk2IhyypXwaD6/QhTKZYbf
1erqzBe+Yadh9LV8qEmhaStbor5sxOiDS79tb7COOFOmx1bxLC9/bBM30TOcZh5b
zbQ1dsERUw+k7yuX+uRBoIRSehBuFC+pA5v568++N343CKgs8dsWyUENRN0ZAT1M
6+QppF1mjQ8q2d94zfE81Mmf/UiTWME6ASBLVEyh8k1HTsbw16vVk8eG74igNweO
kIpVdFntZsPlDhGlhGLbxRIOeU79qJvfMNHpKlq0nBJ9w6JkR8R2vI/KC3OnL3Cr
JT2xoowjHn1eZtr/Xo8XvF+jx7wz18uWChUjrMfQGzI4Arv2TpyJTghn3nAVFIWX
9rOPb5L/A3ddyVMGe1NrCdWvKT43sE9LajI6cIbwqOl2Smm7Ow7a4YE+IKJxoK8K
vrHAeRvq40Mu3rwpQIttmMlZH5/FEOJGIpMqX8s4rSx8+77mGzSTN4u5313mX6kq
TD43AWXFEeRw5xdWAJOhWTgc8x7BpR1oy1CPE6tJVRlrVr/Y+em9ny4v2gAlF+Q2
z2gi1tOXzwfDrn8ciJM02nDn56DzLI9x2IF4ZMJoPo6wJHwxalixFHYHk+LpuSXE
vrxekKdSfpyZSEO5EDMGHdmPzYaiC6sSp6pKghl13NauJ2axIWRCJH+qut/lJtiF
iCtA1Tc0HDL/su9Xqva9I4pN1Mi0oEayPPBDlBMMUhLI7BzZOExFjeO9co9C77Pj
+8YMwPbkmWCkvxaPiZTVquMjkIWTZR8QHu3MTxIi3NzbDYA+eu0l7MeCKCXj3ay/
Mtrf6z4kw9vMsize/wBYoDvLR8OF2eveJdEEG7ef551K65MVuCx8bkCQ1gPoFwBp
aDxw4ZoBWm2NNfHaZtrEiR7Y4UwdR3YpKJkdAjk0kLMFEjyfXJeWVJmA9l3+hle5
d8HzkJK8kf5BgMXxeTVQL4o3x2M0wkT8MKfTJJaDkluTi7l+YBUSzKnPBZhtQz8f
w0n3hpd+kRUtuOLHrzcRwCRiKtq+nlEPx5nqiCz2bc/ZtJT1vSJBwMTgZhsoEjXn
Rbo9pDeuaQMvVecd5RvCkwGd5T8pbRBh8Xz/LSYJdjakxRG8Pu4nc1xcmdmjSjv6
dr8/LthoE13bEH0D/rhKpfiJO1l3nqmdsMCYFCbRhqpFWetQxs+4QCr76EnzIXqU
C/U+jv+BzG6DkZe9TTDplXNfE4Fyi+ty5aJkf9MB0evycm77DHswEx7DGNHaQ4/2
eIZo7uAxf3bGerOE+wJ+SqahVTufOzPWxUsRu1cPIWHjLLsamslO4qIVMZq1iHOT
n4s7eeyWN9Xosx7BEy7yzhrNBCeMFeYUuBQ6PH9tdj76fr96W7ll/oqVKqY0t34q
GCOvw1P8QK7aDyLB+wE7TllReZDfNKiQuv6bW4pltzZqL8a75QyAz2mwhnDP6u5p
VjjXcGMN07Rn0Ot1gja5Y9v9myyjz5B4JjsLpxVt8qA9VuFHDInl2ha4tskCGcKa
pat+vl7mL8ESDZqKz5CZVISGcB8EnJc3qSLdoMB2tpMYSbVI8sqkMNOeE9308jtl
e6D9AvA3uSufG80HuWW5HQo5PaaxOuNcUpbEUaBZykRurEmslVJj9oJZ8rU7kv+f
TAq6MZ6nsy3/1D5sT1wRPVUXV7W2RylxuapB75hUYDeE23oUJ8lo/0oyNfZ5uaZ+
pnZSpp54nIZgbK5koUednU0Y93Sk81Vkfdm08nZxykXLRYV2NkReao9wXnFhktkX
UPmpTP929FFQmg/tRlgLLxWVlSybv8UfJgiyBDcWwT7TrowElv9D9TrxWQiS+Omt
SA4fJzVJJ2abnucmnQNcdkqwP9CbkY7VYmiX5nYkEfDECFsuiBPb8Ndqtt1ipphI
T0DTfExYOW5Si1f/0mldCZJwXXMekb4lJUqFzOs1cB1XRyb5ZmbBsPd6ABnqFMzD
lQkWzyW+tlsCpKz5LqnNk/QAr1rYO94SjTbLTzkr4JKxip01jm/eKfCXJYFKAPyF
NVo2ZYb9J4DtZJkm16E8w4R13IXItAGXSvdPktBqE+77Cxc8HAtO6rtbprzbVwCg
IxPAKJndjV+YRgw3+jBgLXATNJ1Qzv2I1RLxRNk7Lt0g0mPotjn3qiuujV3cjw4e
a0WKtJAyjxmA8t4IPhdqVpZlXFcENxlIFTqDWrmlun8zkxVjKRiQe/kLZj9EmKqr
rLkLr9Hs8aX88fzF4FFDnp8B4N/kazJVnhyeEL17l4ZyJcgd6Qr509+rvVz2G/FH
h5Q5YHy1OqWNKyhFJ0CSDaI6Z81yAM8t07G6N7JpYIYUO192R/viOc7RqUmkt54/
BNKWuTHERrbAE4vikwzazMWlAYkVV0WT9kCXajl1vh3yZnVUloSTS2tboO/kqMRy
5kyyyjSnH48N+i6o4Hthd84DF0/OvUiTebKgih6vU9IonZpkjUu204AF7/kpKAOF
+m/GhW/cAG66iJIaVaJVIl3+zJgMEdsiyas9FZFA6bm+sBaDhNHm0kylkXgFuVIb
gySk1bvtjdYyUbmOfKUGL2lqv8UsFO8h2X8WQ60kTK3Oi0i3tJGnZJcQFoHHWyrS
EY/ixG9mCohDQ7Fh6qPjQRQSdMBIPat7eias9LlwG7L3aiyGJUJuvAc78ZSn7nwy
TCY9JQ3H5poEPmpVwk8AC7SOHrMiCbczMKZhHiEE5w2z0e4Jtrdf/1B1PfnDUgcp
T9wjC+fpUQm9muvT4CVcwL2MO9CMo0AQaPtTUUmUPIBFpUotcl3ivzn5VF8UK/yH
MO2Pek0MhihwNyEuZODLdLkXPYzdi35L+/8swmMIREYs7hlNOPC6eVos2newPpjm
rev6a8FfeWSxe3ioLNbUhMk2cfsMST1vJ0Bq4fJnweCTsL0AGKdz93yTxYtcSuJa
MR6OnB6D5xpb1yqMq5sqpU0rcLSyzxKUPUCaQglBmSbcfPUoOSJHk4QZxdmkT8IV
RTMG+8QoNTkq5O9fg+KyI5QgKLGIpb/Yjn4o/2XyEi14Dvu8xtWSz7vT07J71gD2
1+cqzr1jhJYuDHyYKGSpVTNOBL5wb7W73/I3oy1C5zhQeMdswU2jQQZHy8KD1Upu
g2c/EgzO3I618U6IIhUKZcnMc693uzLDKgYwDwPXPiMY3qV7PHhllye2DqxDIiMA
6F2RtqefcFmwmz0CMSagG/gjoVT1d0GmTGI6G11tc1jxkKuuddWXS6RnHEqlEYeZ
1LCNitUwM/ZKxFTYXcBriUAAuTUONkUS+kvyoAmKLiXiKC/inQASjxzr+G1Q3/9b
BylZQXYwGCou5IxVHFWl15A1WJ1bvRickSS5ROrMgLOsLkHdK+/ZZceq15G25r1W
kB3RSo5wdUevNZCfaqSMZEGWbBh4pxgcJ0moMBHse7qHd/LYm5eJTm+1yiq7Ntkd
oOE83EvHX4ddevUDjYtCIQyW017QrIMtCX3FkvkgaelLrA5jgG3PrB947sJk8q1Z
cwohro9fW8PwTgPNjQ94eMwNAJVrIOhJnCoczmqO8VV8chGWx3091L+g9vwOjOfG
deSC0LcKcfC31dgzGAzGWqb50p4gIvDBmc6zro3NagHCY2u3VT1i1Eq9xIlH9tNQ
8C+RWrIsOoe4Xta/jN1WWkWX8cQe3+nYRN5GXSl/xyfQOHn3TbcFBocqfuC/qj+S
yuKEOACd+xPp2OXgz8FAh7/tFynLMwPv4SUsR+m8aP3Icht5fzPWLy7/hNjrpUUC
TJJ27UnVcrmQf3OKFitvwaPrrm4g4v0beAbct9NRwQCuDQ4ZqXnvYfyBZkP4Ke87
hBqj8hDrb2dHCzKAMIozIF/5H/vIDBb5nYAjOu0vJUTbIEAQhbkqEqfO8b/aVzRO
F+FvaVHLhz/kAba0asNRh27U7IVV/JiDSeL4DMBFl4aaHmGV3KnIJQDSAD7IVl6O
XNp3Pb/JkllBxK5WCf0XUhIsAGudeYPVdvOtSsfcSEYxTCHN9SeUy+RPQq5JUF/X
q32auDju/jSwH9QR0dk9JIPFg2E87lXWROPht0WrCvxFp2fJ4vllpnsGBGpdCaSf
EpVktRRZI8Ue8GOg4LvCtcyyenek3Aay0Y3G18N1YHtYRH/v3huDwccCfvYDRwns
kwlEDI+dddyIPAQtxzwOocPSD5W1VTku/ytLdVkFMQX696v827sxhavUnwZAj3Ji
Xj2LnDAPVCcKBLCqNf+Y3YAzcltVD0uY0uroXOp6dTRaoUK4ytxDz4r2ZUKb06JB
TXY6ncKqmizPnwcLXuZ9cJo4YUXqbo9cTfnx+Z1ffHrEIpPU3Ev3TtDsZOGlq1BX
20bN45tTUMPA+2nllOFl2jqBA9WCVCgD4lxYx80HKkVGXwTlXf9LXDWuM14deGp6
/d8086man5QWqthKyn67BU3KmJq743TaYuzfsKa1giIs580OfVX6/+KqNh0L0PRg
6eLILEMR1G/5Tuudg00lg57euWkcF0Anr7E74RXFZPKtiXVSG2R5VIF2tJqQXI6r
1WqeQZ6bbsZMYSOXsI+TBOcgZ8a8v+rzGYMz/Mejguo13b33ho8dq/B7DdV+4p1x
+MOXT/gGRswrwyX8/SmxLwzPsbbOemTYvMu7/e73RLFpP9of5fnRPNCgpO6T9tP+
pckVd6VAVLhmbenlePfCIvD9ZM0OdkkO9RYbuQwNbglxN4evYSIADSAe3K00eUBG
Sgj45xcsgmZks5a4n1gOs9pv3V3pDwpuagOHDQevBBdsEyFYh59vdlXPowTIF0V1
If0IjfTtwltC4t92FX9n5YQ4OQocOOkGcnF4u3s957YswUj4VyFJB1WAOO9+u1Yc
7qUwlzXTfGj8JSZSQw/s62hRY9rgIbKjjdlNzu8zyzNqEq5WYRkulcYyGswV4qTE
EedJ6gvExisgMQtlrs/t8QkdtdhDFb1qKpX4tXwY2DLq+9Ceptv3lA5X2JwvC76T
dyuLXyiRKv9UG/heSVWcSEszPIGAP0miekF7+Tzfx+EKizFvaotzmYEzbPmYLv+L
5nor4nmFgQjKRcVBbZaPDYXFnCA9VvgEDvcJ2ClVkBM26kbX+wPlkR8F8zk65Doz
JLy5Qo+/cRK+MtdfnVcm0WKGM7uXSp18U0XdjTJ1aAdqrMGw91uxzzYR/OUuuKO2
c/ZRTMV/rgjslQSP4stOFsrradtw9PUfe6jS5QDZJfOylJxi8W2aTd3O+YEGQ4yx
fvA+/0xbTkeCGk0tw9WsEgYRGeh3UsclJOVnXNFASPT+Wv6jjBgSxN0zaKQgmp5C
1w1Sm3LFrifj1nMZfk5tsLopIWr7PeWq0oRIXv0POPNfi7EjQZfPN+Vaw6PkMekD
vfFdEQqiIHAcEa5H1PtFLBAUZD9ynB3PZqzDrrPmePcjICOHhHwr4FvwVuonuyCe
ucraG4MlTGHzS1Nok0YErUgmTJSilXhF/fIZMSWXED4LFK1H2Uv2m9Y0ag3gMmdb
TsygXsLW2yLrE8H7oE0YpULJeavui3sA6/fNRbv5BuUeRW87NuV3demSJFNkNCf4
QW8AwujENvKz3ktrmSmnBJYL5igf5UaJn/48Z8ZyZeempuenYy7/ECzxYGXELzDg
aX/8yWw8hiLs/XuBCx22n4BgdJTGjxe8GEoPy4l8YEdA9D0DDoWl58GetPhkqMhK
fR4F4qAYyOPMLe5D2C/Dur3MYgP5UoeglOV3gsrIxtHdOla0FW90toeItlzrZfFF
tY9XXZ2ofijlZ74wsLTaAt0dpeyf+kZOUAHI/uy2q3iFsXPUMcq4IplADhft0p+z
1Akjvc5G8F6O8UYHI6SG+AkFSubRF18SpzUWoX63gCiiveF8FHOtkpcX8Mry6cCk
iMu/xmY7jACgmjLXegl7wlBJJ2F+U85bLdx34/qWukSnzi2869rU+VqDHwklqzUH
WkbUvyLetb9zF/ecHOUlH/tZSKmMlro6jbWCNHxRAJK1ynKbThrXZ9r2ju5iaE0K
obR8MYuGq9MLSCIakTx79wS6iEH3LXxa07TUCSQswkZ3kuG2moYwIBKHJkxh4iI7
uc0VTJGy8dpW+UxnAQwurPDrlPrw0T4uyqbjIurRo3+zRud1fwJMDfFWZeHCExQw
jiZE+B+19L/MZj0B+9vWfoSYr19DET6bLrFtLHmTQ6yFrVx+mpX7XARFq2DTcQCQ
ipU3g7jSDZYi2l+rM2WSESkLcCdzzMNcrF1oBnCOtu/CvHzjaiBb4F6LAXSe2PfW
x491i+wtO31qe4YmK+I25RcAEL7NS11b+nO3uZgCPYq73pu1Kj8+Jd2kjATrD5kB
N4/wnIiMBWJMZAgp1ZxUVRBwrjSV9NC8dB3BO0NIUCC1sTdtBOJYeXuZUWS1aPKM
CG9XWCVmUkioImZCELd9Ht2JxEQbD9pkmJj99kz8PHp1zy5TxjJ4ezKE8P/13y1y
/YGAFB7jUFhsg2Ee/RsDl1JVcu1RcxQNXYGdfY7YgdasjhYB2u7uz6/VJN/vdKEz
H0GQLqMmULf2eB+OEJllkOCT09GT+jamb3rReCNrBGvwLQZEUo6O3LfnwKKU1im0
38bIQWVeMV6j67B1868ulML6F5EA2AvaFxdnS9A069CfGFA5lm76qKQdP6XxNpzE
K7LSFPO/2tmjq8qaxBnwv1LT9UCDAMUmfXGP/R7RyprVjDmcGPKDbB3AzvdN5UNl
vGZEq9rIXcy8HiMsEAZfcJe5wuXbuBKUObeDBz62VIk4lfTmamCNmq2aOpn4wabV
5NAUdp7GyPu6oXX2prpOZKJBMDpcrYJrRcyOPQ5LCEojx/cpqGwvrcD8w6nFRE2X
jPnYDhZntmsO0f+wmB+qQH2rtoH74Nd9r/ndfTiDzer+vxWxydcpb7xyG2VXVlHN
r0GmmLsngfAJqNtNdhs3IOIPYdnhyutDZ54Z4NsE7D14UUZZpG2IvkR7AB9iZWuk
X1VHIH0+P+64HpZB9g62HY4qOIBf1bXMTS/R4OykCcxd2h7RlENklHI/EGXqTXSv
XYCCto58Y6OQNfN4ycv/b5/MorMVTYkIyajM4u4mLih7tDhFsiiPe6gmAf6Yj7ab
yNCJJu5HB45MroUnctobztuI/A2fACN6pbBuQOAy1IDITJhomOgOu/8gsh5JIxb+
2GdbtLcIVsNeyCgxGgEWeQksJI+2z38KA81mGPcngJw/cvLRVNYFJ8qvY1mWPxlY
ZJdOWQGB9ENLgw7aNAIImJ2fPuY3xkSZEF2+vvoQ7NPLIkzY/AguEOoFyw3Z4Py/
vagXVMLDPPNyr+bNxDiqrwaog/lGKqjrHbyWaQ3FGC/5Ez9NhZVkzijry8c5zguG
0EzfW6iNIRCa021FzcXbUxgj1BqMKofendKBZ7AARCeg04CaX0SEPY0PL/aGfpXT
ipIZlF+OdkfaO2358bDdUsYs7nmuzvA7YRsTMHPn7GqYyHTEyU/rzqiz5roX8Atj
yVpPYJIrimHv8hlvYqMzJQxL7lqN4xYdg9CfEDhCXPCuBKoWZH+ooAppmGNS0AXW
khWJe2sPpL8afFwYn7+fqAVmEbx7DB4B+3Mj9UvqmduU09mbwvu4WB3jQM9ycBX9
0Zj720BUp9P8awG+BusgLMVNcVTOh8KxKzYWvrdTI/C5pgIGeEg4pSvLfbw0AZ9c
n+E+R70OBdoWE/gTptkD933fXOKAbt3GgbmBnClTn9R4tjxcsh8huGG2cWH+ZloX
EpDQbtM8CeT8OW5u1ZzU2xo2atM9BRMyNi4xY0fMDSeZO4QhayPdU4s4msUE/rCC
WcU3vFKDh4F1+vxgGkS7Nw7ZP1IrK244sWPRIbbGhlJh1RM52kHtzMTcZIs3i6Zd
s1zuacRwT9EGrSzVtp1LzZO1U0XHYptudbjj2eo7eRBmkKAuGxycERTYXh0sBJN8
A9zrq1ltCvd+84XtYVmw1+sqFNdMzSJuOPQ+ugw9lZbFj5zUGn39A1A1/QmPnce4
z5NZCFpHAT2wMNGfmp06M4AtDxqKVRJOzgqRZ+EjdTTipP+dLhznEqQbk3yLbcoh
K9tKOkWtgqVvmi5v7qG1TlzO6NJdsWo8Nqpm7wyvKsiGGCT/onRP6Poz/cSnpuqQ
r3zeWtdrGCBzt8aeIUYRZRxyyHBD73tFT7WSuWtGyme3O3Qho942M2HZHsyUKoJN
oyd6xy0rBnDLm9VrX83pzHdSyk8bsVoyzG7jEexhm4e7r3j3ah3cqJjL2WKl/5X8
D484zMaPvX5kC+y9rBAeNB7lboUOhLOECCilQTFMIbQOvH+UGzMJXE8jpzTyYISN
UkAskNIHUwoWgQ99iROdJ1EkehVrij0zWKwYjHoo0DXFaFGcvPwQlMLONcD3yT6D
Pyf5MOCU9NUtNrjtP+eC2eQhKV+aAzWoSB2mbcdxjXY+JzBCWK4/kTr6ZEWfEHwZ
rN27GT4pVQ23bUlSKpECpYn+97ssj9AF9cddk2gcNZL8xzeyVCIUmx50qZaWGTPm
QW/5Qtaz27kOO6X/Epzs3NhBbclxi/8DkjEQ5l2okou92wXSIqJgWyF3wpvE++2P
Fo/0v2noV7ZOJSy0JsFYJ4bE40RTVu6C0N6FLjCA7O9/iS76YmEC79DyMHARZpA0
uwf9VcnNSGtS+dc9MiMECJUprNMcuidisJfpjawjM2Hn0Sn1YSfLtMRRMTKnBGAH
nEjckuGd9axFckwNCDEx2euMYdM1kjEF+RmKlh9U0A8nOwCIJ9o9oR/7xzjVv0dF
oAvayBvzIUtQ6fE5ROSjS5GF2S1NbdRFu35di07uhgTkCBhRlmrGDMy+D8EitoTX
H4hVYt3U/92xOKkQb/jgKASXeO+esT/jThaRm5Lzl7GDRONRH4QC/R9XoFdkVqLu
oOA+zMopxffDlaJE9odO4K+5lMJ3HtZg47oC3y48C4yDydFT3tWP7e3GggDaA6ur
TZel/rdr+5hQWL+cpag+tPuLHuoEhgIrStOR5Fcwjwlr3uZqdXOHEbS1ge+o1eUr
YkfRKAhOmFOxrEIWcSHWZ9X6OM0FrABQ0TkkA1cS1MsSirFSkTbFqHZNelsCBSi+
x1bC8AthbWTVtYROqS6KGPlXcj9cxeSoN+rNXbF83dX8Mv1vd2Jm0Ql8M2CxQPAn
J2wP5aR0TajdPen/aa7AT5SVAAWgejBsmAeETn0WCMYSVx6ER4I9gcugeXpSr4tF
U+nNoRb7mcimb5eCV+UZv/eaKotrEqB3beeXsaIEArzpHV6cRfbMhRr+okKtKeof
2YUB+qOsHictdZusPXcslzZsOHOviyPBHI0UU2xtWM+PXMKgNlppj+xyL782We7w
FWrYQGYCr0ciRzPGQL1MlWspftpIRHANUn8sAxLyPCSGg/9Tx7rQpBRUOsnDe2zA
Qsyev3W3HvySrJ8gnH3S52HyM5YiwdDi0CA8HAZ0YA+OA3iy/C9AdhRUNXhOjCHU
SsUqSsHbZ9Uc602yhYpEF4xuD1XQFr9Oo0BEYbdDEWI4KLBl7T57ab1zdCxG48c1
ftlmZJHwbZBXrWEUvcQOi1pOEgcef8b6UlYC5f2j9T78K4JlFCBgxvlHlerz/6Em
ybqds+qtllP5Lonbsipp9npbtaWjQefNXfsMzxT/gH+XjvW0yB3fBeEoMzWMn6ZS
Z68jaMTSSc5IfHfOwg/UuwsT0Sa+J62oMPFVZC7ex5EzlDscPnGYvxYNFxLzy2Nw
p7DVuT8udEpsK1dFNWDZSdNn/SQa3L1c/0ZiqOpkSEE8chHvuoPYlvsppOWlM259
tYKTXWwU8wIoJic1WQD2SxMeJ6KFGJa2c+3qptAjQj83HbIOGCLibQYvREQHCoXZ
Rw67DeiPkFYeWDQiD8yJvkYFqLSQiRkV7GIDjDEaZfqnGVzciU1YTGkdlQLGpUwA
RhPdQ9yMzp5ecLWvJItVzHP/yGz/gegBLBVLlKHA2uZnwd/v9GPv72icF2hxvZr5
xO2vOUFGoL7vu3X/VLKHivb5arfjS98OgqxoFfoGomQwUqc8Swjrkc6Yr/+fDnkh
9YIlnP2UM9X4m250mibwT0u+Qn5jzYKyZtiFXYIpoor+wHMxT35s32IbbA6bsA4x
C+EfNvZFDWxSAZxaa1ABioUAWSv11KbEfznXSrnkWQQoEvvzPAnqWFsyj7br0Aoy
RNVr7tze3W8qUK8YKMx0HHc3oVILqF7dA3fDk6deRKxMQL4TvF6uWqGIYCxN/veL
GeEhEjtercwB7HRaplYGyXo1/FPe0RN++H5P9Jj7SurfPfHWUNSJT64Q2iT4L3Pf
3JC029Yq9hHjgSOf3RnvPnx42h49Q+DRj7qNFEhv2aGpSdyIRKieb3sKChqFTiMp
EsDiHrVfjFD17UoLy+myIJZqB5QkN0viN3bA6hEcNDwItES0938WD7GPCwBBPfAD
be1tJi9weOJJgMEKv2Waqg6ItRo3IFD2kAVdCDf+632KAuQHYe7PwKQeqvje72DI
FnO10W7mM0HxouO8iJKK/SjRdkvq+RaFUggGCFTtGELGbfmvoUBSgDfYSdnD1gBS
+35SmvrJxlDBCXje901pDgyecqwg1I6aGHPZXc/2mTiMFjMEYIRctAGxJ1+S48gY
pHYAVEsfBk/eL5sSB95uAjrOK/enNHM48tvJO/280zTDRoaODBmrSuT5Sf6fGsRq
Tlj4WBg/QUWzg2XD2NoyiGUncsjQ8FdTIJtYS+7RLGYwTQTJ4Covm1puX7tN69O2
saEGsdqBhQHHSHogNWKOoDlI8ySqnqIXPU3leOvhoUuPZeGsTulLH2Eoz3rOi3k/
R7Ib4ChDSyLXhzzhb7a5eQ4BU7B9ehOGzudUQtL6aFF5Hu+DZ4iQpZoKz54YnaNR
5VxPSRNhpo83YEDRm/qcUDbWL6fuQaX/b5RXWIb7UPwYIJ5+Ddsd1iDQpjXVaXUr
04yYk6Y3zBwuwzY87W0ITu39h/9J+3C3w1jeYxEin9ySMFoEJZDstlCvQCLywB1i
mTXM+Lt9ePJLxy4hS94rGtOMi6ZJkGVzoyuSQUVlS4SEhCoUZ+DeI46urT48mQQU
wxjvrgdZ+CS1atdCBhTIHslWyWYHg686yYt6zv04jUvbCmTOqY6yVFBQwKc3cHT8
4wA+BD7cGZDqq/cig8luFlCsK5ydZQbJFBFibYQYvhZD/jLyDjUBtUoV5Qz+iWFX
TVyrPXHocln2mvUvqkidSDTxnzfhWxjADRRNx37qp4lGU1HQadWPAqYC2nsVZNNe
KaG0JhhgtsqWRFZ9zlo1+gRbGyLYqF/R+aOEkjG9D2l6BrwEog1QLKrzVCaVKYQT
JBdJBxQnk3H60/DcnR5tvp0jX1mfvqcTh+Ap1oz/BYDOdWBHd/Uq7tzgQvI4ntU0
1jMK2+2mRYzOU194bPiWBKrl9MWS8BBy6owEp9a7u6zTdnI53cOMfgcByDufOuDL
dfUXXHW9kw8PYIkzHETrVnolprtlo2tYEozpD8PJX5phAKp38t8cIHmX3FAFsQpM
nIKUCG1Wzuh668/1bJ99Wlwrp6mHoOFHa9G1JVu3ES4nedu8/nPTkIuK3EsdU67k
iKWPGNabO22JnhbH5EDQmZaE/s1NuDghySjeEBz5CN3tH0xAZyyulN41h74QypVn
Z1eW0gHV4vtqQn8SYe8qvgn2dhY6t7r67XP676TEFjwCPayX2vaGNwY2teggQzEj
gp7fc9ENfQPXrrTd/SM3JfgmPTzlNTpwqFZd9FH1PDN3vpqqKnq1lDjLzAk0AIcF
uxWzkYpL+fBDjYWJsNcnaZREGmXVxnKhqzMXAOkzOmam/f47NnTCewjHZQdccXb0
arBspBm2I4x9uCu2SwR4pXJAhoJIrh3uPB4YyWSBYQ9rCFk0jkbCzPf1b2FYMozC
ljf05I0N2egBME/btCaUURW6dHeyCdCmgWS6+nV+G7ck//H/R+Wol9yBclTS1hjv
z6FqkBLfqX9JQE1XblWqth/bRgAFiLhfmHc8gzLFJQjxsej927t99Z5fYvmRfQxM
Oipvt9jCgky3zmNL0FqI18OrsW5f7WjMLIoxvKx8xBsXpOp5gz8ZT4YFj4aHmzO/
pB9kVuo9Dwsk3g1ViSfwqyFFkka/apQPWJt23ZQWC8JzmmcOfhhDdcYCxEDCXt5G
NZrZzaW65RaKH/cA+ruevhthUHO4V5Qq/DWX5BlZYDYlA23XAM3SAEhcKOEGd5Tg
cPlztZTZ2RE0WZ+h5dNvcuVFcK2DorvldnjXmL9g1xaMeJfVO0q5jY3jzh+m0hTL
oxFWNCU1GmD+8Tx34YRXx5jN7pbf2/SGsbWE+RzgGKpgCMmUkgM5WeSL6iOP4++W
bo6+tLEUUaTigDfOUwSpshsP2J20gpFMbxOGFITB3emQbCTu/kJA5+pzaepspyrh
sV6CIaDmmy71th9sko1yP8pigJLzGt6pXt/t+Z56D/alDFavbpmy8WizEFTOBAye
IzrZu7Em37AvRcqvcLcs3aGjRM731Nns1lOjTS/IjTjbntUL2CcGxgI3T2zm3y/Q
VxLuF2/Dzbg7VzAyYuPstEQeHRAviidQ1tfUhrTmpfxaPttIjj+Q33IRsLMxYrzr
UoXMNmJxBw9tBtFGypi/EUlZrl7ncY7dbhce7J79kdC+1bToCRpgmfv2BoiJLEQ9
foGymVTudZ7gNGehLZDUkA3Ox5YhQsXr6FO2M1vY9yoYD5piYKUJ659namFFfi4T
gezMcwm1GFVr0rmHKZXSDNJ2cDBlK3LGDfSsrz4Z0GHWD6Od+0F2HEUM5gxLVRol
RAoaLj17uuLEhtRGbLlcqWe8dgYLB0EHQqq3PIChxTkbRgyms12l0Gy3Jq38fFh/
hZJomqw9OUempyV4E0Nfwe9JDW9gh6k1BTsWcFbkm8fNAVjPuHEKNIJkNgToK+Ej
8bdqkFnn/1zuDRf4S5Nxm76UEl7Rt1xPFA+mvzbSIY4pS2AiUEUnGYan71nwf2YE
/I0IwWx4dGaZi+kBPHohWrULvrG6qYNL6X1JUxB5G2UrDUAhJpW/y7922l3Fnce5
pn1Yk8+MlGMFZICrApB3BQVgN65k+MYJ9+na09vGKOfLkJNnpJrgefLsJKgdDEV1
krFgl30iW9ezQDhxxos4Tf8JVQ+PfeAcpiAQvoPW2W6GtBz+2uW1wV/3eFv/ZqfD
MPj0HPMImoYbxmld4ijgwJkS+64jhkwVVcoAuEGxBabRKvhsgF7laKSk02fjb9Cp
DF/rCQSy1x2gB+yovEJN6/7xDAOsngqumya1Gx8wqk8Wb9ICLmUyCvYr6+aIJiF2
1yff0TAWPPMomAYzs0zHbn14d+4ZQfbxRq7R6xU8bYXUpjE3h/euZtgXQ6kX9l6e
q8KG8wJLZfF3OtpZpAV9+4VH7Iuaaomfibwny+4ciHR6CuErF71v1I4DCZOQNNAU
+CSjM2dbyrBAGJCSxVFcYUvvTyG8EsFlv+wvyWWfWZ0+DAQiAyCw7kpa2/k3maCK
zvF2Cp0WZiCNk86VDO2mfBoE2W3IdcFojjUhAqZ4AnUgax/c1f0146ofoe86kQF1
Wg252HJ/el6OEgnFuOhnimqNU26eZlOl6550Jf7RIjIrmF8YZu1lGelBw0BhCqDK
PJIPTMnYunOqinBp/L+LmYlH7guGzkgqJMesJogYG1ZwolcjOYvBDtMHDFLK3SnX
TEEpOVxBViZTHcilZu5kvW/95OZl+K/H7iGwhHkaIyx/e5bMaxcSn6kcniy5GlS6
sjoKuF5QuR3VqNsBDQPblIWQdgohIr8RFZmbGYQ9khBRAD75BRIt8qlZzBWDZRqg
lYYDYerzMXbyHA5Mlfo/7Pq8rVIZQ5XxSV8Juhe08NEGtL7jCuho7NJWNpkW9c96
D2/KPJFv9hdmPSujSF47chly/Kq41Q56Pape7xGUaEM99Ra46ndiq+wD1+2czAJU
VRwwI7ftnzQvYGi+9ulbxo1LI4XT1xjrBr/PMkI9H5XUIXZz/JaUkmxYGqD8OnBE
Tt3P32MyCERGchMtyY6iDOqGcU8qQdcMT+HNC6fC5bhk+1IZzu/snGWOlWkDao+G
P9ZtF+DshC/Ve3A8XuGGz+wbCzq+tKg7JkSnJibLtkpoGzQphi3lwvLWt9gOZMV4
Wf/l6V1YKQ+R08RJZxcvjbJC2B4BOmSCNyYg8YtAn2448zgoWq2qSLUh/jFrkP3f
+vMxiQofADyGmTIc71VoGkP72DR3QkQN01ZHI4I4WCfHGTuXuSqz2kS10rCHbUOI
BG6l6iPXngpiRTrGvGm3y9C/Am2fMOuJveDTvOsIotPeDwl+7W4PyrFDUxQpoZzD
eKPo9hAm7V9ywbUPmsFnKKviG7ccjlBO47+cmwozq+RRR0e1g81Hi4U0okNJYefh
gRY7BLkMTQqSXcW8aNQ+HToUf5nU9W7uYBw5Auz7T3VaFD1tFDeb3TlQl2CCH2pt
BxFBVZU7Ig3MoN06W0i18un1e7kSAjkhjcfYBNYXCB5OwsP0WuMuuOE2tsUST0DI
bqhTf8fj8DG88c5eVwYG0x9TmZO7m/VIuvoHDj9gPynFlR0W4jpcJyceHsbav2Nz
1LjdvjaTgxkklpRlDUOp8R2oR1q+/S1lMyDNpsk95irx4XfP0JIN3/qbI/wD5mc5
2eqUPLcV1V7OFIu/DAeXFNsOzQ4QOLFP2Xs2/bjFnR7YTnGbRfrGNj/RIutc/hR4
iu2Yro03nUQqPlB+AZmBj9mO0ltdSUwrmy7lC5PcNyUvodrhEN9hzPthkXpqoXMR
D2cOexN+x8pKiWJwYnHByA2MjILE6sjtwJh3JDEuDT7x6RueZ3ZX/LwMbblmlY7J
BbboiE74lyrRxYxy+qqjPu3MbByLunHoghRuLI2I8MH4JkqPnT5lGnMRk0JhhJvB
8wuWS8bludxhvKU7pen80qJSyjBORPp0kGmmgisMR7Gz8t1EHsaCXtn0pvaSRiQW
IssgZ2UFdTTs6xN79ec1FNypYKPhk/L2twRkIjdNIaUtGRuVOpBewammOYsHb4EB
OZQHztAdfJcmwM1BdXSVESELPkmPR7hb73Oc8efAgKn1TEoXa9URBmbpay94Me5x
xgxk1VsBryIxFLPRUeG8AGQND1iJgaGjVTTidpdrUiQWUzTTJtvlOYwd5+DIzR2W
hFuDWRZ64X7PpuAn6wH+dwP5kyFSFa8qp7NoH82bpqDw/huxZmiHAV7CyB7ZxMPB
Ek8pho90g3mdHhp5OIsLQRPE+8wR9V81TIGmE/9IWlrHaCwtPZXPAFBzxQ93hMHr
8TbxxKY4gI6V02Vdbhg6hbdaLvxhIxpkQGhbHmqTaWZG6AGPNBiUXZkq3Wy/bDCZ
bBbzAHnOm9eKT7o9vvPpZOVTtesuVrXRzkeSXM2NC/t2LaIlg/bP7rgSmyukvcNm
0WKHOACgK63B/k+l51OOd9fWiTq1RK711A+8q5MCwyyN2CsjHEgzyg0bXydlmnSi
36oAjNDvr2qxtTwxePj0MnKnNphERpX6AhUO/y/4iDKjO0/pXXbDxprowLqdRizD
4rhF1Jt1Sd/5r1KHjVXeXzIm3OrTYyOOSWS5N8UlrVEUwH/PEU7XExqVf9YF4pJ8
9qnsM437Z6JMz2pKvrBSjAJkrGdC6+NadhKiyGk8km/+wxtLSy/3NmJ51uGmEuPl
FgR2oYRizQdLxqY48JBdxOyXdR9VAmoaKJq2l/gOEaPNzyjvhXHp588mdhfBoyGt
Ys6KuWQJvglZy7kcLYLnlxuBoz5Fam2GoNKsfNDLR7FwTbeI9ZtYYcz2IKIHnH0X
ABMVdRRzruA/cbRZOwnwtV9l7Q58J2fm+YxDyjR6PAMSCABbEnk3q16d2XJ5jZQt
s85SqJGjJZaA9LgGzhdskrxHzKBx03xfttGy/QPgMISHl9WdnhJ2n9hJp25r7FjC
ijSKpggf+JHt+2gj8IS1CbznBKKpzRnAmhNR4vE1vDBPC4LlYzG+DQuHeUgFbNcH
XgB19LJt/do+x9iuzzcJg4fYTXawdYeBlBNMNrFyszh1NoTYtn37J0O3X6i48Qzs
Y+K66be+9mEJU1FEwPGVZ9m/6YjKMIWaRgKFW/YmfcjieKtpg/8PW0OS6j5b6Nmf
rpsmPakH7WQKM5yZ+csUOFEegfP9uLHhwS85eK0pyPsT5w1Xbi9ky1BZNPl8mCI7
mKExJFz6YKgm6miZu/DTDMYrlfm7BJ+IVbrRbGZYY7vlCKFXBXsYzjgAtImLyV5q
R5xGTXVlAtY3qMlxSg5AQoybmnTgMVO/9hW8VXFZa8V6lOBEJcFa3coG9ohUHKCw
rsaecQ7+Hu3KhrdjNJuq1iIop6cW6K7JxXnqzzy4XuAuqoCB83TfYn1YT4OznpnF
v/FM+6qzVUXkDTq/3/nfhXHISx0C7GaCiYu68OeNPGCpudHBhLYi3dQ3G8vKXuXl
m/4WHo7LAmFpWiLX/NNQw2ZKPQa3Qsmrm2wDED2CS4duqLbrd0W+l8l1octykPsp
3pr1tSJw1c7/LB6BtTc3YH2awAdA791vGV4zJsDnw/TRvfmLWj1BpkG4SsEOIQSo
NH18DMcJIPzX5vbX1GfsUBNPKn2Qr1xRHDmMbhbiRWnrTTxxlDy7CNKvpahsXjNV
uiH2DMLvvkJ4IK4z1Ax1QkFDFPfxQp7A2cpDKSMl3VV+org+QOJ3NEC4EISXBkwJ
3EbdkHonyZllGAS6exE+pOco+PO3tJ0hmurRSpZfOS45vy2KGkp10appTJ/OoRUX
5/iC9gaxxWAbIXOiYwT6alRsKQec8g49TGbgMILwE5+XxWUvZoPfDse6sD0Z669s
esncquERjiwnpRT5do3yJ6/Uphk1WOwJ/PFJsHYLYvx0QDRwX4pd7b7cN2t8mpMP
n5B0Ltt5XOK0/MsmkHL6XL0qB2U23u0lXRmcRCmyR17flvdGn+eXorTsFUB+Xlqx
5cgDYhvyiI97B4eCtLAHZIzWs2M9tOy6lH5052RvhkoGboThGAWcUN9AL+Ydl6RB
snLUrZgPVhlBLkesQNih4XI5YWR2gsnS9QFXzwwiYhxHj0/JI3RrOomRQVfrjjiF
1KnyppUsuKW6KBTN9v/1WAWWc/KdAYY16Qp8nZLdANzoByrY6PmKs8Z3weO39Zt0
2gzowqDDW9xDjRuLxZtWBZuq3w7RXZD77nbANinhCSPmkXxfdgl6r9cfq4jRyJrn
yqlgxkzY3L5k9rInQ+V+Et/jS/TNTVRYiWifcUolAz+rKmc84yRUUZzAeUUMNw8U
jbf5nGZIj1NER3XrvMbmzxYnwZcFm1Y+NHI0fvYxvWSwazjWtxDiGHH+txZGrBAS
OMeuQaEkK62iW7DK5WKtpiVHhjpPaU5/Etp/RcDX7GOyuhjgKqFykopT6N6CzqEy
eeUbKYx/6aQl0MN3ArSP3TxRQF1XWuACMdMsPbgsHGoHoB/qv9mlpu30bzoxlKv1
F4fkY+UTdAesDZIRpADtomfog7I+etOS/cyCu22sz6Z3NJlvV+BcBzN6XACsixG/
LNiBUP0hjktKElT9Etf++rwG3YpSW4JuP+gsvjs1I5/9XQ3hTPP9p4P1qLoPSSZ5
qbMCd8dYyiHqSDaIxBFxgmvVBczPPnfmBHP2xD/cUezBiPJc+mu9qbOqoAF5hw2W
JlF5o/RSPp9VH9bZRCbWll2QRsydd+st8PP4Q3sB2TNWTWe/ccHF+OuucxkHrMvW
Gugm9/VEGZxN6TasdfDEd9cq89UsPXVV8ZFrt9jha7PQfPWgvkcOgaegiY0S53p5
/Q5XRuH0FXofNI5Pxp8XlRxtQEqH3rYywcWiT65pmn3AIP+ZGJmhalWSRUxQpt3q
eDrRqLivOSEx+2ScBzjZwbFAQuhK3jaLJ3K8Fz/X2waQ6c8iIUQ2GZrU3E/EhESk
494H31DGgfhseQWaXPzc3sPqQy7C4lVe3II5AjzH5uk156o5TbkPH/RXyOQ/BJPH
Sy37TYc41xahXDyzCBfyoFURBIktIeAP2ajYjL7MKQKZgOMIRafBR0+C1z/xEuut
yBEddOOujkYedcaeyA+d2WbKN7eVK+8Vc7fp0SMlPAwHWdY2LJom4C/W8yH147sv
/QZHF5WQXKqRf/Js4rd4vctIBALTNMdwRB96hVHw1BUCW/BcJ8+/Ba0Q22IICYOl
T5/58c2w64+E3fBnVkkhg3tr+fTZZAiK2Ob+dnJKbGCybbQDJuOJYa7IP4mi2Prx
DCUa32AsxBGTwMvBHNwLuiCxr4vyopj5f2mbUluzkcIlbU+HSZlOVRL1oERVGhDB
JyjtS4v486JIOEO4sCvQg7Mc1nf/dW0d3PGikXD++FtRD9QU3pfpXLUj+ijqgr8Y
EpSDNkY/8duHSWX/dH9TPH0mjh9tkXAKxhrZzIzWRgbps75zche6GW1Lij2M8L5q
mkQuY5/bc+hbbUFzZA1OYjF5QhtfksoxS2PMZjo7DnCpeYKAkIOlqlaublvZ2RM+
r4SriOEun2GWq+E1/0Hagw/94/EHoofFn57ihuubJs4cIpKYVLLC6Ky8uewELlhb
dMX9ib4TfBxrkVHRDfgrQHTuMH6+7Rm9VmgWaXmn56i6hSA+UntgFIW4xk9nN8kI
W6+2aK/JxXFrWVBJVKw5OpsUquFD4gyDF00BaB6af9XPckbvWF5ICj8HsNvAN5Eh
YM4p5v3+F8eOlZpFT86SiYBtX0sOjdaHq5GbKjGeIKFZXyfFBLWsK6Rhnb49YKEk
YJ6b1vzTHZ/vmNDGpNRrHdpfDslC8MM2IkLBXeWVSfIDs7hEd/F/v6XkDGP92rs4
eDZ3ZdldJh5nw+d+Ku4s85xHq75XpseIcGWCmcgnW8scMlOBYo2UDtKBI45Eq+h/
jKQBY1lLcznISALY5LHGbhV7cuN3dywBGZSBIoeUfMMEN+XjHK0uvufGIN4oIKEA
7lJy8uJi8XIYOw6jZlehMqSxK0a0GkMHDmpMoyBA5oEDzgP+oi+chN+kOCCPR3vu
xgQirZ4u56JJciTzbSIfcoF9vs1Fe+aroYcCmj3hJFeItyKKDa6Olfrwq8NuhQH/
xD+JOf3ZnJ8SAxoZ3Kp/zGG9ekX3XhVnM3FjL/dy37nu8TcsE1rfhjenBHGCW6zQ
ZgcRjtYM/ODfiTXEgVBBRjpHC0YnXxSgKvjiXwqEi6dYSekwT1UOD1NAsOMDIhTQ
hD4RqpEGa5zY1ni9EbxACTu/TN0wphUaON5EYI4xalGrqFV5vnHf9dk43fM9vzWv
q6g5pT+RXxE0jVF+O2xzo4zounQxQcxife9OGlYzZBAayAYmwwe8onrPpCiB/Q3m
c0A4XDSzNSjHabw5ZmWc/tw+kvgEIKBkdel/cF+sTVUWlHm0chWyUxNsJtncmuS5
FhEmUMADecOU/xe30DuSYIqBa/8nU9LhVH4Qnja0Valz+u3cWViZr2GVbvFGsgBJ
ihDir5qrv4IzygET3JRpuyM5mvzWKYlQ7Mq0Jh7WUOlrPjFLY0fkpi9EVQ6sUHOe
3Zd0/OSZpWNxi3o3EdI2MEwZjYS152V4GrluLCNQ7X8rde4skSRpa/Qp7P8Zh0Un
aTqhrFP5Iwwno48XNKNbaWuZo4zwkOBQB/JhSbEuFdL1lL3sSVbJu9NMzwZZwSkQ
bckZAaucuIzGJ0jK/FDj9StwZ3Y5wlBtuCOtEXtafvY2JkpqZs6EEWrtBMuoOywE
i8Ehq0KoRVRCvsvkRaU7lAuLEmlMfJI+sdVnSXpbQ/T41MV0AcxYCG5V+vp3p1Ub
G3imvIYUgvC8Fh+z03dfEkFMnHlShzNAm9WI/58zFk8AhFXQS4G/3EiK5pi2edmT
emAhe4YtxijYNqdcS+hkHrjG0ERoQvCUlmEAQMzLkljoVFVR3DvDMdrzMv9YGdie
Lp2drBwCb58+bk8BC4M+faxcWzm2sWxmB67OVF8Ja1NjKbe4dChn3HyASrF0ZCnN
0HPgCHspGYKl92QzlFewDnbwvJaZ7t9NBWrQ5SPXpDoXOunHcZ2NODjpxXTogHj2
sWKhcsdlkizD930n8kSPms1FEzilwDzVQ7xyCQHgP/44wl6uKtqChrt3f1qjeS7z
4+1DNjRJ3Tk8/rDrJZ2p+WTb1wLMlx1H5GwTKHhgxIwAwX2aaKwiqOw+TCSKEBNk
wt1sEOZDZgdMgf27aDqgqBK+iRxK8SpMVWlfef544kxBNbimAB57ypavx8MbW1UJ
c2nOVF3L4DH6KL1UDID7eKDAqWkWP9dWRKlwOTuRpPHgrvtX4ZHI5P2dF1omWHJY
l6F6bktggLBEjjXiIr2PO/gUYnWFmKVzuD/QGhiS43auPbEarpWfWktlPGe8Tl3x
VGxqTUS2bDEvBlx6JLr6g0V+O/K0rXJaTi6Lpe8nBU0S1z8s09Q5UgkIa+HEueMa
qgom0He+DukRkfpPtwvEDYvMjjGqzJGkC3quM9W6hFOkbJP14rZu6YeAM/3eJv+M
JYHfdnyNSEimGiaw98esThGWVp7L6ehecJ7uIdUF36vRf7XNEKVggTbW2ZVSf4BN
WQHMxnAlWsenEEeCSmwC8lS8EtmfWQSEBvt0GM9lfDW8Y7oSgI+2g3zBD1srv0dK
jN1Ju4f/L8EHZ1fn8R+saLK2agjumoVJ/XE3ie/p5lkvRolGkJElcOkvRM990+4F
Ekn7z9WL9edHRVQtAQf8t+gkmeXmPcuAxsnVwridm9K+00gONaHagHAnuRML/APT
xqWabR5q0GiMB1ibzQIxKxs53HhuTdk9xLki2zU4/9pkVQgwKG9saIkyn1oT80Xr
G/diQ5xk7o9BhjTk5mrQYD6RqXhTDyFzXOWpqzQifDmK2J9TUiro+qPcSjWUFPsu
TfR5S9KS5CrKKV2bYGhmMK4Ta9NAiyGb9pf8KV7YKTGTB/FUwtmj0SqxEvztdg1l
yAS3hA7CR0csR+wWeUDhe69QTLJNtz/+/9OA/AtaQf94/qr2UVvIA2UV+TE0UCwE
fUEqB315ETx5jjVTGK/7KGEX6FsWDDgzJmicaoXUIlya/LQy/MUmAagL0ds/Ivb2
/AEUbsbb+6PSN1OoqoWlXwJk1DJRvPHrk7dtpVkNVHeOfxY94HJIwAd7IcrKPxyo
siGx+5zIOe00Fod5PghCxbnRJqLMAirdnJAD+5+8pcAgDVIVAA21pwXt2w/XFUDS
qjnVB0aH7w0y8HPI0z5/ETgw3rmYH3k1CYDiEz1PNUuqzZG3r+0blmngfxPS4Qt5
lQ3l161eSwJSjghGtQZ49rj/ekVM3e13mQlwa0+n0GPHKJDGj/wL+dK55GZtRhkK
JLJduY8TFZrLexe3TagYkwQsysgoCEYEtAHfswmvoXITcinulhmhT9i+ktGlR9n0
DefpmPB9vZllu3lpvMUkZMgiYAgl0eRbwRm1LmqrgkJyVGWikMyKVh9O9slg9NDC
Nu4pdTYtr88n+9ei7X7z0OvTb6WZSu0WqA7ROp0rLjirgDC70uFWPtlUgkbooDaA
Zbc7kC7pmyLlA4pL8ysFklAHcE4fzfvRVhP1AOXrd81zQNKJWQWgX5rA3vZef1BG
+l1vUoM3hvx0nURPH5iC2bcaA4WrKc9yFMUboqxZf2WzUTHnf7enF3bqVitzlA9O
fMatrdCFARzh+EtP4O13DPlqBDeZZw2TiwOARWXGCu7y0ID29I/XCEViwT1bkHt2
09FgDYg+Qd3qk/h563Nd5wDon/X6wlHRSAvLkCNDXAno+9e1d7DYXEPXkEB3u/bv
oD5um/H0RPREvYunn0+NbTk45Lu9cziVYH2s8bmp5Nvuvy14E8xqwfRaqRhPZlNB
Xz69yOW5J9XFnuHu6EYo303ih89BIQdbWGcDElwEntbEaGzpkegKNXV0zgwFSBtK
tj0D3uG7npAqM/bO8yMdn82LlRu9ita2oETvgbGNiQReiHWeZtQ5c1OXCxE/IM44
2wfgZw4C5x7QzNQISFEUX2mzHbgYTGsHw/lJOoXKL2IZ+FYEYxzbt41Npwc/roVf
e2SuChKOmsqb0vetSeMJkuETaxmnGt5qxxHwN5tw26SAOyV5Z7DwtV47pvv9MxKy
6OhPfC67Sw5VsX4HsvupLcVSqBH6IXbhyIJRZ9G1cxAgnVSybG/Hg7PHA2Sg1Wd4
lGjumOwQT+PPQFGuWSU13ZHwArgCowCPApeMF4yZmRb3Cfc20CI66uk5qKk33eJk
oOsP/hy5HLPeG7gxzr+qXeYR18btBo9QpttQJOOvQevwjIKEiXvmL5HfE6XC9J70
zCUeP+Sn1xCMcjXTZVEBdb+3Ys/naZvRu7tVz+07EWzhjksQ5otNIxZZyXzdwqZG
1VWjCOdoZJ+oFyoWqWLLOhowwT4GwMr7nWiMyeAzSiaS6Oz0DpClK//mJbvnqIM3
X9O5zfUtS6OyuBSfLxZMasBlYN6HSsU0q4CnI/UoL5Q6Tg4AZpRm08znyPh9u7Ix
6TZiVspQu57gfsBgnniaWPqBOBeBjd/6g03lg6uE9sviakdA/083uMaA0hrsFpZr
Q6Q7pZ3/qeUx/tbozSRJV3wFUiPIbptKKyDhWkEoUDeNGirndnDAzGtXI61tzZAr
sKtEHiSfT7xCoBHFsCBjW7oLXOQ3f/kNZ5UXwb6gNJEcc8yaOhMJNqtquz0clXgT
8a/ZUxsLKIh6lLZPdP2e4wVOEyOlmei1RJXesKWYP5eHslP8Ysuteh1wHpPINa9q
pp+WlMQ8p62dQYB410JdJT9DcLPSnhaN/tHkIXOC7OQsUYe9edskAEL7WGOXzMx4
ocPwkIyJdqEmkU/VlaY0wCsTQiwK/wBQ0z99nxAZlKS1sREy8zp2S5Uq3A2Hl1xC
tSyqi3nJXyqcgbxO8W5XWVqmwvmOxI1s16pEjUVnKOEMU6CU8k+b3VdLLB1ZmKE0
iEKCoBMLErsO81wrYwHPCOu5SRcgUPWbnia44Yh9w4XX/CbfsrLejampNMn0P3GP
YQjc02Kq24uUd6L0iCf4mqhJvqoiaUVy3/IUSljN6D1bn/Il374DC9UsPKLa6Rw3
F0OfYGayOK+HMwTgKadvCJ3achTvJIYtD9SaNrWYz5zrxkhLj6tb37B3c5dQFfPy
6kH9Cg72FHQUtn8FTglyj+14PWkLbNgCQANHs6k4pXGbYXV16j3NADKPMXRWZaNi
LBwiBIPAmE5/Ny0CQ1ZgsDezFwo0BZ0px7D7gvvWKONEj5zCkJ81c/cD+sX79WI+
7aoy5V67SEEip5MPzV5btaZjklrbgKTfKJRWn5IeJIGLKIQvPzTtjIfxZEr0El5f
j0U95cwq2rq6Bd658ItwkbtigOW3GAGdckLBhdU1sAsdMh/eBdi5bmrsL//kBYnN
deShPuTkzKQoIRoBdOAE4kTXcwyz230Rzr7Q+U0t80s7UfUPFK8kaZq8m6vkNmbr
bYcLnA9jiLWtVBxcbeYawasGs5XVp6cPyzGj5Y4IPecTYtEFi18z/X0nmNUPO/39
NlyUcmgl8vzcfmab9aDcTLA3Rwco0aADDioOU7147kCIkhiyW6yUQ53v+Z6igaei
HENdvu8DH5v9mV/kYTdqbfqNn+xt33b5VilWElkpzRoSiE6m1EDSW+n3oDUyXwEz
460sRy0SphgnhJ2g21jdNE7LfkHeN8VvV0yebRzZCZ04ImAa2T0+6uUbUbPaVJr0
Y4uxnW/y0weYbcB1O2bGXDGZ0J6OaUwCFTr/RBWL8yPaDni3Ms/I1OJ8dE6lt+2u
pkDPuOFgeM+bnL28XxUg2qmll6VlkoBFhCj9eOCA8plDKaq2fLV1NSfhSGvRj8um
k/UBN1FlKaC6legix5vuL/LjoD4lP22syccYzte3xONQZPFHiBL9ozaAktQ7qGn6
r2dhwXUex+yE2CK7CnaK7sqiKUh6utPR4k/d3OZ3/lf4mQz4ObAuabEtCzmcChR6
mnE2uXzfJUCWVMbXl6DD+kG+TRDhzxoAbY9wqs6Gd3g37SxjnFFLEkr2GL2Bebiv
bINlN7Bjr1SGdSOr+5BX2VDr9Xcz3La+bBvBOuxMjXbZmxbPskRgJSHxzSdSWY/N
S0PCDP8kaM1BXQseCZuW+VvdnW4wt1lfc8CF4KMJHDjcp2LbjRv8xneFyx2LmEEc
X2xGu0HdU9cQAaO2H4QUxqR+frMGnWeAyi5Szqr/W3iaFcf/IGtsK1SjtivYtWQp
he9lKVfPIt3To/FyGm+OHbok9vMmmSJZu2bKyFuBh6aCBvH2kb+Xs5YxeMSSDSfF
LaYwIMS0abtwVHX0TSoc1VZy/iJWPnENP3AV2+DkAb2kVMziZPH3pG+3Qn2R7iVK
II7cBbvNy6dOgqUrNEjn4beXTXIItaZ7jqkKHJkVaG8kE3BIrJUOVEf9LodYSNL4
A6CnvviZch2TjkbniEebSpD6NvUtNGufGndKl2sbMLCnJiCVvlwgIEuJA5hB3GM6
AD+Q3AUKTi5V+v54enrO6cjODhHo1JUqiecwaNKBbQfar6wzSocIVx0fyJR+Tc+d
3AfXRu2D2O48Qq248zMbiQseB/qRtu5yXwIVzmiSSquXu4gUSWBpnshSqNNARIMj
iNCbAy7/tt8PE8+nvzLIVdBg+uGAKyilnmhE7rFORGyh/4pa9mpeXlVvW29DrQlu
4+G5ovStJtGNQr3oIQ5kaaDO5tFJOBgAeg5gHu2c0uzVYVN67n1jtaeToaNb6/YL
iaXo7bWxqeUqBOSO3I8viCWK96hELOllhz4EQMOLwCNGucDU3DfIwmNi1xtor/wn
eR+YRBtKR0S3NAfcoBYZDIEoiHvv/YSXInYHi6Glr8t/1BVYoi4lLKb4O2CPCias
lakVkACaHIFvSiBFmNwHjJZzOqVrOq3m7eZtXE9sVzHnudUELCdHDTqKxx77iCVO
VxPFIoz4AUi3pRWze4INwKJ3qgz1ddqvHXJOgp4Y1Xr880kLHxVELPBPDhcEceUz
IIcHoEgy5AvKZJ+vVuo7PejSbTaXmSWuB+PAI0tVntyoIx0Yb1F4gPFyddvyphhQ
evQzcqk1rZ//dp5YobzIOOuzH1PmxKeP7hJIMhY902aQgOUx6e8X2is706sqxyIs
pjeAFOGt/f4C+mdIedC9C0vTc1FnUKX9n/Jye83QEfASFpiyqHz5Q8ALH4kY9yBR
gouDed1RlbpUaNANyoydjuyHv9VrP9Aehxy7KMdwu+DWwSrEhAfr44XJgTA2qw0/
DCAIjtUfLOihvtF/K+JpgK87HSh+z4a7gaelG5X2AqLpzcL0zEbo9D9e+cnrW8w5
sngUhqHkU3BKzx/dy6dVRTEqUckF+KFfvi1AB4iSgSoL0MGE7g/G7rXgNqpkASPC
pNaVh4ZGFh46MrSeguMJiW8p3FBw2HG95QWqPdTlNC60B6IFq/BBSnOb3MoWwhNG
VWTovjlV3YFc7SaOGC3yRgj9s9j0/9bQ1vWea/pcHvECD9yhD+pwmxZbTvDGPAEy
xE3d7lz8yPhhznB6WF5VNyvD4tpzGbm4H+GEsgSQR/E/A9Z0nk4yxsZrg2WapXhg
wt5WX3sQw9rHGPmRmTYhZTFHq5qYyXA9DpAow1s2NCEfFMX9DXUfOPpZ4GJu8xxd
fz32s10AvX43Nw6JZuzYN+K9TUjPFXqzI4ZsludsTo2v+a9F9DMM4Pn9pf2eT8kg
KD8bO9ayH/pylAvSiiPTXFa4k8Ss+KuckCZ2aoXN+KuiPvfO76XrTyJPKUNtHQm5
Chpo2EVUlMNF5q7ZSm/wGoS63q5EbHWTuWaeFLfiB2j7zptnsa43kmFGSO0zToGO
s7p8Y2AzHsbgrWvmIhZ7tP2KZz2g/86hZqycCPxNfxgZ9Ex5f61XBobS5OcjxmfI
E9tRbZnZQ/reopfANJqfCPAT7nr2bMK+gG5AcP5eZMaZjT7NOAR/V4zxg+dChL2x
ezD189Jfr+twBuS0hIKqo2zyVZd+4RtVuoXJxuYfiigJItkcOcEtqtY97to/fFxZ
2SrbxFp0xjfOkIv/Qw5C2Fl/wm4d0yXDhdq2RqUHQVtzSs5BNU6TXH4ZApYbeR4z
81kZG8yMErbW9hH6RoUA5ceqjsUnoQvNbvlXxrh0lJWVCjcLTEzwMaMaUV5LJRhi
QC34+wivTAciTBStAz+9prw7WdyQJrCmpKA+DbO7myr8DW49gn97Q37pN+BzjvI4
G8TyjxJsAsdfYcMIrxQS58esltq1RbDnxMzx5eiM7DiqfX4LA8/YJDmtOIYGWka1
gXNjlk32fi8e2D5NKu6S4MfzGtWAVE6n3DVLY8+ZHVcOOvbEjHcqojMHj9W68Goa
nxiEVrNL8oH0XEIlp9nZd7HWBMeWWaI+ie0R5HcKHidkrDI++r+FEQy3/2JoYvQJ
swGrsS13dm+7U9o5Ozh6zIOjZ6GoTogOMEqlxc4gpZcISSxt2mZNP95HWzF8mXzG
Y5z8mVgVRwVKIAKfajVDGT2pYKMQUEk+DQkT6+MoASdRFBveiatf4rHytWTHr4FM
QMgpfkmVrhG0dMPZx4NiWmQZe4ZwBtKayscSEOWqO/elNCgD5M5Sz+N5xzBL1PB4
BeiV9IXByc9LQf8dhwLnt20IL3/qHtUuUU6FX4jetXL2x2lX91AegRZG94mtMm3e
bBi1q54S4HnWXoZ3VuWwLZIOTx28PSi26ZKaEUihPJ6/unC4Z10l9lq56sw9DHVt
BvRqeVoBIESVALypt5S6EFtnsAY4ujOMMwQ2Wz0e15BcSSEIpsF7bil/KOVqfbXi
2eLp8/1Aq7XJfCYfJjEwvEQbk3/gvSL0Cvn4Yv7LI0kgsZ42w8Qdj6TkvXHyno9V
fbBmZP08eUvmaXe1xAeyx2DZE5A4k4uEcMnkl704TRA6qdq9MEmNHPFXSPvbQx2D
svw23d+KgKoL0Al3lseOXEPxr4c9GN08n7VZdbDy7OE41wtlx703oTvTwegRbgcx
CDPaRj6JnP7SvmB7IxcG34tbk2s7hpjOEqFu8AlEXsEBYIbouh2YR6eSYzUoaME2
6ycv9eWXfLl6a5YzXQfeRL0oAvw5xc5vOk9FySkDxos+DF3dd6ycJN//LNypHjv+
Em4h8Me+GjquyfoakvahsJ+zvog3txAP2Ng42AQ/gnr2xmhtCeatjX51joa7yPxF
qnEFmm8lZ31MinKvxCh9KbDz1QFNRw92iz0jfDhXSwPTNzeBxwNz2rrt5iO77XgK
drua9LP9XXk3yp6ZGTslaMU/1/s7YHKx1u6Au8b8fDiHB/d5A/TWeYF8kjZ8rf8+
h+hwXxo3K39xJFWQ/DEGhleqDaxKhOHjFSPv1o5c9crAPdbC0vNlxw0/upVnZUh4
5aje8SUoSdUcWTkFS/A8X6XZJ+DLBsOf5e7rokJZmSfpXFRJzpApE+xNXh5XzZYn
lA6JU5S3BWNeFIGYJ/bP7j+27z0N+JK6ZV9/uaCWMM5ALR7d/dfm5EMm29pZ59Iq
+3MMrWdeX3AWXBi0S+TpSzWvqHA/LU6Bg+M9cFYQN0IrJ09S9YW6oQoocZhl4f6c
ep3XIyDvrew2S2+BP7oX4zRJvnueY+UwP2NJlzkx6puwwq8ninlGRBPJbFv0TGhl
/qLhIOeQKezxW7p0o6x2WZEsFzIfsRbZhz9NTJXgMyH33hNAeZkwx5MjQir+3rin
sx8PRYN9i99tizGI4HvGHAHmktrtWHR66iV3m1j071+FW7Gqz6tWW64jI7dm6lHA
uvsbOW6NNsm3oVSFX7CJlUQIjoiWkGnuFLuW48RsilpMsDCxKX3wEJgx/c8Rx0Ty
nKuxqkWHjMwftSVoMwAVeSbrxgECyZMmlUokAx1Ecg6EQ8UBcQIQnS1jzdnoTsGc
+FEjbwFI5WC8uf44W6LiXBfex+ZKmhjI3QfAgCRFOdZ8IqM3KAMd3lF39xyObSHf
qyfDw8A/Om1EDrUP0MVicfUv7Ksrtqa9Gky7/YIQhY1Oxau4KaNr+rIT6efcxrWe
LFGgFkZtDFn9iB3pVtcnR9NNHiB5ESpyEk9opq3GnCHktVYnzgFlfveQfO9oX1TT
ITC8eJsHsQVKCXrTwY40gMHIXW0VVFuY3cWmoEPk0nuNaOs9/T4uyKLCI5/HhTlg
9W42yLGiZYSCFcP1FMOOll2XmkpiIMQBqrgL2Udh3vLzrNez5ALzcqmgQ/pJoiyx
jh62/tKFBiD5atwvsR4fxNzkd44aiBmj9RPliTNg1S3vsUN5sErwjtukZE5WE00i
d17C4vxJMI5PLuQATAaEV+jyTruMoEv+9XLHz7SRx84mK5NRC0wCMYNXPBfN+trT
WoseeZU+/eOketQ/dRHxH2cbmEAHzTabxJwFl8mbTcMziKGJteqFboU9VOG5eFGK
LVOykk7o1d709C2MQ5Ob5oYSyRYHk7ks30jAyA22Kdcx4VMTTGUv95SNttyN+cjJ
Cyhi5KkneFN4bfut2barkvoxmbscfR67J3iXYYoVaCdKE5pH6r64yOHUlpaFj9vn
WkoFr9M/KodTzK6ngWEV7LAkhzdV2o4hr+/DUmItsh3TUXOa4tLQoZMqgwfMF6fU
VsRgLaPs0G7TDymjw6hJaP/x1yKmnsPqLkG4az5Ak/grK/u4WhPw0+m2pdUKfWHi
aA3gsYkyxXsCZxGKLtIGD2FbL84MuHJw+43aEZQ3tmbo0nMgoKOSDtixbHQ8JUMs
TIFUKYqQYQ/nNeGvDD3dUyiJHkhfhmOaBKOvuZNR9b6NhlviSQSplSmB9x1iH+Pr
8aknb8KIoFSG8oyt0l3PLP38UtQbbem7qAgpu9OMcM2LL93FcxwrUArpNVFqgkG3
+O8FLYLzcut+2w9e+oxJB/nhjI5iVYI2oO76SbBYrtpXY2PiJMnx6/jXrQo6fM2A
U+KrFcYjIhKqJBSWS/qXwp+CF9Sq2Y0jmnBC1VFTiF4SapcLvBFTFjg9Bt3bMi4/
lL2Xrj2k4ZJNwI9BIkGrREMJ0cqAB7tpl7doHIM/+dVm7B3nn+VZr4WBYiJXVERC
kk/M812QP/dnV22BCioax4Xpfrd7jcAD8t78C1HVq9gXwmGEBEIjZjciH4Cj8l+P
Y0WToX3bE534d86QvMNNh8eNQDL7GywzdBBNnuaxG8StvxqytDuWV7uwk45mb7vO
Ip2Hb28WONHui+7N7Cb5xqS/tbtysFOg1vrLQZvFoDL2gPRkZq3QemeWNOOKuLAh
CodD5tMbeSXXSvUX3m8GQv32tgOQCi3MH/r58HgyWxe4ogvmdy9JUPLxrac3D+EP
K5QQm2jw8dtXIzKLeYzGmDWOkXcRqUGlbrbUaRAc6lrqE5NP19j6DG0IyPwwp4Ld
bi7DaWc3+xAWYwozRl6HOn2/UFs+NVlm4Wy+N0sxm/DE+23qdocyKpOYeMpZTKBH
mMBn/4H4Zf+kh6rMiW6BJjZF71nvEEF2qW8L3Ote7n20chKHzx6iIJK7gLMewxuu
sGCdR42NovypDyv60sZ5Jn3UI1cjk6PJUcJ7PmViyfMjZFImVGO9EgYd5j2dzHZa
KFUctVLYOQDWDDUS0AA37YNIyS9xt1FMHRn0zIjv4Me0SteHlLRf5lttU4v4qY0/
l5fwojD6MD70+zIs8pSyQq8jc+bVj2Oj5iTTduFXSek34n5vHndD6gISfjBSCHAk
bFb+94Y7pAX0m9REKj0JhVQvTode5PdgMm5rxyEV8eEjCdvxVnqlh8veycvlExqp
B3sHvn9cFPnsp9ETzNQklm7bY7WoEruHIp47uXIq6VYr5kv/qd3Xov7cIE/VTUoh
/2QRUyUxRSqlBOIg5uqx9pHwtOo4OoAkG6+qri0FeUzyds4w7pM8eDKqKZdtM5NR
7iLQlBT/TTdQasA+7D/BQajV1OPTwMEZSRPnyTOJndv5BLXYJG+f0/5AnzXYxuTx
hmPHOWDrsoJ4fXrejr1mXo9r1pZi8Tl0bsGT+Pg4EWgWhAqTsx7H1D7KgLDKq5xh
Re8sf+7EUBCDY3zRr12HYAyPzYF1s+FqcvC0B5QCPLJPPh8kNT8dbuvQNU0C4fPw
i9/VcfDDzDKedN2U7p2LmMmUpkz8L9BJ4wv5EPr44U8RTqKtemm8aL0CJ++eGtyx
HZ5hwW5cIxDK9TI7og2jfg6xbWt91IDzT31nE0WgEr8RQbNA3lAPhZyZc8JOzzxo
+ddIWpvS8b/y5PVoWRfaj2eNwe2I2GnbwtSSsCfZYuCEucUv5virs0nV0+t52mUa
d2H5NklUN4Cp4PKJCMMFE60Jf/ItqxG8GhWKG0WMwYompphHCz/8BmES/CTZ2V7S
00ka3GtZhP+Tu3xaN/K69ftzCXuyuPbF58OVe3GD6BczhqRrhSxzRycJVrtsAQXk
RtkiEs99s+TSBn8NXnxk82tU+EhkM3uLioYv6uUxw6zk4AqM3SWGLx9tc6NZalsC
pG3aXDneyCwbU/oE4Z32JN5f8R6uwXqCkS5uuaBeprPSMiLH47tVY0hL01fuBcU9
8ZsHeXOklxwOwFxG/nEU0nugr+2aRl+lOe14LZmufTTjQnkeFcQ6BUKQgtOJoi6Y
8tAe5TvYRMtVOE6/5qK85ME6DNV19LVsYfyl226vH4yZD4tBQbNWMkgCkHAPBE/t
jAWhAY1A1Im+/Js1xVVJNN0pal8T0n5dLfn0wyo6vb3CPH04XeBABXqw0JtzxpDe
71MhS1lR/KmPShDYRfeRkMfEXXTlCI3itGOeJNqsObmW+g5lljQCA5FOISrUhybK
Cpwl9Kp/eSbM6S72/HZu8gPTVZ6rKhHJx5Q+tW2dGFT11Khxtg+hypfn7haXP4Cq
c6IdKECybTVhwNM53zVaX+dWpyiWto6iBkRucvG3g0g8eztcJfD6YTUnkpTInzTd
wfOWZROAUiiQbhfK3vGxayHglpRUl/hPPF4RP0AhNd4CDy7J7Ria9s6+fVSQ86g+
9pda7QNia3rxthZvH9viq9GoEDkOk76+wdLqTypujr0aX5RpLZD/cOnVdaI+7fip
F3mQlyItAxkrFlPFhteM/4Y+uDIkRq2WG6LA/k3bqkRVQM0pBR9tWnyfSwTdh+jN
NdrRIvmpbTJszQZCewQIFrQaf2+kaLwc5fHZ9p4z5+xSs5uKutaWV4ZzR8G0dqX1
Tb2qXYtXZoX/IYfEcalioeykPUkd0qg2Ta8kZcnFkOrz6mnhzcYEe+VTGKvGsYe3
lxlV1vFBjD1w0+YRP3mTEGBbfk4qAJ2igx2zbW3sumwxDQywSHVLEIX5aQgKdZ6O
Xw5E1FO5xC9jp+l8+My5jCBEWqWckJVuJryqQ51R+OasEITLJzAOMmEAObZ2cRBK
tixT4qmKG82FyYHZtaIdK01Em3TWn4PT0dFQhdfJUTTiZT1bq5Hn/kbcZmx1M3wN
LTmrD4Tz0ELthG1zaXFSI7nYR4LIgFnEM4AM7WWSvcg4vMXw9HFJz7L2WMq3ceYb
kBuoBnhEXn03MEsyaLzGcw1n2rua88QWEzGnBXkuzpKkLm21AGBEbIBPrGcg4Mo+
74oa28xWCpp/3MTWx5qwREAJW0cPWYpM7bQtIINSiIhSbuov0qw5LPHHZFR663Al
rhVj9CnVdauMhiEgeRdqTU+j1oCGKzMwguEYeF3YnkFVno76PXFn0zh29Hfn1EHB
OOcLbkXY3U8f5ZDvv/gwMkW7YuH2Cat7LmeokHxUOGf/s11fhCRm2hKBvut5iOH2
bfgsN7xiyl7kpfd+T03/GkTq1VSi55DgrJ8EheiCSItNGdsAb8EpZO5rHBPEQA9O
P7xA4GFdUETvKLZwrvP4X0ySjaKfPDmZD5OpL33cBI8Q7IyECul6H9aZ9o8hdQww
oWlPuVcyp/TiKusNQVev8Bff/+yNAE/uRGlUx9fINL2zNlUT1AJGpIr6PC9/jSLF
Y/sLd2SjtbT9fM2n1OFny3X0xfU6ONKWDK+XJPOVqbsJQm0ttKtWx8AZLFlYTBEn
fBvkmVq0EMFmRNW0T+jO4tEadHDgLVEp0DkbXaGPipeTcNR9Hgj6DoAEgyC0eMC7
D7LCygQFjErnrH4EM0TQr+h/TRReFoJP0WeCveihRIsqrCA3qT3LMt9qe9fDb0bS
dBNjFGtw+kA9gezO7duIXgSa4rCdcbe1PmbQ7bEf2O5SuKabwbAYTq3iu6PLMDdL
C8iYo9FyU1b9JO6pkEg4pATOz+2OJgn1lptkNh4Nvr7cD8IqG9PV+DUI1Exx2YMl
OkjXuswMQFNvGN3fS0/TXlysuRJxq64IpXIBu8iJ/WJt81Td1SdqeqyjrBmYYVVi
sB18otDdXwMkIxEiUVJaoGBSvfnbFrVHDCmdb25yCpj7BitmKHDB/U3lmhadEpWW
I81Fq7DCYR2cvgUhIWtFp9x9PKKar9uKps2QaXD0P9l3U48lP8BahHkZ+oLwqAtU
im1jUABEs+LIscEGUlm4XFDafx5XKkV7Yeo1gIvJSZEt/3AxttYRkvGO5L3NLEDj
Lut7Ufqph4jWsxAFp57byIPzF0yeveho/X46sMNWUl4bQEKMWsY1m/wLbjqVgFJI
+61VTXZefbkyQGdHXHVS6kHUWN3WkRMxrWgKx2GFCumqeI6HqQEgf7hOHddARPD3
/KfT8kIbUBUFtvNtlFISy0uObiiZW3UXVKVWVBRu1ib6crbsFPtjnV2qOl4ua4s5
SbW37LB9KRF/oG135gOoxIGwvkH3eW8OqCo2pw6uCG8Xd7xqLldWGmixKMuEH2Nh
r6gjG5JGzcAYsSjV70GdCpR4P7bKx4GCoSVkTcNF4t6IdeuiuR0JSbhTu1+FwV8R
AOHQJrQEHMpG1JjK2xAx2BNpx7Jns5403BITN3Kme1aL+xzlB54WpzbVtvpT2xOZ
oHwmYsv7qyByeMgKPmmBxzcXs7te9SThe85ZdaaIruHMghD+QOaqFTUy+iUHQDo4
EBRHiNBWV2qBds0DCQXJbHREm/UYIC4N2+NM0Rm7/5YrzA/YT0i8pG6gl8w4ehs2
QQWPXO9zIdgVLMj623NaaLWlnO9BV4Eac/p/kBvFh/I0XXwoLKQeI+2NzWP9uit4
oZLTjzQSyI7EYQBb4nef/Htlw0fTPdaHV7yBf/BnrlsnrbI5LEbPbfeaVuoSJswr
LE31+h5uvv+dbu81PmQm1NhTW2OjIr612L8cxxbTK7EPsis6ONb/D3HJQGdWAECx
2i/H8XohGuKkYNEOcH/hUUE+Xqe0iWQgEub28Z+jAc/miDl6tp0vfdeTasxYQy65
DJ8Dv6q5OrUNsvWYDvRb5sx6NO30Rkokj/4Myqpc65R3clBcMwtXeHmf5slj7j5U
sKiC66tcEpLoA/9ycgzMJ37GJcoHg1aDS53xzinUAkx2C7r5eMxArcUb3tm0R3aB
ccq34sS7aQEG0rKwpOn+EsKf1oOHqoyx8/tgIaloIy4hRWDrHWmR0EMP88K2De7Z
JjR4fl848xWpGWvFLjr4L7zdsq64TF+7M1TO/I+uQso74MCUQj8sp5ZGbWznq6wF
JqiqL1wPHSELThAQmLKeei7NHzGjUMv/oxcmmD+6JgkVfm5pC4NZwq449QWYH79O
QJJ+bmA7xo/TvutSAHm/bfqDRca3fY4jHwxT8mFYdUBMzL67BP0P2XIAzJZGL/Ft
1SufYK4xqIUxxACkuCIe6YEh2Z88ZNShge80tO7N5t+HTugrYFUK3GCzJGbZ9Dop
UII1r+IXyLWE9gFsxquWt5k2YSwzRtUNuUR/GS/2alDNE994H+4PB3Mx2J8wlJXa
v0o53WOUsVsK2mvf/nHS/wB1/tBcc5kba1K5QOHJlRKzTWjAbm7TURVdxL6f0sA6
YXSUK4rD/UZccds5gdmBOnvM19v6ugRAMEZCL4WDUDxKxb18WpeHErKwIw2w8STc
2kw8TrN0YizfsfbE9KZDmggWme5W5O1j9wJ48xeYX366a1ba9RkvkM4RCbOZmjvV
BWDAdkZmztwGerGembPRnYn002qKGOSddKNZiFtMhIfw0ZWVt3HQlTOm9t5mFVlx
faxpL6FfUXbOnycjY9DfSek3jQGLp71bbIj/bCM4HkFobtkwzwirQ6TfjytlbHol
TRWlCTnEZrTVynT793etxqiPBqbpdQAR29x3v9r/VPIsQDTBDlTVA6/0IQYNZlTw
6B8UxUcnJditvNbzAnzMYCE7MWZ6I1iWR5FnY4OwSfPsfVyOTXFGeb7eoZHiIAtw
PYVuQjTz0P8cmrKSQs74RUlbR93zoyNoAJUuC2NNbyJMiojYzsgQ25n+hBWmhNka
SwTgTwaxubgoj8gY/VH8Vxx9V8irJI0ExXf888g3EkDaktY7rsY2ofmdywc9Oe+E
GxNTRMY3IGcN6k/H3/T0mn/HWojAXORHsxsKjtlBFpbstRAD6uc9kmk4wfV/mvnG
xJME4aFlCasH5he1kGCqI7Mkf8qOl+7NluYITjM6cddXBnP8p0kqLxMsVhvcRn1Y
54VZdFC7WfwDiGU1OOAAsjp+ZRAWgSrsX5aUO7cYHRjoAU487gqsJ+q3HJW7y0El
DUkBdlqLEa0HSjT1SqwGaXSlZyfMzL7nS5/nF6qKXerANaA9m2LzyfQUaQq+b1MH
nkm0Iv9WtrJ0tDoAlF6a9Kvj7c/i/Oh65zXI+aobwBQVMYtMV1/zZQp362q8pxCr
dINVkxT+PgA7w2ehbcPCN9gLo4w3fw9COy2N/1+bKp2ww//xdzpWU3viWYH6/EbP
65cZeRiFhDVoA4c7f34we3XBq7WvAAXTrQ4CLJsr6V3iYF1aEHH1Kfkcn80VFNKl
xcQTQB4L/5kd04o5U41/bYFoIUPlU/8bBFH7Uh5wOjyVCTll1zcq6/F5VetLbJzj
hSFxa7eGpSUrCHe95pPYYMR6RS5RpBpcbZpmqY98XKGqfFHt1Q0x0Vitw5v6m+zI
lXBEkZCjpKT1LY13wdbTcJBlwi/hnwqcHeTNrdTmi8Iw4YkdUpWOiXC3HHPlOMDJ
LpWNLBf854E6EkGbT7c+YiBrSOTdqJaB9b0n//X54OPBgyl/EtbsH+oDnxIkD1Kq
sRAmfpYPRpsL206biNuVVz3fUDboSbwkwmyYPddUMsyJk+wg0NTCdMZqWmbLVuGC
LOO2Ht1rfbIMQF96rhIirxgb0cxPfP8TTak7qQqMpcfBMe7d1/gQ3XDuTho4jEUY
HAo6EAMukjDG34i47r4/iSrOM1QKzY61Yk/8jMoDhlZw4iKZKgFsdisIZDFy66K/
roT0iyzvGbFs9Y2Jo5Rgw8WC9eWrGeEzdbS1yxbTyEtusDAX1lvNUZLdGk1wusfY
jiafT7J/vOBRb0mixo73JVw65i1NbGQDIZ7er30feCQbEWZuaYRMeuVN/PjGZqxJ
ne4YGT95TR7sG/vJYkvj2NFzQhraIicsq8Ap27ZVz5GAGiDIXwGw9MTW1Vwa334T
zF5sJ3u/Y3yaO2FoQ/qowPMh0RHbfMclVWVe+Li8YEZyM80ydxjbHfO46dmFT+/i
9mha0NPgblgbY+I1vRVTiGLJJ2k2wSsNPWKAPi9cOjovXxH+himPRSMDikaHh/y4
jRzXzzfPXjvmNhk7KW9IaXxlXuh4RmjLAmBlKJrR+sSmhxktggo0Y2gRxgI4aS8N
oP85FKoY+9plf/SuqGg/+NdDZQ71YmqOo231ijgJTA/Pu1PE+zHvPGDIRouHOeMJ
srNK1E+SDzK/1yH7y3yNcbdv7oa54pBrvAmlAtkJaF29L2+/13kg4kYirwr2hh6N
TQHqwl3j2u85XRMQZ9F/NMVqO1jX3dlMh19VcS0giVOSCerLodIlvUeeeGtm8WAd
esOKchgHQeVUABc3IgkSFLuMCMTYiGkui/GQdW4frS8syECJ67qprN6y9cXnJfjp
xVrQkbWyqaI956zW6K5t+G74CF/sBPFK+Iib58bP0vYFxYW87mdS72XCMd5BcsGJ
u/6ebGhjhCHS8SgyIOQioM7TSOBVdu+uPgwMMm8rjEFBuleFjV/hBXa1W9/rjRhL
wMRsiJwtoLcII6JMXLFD8uU4KMfdoc0ad9yQKWDuh95bK0bcCaNcmlaFbfyMF8Jq
imdIVzcyNavSMErunCruxfb4NKsmNIT77z3KJov/k0UIq9nPEuP0iJjvQC7pp1lV
rKDQe60JRpx5WKOE+TFydJG5MAxvN9Htaexp2Q8emOoPniCGnyuTzu55ujzY4eJH
cs/CsQ2VP5FG5GWO29CU0XneDbfos+9DNwWUFfg0ebiu/5y+X1ifd39yRvl3dKGG
FdaPWLvmk0DJ2CagJBaym4EcgT0kQJQ1VdsQeqAfb8F+Zi8kiV2bkYssMVvA4kYX
nqEH/np9SMlK2wz9504y6OKA5rZV+Z2BRcoQnlfdABxTlwBptpKfzWV/BNSUuVNS
qIX8hcz3z8jVyVlz9sKEuhduH3nGWUYqAUXtOzop5RF+c/2DHdRBFs1gKLELLn/q
FNXZX3rlWtDPWweglNBqqCbShj86qlJEwIE584kQSUzlPL5w82Bcw3/zI1/dFqLH
X6pInJarK/Y6k60D6M7KydF1tXyPD6IJdLtaU3uOWIqBra4XyNnOOu1rRSoHbs0q
lEgV22sMr1RKw+5KyWQop20oR0wnaY01WVqUld8atMSE+bvriXI01Sk3wRZeM8zi
iIiDALCD+4bH8mWY7hQrZloYr15RxCxMmgSgGooBc5i6zJ2cZyhxlMsvLPt1y5aq
l62JChujOQ9/xggkSCKnd/QyVErZ/3Ts6EjoyGMGLlIq4HyTg5KUFn6b/gYSXXdf
jhjgWlnqldFhORe0hGcboTt77JokZ66d4a5/95V+2goKyIqIa/OIHCiy2T3p7F+8
7ie8lSwa6PgLIyTfHh/AMYcRo3jQW30CQRePYKisrsArZSX2QfGoHsQUoJDVa5S5
xQ3emQKvCkZwuwCGW3f2BE5t/UyEt8++aN7P6vD8bi9luV7TXchbCRd945oz1hPv
hmrRxaftyT7GSyxdfKaL6ZkPPuF7XmvA3FNTapeJeXRGyazA4fL2sa9LvoNMNEax
9iapc2WuTD4+igGsGYDdTVp0O5sHY5TsUNvHsbLNCKPLUtBF6m8iLzgbxOj9EUra
rBmMcQFQQHiH/FUaKX+qba43NoN/+yFVECNgGE15BylffmZsiAz1dpPnSnBBED4c
nRrESen8COLH8AvBIlUtfHseullCtOJ0Da3XZPDuoiuxwiNP3CYRpmDZ+dq4LuZj
dl4ztn4qwdUp3uTvsuE4CWmX1rkk8c4qMhmlviYnlzPk35YsdK7vgw1++npD/p30
LA+rOr4cy9TJE1hRShM3RLbV2X6ZSL8f590D/XaJa7aafIhyHlXrk+kii/JbiJgl
1azF51r2Kt9OPMIPfmIE+tYxy8fe/mNwkHNKdM+XtgSqtnyBYil2SIKt0PAgMf8B
qom73SWrFiv2BTILwccQdvtpqBCtp0RAMiCT39esHbMsIXKJm3vjz4ZrC15WiJPO
Qte8RTJaQCg+6xci9Tf87pDeM5xYnFvpDvLU7lOWcIbAk/p+r3xvK0HkSMX1OTXL
d0AjnsaIWxqUEDS3Zcj9bQucjWKY5D7bsr4/37FtnyzoNTnfOnBkrHX9kMgbmkHE
qBjzxL3v4gWH1bow+ZzoA6CRoF6eQgiXwx8uC/0nJdKxvgIGGhgvAtsCprHyl22k
bwO9BuCejj6g382iRD54dZ/PTQ8HENQERIRjASsN1QosY+fb4Oy57ErQHVpuXm0K
xiEFxq9MiKghBOHbFKnrWoIf35KQvfO9b210XTNmsWaOGEpCDd8rdf+b3Pxtmc5a
pO866U0yR+rhLL3xqK/Ga3AoRi53peUZaUT/nLzj6JJM0/6xWDAPyCIRWDq1AC9I
dkMajzGEbd9p/BCQh9Nxy2SQtDYAGnlJO57JxshaD1iPSJDjXrZpT/8CTYHtAZ55
daBib3pyN4KzXr5BLQ5zbOPLV0Rrtfw9fNTugeb1ffwvtfUHLtOsshcM7TBdFWFQ
R6UTl/OU1AvvUjrAeGBJ8H1hNJjPbIskHfiWIS4idSilDtHXpyOjQP6CSX/iDal7
QzAoihO85msGAO2PcmO2vmroxlZGREPK4HuFMmXXw+Fj10YbWrAPCeWOQedP9C4V
NxZjOW1gkf9DMTkyf49ffF/eK0pPhv0PgyISPFrOwR38IW3FRLkTlL1L8ho/NKoT
qISOwaGmZs9bawVY7aCHCz2shFXRpfNMkvKxpCMUm3kCTnTpK7ZAB1a/Yq0Qa5YX
d0Kz9AnzyUt24XLMJ7tpaOlAuhVvcsm5vvzemYEhEwm108VAbdJgKeLrv0yQb4aL
kBQdGkurCfMfYWVqFdAoXXkUWpjq95fEfvsCz8gd7ISILGolTJe4T5pIJS0wIggo
piGySduVXlrMsPajLhlt9FEkk50IzSzA5ppipLPIRbR6bD0z9YxqL6MjFVE//Owa
cXFShYm74VWnc2347N01xkP/pqc3MTMwyygHC/72vc91tZ1xI2VK4L+mZDrnHcpE
lac4kCTTyKd1xXcT9rXPBHcQTXoZ54pnbjnIGrspeTnQjbsxiAoGPAkKrGQuc5Kx
C5kBOgizhqcZ8BtyTktolO5WM3HVxYZPFuWM4hkkpI2DO2EgvVIBE1PXbOsRoh8+
YwxRZDoACPZwiSCXMvFzhHXWWROnh5NSTzwJd9v9KKd5XanhGoYACk6dMqXRDhYC
gkqAI47uGd2Q+02pQF4KlcmrvjI4YOkCKrWkqrziKkmi6yO2F0xUh14XH6BtAGmz
uJaGQ9tHp2YODr5CERxabil9tP4Dzj6/MfNTS2z5vO9JoOoqzW3ey/T1cZxvArl8
NsN6tVO/OCA/gUpTIvuJj73KQkDIkxoyVzYsdIvaFJQ38jFb+bcWL9NZjO6Ikw2o
mZpk5b9BsvCYKhRy0ABkP7hZOf7FUlW7vFJwYBENhkgXkNS63ilUmPf8zqx5zb/M
6yHx2PtCfivwWVQrgnw7FD+zBF6HzI0m46Wmi5guFKsPzPlUUW3BTQcwZW9FgXT+
qkZfHNppZj8m1ycQj4K6+kt910LfVmBnZ8Nvf/E5Wm68RBCrBOOuN8uMnDK4Fmeu
4gzcs07V8LRv+uqSN+y+mAXDZH+PfOEdAGfLhcceBK6YYGAAx0+g+l52wqLTWPLw
lyoFGI6Gk1J7qsx5dPGkycOp281+lMn22k2ojFAS3R9bp/hJuO4JPerrQkXwVf0/
g3gaK7VJ8EG4LlW99GEKXQ5lShXw5Li3jon8vnQ/S/vsZKrI5vNKfomoN8u02mjP
DL/xg7u+1tDisw4xAleCTTsslxX8nELSAvu4MdrC2kYhki6eM4MAGV41K1GQkULg
T8gnVbcrbyCVsQBrQOVgBxqFYyY6oZ379H2uj40cqaES9oxHh+qIejaoH4pzpL67
Crgj4FRxmxMVzRl4YExpRIbMaDEVW2sAkeMiBi6PcyVEsxYXfF2g5Bdq7UTNbzhE
irkwNhByHNzSGkudvKBfbe3MgbadVYFEM/gZBEfDartze8vKjTAoJyfJHLB5JTH9
jXB1jcnG4rfz/fRDZOPu5wFfF5bcvjyIa7yobT4UvDztnIFM8PgLlqMnz3gugZiz
NpesiqdnWMvH5F7bF6yqNr6Y5KYhzNAbT33B9hnvh8cqnuMRfKTe0yQ3klHnImt1
RryJUE8mTE5tM51ZOWhTd2TP4yLe4wn36ENR2KvJASWnf486bTg2JbhoWdbZ9EnE
Rw6ZaS2d3s6urBSumoFu3tym6I8T0cdX/tnfg4//AzURLxOpfxcAzErWwwib9k2W
ianaDMOumh8R3mKn0fpHhL5znnVOHjjqQpF0eTnOf5yPCIx05ZPuC1gb8XVDs1qX
AKp3VTckV0PAVUSdVMsCp43BMOT4QDDiyjcsoGI323pMkpHJ36DDMute5oVKbIuA
3b7HBJky4++x9iHNmIHsOBNPdyf6/P7NKDB+MHyrs1+b+FVcCrwH01spaowS3OGI
MBulUx/cDx0z2N1STyIT3x4hbrfaU5Vpw3tMkRCsNtMuj4JvtVPWDq2XQx86J8I3
YVZCpDpbE0RkaYVL4urRGNskJL5knXzl74K68i7zwMTZwvDOSrl+0WhqijhNunUE
zL5T05njhbLPyJ5u5QQlL1EkhQqxBcmuAwoayI0zD8evAflfnfTcQ1emFgxbfZvX
HebNSfY9S8/BSIgfLb7RTmOdwR9jIfz7/n2hmsRhWba+2D9bggA+aj1wixMi55Xv
Z5gwp3voc40Bi3LzHs64m9TVV/iKgOpc/WHvAVNc8yGrfDMInx69a5Qsl4Z4exUz
MTZrv0VhPUhZSGe97tCjriKIp3FLkr8WvoFV0quf71DAopAWjsWDnTbCtBnP4c8J
4+15hWDK2fPfL4Lo+K3c8uC9dZBkqZa0sZUDmv+ZqUngQ+gSiT5rr49+6kZZk2l7
DNW+WV4iUbELCOtpckXv2mqY1SrFYY+drdIwSv7k8ZcT6FztoDrT4sLLneBs+RS8
D5skNS6kH0Z8I/h9gPeasyr12mCLXVrCFg0alnWhYH6eDeFU9yBC5ORAoBsunsDG
kLrY+5fu2fTMTx46df3Mvfyz4Y167QcnhDixlq+/BYxQm5OuyCLAGxUlkcbmTBjY
ajYlA0L5G4Z6xAxY0x52S8k2MW9KvVLPbjhtUolc5Tj/hPDowSTifavMhYXzubbI
xgH//w7RezUTTVikgtZ2oVmqv3AtyCkIWHKTb4LZXgxzqNQMcit2A5t+RC8Wi0Q4
W/JQUW4EPTi8zvazHygznAAcjo1wFBq8PkSxQxXBDG0zDUHxWsQyh2LFEtY+AcRJ
a8V0VT3wRN5jrq0kfxEiP21fiBAWgcBSczJra3hcOaZ6xj+0f4fyawnaSVMezhu/
ysh7yTth7wq4J1hesQ1viQOKoeQrjozOFOR3LaKbUQPPvF2uw0T7DhTmCMsBYCKx
YV/9a264yFuHkYvxVRILny8D5Au5FC66zLMgqBzD5kPmu4peJPx0lvo81fM9Eyek
u81vZHRvFfIw4aKafA80wQUaclwjnwSwvyOMNEV80lczRqPKZ2oLlRZu2Ehg+Xcw
N742iswGPZ7TIsxnkHcN2vF+VBCSl53SWvFjfTZDCm2jwqM8/tR/rkL/92B6YTWV
wZN9u87q5c9A9Dn0Mn1tlRr9GfTvOrSbep30SGeIWBtK6O4OiQI7zS6Lw5s3BD+W
yO0E3QmJQIJPFWWKM7snqF4Pg4OjqxEdXv0GdGWXo7KtLRuFPtu0OUZFq3mt15f+
juzyY5Wtou/6tqlPcUr/AGzEUWHI6xRFhYZbA2/wHchfEwksL3i7y4DcZjjnCdVO
cIPpSxklcSJwWNRZ0usBOptFI2CHjPw4lUf5X65s9kfN6mFQNvjLUNuW7oW5MjoC
2DrhXlQ4wU8fpvoXJ9NBUrBtFcW8Zcvof/dmzDCHHZ+XECNXwspQG3wi3kAiKkBB
7/74rSEr4T2v3Ic76oKTTkggQcVY+LcUlWZU+gJD5mAfmvuUVludXMveTCau0mMV
RYuhy5Yr8/vc+iFvNehrZjs8W8eElBG3FH3c7INBU0PG73iHCnMtSer5eIn6dfTU
7Fiq6dbYp0LaQtUUsKuVflOp1EkQZOKEtqe9BmBeqtwI8j3nVEeAiF9/KRMe/VqP
FOA300+wVqKHveNiiBNsjgWl7XS0PuLr0esJtRl3Zm/CtQRRfF413OgLL2rFNevU
SgKRew9aLR/QhCc4knHVk5HD+cut3+RW1V/SWHKFygJBkVPIkO4poLkkTYkuUlJn
7f2cbuyItkacSM9VeUbBer02rxpgU4346SxCdPAobfl9y4S9/8vDZYfUyOZ8MFIk
gPMSx94mCu+F0clnjaRIAvXQohbYh1K+oMSjZwMygwk9ebWOcjJO0HdnZ+gNia6W
UuAJqIolkFOZRkct7jfxryQP2r5AW5yrZeDf4WOGlAgX+e1Q0efR1V+SEMceoUZp
oLYD6/kr1Lw54+SNt8RG4EtFw/N/D1MrcW4yW5ITqz11TmWX2f/jGCHjzUwWwOSz
Dop0y6V9NnJ2NzL9rxVD9n4Vy7o3xgHeE9A8bBDBSEChzKTl29sDpyrx+4Ln6Yuo
0Kuqgpk0KSwr+PzRZgrtNpz14sC3SebA5we1ivG6QBl7ag92vXpDwqTGwhcSHvI8
IJiEfSMTxsrVys4DZBp8LICxhSuNdhBOHj6wA/xDrCShO2oWgtpdv4A6H/VnVNEQ
rw0wIVlOH5j0lCJ9DuHLVPhaxbgmo/vJhJMG24xMMJYmJQ1RLIug7ILen2lGdIqw
BJpoY3uBGky+A04OTYfA3ISoHQ4DzqJp3410FFAErdvLLtyoz4DVsN7bDRPPZPmP
vXsDw95rVevo9sIqGWbTDZv5Z+M/1Q+j9g7t2i+eMN0puAlrn3JqIr3eJT/LD1n6
9AXOH+PdUYXKVS+9USB7zC4fyHJaTVlWFCNXT/4lVkYmydPUPKXEDhLyDecDcMxT
MPZtEy5KBdglSadAOL0tikp5fjp/lDR9mEhCPw124Q5DNwMrLOc09bTrxQY0FMqq
9O0QacePJS+0FxcF+rFrcUSpehKeQyQ7EZCq4UDDm41KF8H/311bfEoMciM/IVF3
V1/7h2NjXCoAxvKcdrykOEuotQFVNMh+dhFkRp51n9jdMybqvJrR3UcNxqx4rbQw
Vwiq8f9YPytFyeLNZ78rDtRzKvKyC5MyF0MQnInKJvnvuRx4qn1JjdzjSmLk0WfR
gSL4f482MILUSmcI6k6k//MavWm6h8vPCovMo/Vsd2xlNTCwwqK6qTDg0Mph33OQ
WkBNr5VdELauCDe+LLawW/6Mv8wVd7Z09v26vEVsijoTnCexQMBrqo3EFWhjfsA6
qkEsq0HK/rYgWgNjI60gd15T31OdYivuuJOxq5Kcbz/sfniSHBYcXNANSysQGsuk
Dpy75qyWSw7PW4/czn4r23dFosM52U0gOZB7TqbkHXOtgAALxpCR+kcSZC4PNBKL
uKFQicHim0hYmyyaPLkTn9KBbyI7ee9lFW2SaO4qS+rYjRNyp/M4II+uOnwQroDW
Wleio+YhG8NL+7Qq473VsdTxA0nxmAH3Sjfu3BgN5b7gEFPwaxbaxgfDwqh0vJuA
Li1sFp9nPcNqU+Bmd/omnZqfB+aCx+zXRC/bezQgehr8D7X1SHPVtRlP7pOwRkiY
iap3QE/QgH1XaG8PGcFOJ2h9HOrZLpkHcfDimjV2XRjbUU8/uSq/zO4rOO9aY1Aa
M7kfpL7VaHkkPUMxntWpg1I/GNjIHq60RI9uIKOFDb+gWo/jtrekC7up2MlwA5Ey
KZWnnQTVDU7iIlP1jLXn+aLg1qZLulL4kbezt5a2aLialpvc2Ey/Vk9yx6FMeEFK
DpeDS/AZlzLbgMJ8QCNfnX5sZvMOv/uY1CuzHl8S2zi4lqtN7HLwdYEryUtE2xZi
TQ9KCF3EqmIr+5Xyub87vC0h8XK76qRl881w7Pasd+2oHtn4VBQjwvHsDv5XNLXi
zSWuU6n1VBP7EvykwEaNT75MAO1dlv9XcCy0HjLR+J0rLl/dFHzip8KTm6r0euk/
oz37OvSYrIuR4+kMmhMUQiVy09Zxqe25oO9HRfUWGyMKSyblcYNtOTSvqiwzDE1h
DGQYiUEh//iRQk9gP5UyVOkgoDMhHbZ1g3Wmyd2vC6VWhT8GxDbQcSidg26dLNqI
N/zjpUfeLOFHFwIEOu/diNBDO9eIJekNkCKzZWc/UN31rIsBraB2KuFtFD4GRxI1
c3NQwBHWZv3/2w90WCkXNya3BG8n+K9+qEztD1kjgCo+27ZUpG0HpVzrK/T0szrO
b3bfbMZjpp7hHruzycTRmzppuKSqTwkKJS3Eg/LbvbDeJE44ejCxfAWygHUy9V1I
KuGksnXpXL5YJyHUmNlGjEYg6rsaeNBR/qFW22ONXzVrp6FIhccAtmhVEzUZ4T+Z
/XpISV2ea4unocXZJojgJrX22Kg39dIeO1yw8m8aVV7sUp7hF2GTmCmELxqontmQ
lMoVdih7py9cIQ48vox6Yym3chGY4Ajxj7vh1rx/9/ThhM0SJwU/TcRfn9jk1xS3
5Oa0i+ssf+iAfC9WJKojAAlJvw2Jy7uac1GgVkjlGB7rUk6Ubfak32lyeSjWCbPW
hoRBebocFWPuWsS4WvGYMsz46sFrKyC/pIMfVzBE0SUdbPFRhrbDtOSHXqlEibjh
z+nzXNhr8YQADwFoPZumk2kY+pmG5XLPhd7dAwA5xc/j0QTot2pilMFgEPJ4+Oqb
cdXZIvckXH/vMddcro264wON9jCNivYycjQTBLUF+Pw5JL+uDAtZjK/anEiAjNGy
ISznxro/wfiwKildoMxKtJK4u87IP1X5/fDQ32yCmoDqlPm8PV6vA7n73kFqN3It
4gdgf7T6pE6XjE0uB77NrWDXf/Hdm2vZXNwGVbKjxwn45xQ44JuXQeC9phZ2yaA2
iqm+Ak/VHb4PtdBdejZZuONxIaEsL5QTSveEGDgwqW1hCMQl2y761cSqGYX1dfXB
1wY167k7x1cV+uvSBv3GpwzCdUwADj6+fFaTZROPGhI+z027kTjPg3pvPlq/3na4
Xo0DY41aXZDL9puJafIbVU8hV7JDLSx29R8rfowra8v9fvi0un5hchu1x3dq+ZLg
BZjI7HZ2H/ra+MclAeqFB/99/IwXmD8rx2soCmcQvILNZSGF8Qoj4WWqrIB5xt7P
kpK+5EeZbSjXx2NX1uyLiGsP5hHI1tOQUU64YK1iVmsQhY7KxrHwQoOs8qDcrsSj
g/+67eGeZECK2EgZK5Qjqi9+t5PvjYYNEclEdGM3ldMNyAdPumrf/FlfxIsniVk7
ShAzLIGFass6ZMpwLfypQE1yts2CgPWDvgorYpUAZCYQzsDtjRXH5sCzmr/gIpBb
CN0yWo3w3HI43YaH3yg5i5Dgmf+Ogn1cOPLahcgCirptOEztHkTgHhegbOBFLrsy
0EfjIWn4ZfT97Rwre/S/EnXj+rLe0rPtMuhWLdolY5d6BW2/dzbQ4UBszyHVGlTg
SiXdW6MM56fapHlwDqDdY7QWH6g3an0ipD3klABIIrqpzSoUrMBd3aZ33LW13lsy
2aVo+KMCUIWuusnLEoPgIagqYd7xNgnvI21hdCL/hzw4GEUxdMOStKIjBHAlXIja
A3sd3Vs0JCti/ioR43lHGff+f8JArJcubKDg0Sy08WpiVashF4lN9tSWDXisr0RV
jOkjd/lotMcorP4SM/Aj9JW6x6fq2oe85oza+RvXCle3psGGUYbaKXQZ3e7c4GzG
RPuccfp8Ydj/SEZTXo2Cbd2HOsiqUgeBtbolCuJ9z5qKzCtTrp+1Jj0HnjoaIVAL
0RLY9GnM6YkVX73lGCPbUVEBHI28cDei72WDIFuWE7T8XWr5KqMH3pnGqEEkckuY
x/2HrsVB6cQTRsoKDERVfvku3XtIo8AwJq/fqh0xZh4CG/4t6A0qicfnlatiNfnX
n5X0PAhHBptJrSs3VAnskri0I4CTvc/uZw8mZ8hJ51yX3fUlfJjQleiXU+5IaerK
bsNdeFoM/FCIwuc/9RmukW2efdem2ueUg7uwkquJp0ZwhLvZRwpoSK7Bsgmxlfgm
NZUB6LqZh6RHmG++YZhfhllQnA3I6smyjhfarVpJ2wIMtEvJfenl7tQrSZFxHq3S
zyw38xvQBvYsz++FzXAXlX8zEFrL6NDy+QmwyUmO4tCjdwCdqW22UUBVXfDGy2JJ
5iqpDsSTgSgbT4psmc6z5uKfnseOrVuZDuFOnXI6F3VTHpSZ69qaM+0vFyaC/YN7
QjLe/A2YOnGEpEeeAN2VxVWOT0XIWGGvG7zlNiLMhkJsxbf/cyiB1kKfjPnTKR+n
NgJnopiTOVpEBHqV5REZolqRyu4DmXYD/EKl8GKBwolPk6DmLqHZY8nBf6VIfDwg
duBiHVMnpr69xC8FCEon7kQC31R4Uz97W1IT2Ww05H/hR/hXjuJqW87jR2ftX0QN
w4DQlUbkBpHrTbaRlKLKQvKBWjGUNGBcfL952AvJE6Szm+Kt1vbPTrGx88nRycYT
+oNeZRkjZGLwgjKl9YO+AoBOLXZL/Kmmfi+ZKpdHlCHxx7lOYBLwI3nSqhxis+z6
XzR+RcgNH3iHQ4FWlB2LBd5TBKp+3bodiEnS6ITIKFmf4OrLVaBH0YG8YpiDWCDh
70aUh02qi2/Sq9GHg+6qH/jsiiaxE6jspVU3x5N6unFXjni1tleYvdZ3CjsU4MHm
Z9uRe6Tvk7ZHnBOm47/i7WpclhVXjeVXUcbBEZJvd0egwNLFKmirtEP4lDsqWe3c
8urCMZET8djHIVWqyuPHw7zqmu1gTNxc1BaWUPubocf/wmxWNQA9yTVS+aw8iTKN
cMIirzIFn3iU03V8CMld49ruC99wUYeUd+Mlz5ywLDDBa6pG6J2SphRtGNa9Cb1r
le5uFwHtgqRXGCI5AXf5j5zFEvHwNE4ufjPktL3+/AlYkr6VB4AlVZ6aKCJ4HPgn
er5RdfIll7gOgTxo20XTgRI9Ur0redpUrfRf1DgwXlcPfr/U87KMnGn0G0igmzk5
Jk59JLuRqDGrhIgbqbdf+Gv6mHnZCYx0fj688YqxrUTLzq4RXLhJvOUWLQyypEU2
iQfbv4bcOerFybQm19xg2ALq2I1kFx/p3WEI1KHVp8dwnvGLDQ45dphnisIFyRhh
ok71Rm3T1de8BhvKjD0ufcOV4SmD62XUnsxPB4enT9ZhiGT96LkBK2g6pF1tTFH/
pF85Xr8M8bt5NncNHUelMJSM2O9zIObgpPXPKDnaYj6eYBkOVWNSL0n7Z7nFUvYb
+a4bnEn3VNqv6aNr5bhxNfk1fs9D1sa8I7Kk67znXaRR6+tYXuI1wG7YfrNu5oe+
ifaiZCs8gW1oqTFtim2fxED5SIdy4Q5OcqO+R6aowOJrU9LcvuDqR7kmsiu8SCDb
AKv5HsyC7lbYFBllIZ0izBVeTwrF3SQyuuwS0ZON8zjx0GP7otSV71fdzRFdrvOK
XWX23vQGEEPl58sYlbox4IvlisU6oiBTmazHM7/9g0hxWE7nmR9mdlQZfHBZuO8o
/EcjJIYB2XcfLkmS2IbaarKZziGHR2GIYPtrfQUXYRo+XZRPgdygNKEzRx2QZfM6
yELeF/+DGeLNYXnvJjvzuzPPshPWK/9uwO88T8IDFf3OboBzT7OGeK0kCFziawx1
htsDLdNdqRrm3sggkFKqhpO2Bq1W42OfEZs1poAVwLzr/W5td+I4Ztc+ZbC7Ew39
5LcpNpog6MVVIhMWgQLbDgCZGOV4Uqm0lrGwDsRTJZh7DBEeFVsR+Eozf3E6goOJ
cTrbL0R7S6GsY1UCtCTfnYzF7q25JnY6B14zRlk7d1S/b1cy38kKorWbzjsbELS+
bZLAet9F05x7Q5bVW9vmmzThYq36JcGLLuQxTKyChJ2gwquTxlMKXtU2b1j2NlZd
Gqq9Rzf9CGjPRepfZmqAKpmcCRgL+PYqZi6fwNHkKmrFR2ev0f19wjPPqewN/QYp
Jz5KuJ6xQtCGEUTe9PytsVVkOxmsEnKR+hqEHRKModvT2wKjL3wDY/L0Ks+qXinV
GL+XzvK1r43CJFqKgee+hDqfnlHA2JT4ZeyHtwZqguZeChVhTioFcMPAV2va8aLT
bEVo/D6vebyOuqvS/0X7PpPUPyMgdkWnMlGSWmn5Ud+fi0INVpdVaCz1uTBLhQWl
LRhU1xnHQm1nC7vuD+z9OckVWmV1IbgZUxnqlpoPvRyvPGOFSrbh+kWg+51MvQnT
uZ2PcyQNZ6tZNfz+TQI/wXYHY1/sXZdTt6czPPjNOaSpwWcDOQZfd/vLI+Dd6Z0c
95Ne+B2CAjS3QZ8ah+6HWPRQim1t0HEnzFPLR3GdrNH043+hRmIB8zScc4adCb9l
i3g794bXF4EZhnAtANAyj9iFTfZq9MLyWoGjnX/5Aehf6lcKkvapO9cBY0gOgORY
vYfP/NwJzZ+N+GvF8Cl0C4ogZvOOWMvmD+1FeDHuZFN9n9ix5f/U2VbV4WWsOclK
fIQTegkDCOWOeo8wipSiKxB/ciQjlBwYNPj0MCT8X+uzqg1hTGOOeX/cuBvGbSl4
mBG6aUVGrgwooYSjESqPd0Oje2UUhvNSHxKWaJN5mJvFug63zw+Z0ReMJWjttxvW
+6yxyRj3kKo+g4EvoWaoMP1TfM48zjsjref96zWwmv3cQa5GL74glwUIXWr+FDXQ
5rU5E54YFnQKwgTaI2AdoFQvCXurbLk446LOvZ2Cq/MS5ViCNqnGeftem3g30JOy
AVglybXD8S55i5lItNa5Qi+VyCXiUFPAU3hr4pVnbNqM1HtfWVIu8Ar9GJkJ76GH
DF5QsU25ZqYYMaen+ZYf8WX9tHfmvjyEUI8B6PCdNMDGaZG/4I50CaDuxC3/SEJ/
Xuk8gkDyIyeiwqGVVEcYddMfyRTsFRru4pD5iKjrAVFn2CW336wp6kQJ4smp9PM5
gg5Ped8JxKDf69DX1dHA1mxNuCzIybyKwhsM3Qn7VDNOJkwjKxvQ2PpJEGGe3dHa
w6I9p5j0mFpAk1qO1Ttluf3yUebKfR3L5IJerk12/uPIqGxjGjJjgk408Wl70DqO
DrczRNZlDvgBGr4274AjZP7KL0dhjnTke+egaxUQmnue3Ah1nCVScAaorDt+a/oe
/6gAEqi/IP8X3ho4YwZimCGGi3L3DSXhLS2l4ZiQilaM7UKJ7KnB6XzLoORXysBJ
5q7NgI3sYx4qXBR4NgVs+wUFkfaDfYGUdnB419eDQB4vYwaEbtRtxatZP6N9J9zo
zrwMCnr1P5u0hj/WdRGCQUTPECS/sDrT1J7O1mK+dJ7FBaPthSsLgAeUhAsRc3lI
ZKOUJOY89ztv8ShD2IEU47tWcUoxOxBOIqsDI1W87LgQ/KVL562/40B21au9pren
m751XsnBtgC9xLBl7iun0AQ97eTtTwZOsLJZuQWOmuHO81G3Isd9QdYJcNqAVCIk
kObbrDS+K6RErbR3GopWznknW1feXl8ELK2aDDyoyxC5O0WNQHpc9fRqYNpwCfK7
LvCcWF6PWf4q96vOQY5nFSp16lalPot8snd9jFdMp7fhGz+4QBCE6bajdUnxiHI1
z7Ve7wOL5AxrWH8TfTN7+ttInIEKgimtfNNSUiFzAXKCZts2c7RNDQx1dcvby6Tr
YlMrrM2kzQ3A/8YQsIya8bR/LCEqjkcApxhJRFHXon9pzNkq5UL4nN1R4hn72PuW
jeZy9YTkkxi/9HdJMtlyULA/eN/baZWs2ORDeuzIrYAOt7vteDLFkQaoYvwJ61LO
Iel7KIjEoTp0mUmvr9z+XRR37PvN75WHrY5JNFuX+Cs9DQYqW7WMU0gCNfLuwbaU
7XIP/XeTDLMVINhR9yovEXpGIbV8GouqJcDWWGCiXr+vQ5+KsEIa85/Ox0y6EcN0
pA+LeXUmEAaIv5qxXlu4BYpM4n9KQBDUWlSYF5kjdoNboJwyzAmNeLu0ot4fELOt
lxbcUSNPXXVR6fI0DcfLw632VVCiMwKlA+zzxPbblh+bYMseq4QH8BMFssMU5W5o
Hh2AHqLAI/FPDPzC7zqsNuG5g26mj32i7n3CKs4dHf2yuYCz5mBmKYudBxpPwdkU
b5CR0PKihwZi0ZYmBztV/o7AdVNE0aYMAmQeXK8FB/ytzEi5RCxQWxAnsFnXQhd5
WbzDrPYeboeZMwaVxpzYN3aQjMKr/KL+m4bO3bcG+gQCkYsND+OTdB+/ySFI5ch2
wsB6/F0OaIQvInhKj6av10/1IWxkq2sv6CtlKvaT0BCxFAZsVrLXUlksZP381MMv
odgBqV5Z2lajXfjNgSPUaF4CwMFpLnF81FCV18GaIvx3VWxGs4j0tq89JTyAHLlf
ftI60APua13gGN0Jde0nwPd0/BlsbOSScZcIGQL8HdhtCEMHXa3DABHl7ej3ZmeX
k2wheGN9R4x6YgmPldbiM0UE+aGDX6lZEbN2+zu+u1CYRTSJlkODGpuMuC3BrAIj
5YYVPU/FJgrNe1cCvwFkhVtB72Rl/8KoGlantClfXcX1xzHQpdsEsNQjf6df5HQE
xyOgvrnDfiLQgsqySC3H6n+E9z4GQ9qidZ0Wa7B5RtrntY+vy2kVj7WsiX0kXP5T
JlpIAlx4V6BYCK7P+PjkQdLQb4NFer5LezNCrnBdryLNDigRvIEtgwXFJenDpDZp
jeWCzhU8K8OxKSj+pTTb9e5wBpDYmWeI513CgVWRv5+l0jT5q454YYIsqHsgPOa0
VcRaWldBdXwIaZPhoj0INIzHEq1tc5AQTO3BheOGEFSeUOtW9sEUCsu/1eJrZo3S
pJVWDjKwdh0o3An9m8iB4414Tl1qSdW1Mwu1vwHdKuvJ8AXhqqK6scYfnxc8cG68
0uoL2Y0UPUysopp7EO1wOpE+XRmp4Wp4sEiRbNlbVLtD0GPqXYA3HKWPjn/iHR/l
fQeRih0Q4wXFjLDLb/9Ie8MSqSik5A9fYDxHoPsYeiexf8EUm5M9S/JkG9LJQU01
b3uAfHTedAPKSdZP4lH20cD0wDRN7qULe1e0TbqeLET4aVMjQQUrmB/xM2zFxxfj
P2WIzRos/tr15HLQ8KdZIx5D96YkrlZxlCbWTFRd94TQWOJfM0F/EaxaXmPgrt59
+8hIV2Vs/0RbWGgTD8lUgldEwU1DcdFyIkfXpg/1WJY7icIZuLPL6UbrayNXJGRL
ecjCFuGmO7IrCNDyHFNpqBBR3X0OukokINFHc9ZmM912qF5neuPlcU75jT66yLhF
DmlRrNX7NiS7JOOM2reExIxtGEcIO9Y/NBXnJl94MjZX0FI3DnWfHDDhh97EVJXj
xiJJugAuSH/mV0iEdoYQ+zo9Edi4rsZaNEbgeyp+Boe0S0o30Lh1EJ8FXgZhKuNg
jO6Q6PnJXs8jxU66m0xFl1ZLRljz8GXOjvPXr9Y/BJUTXA9FOOuqy3+TdUPCBDGw
HL/sZCjF3JPyrOL+tCNwTKe+Mjy7j1dJGi/RvoSw9nDKYpvXqKLYcu6MqJIPoIwt
LNKF+OUhp85+ogHH2bT90dARTGJ7VPl6znGWPSx8LFtG4gcSK6/zjYvjm6ZUMBfZ
EiwDl0Py4IjQmYLH4eErtaifX40q8WgcaiIfqZ5DrhIfGQ4Wrt3yxKstXJiQRh+f
mvclF0u/ygxBSnow2kRR4yxnRhWMAI2yW+560T5V+UdKj9qlmHEWGiXf8BuR8jHg
rF7LlptL+kLU4fyXDTaHCu3GH2DsrtygRL16wTjG46iPx6k2kODM3ZwbEqrWj1+n
BYQm4+9lw4BNty0TeP0XO/1DnysDZYhv9cBwhAFN9Egum01SMo2/sXVIuQ+0Og1Y
nNVg2LJT3MBGy5SjK/2hBgAqdSkNFoGZ1imHLy9+4Hs1eWIJoW9oaPVzL6ODxRmG
0emVLp/wm6Bwxi3EFgy/VJMmbc+HobivU91qYZl0CvXcE483V0IHB9k69+fVPu1l
qxDdZGF6KbYQKHrWauwNRzEfvMwLyiWW/opKPCTDltydswb8Fl1Kyvp6l1XAGRpa
ObEuqkfB3ewpX/OkI/oCSnu/JG+vTn4/OZfYSgsH0h8nuwzzgegVV4a7HeY7gnZ6
WtW5mO8iAapBKRzTCONcsEegAYAKRX5AEAyoZLeN6hhPVMBmtN6eWwEVUmvTGt/9
m2VvsWdBE9rfPFtozHdcwbTmHuVPNdlyI7wyUxNWfZ4C9D07rOAqwAn6f2ZnVCed
Yk0Up+KUkrBvvNxbAz6AQ52j7ZsnzEV9npCEoFUR3/tVS3kOKULO7sFhuJghk6CB
VcBbXZX/OtbVXBnZRGK13OFNj6luakcp6SesfouAe1jm76ekvQdFWPgXzroml31F
5w14Wb2rD2hxtayIkwSoNyRS9q3HDLtWAf/5BJKTvgWdO2U0IGgs/pSSQ53c+9cS
tBiDd/NgUfCBHW5uEQqLvLXPi8WSlC1YjNxmWvTIf59hH12nv1AWdCzB899BRDm0
2MWprPnUbbghOPAUGffRW3bTW8gL6sXsszywjcI9T3mp7KDKDWVh0hqr1esUXVtX
0YisBKup/Q7F8DtJCP05E9qh9y56VoWRBR+lkAvvOQB8dq7Px/K0KTUaTA886asn
sgMbY6Rj0z0brGpo7JDRZXLAX9WvQWUP8m8+dVXpat/KyopYTgF89OvEZnrcSewm
k2qo7VngDcAFoM0URnkbEmMMb+P/U/rOSUay/cEp8FCASv4khY0kVDQUUvc/RZpx
eHQ5kwX4iVdIMKQbeNmUsiA7pGBOheTk0Cd0ThTCKWcbYbzzu6aEyJLKgKnwkdOe
jBTTeP7tozVh8ZAPDHy00AL6oG+OYh+uGC/OLMVDvTblhDrPeTNdfAmsnRXVTb3v
x/b71EUXY6XKGLa63puhOvTKVhnnW0tjWqexOA3MXq8B+wEhVoCEIxxzlCPl/aTX
AHQR5PXfhztCbTC3nNIMQoelm0WH9ThPNtFc5dg5UTb0OS13pIN9p+u52UNqst4t
UzWoSEmL3oZXEK6+/2d1kMD16OK7eg4GyVXLmFaMVSYSHCx2W/zT/fxI1My32uaU
U5oYOnVsw1okV6mXquhZSyK3Pxl0oFCOUJ5yLi6bG05N0o4HGXJZo5qrtXrAVIii
0rYKrGvkkBzRiCzJhkryu6CaM4eYqI/2I3G1yaz+V/wZaPVM5zIKnzDLabAfw4PT
ujBieMM3n//qoSbhpzHjRJtt2Qfnd2Wwa8OFr0rH1moo4QgCTrVStpPcwdX3pxgh
MHPaM4JmBx2e76GamwjcGY59DTnY9lHLBkryUtXuU6k93oSzgFTG94x12FrIO5o2
9RFgtE1WiyaDNlk8tP1QQm3aoEiZRje4ER+PQh1owRFHIFGKv0MpwqgW71miJS72
WY5XEot7nRByj4ydgpeR65UAK3IhVUzoeZQMNXlMaIBUkYWhvvn8OZhlH9ivgRaJ
HyNt/uVQojoFfb3dpEvYFA+My7RNAqnHfENPsubYxd+RXG27QrIaVlb5rTRTfn4U
FPm8qScNnb82mwL671WD2v2Z8G1oyeJhL3lT3rEHilv1pjy1M+mzmU1oMGsofFN7
QQkHhKNxeNflaf2MyD9Au55Fkt2vVFLLgSmZdcVVSDgKtOAH2lvUMcDwVB7XEYoa
4SWLAsf9DjfoeC9v074/Wv0nv7YjzeDdc1qVrrC/yNRmXyN56D8Xpjjg835cmPQi
1K90d0TymLtr1QjsIfc5p/LydMoUfxzi/idwAlOUgJ7uMzBvu2u1R8rMncWnPCq4
P/sO/LgGz0ec00EWw46TUMjUltx/B3610PpYHBU2J48rqhCv6EYcA0q0yPstcjOZ
XfiXVExE6eJcvSmtWI2jeTOqZ4TVOn1sZba7qTSaf5mBVQJsXvxLygoAm+R71jTr
FbCqXtaYvhbUewrqX+OuZDCo8cTByIIHXMHuBRNQWU3x2s+9y4mTD6kBSfaLBDNp
qDO7NSCCqCDhsDJ1WLd3yWkRDDM5RM85ZqzUztjYIDfCeiNHkmNtwWhQBPclvNye
hI2IEPpEbIra+xapckvTSJiX9GxeItnNalNY9D0Q4iUlcNQZTs6REeogzSU+swQq
h8vyqLtRrSi8Qb9FwIcJhIpYybfA1bLRkBYGyO2EUbw8m6EFWDFR/MmQZSBDa/JZ
L9U0SBh/bKPp7DoMx7O5YvyXh0yoD8gv0IeN/Aie70MlJQJp8I0/WdiwwNuDEL0X
cZJ42SUtksPQyumHMbYJrTtB8QUHhAKw3kuniM/VXKCwx60WijoyRrbmSArroqKH
A/9yEGxxekdXyL4Y3ewzSoYNbGRa5gAbP7CvUxmTCASMr1QyrHPgmPt7It1qK69C
cSfATJy1qyBxZWR3wlHpaMqwccqpwP+D8fsNYWyHR9WAA/oESM6fr4E1qOI5Ttcf
pZF2gPoO3tW5mozd7P4ukH0NztRS8aPGyj/3+ROvmJqR+ilqIjOqvoPVDeMcTeZI
wW3YoJxGEmEMsnJTXLhCcAoZuoONN9KUaxtu/1DCoWJQeIxaKhv/k/77OZqp6fPs
GixWBPJ9r+Sv7+beTW9xk1HBY3gNz97USHtg90Ixo3xY63SekWrJP9kNkUSRnDDX
DqzGoTuvQquxnZxnEciHUEcEle6i/eKC3PWqzvssszaOeIJKMXDnYVqBfasq1Qwh
Pxn+9YrNja5GVVupbmZNwbA/mppPmm3pu0p3DFfHs5h1pjMmMTT2tk51sbmb8oue
WW/GdtP6b+yT3HJfdqzWce1Q0XzV/7tgfcow4vCkMT8VMXiOIl9rcfJOAKU1IVeE
H93Kes9MFA4e6oOURmwqak1A834uOadoP50/SNJ6v54sC/9KICi5epf/eXJTajwy
l8IBy7rdSk/ax4BdQEGG0VY+AnjhLsRSemaFbgYGo0+q3VHqhIwMGnYl8GLyZWKq
rN+jCwHmMOHxneixh4a1SPgk0RbK3Q2WjFNvYQ6FxxjfquTOt0kLmZRV5iSQ6Lfa
DqxFGXt6eMEm8B2Gj8GPfMA27UekUcbneb/4LSVLEPaiQK+7sPovc0kuiKBCCCqn
kbBXGoYNI+j3uSulfhEocpVzwOR67vMMYCOEkSns7pGdC2sdBrFIeGY3WnNrDR0I
+Z1mC4CwBK6ZMx44x2ET+YIeER2dJWVElPtUtToYalrZi7wgao4Y7iKTGPW+Utqa
fkHx1+rlTEjm2fN2RYV/rT8kSEfJDPGKCiirbdmmR+b3RYiEYfYKC4AzdJdL/tvj
qSNjBEs8Ve5hz8FEw3qVQgeF0FPJ9KKaS/0capZyd9JeYcGiE+rOivWyiwolZ7Ed
R4bs1HhuIHBWHkpJeY4xIIvWGTJlWF0PzAcsRrJyifvnATGY88YWBDy6KO9WOj3W
yWO5g7SeMNbtCIo0hc4NIasi3azZL0YV6o9bVVtFv5f2+k5O4ZLeYED4RifAYS10
P3rvXUTf9yAw7Zu4u8MqZeGyOUETE8FHM9kVgQDiEpZ8VqB56hUAnOhdboOd+l3f
ztMFaqZbEoidz/qOKiS6HlPcVn3YUxdasY3S51evFRZwxcd2X4yneV+9Gj2wK+kM
LyYzeNSNLuroP7dbm4Wt4flQ6cJ6WpnxQcpxhYd/uxHg5FuUlGBQRSgnmHsXfgSK
13byxlhqumbi3qbC7YlIniYe7A9JOSzp97YpPP56w6atpsJdtZkO61kILfy/275E
Vfvq5X8K4Vl/x1gnbUVuhvDqHMDHBYTsP688l7BlZ5F6WXym7B8OTlZf39qXBZlS
7D5tdWJzdmJnl/6/pjw4HawHhULfoML107QjyW0iEOQrTkccsgZdlyQdjCdo1Y1B
vivaPEMxZG83y3Ld+Waj/HFVJwaB/Xwyq3n5NTYvsnyjzPJVvmXZxBdeU1vNfXLM
bGqKYnZDkWm3JKQdycfh/MeFdl6cX9rcYBuYqViDuzdcSppNZEomjRqZUCY7wgnv
Vv1Nv8DTZl1G7LuUVfnMkZK3EarIJFG+GGdOIxuzDd4aAwGg3w8+be4S2OICIPgn
pAoewE0Ocf45mOYFioEM2SIyZKaXmqLBUYPbds+6MxVmEz4EH1hjDa+bSe/PqzP8
7G84E1VQ9zfjW0vdXIYxgX/kp5YE2gd3C+YVMbU//PaJW6cuO6GarnY9jNp6/R12
8EtWix42LmjDKK7orhv6/+PP6uZD7hQwvU4k1foikco3MvU1Ch3th9LRHphVJNbM
kAitbrml8sGZmDQV4Va3HzJLKCPmO2SVq/0cB9jZtb5puQzUvq9CbCp7F9V/qpAk
5SpWEV0tOytur2Y1KCt4uJvNCyAhKP7f06xTzgrt4RcoZFPoRqwDiA4DVm/7LXcN
mQCuHoEsv2WDKyhCrWHPPOYYsvAIrnGvxxoWe/arNjq4USp0drxFAe72MHOdl4+M
wBOYcmNkAw6LEmTc9xJcaDhw9oA8tKMLojf66W7mLfIXE4E6F6EWrEiK99nIPP4P
GvHpV8nNxCx3petwb+4UUi46sn/NXh15ipkJ6gwwWH28FG5233h25iOol/FmfTrj
+VLeCuf8v9LTYzm+tdBEmNot52gjnVsHum6gi+nOcS21RrS39LdxvWcHq+YHpjZm
qVPgJp/Ekal1kIZAhcQyyFtlf5wtgoeLDEeEPFrb9DPYgNU+p1ordQZdxKtSAufk
TIlS6EsIQHJ7vYEw0YKAgb0BXmdTbh1INEkjw7iVwM0451MBpdO8/NMxklugabVu
j3f5d3vaIXXTrSSHtDQ4PTB9ATqqJ2dtXypbJYWfiZHYebM6y7+XUzz/Nj+3Zeg+
NfJTVaCOd1aJsZ+EN3xTuAWQfwUpLrjwcC08sxd+ZfGly1RJJLfJf1uhH+hCNi0j
c8QbY20N9qrP9P/OVdxR4ZmtEzq+p5K0nBJGroKtM7x/vkVYHD0jNb2rBrUNBUrM
RFYrbiyhAR5NqQ7CBKonEzmLeoOUi4yNaDIl+KErjfuR6b2G9uRhM4vuF9TfL7Jk
zl98uHaEuTETCAQTiDIHD9oGldo1T/TebgY8ZEIth3GxlEaXO+lDvf5Ed6Ipp8TD
6I0zgmvg9dYOTp/m5T4GKIY+a90qihkzw9MyhWVlwLhYXK6qw+ojYs5Z1DiJrUJJ
LKitoN+befSTFppjIR4X3M27OK/6vAPbQcOWioWr3o0t/+ff8NXXG0SyGtc3nN7v
4/Pz2yHrV1+VYeYvx0eF2yPglwrOYopWlZ9vZ5BM2whsWMnvdIT8EF/auKb8OzFS
hNrF/Hh1jNocB5X8H9LnGFPOFjM6cRvUMn9OIocXCM950lIv4dGoKXT4g7ss2vFK
62padm5u8OHcE8bPkMW2eMeOk34N1Y650JcyE6IXEgRyU5rMwodjSGuOdWojKRao
cQb9ZgyIGeaNiLphD4Q80P0ekrtQ9mNl79VzcQYnneFB/PS8qcnx41EcaQDEkpEL
/s2K6Y154xgnX4KK0mD6Vdi7W57Xk4gOG6ERFQRdAoCRLrdAs3BPd9GmV+OlafxQ
4jB+wKwxy3sfHV2xN1tUMq/t+Fifc1V3DbzgCPM3t28Fok0NuZfHMTExlVN3WQUH
BTU22L4QolDQF0nLpV8zh+2Kl1f2tf0edaJtyR+vUfoLMJZkt65bDzz5Ly7FbSlj
EcaIiZzpXGuQ909erCctXQ+pL/TEZw3ruxjQZKpueMjXgRye1DlutL1TiFOidPJT
aL9GfVE87sAmy86WKgubn8qdtDnxdKJxGsWas4tABD5637vbUBg0p9yVvwjx2Bnq
jtS8Hs9/qM6B3SZQGgZDcQi3H4KFFAjCd/7LEUYYCXjzD410HjV0yS42Jl724Uac
EfxfpAIurL4uKDv3r23a/ndxQg9rBv7SeDCnoz71zkXRmCSwNkEe1EZe0+AXs7OP
OuuuiatzFDy8uGVUlAFPh7/0pC8GNXF9LVq1f5dMEiZgb4YkBT2jyBEPHQDapM9u
OzXL1vrX5YY0UrgGrID/+RLnImtxzsgZyr9fWa5+/4G9fqsJBfzkJnMz46xBNEK1
qflmVWBCU8d1O9mgaAgXMpemtDsamYUev/G1eo2zt/T6Pdr4YXD+yk+O/e3VaeQ+
7ntushNHYEAaIlJUpM5+QMHnZyvguXjZNGWV+3OT0WSTmzESVAGUNQO+NCUAz9Aq
Y6uofU3h+nEZpMZKwvfX1PxMS2JW2o81BboYlKIEyIuY8yfyKNJUSuTIInnmB3ZY
lc3uuY9olaT4JQjnpbCO9UAHR1yrxcIyakYmeWA/8s4KIvpiEham5hIrfvGpbMb5
84mA2iR2ScL2hzKHfLdgNppLd+uM9Tq6DLb/r1RxmLcyiQJwX5yvzK3zG3lFGHud
/W3lU7S9UDngNO/920WL54RJOB3ZUiHIhPvKWUUAjijv2ieR445Y2fcsDvJ5bm62
zFCrk2BRDFQcGX19fG8f+5cCv01sBsgRFt9vH6l4qZdpy1njjFSEXLZ+ro9JV3Dx
FOA+rxc9GE6bwiY0E5GYt6bSPxzlxxVsCkCMk2XRlR1cRdMFWOEFtGd2DU5/T4xX
VfC6xPLZhzPyIPUW6cm0teddbmylDmZO79KA+FqI8L3u6TAqlbX/+xOa8WPrBrdw
YPRLc0QZzlpN6rTbLfwHXoBJfZpH64UL52Wp7IT6sC685aT2syY8ePjc0pQv7zef
VqVfac/vp4nWJ25Alj9v1/YCSm+v9woLhds2vy7E4ef6HIfglilCNGQktdHVCi5+
W6x/dDxphowAMafAtpcMZAA8J1EARpJk6vgqu/7OgC+412SNCDc3baHrUTxmVWGg
Enn/DCFdJ8Lw+V9dKuHX8KuiYBEzAG75TTpq9ztJMAIppUzYIMESqrex77XtEVAT
SCwhQOj860eLyjvBj2ru0nOI4UBxpvCvFecvGmoysKxsn47u2iW5V4KFZCrwjS7m
o1BeHuIwMlmI+Dlg4qkJSKfledE71Ui+WGcyPN/GV4sVTM2d6XJbJy0kzT0wokZw
VhyIhwdMuXRIj0qS+rsBZbWwpDRbtMbhdTKUw4vLCSJbwh8/U7W+haLllsRkRsB7
X6VPi9WXaFVndBwNEE2m16o0iber+9KtEPmxSdm/Kzdkn4f0NG1oQvt5YZROwJ3k
AaBH9/SMreoWFy2hmrMe+6/Wwzg+WiWhixHICeIHFKjKNcejU8Rxo9yuhPVB4Aeh
5zffAoc4fn2qCrpT84EYSKdGSpz+p5Ve3cWZUYOZrSK5aPFXbNFupI8badDbrKLK
/NSJuzLEGrIzk3ZqNsIelniOpl9+Rk3AnolA0DVhUuVb8z7xFyn/4F/F8TP6Yufp
HF+t/LTxuotfq1wmvw4RGfx6E8f2CNslJUTiAwgQ/JTMAi31GyrEFRjspz2VVNvN
KmU9pVQFwiTlCZ7YJvFxcCXhPmQ+OSiGcT32qRUndrH4vs7DCp59n2hF4basYUGm
o/oZNaCBGaE6IQYCLXK479/mWnseIZEsVFuOiTLNEGw3WLTK6hwiVxcWxA5sAvy1
+UFh0COPCiFT+5uXHcUTIZf7tnIOOzd91Dc4mi1jmX9mfZZFZJKAkpmAAjEkxwL8
CmOYLMhHgPkIvqGCtHELg5mkxVcI9YGhOYUn10i1ZXK0c2esZxAdk4WqUT1d2TKr
5t2ItxWGHBP7TmxJzinqEliGVSnSEqWzugXbbRD0pElU9AtR1S+BUaVh0xoFAH2s
+10vzA4ZN+S3hOFDtY9hy5Wv2hMjrV9lDxAJ2H84KKTL8TiwfGgURjs6lENw7Lx7
aqdkfwogJIWhS67n45eKMVT9V9Z3JPndRAOCTGj+kxSS3/Cp/pGx5+q/I3LbO8j/
Ys6o2jExPfLzvN2its+JNykkjdtEADqnqwKbCMRsSkwwvZSOuByAYBxbj+YHNwDN
lYVXLzDADEURBzCTe6eqoG4wVNB2RUuWAUqxkDSDzU4kwOXfTGylHXnMO/Z6gyCf
Y7u6qeKLF72BYHwlHEWGZF4gv1kZRFX4dHVPUxpcas14Umh8+IszvYgTA+lA7PSw
IlO62l7UdingBt+oJHgW7lt3871srNsZNNLljiq8/6HvmENocBMQwas3hdMdVdHS
E9DM5xNQ3tLVVPn8wd6jHh0T8eRb9J8xAqWn4lRc4xnwWssW/q5aytZMqwGNNQnd
H0js1SLKWFsTopUOyiIKEyGpPyCbd30o8W4w01Kvh59mznvoGvteBXvEjqT0uKwT
XFfQO/Z/9ir1GcgVHYw9lqI9FOWLn0aV8zUXq2mzK+jHouX1VHK16RceX38J5Iba
szHUZZ0D1kmuj9JfcACSMb4Q9D+TP9knbkUAh+FlWaZbmbuAvBaSQbcEHhPvKyFE
6V3vclbO7hgAN4/IqCpLV3yC86P9CjPDnGyCrG/MNZjH2DK0vkFPovaFwCFH3bjW
6Yax+NygMydl9gPxOyjsj9Bq7Uc5jScC67DfteFHr2qxxqD4TE/rI/YQGV1u7zzh
WaQvJEDCtx22Hu0nxOfwoH/3X85w+EON82oOdI37kLqVG8v/RO77Dnb17AR8OsFf
FwnHZh8SMKejjfXtJYPfMqQk44bk0XFks7x/y6ggXL6duzNpKTq0n1lQQ73Plhe1
SSryELssYIWy/7xLItvlZ7Jfp4zwOn21eahEpwsUHcPbvNlStQnFSjlvw9C1HZP9
zF2+ScEHAoS1YAizivvmLaKKK6PT11vYUI55Ziuu52lnD27x4Ss5A1z7W9+wUU8s
d67r0a8os0w+mperIGngCOa2MvvVlKdlbpieC25hDrrZIc8BKplGq14Z5oZXUKhB
I/3jihfTT4F6RRqp+t1IqDXsUH8u1bR5PkfzCl4X/N/edvzK/DKbu4Xf8IV1vsz9
3Fky2zGREpDQL042Ym2cMrf7jk5jH/xEtINR9Gme3oyQAw0r51Ec2B6z9vZ1+mFS
uDVLkrMyNMnBFyX7bPWP/F4r2RxNVa5o8v/kVc94EqzJOLei6maxvRGo4atlSwbl
3AMJaN3712bpUQodNUsNSzWxcaQqehKgrdW0As97k0g03spUSiIu1i4mE/pLYGxl
NvgqUrFTd8u/33mdj5gNACLB06qLf9ws5ib/tr20Fmv4SB/m8mD4lWoAcjg+KNJJ
Rutxm9ofRe/3ASAp99gfn305WUSGmYMs3e9UzuIi/N/7xJqLQi1f4dfdTZsGm6Ig
h+peJ/FrdYxpaEmj87KjmbOFdosHiiMKCZI6YG49iemUDo8wjuC+gTLlE1gzxC7N
hUBElkg0J9tFDGCdeyMvjWcZG4tYCBO8R4gXkeCRhuDmEMcV9ncnzJceq/Di26g9
X43jHtQIVVQu7oUc+d4+/o30zc3FJerZkaoAaB31GyEKxLRNZmzCNvYw45A5qtli
hDwdGmacFP6UEW5/xUaVoSaF03NQqDA5N+1Ef/Wv2vihnsnrJvbe6RYvOIY50cF5
FLC+cUQgTDzjG3jtiE76Nb1SvqSYo2V1OaPBTBhn8C9kU3O4N6Z3rVrLwhJyIrCB
aVqz3Vlh95glnx1sgo1ltf04KH83u9LMte6K6t5AyGJ4D7nnF9XBUteX1k9LyJ+V
06k3hjQ7yQRNdsUiihtmYyHdvdp4t/kEDkSoRED709pjc6cBocLxwk6y+1A8iYkT
5VAcPvSeBgW5HRCZ7xdTff6XoQBBsdM/0g7BE94naaGjoAuhZquDjdLCDgihw3qr
WI5nIAxNw1I9mJwQ3WvfKvHKzsIWSiNnMoocDD9ImGg5GW2kHeK9e42vtzsHKyNa
8ZfDQiG1WzlnUpuNoOUOWWoNmTITpPo/TfA3sDw3Ay5LbOygwYdKZ38VOY2r75tm
b6lfEdDXROLG+5Swle8yPpWxxXO9wvQIAZLDHQSyFSm22B9cl6tBTWXfBZzYSf5U
0gODMqjwsbQP/czZGFU4tu3SLvdIm1E+CjB7a1Wto2Oe1gI4o2g5cnyzrhMo7nO2
RxZATx95xFIz5ODvvC4/vUL8hWPAblRo0txrQzNKKMUDA9LzapNpImhPQg5VnCzs
TFm1JaxAhlT9F1bvWvrsD3qxxUuQ5snSkz97k2WpSYI4iLJY23RupyEyVnCih9x6
LJDKCWw7vzouinGqM+uOEuwURxYEHrKa8p/17p0V7O5ZXpxaf5lGjdQiEXsPlmcv
gmkBqWg6rUpUH4i8A3HUeFMCOgRNmzMXaFqP4HBTutxexnvz9/Bw2bWIVdsRpVMJ
zxFIcAUzFot/rZDfDRjPQ1NLetNcNb7cVuK1cwFby8xGRdPcF6e/12DCB5K5hH4i
Axy9aPKKtmtgJkXGeBUfpDvVEQ4YFI0wbt/s1rZaGzGwEFZmm7GEo4X7qYWsjLca
XKvFucrUkklA6+rfErDYUg==
`protect END_PROTECTED
