`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6pKmzPaMZdBFdDXFe5phZI2bMW5vmWRES1glh75LzXfXk673DWUoW7ejLOgc7nzM
5bRzAVJYbArMCHVQeTkGRMBZgW0hs4Vk/WnSuxXS1AcNeVji2S8YbM3JjyKVWOzu
0zOOoFmF+Vxu0i2V9SmE+WNSATP/+prcmN+5xQRo/kenEIV/3GABrq0ifz4V24Dk
zq64Of31/Ur53eqeD5ef19JcbjpifgT8veoHhtXNOdFhqa9ET63Mvin6jNDmBuNm
QgrC29HHgpQTdcQwMWzQZdWNQRuWZHXH9X/wX+HatZj6ZzSgwoh2a0TCX6J+1jQb
Fik2j9Xh5DeC+16jEV+y6POpBUy7kl1OqXpjMu8xg3yRu4BCniPBzeUCIYZW7ncL
Dx6Qy9nBGFRiuZI9BMjbr94L9EuiY18DiBkB0i7ysPccCzJglP8ZyeI/BkDtJhtY
`protect END_PROTECTED
