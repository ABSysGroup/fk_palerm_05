`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CWLywKJgQtefcJYIInzMB0GqEb8w5/oxwlgPrTPQeXdNzaYl9bE0Eg+cg+6MXGU9
siNYLXJ4aN5yWD30NU9Uwf+fqoNBOdqNCOU3JlCIicK4l286LTScCqFqo1CEEfF0
b2Ib180KN81eBemZm4YbJFhh86H4Xg87iuIlZS+a4YqWz5IfArBmUJ/ZyMs76fLD
YR4ZjRn65msKRXClmA8r5/ohJ+g9Ae5lIlGZiR1n8lq+hdtXZ8XPdanxh2rEnpm4
WtUNCTbils5ymj1C+Z8Dbw==
`protect END_PROTECTED
