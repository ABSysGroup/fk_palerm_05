`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bEPVw/lp5Jn8nXZIR35ND5nZddMSPlDzNUjeDLURQarU3T1a/fPXpjs9sDh4//Yu
AAKF+Fj5vtB5v6D6RvqVlYdNDg8iRqu6XswKj8++e+2qMTw7JRMKWOjiJxC3EgOH
l/NOLX9Sp514TEl4Mp1UldqNFzYvsdAeBFvYcUs8rpMyLphKW+qeA80cyIOd+sDh
blUyTMK7lIAcdNtPCFevXlvyyo5QtTTbaju89Fo74QsvwIiuJZQ1zWIdO8soNla9
U7EBo308KMbAeu1FD2iJz9mBiDbUuECaG1iChmzTGtfX4xA9Hsf2Q9IO8rlv0AUD
Z9Fze4srhGw2HT3Pw8pPq1prFqbTb9VMcbIBe8JpyzrnWW1ckPNZ25qvlxRDn2Ct
`protect END_PROTECTED
