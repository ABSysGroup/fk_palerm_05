`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4yiZFdrDps1d3Y16Ve0s+Bue2LQLfi0E4L8GkoCFghjtPX5QMM+lct5TJ0XuTTbz
l6G3X9/YpVGGY8omatYgvWjxkl4sset7Kz7DskmK1uxMDO/GPdOY+1Xw7JRClokV
43Hy3ysNIA2yMBPnHXF0sTD27VcOszZcsKjzTjII5TkQ941rQ3PAubyUrlfYWGDc
qA44lOUk4palCCcl5Mf3/YAX/Un4oKoxdVsLn5QoQHpQzp5DSa566Uv0N8Yx+t+R
8qSrWl0MzfJwkbOpfLq5ts5aOcloKGdTp5BlLmH6p6IHMSdv3Nxytr0vLoFsz0zN
3X20ltquxGaCxQOR2jMHKqiZo52gbxKjpy/rR02+g6uaJuQ0MZhRerwq2QRLJPbb
`protect END_PROTECTED
