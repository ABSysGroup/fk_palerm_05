`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZoLBKa9RMbR5ml/FEEcE3ubYF80ZWwceHptCyrg0VSIlJYPctB4SpBV3SCkfmIga
Df/8DcD0Ewi2a/ywiNn5ENMZAnq2IF5wwQq8g+dcXVSGixAC324zsAaoDGoIUwbw
YfSgBcB5Q2YHdW3DsNz0+TD62rCn4QkIEvbvw8OzBXcVjCgTgZhfFJTfBMe6SAXd
h4cwJGVOQPgRzBKmVK5ecspGKJHwNpd52cr0JyLqNQqyVjH3QbrVM/XIjGL93tIx
047CL4JV4yd1hidjygfmxOMShydbFxda/YXs8v5J/bm/gCqg22EaHS0QZ4PbPwP6
dtkjuw92b6wdb59jPmgjnkrKDtWOV+tn/2ZOdKDLzEv3LAe3y/K7Dyndv2/abw4L
aWc8HCvBTDzjuzEPV48Em9mPMgdoIIHSA8mhd8OaiFz+1Jon3lo+vTSC1ZctfNqa
DCGNEib27om94aILujBp/e3sB/CJtPyBtkHYPyljOJB8kye/iFdFDdd/aosVoV5h
bEJW6ZWZ2W1/vJ6K+uetyCDiKZFX1JWQEe7W/1OTEfsXhxxnOzzZiF4TAN1VV8jA
uY2i0TyNKGx13+Irb0I9gnxriwlo084lyPhuI1OdKbyFRHnsjH4NaQ2nUpSM6YZn
DFGi5vaZIoaVuxGFR3jy2a/3IAbmZFMhef9W/PVZbWOy8S91dbEuVqQbrxwRx367
ZhFXEpK+jWy5cm5wvb6/24WhKN9+0oowFdVn8KCuoAzW1WzZtTTN1T4b9hfovROT
2rOmuI7yednV9kQ2/+MmORMqiCMCz9WrKCpOeVGymukaWJ87KhhdFRLUnRSCsIJy
hAyoR9cvcSi/cRqW7roaf7aZb3onNbIDQl8z9LJjS5cPWg2JkB9ZbmhN/MV/77c5
UkK4v4tSagZ7uxnQcsZfY/jv/gaA4S+kI373GFjUtPK3cVTS+MNL1mDSdeFh49ur
GA24KClv1GAZ0qzhaWb3kYYcRGS75YiMGY2yBnJkPMUyU0GtgPp+NxJJ12xaFl02
0CB0P8WNTMPSUOXFYi3EzL234f6a46ObNaO5ul+Hw4TADIbIab5peWi+uarVVNne
aCum9z/pUt1nO5H+Kem1BHFncFxshIE27SCDp5GKKkiEbSTBJuX/YX92hAEXHrGn
walpPAfV81A6xBpIveLbZ5Vnur4tkIWCipcuyFfqSLNpuDxQMsxOHAAgxp36n1Lb
QjyHx/FEr5lrzKxQjjLEHuy2xhqUvO42uJ1NPrxH0usFc+MkcXF8j0cQcoTS6pSa
KrZ0prS4mNK0t2aH3/HWK6AGns50dvz3Bgfq8AozwU9JEMEiraygO8rgSESY/sCF
hont5nIvtXSNnp0iuc6tEMxEdkZcoMXlbPszAfc399IL8vcj12i9z2Ez9jalMnub
tUZdRsyVWdf5UP+s69IYILR7zSlmc+YvtQEOzQ6CYTNMhO5sEXSnEZhSX8l77dAG
4ll1Qfva902XwPClTws7wUSVDNBdiEMiIT0m2V7wKLcCtQos+vFtL1PrPNn4cEq3
lQ7KNsl4TMmU9qcQKARI5ejWLqsULRG5VMUWeoxqMSXzPAvIN72cnBxhZdfnNt+t
3jr8LbJclp3Tk3eauvkbyUP6zi8V1i1KPypNFfrQrJjdTihGoP6ZU67QM/HUU+7K
sYkpeprFBltvZr3b61mW/w==
`protect END_PROTECTED
