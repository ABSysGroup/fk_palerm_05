`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u3BRy3Xou/FCTArwPI58+t6vspUBOO4A8uobMfOGsmrmHSCnnMxVXs5mZXOaOKc0
6lGTUH8fXbrpuknxgyYldzWlnPx4hbz1zM4K3N3DgFZz4QDFm3UB24b2kci02Yie
skp2c1P0AT3jA3f1Ki7zO39Xz/7u4Za7By1Z2bJKLq35rVZ0atkBM5DLnW4qBB4B
SorcCQh303zYqgJMzGw58nrLRCxbPndSyeBnjo0p2s9xfgMZPeiEhCgrIxhIuNuL
iZz1IZg2f1iSdp6YlbQJ7UBesnPK8/YqwjsxtDLQmUKu0c2Jm45Na5H95YKMpDnS
uKiKMrSHS6PPfBns0YjS8w==
`protect END_PROTECTED
