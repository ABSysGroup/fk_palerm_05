`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WJqGpNji2R+WH7t/ZtT8gG3k5TYclMNU2eUO2hCqvSnT8JwHvYDdjoJIo2lB/qoo
TwXWpU2+AEokz//ciMeyTRwo716DY3fEqCsJNrl+4U5tqWo5g/eYbqTAT3DhzjF5
QezKjj9OPnzgO/9pQWU2W/nKYbzASGUYkQdh/l8MPGYXo/tgvp9fahgkj4VCKiby
l4COm1Pes1PJMLMygaImh9nH632FuQ8PAH0Ox1QnL/HI9wp9foL1+j4sQ6986Udo
I72EP9XbgOcLfFdNU8PmzSZpOBH/xHk1ickP+/j2xQJ5I8kmQyMV5Y6toa8o6Hcb
9YAi//7FQOFEZ8uMb0n9ZE3KyhWOZLpv5hiYyovpcc1OrZg+y3eXYn/BF9ihcRl8
d5sUNwwtO2Aypw4U3Zu9Mg==
`protect END_PROTECTED
