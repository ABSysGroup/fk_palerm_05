`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oUP3HHg1bLwT0vJDgVunPvZD1yPT+x8kr40a7Ot5W0uZU/2l7knty/HVV3yxWzS0
/SuAXwb5BYjOu0k7tenxn1Da0hCYcfC4KtZzpogCVF3PuhdLPhjaUaT3Q8c3nj7Y
Wjz2MBps9BChLAvf7O1K0t6K0Ypxj4K2ooqRU7io4MHtBg+AbstmgyxG/oLq1gYM
dMwVBODedO8lK5R5qi3JNh+3bBAR3ObQrpG7o+QN9gtUMjv/+xvyu1KL4WzOvQ45
vqGftrsOM3JCbYH8rpugacCTQdjeILGR5z5KsYnCaVMwoFnbpvJ0+20o3AItwYRA
fB3E2cXpfIkUavkHuUIGJlfNHJlDAHLnGAReumFMGH3Wf8mTJ9Gu8zSWZRec5cWL
IfvLSUNCuCi1f7UrSu9zhOjOBwRhpQGVxzQ92R1AbdeaZgKfekNx/Fo8Qf2JW0pG
vzzV/2an+Fk7FhsZ6tP8CDyPolIzN7A7HBVLNJFLMLA=
`protect END_PROTECTED
