`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
thc6mq6qVrJc6UsJkvFhWv3XkFi8MPNKHsyY9IZqOINjA04RH42i4eK0+l1tBbr2
4jwKopdtXb7zRtWb0RahpOWhz+tEgWV5zxdc6uKTGQPexwXW1wGIu/XUU7+5BqCn
N1h4ycjDvc/iVPTb3LMCexOBIv/bnzjYGOImTC6OIVI+UOac8oq89vABLZYcZEru
E4FBZWSShx3L+niJAr0T0pmoI80sn/OARjzz8OhAx4mrWUTnYO08fblwdej9qtoT
mMcsYOiRZotV5qoz/I52bXdTOHJ7GW0Qqj+MGczV/QHjvZs9bU8eAw3BLGHF6n4x
I1TLGCzcgRdcAbXXVPHEUcCWo5SFpu1SPGEsmluNxGXSP8giiKLLx1azDhJXp+MB
viLc/ltG3JJZebxfDVG235g1HeKfyS3GTKuwQuNnTeYerHjHvmFZNL1tpdGCzUzG
ET2DyBYc0SpZq/eHMFGANb6kEKAVwwM3GmB0zVaYr9u+k9YbxT6Zi/rThLAN83Q0
tGwVjwkMPf1awQGClstv61e1Kbd5bisaqmi/OJUtAoAtvu0KA3W+7XsrQvnaWJZ2
4JMJUdn+DZuEpYzUlGmQr0YVjNxY8EmJqYjoemONrbhaLTjxrcni0gW5OJwKIWNO
QdZPMYY96GTRD4jgRMOVLVdHnlOBpam6LEFwQ08wc7M=
`protect END_PROTECTED
