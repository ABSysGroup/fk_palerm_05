`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WpR7o9GoIjVarlVVNDag2QIoJv+/RCvCUH2ZweOMQtpAnQJZwrG4ynFrQsexq0YZ
m5vWpuo166ZxprPQn5HV3DqVi3TWpCh+zWoa703AytdbrE43Ai1/lJszwYl04HPp
yNww165ugBuxl+NlZgFs+pJjVTYD8cAw0jcEkOCndMlQy2/eDolO9sbYbIL+DgIo
R/Hdcp/yAl6f11T8AuYhaPMokG18YOr3bkyk8lmYm62NkvHaCg3Nw3hxW9XOlie6
npKdYyp+bAFa+FsWQJ+1Pa0szszv4QJ/FqEUvKl9GdilTaJCEQAH70crbrCWxls/
znH27e3QmuhGRHsaj3Di9vsRPdZDM/X0scDS0uoAYo8RTQaLLza5Q9v4kR/eoJIL
r4941U2tHpez5KpNnUO0oQ==
`protect END_PROTECTED
