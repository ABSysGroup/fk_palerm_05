`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YS/5H1D9uy7TGhiiy6vAUF+7BPZqAi3/QC+h2GS2XwvxP4qHldhdVoV9TU2Yy4W7
6QvNsvlGTM7nX2zDX9jRME/ceJYtc0UY8sqZC8IozDuGmRPebEfKPUgVrr/BU1L0
QVYLINJgq5AoPzK7BPtybUlO3IDU3bg/y3jxzueX0RaQGBO1zlYPpx/FcmgHNX0/
kiGIoYRd9NsgML3+BksOC7PhtM7v/2kKOkCD9qw/1dwV3+lj+GBLzUBay6fDBFad
YoiDjpPFW1sNmg8Qcbm+R5I+fj4/Zd07NWyR/3AETMZTaQ3PVlbh9aypfMpTCd2a
00rQnNKdOZR0+5xMfynwbrMAkCI4mqCJjgwP1IZ+x4HesSwEl4wgBhX66Y2wl8Rz
`protect END_PROTECTED
