`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KuL/vZ8yA2XfjndljGt8fy1fbUCBH/FNKQ0WQiDpOo07JxTxqH70jVVMKnwC3kkX
m1TqjPn3rw8vzCtjjvRMVMNNFUg4VURKUUf0v4Wzyi5aww2poGIvqUYIld1lR9ls
AuX3sFsN5NHRzgP2agxjP9sk5+oFrDPvxzISUAGIQThCknqTzpZf9U8ypwMtXALs
ToXv0mx503nyDopxT927E8tGO9asJB7mgzgwwCtGU5cwsDwsze2wqc3PNOTd+5Mx
Y4ACVpKD/QStMnUL31lWB9szG+6YQHASm7tXvU7StUBB7trekRWXYV/SUlHQvD9m
BipbalmbbgKtyxLNNj8LTeiW79E5cUg6leCl5kE/ThEV1PM6bRGuT/z4qVmOeNsD
58RmUy3X8R9gZRKXRN8CKAgVtWZU3ETu14AD70jF22ALl/WxrzxXDZ/KAAFXRo1U
3fPjA/8/qqCjtGZpK970LryTeX2knItCQo+ebCfEQZLrEUoNvlnCp40QYvaFBj88
tYhixmeLSG263q6JzvU+0w==
`protect END_PROTECTED
