`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
swdhG3vHFskR6V0Y5pB9Fk25/yQWgfdp8A5YXVT1g2bqt6XLZkeVpWV2sfoFw3xw
HrfazQLUs5baESgb/TCzy9PYbfZC91lbrr/IodT2A6fqpRGVq8lgCBS/FQzYuUdJ
FabMogGyQaHpDRQdM0piLZBL+rTxqS2esT0TgqsIkc5FvWyQwwgcgZNU5RuUPlI2
uykcFykwimGOGWmOdXOQnL5KEZZq1VTs734Q/72sXj5Lb7PuXo6gUlwMqqB/qGWx
OLWpmpyboYM2R7quZEW0b+cbAdSe3WyeA2oCL33/axWV79F+ucKBq98FoWKt9V+J
hPd4JN74dK2tGaQO0PvzWv6KupX2z9HInsBTM70opZGz/R0HVtnUZCYbrXxteFkY
WZWjKIjukw12ZuRqFu2ImBDiHai0qGNXVLiu226XM2o3zAfY6m7nInQ1nArVLSpZ
YLeS/7JxoCFHPofM8xoOCvgglTPDfNuKcNdTb+tHzTABgIfoaRvkKsC7zbddYGxr
ESnfpijArJXUBWwCCtnb/QsLf+oesDxdwnlUprtgFlUeupNk3ImRHETkB0TglHum
ckWjXEXrcjs+tUNToBd6Rdex3HWF5tPMw9M/6lUDam3iDNK8zOjagoPU/J3BQNvK
WcT6lOONrSw2mkO9BcdcMg==
`protect END_PROTECTED
