`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O1T5zvn4HxHdl3lDXOvtjp7qDrDhtk35qZmZRSHaSYSjksl2xCfrJoYKYRjPHdnU
r1QdmV3UED0v0OgHXAJPfgQ1eq3j/v4aa40B2zIKmEL0eERK9xvwkUFWiY3UctPv
gRC9mbZneh/K3wT9aDWcNi3osWGDVB1afcoOiTtI26fNqXbflddTZBHlvC0M0R5h
ASqy428r1yh2cJx6261NllDTtEbCfmnI1J6CsxeRQrwst8jtvJ78jbn6hRT7vhux
Yw5xjux9HnCFsN/XAMXSwbA2ce3g0AukC8JXwn9jLUBpq6MfiWJgtFqC87rAVfkG
UayJ2b1Pe/e3u1U3QtYEYWikDmnbM2tZUAkxGxBwOsCFqh9XgWWvZFZvEMlhw18F
vRgskT1hvtE8shqXOWOfFO2Eu7WBEa1k6yY5sWEsQvfiX3PIg0n2nm0xGDhn+08V
jiakTjfwu5J4gRT6NOJBW0bAOrMfwL/+xMr1e1rEzyTrk82pJS88PURNdOjPbGf6
BMoLFlSFonHeCx1otjnUTWd3iXQBjnerK3Nu3um41YvJC3LtSilzsjcC6K+JraM1
Fwh+9EoX8H3ZaIgktUdsPY5269R3FYox4sUGv87Px6xZCDlf6HDiRHAeFVP0XndI
Xc+d21euJojLC1vKQZXz4YUO0bc3H1H7eQHetNvzxH8npmpyDE6TZ0qX4gl9xqBQ
D4w7YGhOK71gzJ7FbteMOJlfjW0fceWfjlteN6mdgsgdQoe3i6Tn2i50iUFO5X+S
fjVTjUmnWoo+6kS5yyY63m8ZAo9N+ktVMCFFXT+z8pw+8HaGmBh0TxLBUrnQGDNn
jozHIset8csfUHi3VenhVgfuAP3GYaFI1OK2JFSAou9uRSG6tZWNJkHfCaQ1js8f
vUAtMKxCVRebP+yL6W+lM4uSaz9SS3xaydkuaIaIXY8trRFEoY6Do4liFDfHQhSQ
xZEkUY4qdB9dovsix8odszJFmJowQexR0h4seE/Ycw5rhrGPnyzeOCrqY0DFMt5X
KCmJQajLWzh36kuik8AqLtTOwUDtjkEt8U/K34u4i8oJJFuLG1LDL25vq0eby5+k
SwBsi2BszTI4Xl8GU1ZFCZr43fp1nPQWD3MmwxuVqAyBR03qgy0xG6RSbkMQQo2X
YCHvZ4wEK3z+Dw0vEi5C71uX4miPABecQnXAz6n3bXTkBPEvtuWwtugxce6CGCAa
7QUkJyLG5UNmjCVxst5nU9PZDIVnyTJnJqZsvnCfCv5T1e8KCmcpDtUX8YGGDm49
NBHVal+nbBCYLt1Rrpx7tZN5TM5m6zuJ7VbJY+4/vMUiGTmF9Leh9sndhxih/pFs
CGUVN+bV0VzqRHxmxLd78tMU729ZP4BjygOu8EUUOATcwtH4+bRqlw3kgOAi9FbU
WnsXRO3KkB+nYuY1MJW5L862vec0/HzVghJKvMlxrGwXHiBdvXFPpH5jWMBmCxkt
j3Z8EP8GtRSJKsmLWPTJ4Zhj8CLCPlEa0GB5bnNUpOJ0cDuLdyVU0+Loum7U3pjI
SXzb0exmF655mbKftxbAucD1lRKWt96lwxMBFOPKcf1pHc7flNmYoQyPgwIP2VFH
v0nUfCeFBNrIrdjr29sIjutwJ6hqk75bnWfHYCzTOJ5hNfXqkl7/lrUrA8bKJ8UI
HrjFXQk/VgSlgzhsAKl1k/BP7P8CxIJ33FBgwyZoF1qLEVZliBFRPtnxGYGigWZQ
JRd11qTDYGlRsoDnD1vVi1DtPKQWHeTJ58LwyuLcgsoLabvrW/U3J2pHLQAjtfdW
xytPAeZWZREJfhuvxvH/6Bcs1scIFM386TBlto+dQ/YTyAAwhQGA+EA1q5M87+/q
U4iPAZNBqW0fOnmlMYan+iKzC0a0uBiliMoLYjADSSMhSWSIQn4CSKB00xHVvlCT
A1LvjaVXynnU8LXYip/0kN2aV/JNpCvzMtu2lxIUTnP44gpK7t16Jkoq98UD95Yc
ayYaVTPSRPunLWjzTkf7l6MADJpyDgX7s6IAPOAcrgAV7QZO7A1jwKtWjalWB/iV
HmHId4IOFKQAW5bIxslHHOALZy6W6Vu2P6k/Bm1JrUgxtZ54CymAfV6ljoxaD4NH
1bMKf+FiFODpiz+mg2hVk0a2SBCM84UtdBszQZTNY8sG97GZ5kXITirgrMEMP/fx
VQwaAlKBL2G62G9cZbXkItdTILwORrE57UMqAllg/aMsqiYY0aevjsCt+uDi42qM
SlgIMXPAn0iqMVtxud+v5OGjgcGOHFZC5G2dLvUs1izj1QD7t74pcG71Pi622jAq
Zz4PhcA/UNs47GHe4GTzoUbk8Wz6beDNoL57qQ95wX+SHxZkozdomEkmIKRqwbsT
+KqKdguGmlOH8ASJ36dlrA==
`protect END_PROTECTED
