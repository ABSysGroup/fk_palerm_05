`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SwqzaPM2VYyB9s4GNklvJYgjsgd8D2Tj1gVNQZqDe4kN3O0QE5aPOfAGsJQ4YnCK
5s3xAtBSpYCblTCnh++zMsQ6nkX98DQ8OXvx8WPvASSnIfLVJ4rrwHXy4ShaNZW+
KcD8GA4f3g5inqPDd2KzWnRsA+t1AWNScneVS5Vf9LT/TjGuR35Sal31BIc+Rfc0
JqoEZLHG3/tVrnFZBO4v4g==
`protect END_PROTECTED
