`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0ei9UijzqtksMPstHsYahTuQrBBpjXOQDVPa2CfELOBsQmzx23PpevpnD5HUOZqM
vp6feKpR5QYgSqT07mmwRIMSGPcAvzPhKlCTgLQy1xIjVbotKwjGuHl4noVsLWi5
NxH7C1Ca2xOkVWM1osMAZk8bppLwD6qJrULWLz99B7y8+lnkFaiVor+l11jIXs4J
XtuQ/4WntgyBOT88qha9hfc7PCgG8D8ckFAxrdQGW6V5Ej7sUg726ZI1bl5oJoC5
SPO5pXjyIFkbjKtodaw/jWnEDWQliUg+NaD2UU7X/YkxRmvCP1cdw3Dtf4JXzyCF
ipumd0FLu3B+eeciGfIGoZCmcZ8Rg11LFBaUDQ2UlCZYFQx1rGAtLBFJ188Sa7OO
zUp4ekpcw/hkwu8grqTXTKczfsA0uvfdr1yx6iv6w8ZzQxyw2dHFvAId4PRm1Hx7
AOUxjXnmai2y3EecfTpWeLwa4E59vX+2v4JmNQJy3rIp0cTYWTMxgfwRGEpEJFao
wPFWkLnkXGFg3EMrJ7aPxFEsHFlZOB65DQcNXF9OhZk4BJdjhI+vBeJXmhmXn/Ts
JP4Xkz5TtstrgG6jD6D+Ss/vFhJpUqJ0CaBYpuYqqay0LIIdN28khGmVQ6SSu/eE
3D+zL8UPtpeuRIErgE/3WW1CSaQ4rW1c8JGVW7A9u2bwpaNK8kDn4HCgV2PIMfS7
YbN94nQ62TpdQh6JQW9B3P5VpRmqRm8UziD09848aMcqaQwOlHX9c6ePfIX9gLC3
q3jyrNOzyOku6W/Wd5JGRA==
`protect END_PROTECTED
