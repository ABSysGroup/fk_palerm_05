`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p8sFrYBNXMKohVfw1O3q1LuG/9oYq4vSgwcFH4mJSJuTaz60+UH1oKr9QNjcMM/F
HYoYOF+aFoG+MytkoIJIRxRTKxX5tY7Y9soDfKS9cgylb3c8I0E7s8azALpnmLJz
wYC57/L3Iy6xmTlrYn1TRni+G5CQ2BP+6btRPNmBzM+VysiGyY0DO5KggjNmelAp
B8VFM42h8+flqjBaF05XmbAuz4xMfC6SCJPjPhbfM3YQfRiDY4gFmxStxjHioqcD
Br4MDeBxN2splRdx47Ub5B7YUul47vyvRizSAFpMbpAG463Ge6/DbNJtkdTjKB/e
tauSDrNfndQgj4114VPuGYp9gtfjMphqC7qqDK/jusoevyYoAzykJdKKjOPEFsJL
1GXT1EZdyQSE4dQNTMbmlck+l7KfZzqXsETETfTYCDprdLA+WKJl3SbqFEAtG+AD
6Y1Zz48cShVGC20YQG5YE/bhj+w8K/P41o0VQ7Q+EjK5mx/QcWS9OHyH/vy3MkTs
rkENFcUscC3kOZlDwra5f/wRAX7ZhtG3/Zbh0KLfiPXfEogrcq1Hz5FNs+KXsU4r
sIXkgR7QPupX6E+IDj0X7027K6XpW6SvYTbJs09IOUosoNrRB40USWD8NyiHcz3K
Tlu1iTe3umDt1lL/aPzvpIinWP2pcllbm5mrK75QZP0DKCVKq6wSxCoGrV7aVcrw
tDhmNOpo+ayiJ7uUp/ITb84KUvpXA2GDcFUQMCEx8s2y9SXnbps7s3ysP5PhfUn+
2qKW0ikpGyltvRszRIi31i7pzxqDqK6Tw+J9Gk2pwkHQ+HtP9njQ4DoPEAY3AFu2
RCWQhy49sHcv3zv4B3Opn2oO000Df4hxf3zhCqgDxxeE+1QWTEBRU026GvqPRrzz
MmxA0hL5BxVLiWStRJghhePwnTyQvN7iHh/VMicyqGzpIVbAyR43xL6MgQB9ObCq
ESLDbcmivPQzsrzlZds9fOwupXKL0FUYCfnnGBttcFKzw6jKgixGh8J8umzh5uZD
fFnsa0wmfkULdEkorzGaU3It/09tAIKAfUjuFUkltToDCkt6y6DsDy3mQ/Khcrri
m5B5h1F2S9Z6mikfR3aRbrXD16HxS4gRVhogSmK4C1E860pZW2H6iCVS+koyrPke
FYuufyTUYBrlwvEUz5S4rrWXcHibfQczj84TYiAcDoe4Yrkab5IeMyGbJztddNZs
DSvdB+w355dtiyUnoTu1isbfZPjndOl/UTWlXLHmSzLw9a+I7alUVxBam/RO84S0
V89E5QtTn1cDFR/qTo5pRG/J+fBXxCEkNTE1vIwGCma7NdqQLXalZh7Y4Mk6W0EQ
3TFlP3RrWCNMBHh7+aaw+kvfY+HdgabIwxEMql+ZPg3IRo2g5DGsvHKDrB5s+zPC
vhjxTOatXV1uCqrccHIljdHbY3U8TkTm/l74nUVNnSnM4GU1IrAw0WHU3HlBg4+1
fCyM+tMKj1EcvsthZ7paA+IjABxrrzNuQhN2ab3w37OZ8XV/DZaZqT4lcY0I8WVX
2ws8sLHHonubt4BDpZJLdewOeF4PJyk8PHep5nxdvGYtzlFBVpTTLISqfMZDx+kB
C0z3MqXbKHHOVYsjdsTL8CTMJ0EhnEBn+ffAz33lMVPBeIlKenU0/f7lCBppFEZl
Zq2yC2KTnApCvyonozt/qaLl4BSu3P6KfbMZSUz1J1L7qmClxAUst1bFxw5iMNdA
EZHxubCxtC44At/GRKqMVqg/M5KxdeeQV3roRnG2bRV1UUU2S2bz2Qa0coJEOjSe
`protect END_PROTECTED
