`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WVNV89TFFFvFLv5GW9bHNfRjEn55yEwTXgZj/25fNPiFJ70Nsy0P69uOh1WV+Xdf
eISeGw6hRMBQuy70isEJqdGPMy1sqoQnrVxWrbid0g5Ho1GCIrVh0VV7b7mPkl2f
9pHpw05f0RIhwL80YwYpPe3SGsUwFtFpPY5VP7rrfKzZA4t6yCOf81o8uqsozGLK
fCovsXzySKwHG41suG2w5ArEkfBG233JeCfnftXkWZXZKQ/XEZRQ5qgt5IYuxg73
U3FfCPJyUVhzzAqiq8pb2u25KhaahybKXpdip37eSRyXMwSWtzQ4PbUy5PRzkF/7
rPXHbWTNWTV5PPt/ttBVeIc/Z26ebfmIFce+pyL7yF20yakTi+lFQAWcIwxoRCfD
CVuc1BN28xTQ4VoDFOE11IP9VkCh9C3WoMJN/GcpWdpvINI0I4iFH4JL5VOPwXGH
Er8NK9KlmuPaxl/aMK3es21Ve4YtF0e53M05xMi3Hj56B0dHeG6OguoARnjT8bX5
RqUZrxT0GKtOOpO3XUKvPczZCfZJ9MDSBG4YOgPRp+ZMy+rvZ4ja4G9TgYkjwTXI
rE4DeVgwzce6JAmzPAlAUkBSGMCr0ZSJLzM1Vb83OcotZroY1pa4wqlFXyh/qSUH
SJu76oMrTgAA6H+QrERjuIF0qMaJdbOEYXf8lhJnLC6R9RoA2U4ndnoj+pCKoUf6
YWkZSMVqABOY8qTA+d0nTw==
`protect END_PROTECTED
