`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OgFg61hw0VUknj4PwJCi/Cy3XksdM65HHvqDxeFx7p9sw9zAc+1VO1UJOutKhNQO
dSReuISAws+mhDizBPOm6OAvp9E8l6WqNSy0L93Jy9qFUapDJJ5NW/WsrnhnfEDx
oEFeP92sx0X9tN4L+0ctCHFnT/8YyU90KuwWIaBOOtnTQbgweqnkv9b0/1aZtp9e
EtwRX+3JtGZiW2FsFKSh3Ln66vA0fmVd9jj5WaaW/ooLoGAHSNTyvW4Y9vlqPEVf
FZH1q2VoZLLsFEPTSxbpLdSdLpP81C+ehYrQp/wz+NxvaN+DhYyf78oKkIgb0Um1
S710GJmEwMmyiplZmfHDrKmdc3sIp4JMEX+A8f4fYAEbWZS62m5rbRxwXRq3E/v8
dsUv1FjLFidZjguSI7CkbkaMmwrs7gTznbowHbruYNk=
`protect END_PROTECTED
