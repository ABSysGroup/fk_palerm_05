`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZDHYBSUcsai69RQyeoi5Q0HtV3HIP3n8y1thcu2ojmBe0b1BM3jWzc7nmQt1EMVe
UjlgTNL7xuMOfRZKJhnlFBXAiWQhXb/b3LMRT+7f2cy8RyUY/ygIJzqXosgc9jd9
v+TLKPqk2U0/0YrXyqXc3/t3DYqavwugg2tZK/4aq25Wo5M/Qty+HKPMa4yXlYhW
+Hg8gwCDqSk2Vw8JjzDqSCBEJ9+PmqNE6KWvte7AmdP3s+x4hmwApfNcRCQ3pc3l
ryvUU3+g63Y+prszI9YQ0h/BdRMGTi+0B3PdnqKq1ML9f7huty6a7POTG28SN7fu
cIoig6IRguXv2REyYL1IFDG+EeMLUtA+AVCQrRgGlDi3cQWqKGHqb+Iv2frw6bZ6
R6jF5OovCBE4TSqaeVmU716eWJwT28/lC3ey13thE0OXAj51sfnNd87y6MuhdPE3
mlADau0nZWRps0tqcTtF7r0R7q5tWz0XXZxnqEUkbiiAVDIqnTUFY6CKJy2E82D4
bAnxk07Ce8dsvMR/dRuyvPxDlY27H4Z6xuusommm+NuoCHj897NQrqNTJpxfNG0g
CgCZ9QcKkgTeUauwEFcg3ohQjBVjv6dzcPty9Wm2dT12Oo8RhDzhH1gZNHvleMEl
Pi6fmna4i7oRFFidJ9rvjK7KydUM1KEysXw7O9SluH3dWw/s5vvfmZ3Z89Hz74EV
t5KQ42fMoZnm/L9inHGiH0mf9nW9wGCV0NK6iFhW5rqifCqLLhnK2vJKPffQYAgC
h3+hW96b7cgdZrH76iDVY8mlOFjjitYShoY1Jlfa1Q0yhidT9er0O3kfEyeekXlO
O3IkgGNtbRyCKziMmS4qvrwd2nrzRwOkKUTPWBUI3terf1buQfQONECqnYVlvCiT
Z0dRVhpe4oirGnb/Q9ZtdEJ807fUel53N3fWLfnAW3wgB0eyY/7AkPaxSq8Nh/t/
`protect END_PROTECTED
