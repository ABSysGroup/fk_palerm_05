`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G4xW4L2O0KpeodBtxEDiU3nqd5lJdsjH2oeWUAF6AiltTbJ91xXLNUHnj5pRu0L0
2b5xk8HY3oV+eee//m4DwFZSn278XjyO0WNxOva9ImvHEnsF5uIFqXy51nxQ/GW+
l4WrLw1Rx7UPefeSWo5cZW+swhZOIspH+AmZJwGqdunkrCI6zTsPPVeMItZmsNpE
30vA/rIOePOxZbyWXvY9c2xvRDf4DTvhDSpQqsNV3r6FFrR90+A8mk+WOlStlRJO
OmfTK2B/mFppqcmTY3MFqtZ2eKCrq4uIDaZnyl3HaLwwTFKtrTDvGs52D+8gFDeR
HPhk4ILBIXzoH73/bUZam+/NGK7w0nGE06iF+XQv5UmStITAtF6K2mHGuUvy7wZW
ZTjxwis+KvjHDO/1O+ejsqrDf150oZaArVePnAJ8hzjnFA2O6+9ehLqvWmn60IAn
Cg5wPy2WGb8MgkHbhJmWW6v+iLlUIwFCrHhoFQtDb3H1dQ9bK5G7Pr24Wpod702V
XLSIWaNJ1z+IB6V5zNgvrVPcC9MGyUps5UXm7w51t0IlyaRP0HiWdQjRGQLfKyF+
oo6HOtZM1klZPsEau8dW8Ys6NrRz//lD/SjMg+mAPCpMO7ZXt4+GwnbRkkVxOGC6
gu5IKUZS/1SUT/7uAyHFLtWrsJ3znpFWiWcXwXQLvNg=
`protect END_PROTECTED
