`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qiwRC9x+cPfI1rOj/nLmF+fMQaxiBjaMoA1kS6xiT1YSLCfC5rSmjO78PZ/kmxjX
ZfpfsA05df+T1pZmWO4zSjUTag70eSUB7xcFkYkKfN2s4qJThmosC/jOAckIvq3J
v5BzoaiLcMuL9XxTyfEfYb4cSfCwNEchU2Iyk6vEb+7Ju1sX9T8e2amKH+SkL5Cz
Q2JzBM++SkBUANoEQ/+K9CEf1gL7jqfJaKYETcd/TxZtl4z+hnutJgpWaOk/UEEG
o+eVIYSnep4aOFDm9LsoPzO4WHg40qAi2vHdk3ouvUJ8FOJFH+nWiQGtoTPUvVQl
nvYPioD0Wlb38B0BQkOoqg==
`protect END_PROTECTED
