`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rmK/IBaLcTwg1hNsh77q895cYy/gltChuI5XnSKmEwZbI7AEm+LoiBkujLHu8VHl
lxaM/IEZziDPv20gsuGJGY3ne4gOYsQDFmvtVeeQHI8HDWAQks5bjTk+21Noe7SL
30c6s2+WMHfGCpslOh4J2U9/7vThWqkJkEB1MJVdr9RYsIivm1A+e0ZfeySO53Ew
5HL1J40R93vcXbiQ+l+xBIlFcjIfbi7qlQJtYHXWRQHq/+tRu6LNyznfLjbwRTvw
IZp5GygzPewuAeGOExt+uJoGMpSiFgSPpETBz/ylAi+CaswphhCteLrFCIcV51qO
rxr2xSaqN56xZsbcXwX1n19FvsQnxZnGv1QqGTULGgJ6kCJIBPpDz5+9+xj2FBmB
KNT5iirEifIdbG188Ylz02obnuakUQNCix5HGMKl0REEatjKdD6wZgHnS+shpEZa
owgv1JB1y4kCXw4etUYayxOhdUtSV7mS+zhZN11/3qvz0fAEPpauNB4VwSreZryL
Yv91K8DJFCqHMmO7zv1cqPKIZtriLBoc09qxD4fm33HRDnq50Kd7wx3yKibSG8Wc
FI07XIb8+9ZTsh5KZm08wkKyUAo7zXNQ71lXwn3At+Q/+apTpil3yvQ0YCRjZ4ve
r5JROMHIGaoMm7kq4UREHRzJGwntlQ0Yq1KRz/NJbhT6de3qtb7CW/6owtrDpRJj
BLtnn/s5YEEYk/7KnVo1eYiTAUFDfMK9wmYd4Jf1d4eQVcQL71sl1CiHrB8dvXgn
rd1l/U1pYm2oirG549km3w0hmQ8xKTkvd2Zu970Stz4GnzkFSKlf0oVN2eGhwMDo
sByWxZfBjinVkkdMMkM95mZQWWQm2xzpYYXNxOQWcrDc8HVUvif1qVMzardUfRpL
LRv1u+Ft/N3HaVJ+YuPyMgCV2/tqJFCvK46Ps+EC+pu8rqgROTPyk4f+CF2XRi88
SilQ7SGq+uR8hFnOeYlBbHtXU/Cz60a3+JbYBkKuG+JHOT8Z+6b2UZ9bI3/Dpg2H
8XYord/7s+//e5y2NBcIPBL6STT7fkUXtyNecGu4pnhBKaZNMfEGF7oYo1GYhSQe
LS1zLrSfX5xGVYKF1hgbapJTcV7urvAKBVihQP3LlWe4/dZN94rm1FvEDlZMCGvq
PNpNdhnbx/Esy9vLjLHvV6silBUmXjHOlynTh/4E8gXlIShNfSEy+d4eh6iRRV3x
jZVRP2IQEHW+1LqZWfe60h9bQEJc6boBG0109DHgDI+Wv9GxvbKgVxHaWRUfMKts
hlRTa5P+HiAuC0iM8CLtQlWMMWTy5RnYDHk//QVh0/XzAfh9cmi8v31vZ4/D1my1
kHqocPO4o6rd76YvYppgus7i03HHbfg8VD8Ji8gYsQIpFEkev/eut3pITE4CVA+W
MGrPqE0L6yi0x1UkE/RUyVTHsB3HO3lqt9lN3htZDCptZYLO7KQVzQ1aWCwo4fwP
VPBqdYP5d/8Mnxe2gmUeLsqHOhJXUWwpOlZtIyI5cOm3ECazeYztgjStuo5z/Dzz
BZ8h7dTmqeocR54NoW67iYZzX157+jMNlJA5d1n5cRsXPLDahsBtRobmBEeVMgne
ZO/jdj3fQArh0+O8O7697GySQd+T8GKBNg7Io3NqwPLFCQ8USaVpuj2/UPGp4uNc
gGAcW5l2Cc4cArxKsAFY+K9V0X7csCKpAsNSwFmWpn3GkE69nNEzdBmh3NBZFDcx
fsTd29CeTu6kcLDppTJ17Xk5cmWNSrUPZxOBlCE9JKXT+QPNvdOCzKiynyrw7rNF
/aiwgIxlGuaOcHdxq7q0MCA/yDDG86o4oO8Qwdq7v1eEgF4vDKSNmotUiQnAd2h1
fK2/XSY8mhdpdfcd5tI0usSahrjGvkyPRWSJOi46L+1z+kSGsNBij8Jlh0bcwQpC
KDgCJUqAc2IXsiowVlY/9VAfDpNXI/NEbQzIz5RmI8Mw7VkjwPpRfufIh3vqCz+U
DOd+KAJMfsP1BoQY1+x4KWpYBvtoJhMpm6kYTFE+w2B0Fiviz+MOeh8WoBPbIxmo
jo1+ON61T6lTa9pdZOccSTVD3B/gynwOWHUWB/YJc3Ygf6E/x0VpN/va/taMQvE9
wrCDPv/UBceUReThnnou1esOzKkakC0TUSOF07d7Xpvzfv1ttIVn2Jf1tZYMunKN
Zknv1BiQjdnEWinqP25cYs1WvCQDWy+F0q7f6NopsSqtXw+Q93UozAscIZ9o52KH
kpyVb44DW0+kKY52Ya+VX78a12saa1FC4hG262KzGySLxIchPy4nymqFvhsSAa4o
SNNhkFrUV8c6CXYgNEvYVCTTlWBTFbfDy6pdBF450lkE990yfyw51aGkn2SZh2Nm
tQOykHLDKAobHqdmFqjV3fi0aHMim3BAaTBJdvnG7KFORV65tv7RHlByIjIMLM8N
IAajTs8hNOe5ykhO7/ATs+MNaflniYUuMUpB9yQ/DAqyNH3Xcnsl6O/hOTpJr6SG
uz3W9dmyDlbdMdLKwXkkJ3meuxKMJ5qLvzfsBmcdtnbObE40g0qGWnCruApmYVwl
AKelNjb2n+yTze7fcfcPbLaP/py2kH6Qk2/fRvRNsCuyZj43KgTkEBu/eYJlXET6
q8GG3iR3xjy3tWf7KF/oOwn9BTZcYWUf6GuPc/9uEtnGliobPZ7jn0i7TxqE9TKH
gWF3kNlRYxYipaxBcgRCnaBLyL79GGNC3L7bOH+cS7bMJb0aSABv7uXjTw3FXvyJ
TOAxrxIKMK3uE7iHmbHvp9U64Lqxh4xVB3rZCRl9XBJC02FsCyQs+YE36I8gn7PM
fjPertXTfd4NCDRt+S250fhv+G+IK9omUHsn2EfFjpt+8RJbEqNPzp6rbZ9IV5Jx
ITXPsSfmr13mGnR2f3pUaCqRvfvFRp6qpLRhdGbwS69Du1FYCpBdTheryHiBCAqc
Uzu+5MoyzEWZRiJl+CJtOzIjgLqdwgjAMG4+/WldKvZUuvwHFOlmjrpIdtJGU+b3
aARvSeeSeSkxG/tbSZ8SeirODej5ngHIuBvO1Q3BjFN0VbQZohhp/2aeBAfsxOq3
6u/rU0LaYgoDeFaK4zM5oFbPp2SvZyXMauA7myU4mFwph/SftDiJPsK3JCuzmA2Y
+6FKMrxt5F/wgo+6lquvvH3l0RQ6PplP8OYD+kZs4KE3R6bHqUS3hHixKLHtYq6p
Na+4GX7i6rVC9OEKN2NrmMU1pep22u58AV7nP7xLCmha7x6v8wdeiKLTcW3Evo9x
Zk8ieAUsXtCD/7FQyVY26uOx0k6Z6ZtBN72qVDemROsCOKkk1Xnxk+H4y1lmbM3B
Ev8aWNvwZrJ03bQARmn6I0m7Nha9lTh/9xALqKoM4DCNlCiDf75O89+QnFfQLJji
F7ZNigRHAdPt+jFG52SXBAT1cO5+/ZNLP1MtjNaIkRqBaV8iIkGzaCMQSlM2wiM6
iZQt80RvvvF4RioJmtDGOrtuezMtEauMtC/P6jF4Bmgdly806rkjIy2xoGNhx7bb
W1MBo+I4rKaGJ9kJIejfbwHYpM9jc/ayCBGiH5tMglr7h3QLRvtc2Hq+xuX/pf56
zHjogAy0Sbs/RuEy9WUp5bU0dzrKtuhzS+bjZFR5O8L/RDHsKn6ajBplvloTKJBQ
2KPcZWxnhJxdXBcDBPc+pbRrYU0oirQY9VBXGSjJIe1/OJLKbZbTpwaD3qXQOC4F
X/Sa+UvLZgDnYuZGdaYclS26qNz4vYNrbDv6JYBm5SSORSiUOmr1sW6Okrn0EYJB
DJYYyBrGS+ML1abF0Ff2w2iiYj64kFigJYLqoM5u/hdOZqjqe2Tpfx0ODu3Sra00
CdnqdiHa8Adhq7UzCh39iSraOd4xConyGv78sIjz04sOD2afgl6QyBM0cAqpnV21
HLDJPUTzaDzGU+VNz+vh0f3avHDkhVBPnZKc2GQw2yvy+xJx7JB4kwgKG8glrdED
zrv/QuNRjlzMA5X1yIDO/Qs9xW9uanvVi42bF6a7pmgBNxyXxY5JlYigIayuP4VZ
sIHkN38sPcsQm5qsey6qjJQ62xo6gnToztBQA+pGv07evl4ZWfCLgSDncRVdhd5k
z+X9H4KhfJACsx14cgDGKzBkinyhSfhib01XQ8PCtE0qpaTvnAgnkQjTz2AZRoYj
+R0oWKBIPbm3K3RHhsDYiyam6FP1RM6udGms+B6DaYn3dF9w71D0bv4xC/xtHqbE
SeZ85jySmboST/Go05jpa/40b0UT3kxK5wsA303MWknfwk1u7xOnP5xJLS2sptj8
IZmIshGDQiGyuJ3az2xi469NlP4d7OFpJUZE065iohJctwSI9HdtV9a2RornGNRc
kRORnCG2rFKO4TTx50ObPL0+fNUojHurr/CdO0fPgO+QxX4QX0pHC+NCUWprhLQc
xk6VMYlzZnfOM/pekyhN+wCQD4hqysMHGzwAboMLkmzs7XK3ZKBs/LyjdKwg3YbI
avdvlnp8Lyq53a16yGYXBGOcj4Fxz+Tg55kJINIF8DG7hwZklmhKrX5gsV9fWiUw
9PS+jsJ5cuc2EmGITEyXv1fh20tBWADv2EXuLaxjbPiFOIY3XwEwz1eLw4AxR9Pv
8NK3CJYFlPn10qq24QUfnbrv+CcJ4Tidp1xd4ibX28Xlw1xM1S7Zkkx82CTQOPE/
BUkxnvvQlh7MqdzWFX7AdBsFQhyMH7b9pLWQo0W+YGog9pqwy32XfetVSq2U03T0
1jviXfbMXrAm/m+MYErUqsMSl+K4oiZrhHzrbWe484nvezZIsrDauhA7E9fDSZBP
LY8IglmRI3FFmEy7WrIAug==
`protect END_PROTECTED
