`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DCbWnq0njwh8BeGSOJceVyxlgMFqwn/+Pbo7PLoULL+OB9yjb40kHegCXHE8B+gq
i8kvdyS+mrKGE6t9kec7kcvDmqJEL98f11CBytxKfF8iSItpxtEs36zUXLkFog1x
e6JUReAKvCEz/QqLtMyKB3G1Iv6mJUCUdo4YNQFkXAq1ifW55V6Apez/eJwLzzBN
xEx5S7ogisFsQAGjWtoemlUhSSPHVDQkEXhyvh/ppynoh8aU8qGX+hVlP1NIG2Ew
R0pre85F4Qy8vYX/Aq4KdenjfEkh2FPAOnnUxU81sIYIyCcKHlUIJhSSGC2soA+d
RdnIO5NVHKOnCq1Y3wG+F415Up4IG65erltt2vGczPNZ3cfpxRcVNkfbEascpZfN
Ao3mnDeEntAWPTcFsa7CEwAH5/YdtOQMNKnvvkOtVAEYocaZVKab/xCsl4E9m4XK
rnHB0h1n3OXWYENl2UUbBZWWjGL2XrdDU8z23xGyJ2+Fw2BuWfmeOuKR1Is6ZyKU
tYAeOw/Q93tSppsQxLPAGLtaO6wUOAYLENJPTEqAtOk8M2vIxYsIRZy7bpBB7fme
3xJQtKlCybjevDn6agAfGpSw/PdAP0aQJmkIAIvcPVYc6AZDuGEQCriTZ/TgCRWW
JZjmaQaSByxFe4s62CXNIkJYgQLsW6uWJ2xtt8BkiKu21kKbYMSHw2a17/f+hQy9
zmXlSPIl1/oIAbcMOYTAtCJk+LVCcselBMXHWBwDwBtKFbi2IPkTDgGCAjaydsAY
WUQrxGvLGgHcBk7YyYE3rA==
`protect END_PROTECTED
