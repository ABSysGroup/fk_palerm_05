`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nA0K6MRLuJAFTPp9tfo21n8S9IlhLU20TUSzU/aehgbrDYdsU96lPXTTL2jyDlrJ
FzVJxV48skcA4jPt/jEuSwY5mSev/wFcev2Sai6IumPTFLJFL9hpFjnYWwCItDpE
Hl/Ma1fD7YfozB/0M55nNo9OLyN9/jPbIFF6jdJY/Sms2+6UaJ7eWItxjXnW3PoH
Q/nx+b1jU8LV8GL2gJdx8WKHRExpZSNyieERrOVjJsNt/880/7JciKnDksPVdP2E
nlXFUbhA3ztmExXTZThwHLScuQiRw1B/1fAC2JHeJ0jcpj4I6MiKT6ejO/dBfd6s
ydNA6E7sQxnvMxJKWuO9rhOG/q0hGBS1y0L0BmtosKtaeQdj1AtwI6Hd0OBRVMj+
iceRZVz7JhZVakb7slZ3gjI7LX6iHu2JbpkgdbP5jNxOfg76ZjFWe4pRnSMhXwD/
zWUbLv7sFgX1iayjBszZov4bB71b0hR9dREiaIEglNERpOvS8TL1XFU2KotBwGSv
S5OxlHcpfu7x90Ht6Pb21kTzSiWF4jqqmF3GnYXb4AZxM815wIuWwf/fxVedmkjL
GpVjbV8QvaphUkACER/mjEeSX04Vn01oZBIF4I8Zzgco94l5NQTxdtfjScuru4ED
nAr068mr8exef6FH7kXCkh4j3vIw7I3saAoDeYHqq4MRModITy8BLYToWXWygC5O
EEvAqaEc0KoviPS5EOmGGOgRvhkvAHQRSODMtfNwPNydTxH6JpV9LEiwGY0Oz0JM
VWtAJQyIE+j0Jo1j1FxWcnrmxzguSJU/bnRExeQLG+83bdUi2tjY3Xn6vOZkZhYB
JliO0kf1cNRjafCpBtUMzY9+Cf+6bvNlNVnn8vHagRHa9cS8orJOq7hQl3OZQwlA
T44atET/txUfrBLORQlt+uIRNTt9YzSyBif0ltVrs0gZ6YWX4BOmu9w8lCxPU+xp
GcCtN6pc6JwjWewAEgclbw/w1SDk+dQa8u0QnGRhZoYjw4NTKuJXuvSXwTEKGO7G
vJXaZz+Z+GdYY19GRMgRY3/5GVenEA/1pRTd3lGwbQ1jFt1ZYBxFOKH671I4MPhc
kuY0906Sy2zwdqJnCGZNdEjfDAAB3GLK8Q/w+7UsJxLhXarug6hqOp/mwjSnAfIC
B6E2ZMa8DUC2AFiexuEI0zcZS2tVUlCXdYejcVCgHasEP7dU1y8yM2957yaCqGHe
apuRO5Zo4qEpg2kboP56RtDodEcfRc7qmt+rqOF9PU+PwGLMFq6Hspx2ouTlV90E
pkFJiTsSt9cXIRAL0HDAjE/blqDPE9y+S91q6YAPmiPje4VF5Mt6I547OtpeaHt8
nwRfSwv3+82b/dEMP+0tnME09Vf/CdwtTwsEPAWigwqkEuazANrOmDrNoLespG3o
6W6h9smS1CSrbuGG49WaFDLL0l8nqDQsPlvVauqRKLU0q29Wr6mwVigmgkEoxAu3
TtNsuO5f70o3ttNz2CPoErGOsAo6gXdSKUbaRL6FVljwoWIJbMZuDexc70H+z5Fo
37rhQq2eK32qfe+4tT4eYN1NQ3p4+Wbk8AclnY50ZK1qMUbdIONOubnk68BWju2/
/c9C3i2fgIYbANGwfPJ7D9QJtOOg3dDYQb338MfzLZma/gT0gQTrWsDNvcA5JhOX
hwKTcJY1sRDdGxjP+HaqLqcQ6dYVzAj//9yB0bZN/mABiq2qVyEpE1WR0gxkRk9d
0hqMRQNRsUG8F2hfz5cjvvABFlHIZXqyH3fB4obR9s61kAUmijFnBB1EWHjMWtap
xTqpUSzEvEDSxxYi0OusYe5pfbyyrvwqHpRkxy16nYnGAO1cOmQOQfb01RdnpBSI
sq44x/gcTK6+H3U7uJ3zc4Jcd4550gkGPjN8PNJdtBUmwD+YbaXWBHl06lrlnZi3
fao/V5pI81YmPRsx7muWkKQ16044vZwOh4Sv1d9SRQ5dzqMFmkIE92OC99bNK+SL
Ms8xm1SxG1uVAxBs9Tjn1OUWdQJy79vvta3N/XTkpqBGtyJ4Lier7AMmfG05yRbd
fpn4QuxMdK0/M0RysGdbL6jl/XavIfBJPtnNOmT4ZTQ6kDLvoE7Iz11e9Q8QsttC
wWEFynnJSDdfkpAWv6wYU2VVdYBsuafnBEucu/q3Iuzz3awRT3BXSzulNtxUm8Wz
LJ0HNJm+Wr0tv2ie4DvdSNpk2uwCOosx7auhejT7Y1TO/nFU0cNr1WMr9u+ec6et
cWQn9QIwSSO+e+/wU4tnaBiTFYpcFEn54J6MT0Y+FO3dH6jpEwF+gbZamisyOBbY
PE5UyKeM0xU47u1M4fs3D50Gs543c2uxWBDawA12NUM3L+LyO/g9AmcgUnkuAG83
2mDmtBxb06byOF7Qr6o/A/Vqrtntgn4UA8YjlPJOPDW9C0INQULDlk65R7tuLIFM
fO2r+7R0S7A4VSup6jkVyURzSxlOxPbe1HJdPrwY8iJM+6We4fTtC1wa8HenCbO7
CEh95XONry9G4k4YxSFsPvxVL8fXM4qqhy+ILuzqR+TKEl/OxYzOZ/al8D1wB6Xh
2iahT9L8mHLU/o0WyIpi2jrl3+0er/Vs59I/+s8iG9kHTOu0V/EUIIlOYVKxMI68
BZV2SFrJMJPzNdtQ+w9uuQuj64KX5AYQBge9ocx7Lf2Lg5sRGdx9F5o9WbtmGIhl
0QaKOrSKqIxWy7/mhvtb/qK97UG97b6h+SCE5w6nar0VdYsrUAN8UR2Pg3uuiT0t
ypSLsi7TdI0RQJyzGTTCOakAakFYYOqO17g6UAc71utme9LOM51SUlXn0o5jI1B0
1dHnIeGjp63XvEkjxc+7sHnrnN4AXq1ZXdhCu7fCjhnG+H52QdDmL+rhBTZEysi1
BFFr+FUI77hRB/YliZ9AWXbOAZZtMzqBKEXNd7+2gj68XIE6x2ivgkB1Sk1oMnXK
7rK2XDq+BO0UmHT7E91emw0mM52MXTu2leSfUlVPV/10Ffe9wZeqWMhfnyYyzMzT
0V9yM1I4TtbZnguf3mHOEHR7Cy1QhtjNzEx4eL/v1LMb8/SPHPN/e3qMv38AP9A0
u5qOXdpqN65KlB+LN3FHRpCeA/MCsp4BhU68fbltsXc=
`protect END_PROTECTED
