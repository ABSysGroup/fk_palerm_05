`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oqt1ms0yWKAUyL718luMwyztHrVSvpwmbGpaxwaqWAM+I7utIFRbWpDImPrc3AZC
Uyt0tRF9utkUT7ESJVY3Vdw0GhWSnPTbNRhnrnN41I9m/pPkRo5EZexmyGeOJtvt
WwOKVHa6AZqYkuT5qNxpersKPO1m1oLYaF+9zQ0qscVHbjqR5FW5VVskHkwrSaZw
Zd/A7cHwBh8UfPNabvaN/qeJSa1DSUILq5ujpstL3YlNzmUoaCnhTuCc0UbmVYrL
DFuQYOGuuydKAncxsSUFbFJfVTJHzKwXCL3U+/stjhE5jeYVWwsbGoIX5T97K4Rd
rkEECWfa4hzDjOOGQsm7pXAEi/HCbZL+SpDN9uP7+O/QxOSvUc3uLJ3GoSgtbyHu
SMoJGehXCs8IDL5bJksyuZir2A4NR9ZXndc9TRTlMdh6yLxZa+rknkNCmaRV9dxO
envf/jU7+2Uk1Un8uZQ+Od/TDHOCqvGbp0mPnFaDa0atXcjAG3t+qk29qJffwgoH
X1qwa5uNoCcrafBiRO9r6gJI9eq02AJNHEaHN8RJXwtvKWuS9+ZyZs+891qjWfHx
3nPnv20gswRAz6gqZoh8AjX5YZ/7sPei5CC22DIaORBKgwXDZOnZktJ90S9V4zxd
5zMOliQnDUuka/0Gfo0kZO+H00Eh1x+ASyMqA53vdAXMrnpnujnN1j9WTStA/d2D
KOt1uEIngFTq4eTnEUgxXb/LAJnvBRtHAwRIiNHhVJI=
`protect END_PROTECTED
