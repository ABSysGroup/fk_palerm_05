`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VnM6Vvgg7kfRFxxgjIuAZcQJN6bawAsoOaZeJ5egWnyAqGoDV+iStZeuApI+AGH1
hhf7meEtloKHH10z5g2CymfZLronDpbjTwo4F5I3q1CgTN/CnWydMfywpYlwATl4
EcrYGYYG+mBSPHmBVJHjFRizw4mPeBeKER8tOIjuvjIdGZUN9/ZUeatnIRchWwg0
VHTa0yr374ZqR58KwajCrUsqWX9DVN03ksCES7jff/GkjAFvV92AziCLOH0RkrlT
j/rT/91F8Ui0ZiPH042p0i7XMB7zxxvjReK6tTGUIr4fC6D0lmntYiZzbPUcLlT4
Odzq2oRjEdMyv4B7Iw8QX4v9waU9CK0juAUjhLhC2isewk3P9L+l5GS2DL8Q0JqD
xGFtX7PYyj6ghZawSef0Yw==
`protect END_PROTECTED
