`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1VfMK6OIk0Nbi+ZbiL3W77b5+1NZZJrYC1ka22H+DJO38XVKBPWxLyobMG9fYNfM
sxDl+epTtXKcnpg5AeYjzSBloeGvkyA6GTQuAeTOxkktf4zGHAUToEPomlPdgDKk
7L2Qog29U+afBRltIC9vKaqKiBSZOtS5xc2+VMqjdOHDc9YpEzB3dl/ZzYO+X9uJ
XsYnJAdpOqFO7to6aKfxkNT5aHPW3mM2G+bF1f2l2fzuu0zx15ZyfFxm6yI3ar6A
L4XQ2mBxnsoF6hTq4ZN/nxjaM8kn0m0y6SYdp1QkF+kLRz9VadSLZuPfE3IVewol
Xtcit0+kQrUDkF4Wxyeo/A0DMTCMlJFDmquhTcvGXCnzZCsbIQKl0rVspWPhGDfU
fXctii2rcBEHemb25n/ekM9BZFMSv8jOUif4xzaAZDzWhaZIvDOetk1XO77Grsd8
Cv6tnFzdZHQloHQmKM11Z4G8Cg1xhYi7nneOwxQnzIJqSAQ7mxoVOOSN4FE8a98E
QWM4N8BPWB/gZ0u1ob00edVPLGQHemzWvBTOJJ0ro1IIYsEb4FnEHmusAq+U8Ee9
fj7kVIdgAboThmlUZUGuq0kT5qtFqyzeXmBomuN2dnuwBlUI5w7VDFsAROIIH8Sd
3aj0K2vsC3Muc926H1DOskukDePPyQrFH+MljLRT8moC0CR0Gvv+KAscFsSIvc3f
sr9f3E20NdRMF8wZou2L9AoaJB31nbLqcxA1kaJKaZDHzvAgbqa2wA1vh/XQzEX9
NmMKTID45PIMF9ld81kU4qmVbr0qaV73pwdN4UlvGLnT77+CYemdIXOdr/59ABJJ
wEYGBwRhEK0NcCFH4k762w==
`protect END_PROTECTED
