`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P4cBbzm6ozXSVBwJHzoTNA8Qv54D5VGz3mfN3nRHlrxaRpT3tvG9d/c5FUKUpiqp
/uUrWw3BptI0Po2p8y/bMc+BeuwQSSe+AuqmM4hQnFkG8qavkOKmZnvzuE/bOT7d
4I+B9JfTg0QBMzmd6shXPoqwdGwxzsktVwGtIOKVK0QTKdAvoU8AoA7xf09JSlbb
RauTh81tuEhq4Iska7c2OSAjaRvWI1eg/0qyTffbRJjI/kVLBdLta51MnRde4tEY
1VJoI6una7yE/nWumbXFui8CGNQ4oCD7tGroz/pGjMHh/in1z7j3aLaVUPRDTVxc
uG+9K4EoggZqJipCq0vFpVOhUHrlRFQ9c479EQDBa0ZF3Hxty7+tHAFw2pv9FmEz
Yi3V8RYuDMhlE7DhyHqYCkGlzv791sYHoVlnLdQ15nw8ABvq6le+cRrYKAMB3fPl
3USdvMpc7m75umoJerc5go7wnQ6o+dpy0DP75MW06Fl5uw45MXKJ9wgPCuQqz2Th
s05TllZSI89OFCwNOg4jBnFOQX0EtY5OMvfuHyjN+9y3nCD5gt921NEKet+9Yyfr
6UTd8T6m/UknbNpu6Tj5dHyCpCLS0GNZbtUqFsRkcaxSyR4KtcZ2ZeMt0/+gOpXT
DYKrctGWsnwbXrejWKRvO0S0MhlPKS4GKg8fdFd3nuZdN23xLlG2S/BKKJFfmSII
7SQs2Nzeatv7zsfw1Y6o5nA0w5bV3lM0h0SF9KgtWB0UbxJIJtMQ3/Q7fQtH+Z/y
VICEIPOvhNrguuCm7x+V2WjDQdQ6S3Or8W5fzI9yQs1QkEpeiTs6K/bRi9pmNhSC
z0IxrYXc6pNoTvVq2Ox4qoqgM6BoKBatjNTUEI0oNvNFlwzbFe0j4RyBi3TaSyDS
yvXDTCVnkqQFKtfxAllm/BVARtmH38unget/JOgDhf1BYlAViDbCR1uj80rxzBqA
vk/70v4O1d7LLKQFHmnetG1oowhuyDyVgI447tg/hJvhZsNAzWzmM80rujy5OGdM
9vE2YiUPzDBHU56YmSeyDvx0F7wELeTWUFGDDizHBxUyCZqFcd1a2FG3F+ksmABI
JnOJOkUdXWYJZlsj5ltcSa0sDvywe8T1efGh5gELbojnzVNGUOwx1WAUlZPMJ7tw
v7u9Faun+ip7g6zN90azm4ohitLvKCIlLJ/tSKvd/yvnClXzpYYhRRtf441mW7gY
Klzrsxu6OkNemfAOm1vbPKTJ8g0a1E7vnUn4HCcpwxiP8B3+vB6Zij70sW2XeVUz
M0VnKs7B6Ki5K1ZAhUnLtb6kUwZ1KonEOeBK3zE4UiOac4OFmTRpNhVr3Cv1IfUr
`protect END_PROTECTED
