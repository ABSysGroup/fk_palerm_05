`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qh0k2pdEdPNbrsn4v4kCdKWwKcX9hov6pWO5l6eDucv1pLuwlkFfbaXgJZwO5Y/d
KrWRW2qy9iBLuA4SDImeZnjWedKLZ1KNjku0dYO5t7Aatc1YfUD+AgJT/4LgGGnf
unNkNK3Vh4i8uKbg0aQlI3JH5mXdSL5VsdxFTxqXGZNN9+sXiSqSqq0isqojFe81
WA60EmnQ7jGNhfRIsLWIdRV6uO7ELw6rfCest9/UCHqhhxOZba3+2XdPGmjUJ8u/
rv+ezcjmLpa7dQkSFqLBNNEj7DdvqJBTCxNi8M6pl2hBYFaBR3rog1e5sn+uLpXa
l7nKVm3i8GcJOHOj+AkPKxhILUXqwdTIpROMZZbdpPqpDzLZWohKjy+d4AH2sMVq
0EYNiH8Gr91DnUTZKOum8XdLe5UlWz1m8zQolGBcnsv2+Em2Ig78qFVtFdGQXI+E
Bg+l9gvowJTQhG7Iv+Iwlsvi823FxPLvzqJ2Jk2NLAbGg0r9zE7MwAplI7hxfkBI
8ucsAJY8Nf6m1mTfqmSK2GqpOc3aP8ITyPmRR6TlS/yOKBeTvy7Rlcm4QdsHL/kF
7hfAzTIKBCq/Ga0nIVqxjEu8+gw6bLcy8vYlv/SYjdMqAyieeBVrRqPs8y0hRNe0
nTvxM0j5rH06Ho0FLwdPXL2z+UPxbiscWEK5tzKiPWVuWloSKRc7Cv1PqPwTGSBJ
p230ECo3owUM1CzbtSzxxlmdqb5d/WqFaWgGh6rC3SQ1YpfN9bPikGamXTMmRzYB
tGTkLlaR/QeiPZILYIx7f5YmBZ8M/VF8GJsY7YHWu3aj5iRrkZVAY/ibf12aX9nt
dE0BoxocN48xUKDLWIVCK4bsKUqd5tIt/Sa1ZK8aY9dQKM75fJNPlXThZm2Z8Lss
ubq0PJCOjeL2SmfrcQej59C5ZNM89VxvLXInQ77DTeNJg5PzDBmGIUv3LicjnrYf
92P8923fbGo9P4IMfGcEmt2FuvYBvb1OQoILEKuFAAMlk+QxkrkpCFYyqZrnQrEP
ozbZKJowJ/wqSRgoGLEppezFx2MfTjA/ThXD3D3n66Tva498gRTBmwd9d1jfHnf9
LRQi4bIrzlWVGM6/706X3vjqVj6u8akMCdAry/UgwHiOGLLOHbx6wL9bEPHgSPBd
Q3/hpl01A0mZxLEGE2dQC9t5v+xJwmzcrU7U5NKCBN/isYXj3giu5mC8j3eL8JnB
gPfmFQ0HeYMIkZwhaWO8nNQV1KY7ntR6A3CfjKOM90mADzzLlk2psk/0v1k5asOh
xDBENcf1E9ojJ1yPDoyGZKXQoWVUNJ22tx1rHpEynP6Hox6NQ4iYHiwCzF2tiOTB
mFCbqDe+eFuJJeZtfyL97C0lrUG0R0yhJ/i/GQslfITuOorbE8OqrizZkXFDLLgy
06A4ghctReOX1S2rCm6U+9yWiCNN7MCGM/c6JwYZsJO0JRKEXlpXOUYB9IGuw/U9
hyXTaOdP+ksddGTqPhYHu3QyTg05yLMnfU4IBpHup8/4WrVwrr4WFnAms5Q2M8i6
rWSyLY3PqbkA3mYjGHD95lNuiXUpZkwbMEG7Q2TXipveiu4ry8tH4OeJSQl7ELe+
wgZy83GP8GBeZnQUvdUJD2tPYALQev16fyNVKqXJtqCRAJUWgnQa/xA8IGUPVE9T
E4ounJ9PzYONrKGdiCrQKcSd0QI6ZFVIuPErfqKLNqLg62DRgh+al5aM4EX/UxF0
jwCYN1RZ6ODVJcKlPZQpu6r98vBJJJWV4b1rY3lz50jTZKvq4WeesJAempTrAzq1
5WXgBByqNxaDpQ29PV6Zih4L2TUMjrGyYkvs5miT0kqaq4f0BwOG+NE8exehENkJ
9DubWOfKsL/A8K7Ho7i5QI0tmmBkbSrmv+M7Cx9yOcR9xMAC+A4OGnEwfuT/pKTf
9JFB8xEseUCSbcWDtWTsyWJvqX5xA8207C8hLhfifgPZOP3ASr2q9eX3Ng/phTJE
abfzWDrE6Maig9dM+ch4U8tciLjPr2KihJb4c4o07ZpBY3Me4xB2B13zxFWg4sbS
Fl1No9a/EyLEkJwIFdAP04se6aaemQxsdf0Vi/f8p7yP1CTZKcOVe5mywoR4lP5c
AnQvfTw9egKvcUoeMffMkvSpWvfqcFg+DRcNsQFuAqX0aGkhklsPz/LT51BtzhoW
X2SkTLYa7PRJhydPtMc57RkXtdXfTc7J9ahmt6N/i+AQoqjczCBDw3cQNTjefOv+
k3NXAX1V6eZlYnjXcf+IkWUrxpdqNAvWJixoUafUASoh37VbaTPo0a0v3ke1uEJc
MK7VFNV4gk/FFIQ0lsLemlZWKKP7ta1kMpqZlmiAkUQ8dJX0nLEorc9epgZbA1nb
VCY+AIhTS1YPTwSfz8YHTNon6keOeL9stn7qQFnPGiRY6L6DMyxlSc2ACq4jGXnU
NUkERFl7gOS2A49It/EeF3D4Mv6kRI6EZFc6NjdYVVmUEzm0XzO8kgG71OxUkJCk
meuAMcm9WLAxdOmjwGZ1cBJAFPQgudSzSnV2qjXaRFCBKPu2YpGl/6pEeqckUtM8
pJVwwmwiyeX55MsA/Ymibts+3mXbtUsDMTgBQBOrIA2JDDlHw8+kadIUsTty4Pay
5B5tTW4dLS5a55yXui/B8SKx5Ys4LvVpH9TV8Db3oxfxu71lDhzOyTB3fug8ILgP
OhaOAxRl0h1IERw5gdyH1nNjZaf+3ZwXiDWyJ0faGFyiCFsfHgq57wyLsdR0slWD
AnG+fQHjnkZPvUO9cMMvnFWEDvdzcw0FZEbvsPS9cLiRoa9di7BrcvtE1cGhhO/L
sSmAwz7ryB/s587yPNXjxK7uVCQ+MAckje8mwquNEv3mP0/XSh5pi6jHe6L+azI1
UUm6jcBBMPlFoiOKcWjzOMTd2EaoLJ8GWquh6d2scUgGqN/LFcO26PQp+3MOuxXp
Pjq6PbUl127hYfeUmQYV2eP4gqssjUG0P63OmAwYsOfFdlkKFwdX3DNxpOwBlApb
2j+9wFijJRVsZw+Sd7bIEesd8A/BuTpjwp90BVAAehG6KK7WCMYTTtaTCI7CHOO1
gf3QX+9eQ5vIriUHz9MquaiREosJxHuyXOPSNxAFy3pr1nWAQSlVDFIdeDhCfxfi
RZg3yDU8GVpqMnpnvOuf4DEUmSIlFY9xRVgmxMyAvHTCwo4GgxBLojjzUUB2PMmj
MgeuJmAdx7l8ZKGFDy7LRonkacdsGLpisxWrBr6PhpISHpXQOz0aS0voi+E3pkoV
mrujKijWMhahTXdYfunaTq3+PO5zfd8jHxFPuaOUqFChTBRqxTMvZ4c9OR2GKZl4
9v5U7Hs6M5og/7FZq43XmheRVb8CiW7nkUGgzgQoHs3FiX8kpotk0Sxh6QZsBqvr
CXzO+d3K/WGsqA/+Wnzv/1DOf2vo/iVo34IrxnlfYc4+chLU0z0NUxskgtsCg8Cf
5krphu1gdIsEB9KaGHAuFYKw+gfd/U/isFt5Q58QP/TELk3xxYDnH79Bh7eEJkcW
/NDENA+VOa4sn7GHNT1O4yJKCoibqlkJd96s9YLyAvnV56KxWXXtS3uC/yB24TsB
fZl8+V1T5soOqck8Q2vsU5zy4vCo4Pg2BJEHxeYa6jrznkfX5mqcv6GOVEv+o5nq
xeu0qe5OfLvjfPwwt/JFLZiWCdQwNPybEEcAIGbLEEE4FdDZiIe2I/JQcNm09K61
nQ7xoWIOPL+Lb6ezFlfZfUCRbh3433kzlb0Rs8kFQbABI0Hb9zfhrphSnQ2pkPNW
8twP0wdkCV+cyLDPQxQCieXOFp5Guu4+eMsBOAsSY7/XXwCc9hyXd+4rAaqc/VE/
Ll5Xd3ZqXygNeua7KYFXt8+t8MHytli+zvrrhn4EZPF0aHwI9AYVxAsdpXa3+vT4
ufMlMjvWkDisM+rNXHsvgi6m+GwlY4U0flDALGy7lkO1iZCsJDQteJpqWG4ERECS
lUAAcTPhkq85waGOG92284vDoozWZds++d1r7WjY+o3W/EELNe1rCcWn5EIP0+ya
OibsgM8lwMPrm/X/rMBSIYPPfn42IC6wK1cvUJwtPv1BX8ba1p1Ilg5lZhHGGTlj
hTcDHvSLKjcdA5daU22AlNCh/TLIjx2GfnGR+zRyoVLrr7mU1XXWf+f7Apbax1VF
yW2biQ/LIGwIv1JEO7P7az1cCnhoTQM1UlRFimLlssfAG8Lp1hHpRA2TBt37KnYO
n0oPpha5DA6RFwgCcBrj3oQoCwdN+ZTevciFy+IhB+BbIyK+x59tqxeiemtgoPED
DRTdg8Xk69soX23WNb8DGVnJUg4ae8qG/LWRRj3qKXxZxWpvbrowLuH7nU3mnB0R
UAABDfs4zejaoHXHGisKhrU/7sTbeoOKDWF+onrDgl4NkDNbyuQyqRQeHyxsUM6I
3a1pY1T2KRZoW8wgHRdS7uB9RCjRjJivqblf0V+geaB7lU/KVTjcYmEBxB172tao
UxH1v+O5/ogOKP7xqSnwCp8DhOtnNmrEZX0DtQqlk99F++sHxlxc5jR+KDRCHywT
hLvZ/Ts0GU7iqqsmcmble9u3VhieNy9428n4mCu81MbaMjaZF3UWz1+J459naJUV
KSn3Z0b88AxZulRlK9nwvHuAC+FLAztT0UUb7n8qohQFkkGG/191AmXS//K8PK4Q
TVJdNrQDbwmZwO6rKbRU/nqDwFxzVA4woiVH+7r+Y9LdPfcJc9Eo72lt8jshHmd6
ko3AIu2mHp7VfcaBm47GX0Tibd56m5h9V2HLiL9ZZAWAW7AGLRmiTLKWy0X2y5B/
0HhzWOShuBqFrr22L+9AeFZDEndSduJZZWh3We/z6Zw=
`protect END_PROTECTED
