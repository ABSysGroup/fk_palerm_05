`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8tBqDKhksMIe/zYLbbUg3x4Cckjonnmh2cITq9sTNne/fe2YilpuSQmMjY/dBLqf
R3LwVwAC5Zx0jZzSqHLN6reePqFfgYdlucAj8SdvMnKIKUPQz8z4tXzH0b8mgCsR
M+qNnFXgpW5ZGtImBI8GRinR9Ufp2++DYttQO8vr6dHx72ltevUnfksceck8KGbi
TyOAVTvqjg/yG5BfvXgyWEh8NJze7qobE5RLPrU9Mb1kUGtIe5CNj26c8ue5lOlI
IbI3SwgHJtBrtOT+Z1G0f5UJq33FjD1shWKLL74STNPS4H6zG9tJOnf9SV5+vVa1
5nNo2uJSA5Qr/2Jj46F17+sLO24IJfOsYdVVohHyG1WSIktk+2MyGrGxBZeKk4Jt
IrKERT5Pf5a5rQ2FrqUQcAwc0QiQ7H8yAeANup56+tO2fNc5s6kDkbCQuUfII5ee
AsAtay6OWTgAvGB4vuHoh47oIYzwMDoe7i6MlmZ/ANj6n8U/Q46BBq6xGiua2Gwv
+K9cBlWEHcOuZ9Qk+g8Z8kGoq/qEVZ7aj5DQNcW3gu/Dag1u2q+JAkd1qXkVexFu
hXmqx+Vzdb2u1Tlbm4TTpGHAtmrWwesXXVuqfbrRiNfLfuRPaWhEHhwZVqIaIJfl
Qa7nNK6fp+3gN93f4pkFdUasprvSgcjOtnf1jERX8u96E8XxyqiSmcQNZDf6TdJT
SyilJcPG3FiuE662bIitYtTLaU/8oSGo+OZqvfszwyVKCOxpf/rBzO1ijufs3F02
qgflo7FQP4MBctKNLrNYysSByh0rEEGowNipFwrhKJVNTfH1KWIPHCv3niwGbvIF
LqFP1EDJFbtVzpa7eApA0ehP3MeDwWCrOrudxALQAEEwCpp0PU9ZjkmDa7zVZz9E
4DMC+KpnUKWjXLHTx939+SeVW/khD8elpeD4r6lwxwBVlyYqIvLXaDO62vmaviI8
S7tnT6MnDiuGqwK4FkLVq0zc6PI9V2V9wi1FZijrZzU=
`protect END_PROTECTED
