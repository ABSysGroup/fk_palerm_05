`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
30ar7OWuEbbS7rIfTyT+mys3JXK29Lt70kTFDQVKfDHRScJO4yRxttE5J3lgBMhd
0y2ZaBdeUrDsljTiys2uOJDYKmoOSJVBNrm0qIRf6753GSAaDGav2MQ5LMZ5Ncwj
KwEmpvjpdUTfGlAcBmn4AoFUmefUVnVGVzCAL9+wV48gXzrBphZqUAz5hRlXbWfO
OAB3HIbFUMzdGowbfOmLE36344NHcUJt9aycoQfiJdIJQsPhvuFJmlOGNTnLtier
DnVyabQNSAN0IajwMbd6JMhFatUpXcm46CirwMnHqHwSDvFkJQ1zzKkdMVOleM6m
t1kFGIMeo4+XMoq9Xun1dHSJR3725bCqIDTMx0Zm4Ibx3vJJoFoAEzGIXuTLSe+0
CFW7AVunnLRgBy7+0lsbTHNjDaPWdll2yf65U/idp3E0zYTFbgx+xLRtHzR7cYgR
b3a6fao6vrJ+PzR3m17hvha1uWCVcpGKIBbr07BelFkFE8FrFiIRVtDL2U49c01q
5YLGSj55FCatCr7bGqTpKQDCiRq0kIo7LyXxtqyGAIjCNWjc5XA+FZfcxAXU590X
f3mGbXNnmdS8UdBB4H258aKBpP9rAkJes8ZnqA4H1d0jpxPXpv0oMmgwBWkGM74m
9bH6Gisf7I3/xqsfve7uRYvg1HHNxKudVnhbSBGseJ1I+HmEiFA0pR0Pchgq770F
lSsodwIMnHsSa0z3FJ7oHlkS5WYs56ZBMDCoiSaRSCSXyDk54Zfu99KSZTFk03oP
kdf6kE0yJ8jQA/OqOn6Z3TOXt9lmMSpivfbhGOXXmeHQeCl9TaMwZFFWxyQjFYih
aqQsyBp8KrOyWkHdx0q0jg==
`protect END_PROTECTED
