`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xlLn5LyUHeurfYO09WFlJvUXTJD2Y/XN3FkFKPTGCtgSZDk4KX8tTJfeeygPE51W
pk4KNjr1mLStejD8RZ1PAVI5yQG9pKKSWtkGGICwGWGEIA2z5/Sqyr1WraDfn6uT
8px4A6yarpn6ph+Y18eTxxVZvm9ZanL+kizaLKNrthZM7IW+m6A97nUw5Yo6XGKV
pGCWHoQ5hfQdGNoOOdqXigRNMNQC5OUqVtSBe/ttXH0vtut1kBKXnAsbIC6um+py
cvQ5vV0qmK5WzKGYgkr6JJIXAI4Ntq1BnDOzb00QEz/nL+YuixYdb9WfavUmdie5
dP1SAC82yFk0nlgbDzYSJA==
`protect END_PROTECTED
