`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mU0aSlhs6+AJs9Y/WiOrN4NiifuF5QWWoeM/J9tTPcRpcDkLGucY1+s+P+6UGppc
iyDEF1DRFB7KJhZzrDkHPRy60kx1M9OAhF7XcssI8WyP6X9ppsOpTThvy82fGiLl
HkQP08gfqZkKOqZk2ocNha3IJqtJqq59VdPF3F7flkhQuThn/vq8bIV9vuTXN8W8
PDJCe68u3Qj5EiGak8vxvHplO3OhS7iUBPMRWzFRzqBxtfUhauOnlYzl31R4NK4I
HzS3DiqDGKWTQUFSI+haEMvTkZmYWxo7iv+PbcVyudPacCmMuLWXVt2FkePP/hdz
s40MURWtXj7df8OM5PTQha7TCaSFHA4o3nm2HFuZHwPvpjcZKOWjBA6KdKPgQxUD
3nzMV6oiZhzbvyOyC2iYMKo708AXKKFCf6McShJU4MnIPklIDmW8JIjp+vXR1vwS
4ZYKggL6ChAzhlQ+WFepFs/iZRLHRZGQ9oJ1CBQx3s8CG0c8Br0vyAcKeJAkXwM9
TOR1cY6ZgeFyBOxTfKFhRSro0lC3u7sb+2OSH76s9XP+kbiEZC1yKUubTcERtsyp
Jjg3MJodvtYXrXasjBxuyKzZ2BPh+BI3AesVdgUcB9luSMN/MK9E4TsaLe4F3qdO
YiUSW2p+luY9mYBy7NeLZvOOK4EBe9F+o5J2NX+K3Gm/wr3MdiD2qlTZwNGk/FjJ
JCm2UhCXZyav97hVpeXoL14G+iO6xCs0nI/jhOZpaypkiYEDgmjBexqB72sA3V8I
pwRr8hwKEwpKBD5x3GBDkA+B5voYnXsM8jlp+SMYrUR9ChkwIU3kUs4OylTQWcj4
4PIZBUN2dHUwAlYcWXsCA3Z26OVWlELR+zmNWd+BevCtKmxkQrMvKtUiNjjq5lko
JMBlP52DJeH5dPcLKCZTdS5Lz7nQKddD0wcKwTSTzXSArsaBHgi1WeaPx4M4ODff
D+QM+NJtOurti6E92Vl7c3E6rMYr7G0wgm440Fgajexnq2Z0zO4o8P9wBJGJTX/u
+TgRuDtH0jtV2RyDik6RzE1Z7ryQLnhxBPzy5A/tVfuSt6HeFUuwAdwwBy+4Wx1Y
tIu6GzvWjdskrQ75bdwpsUd0/LpXmqkBRYL7VcVFkeO2/oFHWpBGuzfFjIfZz6IJ
QjPHmVcW1+yJb2ySB7sXkHPZPtFdNwZcXc5qTfolKC/Pu8l2nlrsk/PIsqy0qRxR
p2eMe0dExlAFUivtU/xHLK2kOSSvA4JyOmEFs/CUYChO+IKtAsBaALred8TbRKwx
XdGBLMjJiTtIpP+ahDld2oXxZA1FfhoS3Gny7hFH8uOPIz7n3/AFYNtOB6IOlZfL
pKC8uBcl7do7t8imM27aTPYMwky2kajASPcSpZrz2I60tM3SpVo9JqjHKwdqTWv7
X3e18SrG8+DEu/bsrUP0bKSmERmwKjf4iLaobUg8Yb/KbO3HHppFzzDKb5aiApnC
lxccDaE6op24AfYBU7ldtAJTW7ItzY1ncG7l6ENNYoZAqhoG5kYRyg7xbb4VcwSH
qwzys59oOwq8xCpjbLeI/01jjYPpXBaol+omEvhOEEKBlH7qBZfJ/2o8thkRGQl0
ES0XX1tPP16xZiulQHkPlSV0xRQM0lgbs9hLJ923+RfJwtpKSisko3TlVjIhvLsi
xRMzlHYOX6qOWP+ZxG3ny3h+CV3EnBCwvHjGhqxh2gabWGpSziftTp6LCp1Noqqz
Pu6f2w4OnEkAJBlQQG0/Bop0SXfLwVrTevUhKwvuUaPaWZ+Wv3y++l50pg/qTQGq
frq2eY+j/b8hiazLFTbS6PIT1SwXIj1hU7orpY3QO/yFa4XUlmRXN3MbQs+U4yxT
wp4eN3sLdDT/TQzt447aFyjJQnDmdG+o9qLKJthvjmWW/BOXY/ZKnt7yusHntArM
pk3uKDMdf8Qmol5LYN98WYypYGwy6mEBAaOXTTKvMNBbMAWjOwoX4mLiTGlgTSFm
VCDgtPtezWyeUDctjwYzN4EO0zU47QB5dUpJOKcx1t5IQOMU0pmS6nbnaLXPIs7Y
aB9x4N72ZQjACi6xNLszI/7XLROIt3mcaNxbCHEad4yYLTx9mMlQ93c3jBeg3FX6
kj7SIPNzd4Y9k73gtv5P0iqO5O5fmLci1eW3cFC/F3/IwrOXc40azmH01qobZyWC
6NV3dvaiCM9x4O2oxqd3vt3UvhKSdByQoy6X2q0Vx2D/iLHCk04q/cHxDYlKUc5I
oyybX1q89SPbziBKs38soB7vrNEr3OufmtxVbqqaHpikkTf9mxLzxfyMxVswDNs6
mhxEoDPbOhnq6fVBssXzCjFXyKC/+krh4DFBx/reIqz2fpO8g1uJaNp4RKB9lSid
yJN1DCEcg9W99WC5roQQLVYY4NyP4rVXo7tjp97jo0rjgA2JZUVRjR5oRJT0ENDP
3cWyekZUaVgPqJlXOVSK9adXikVevTqNJlHNKVlAqf0tZg2qEJnQuubZ1YWwATSv
n44HQchZKldzSR4R/GRZXJjmjpABcU9iKHO/isVrgV/OahJXBIdKlNxVI1EludMH
Ki4d56tC0f1xSIBo/liyutUD1GDe7tDHQngJ5cA67oFrd/9wFLbLcBxVTnzIM+pl
s69MbUTJ1nNykuIHyp01Eo1v889MT094Gmd5sxnI/FZduREeQ4NtXzyfag5CU/rD
weqwp58oz4HnNAlw5VfoQMpCVqGSvxkfZNYPSThZFXwJ1GgyOT292y6hQN4r5Hcc
ryrs6QPjb4q7UPXl2+7yk8Ux0wLHod1s260HEmDZS+5N9cIxzF1Y107CHWmqOpnz
X3rZwvXxNprdvx9nakuil4rpkJVqsNnnImk0mVdsii/LyaTM7Q9P16rk4umqiMi5
6svmsnN8oWas20D5FDSFND+vt5iRegUsO3Tt8S1hDgfUpKaMmMmcbcEeuzEAjtma
SV9n995hpbhQzcONdNLyfQJoPh+fPagEi6QOuUztIAvVST3dR8/iA547KreuaMOe
96mJytAwKgjHXkJDLiHMLTWc2FgA+3nnifABRQD/YwwzTmyS6nyVddyglcClDFr9
Yf8UhyGpFZRGKVV4uc9IRk6Ud5yfYyJaDmum6BzAi97v36Cnc6IokH/zX/68+7gV
nPhYqfec2ucYFufywWgMp0+F9W07J5tRivmmXekd9esRiI0Bozj8sT7cn58Uqwz7
tMm3uPQXpJQveXVGmRhmU0ZtTdU1v+63IUn+TnZUhxGHeFx7a70bs0TuuNFV9OYq
+4UdqCcKUGNQDPrOf+mi7LHkmlHMLDLCryzPITM3mz2JBr7qUBgj4yfSszTl82Bt
Qwp1FcrOrqyOKSL/SnqcQGeXeKLpysf06LChmAPeKF8=
`protect END_PROTECTED
