`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sJ4lGhaMx0wsh+tatkZPX2ulHrfqd8xyU9fFdSJFFv1AeXyFgy/uKMC58tY6E+No
sumJXmzeEKrk27ZN5s3p3dw38kNikqg6mmEKRqM8GJ3S97wjW4Ea4XBtl1E1lWS8
d8LRAPc40FWLY5xHmYNrtNETdCVIZ977xxHUfnv4jOy2i0OnrnXjMpbdos0V8HUg
PIqp+SOK/wSSgdrSxA8Z7CknRbHjgjIRAw3pqdqxbpsSFaYNWdj3ZimBhHIzQE/+
gbv/Y2NCpLdJcNrzCFR1fA==
`protect END_PROTECTED
