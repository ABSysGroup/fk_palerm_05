`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uEhV/KwTb/jh+/+TQfSlViZz+GNd51XLXpQauqnqwpKUL81iCtOl4XUHGY4OwLGi
VIEHLX/u5L7oyyE8SeS/wJOTq3mNspwLlsGwFrtWLsz9c5jBiSsLBnuioimIvOGY
Kcnwz8jxgEPIPm1B18185SR8sflNVR7ho7m4/YuLpVYLbXoGUP0vkwIWmdSQXIRX
gb0IAsKbh8Qv3+QR39aiJB3xQE01hJiHmJpTxASWhdm5xvtO/BCyHyo4++Zz9Zy3
c3t3AbqfYDMAwJWzhk4Pa2tZcnGM+tFFZCN0TLQ4Du6nA6at29gQ3PCiezV39KPG
mfvP5gYxC2XGiJEMsC7V2jNcK9+PhjqX8IdnQbQ9SWsoD1SexgTTavf4Mty5Kdx1
f1XCLAs8/eP5eiBpKWWMu2nhYrt3utzFmYLbCxJ5mogyb1Ag5cH2LUs8s5XiVVtJ
/0jBHuzI9+Ty3ztDWC+rGdnOOyUVnlDGaVR9FrJB5vySp0aY8QlB1M5dwbv0YnyA
rYLByOgUY4EgvBWovucv06CYzb55L8yOUys4OEYTI7+gW/VJThZGU4vdiY+iMstX
ba1lGQIK9xtRGkBIWtvdfpDv8G7w9W1zm6oEncePsU0tFoz/UC8LCqa84xJ5EeYR
qjF8GrKCVZo/YDOPw7p1FHHxErnJWUrDtxmQjG2zoRE=
`protect END_PROTECTED
