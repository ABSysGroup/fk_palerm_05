`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PRMTfFWvNXrWjFsMolqs+cEc6b3Ci8NXPkmizdewXwignL7zsSkKto7OMWllva0G
HoNMrwsPvC4Dr8M0jn4EX0b1tnUa9HuOBkgkTEevE+nR/cRvE5iv/uaPMKFV38m5
P146uzlNyQcqh9I/Uszwsrp/GtcUtsj8ertophpZQaClUYBE7flEYAYyqa6T7S4T
GrNKYNL6lfESMwgnEMlX0K55+8Nmxbux+iwM13tyIv74vtoaX8v4YvxZzQyY2zLE
x66hrKY/5omPLhXw30u09MrDMqOs9AJqJG2b0pMeqhkzUnaQb6PnoVyVv+PmYdhH
SZF6tqNzJTAiqbWSqoS9psvn/VL05oNyYTp8lexqWEvXlj3vqQWSxMoEr5K2jxiX
d4qlMKa24YxYyYaHX6th+49Lv2wSFYIP5JPITc/bJbwLwbp4XYZ0jzZMhuuKGx9D
VTMOxh0azqJ8ucvoV8HcSEWCZeQ1wxZHgKJSCDb0ONU27EMbJuGVh1VHllxieTFq
haBvxWa7TmSKyRNAzm9bTTIKtUnhq0VO8sgAylOMiG687mLxJ+kYJ4i/367fZvsE
SmdBSQ33C2WFezCEfejppufB1JSKhgG5vUaEJNpgEy+N2Fhb7lLFgNF0yXSRb1E8
`protect END_PROTECTED
