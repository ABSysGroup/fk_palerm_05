`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TsePXNbm5rjCbv7EEvNvL3mk7P0o0OCiJ0OYvuuBrl/P2dL0l8gmifcJu6JBja0b
59vSxK13ZzJVoFKBnftkAJ3uHRp6rLOBTVzpBf00OHb8A0KR5BNWMFckZ+6jgwyM
XrILKIbFbXedwcOQX1funKtoXcD5L5+mz/OM+SjxXQQC70oWvOnbMm4meCg7/wii
6CmLle/nENkk3f2AfVztffKnkeyhtkh13RHPsdrKKHSSPbfb6P2A1GNurMUodUT5
YW7lNK75TvzTBysWNLahxlKJeHefxrMmXXcaOx3EUUoJB9OETU3mR8miFZgHZLeD
OHx/u/0t+0xC/1gOVs+muoNcqPh3i5i8n+jS+R/+6Ry2JkRbMwZejJA3DZD8Jme8
tvVFauJCvLKoWUDtZf4NSjRUQK+uxx53TKQmk1NMDvOSPLaMMWV7ALnj212uPT5Q
V4r3MNc9W1C9y4mLsEx0enYPVMKRgnFBQ+VE/GFj3I4YV8M0iwsT1pDQVSPPyBUa
7ZxrO0rmZzu1CMFngp2qa+pKxj4qKYHSJDsVrYvQ8gzhd2BuGzoJ1mgI6iDCGNoR
3sSfbzRKqu29XTnwQ8CT5lwuclhCdxfr5a/HMQbEk4Z/kH30PQmEmna+NgI5QJhg
qNsANhEt+EMNPDQNLyz1L7GN9LtbtdW9F+A8zmGBahgkia/sL8+JIxkeBaX0BOlH
9hp2/WegZDXJ4g7W1kDux/XNC84jIWnkCPnCJa6SzLhOd+XZx9H+F1ekby78JzYU
QkVtjSl4GlmCrqWwbCOtanEVjyp56woN8EX3DyC8PaPEFIGM2jbhfhjTKlGU9EaQ
d5HFcE3AD/Yh48ETsMVGe0oBwrfVp96WLpjzYFjbOUi+zvzKA+6LNnzWyOqj5BZ0
tnJIEyIErm4UPwZqVHQCS8BbwiScS44jmdeaQ/zPuVGzQhqvPdVJDgEVljn8iNRJ
JTFBj9KxsuSKHMpw3yHMtxJLlvdwzqOwUNIffKg8uqvIhYkd4WKzve/+KF0n7KKi
Pm/LePHI0hqsjYhBadhMCmE4YhQeUKURy8MfdukLYMQjkNpkDzWy77OUss7Bd5nn
L52jKevR1xlrBY9LPFjV2ybPJJDngh8XSM86LHlu7aXo082F6Q32Gj1g2S4wpB3s
l9C0gbE7/qrt74kfhfgu8n6iwpYYY9nSVdZE3DTFolc9WP0LwgWGr9+ZrF1kcKjB
W1zlWP6AQ+H3wVAK/wAN+aWlJhBT0iA0lvcFC1TuU3NAD9aMSCb21N//LKrZuZAa
qvPCiZHOfoDxwWct+YfM1Bw2JAavIc+TzR3BO6lr9QMFbpwMP+kcGEdkNnsxIzpq
z0vi/V/Gk/WZU32lBNghYFy4gsNVV6mFK54uz+8TLZM6dSFSc0Tdvq+q/LHkupXj
4GF/LJURN1Zu5ZCbMWDu9+O9olOwo2EulVKi/6EM5kSW2LEmjcTNbFAhj0xrqZJD
7MVMOl4BfcupNuYnX8eEupRsXJ9o975xgziqqUGitcg+lpW5j7/30IrwYvc2M3QC
jKSeeVt9EHkAKmINYI2H/kX8n37PYNfuF/nG64xrGzmqusmjYKYMqoNLjqk3rG+5
3o/oCfWcFVZR1+EuqK5wRRVBq07Sjt3VmhDLTh+P3EebPF+jULI4GBgfUjxblc41
dGzYQkgBqwUpU7z4orVvQkfWR+huucfo4EpHE5EyYESzAxrC7ehr/sbUYeKkNrJM
Be+lqFgTi7eJSPCazGN4ROrIzsbKTS+5r3E+NyjDaSABDhpkqggPGDrnZOv1cOIw
ryO7v68xIyF61JEDqZuNfmRo8gQukW5g5AX/ynZYaXmCE41fLShaou8IgZm9lZtF
iUhCQudOow9GUKYuCAeZha4VZ2AsLwAK2rLkFz+PdizjW3nKl5I9fRkEknhWyd1S
e8npBVjq8wy7h6kjHrFjbO1YBHYvYRBQJL5D2ZuOyIWiGPAnUq4PZCrWRUF4eWye
A4zr4Q7d2hwKzDsnzKDQdJSMOT1FTKx6XYIAS7dRgEhDBuXDwcRS+tZ85eg4TjTO
W1Qf/Aa1n/8bGKSt0XAUF2sySjJbw8JjKBYfW1DJSooynbkm9WtMUImrUTWQ//T7
ZtN2NJ2ZImilMzbnZuMIzBqTo42fWS/sajIn8j55EZYSbhVu++mPsgqHZxMQFKQN
w4MIRb3SOEduJeMcNHfKs92ZrdEVO5PD95uioBYYnGx4+s1r56unNNh2mQ75C9AX
oWeh/J3jZXHw6cU1P8LjGmk0G+qwH1f83TF33bAcP7kayIs0sd3/YWcOAR72EwSV
s4M9rij3M9AnZFw/0YMJAIGd75dx03IrFKXKZf+AdODmX6zNoviyH3Na2Pr9tI1Y
apb0NgI+02lchKs42+2gRbUFXWh+c79bsG0vgUpNGwJsC+2tK01iLkLcr4wRVKPN
jrn5hFFaHdqw8g5TClO1pS1kcoQFesXJSD4vM9G4O8WCWN5zXXy/Yd5UkUFbK+cp
jy9zM9Xew55EKy/WGOtH6uDNzwmIHpaGKpOgnS5rrH/BXWxXh06OOtOh/V12kvLj
jysRbySZ9fOxyXxo7pnX0f6ZfBx9I0udvjNgoIgIBh/2TKZqtnNkG9i92yNb9cTM
CkQs3XngISW4ujlog+nPS48cTMoQSbIF/uXKo7il9+kTlWZMZfTmy22Hf4Jy3QCn
T7ZKKs/vaOybX9k+QV73+JgV/i5xTsEU73On21Y4ZeDsJyWzAtxdykw0pS6HXFe6
PifsFi9Gko9b+I304ue7To9/eOwtfslzlzjefi7JmmzMCy85TVP5PAM7SVVv0Po2
gLUEfSxUeL6rLkaZPfxQI067SwJLLfMi3TdmjI7TEVQG/F5rueSSVg52dcj/tXxA
zMGUDxJ2mhZ5diyociuJGrb7Q/5WFrcLNOnvw6AiN9UD63491JdmUsVlG0+qIaga
DRyNuz9TtdoFX8mvDKvlYnnWd84H4O/nWz4Umwzlyit9wPlJTnbJ6RPg/uoWfEhb
Ei7h1bC6ee+nSqbkSpQx5DE11j+D7bElJ+iooVYCY17rDCY6KiMMkGKuPsxf7wxg
yu9o63V+fTFkkwK7Vtz1NhSgVLxFBiq1bf2wSJMLuhoCkjpKXsBZzblw/wIfy8wF
7cCEYdkpPMmMqahLTcUTOhx9jFRZJqmXxr8SQtm9gEYhTh4a7TgDsHqokeTVatyN
4yYd3EX2RWb8Dr8iR3wHhELIaLLL4vYYOXLZQmxUgR7T9X5mju+fa7YMkyjeEB6Y
3lqYjjGXlMT7ECc2JmX3rJ1oyo4Y8hOeLxzCSCPX4pZs1yxl5iKtdWt7RjTXJj3b
ZOXLDLXtP83NR2H5IEaqb3isO5IRvQwKNJaMdGRXVNXEVHcZ3lGTPPOYis3leBxF
DLpfhuYImpMGwZdTSVUekSXG7rpQpo7XyfY16TtsWFskXsvK0nYwm6ItCbGJijkG
+1qwO1UxdqBUQ9YA5cbBYNFW7Pec23JmT7g0jp/Hs2RFT+6JnHrhKiwQp7ag58vq
sZOiZgLn1C8vfQIlRtNZu4t1O/eqfXqF9mRdPyPN53JXbh/UQzCzI0aUyV1O0FEB
c53onJIDowKaj27GG3sv5aKgeQLm4ild8uFIt1OcabaXSvoOoAcgbI/FhfTxDMIX
aU2v0J7efLO0UuU9JjjmyXKwtrsDaSKa9uHeH4dBie9EJLWE1blB1oBYQmEbpGbk
n9je9/eKnElLqEOV6ZMcC5ruD1uScc5DN6imyUvnYQMFuaM45MY/fAKEZieRI/aM
vez/hIXTNDa1js3LNBwCfd45fducyWPlQo3RoVKJY/P8tcXSW23iTFl06hnVGiFd
GNLiENxG1Z1HAypqg7UNbjpihxH7Eo64psjP60AzNwEJSrgoSK6/ckzz+j51IwzL
IOZIsqtlcYFpObOJ3lyh8FQ1fsqhVITL5mxOCumt1gh0NMp7GE9EcE30+1xqq7TJ
HkWwvLbc0JItbGCUatU39+J+IBS0HqIlHwsd2bvXClhUo1HvyZFsFQJOJnhMqHmu
xPrip2VnwdnVaNE6OFRMBYEGNpVlk1dGwA8/szwfaTvNBVZUvt7pEi6/2Du6E6So
H2CKGGtdvsUTOyQuinP4W92dQSVKKSX/tnRYE8NnbRzOmLWJTxWgHP5sX+38ZlL2
JHb+THcW2Iq2uRgGPYqgN04VnvYPDfueuJFEA2v1H9SFXAIHP5eJRyMcA5d3NTZB
98a3msUbZn+sUKjws8fh672O9Ny/u/ZasjheN/5OK8Zu4TVvXeHgMH/GYqGBSqUT
nyEwK7yrXvd4JJxW3NQEva6A2RE7JrxhgTmJDg14K0Zyt8mxaVBknEFAWmfjD/uJ
Eyx/uop0R9D9OKdeSiUxL+/5zTp6XJ/T4VEcRmXWHNCHhrxHKIvqevSCDC2rJEFU
p1oScRMpbvyUGuA589SZndRXhFal51wPlnoBK2or3wKRkBt74EfL1HnE/QXoIRSq
M2btfOh5Oox014GWA7btxBQo1qoo7ZB8MTe82QlQz6pezqeHMkWelS9Yhde3ms/O
d6VawDwGLKfOYgwO6PMRtgtYVDhTxIrupM97ydMHQxAupITpcVU6fdMoDG42gdHm
8WZovz0+4TLARR6WsIE1mee23URvjcEM8/gR/TCgX09JtzLqGAXppI2WRAXkgMFA
a3D9MeOkHnH5viyuO9nz1DntdKt/EuqOPvRwPnhebOni8to5uPOecH5euG9YYoX7
iBcMnkZOmL6E5ruWZicn89dnF8+qaRPcNKppKwDuiI3srFwVSACCUQ+ZoCZMdpz+
yJMtxOOYrEmFtl45Ny3vIWpCe8aeX/gZTe4A4opWclhHBItjT855CUkCjlR5Bw8h
Mho3MQH0Y1jQ20nmh4OwOj+frJtAJSuZ28rGXSNanrLhrnHGPK6HGeojf22ahuD2
LJXRTnIyN7cv22NeTFciNN52yBQw8ybIcq/t5kCqUKdQ1y5T/BaXhl5HGe7DYtJA
kbmufGaLAqN8tepkXjr4ZfbVVpG0CfCumpkSrVZbRMFNtX9HswbmwD4LboPTRmpI
sMUhgwURa60JlSgY4j1MiAoiEjV83O5xBb1jTXMN49YrHzjWJ+Se9af2v5zH3bKl
OJ9Vip5JTioRUrK7HpfbY09F3wY1Z7Cvc9a1E0QSN/rgzSQASUNwkiJwQBnQ0040
DNAFzaerASaF5ytgpULrXmOxRacUh6zCr2l8X/fDI7T72LS9wA+mqhjciFXwFLve
T5UE2Kki6+U4ZPEmGxgnhKCNezY8RCozl3UcF9o3QDS05+Pb2BxDl+IZHJuwRbAE
5um8s0TPS41Lr/ycLjZrNDLJTwQrqvtSzlXBNZbSPY/KFLBB/M3tShlq+caeFIEB
/F/t+cu9LI6f5B7wgSsWbDt016oejtVfmxoEU23EEtjQg+8B7cQuX87eGd9A4l8L
sY1PSmgGNTipO3dpwy2/pTpleynubFZS6Cir6dCaOYjYFsOKJ+3V2psl2vuu//sg
NgsxAINuQ44TwfLAvXbVTlm+jP+O6etWPKWP4Xkbj3MSMt+0Bv4d8zp/vSPoXKSM
0VfidG/+As5GkjkhieSytl0b4uIbUiAD8RSvOlL3nmni1+8uRMZiNywTfoSqECMs
kC/2FBut9rd+pdueMgdDATbBK+BQlYSganWpogCcawf1+RXoaPoEKOa0WIq5IDNL
z9RBHGKvwgLgx7cqg9Lc434/9IxBl7LS3jopp3YUSV9/lKMntJ8EALIsp/BOwu8T
7rwk14s2ZmsN9HIov5Vr5Tl5dKv9BXuDWqSNkiLK0YX/6RC+DehjZK2HFQRVWbLE
h5hGrW25aEtVjT4yGl249lKFLY1EIF2tPKiZVbxIe+pZ5KKTvbfTY14pfNqBGlgQ
GM6dF6hcQwVPuSbyaUpKKS4YRMQ7bNz/pdZC09ca3h72SscHL67T1HnSzGYBxYkw
EP+CQLE26eAj1LJhGB3lgJ5bKDaodP7MdF0ouK9LBr/EDJ/kilJRZymy83Jbdtpb
X4afpwPGrrTOsWdCjsenuqgDh4ZW8ADYbY16VFjoqP0U0DDTKcSSp7xr1XEdXfS0
OD1myVpRJz0Tj4Cw+W3Wm/kw1ROU8HBifToYc5UkuIJeAF4jLpp+pa0+OpkovIA4
HHEmLiQbXtg7UAV/zd7kXVCHT6iAxYGzPHDueIra7wwBLItoy0HMTFKRwECeWeZI
GVNpicZDoyI0yWiWy+Cmk0gDDCBGTiP0wwc0ft1XlHaJNk4RqI1UCoQoE6lDApAO
mTa8WIxR0+rxPHwwO3M9Bczjeu2zPJIc3a8oc85ArAXsaiOlqx9M02xqtC3YLokY
FiqBmh9pF/Q9OKYYkWHM4BtFZ1zdNIxn+UK5YltOLLUoWMeYIqTaDEK++nyju0ow
Fd8v9gqiFYhyLmB+XJElOAy1MWbZqjBfyz7ox1ibtTUvJy/yMbRyBetUHVxsB4sM
T7IBj3TXJfdtZ8TdOP0Rf7wHzZrvpd4HtP6Sho3qHvQyUOY/XAxXwhl1k/AOepWz
ehgD1TYx46levDnIJgJnZFScKg3+9JFFCeegISwpLNdOjU9/1i++PshrOGBYlQT5
q2cSB/qG6YwYVH2G86RWKbWgDGFWpc6khDJMd2mZDa/HFBkN1JtJrAuJYpCIjIaU
sdC+r3/YZfvpOV789wf2rfhg5aT8s4kWz26+76h8HDLowQ32pz0PywQHlVz+F2k6
FHwJKp4kJosh9BT6TRiSOhnU2HuQpLr91U7CGyWtDofyJC00LI7cMqpuS9d3qa49
JIxCvk4kb/DP5azceCCPnf1lSmWVU7n3TuQ3ef5UZwTP00byNxDUXQq/ihyJNO9U
1x1ylqr//4mn1yf59n3RmRd1PUeQdb5Sma35ySYWPotFPWp8y/Yys2llBw2Gkwq/
QKQSuSac3NKqMf0LtsBB+d1kft7Q6xmhO3WHHqogOYUWc1D9dtoRSKVQ0HPulEJf
bazCojlAxptJ3rV3zzbHFEEiUxVGgEDTdR+wkqWkJmkBYGHPTYhP6fdh/n0I/tN1
ggn/V9qbpQZ+EfA2L1gocO3uPvVMATo+FrcUEwwukTCaX5JPfhB/A1Pp7WSrsgfZ
JAIIK9OJMO7yFUGPvvkmwjv7yLspOj8KGuWrdVdSzB8oLgTvnOevCVmCjCrDVj4B
bpX+fRbWIpo8ULFieQHpE4mgy8E6T/8NX0cvfCu8C4Oq0vpvBR2B8rU2Q5lvAp7t
OkxOPaKuvoOvQUSVllHpK5P7M0NzFSqQ2Bo2hxm4yRYS9uI6G+ek2aXyzPQQtUY/
vXCMJ+HTPAo0yxupiBDBNzg2XKvTjBynSCJcpS7cFlofpsyDy//fhKfYzuiagw63
ZiCjo+YkelFc3Kh/CCcyiD6h6fykccoOSZAsyg8Ah9AU7voVrtDId5Dyl9Ifdlbt
rtuhv1dBl70dWbE30IKDbUoH5Bb8ii67/ojVS8yetdTR7yapY1et5gD8V7nfSZuB
Ime/uE++F1V+rYWHaXAJHQtDpG55Tau80HQMXXjIzjmT4mkFdCtMf6UePmQbG8Rm
lGQWq+O72Wf/KdznXDfVAQ3oTqdQ6vWyFOLjWJsbewXIBxPvWiWOfnAKyyB82Vfl
lGLBY7GwlfBoXl0S0FmFxnBZz16HtSbcodo8gOiuX61Q5kntmNTlkDmOpbHS3clm
smSGl3tEzZEmS2Nr3St+NisncAqaRdBkiWLDwoPxLUHkA3qKqaNl8N7gDOn9cBIK
aVTDt9pe9SuYUI8f/lu877KQZZK6r63/nhS/1AnpaNT/XiI7Pv0ULdfHfhgxTuja
2r8VyquFpSgxHCGh886AUXDK2Z4UfGuerFz3wNt8fFmQ6McI2BPTGrwFZHxkz2yS
L3npJxc/t/myw66WDb8Yh6lk+fyYx9KSim4zCRbcm7zaB8xGLv3B8A4q5lpNwwKh
5z5vCNsT+AKPO6zyRFFrc24Spo0fNFuZ6bAGwMDwI15g0Gn81W9heM1nJOeUrXhC
XtZrlv4pSoyNHiDYZ/1u6Ymow51Vbk3u2hB4HSrrV5WmGavLi2IWdJwJSdvbJMWh
gCj+32WyxsNzQ5FD0xgCIesFcPfRzNnsabe5i6pumWFyBQ5Z3D0bzSEYZQ05Z/UO
9Asz3eWAuyLDR+jHgP/LgwB7PsZLHRcmiw3vjVZJ1coPxuxTN2MmJRwMN98TuORe
S1W6NOg3IliJQbsySzzRsBYtk+PHCgUzPQizIGLIfD6CAWJDGlOw/BtedkYw7cfQ
FcQyCMkJRC6myygsmk+vYb+J3cpu5qigCF3jNrkFEz1idngEaH0Hr1YksNi7hXwd
R6C7DuGMZBMbnWZ213u2HCZfLNlv2MDr+kOVDOFlwKhG0Ta4+saAGKCp3amq3A79
4+7k/iBL/t6yYZfGwlRLVTqgTFFaBd38acEk30xhIHcj2a12Qk979lOemedZ0SFE
i18B1yXcF3biU3lG5bzKiq4yRQuS6PqL0GNE7TyaiCGcwM3nJkypfeS9F2BRDToE
vaLWqHJOlMDPU9ICnaOBpJC5yScuc/niSlnevFbqC8hGVc5a0XHG9AWSL5rZSO5E
5NITTAkZ2S3yL7bnkch0rVI4rdhgvHEjgTB9tfrmk+mwX6R/+8TLJeZtK3AHY6v0
1jRRezQuYOWc8RqZI11N+rgADh3LNZEpNRbYGcIcjf2QVwjqVqcVJNQeGczeF8Tg
naGfegm2tGBX4hDHrZMMX9RdEVGzqhYI/HYzZePtUmt2mroz/VZ9J3+FZU5805D0
6dy9Cpkc7k4uyllGMb50bV3z5rAj+VzTpY57YB3PzOEdQ1HPpPXEEz839koOi6x1
PM493Fa5BnBwOFoaFz/oDSZMHp2FUScoEE3Q+myr/hTFDt8ul8w8D2NCGf7ZHlp7
KYmpeqBsX8XmDs+6yiUiotLhZoa2jKmu1vwH1XxyRUX+bgbBL38SSUnTk9Xkg5kz
eNDAcw6hELeVwbAiI+LzJuM/rPu+WwtUnrdKT/TyzdHEWz8VXZrn7y8/kmj9+ybA
pRj4Yz3PNr/Wnh2fURVewQrHzR4IrI5eAco2rMhiTaSPeOBynTrxlSCLYS7pxYZX
S1WaBH0FBfjqJqVtunj8q6HZ8C/HeStxLy2Z6Dri1vUACiRAEjgW/gKYkiJjWBkR
DJam+yya8DCxYuezvnZ8D8lEJHtbPe9GPPPb0jfn1vrcR+gzGQjapOTYw8Gv6N5g
LkT8jDC2GlCDNPvwJoYybaAtaXqFG8BQbnPDbEAi8Pnxul6ZhKp6lYEppyKXlD+x
fgPmgFbad6hqN02PffoFUMQcjhgPU5Hwuxdyp6mwdheUpnhknv3cWrEnzSmAQ9a4
8HiW552PnAk6IuHNTCTGnNF20Dl4SPAWzDY67rtvGlg=
`protect END_PROTECTED
