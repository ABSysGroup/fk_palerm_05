`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t3OFY9IyncAUHw/BIxTa3Lc0Bm+I3VNWsGRiA0UggCLsc2pWK9WSVKhE9cZv+lcX
CpYUGI/pBvGiZdPYCNEk4q81uEAug/dk5qpuqokDySt9zAgzTjhUjCCsyKqluggE
740WKFL46Jc93w/rEVZ/btZyXncVEaBf/84SOayKGymI9W+ju54KK6FHHq77v0pi
B5ji93FpV+hDSazVKb5EoPoSHyKY7P2iKkfEmUwmqUmBT6cRxQZ4tMAOcCfng1a4
Y9d1/+HLbFFgsJY1vb+p4PC6sjsCEN8Tt8b9dCktaNysKJGijdl1ASKM6KCoYV+g
llzoUA30FqtYFAzJEQOZtJtESLQbSH7EH95PovF10TgHRS1kBQS6FAp3gCMMq0Jc
88g9S1fzgfwLM+rwcWK1zxhApQCItP4XEmpx2HFpZ/V5ZnQRUgsuDG9Lxx1ZsmDj
`protect END_PROTECTED
