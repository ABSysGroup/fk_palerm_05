`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XxMdn1kpypAhm8Uh9AZE9MnjC3Y2HXzw1L2GrbF+CknTKUvhJUys68D2VcK5m+iS
t0Z5IhBvsBIRd7z+qDLnNzwz92eUG5p6FJo8NqF24fhYB6aIwB1QlwFKeaaBx1d7
CaQqHmYk3YmAMDgi/b8gZEuJBrTZFYsBeF2+XjpZdWJunl+rLRuT2LqpbMszIA8N
eRFcclxERGPy7SUL+WFWN1alLS5jf8eNhpRWgMUfCIx6kSkciHWnFEyza3Bd8cAn
nHOClzsF4lM07iOrEiL3uKZpI2hHn30t4vRMj9xuOWvEE6c4871zqFeTEU3Qrozt
gr1QMaQQZzTAnkJzMqZlHLW42lMMPjfYv1gY989egnlyZcQg457pwfo17+Ut65Yh
ZJ5G5xlH2bmoIao6IvzDJiRUJhF8yzHZ+VBWPWrN/PjDB4wkfTsfdNu56s8OQUn8
OR9yGmwdtNS+/gpQJzumc3A2EJ6jggbthIArk/UoD4NBS04ncCXvm4dTQTVf6P+Y
IwencLRp7CZmNF6yJe/w0GL582DGaj30/wxAIgkNm7S29aAZTI3R84aFUHU3u3Dp
`protect END_PROTECTED
