`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fOfggRTUFyU3sLMsC0hotze03oNNuSnSJrr/L9LVq4GVK+ATANxzzYbPvkQBxxWT
TB7TU53EwgnGGn6KlpUDWbqrPHG6ahZgqP9Bik6yXf1LQeh9UPxMtRQK0t3YkI7x
R3PHhnXcLkDirZdHR7EnJrTVxfZ764e4xouYcnWSuU1+BXkfoXtNNYLav/PUSYOs
/ERJQhsL3HHxTDjr8AqpLccIlR8Zh8aqbGRrHqsv+qGUxSOlnDNg7UT8JxJRZi9t
SaIKVfOGGgC8ddE3EXJOtlVfDWu/HDYdgevXy5+qERROCmqGOVPJQVyxNrsY0G7b
/nUMEh9e/omLhpaL9ffj9SfLNdk6rKVglvHMEBw4DrirJrLaw/v07vRJwptY2qeV
bVJK+cbVI1ijMQMQISkVHKunnE5DWJ4EuuC6+OT23Wj1xV4i9xNG/pJwpDra+zIb
/iyn9Goi+M9oRQcSrSQAUlH0RPcMAz22HtcmC1zgO+eKi8K8kHgWbZQDoNRzV8WS
BveceMi6mmXpfcT7jMmxKH7a+QZ0SDkI7R+kNf4MEOofya4JdXzTOFSxqeQ74mrC
/ZBEmwgMhqZnnt4+TKghg499YbW13kGL0kwZadJtMqr6zQckm7gBSjWec6TuVMVx
NfBeTK2PvXxeokNkzrCLKWO5Hdz7crhiuvms9ihltW9aBjNyMHHLZvQTmE2Cq1ZI
2chnf+51bghaM9GzHyeQnFVlVsIN84rtlgA9uhR6/aikWI5At7uC2CcXmVEPfyiL
5mDul4JpR9YiD08g3QQCcgwmBI7O/NXUOCXDxyrt+exZDdqXIsGBC7NaCxCasGHC
+YV/9xcyGpi6iDyo/t9CCzikKl1Ag48Fo+yo45GAan8=
`protect END_PROTECTED
