`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YMNa2wtiUCIMfkuhekANTl2OlAKG6blow/0k7thi+GJgjhy59ItnNXS07lsDNJFH
PJxGboIW6eG0kG5ykQkubVVh8ycwchBVHMc1Gi9KE3PFYOGmzEGIbobb8XYgby7M
yOzrW4zfgSs2bD3rkkpLq6xecR2kTCXZo7SfYEbBevsN6Oe7ouP9SD+XEURotQNN
srORbewrRzFo7Tf6v19euobJrsbVhaUQEO4kv0SgH2/iu1bDc1OpvMfmOgrVzLTG
+UEMwrdGhHiB2tXntQvBW0QDX3MuZHOthuqrbiRrdQM/yAfSBpTANXAb3a2O24t7
+MMyCLqA4VBlBTpAi7HDjr5SK1Kuvb82p9QNwT/833b4NsU9frwDXEZsxvzFcKH/
d0S7nYNMw9xe3UOIIzA4HQBQDHfQDO5pbK+zkJolan8oTv8PE/01beW7tgWBM1vs
AQ/njo8v7U1z+dX0nRRAAoJ28PB+Yyz1+pDoBtQM510e790Pixomr9wUsFGfmAY3
WacNZmHvDNFek7jRryJHnVW6Z1aXQtDpokPt9zlJqDVakrDpAP0ma5alp4TBLawz
mV87rs97E/QGKzLhdYeX+sFqd0vi6gWP32nwpx/5NMuR1B5JrHcDTmgK5PvZY+U2
JJNJ35u63YRxPn3GWbM5l08MzYai8neQsyLKPaPhlDdD7YWpFQqbC/YpWRTTzHHF
vaMicQx3NPefnKauw8wLjaq6yyt85waNDs4xNBRTE4cjWbAtcDvDvCx8WezsIh9X
8NS05o6usUIPKOdaS3sf5me3AtI3TfuCLGtR8xnh8LK2N9TmzbfCDtZfWUuOddR+
DImcNZCgyuxjMWBXQqqIZ2lOAV3wexcEY9CBC7iqzOzhRg0Kg5552b2HGQ/xgtuD
17oEYLy5X/ZSkaHWbVbS2DMSZ9XXGTYQiJw/I4QDofUH1IX9g/RwbEw1x/mvVu+R
l26H2BbnOsOvXx8fqtkGWLkLnTB46lXwvgCaE7NR8fMXnva9mE7OPeTWkNyjxFNB
WRzfCIXBNnctsToGkqne5UJJxEmU8XCvZZG6hk9oWGLIwODWmbyg1NF+3+JkRkH4
yFqEXLMotTP6nJd3q1qOUWY77uXWE/feENRHg6xHAd78Lep5bAP6JTLJGheGkZoN
gZXeEUXlqzncG+Snb4xK0omzlUIyNboEVIrvxgbEntivrf0xylPje+IdSWqUGgVE
ZCiJV/sCgAS6i4gzLK+jnaYInTNE7KgIVOBDXPz7ItPoRhVtAAi+q0d8DXnSYeb8
XGsNA7JDRSC2msuiAjUNftv4QpRDqldcgCbPM6x4T1tfMolmv9xVv2IFWI6TdFw1
/usKjzWctLlVBujXR25MfwjfVuHvTl2HGvvF0ksMr41MwomiVw4wY0y1/kOLdSiL
5OD5RShYd+97Jn4PJ5Fw8mpePTjq7S7UL6QuEKlCj0pxYDexRJbVppvbOTq3rdVO
AO2K8kh9QgPlB5VgjY3Ws1PCSFoyd9zX0re7dgEHFmzI/tuvxOizPZWt73r9HFzd
vaKOp5k/O0Ewn3g85vVa5oAQLgIaV538fwzUkljOX9u3QlZicDcEthhdM0eznTGs
dKl3/iuI3AW0lWw+890FIhILSGEbWZgSBqUyxQmuTFqNaeWeV0UxR0ksFRMPwrcy
5aGQpF++1sH4mT7p7bYx93RHGIYZ9+LdKETM3z95RlDnJIcIiNYckPSXx+h6qZ34
KM3ckv2tVgMtXeRBn3sths912SRvXINQat3f2zE8FlQrURvz3I7SC3mOt5WV5d3n
UkHkMROKM7Dp8m/q4XBpxvy7tyYLeDigmoYv7YgyGYkA+LlNdJ9HxelkisyzFhbu
wKdNrEI+2Z+ciEejAITcF6lBBZxGfSnt3clkd5vgE+pTYDb0deDheQpmH2g9Y+Hz
P2wdVw9v3Cjia/VKnqNRIjnjXJSclZ46A26RIdhE5wjOQ0IMsUihpVLkBAVh5peZ
4YnqIn7qqKZq5iuCIg3t8csC4ro9OQdgVUQBeSOa1fPDKhgkDmtntz+pgyd9dF31
GecCakk86Feqzu3g9sAhga5qa3zlu4mmlSX7gDT2K1fnyFrzHVALI0D8UdQZzPgx
F8ZaufurmjlqNRKuEQ3tx7n8qmd8aarDKcNrI2d4ZXk2XpF7B9uULTNYrrrxvlGp
zjRmSRYe5rURcmo07bqPNuISl+Gma8XUzJVfoQWuLwb/RUzKWFdCeC+mxe3IJNhB
qjV+mCalG9HdWIrE42YumlGHgCHWAzhpbyNaPJgiDglLi8wjm9gPOOTeLa8b5X5G
XlKtCZ+gbEiXGwMLPLCcwSDCFy/en2uH9nDsElfrWuO72jWrCBSxu/85XEf51hLM
yy9g3PJ39rJUwUQ93B33kRQBCvwYJVCScxJhohibsRRVld06Yfg9hJR92USwHiEe
+j/GoymlVkU+R/mgW9FIS8QPr402LH/irCPZ5bRIEqv5AX+WdVP9T0dY6SlvOTgF
4JRGuiiD7fs6xjAIY1/b8b0ua8mrdwjMMO2aDx5l6O4BRUgWIsIpv5onZLrVtLG0
0tO0EJmAqqhZ04tQSLcQ3WOVKJJSCjuTpeh95O37zkwmHjDCdwb6xwSgOJ1wejlO
ok5GyxtVkxqeZNvjolxiaZ3z33seXTbZ7MGWx+UjOfeUdzA2osu4qHgfICCwpCgo
trQ+mGMuCxlj+spxQfFUlC4/8sX0jSZBWLwH0r0gtr90q2B0hMZz/h9ZwUhBvpl+
QlKkkU2Bvzw/DlNfK05W4ldY8KnOXZTRHwLF/4anr6tXeXUV3etEI6O8ySopM6ha
ltGQvzbX/Y4V0s410w9TjEcr2gL7rdsrYgTRkzmuFhzZT/1T5H67plJn9uEpA2y9
6E1s91oCDYuX8gZMy3aFqg==
`protect END_PROTECTED
