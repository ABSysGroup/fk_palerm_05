`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xYwWNJJv7u3hL5rLiS8eCeXHqjLuYYEuyedTtwFhNruC4OhNKwiJHAxhRF36YQM+
j48CpEVqFVhR76HnkEQI/8Fkd0U43L2YrleXH0SgrhEj9Ef6XDza1gWXRh3NMmCh
ChJu7uaQ4SoS6CGnDUSrZ/MrsG4a20DEJKQdV8BG6s7I/t9NQDrXHdvxKlpHy6iH
Z1YimXdPHmBWaennSy8G5JBzM8ZZwW2i3fEbrfnQCe5VzZhoCoO9N3rSM3mdXdQ1
6vM7aKXqF+1ZRYF3W5iOL3DR/ExcQwOp4cnCyXiuXBwd9VffHsxl0dTCSYcBvCHR
Km9sxvUo+yh8RaV+Tu/+7ejRfW6i8zp45a+JQpGo9NmWKnRJ3NjnAkZzl2oo7D+/
GXDN7mfWX1txs5WdluMZuO8MhpApo50hF49tc6gE0u1oIVahJiguCYh91zB1ZbR2
NzTix8yW6qBGEbzdSXBwWdtE44xZJO/PBrqzxFaf/XyW0Rjtr6EstB9oUccTWHkn
`protect END_PROTECTED
