`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aGH6kpkT/xl3RAYRMNnxwT12fwoVW+DbVtsnwW8X+nAtIPetb4MrgbVZbhRKg3aj
g9+GcVn+8vJt02fHNcAnXOaErZdcvQ8L5+Js36BFoeeOFG+L+aBKnncOOSiPj4/b
HNG3yKKj/DGRyqavStNCC1Vf6rbxtQxwLvlvvsC0W9omrgjLg3veym1xGD2ItUyJ
If2JWJxDMZgMuQVmZeVuJxOSIHU1dARP9RyRguGfxJf/R8D1FrNHAbXYhzQ/85rJ
u6a/b2bgjRdC+bVCG8GP0P0etKpfwrVKNzV0Z3CDjfUPCUA1YL2Ptkw3C1+kCXPl
vbiWi7zJ3yZxdxSZgeXf0OMpWUY5AZdFfI4WHrDSlyn7BOVLevKVetJqMDPjcCB7
DyqXA6y6qCVt8W2yf4cuwA==
`protect END_PROTECTED
