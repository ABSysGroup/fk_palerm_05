`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3eSx24rtNqI70GAz+6hlfy4NbnsNU2emO1volbebFlFtUMQ8TK16Wbt5OGRfcBpR
6e9TN/Ln/k7lfJyIi70DijCCEv07hYAZHhevOz9VKVfb7wTbLTR/13GY8UhnMGSB
a8lYXPM8t4itOAchDL5dZ7pxG9LIeE8AufuubzV1gj5ABKshXd5zmKBmLmAo23lh
aR2ADZDJfUb/5aVLPTaDtlR45k/aA0mkmBo6CUuMg39cj/jrL1ki+6nuPyq8+jbI
RSaKz4hpAk3nuf5zzgxeNgszCu1xA4ihFJnjjlB5Hy7OfJbw+IDYXweESGyTa10N
wqjlZGer12Ky7hosmnwSJPOWu/a6fvRQCGYH/FhCyxEUlrfzlzCg3U0uE8GFQ8Eg
YmIKQiaAbXac6u2R2AMJTEZY+Mv9lNbZ9pezgovN0i51yesWnGwmERmBLclSp2Yq
H08BErFCCka3PbJJ4a/ABU1NVDlnbXhFNq/NB52Nd9W0VgnqtvKIEjriQ8j6HhRc
Xmck1joWi6+lU26mWNf61y7aXxEMM9Wnj+9L67DEgOQn9Yi6F6c09iCPcTh/N7jI
XxY0/KtOZUoo0D8f18bCl/n3eJXbHbAcX0+1o5a3qnFjx58ofl/DXJcy9MVYcO2Z
obt7Vbk6VkYinBHmRwtZf03eXmX76rcrBIjUya5gRwozGQ/UMMrz87LzPo1JYnAX
1PdUXcGKWV1Sir0Hfdk0VxDSBPEcnJKMVySCqljLB5MYQ6z/9bNMbBT+TC7f9/Zy
4rt1MUzQJ5JsGbbRDx+YvbPIH11N11t5ff4Sq3woY8UiCqBNQ/TNX+0l53J6J83g
Ipzk95egcO+xS2vXLPHBFOksOmdWrVGx1VrqkvUjl61TOSB0FvgnW8FKNFCBFn1q
0O5Gjgx+B+9iWYJaWUSXQXD+R4HqH2Ybaz7XKZpa5K7IUk6kJ1cSjIOr4ohtTrXY
XT1m9I9wtV8bXJ2+OIjrHSQR/4HPunMPYG8pQvxPkyODrG8iGnLS/OO2L2HlWsy1
qHbLifn8dCay8ODowDOE0ZbaYomTVRPeh2Xk+U+Q5We8GoEkONBCQ5YXqGcYXHhn
QfCjC96MsxSZq7+BlPbY7oK33SomWbpnXAV+AzM48UNBXsuwTemgQx2hi1Or6MGf
HPlDr7aMGDvS9ZrY5BDtF35YSMtkLUXStu8xagstkCra70qiWmkJb1sHxs0Gy3hz
NixkBw5JkbSJEIHigiFSSBqvhZhtgEolq5l0Y32OV+UVWVL3nBKta5HLGu560lrY
`protect END_PROTECTED
