`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0xBXtA8O1At6lbnj2iR/k08oFMXqwd0kvSHX8B61RFcOuxxA491cM+vg0c9eX26i
wIMrrQfzqiJ+FeYYHHvgZGG7xlg/qnhRmn3pKJLl3v9IDTHSm6fQwRwWaSn6722F
bamfm22l4m8AfrhuG6r2QFvwiuibEz5KIJz0dKog7FJ44V4/oR7jSRmoD3kRQTxn
lxUMV+t4qIaoH8XvBJziipWrRkJ6/59iP8gTzbzBZGKRlvKcG1CtcNeusUrdQ4G2
HzX/Itvj1z3aFw5tnsfBzmnpVeibR8lPPXeB4lZS+cqLH+oM0G+Yp5McGyrxgytR
nSrSZ8IRnxX1+QjuBGCW3IdY1TR/2PEJJGFUy27MZavOqHaYO0wAVJwi8eetmEbY
n02q1AhbBIm8hpRG97GrET+vi3IAlRh7d2zbhNfsKNKfRQlvde0RFQMSr98stt4O
GyVaCX+LC97aao+jdvCQB93mqMEx4hEnyJApmF4zif0X1HnHtP+ncTmRcK2tMaRt
BhPoZlckcnXOqhdgsAWcpOTDnlf/LDK+elQBSI2yMpZlPF4hY5B5zrFOzzMxi/yd
vZpMw6XX/s2XYF4Okm6yxsO4wIvH2/V9229faG7NyA2cadoTtUrkO6gQCA0Zx30+
ef7uMW46KR/GP7wvBWk1O5bTUzuQ40koEUadb0i69LN3HWD7kTFU2tZoxuH3ZqrM
65iuV0qAVO+LVtihLDMp7oMoGFfKlamr/HojFeQWpEqc7yOR7cJ5KEaWOO1qSMpB
lGCtk6fTvoDG4dio9LYSvjb57uzzWLdPiluoBhFQwuXXQLbPZJBgN/8UW8eG1umt
+HA8UWFKuDkZgKEUPGmcdrBVBUuOm3M0rJ2crB3ZmRC4jKwgtdWLxl+UAXkMvcS5
mEd4m8wER/sFequpvsHTPaE+pV1dGU4A1wgIsJyj+qm/QZwaZGNVey6cR6p3mARC
`protect END_PROTECTED
