`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6dvx7U17xx7UfZAcBg+OtQvKvGIbYDOZcW1UrodwoMzOnrk0XQgB85UlLR2UyX6V
EdyPC4C6OXP1X1AOfki3kRTC+1+5jOBtMcUIaxBSAQiv+MQK9CSj+8CUyBnib5Qa
sbZx+iKhQms94q0yBfuI29fYjNHaEbL5x2RD2jS8+NNPHem1vC8td4ypsD35K35t
3op85egfeHfBF5CAy/LAMEgL+HR1A63gHysOaUn9149hzxObGyVGhfckcL//y/nH
OCb/bIqMoEdn2n7JZhoZ4IF6TwEuDHWQzHMHaik52JaOUdDfEwNrqLvyOEg42sRW
FBQiTwRATAejsrDZC6ZmmFqAVnXI2e5EKAjMAGCvnVLfMVDOEx+Lrt6QN4MCwBpU
MAPYw5liSR1sIdmDnCEJHl1CEFk161ixxyol5409RQFwpAQYwa7375pndEGEEgb5
apebrLq6Rql8sXPixgHSJJh1QPXSGtspGEgBJe8C1kL8GooWnedVsXoGosZFR3ug
Fw95BmboW7kSzjuevEorHZ9l8k9NfQ7wbFUMV4FLFy9LqrcX+/AOE1LSiOJmTqGE
6O7ujyM0G+m/f+PtpzHitnA6LDKZnN8VcKOTdIw2RKTSK9+Nl5LXfYVg9zb5p6L0
5zPr5qih7fVTib8Nxh4Ty/F4s1oW62nEaUShBgQwUif5OIXtomCQSMcYvnEWxd0X
XYR9GqO0DqOs8zK8HWR6lXUXKKHfiMUmZfaPGm7fjGIfKz8uau1ToIXMoe68/x0A
dnWMi1U98GAI4OD501LCAw==
`protect END_PROTECTED
