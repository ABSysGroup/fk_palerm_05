`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fNdCyAKfq/PvjAMs12PNYB3Xi9T26FDgD6oCby0cBABjXqURG43WmupaRU3RlEjW
ABFkI+ngQocoCRgTP6lYiFyzvTpJcNIKU2XJLxfu0zmRVU3sEryVfg9vWhzNpnX5
amjIJqzCzcq8kHPsLBL8H5+Gj+QcN7jeCGmh48Zxb/E/RcEOBEh+I1dpYmi2WXND
TWOZj62GPQ3WfVxnR3sKWyEjg+n1nXJQidXF5JudvD+18TF5CwIwGi7uBK9hNAid
mmJeJDGCiutMN1lzY8C6s4fgJFr89WWtm+E+TARXvA23mK3DJHfG3kGCjCfCC7Vl
ghsKg7Gh5hKum1ufJMAl+SusCSqgMTugpWwhlFxSTguecH2yRvJrA9K4XqkUS5C0
kDKZPFzwo3aF+hmhx365BHUsxsSpguplje5qakmZP/SLpG7M4p3gMFJxzedPv7jY
`protect END_PROTECTED
