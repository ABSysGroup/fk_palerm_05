`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cEj38xfJYEL1aoX77wM2vOjAY4R/E6Y2Z4H4rjIdQy5Le4E6tmaV/QeHXrTjQi6z
HUmwcWFu21Y5W0My/gwmJp8+kmBlVqmnyBZeVRQfZaKG8kLzYTFUuqre1S4xBirv
Wlzj+FUSKkJkfJyVnzo2aAm7gVQdutCuZvTzaRA52mlQLM06NQ1cD7FZkW+f7bud
8B43Pv0spEdphiaDABYYVmJq9vjc1Db56JFc3pATz8VG4zl5vE0UUgnWOefIa8y1
X9vGOBrfI78GIpZ8evKMS7HukplDhbj0Sf4j8Vi0BW5tv74gpb5N6+aiyjmvgLoM
FznWUTFzdXaN4c28Re06G5Drqq2tsLssQ6BwYRdVwqf/nhZAy/w92fUqAgwNAXWJ
A9aXjB+SXFENkpHQS2uphLnqtrr467X0vLnzBa0jtZqm0MhKMi0ap1N2yrqiOKO9
jwwrbzeyv0nszUDwmZGpoSdna2Uwz03ji6iyNUo1We4nPB06ffEy+F+a6cTfs61+
kEQt8WS5UPOndazgctWP8aNImqDJBBQuDcf5TDh2Bq01tsS7POzNDQot5ziNzGQD
INVqfruLc4D7xmxXXwGnmijY1RyyqVLqLbPJbQ6TLUeAUTQ1MD9QkxpO4TjvGtk8
mOrU2m5G60X5o/wPfEAqMM0KBjS+9hAe7g0blSxe2IKkC3VsCFFR5TOurDp5ubht
ND67s5r6wgFHSNISRTW34oaL8GHaU3Tn2BtxdThr8byuV25LdZhjlmxm3ApNKVeg
iKKAiADN0LJ/XG65z/Z+XJ/u3Nj77tQPje+vsH/2zHBW5pjaAqi+BTPUTWJQKaHF
28StgcI3NN51e3myjWfTn3wN0QO7XyTELqqFzbfHS6nTV+gy5JtUbdVHee8PRuK+
dpaMj+1WkrPSkJ0SwYe6o61GgX2h7dlMhw/tDIlq+FZiJEKZwiQhapoX/LA54Lj7
BHAIBaQZVsz3hGMvs/iEioiuNvab08myuksR4BHDljhFRRl24Iw4N3NtfDs70Usy
E68rvUCIJB7ur1W303yQ69XVOZ8rk5DxiwM9VuGN7B+SJ84YWPZ0O7vTaAr6ZnEJ
Zo9e2ezv6a1RnLcU51qxUZc+dB9Q/ph7yNMKzteyxrrv/TA69gxOb91hbJfNndDD
QYxkB8fbQ+YHEb97F4K/G6ScGlnVqaeo2E/MHhIqyubZSbGgPtJsOCjjbUgk0Ygb
MAD0QzDM2DjYvPPVZVtELr7TICOH9t9sLsmWz94mG1P8USYOpq+dGGJ+jEemvyko
cZ2DUESxW5uskEN5ZCWGPcsqY2fNKOJ+fh1gLVcY736T0mDFdSNIhloKGIndCror
tXv8zofdhniWfBjssbRQvy/sKeFDlKkoF577m1b/eoPRVX5xAt5H1CgomUK/X2QW
uEpdjBkbMQ3r0aNH1jeggS9T8zwOMuarVXvHCWYpwV8P+FVpAvN91h403A081Gzw
T49vIUToH4Ys+p+W6JpVfqqXdv9KjO7T2N2Mvwvm6VUJ2OsPBUs4+YJZwKNx4MP8
+V6yVf8gjXktS9XGiInFicYa8AVEgvG9RfWq3nTErs6zUyeYoNsHEK0TucJAWiFb
mzvqNbOdbY13hQCcOjaqY+RHRLLRL0wuUUm8+9o/vnf4+PfFzaEvgbYqv3CBe62U
dwVV9hnUYbiWG6LU3L8X2V+lvc1UZtetpSZjKzBgJB29nShC9Bt3GPuOqUn+X46F
GxWnDvXV1YR5buDmf19GcePgBZmMLD++AWtKT9dF5x8a/OkuUJFQ4dTUnIeFk6y/
L081cLkYy2fPU10vfh29CzLkSOHp0dYKsuu1H6vWYn2hqtbDm/pv3yQ35TwuZEQw
7IxQYdpwSWkxglLuqfIIJ6Hpq5EzklQyujw5/iScSwddFLIGJ2eqX0QS7hqvvk2b
qXsGE4pBGFZLhCyGzCxozFTxOf8U0QXhAcJwwORF66ejTsQE/EEsU1ai8dJ43J2E
41cnDXPWy8vGJ+icWpuUjmc//q5FeT2N5DWlsGvctvYw+2/GwKMcjQ8QFtgSFhVc
bUs1sSaCdvHGJe/mMR+uSnDz7Fa6pzkwuFLBNxbp2Alj/QPvVdIZcrkBL/3wQgZb
hRAk/zw3kp8xCVib2UPzQLs+3xa4OW0d74K5s0+6NU1GIidt5USTGKJrvxSrn0PW
TU1E9AAKZnAnNPHjLVbULaadtPwTiI5IcWNtNey8Qalx0f6brzOJIAUCtI3T080F
sAyqC2YJF8ReBLrDJAfIXQrTnUa4FXYid0fkyO1HtO3a/9yM7GEwjccTgq5YcvQE
5zFZu4Y9nfCcvR3vphF8DkXNROcw4+Aiifttem2uiv5UnduFpO4VIrsTzjFcAKRy
ORVEbQBSKd07PaG13SMt1+m6QlNTM6PNQawtV+nGhB6XaWEFX8/b5U29nJq2/nj6
Kd8pv9bbG+PLalajCoeILqem1hUtplwpfjEhl/6shUO9OzlGmXU/umcIe58z6csw
tF01fN4DGkNXAWUt88/HMdoBoJ3E5P0unkxHFvjHLcxODJ/+/JhJrGYRI3IkSk11
wvTwVlvsnGzn5zFm94F7TPWQ2aD3Y52TF7xNL7CHv8430jsc1+JAcEj+cjFu9kav
MZJCaq0EHalhrxTX0Gdou/V8ZV9JNFHqgQvGicv2EvPLE6h64uHazJYxQ+KBPnIw
69l1qy9mUnCPbUZtvkud/XajucSX7YcsbdUcEfLwGIdBYL7VhfgIMYi3MOaEZQRp
fVUifCuw+riSPvUKZQxnFrl9HCxFBSjJgLHshBxolP2i4ASJFX3cLUjL+tNz8i4K
kM91gq00hmJg7qVUZiEwC2E+pSWy+V4y0a/g9oDIfShi5WBY3aogodanqM/dFWu1
gOwT9EkPgXdM2yKZa6VloSIEjkfKvcOxH4YHOpMg5ks3scJHvd1zE3GgCOgTVYtR
Y9/l6IVCaJarLco4g08UypQRcUa9A+7iN6yy0nPfGm9L+MVtHoaBchGBh1mx+FJ4
`protect END_PROTECTED
