`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a90xEBecgCIvXOLKTc4IEGy3FO1Iko6SecpSGDZTXYOWUBL/qSFsviJdCK1y8V2R
PQ9/i/Sk8c9nmA33c14oInTvwq6/JqR4dlioK1qlumjsAgl+NmLoAbj0kxqh6GE9
5dUtQzmH1wEfcCHWtULPRsoXQn4slMg7G0Y0WyzDRt/2hi8u0+nfYG4w9FVfL5S6
XzVt5uB4XHWWZrluz2UCxHKuQnvPM2grvbslzNe3ZsF8j9Yyi9BcixomsO6hWWBc
0Uo5xAbtbpeoCNgTO61F/yztPSe5+JWXWkWWLGKbl+68+KUCrrsUeV6rgXGAsaCF
jc+rco2eZM4pfMxFFCELdFmc8IgIycuLp/z/l+CmC8SLqFKaA8ZtpCYeu0quDGeK
LFMSBYEsY50MkL+qTsfcBBcry+6nBxhhJxntItb2VVLJ3h7Tl2vlAIJLA2xPQo87
M4cnZUsM2bZ/sKbMowrhjmRZQcQtYvLgfGy8ZdCA+V82Oi3xgwqAgXzxBLoA63aT
k5pqU6/Wfy1PYMIx5qhXQOhbEKYNjs8J58U8sDVfVQAS8OzWD+QdQY62VYEwIyLb
eAhyC9D1OwPH8oilVO+kG/we0X7tdnF3nqyivbj+6U3NU484fOKt5123iotzCh6v
cLlo9Nx6qB1pSPDPwUrQDqsgMebfh1mj4ilx3Z6YgFwZvFZ0eLOLA1dVV+falQKB
vHc/WSgYF5WWyiaKatw8YyPzn9gCvt4J/BJKi8JkhlWDdvibNkJRl/qP3MWclOSP
KUpj7zS4Px8zoD/4ErA+cu3mHz9FEmJCoDAhigXMKA3fhMa/4Ghmdw2ifXdrW+DX
eERMQzUDv+GhbzvDQDmPVZxL15bOGJKkTjbBLJYbHymuUUjoMrrsadAVqoFZzqSo
0TAi0xClz1fSnm07ii7KvfZC08ByxAAVdoxIw7sJkgpU+wrksA1dvduTDzUj71cK
KvogoYC+LlyWjd0ans6ej1zQBc5f9bzcta5i4GQVVXkXrJuKwlPxx8B9zdQm0/CT
KJxLn2NMDPG0DMlOfjFwPxnVWOhiP97TO/oReIi3HccwqwzPfPQzItQyh4nzz3Rl
m023KiukcBdrRl/z3LepMG5dZNhfxekfUs21u7aQyXJXVeesOaLQdrkk6Zm7ebLk
TSdmS9kTbzMStXelApBtQZN/wLYatNgTaIJwZKwYs8ND4UZz+rr3oFuz/VHlH6pR
AwLQELsVpx1FplEA32YT067f7wRdCBWQC+B9te6tC4SRiMU/ebSFp/u/i0prHUXc
8m4hRSLClWSji5Ktk14H7FbBI5pDRuWTLacKVx801INzOOxR0phjJkvWsrgn29wg
YTvMqUy74wepw8ZRt8gHW98km1GFikGl5dHFln8zARMAqPR44CUxAeA5CpRX0nKD
oNHD6UwegfO+gdebYzPSHY7mPYL4XyVugOnYgMa8+AHxOIlRvDzIidUELqeFlPGH
SWNF/yUckj/7UTjFBcZ+mYFxOk4KZ3wO3f1JJmPQe8dLvysPHgpiAbED4rndkHQS
eppqOcFFh8K6Qtkhp5gBNjmnTZCDor1hoMRGVYG70pyJUTp6mDzq8sUXsj+4FmR2
G1RAKkIIBVa9EUj8p4fUOx4YavgiP/GZmUh0YChxaOObLwM6PlPBobcUyv/FBNBS
9XZTOMm7l6TsQU9MX6+VVNGc6Iwpr/IdrgNA2fJRD+pn3ZxcmBZHnehzvWmVqUjW
YiEON+IqOrg5ih3u7EFZKbbPoq4DtrbjlKgSNft7v6C4rLzihnuPJrv43rML1K9+
rQRs3J+nVL2TqAWVV/GhO8hLj1wZ3OVkOqMobGYvdWx6qqCtlnrfqqxoQaDG2K7E
Kgv0S8Aze2kcDD9yaOFIOkZs7V2u6T66T55w1RsNYLLBRkxT1hCwEmtOyKR86o+R
bbMJ2I9qgy/lENpiTDavjpW2y2Bwl2LOTeduNd8Dd1QhRyjOLocw+DWV+gXG855M
aI9CVmy1sA1AEzOLCgt5LGjE/DZH5DkZWTAcr7DXXWQvSYO2E6hb/lg4G6dD8meJ
+q9W7dChy0R21G3s55AeI2ftJN0SYUz7Y35XPXtOn91jhHpiWvN9pGjmo3UDONwZ
1tkkWGAr4p2rjwvnTjYqIW1qoU+T0nLHOfBwioTvWVoIms8f6dtV8Dtn/q8vHKuQ
ENFjk1/f6YgaKUOlnRRh6OpTyzqso2Q22XfIbJ6mAwdVH0aXpkV1V+8OYHI9CQ7+
aHOYUclqlzBkQlCd/DKtxyx0y++2s8U258tSwXsxpwv8fTSM/X3cYoz1GByP7/SZ
p6vdN0ReFg/lBFP8LOI839amLavnkbCQwn9obz0tiWNK9ad8PVO+GGCvXonCv3v2
qwFq8pYU+jL19LdcjOeYRD2S8mD1YQ3zRVw2Nk88Wk6/hxSFyM67zuyMojnQUSul
7hPl3pMVqxO32kuZWkSnk0TZHyg3x568VnJdAVEDQCk0jlt33A0L6OFJtcIjEgcP
Zqg50UFUxxdnn0/LqfvT68FI9rebBDPLFH3ZphiyCQNPvP44v3GseOBCAPJlMlRz
B67pAX64A3ZUt9AEB0KGj8D8Bji3SXnKgxIv25PwkD3ENUZVYKZeLD+OGsZT+ueL
UiMI96cVue+1HkkrA7RQhj1R9fMDfhdhYPI+ciZEw5zxq44jH2gjkVPDM1z0yOHs
ABsetvNZFU2DRWFWAGhl9soK4qbzpgzvOiMZ/9hzNK0QNxrFCGjuxEScMaJkYiss
aQZlLxfESsZB6WRvyQMzFb2Rr47UPp78Ea5rfRIuKDkFerc7cv4wMcu8ICchWgM2
V5IhcJtnOXIglfJkbv7aWsFeK2FF+JEZd8oNBdyUeFSMbZfw4iL0OR+tNdBOa2yc
OimMVXxN90V/UWJOoUh9ifkO5QB/ikRTykx/TMypEXY6nfRHLPM7CIqkWKxm4HV+
hU8vAL4fj9tBlNQx/ApbArGOw/dMoT6tW6JBYrBreUD686Xz+cr7AZ3BhAjPzTGp
pvNsqC82qn4Ri4LXqCKCjZJxHccQUXBUNFYvGHHPcZK+G8K/G9GBqf4JH74qpNBo
yJid80rfLCuv1yZyo8Ic9kpe+bFkuwkh/hmbC/I4FlDtx0Kex+fU9dRCSFl04JSr
6dRd0iV2XVHkmkxjpHessNH5ULBBHOJFU5H6RyEGvrYIpJWRCFIfv4xNZPy04S8z
TvMe1MPixxClURhqmyEOqIh78AOhFZdjg4LsudORjW5ZBN/Vidv9j1FTKMPjw5o7
CZ+/EVhS25vuFG2ByNn7YSx8tyhypT0V2GGs/RMf4p++MJFbpWOY4JZFnqEeSWh1
T4XCV3Zqz4JtK3s2eFHhWZG3zRLW6EdFwp0JtecexkzqY3pZAKxbwL4agcbn78jB
QH1742ZyJw4+2XK3QeSEu1Hbl64pqIFTqfEO9jchvzxvqHdihAjzI43mXSV6yF3F
x5cJ+VQGuYKlLrdKH5a7MgO/VQFkSYf0ugsEhd9NVA44L/hZh1T5k2bCZlBSVKv3
Z04QbPLzKqO7Hgr6WKMKS23svZBuS4XziHUW2iF89/OXoOzXVa3eN5az53eCjOUo
cOVKPJy76h3R/Tv8lPjSZLlBtAsUUgT3DwM/vh1k1YW9kNk+ToKvnKDKLJDPfeNh
2DeMoxpZw8tgXaV3TqeAbuRXl7r4kWhi8hYB4weHh+hptWvf4mV+U3By6Oj9xbtp
ZUJr3ox34M/IYepzfcg//ZJtwMsylGxT6fxaBCt9OO9mL1lHkgdzkBDaUYpEIhHw
rs0BCc16dz5Heg6VY2CKngi/tYjehAqDLA1VQnFF+S8H7ZBj3Opv7LaGTl9eDQ73
tEw8S5jBPId2tb4bUrEM1sBnIq4/c4/ZCTG7QcshgT7BTZR6ywMQInCpO16lMae0
nEO73ZrD6q6szHWZPVqZ8ucMylV5XUPtCqypMdpdQlV0IOOr2USsuZaQF34EvU97
aCSiY18bQcPOiscAf+hSwHIidEaqxU2+zOTclVxgR82T/6TrQgSiWuRbhN+R7zN9
MfHBzkgIv3hxmQ5f2Hbc2H1CiNszkvX5zKwlQoBoyCYozqCQaKpfXFgR5fTUMWQ5
h8itYvD6ae1Zon1Pv7Ch3CpximwJ0CMej0ug1KtUXTRk91NXX9R42kTQMBzLEUsQ
yxsQ+9o90ailTOiY1y2KDmI3iyUjTP/w4qxiWOXP/Ykls3Xd81lhz3UKiMHiLVlM
1jtd93p7m/xaIm0FL0PC3hceNi5r8djAxMVVUFZulhoV3rL+8TeL4Sw6ZylkYR7p
Zz8VnZ0JiY5sBROBEW7XlbxB2csVoJgHMBR9nJC4httCLadNpudZR2Zo6n0iPR0K
OWwfEFcochNwVOO0Icqz6FH2rD/8GcrkULvPoaSaBKiyCNIZv/jNf+K6QwoXRHfn
7ztNTgyyiFP2/bNSTrG2qUFtcNbUEJgZoviNS7rLhmWMenewOmCRFVWNSF41l+Tx
eGR/PCTuKxpJeQIJ2ubxgzaLbErR1p8cdu+fnJbJjp8/sit0mZEJHTuN+8fwnVg8
nxE7jpgBydaZ7j7tKo2DSbOycFKV3Un2sthzAxL/E87RoPUm4LVOY24JUkLxEepv
7+ElId/FX817bDdh/oSCIrFOfBM1LeHcW0kFIw7zZ6JJf6KbbIQLgI+fYfnMWglD
qlt+kKP1gI9xkkBqNQIjVscWxHpbtfawIL5jEyaGVq6UGwGjXW0/sJDjfaafexfJ
fRCdKqlttS7aFKJuflTo/j90xYRpkPaQBGY4FtSYZ1U5KVdhEGjih+8NgtcN8VEN
l03l+7MuNPRWed7NyaAOEqT8aJ0qx4nG6EHhMqp9VptI78FVs2mhN6dG1y/Jrhdf
oq8VJmU8+jFFKix9LjL4LPlPUftAPk/lPQvZtEpaBVJFOJ315yzaIvwiMKsaYF+e
ufTUzykxMD1xtVMKdekD8xCOR6vC5I7SqIM10K5CmWZ4lZP/8NET6p5xlDyxjFe/
mQSb5yjmKOWtYTFUsIjqT9zElU/jdLAxt7ZzNwRHzmQTDJtyW+XqTIRyF2h6izFt
Zq977/WSNYxg71fbhdlaSM/81Yw1Qlnts+Hh964LqUKjuOUcAeOnZ8UaNQ5ZTZj9
FkmTSYCnFY5dbhOa0WGzw+vrMWAJKXBVZsfvI0mFg0AUIpOoGLvUW/0+hsjrWgGO
I5tMeN6TVve0b2HCnqnvUrA0Iccx7rEtaPf4xXPquE/oLJpUQ8ZnRmqWCVmzjdBo
S4BaWPFCFQww6jobSH6sECvroNicg1vG0k3K4HquaiYdl7eHh+g2pqWFDa3NLVRp
F3ujHzNESKxFJB9EuMnqaouAAe3Y31lqj3bh6eF8bbId2gWKuwOUjrHQDInuXHHz
kPBAGM/YD+QvHh88Ol2qjbdM26Nl2J+YbeFVCC1s2q1oYdF9y5vO9hpbdaXAgci1
fs0sXiaqSgPzkS+PX/OiB4Ls2LSuIh+qOot/MY4PwnRKTkSGPmE4P/srhqZmqwyV
FEm5pipdbG3IqJ0xOl5mrZcVtvtu85P0MCrCBTRLV4QPyW2m4RYYegwLh8I/l2gy
3nZ0qv7qlNzBEamurvRRkr6bD/S+o6Tj2Q4educGQZTcu2PJGGVUrQMa1n3rUYIi
WGPx5DRmbZOjBPZy07WEbRjfdhyKBil1+ghIQCmFHrDgS567MWcmHmNReDmeWc/L
ZmXtAsKCuYsUpuca8YrzCotKe+zQX3rWWeYNiHNnLZc3VAi4tNvHImN9GsPi8Kiv
o0w5cWv9RGkVElpdqwM7N0mQwEmrpICvpKhi0+sIBxJxe1DIh7OmJbLpa/hb5ojp
hx1kldJQWAlKIDqZxMdj6StuZHUaoRg5pCW3geHGHIEIMj9qxLexYaSR/01gI+dG
XXrdjGdQnHG7crKesmAf1gmaoylVi4apbGjsLQ5zCcqqn2lxGzC7PK0KrhziZ/QZ
bBqv4aUdNKj0o9DIVKJQdX/7MVCTjbZS7soY4rFVFzY2d1Mjq898rRX25pVhfbdr
fudUD2NluzSpwgkP2J0nhATY8O292p6xSXY6v75OrATxPgGhPFPiizNy7c0OAmAb
aQYh515x2ecDijTu8xWUyDEb3TnDZOyIw/PqxkD4klD0PRZvX+fa6CcUC2gaKRR+
CIMbCSzKRNrZZy/+V6b7jz8BXhdYnRCrm9V0g/2VLtWzLYOyI54QoZ4nx1LYN8LK
xuG7IsdL8rf8tIU62Oec/XekmSO4HGwoEbaRX+vQYRbtaiN6VpPPhWbBgwns9qOn
SGWgMrDiep2jdhytnO/IU3Z88FP3OmzkdQOE/2P7uh5Dy2v5Ok2zo1h/6SFBAkcJ
TOaq6cHWK06rX2JcztyG+OGXWZy9kY8VKUxhswSW87WiRDWz6PIIII3GZhSCHt/M
UH6xOX7Iwhc3NDsxlP9fPYj9UjiFb4fe3/E6x0g+lqspX6FBXsJc8A0iSOR4Ib0e
8YeaI1TYi4+4ppiihso5IB7r2HRhBMCmLEbPkCsQ1UPeliHRsK7ZxjM/L4ytX0Jk
/kC6rCc/R2YlU65xwAIF31ijUE5HC35WX73yAbdjhcfzIHNpgnUQ4eU8ecM9J67E
GFIoL6actxbpXGuipFWmIHkeyiOsJwBkiekCKp5hzLzUEoppFwwTUtCYS0WsId0g
ihlUY8Gir8OWxqKzKpd89WZ1A8qTCS3VXkai19HJUS9mFbb0Q78cvCEbUSH7zWb/
y+jAYn11RcEI0YCfkn/+V2FcV49Tkk72BafOGsLDs/xvmhjO/TWs8c1HLwh06Llj
m6Eu9Cv5v/n5YMbaamVuiAlCtFCfKogmGN4OUj8Yh8n7hKDhNuKYH4Lgq71XkSjT
GD02rpYQZUH4TweTiv0LWGEPMWpeXquJZ3dSO1QkLTPRzKQf3OUXCFdVJTftqAah
C73rDGms7SFblQAtf/dUuRLkiLUNnmW0RAuC6+IeaP2HnInw4GAVHnDr8ns0EXm8
r8GP4r/zVDPmvVyRhjWnYCKkdkH2evkSyyvXHJ5uh/wxtzSU0sWckqXS1UFDnA35
7JFHAaAYGH/U2VQK3wGqHiPtxo3sDdTstN/GQHuwzD87wRScpblsj2EwdoQbe+31
Nv2xZObQvg2ADZwaQ2mUOvMJqacDlKuFlAtY4e7K2gBlszAsF+y5cMj/k4/5Ttrj
SsJysMM6dnW3rNHJmS3EtrDq2wZwd6EzBv1cYFr/sE+G/PDbAMz6Ap4AnULdpxVQ
DhH7ZMoK5co01no88R/6udi4jDko4l15rt2EkTQChVkN5qdTwMemDXHiQYcFc1L5
dtp95fCyrM2pFVsetfawRH9++XMYzNBM1VG0zYEqr2dr5Wpp3mYLUkuIn/s32aAe
VleDRa5l9eURN31EbDGAYJxEBZ9aAZae/BEQjDzZ3ZIysEqF2nZftmMlZ+wmhg5x
Y1zWPRFkM7Y6ElrNQ+vdJ7qCSmeNM4p7DyLfGDOiYBVh+3uBnD6nXmKKZijlYPCg
7DF2nQmtMUeGmy1GYEu29HKdb2TAd3kbNxVvxkOFVfCB+pMlLSmEUHobPBtmFoPH
IyzUmnQw42IqkqzMIXYT6tDQbGzR2Ee3MmTvEjy5zbXL/BUvsgzWP6AGZ0wPYfUF
Bwx0Mmuvyqnbyqbvl1NagxpFiX+xmyPeSWZCRk1GT3/Wr6MzMqH1HWKzSV2yaeMX
r1xpleQCdvRlJYtX8bTHplsz0rECJdvIGUvbMWNzRDcK8n4/ysr6SMFKKyZKK29X
wIL5qnCwO0gbc5Eq+FZGbfpucB7BqciHXLUCJSRRw1Yty2CfumJF0GdvlOXS32L/
Lf44jplZWmmYLdajxIb20KE5uqBB9jLzLYpkIMqQibnMubKRYuh1hhXpD+38arqm
2psTATTNXWNY3hQxvzmVAA8d6ywnC5/zrvWT7CTyDeqIRLaWpc0gjhPmM1cd53we
1iv5zBFrujl0oJjchJyBUrgmmRuw6F1Kr2gGZdhouHsH8sPZLytW5kzcXAk7XFFJ
opcjMkTGlmZ7kTBHjy7692W+6ktyzXBzvFBwDeRAMmW1Vv63nAF/LrniyxTyxCJN
F/4MgaNqt5piquTnlgUSw/lEgi0XiY87SL3mM3rX4QMctY0RYuEBDWow77/Pkefa
3jgRrPVYvoKbOEpttgebKGwZ4K/d8V/rduVvcqJJw4TD6bLe+/hc9G5Y1Yp+52kF
DrJbxf4U4B/hLWJ2ja+a8KYR414D2BmfoGti7/oidRYD17tQFXAekVIQD4Zc3Y53
zIMyZ64TF+NUdPrXs70K4+PcmkcFXsuhy7PPObuUnLjM1Ji716bEs7z6oJCVGqSj
0Nhdqp+8ce5WfHC9Far6Ip6QHGjO2j6zb6GE5dY6i/qERHUo9e8AYDbTF1qu2ZG7
Rl9xXFXkdZBshSqwlsVWIBPYfRJaNeVvrrKQTWMVbZiTzboz7T9hkSzLDMcO4mVN
82FoWpdKDGdMn84XoWDaENEArnh6BOA8MrcK4aZ/Q/cif+WVd9UlRjgs0SQQvAXb
XSFch+FxeICjPAUDoCd2EXhIKWRXA/4bYn+fZa+QevdbljKNweZmTqCePCWcAego
z2CjjJNutbDpksSnd/Gh6XnUaUS02FLo3XhYreTBXidPgezVXAbL88rZmDJ9tkK/
c6wMoFRKs2GZ5i3+XPWIohKD51ml1Qf1CRmseWDrvIu+0d8/WGZb194NdGoLNpcM
XCXBNb8vWuPG4GZcnjvRKOU0M8ZnUbvC33RES2xjsafkRBRZA1n4xogQTZ+IVDFR
yhmGDGERqrW5+m/TQ8E87aml8yB4+HhBbF6zkbNBvaztXepQJSqEPgqSRHw1elmY
0clYvAeIpIYIpVposzl0prSe4DDwuOQw3fRtUaDRtSaarQwDIA7ASBs3AT0Nuasc
AueF5MAtsyt6xEFY8ZrTJt9KYqigKpSbasa7c33t7/9SLYjA0zUMfQ3VTp4rgBCP
j1Vcg+GqzcnJO6U1dPlA1vrk5B2TsqteuFZuQja5yF+M31Xo+9idhVzquvKQ1OiS
R5gIhRnKJHRA6e2T3xYDJO9p/70JDoGsQtFhHDdOW0NFsPWhwaD/ijHoBHLYjn9n
3I0Tqip71fXPDPu/h6fDJxTAGgtO4H46jD6ykbHsUfCZDOwIVoI16fQ0DTIEYuqI
cRe418cScp7vWuv7h358Q1La2wCxKYgClReypt4ASfOcNryNHiQ90l6aQVKnG39/
emh+xV0JtlL/jKYbm8jtbsgE1cxwIEqgfE9u0a6H3w1HMrfqwPGVeWnA+VzfvWrq
yuN+WvhaLdgGlEG2Y+stJukd+6rEpGEnHSUFWV6f/sTJSx9shdDIGYDbDAY3RALI
DHSystCr/YQEggNJOw0j9+/ap/cBa4JkJ10Zd2Ury3Jii6yicrIrei+zLmHW0py2
GaOoXXI4dofgZbT/IalGa+TleXKcMRhdd7DXnITz3qqnIOURgF9w/lpzWTSCg/4M
L7svCP2awQcsknO2oA5kzCMLzP0gicJ4/0GuscYv92ezSCX1VmJVNXzaoYbPxujJ
q7U4aai/STp87Auyk3rGQezSUdnS48l2tpqbF2hxA4FkYqPshKPRz3aglvsxUBZe
EjfYq5GHlnXjgrLKYp094N1RJOoStjnuWqpXBRpPzhLIrPrlcLLWVHVrJRDaV65D
qecNQxi9LN19p0P3KAcZnAED+plGDsA7Hxc2jaSlr4gbK4JARNKNgyoXwn3AcHaz
GMyFjCZhvby52Nzmj75qgOorkqwB9zsKdvsLhYpClvkKNEsmHyB+gql+XRggMaUo
+o1ijWf93l8PZrXNsCdqqVye+WYNZCdPEfIWu0PaCIdPwDn3peeLnPO1Pj5UJG9D
v28pMCrYqtDLW+DXb7dEQK/AAsnZga2fUkPr4tb7hVWos3pFPW03ZVaM8lAD5fva
f2GwceLg/O5oCmApjTAUGp0LNl4sA0SkRkyJckVEdjNQTTXzuzWTp+Q77wRJz4Q9
07+0pNJwylrN6E8q2BV75z0NoBXBQ5GdM7mT/U7Vu7f97Sh7EB4TrhoAdBBCCu9q
ZOFuRvMH720yBfCbpKi5htwMMRzv17eDFR7AxbFrjl/AwEGYnzo0ETz7yOkFNW8M
LQJkGwW8iKDlP9inqmjJDC19H8/zoClKrBny1Au62y3AM461HUxm4fjoNFI8mHO4
e2cufMER6PdrRMnoDRR98N02wB5hOVUEad8RVLxeESt3XUUV5Ll6VngcJuBgAOUl
td2qf2Rld+QX6M+ZwC41HgeibPuWDAAyVC0mNVlZ5TIsu6zPc9sV5tIhYzRJuKGc
QQjkChOUguLAVaoqk33Wklly/wWVNLcOE6j4vT11SHu6zyFl5jusA5GF4FpGWvjZ
b9XcuHVyBopHMU0epAiSvodRrFaTdHKuVTqwJCf1kpx9RJLXqk06SHuYbEAKM829
SH8VitKxBMseM6noHOuJLnq75WSlDj4lZEBN2yHd44Tq16oIEZM2tlgPvQdVjzX4
hNTd5aqtyycc6hVv71P93s/zUaw1KP/3q0XnKVE/xUb+p8kGZ5nsnjpzU69FXgRj
z75SnkwfqvNot8OIOEeRG04ZsCba8zWLaUZ0JGzXONUr3xwaEyfSNWVW3Jt6ZbVm
a2oWmcWB2l5+Etr4qezo7I7izI5ID3uur8MRxl7AF14a1ctcvf+7HozRrSdg45Ke
zUzS4K0plzFWNYS8yXGQrSFBN4jFtuorhXZ5qBgvNV1WskuSFIcwjZV1lRhc4TF6
REat1sM3rpfP/4nzofXxR6BbPLOj8FX2xbxrjg1maXAc7VF29fRf/WTy9YGxKzWp
DGT/bYBCzm+ANE6gWuM6TtwGelbapztehh+xr7b93a8NXSYEIyRS2ydz8uK056Bj
aegAeBWnV6RbsJCmjan0mEQwNTEI0LomW+6aqoULiB0GXcADu1qbeQ1dqJQLJR5h
6sN41hzls1uYgiBauwA4h96OridVtUA5UwQDN2x+3MrmP67mP7BkyUuws0qmyeI2
kqiGoIGNDo8ZbEaKj2f32Cw2oClUJzSMEexFuCXz4AAh6aM+jfulHhfCUzofd6rL
V7+YzItUoJHIk47eHvW3ckXLw1WgjO3li/B4YvScnGFMbM2DhZ5f0U+jypChJNsx
yb5iVsID2NIDvdEfWkXMxWft3TFFuBTRPZMjyLSLn5CqV4Gm9RhQjdUoW9GLXqTR
660ZfwgurzP8MsOLiL/FRXEn4831bhWt9qZeD3pMqTAKKrjrgS2eJuIm+L1KJFd9
OiK92Qd7kuUC07M651oOYWHaFmj8zEWbXVxfVoKNslbMY03Ex11hZFCAYh0ZHVis
3iK15y+YSvRMNTvFpPFro9VEmodkO6qF47xD1nCQ/jgLuPjWSlFT790Ii8QjFbOY
gsBrYSyYc6wH67fCDyYZDXWf9DvlTFjRMru+RBE1e4GJxuoS2q5DyUxNx29iK5ND
Vpd31tOvZv4zUdekx2yDymfwPcejChV/QN/4gM1avEgwGccpnLfwerEUDR5oHS2Z
sGKSTzH+Sr1uVq0bxKmn8BFma0CSu83YMnODsomxueNvWFuChFIeNXlyrc9ymjLq
hd33PoRY2Y8jh8huSYY7nPr9gZwqNrf3nTe7Fm40huw/xypIQTIh+PcIGNyy9t7d
56kYkv/UYSknEVGbgFr2nrEz6R0UNL7yAxa3ABVzRhy5k1liyp0/txlnFddsbt8a
7/IJb8hFUr6XwhGo9wG1wuYuYPUctp4X0HXclRk7+3eXYLKjw/3qM72d8LKVld0b
+HrQ7TBpjE+LeklnSSw3KSetznHcZJo0yY28AWPxtDHo2lckjUadxWmQfk7Cy5J8
8Tkq2Lg49wIecSHaPznRw14y8m1uR4jAop7HAT6WuFnOuAw6spM7mgoA4FAzPFY/
NCpDg1nNjYC6vPZB1SKedSXNsUuh9PX5xsE4SeOxyiZlR9zhcBAfDi/rIY+jV8io
GOkX+8bshwh3CkoxEKhzDQc+kAIe9nwICPlJtZIJfsRZtJK6QrESkxZsX2dZNv8L
7TmZs8bTaz3c47hXaZtrn5JQAPQBczfz7wfeOb2sHVpQs50DtnkzYgM393gKscLy
6yrw0e9Y7r2RAlPIlMqz/2M6wCoNqD5CWJIyBCGy8gGFpVNRyIjEvIH7VBhk+Hwc
pDTZAxTH+yiAOT1QAzYWowQ4cSrocJzVbG3UazAaNM55GEHU3QpFlP1J1DaQZ5/Y
IO35jrGUQGA8CkQIqqBqwqsSi5bT2L3DNCLzLIEQRAzAXYDK+3f4iTEyHYhMyM3m
tmwK502nYq4L0Qgqf/3S0AzYgr4mzUIB7EgMzzRPqpzo+Wcfo1sTAP6SNjqoxl6N
ZOtTC97PATotdOCRmu8yBm6WO/qIBRrOMbUoUUpOPwvTaj81Esbd+/ADoRYZmWwG
ecBD3WRQTN2T7DONCAr8Rm35rz9ljThn7VrOGBf+wIePEV18sfQI2fw7IH+18NEq
lhPOR06LoXjyfi8SL+kYnkJ/PAIpAuv3sQhwjgvBhRrEIf1Cm4v6pOnnzG1MDsUj
/ZDEr1imPDPYbrnpwcZj4yNMUM9cmeEhPt8dqdD1yBegjCIJ7V6/aGJCSNgW+87p
sO/IIviaWlt8TjKBql5lhy+9wndaT621T3au2JMdEbEzrNYpweUNJP0UP4w8iRg6
+cEXT+nCW/7w90Bb/lETRreV5UGZs/roift9MgMQDzvOTB91pzaJECA/XROLHMhd
HApUbPuMu9CT/aOEgka+VVjwbEtfudSszxi4YdHDnC6qBhTTSET7feREGmcajohr
OomycMUA80wbTGSFQ57kk28+5HK8jzFNHNlL4aOtVmxPONeHGPnnF1z3dowkJGZu
MCzDZlXEKukTJ9lscsUS/PwMTS9+TclyjPZcbnf3nrO2fFwAOL3FERO1p06a1NAj
Y6vFT7ArRy9PWkjUL5lslx+qHfdZCkY478J1tCXxwcjqYIx9wjJzNrf684u/cV6h
ReROyc66RCZKbqx2qvQUAYXsFzzLgYGWyh662kfTBMbSjH/w9ISN6njhzNHPD0R+
HwQBfjJGfwM9jiDnS4eAUe4j5pITJI6rj2AR88fycFg3c+h4l/LYv6LhI9b23Jr4
U4PyNFYaj4rwWo1Cil4jM/Lf7t93mnlvNTDTX1O5UgffflHiE+H1kIHlKYfckMA0
I3rOYu6F8x9wICHe0G2O8mUaNuJI8mHlEo/eHpTxiLeuxSGa6sVUzT2TGMJQHq8d
XaINBxN6We5OSrkkmelWvfu7ym2NUZcndqeAcppZoLlmcPb3zFlj1S0wCtYKeMuB
n+efazxmY6+unptEDN9MGcW4q8sHf6TT1fwZ76TxoeZ+M9CBlSmgTPODPXX15pot
aQe+A6Q6Pu/Dp4J8ULDkvKjvrQgLMlKKyOFTSJLOM/dNNiq2cp5bBTjj7zRWQrL0
QTBZnJy3fAOAwQrvLzdsn3XvRV/yBQGEoIA2g6XTnTLkJk0XOy01gFjLlifbmIy3
uK7kel6tldlQ9me/ajq5gUbTPTAWwlI9IdctbrVQQuEVzfivjSIHp4/ninic9vtA
vqykJm3jTF+u2NXgb1fFYnrJNKcezi84SmIzXEUCOfg5ECyQ6VFxiIblJBMEUVj2
aDJ6k0g67/HDqhKfpovwCzQRYxvjBGpxGE6J2E1DuF6KMSCMOZwhHz40PIuLy4+r
tiza6a/yDrFzTjT1TgTNRkeTf7/SsrC1tPjfAGdoIfUHK210ZiGti2xOegaI7PJV
XTCpyM+SANMg8QjAyr98w9iw3wrDD5/NL2wTs7NOeZmm8WnpwFUAFCUnITyYjvsh
fCIA8cCOvxD1r29S6XMNHLaQGeqKK9i0FGERyfjmldXUpJDST1jvZFdjE+jSE0yp
6MqIEWSOFJu368CCUABR/gIhJro9AzNeitqEjEKYeB0JWw0L+l3YuIx8YZDVlda0
4poSWT4fvCKPb/a8Pib/BfvEAtQ+1odG+FGWAz9y+Ew00xbYB5ElFSI74xZuAmp4
tAp8JNJibH7zNgXLWROPmA6qN+vZXpV5enVkzznHUFaGPBqthTyIkHNO/jLzqCK2
wSibKOpMvEDC8a4iILRRLlVRA26TCZkwJYSoc2uM5oRnA7lG4qG5x3bG03rOA+X3
7E+Q4kqTpQKnBl5jlGFAkQL+gJOO1dKpNrZ2l62ZmxxcR2AZfBMwnn+AXl4DqEsL
xU1AwgJlpgG9rsvLo4Cl2KsNdNiNTQECeffLUytWTgeufYJA7p+/g68+FWcP5VJO
r7CXzTidvha2DGnAka4eZBTrFHZ0S7ezX7NC2QKWrN4YZ8f/ReRFLFOK0xSNreaw
q7fucA0EVDd5HnPM14sdHA1Tng2Rck2kcMcP/EVwrOw+EYlo3x43EDzjqJuEek4H
5QvSjjXLt3SIdm4xwun2dJPtuL8d2daBiSLh5SRKYIfbIX320F6sp2dWTNmTH9JO
1QSvfeyPuG7rb+Okb2jfRRB6oRRwGhpaYYeKGqddvgFuM8KbS9Wvbs81U1ldZjyU
YGfO50JWmNargkvUKGu0Ye4/l97jiwdodmkOoG3xcBYC6+r7R797VmpzIXcVsbbw
xCOekTdc4YHP/I9WYnJdsy1VzUWSaDPjFNphorcgh1NWutHwb+S+xii4aWOL/ddJ
+bff4qezRL1iZQwU4pUOoVMGXlGOZGZ0stj75H50mAuz86Aez7aWkjdzT2AS7k29
Egm63ZupO7WucNSeX6hG1oaPerUj9HEIZjAPZnoHG+y+H1RAd0LBrOLu+7xGP6pV
j6CXpqpRrAtPEp7jATq75vQ9S2J3dr/jz+KKt93AjtvkbZMLtMQ162qZxqK1O1iK
sI7GWawrt5HRa/agMgCH0NT/mfn0o0M82amJhri9CltkntK4Onm7MP6CapE8JXZ3
b2NROPshnpaSLmvBrfg0l4XkKAlrHm6gLrILHI4sS1Ri7RNhWH9ep5MSe5pjeIlz
SsPZXkxV6y5BDoSFj8D0aiBN39+peoMffv8KNa/PL9Jtc1q81Md1mfOIL2jigaEu
D6Bd99/CPiEytEvmK+lo3C9X8LEBQiQGFe5Jgn+faahIxjuQ0keDfarjk7uN5RcK
UbeyGfAR5/hXltNFtR5PtuNYUHEjqLpHsBHnaU1xzFetxRYj7TqvNX9t1EoCIJqZ
QTLg/Y+qP3xBEghBDtJTPlpdHvKPULBtXIM3x61nlXknN5sdvExjPwckaaGdKneB
Pwy3S+dGMCqaoIKJkoTZY6wqxRHFb0228wiZGQuLJ3zqhiyy5yDT1KwidB9J2PBj
auyKeyujqi9U7JKxZ1cugoGLFDJY4zMDjOWIdxLoubolRH2t7epB+B18il/FAzUy
r6biLimReFFdWSyo/bkTNwqsff+1ozrvcSL6LfOkLWM8A9aurSv9Pfc7wzrJGx7e
JIUlutQJQEvvoW1HmYQQ3k0I7RvpWA+12HlelZ02kp/oG4fh7CZ/P0ZYLSX3UBPI
HjmU2a/vw2ij8xe+QKlGNa65Ih4VhKmD4FB0k14iHGzAPYSchpMlAdJndogsv042
e6T33sB/RGo/X0xkJbQSxKDeN51lbgWqBA0h9QtYgYReGXDscZvlo7nDHoFGQ4xK
VS+J7VuENh1pmW4MkVMeVYgVAwe+6AvMlWy/HNljEf727D3pJyO1I5JBB2KQCUux
oA/xvaAEyvozfmZ78fTugcFi6vMJC1ILbfexUkwtwELZTXGvDu7D2MlJpaYBEMfv
diYUJPu21sDpdur18qWRlEDfrrrG0kqxlvALVeQ5YAIJ/dpZWk2yusD0qxQaXl+L
2ZhxlO8wcifvvi5x9v4raBhex/MQtfd48VzpSfPCBSOS50qrSqt8MREBWrpvIj1w
OTY7bd2tlTOoCp+Nvm/+RHig9E2J1hSFBjp2szR37f60707yoUDgBxoo95gRlzpT
VN6CX01NghWemhHyTSh6DMK3bQQ8ZO2V9vKzSx5xKo5YGCOwDyAth/Ccq+fczFta
i+Z/IEhZsB6tlQwrEbBd50A0FLubO1TdjxAOgjLhCGHiDWA3qjOZZA4RUTvmires
Vx4tiU2BDsRhMf+ZvW88BZd6jivv5WqaeN9Rau2k5DbwDSyo1ke5GBGst95bFLJF
n5Ol/sLxpaM18GoyIgDm5TDaU1wt6BLqpI8FKPpmFSBFE/AlLja7l7wNNh6PAx6n
+/7Hel8DDPl62jMZKWKrh09V/inkj/CXga4nZCs1y+SWu2txBunh5XxZEIUZbW9G
thwk3jM7hb7YLfPKZwx6+R2u5RjJnuHjrMwsXB5EU9OpoR4eYyBHBCu7aUKHNA1I
z5R/XmSWuymmtfgSvgrXMc+x6w+w963DeQQzM9x2jXdnZiuV5jvQR5gOQoRCTwHq
K0CriyFhN6yMXeFk+dRqrXr6Z9wrs960Ow7SgCfM21ViwrmjqvrzMx1zj1PcNJYy
ntNR/7/pmk/L64ZIblxURC/o74WFE+lHvDLIetuGP/SyKaE1KLAzOfRPL1HjOFE3
PmoJR6nqsiZVpzhMV4z77HLEkZabIQEImdDFx6lWugsNcT9aZ8QMq3i6rP99AU5o
LmXcp4+UQ+IGyalSxwjsa9gWs9UTc5teIxdV8IHCVYLq6nw95XWQ1+rLyqrE+C71
ocRiiOnDDhhlNbU4TOfqsLWVmcMSyuCodwl8ELbnFynNf8CzeSMhM+o98byNT26h
uH6eobmbSqEHcGkoLI0HD7wxw/H/MkGxtjLQQpau5quZ7hHujdSBlG77/hkCRhnZ
ALkTWgU85QQ4U3Q+LDYIrr26D40/QM8NevkF2WKmE+P3/7v56EMVjU+9G3zrjl1t
VQI2akcDlHe7ZGe89dbwudLmExNxhmfFlNay9w5k169VmJAHQAHABe0p/AaGv8Ji
/CjeCPcgbQ622ygJkYkOh0k8r5DiP+PGyGLY0hQmMYITjqMaUoG/pACs0KIHDLv7
UpEPXgs7klt1F6s2dvOY2trgj4ZloNxcFgsIHelC+kpre1mNRFlopNznsGoN2V75
VBG5N0BwNiq2pv3lo1QxVhmbNMme+xpTf8abhJi7Z3OmKqm+kKlekusQ9WWW//2q
t8SEUQSICC6Le09qvwTSqpzva7F5rqz1FGuN8P+5DCPB8vZmeYeickZPq6QBbOB3
SbdauOS/H/qS+9LUPZuQE/l2RKF8r9Bzav0Ns60BX2gX8NEgYYhpVTYTrHr9bcm4
`protect END_PROTECTED
