`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hxREFxqb7W5R0SP+YyRbbB3uAU7Tk+s6iA+ncukMdwxKU0VaAgkwdUugIDf1N9aC
gl5gH4P+WUW2Ypy5mW+/tBKxE3nwE/JklBPD3Gh0H/iXXL3i1CsQ7Gfl0wGMy0mQ
jcdckHrCzNtQb0ktm0TjX96cDGsA7VOtXcaUhVJEp9gfl1UmWD4bpCoBURAv0fPF
oFZDwLmHXokFYppgSsQFYFWLvJySfh+3rmefUJVCkd7BDJBy1kD7fC1ZNVloc4/D
4IsEYojNHt4ZNjEhvKIm7GL17fr8/x+XHXXBXptYHqEl7y5en0MD1W/wQQcCpN68
aMjGJT0r1jxuA15jG93cgGoMhQ4YxtR+wX7D/7Ii8Vr9Zn4cT9iXGYkyvfGmRPk0
kSoYPimlFA6cGRBgE+zE2a+st7Pj4gaMWgwjwoso4092v0HZF1nzcRUXr7HNNiZi
hebid48Z7mk2JLzDodYMEJsIpeV52HkxPj5IHtUd4m3NL/GsqSIGvHjR8bS6EEzd
6a1VMzyBfXa44TbXf7A006NVzC150RbHp4HC2sIsdmIj7N4hxKKKgYNozAtMKAdJ
IzE0TJPlODZaoJackl0t9fQiat55wnua0TitDNoOOYDqGGuiQvJJPs4ux606hQ/L
Vk0B+i3g42g4StV+2P8ZCMr93Jw+gezzlZeXRcvIe8IVlKRxOvHGxuOXsppGrBqP
1q4tEGnvKMSfzCwF8D63TU+hNd1QEgFEex87ezb7kNJwTxZ/IXiKIKDMuLpSBZd9
HZfbIQ5uTMV3Hb7l9j5OYs9McQQsqNF0LeoK5fKqZE3rCrRGEUUA5YDXyBZofYP3
nwJrSm+4EpDg2HFy7nPafWPT4Beo2cDpmBpaVn8IiX1FGDqJWF0D3MUxIWULamqE
E7L/7A4gAU8VH/WDNXuBF+Tx6SQv4qTM7MEiSMZ9DsCfkd23s3JUQnqvfNImUuYS
0GgVGXLAWl2DOku8WIpvIvPfIx8aa8xiM5kKts/h7GFA6yOfqtLQTOXLMO2m8icr
h3F6oZT4jEVGs9qr1R7qSLcud+xeGVYGNGnKSaIpva4s5sWIA9vASFSg8xTBAVQG
onO6HiOPzsFipoj1ctHm98V9pBqrKVJtkjFxh+sPctb03w5MDeLuc5UiqBgnAP1k
3kruhIRGfC0cp9MBQlkDnN4k1sED7IOKzrJiwpsXiGz19Ck3QApZGZDZQ9KvqSy5
4FBHBBYuL7xWIC4lnyp+pdwMGEJJJi8d1IBCrHzJr30QBozK4m3qVmc2XbfKa0IT
mX3T+8a292lnsTXpeLVRq8dKKYgANZlVwQgC1q7XdG0MvcZ/aSbGURRg8AiuUDmW
B1XHKBk3FFJE1lo5MAdGO59P/CrWo1shl2HosYaogEShWfYfHVsVBEVtrTD6bWIr
2eTBpavnMCkMEZ/D0EDKb3H4s5ghGs65UmCDXCtupROB976OzRRsQD8jI2zCy8Sk
n2OhNrEtxVK7LAgY27EKE/5n03yumwIAWKpruCgWp1Obz3/AcB3zUnu/ohpV0hIm
Qgc9bzkhBSroRB03t+w2aCsHAimoetmAeVEWp7iZxmtm5imda89484WdzZH/CL/u
TiaTiG+qO2cAq3oycojBW70RzO8G7okK8sHvvDX1sc0X1ql0nCU2l0z4f4wViTRv
uBXZeer7wB5fqQkjanCYv7p8yeGS7uFz9GIMuuUeijpeQLn8A0DR5qmhyl3kaWAY
S2ngRC6oZXrFacjdklZ+JoLHMSjo6vt9TPbSFd1jB9J0UWSPT+w1/oUqQ5mVYt5O
+txpDebonsUP1JEgwpSdvUg0qOJL5bmSKjsqHoPoawFS3Rqe/ix8eoicBLtRZfRW
akp+vLMorBVIqHpTAj5R23f/ooDP7y/IZwV4bpTkbHYonb9f+LUwl8DH9r5izW7Z
Lj3nSGbYBb+loR0WjSa+gA2sckx7oFOcyYyukQGPhyqcyM3/UFqNeRXHQOXUWeGc
WpT7M3aMBT0mhpNKFfsDSoT1n5Fd5Wj3SU7DejHm0LFzuj7NFtPXDT6ihey3FsSz
PErfrOBGPM3TueVX7XBC4ugeK32BstSrW3qvz/sgmccZ9eaDDdYXC39xcyE4ZSJT
LjI7Sa0VOqR2PowXfoCeNY3zLIijcDslER6tmm2J+KKUsH0ZF2J2pXZ2Zul0Rpko
LHmmdMkmKsTt/L4Jdb6UM27LZyONJ1FIH0AKqsAGHqzfHT2y2Dt05+3bRa3IDm/A
AD80b3g1yv3fDsSRMhN/GoVGdNiP/q8ZGaA4mA69NHNGEW4CRuznPloiunc3jWEG
/vAlmNGl0/U38FvfyODs1J9CmyEAx7HuR2/OjIftUyftKkBSz9/dx0HFK/+CbjgX
7DAbpNf+E72CQzX8Q6q44T33pzS25moMwBL2iGKJswZ+FKz3DJkRE27T490H1Z0f
GZlOmFPlM2wiVddv3tFIBLMWx3rDnUq9LkylDsn+iSUyoJJy0R1JHISjHyqKkvJx
YGu8DIg0BGEeScJvcv514GGXLNIZ+u0r92enZ5NQnXQrl+KR3fPFKPj7vUYiWKtz
5TG2qg7d7dgHoHhGahgOIM7HBq8H1lYC90clGfTDlgo+J/KU0eklHM1VepBCnEga
6YYgANSE30S8K/xTd9HiHJRMg6OPVyuR5nQn6StZfT1E3so9+fzAM8ETmwWc8FGf
d+VkBRksJ9YPq8jj7aB5exmKaO+qcYPEA6ikjknY5rA82jID9rlrx78v8/CnDXS+
yHJBRNllHSHKyzzxSJdX8Y4IP98c5NK6myVeY3Ikh7uGBvM3lmiMJImBgpTCUjcW
82xGlyJ6F19fF+TY0nUH+OB+IQv2pEh1g0MvwV+O4/xyKaCnFxvgZCjZMeHgeBx0
lFB4mCrxMN+8l01V3/QjwZkLL5mBgTCgzo5DFJ36VFG8z3yeD7zY//vdwYXfEVuT
Hj1wUN5jKDJYHfbNg9/hHWT3sXLo3K1o93ATte61YJl/jWN1dMdRxByjWRYKdrC0
Rbpswht+NGi9Og3TF1nOtZTYuoRg1X8t2l4zDBHAOWTZKWWpMiAiPcuiBs2aH23h
IxwqI8BgDVFOXOSHJ0ceOE5+VIIl4ii6gqVZrHg3p8Y1HQGpg8LKUo1TTaLg47ZW
9LAVR6AGqw1kqKzsJA8D7xn64dMxcasU/a78FxKWYEnxQFxu7rkmfSY2ydYEBeCq
ksHfBPLm6+iIFTB0nQKCZlh/4nyN9wLBczwSPfrMzcEcyHm6zVdjPOrnp/CgXCxy
RadvJC0nOs2SGkxb0QqNHg+mlqyOA6+05bLEIbWpJNtrrCQHTpjw0y1PIrpeN5zW
0A74wkVmLhCquIWoFzSEDxJkrmC7N+Hpm+q9VPiG7Uan/Zj1Joy8OJisnOLGu0dS
XQtFBd9Xa96EboVy1t7l2kkK9GsLAqenLimT2I6DuWYOx/KngVCac6fJO429qRC2
lwmaTMrNVeFFeafOrwEhVozaVb+r93irC3fC+uTvVlxWkACGesDrxTUW4r+zmCBO
1m6CLEWZT5wpr436jX8Sy1aKzMicUG/cUOKeELGHWI9YTb0cdJ63eat8Rquo2Bxy
kXJ4Z/Sy9FHVo53thTPLeynfENx7332qt1/b5X04iNlVAlkooZOGsKyYW8ziG+HG
GBh0k+Xtmeg8jIInDfy/vNPlX9Rdzvh7YgRrLEnt4d01IqMcRQWxezcZigqiGBXK
V+h71qq3r7rKJVzOVEWtSCoRjBnf1Aq3gAMzbj4x3y2LL7Klj7UzxWAlZZra/9+2
CJpq4WnDfvIjpi8vmSvd5AQcDXmlGI2UJIOVBMM4nf0WgYBbzEBYX1s69cdJ/l4p
KRCPmTT34BFyoFvkfbbFA+Qbrm8YTLVWiod+i5Jz/+X44/UWhAVJ31/JoS6k9RVS
6k13z/lMyhNHh9hy6qFfehIHS2k8xkRQKX0HgXdS0Va6ptFtKITs/p8Mt6jxxRfg
P3vzarD9kJCU/RJ74xru7IbA3tgc6dP92J3uo1Ub0SCc13dE1fRAnvrXvPOf1sQY
edQw6Ql9/9TbidhtlOWYnp4/dD39ABpOP49Zfj87taYH3vrA4ORvB0oZag303U7V
oce2df8kfrkNO9dexvoGZRJUWwm/CqI/7kH9IQy/gE6s4aKFvdT6JEIgQiPGCFHZ
sG5mebJ3iayh0jNBvTNVQN2+YfyF4FIHmrgJRlAL8Hpkc6cF+A0wJV2XiCg+f6u4
C74BBWwMeJQADfZ/3rywP+remYv4cfYAtS8AJOsW7zj4wVeCqQohS+0SO6UzZTh2
b7eXjTsZLD5DTbRZco53XG8fVJIyxlUNJ+xmzxb7M3uvhghKxXLxBERTeL4s5OSg
yxYbgHtq+7VHbJbySM8/xJP0XPLmi4Hmd64yud1gfLSIdhtdDE+B8af42xUYR5Rr
gL9bwZHm+zMRvts5KRcXBGyiiAZCIIn3mT8cJ5xE0J46w4fYGHHRROCQX5rUDUaX
d8RSwbnbcaAOEVO1wtBP7qvTqUo+NMPvQRe9g6UflaMgU+WaBMnVQRfuQYRz+kEZ
6iKK/6sExlTXvkSKB1J6K/1GCIHZxcLuV82q4IL4CC6CPlNKLzgoeoaY7NhAQGq4
ihWLGhGMPjMeZ2r/L4VTqPGqCRNSkdU82CQ8NCoUm1rgUxEBuGnRE20zj7SpHjBF
vyhvUi/sn4ez9xyEFNHEPX0hfYMF51/rSNFz6ZmFZd5M8PgevMmi8ROWAaf2BGiv
+/z4d+iE4eHSjh0+DbVkxVfx1nBTrAxYE9ZPBXHbP26HHNnrU/lCYb3iRm5qa/VU
lL5mBLeS3ywIQAXtBxnevjWkdBgdrsxPmaC8IjasUuyGFxeiLOLcwvQloaAshuci
JilbYCCNN5TRLb+bUoWGE9sl6WdwWWNMhFzGU7rEy83VmYuFNwb6TSSQs4luCRBh
RND2f7S2pamvpGbIvEzDor2K15BizfGq8UKlGYFUq4csec7FlqRHgV1hllCs4eZ0
7NG9miw7DsDkJqyqauXDlz2oK5rjUQybY6YHCj0uCfSLIAPOwm4YXa8vmaXyq4s3
M7dUK7QtcI9KONF5/LcPZagkXG2t6gD0JERlJjweoKyg/0x3ufO14NA+7hzZzgG6
dW1IDmj0cw8BucSI4gzibgQn6pDd015ohV8C0frbQiY8jofcfA9kB9zqU0cn3sPu
zl8QG1hUPfGTX3ZGhkEr7/aFoO81HXKwofB/xPisMsy+X58dFzcZz77r5g1vEcpd
UOUj3zUVDGFhn6rEtvcxBjPJMFkBDiFLYnbHXPDnzF85oQLglZiW/cyAjKcN2CcM
`protect END_PROTECTED
