`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5hQT/T1kxDXDDoITbelM24GV2RIEsI3tKW2t+m0EJv1x2ukpH9Bg7cC7eq8D18D8
Qjj68Z5i+qbCd9WTomnHph5Te9+PoOQtr+eL3BOJNGgZxiKQ9oBppRCh3kBqNsHp
GEevWW7c8sJr6NltplFg3tt7f2d1zUZYdAR5iM5jzV12LgtQUs4U2/xQH/dXwn6O
sa5iM3xzKwM4Hdptlne7125wExBUSHpEbnXFPpbE7EbRTMShHCZoyudcsqRM0Heg
qltDB1BeOGlid7u7EE5NgLTvoXXty+hF5ZGFCYTFpcjviXfwM9aMaQJrrH0hfNib
V/0Y5nJT67Heay55qvuq2sBpBPx5bxu5N6obA6xNKJP2s+dvwx/R0/UxSl6Am6/+
/4/oS47+XCy3DGBJqj7NsdCk9pcBWwivI8QqE1zlyEg=
`protect END_PROTECTED
