`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yj8kGt8a/vFsohutpOF+6Jl1HBL8Sjo4awqz9Tekr+DqbbuGLYTbINK2AtWlocVe
NufLRISLQMd8xRLoXIzm+M2J/ODHg3DwG3EKRcfNCQkRDGDWBKjZQ2Jt0X3jedht
EatXeLOaPr2P7B6tU1onoz2KbwtuoOtmnU1g8nHt+T5HDSXiZ4xdIBgonkqoLi3k
V4xonI5ybOaxKB+lILkzq4akEoEX/bkCwCquHG8WHH8KDkpaNgrF0GFRmzJcULAu
L60/PyQ8CFw+MMWF1cK7XkwmcVCqUoEwU7ROe7gIRwk=
`protect END_PROTECTED
