`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
25lbSwSRWeCnrPv1+aj1dqJNVvvq7vnTsF/xB6Yk/xfkfQPpk7kH11OLF0iGK2K0
ffAbQszUVhea8JMrmxQ66hjfbu1lJrcvMXb+ma1eIWX1PUwu8yYChK/WFfGsCJMh
MqFn4AuHXI1hgGSfNSJvPhq3liqGdXYTkJVBNZbAOm2rGj4Kii9ko3RXqvU/PM9d
0aHeeZdiIOoZZrHBEWzd5bNiT2T2Dn3PK8ysX4Z/xq8D4HZpBBpUpTFdpXkie8v0
7IrEWyBsK4eCNIv9S1wJLl8CrnUZzxceBbJ+BA3QP8n4kNk5F7jDNENTV+mqjd0V
m9NDvyD9GLI+7H/wZwm2CDpy3HVCaWzq3tpFuNOwOBtl58Kl6x1Jhl2BkBHN4Kd8
skmqLNzGZLc8Qa0D+YKMxA==
`protect END_PROTECTED
