`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9X6wWUVtymKCnLXAtWdLMSUt+7jdUn2x0a7/rO4ahHcE/BYUJpFD7+y0sX6WVFuW
3xI845l+RnuaBtxsOtsRc9tjv6zCHX3iokE5CwVaILJR/Yor2PTl4NvSXkUvXRhG
feYpHC3PATQ+ZVfcX+XJcuR5l4nHAiXKdWcMrXDrM4/QTFVtiQmJh+W8zLItANnZ
C3XG1TLQY2Hep+OooePd97YRgDMovNqIQWzkikKUO4rBPIZPpOs1Gk/VqOvZYjdD
MJRu5rz+oSoXecq5UYf0+hxk/ZcnKiBC27obfjFS45+D5DujrNoOhJR1SOOmj9uI
DzW42Q/3KYOe7u4WgIpfvDhiQpwTd3h3ispgv5kb80UwhCJ8k/a01/BgftAASgjQ
SNlhXylJoH4fW5yov3Vs18M8sRz6jdJuxAzSY2SCuSY=
`protect END_PROTECTED
