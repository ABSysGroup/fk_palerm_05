`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T8LpUM9lnwaZtsgdu1OrMQCEAckJidpKZB1fL3X/42CxP48NoUSDhl/Fp1oDZ5Cs
wHMEBB0dbp7uciG+jNYgH3r1LXVNURCpvbfGHNgWpH+c68I1LOh1ezo7ai9ysjpT
dEoOsvl9DqJO3EtvEy6vDQ+4gPPSJ3z2tWiDwFgqGqwCWqMqxmNsZltPTBgWCA9X
sfn7W2WYsgIjgxCCjjnGNs3mzgx7VhkPpfos83IquU/SbzefEYxxfr0d5lz8g0Zu
pQVfy+ByCl07AtCQy/UB6P8m0GBFDEhsaIBOa74dCiPPacH6zD3hbmmdqkjHyXJc
/xXO8+kl4ZgFovYjXrJPt0jDUqOB7aDjKWQh9gG+bUancPRQitlbprkaqrCiTXEx
K8vaVUsWUOld3cgMySbOha7ACwVQCyzK7Pl1IEGEd4WWx1B8TWipwKzdZgkgfIkZ
BZuSKjOFX3suGfwnUDfobnW7/dmrMmTFAZY2XA9c01fAXRFSJ0ZCxkdG94fYYQqz
orHSe1Lwfl0AeQr/FPEFEfJJ0dJTJ0FpqabBTl00d/u0dwY09vAm4V1tuIgxmPJ5
`protect END_PROTECTED
