`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VJECWnis3k+WoU1dyfvajsTzd7Y9mpry+yDfnWgFjhCsAphpVW0VWG30Re/V7t+9
LE5rJsZfOaBYYyYl868sKLyH8FDAhk93c749y2WTuDG7xJY8fR1sH1skSBcKfBNd
iY5sjSUYj5Ud63MlRoR9q7K5zjrda6gM5m9s1QoVgntq2mb3ys/KoGRTj/Jwe07F
+X7oTt6AmUtPl2eidWY/QuKYHIVdq3oNXfN2TE6tY0wks6p7JqP4dipA9ka1uJvT
xy2DJZW6QKn746NajG5hf2pkmldWlK/bVM7O/7USljJLPL6ZHoTX5sMt89XIZ7n1
EZge3zfgfQ42AENP/HJCiH8JWRaXOB0/i3xHLY/EQe3AdklWRCihiV1eG7MhIeN1
p6YzsAvPa3ST6Rth/ZHP0c/XvzvhL0/qsFZw1tSnJryOmeb7Tac6SvKad99PoH4e
dwBVXi4fMQQUOFe7EiVS84J8fyl6xEtkE9BVeGAtC4WX1lYlMfnzT2+6I9kZE+3T
7Z8ZwPBcZGF2p0LL2QfglhHNTH8sDU6ex3xZYb9YUEAY2MFttorgVXSgVC4dSgAL
mlEcem2IPHnmme7Y1tfGRV3yrgNCaxxlcKrOjdk8kdzzRi4LCyaYKgAhpmvA6nbV
0VbyVrZJcLRmhxQ2CffAo/pHvDKUEhfm3bOqkOB9fu2K7/4WsAEFoOwnpkCGPvVu
Sb/Fk/q1Gm1LCorapWZfdVu3tZYluHuaRVO65Z47g/Xih5H+ITiKSUXFG3scL3FT
A0HBbbrujsCOpxU5yr4UWmMxJw1P0qupGeoMn7Azj0Ebh6EJot98iCmQT6C627uo
hTNmBpTUMAzzx7MyvVMVKniYQ5gfRfDsxDHDsXHc2tE=
`protect END_PROTECTED
