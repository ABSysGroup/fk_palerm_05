`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jduesiiqag8g7QrvTmQ1r2L2hPv9E7KkDBFiien/fi2LzdxUQljgl1Qrz2dik4fu
ulrVPTfe9TY0WRBdtm06xplRQReg36vmW7DAi4bV2DNS9mUUaxMjMZCLNl/6fCMq
24UiBOorRQ+pdGNKVmRms6bercR4KwvO4WCnc88pscRY/6Du6eclhZoRr1tcBJw0
bjMYVjW6ij/P7RuRz13ZBWf3hHSyQFigHeghUtJJVe+TaQAL08gce5oB02pVE7cH
b2J2Yzplwomq7okOap37LiuDYfqFmaml6CA6rR2OH6pbec+vY3KCtyim5HbLK1Nc
Hb6VXKg3eeCPNH1IWyJsPDLXLHWJg2WgIiMEreuelU4r6xmv8VlXIQOOHMlV+GnQ
`protect END_PROTECTED
