`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZUx9rM0jtdPgcoe1avbLBb/r6FnEkWEFMIOJ9hvNSOsxV1Jsq/fiZBxYcanozYSr
nHFK6JW00jTbjaVgY8fhLJpUvcJeAlMDg1rjuMnQiWqd4iuQ9W8Arj8SsgkafPOF
1sfXMRbJ0weT0pPzo5KfqOxy/iTQw05JtSLDTH/tFdmJMMDPHY0HqnEacF1h92MJ
xxYlgDippvwKfVratgdOG1bB6uO+BTSfz8QY82blNPUJGBCo5FMQRfwDSmTf2t65
uHjzA5WQ/3ZXqNl4UdJ4xQ==
`protect END_PROTECTED
