`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RjAXfrBmrqJKdNYC+OpFFNAlhdQ55BifQzkQihHMdy+LTtEOnBEuncNm5NRlDIiZ
/a+At6C7vwB/Z4wC8jxNVTCbi2g+vDmgW/dnY7CptQo1JMgZbPP3bSc4BAIQ480V
tmdhZRCNVyUUlPIzRo22q1oAiGijn/JqmVm5pnDrTX8+IddgzbMxIt9cb8Gw0VoJ
IKb+Q5HKriI17T8hiszvL+IJbNNiXTAe3G5EoPFzDPIOGvjSa1dmJx6+EHIsXUeh
2OdbUp5g8R7mA8dDGN1gg3OhRDGsMgR81r27/KQofEHiMaRXH+KundQW97/f68Ki
/sLLvJUjkRL/PCiGkLNp4g==
`protect END_PROTECTED
