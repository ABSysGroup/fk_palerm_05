`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hove+/cK2m6Ku2HbbWQacPNVR6tXHe4w9sAB5VpUhtbQti4jKnBy2WyqaMUrk/Pz
U2UL+9FWRWthcpBusv6+y4ushqEbkNO9oTk7xRb2v9PovE/L1iH1XFjlFtLWFsC2
13skFusr5VpZJ03Mejks+rXHj1wSD4EgqUsign3t7cU1jES0q1qhKuElKu1qAmrY
yNqR2TQ9QYWCRtmrauQdpRtC7+Rne5aHwSKEP+d1EY+fdTTAgyG58Hv9fDdAPncH
iZxN+BDDiwPp5azJXi4AIFQSQRVoHKVJE5wwtEnA6Tg3u7LlXnzeGuRU3JgsbS9r
JuXuocSNaEhPMA5CzA1Plr0dDniNZ6pnC1QSJ3IH9oVp1K4U5EJzhxCiOgrujhrp
EIr8CEgro+on5YiLKsjpNVGG5EUa/GEAyQUZMYSyRTKhFnguiAfGVFbUL/191fiL
9FmJdNH9A8Asz3dgKwjeCUz8CLi8+zaWmd6n2ttqvl65oyor7mkp9ZfKYAnw1ukz
UX+s8kNCMENFvSSngXTDgblw2ZB0Ms6nFJKp1AaMuT4G/vT7Pn9EOg2BPb8aYUXQ
tU1FSqOJJyT7VgA6FrgzHYwM2hOAorDTqXAfeonXDre8yRTG0F4OKrs/sQV3xl4M
RkDvUUikhydAuHL7GutwUVNBlPN+XzbUHINurBZD+I1DTpngadRFHVH6VLYIcb+w
zf7a+3dc7q148tC3KJ0XNeGVWSSpwZRQJVmgS/IVj+c0vzW4TLLGqHG37l37KmTF
Yc6EarPp3qp3lQaOZS1V6Psj3DVElp0PKV7Oufh6v77smBf1NBf4wdjFWGdrew6i
wGb8k54yltqrJsa4YsYD7MhdLr1Xd7hZijmKdACyaZHo1JLR5L4rqSDY6C9HwTVE
e8MbRmlQSGhv2fLBNw0TW4ULQrXmoudx+dmE1MBCB6XmNe+oslJ2DgRWYyFjBF6Y
zk84MXQKZDqPFiFOnaleuafg/Kgh4vP31MWvhv0EqkxIxNgO8Gd+kcieAvK1sC9/
ZVtif/txwgiBjtKa9Yp2eEZ98+3RGiF1VAottbrx9ionK+CVBCyYAPOD+5R7tj6D
qzaLUauMXsp7ahp77vOqkyiAqWX/R9OY7KaL2rqhiv8m6ELwzNBbG27BQ9pIYueR
tkh4A2HeexQs3UeHbQMR/nBC0bdX1Mse+RwPfKILlraXN+0LJK2PNcuLlko2SpLk
nWESSZj9RD//zfq2MUdq0Vk1ZnsQ3sYjNckxlm9047JACCF0uQBXlTXnBXJbEgyl
itL3+6ENyrSSAkuUcaglV3CHvTrzDFuUdCT33aVVDMBhmEBqmlOmAAleN9INuoNo
xI+oiirDVQe88agYfuKquIOVaQRJpArUCjxZmYwaAkK9Fhos9vOMtJQNt6KJG2eT
C2206elefXkHHAeJIknwe9ebJIkOObzG53W94QnaxS1Lg/aY3bNA9K313GydhjAg
VTJtmJ/r4VRN4KhwhMvTqYbV5ABqs3HUqlmH50LpoKhU+w/xZw1xMaqPpftJ7VCC
+1tqiN+7Tp0ug5SOfwOroJP2kSccH0ZU0BaBnBCsWIPjTqCLZnZtbnIulzJDgSyT
aFLO/OtVK4nAL++y9tF3O4nIhBIFcCuITUNhUlCMMPwc0VPJiapln7TBSV3WTnsX
QxdgJw/gFL1pCV2J4RJxlpyzkcGWied0H13AvdFe14xAs6KT90vv7HAyXuKMnF/6
0qCuR2w9/B9EE6VBtKPeP9U6R1joOrrFnguNqWHb1AC1jAwmSVAA6qvHqCCdmjJk
uD2acRHXape57cO258/uHN54/TsU9o9eTKYa9PMA+YBpdSDFYNPFatXR0AH5fryk
Qc/RwSFOmclLmjizlG94th5NM6cjP2LxH3+BJ/0Iwes4PsPnTIFjaZOsN/0Sv9fc
suOTK/ojBCAa9SjPyBefbVEN1TEVG2OfLJmb+QZutf3vSUBhbgdsL4UPxd10sqyw
YTsvPr4IvRhYiEO4wMAyqrJn/iUEaC/4BkgaTNCEpHdxvK4xHXIYh19I81UwnScB
vGkVzPmbGl4JAIyU8n1p2ZvdXnjhpqbfB1eiTwtFusmDKY4SmpdHdsxb8SSF/lsR
M95MUHpFs8mcB0NLimRvTseELa/V/SlAeJ1iRIt6oFKUv09wRFOm1lnufHdDvkjd
h/aFpv5XmDHtDRNpi7AOO/EPDu4yEyfWJdkLXdBKIyPBP4I8pM2KBzeug8aPjOnl
jq5WvmLGv3ZvEOYwYCwp1EYVgtluPYvzMr1WvuOfbbtr3AAjzt2vvgAIkqdK3nwg
LT+1AMLTJJRpQB40zKLh27XacTXYhWk6nJy92TcuN28j6eg4Igb/XRPfDqodMoXe
0yDlCQZDH+9JznFJ563AfIQrFJmb8WlVKIuEF1CYRKcdAD4fRfHPlYi2/fJ/t55B
9KSJTOlX9qL/6Xh/rQ3y5IVR+Jdta9wUcVe3VuN/DavKKp+WEoImbNwTMG+1l9pK
uIpflY/hH6MPgiug1yVqhnv9o3T67e/aIahHVqhNo+hqc77ip/ITcAIUwEElpGZ1
vm1cEuRUVel4Dm5zCHLOC6NiXGvokv3leEaxIBtDuaGvX7ZFlKK7tnNj+X0JmHDc
demMZwGjSOzIM1EQ9UtTyiKF6VfFUT1j28NfNeg2lVATVRL3/CCugL8GaW8SnfXK
MHEsTL/CWiAVNR5R4lPgECPAAw0P2T7PZZOuMLCQFjjDx99yHpjJnlOFvB1+BJLN
lp2m9l2eMjiCePeaGuOUI4Dm/o92nrJ3jAg+CwJpsSQfIYG7oyZ9XggR/gN/eLbQ
1ep8AAv9F0HJ1997QbkibQi6/JKhqfmojbj27aM1glJu/Ix2gcIOGU7TaW79pBoG
Tl+G0hSyCNL41A6xgA4CDbFxMHGw6ASxbig/kgrUn1jdw5lBfMwZFaVh4E2pJcbX
pt45yTE2oePyaYIpR0fflbxh+KxU+QJ8c3Gi93RzphZDBeQiYOQikQuxMfPjz8qk
QUKBfd/U1mM/Ykef9TAjQD0aUTUKeoFX4rDwnArVL1seiShqscTOxSw84+sP7ZtU
pZAxueGJAJDQVVlLS8f9n+zJsWu3naOy80SVPRxQ3Tryfm4790H404wboCNJOAs4
VKbWIU8AdrwE+0a7ZhyxlXUEyF05qA+sF563FCuNwr03Zohn7oMl8k4Kl9WJFstI
CsOgQQCxBO/Zn4AWAbOjBEVvWgNeJ9w0Ix0iQS9Sln/QRgBjWwpFKXMj0+YlX3YP
CUkeaH54xCC0ouNQWUNQ4eYlssbs85n9sjDwyCCYxjkgpP+ny6wI3iHv57Tb0/MV
ZHFJzgn8mFx1xGW01cVxbpZmTor1pePUHDwls9oKeVeelp8lpUnRQLM3YOjHm9Yl
huMbt4JLq9XCc8ywQVnoW+DbX7bc8ZKNLtUrFKFhwN720h1P7FIIWiLXSjCTKMo4
+WhXaH8/4Re3C+kPCv//m1yFmiDsppnxHP2A9IS3gHv044UrjznyBy3ppti2RH8e
wWq1Eun74TdXULFGW6GfMKTPYclGtPrShu3tx7ybCrsFvf8RpQ14KHDz+J62snZy
OVh7fiNaLIKNB17m27wlitqKu8lnw+OSrhwvWuimlm0b6A/pL5R4GhpWyWyuiFvi
Z3gRTaQ1mXlxVuIzrGl2YOoPLwfbqPF/kzeCgHgZ5QaM3PXxD6FAJVclEX1/VmBR
vUxZqObKx/8c5Zq8LM/2UxqDPuizpo48I2FHuOg542y5FNajd/p/9zpIegEH5X7n
gk7opUJvZleP4jMfZ2jUCk2cn01G1MpHevEFdammvOaTPvNMQqph1eZYcBJya/XD
bWVumFSegnaCxXaobFG0gf8NOu+KwelGYxkWbpe8rJpqmSzwyH32eCC2IRfKk2ke
tkcuFtGqDoXsOLhdDKtw7ZDz3NHjRbfBjcOjNjdu4KNu9dM1q2zvaYn0yzepc1nq
wZklXw64Rpmd3q0sU+wgI/xFS3uZI69Z5QX80LNdhmKYPp58FPaSNCGkgFgQ30jO
aXHZNUZt9hYJnrgep7I2bFgu5ulqwBAg0jlpURX8pHGuyw9iT7qCJ6AFRkogbPvx
u6GwTJkfnIxr3rNHt6ZcytTLmmTTdHQe+lmECrOdqB62JXN/1z/BBtUWNcscmFJh
ltPJlCd2CcEudtJpjhSKO/BY5koKjzd3J3x0XQZBulJ8gz65ylCrMGCW7gfA4/2N
ZqQwaHK8r7A+yNq3BTguhl2QE+GNI2ROlSOIZ21aKRdVBqgVKXLKOBmXFm+I76Ib
ganl5eyWWefGzjtuMG2sPbKcLx54L80KiiglpAcuOH8s5g0ejM817BCbjo0B2H6w
aImMsQkKBEYzkyg6Wy86jAsxGhRR2Aafw7HryuXdQJcLxhHGaU8NPX/w1NMppq6v
CZtAA/l6oEseps1742SdceEI1WK91Dy6uOx7WGA8fcdq8+cZxEuIQcRNi+wCfwbY
fcqJU5EYac+AbibPCIvc7Y1Lz2ghDEaActVpCyc4viwte4j4hyA93cuHHtW3b8oQ
dSjyHAydte7xuUcPbVWq8jXppDkawKD8vek7Oz3pu8McVQJ3hlFhGBU0o7d0FMe3
/bR+FluMkuMXEEM4GlSL6ejLWg5W+8PNw1sbV8dJU2Sury15QKnVaUrhzJ3ttLJ8
S+NXgbhKlGeHb7XNosO7p2F8ruYCXdFUpxcAd32VfoZ3afiUj2KCC/xBV0+xQkpH
0+Ki3oa9rZgrYuSimteqxTI+etr+ApfrWXLgzsHT2xKn/b7Nmmf9ej4QJo6lj7gk
D/Fal1kshiYjfSom+u5CZh53v9Fzr/TYXWgl1WJY2vL8iKnRwFKRMoLMtb8RaJsu
rc/B2y241TSUKEf5kXYB4VDsYi0qGWccntoUoWjTKWPVZX+PgGkM1Gt4AbWfdrh+
HJSYpSJYZzvi2sho1pvUm/EwURFxuG+BhRx6akUMm7jXZ+icYdrych8btscEw9Va
RXrGGB73YGs2g+BCJad2/JmrlDJCtJFI4Eu0aYMtQn1DltpHWMFRupJmy0DMUDtS
0+KcdFH6pm5loXNYvnOpZc5yQhyE6ys1MIeFf9+RQQtNDG0BttnZIDYFeMcnaxtM
uhTd1Tp9HjHHcfjoNmeE9SJJ3p0FyWZCpB92mlF6f84MQyJ6GY2aE7gs0stGbCNF
PpIQgzjfkvpbNxL9D8FuBINYe7IV5lOhlktt/23PrLg4uvM1bj/WVoG1eRD8tWfK
VE81EbUHePe+xkW4wzDukwt/3a8R2QsRh5tocKRbefDKvhmiF1rqLYrGqmbuT6uV
yW7EHqxCEf/UnrW/nLI+JXbjNjYUV71wS/uIM1z3L7b2LkzJqwUbRCypbCGYaHYv
nJCWoX5MXqDYNUQKMmLcbHZwmNj8wSQDMQT1d8Rjwk/iW568EFlWBBBW+Xwclolk
pXDvV1sLFtsVfJX8N2BfkORB2gNgJGOSB9993zgePxa/uX9XSQ5zHerFfYA208L8
TKjfDeNpGNyf5n7LYLC4lXjH606idPPLNjLDERQdjDZgaMoW89WDGCF7d34nvCDy
lmsrvxmk1ag2M7waM1SRIP/eqOa6KoVKiOfPbARGTQXExNA5IQ1eabSfkWmWK2uy
xBmhJSh4cujEtOsh/Gsv/l03OibdDRF2YmbsQ2VZtDqV6ftkDGelAru6AX0mEqsF
iWF3JV0hjZeQjtnvTG0kvKFYpkA++w4dChS8HJKP0HaOxZ2zwB8jE9E19jTVYMQP
/WCFUzikuJ7jH684prUdCDQLur841jrR+lA15gRFjgtPAd9xy7NFRkEvdTgrTwyh
P+1YjvltU8pGLKH8ig2Qh8RvBDj25MYCMSlePgX6SBjk0ufn1VW76Oi2UUDVYYas
biQh9KN16DDWhtJOpW2wuJJVfiwVf6mAA1SRMcGzjNBQlPHClY0BHNEIcdxk2JaR
t71OBlkLi1wDCImcRH1J3X6qIGk0Jdd6HrCyqZhb5FZj+tTtbhO2Bqq2BBdfXzGo
4OVBotg4bMh5f+Kdqf75YPd7MuRp1yCeWavfhKj8zYd3tXDRwIhR1kMGB38yr8/N
1UrVNAR/v5Vhgoqdi8BQbnqdoYxHNlCZpmfl2SLIG5g9E2Ic8IwYP8GnZn180Zlo
i8Uy9vUB+lDddic3paa3avywUBM4GirNlG7ya/nYN3g9LNoW/qN7U6ixsQPIUdOb
T2L7torMqcomXbJfXU5oE7DU9jplivrzzSecwnI56cY3+YdFErnFoie/y2ttZ5p1
lXOgJmL8+lRC0qOfDlfda0cxMWzGjX2MD+kypa0goc9ORXZV3MsFWrYTQq1Gsrfg
k7BLSTH82ab1cNAsjM1mBTAWideRMhCiJWWn5FDax//AI2Slr4TdHw69bStjvcz7
uSlAeon7gFjD5vxrtwS0USt+ehla8xY9oMrownsIGFfqeaTS5SuCPxut7tCmljPM
XWc1LWo8PEWJ3Ct4fC4+mJzQgL7UibMxJkZLavkdJ6nm0kdR0Bmvn8s/5AjkE6XV
g0DsDuf9BQPTkwwei2QRZFhP1SbszK/6JRG22JjN6wAd7p3z8LE722t/Y6hFN6tz
JcTOTYxW2Gwg4Od8P9/6Aw/trbhu+ggzaGOm5on3+YMXHZQMKq2jdKYUCR7W4t1F
y+qq0KDH+yxAT6STIMj3FAWqidPq1xokd5mQ50H1IFpRBmOcHYUqXpdL8Au8opgh
u+zlsjg49AtUDnPie6K0LARxi0mBJHg+f/T4KaAgQP5gxGIcG/rdgXDW6y618ukT
kI6cpJtlU9bXSW1Hxwpwm+f0p6TzGu6MD7U5z+X918P4Ruw4x1aE2HIcc6S/8xCK
A76YCjPxYNTtlPYpqQkYLstfwm8wCgTqY2eIxlvNpw/WS7OFG7RZrdLn8rSsTgC4
soChnvi6+0XyBslefkm9rZgxCO4194xzXI1k+8rawA6v9AjadVmqkAavtzo6IR9m
tLDrnasucsyclIA7hypN+634FKkY/gI1bMK1vPUHg1FAivIxbGbYPdzKgb1wYhvO
zq/EAtJ4Qo4mzD9B2W0syjWLhaWSxYGt4sNYkXU5VuVhob1ySqDnhsAGjFK4myeq
3/T5iCbAAGkAEBz+Pnhh2LJGCsL9oCPOfcopHWjG7pbhxQtXGiJ09XNfKyPzCp62
XX/gXDzgoOKVLENxpjdHJMpZmhYW+G0n2eDp8+yH5V34lgL+4/4CxxGrhPkU7/pJ
E6UyiGa3tPfeqEQfynL5XMmpxc4XvJI479Slo3Yly7jsv1Fw+V88SYotDWcMDxyK
MKWJ45vtyyX1pwUgZQUqAPGPnRGlh9xuC+TqydYW2k60lRS2VnDxcL+VRcM1Y6BE
CCH26lCWGWO4NQWZyP6llwF49CJvw7TPXn5zWiC1Nc+72Wcf6+VdHRrqF8xUzwuk
/nwVhxgw8Lq/9nTbCFf0UpuLplGJqSkL3S5hdVwXXtBR9ixlUTSMvLF2ae6MFIn0
bNZdQnLqvhL+MO3BbqJzn5GE7jjoXP53JNjAquG+WG3Y5xDG5YZJZKaGPcJqlQwJ
+9YKidgnztGZv4qSQQ/1D3TWQCYMTnbWO7FcUzDEyTRoUeMMZnvSFIb3/g7F6vox
NGh+ajpEfjDWqX5EMCfCGfHEuxTSvMutm1wTKegesn8F0/lrhvLBibZcjKtGW6CB
w51uACfwib1Aa8SDjUGGQyN65uvmAwZQWffExuVFINMiBJCrm93BgZvimsRD35Iv
TJz45UVZg1WXqT2msxFHOmzqw5HMUrhDQfMdPPyJmAWFUxvjE0HBKsFKzUgWt3Kj
BxQuwsZiCi4gj0CqQ8f3YrtCT6tek/JENxwLOtPBnUDD+8OjSRJKG6FYjjn5ZJ/H
TVGPR01reiMxMvvh3vwZmBqjwQiIztajUn2ut+/2lgANNz2KQtaBjwjKXtvtNFK2
LD69SaAdGQrr7uq/iN6jflLplJia68yon0+5mu9KvKeB/w1mPuNiFMKOP7Himxw/
kwJuaTP+kUyNiRlbz46uwnswAEETn4tlJMReMRXAP2cV3+XJkBsk3X1i1/dgMXzd
1ejk7JOByuJBHxC3oE2TdsyoV16AoKfqC//HyDE0W2IYgUm/tYXpbPeKGY2QEMTx
9ZmDAj0fZmBeFsaVTvU4taOFKGRum8cWL5ccCgxh2iAEpaPjLhLRtmJbIL2MN1eU
igjrysAL9W8HGWnEw8jVwj+/MjcCWdJ6Ka2VD1gT9vbnsgA/keFuOFcvFfdGPSoA
yyoXZLFMSVkefms45i14cBmC5M1s2Fd8uAGbPP1Z6HMT9g+6t3+EtBQEbNxITSqt
I0klKiYFNMioiu3mxAK21NgQgzX7VATpzmGgjUHcY7iSxzj4lCRTZmLQAz9ihL8a
ey9XTFmedFcKQjVnqC3DIfL84ZlRm9D0RHbTtvzWGMmXTE4hwyeHkoHm4eI2KIE2
iucpsGNzIL4j0pV78FOMPInTEPCCyTREptkbIe/e5Xr3UMtLbaPcpntkyeyeFR4B
le8CqrpAPApkxyGGQVs1uU7DXgzH8l2x1HXYIsg1+I6qTxo7Slyg7S1shZH+f9Ox
FVDj9MUkrcK86qpxN9vkSlIWU9t2ZEcHZ1EO91m5GWUKYfWxaeWsLnAdf0L3YRGB
SrbHKJcBRZMvJJ4WoLkXEYzhFGQyqNYl9Br/3hIE5lc7J5SCpZn1AjXZPv5wR9wO
yhVypuVgwnh+oQeAt0Hj5RoPuZVkgCliZ4OOxbtnALsbxNV3rc7zd9xBdmTjTEk3
H99AQ5FJJPVNFLfW2rv5p1+hCsBG5AdDc01GKCwVg+n5Lvt4zRDVU8CTDyhAlln+
jafY5rJtvjzbNAKBfjZFtRvH/IkktnbJb0flBlphlQg+urDy8t6df/rE0/kAs2B9
SWH2KcC6zXFX4jMVbfsWug==
`protect END_PROTECTED
