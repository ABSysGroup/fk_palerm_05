`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UOg83LPr1BxSDv0wmAXi7KQC+zOxfm8EN5hJkd7CR7bGmsFKEp3zLCQGt0MPsynn
AFNuAG8k/b+eBQxGaPCoS6ivbtASVaqBxsBKPwUojTiRmkAd2ytknKJtEmHwgsn1
IR6crK+XeRUdJb/9/zA4tOgUuLYQM8nmGt+T9evRMSoZhxn+DQRJNMUi8Rn9+C+N
SjD1kpGPVvex8YKjXoFLVxccuK8GKYDFVXuwMnLY1qjq5gUh/fHhoB+qeglzm0o0
8FGfqV9Zj4ltftihLEKGog==
`protect END_PROTECTED
