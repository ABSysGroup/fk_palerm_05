`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k7acXoxgXDiA+SxHQlLo6n59sIGp5kf2ixIVU/CvQ5gOD6gm8hLCdHBICrqVXVRY
++PrCtASFCUar2bDbGNxcIbKix8l8htAQGho7jIJJ1503p70f5BF0CFHzUdWknSt
V5XF2gnb9rTelYzLmogbbex4pX7QbnE1Szd2edAP19eeuYlxpwF9OoQ/qKJCdWqx
ICrJWlyxP8TnWmJMpQ+xD181rzddZSkHpvz6bapgww45BKOxh8EqUAdpjo3HwKUo
XvQ1MkyCJPZxp4vVMFwpQupPH6iQPS/7J7piNzfLW5u0Ix3PBjYlmYXu0WBgSK6E
lSk/DtXwsPxPDtXix6FznDS5C8oILwXX8bBeZ6zX5OHJdvSK2OuLhnI3NLBPHEev
CEX9b2uN2q1vmi/9oveX6WKfKPm/E+no0Pg9yUpAm9fZEk69Uu5MONw3ho8dy3JF
Y2795j69R3P0TWc3sKZh6lewEEHP1QxHCnCIurqVmy3C3hGJ/rk6hIm45QGqOHCr
/XzLmaohyuicqtBWuX483HZJh5ARJxIcqCPIGqw36XvjdHT3PD8+Tp8hTiiNI9N0
sBWyBmmo9qJisENmBij43ateIfFG9qSv7E6X02jwm7hE3vVflCUTiwZA1izk7yYc
HKqG7bXd+Xguf/eVFnKM7wfId8zleXkQg8HBxotHnRI=
`protect END_PROTECTED
