`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R8CeRE9GC07Cw7ZFDQQ0cFhYXlLMMoZwdstRVbttRAhHSpNtIoTQ4TgxxIzEP2OV
Wjcr9Uhmokb0IL8CQR5Do/1CVpmmYZpj3GnZILuhVyp8qxdxZUbIDSjapalJZorU
JY6AvXdhXdGETUYuSNh1NNhZUBb4YTaPpVL8jwIRSENdwlMDSAHFQGycka9AGFDe
ilfG5A2JqIL7QrmmJNFnZKR7KQ+xVUyUyNb9uLFopPnzonVwemhVs8/sWu2l1p3c
pnh5K2ZK3ekZsdjoFz+c4rJEXd8ACOsDctTum2V4hFrenVTAD5WABY2VisvBsonJ
Yd6hwMnKWrTnSGnDZLITzt4pjw3+MNYe3RQ6pfdJRNA8T679zAUXOsubdJox/uu5
+iCnNoTd37tLOFCId6drB5AaK4PbqSxUhkR17CirOP00clsUStCeUHfqb0eX86Qr
/X7XVnHs7u4WnK/DgaolObyqZbyo0KsA6Kswq+R/uEXnemQPjrDS1BJE8ylOi8+J
6FRMTA6E0fNXIhtM8DD98DLDih/25VDMGppzTNJ3kHL6imD0FyWqSpXR9DA6GZ7+
0aHE9lHUTvzDPB/DYzl4DMmoQdFr1AQ5gKNttssEgu7Xfhr5vjQvMNM11cKLnwca
k9r+cbiaNWr7m9NHICC/7e+FMgomUNqjKYIkrbFJf70Wzlvi6XS2/jNoOsJHo3Xh
Eqo1uRepSujrAL4mesgih0fhAEGolX0M7wZ7FQAhV7oJjk+5oZabZIZsUsf5QKfo
KQL2NkGo0CjB9FVVO0cYBEFKINjzePpyYbPIKW89LATHo2th/cVud9ZcvEnPSCG3
L0TOLItZah71ZRMuwrvZntNn/Grssq5fWQlUQqhgnXJ6AcJwTBA9II5Aukq2A+Ep
/GMbFaBZGCTMEXCPkpaHDFScgjqaT9qq2ChBszXDLwmRg7EtQJFxKmkiC7xgAga8
TIXpZqgvlUZpzXIAKEh02AfZFSaI69C2AW8vudiS/cV2E4cHSRn4NcVKy6F93IEA
ZUjZEmBVX+n3ifBebBN01t6X2x5akGVe+N604vsuBrzI/AE4MhlyTCG869OUbMlu
zP+DKXN4GS2cVPmy/ubfw7RqJW7Qjp6ZrauZLoaca5I8fMmwkmKQxfwbCo3o2b5B
Gu5H12TxOrY4j1bGuAft+GBzPED9mDneftgJivm3TbLI5GxcUG2ph4eDcm0odsEs
E0dHI1UGBXmJfe6xwJA7foa+SRJpV48JnNiCyLt1dw49SqR/+fUm8KAeMzC4sDwh
GOVHTFshAI1F9tCgOXWAlBEin5sfr7FkUo1ecFRZ5iwiGeof3CCVnkBb06h8UKBJ
/oBINTO3Zcm68dQiAw5nOSBk/rb1RhOl0GXWbJUUK56u0PTUjwCc1F9PyARrTuqa
WO4/XIYnMIfXRI0kaFipAciib9HuHQ3NOWW/r6LSHwRSGtlF9eK/SYENKuOHSzpP
wdspSSASZ/6QnCMDhlUJhuQIZ6DoUAhDz3ovLNhA2qWQb24YbovrUjxIlEhvavWl
F/RZbTmpaeHL2UIuqwk2deIOO6UThTHwgTFPG/C7pqSwZNmDhfvUmX2qVObwbzFI
QbgntiiSe3AGIcOSuCpRvR8jGYJZT844v5XKiPi5tGC9kzHXe/avUyedGBgg7KAj
j9uTPFbUlcC8ukwO9a+PUswkCoMVAhCFhGnD84Dn3uVTvaGAGyvmTENxcUzqAzX9
h5bgzRgUnxmUqev5thEittDu9ea2Z+N/PlfjiSACWV7BDb0zgm46CFDgpb2WPLI+
QGNlU0cvdzXZ5hEae9A9cl3lJZAJZm4fq2wPAK+KlG63LGiZ0lMI+0v/aLFvPVyq
2U++ksCHD9FU/e3sx5aKiqSVXlJ+7INRDo0JHC0UiWxhkVVsZxdpDpwXnGClfo8D
9xKDyRrEEV/QYnG85WKuXmoPdhrhdrAkBrkhDUYnuBDKgHF2j9fhxdM8iUlEsjQc
Bwt8xUTKQUAZllGikqEdgypuO1wx5Ye+x8cd8Vx6lJSdq7oeKUOb4YuRpRFuaOz3
g4wyE+KQqHQTJsVeMRGqnMNYwzcEfV4nLClVUAqNexhbRbwnzJI02XvX015xemJ9
lIZyOwMEq91yXiqExTVFwF79tu5e9sUKpC7b0CYWXL+Yqn5zeBc3+oPEzidR0ea1
Q2Id4RgEd+fj0ODZ0FPWynPmfXuQmqgWiTlkkHf/Gc3/tAgIRRpOlxRWCBy18DJx
F7x9OzqgTlvytD4AXUI+fu47gGka5/rTRplAx7bdJN5T2PejsjPK/2Nq7nYY5YVd
lX8wMwIwZevE51psJRZ6RdHX6w/xgXhwk26sz0hWAS0ItYEfQdwSvmXFUkC3V1Da
zsEhWs3vyEeImuWpm2CPPro3u5T762Iapd16QtjPodDMx+Oa1W8II2szBbxYsku1
lG1xbH8hSE+iZQMXqW1pqlIwcODS93SZIQOCM4D++aOrsobGxcdUmOA956tdL3Ni
vSC+uoGee2KXTQ0OY69HIySJ+5jYT3xt5iFKS2NXaNX+0tv/X+jBS96PtQBNErOY
Yz6rQKkR44b00FEcVD7qX0urzmd/zTOPQ61B/JygFUvgwQLBqG0Oye6PKb5OEz1f
aThnSz/UxmMelLM7VyBNS5/AxMuMXcsMm74ESbS5TInVvMAB9crdqk2Y79Rc/N2a
T/O7F69ovLj30r44lya70vkwQ8oONZ/qxBkyRIAHSdbEbfOGV0iZUq0jlZcU1Blb
lcyUYVz9dLPDoUjuXIrK0VrqezjLwlDozOLDnDQpbvQl2OULgXxnCUMBHXjYimMl
q9UN/0uotjK9wC+ub3y/jzyPn39Ri5O2Vsug3U0dYWufX3FBY/AuegYjgHWS0r1X
ChRBxfdWuxQVngEU9Sos6//CQctR28iVnsUOJ/IMu+A9RtVmtLS82FSuu+qvAA/8
DE/ydmNrDkOx/YTy0CwEZcHSyc+UJG+IinGtOHtjEfsFl/G422JW1ezUxtZogTTk
kTKP81qXgSuypujlSHZfeztyMYrYjfvKjTYcQBhzKKoeogeQ/JY2nFgUA8J8Wwbm
7dra+U3KcGdcdbOcr53EYSEZ31yYXJ+EemLFF5aJamAofi45x626LbLwmnFngMub
GYkKwFIi12lOLpE9GNo/sz2yk438yUO+68gU0P3USz+ISsKK2FbrSZ2yB1kBTgAe
vbvKzSHWI7UT81d370tEbhCvSNTIZBKxa6Zhe7vOagRl0C+XKjdrqMMwaVxEDCSk
v/+25FCKKdclxTJo5G7CAx8NOYORkNNlxB1VanMbEkBx+2leDHjGoTPBBa4I32nt
STYqen9rZLnjUpaLRQkG4vf/JbiKzRVNksXhaObz0BH4kCSZEhrY9i0LDiiZbUhw
ij4/lShKlO05FQ3s49x6rOiFmmeRbxFS/66lrvfuogy56g/zfcBE/4fBRiFdB9SV
eLIOa+eLDdQUOWVwLO5o+Rc1IhCC5vytMP2Y3eLFkoAMRVpFBSw8RELlZa1QJyFp
eyEfSHIRxuwIyuo+FxvigDry/lYwrM63UwnfWdPUJrDpnDpgOscq34nyHtmYrBD2
SkzOg3Cs8QuHRkqRLYzQcmNzFaTvBvphjA0MNUP4HYj5C39bYOQqXAQzeWGiK7Mz
kS78W9WeuFG2OUjTOPR0Z2T5mYoz4Z/CAeAkYTpogEeOGMZBieY3j2MPtFNiTW3v
t87ydJxjGtQ1YJpXbhDvg1HsjfEVQ3dwRhypS+4sLBT6srBpMBvCgD/8BIyMjrvD
kDYpWSGUpeBtopUWhQVZZfjCsm6lxQi+ldhvkMrIGnMPk9xYMLO4xkmbWmDjRJRo
CxrUhISWfstcwA2LRWkM6qtvjWjwm/hZh2An34M19AtCoAdwDnp4qpAmEFgDTB1g
WGkzOTz+yJ1nnJ+IBYFjVW0vOAy+Dm0ha6iFWFgIFdHxTP0E+QmON9gRTsiZNdIr
ByKqTO6u8JP9lQAlAHmcudOAmtFw/326gp2M/mnlkHCv2371T4BrtE8pkckGVeFx
8SinIWMfhbcSqNdNo10DwlYIK/hwMVVA0PTUn7uEFCDHDpP8h9+gXb9PxWYb2aBK
Va8/GbXvz0Hw3qboPIt9zOwvf7MxjvZsk8FByqAp8LlR1UUjKgADgeTkenBr0IwN
V6yTEdYf8BMuOT3Pi/I416+v7Py1FT+/kPoylOE1DLmu8UuxDie/xqmeGTkPu6H5
yIaa1EHRj5ffE5VmABd5H7w4YtIgkeRaGngOKCqsadKBKSOzAx1fIf4N1YtuCT9s
fUBIynVGHhTYACsSPu+5pf71uLueEVcM9MbZdR6v+2Xd7YHKNZXNiJeiLGF8dS2z
wM6F3Ma5xSFpbEqf7rRhRDEnzUXBtPHWVFnGOAGjkHSREnaiKAi33zf0HTfXOszp
zTfozq/x0GzrLBHXcIPabNezE0czw8FIRXSA2mu6WlIYghW+YnqF8YYk/N54xe1b
KzUG++YDX/pqHOrrt4kbuPz9dv1EJkHDpnIyr2/w7S6uADV7x6U5YnsTMU5Z2ui5
pLGi7Infx3RB9wIeoBFCoxiPPY158WwpLrGGJRk8JVrLRkZR0hhaYXRWdpes4JCN
M4vvXYzOMtcKdiFhcXBbpVfQs+z5+1EYu501aVg0a3O7X8OtHsQJtyX8lRxFMZTl
QdShFuVGBmUrjVA3V8nw4rS2SdffBUXZ2QhOKHafytnF+OUDZq8RN/+bP7nwOj3/
OD7FHaFKFpCh/Kcd23tgZ+rV4NoOgw+HCRwC5Haeu/5b8wqnGHOiO6xAbayXe9Dg
JQOy6Ao5gggDveJnJG0kMuKbEV7mGcDWMTgCtDg9BtDFS8X/RlKejP1+77qIN2jC
1tSOdTdsf8ePWOVqnHpJPkB7GbwE7jdodvfh3L6dGTnDzNlLmhf+IeWorgiY9OR/
7wh8wAUTO6jhz6eHRDkeo/pH581VMYb8mXWVSJ+z/t9w7LxrwP7LlmkxoDAXAH5F
CuvSFwFdNvzdxsiCOwwGMUMVcRf0WS8ceGhc7NE83fw3Yh8+ZGgHDsoqEJgVkjQP
/nx4QxDdxamE8gH/BTfcphGLxGHH+j0oNVpPpwFg2S6xB28b8H84vbQhfy6imU05
4Dsyr6nJz95HcQm+PH6bjSkbHaC6ubgshCUgYwYckXpNfxSqdODzdn0P+6g7lhNN
5jNQqiDt6k5ynSkD3SPUIgS7s355DELl/wkdg41tSS9FXl6bZ2DIfpOxGC9vXjQh
W0peJN1Wc0vwy8YOWEEKFazyNU2VFq/KFArOJ8DrG0DF+eyAMtwzs+vq49j6BzFv
FF3SCP9QtFphlbwn6wQz2knBr3KdD3wz6nuQsd+0Cv4pruTZjc46PpLeKRPK1aDy
MqjNtXWz4c+uIFjnKzIvJvUZQbaTrU/jiqQx9rjfjus=
`protect END_PROTECTED
