`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BIZ3iGy5Sz39zifz7zPSzBU8MpLdhWEQQuderkkb9TYgpi2B0iXdPPmLnM2XAyrb
CiIIxr+nhFEIxvIEo9sXz4SOZnQ61Jq+BtK9jMl3fJXGAroNJiI7WRT0w5spUGjj
JQTsnRz0EDFyjSYeCT+Z/lxVm3LwLf5UGLuTCaDOloqVG8SxaiaHyuRbZDEPfBl5
NBsuDiKQAWo5e13dvJoTRFNj6YAb7g22CLFAaxnSW1JN0feIrLgd3i4Sd0ueOHF5
/UZvbWa2w/I0OXjwLtXVUOEkHb+PwvroHtEojBM/0xYEmkgU2fRaNy64yA+BLgaG
HNXdACaKAmvqjFjuPya80XGbVG+bgnCYccVMVOWg0MMBQbM/f3b0I7/y87bafXlw
yCIa4iM+g1Zu9J/Xn6QfamLI7rG1HQCFnjXz+OhvqYkxF5J3jDAMRR1j0CAouJqA
`protect END_PROTECTED
