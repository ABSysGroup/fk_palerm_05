`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vm4rAd2WXxqRW/iKHst0DZjYxH4if9zWj3SDakP779kyDy8FWN7y6rzCSIIqMxeK
EfWlOl77FCCuoBvCa4xJniHOAQ4Ft9InRecPQRe46rVQ3l8wAR330pnM5eQjO7fd
lsVtdrc8yQpL/rgb9WiNPm342//PfLGcE6e/oIBLshzdlwpuqN/cYex/2h7pIIkV
35su9CosHcD+pQ5XpX6qBy4SamJuuRDGDf4tbM6eK6S66CZQPpRfmE559XpGKF6A
J039HtmurAlrWwHvFGOafTlx49/K9VHHJKifxOK1HfaaRlQE1uosKFLq041wCqVB
m/SNEp8QGomh/r3LW/L2QqW0RzefGdzwwkAlELYzchDCyMnZL0IBxbATonnhtOkz
i4ihjVvb1Fz0emvZnzpq1ky2xZlhSQHjIzeKBYWN0w3+BlFXqFku5Jab5UrvLyyB
yx37kQFQeHLtO0hi5U6Xa3BmVLKfT/vxFvSg+K/y0i2ybGoR8p5unCYNeXpRYTjW
/Ow8DhK8j4E46PAmW25jU3n+cBvBoP696b7Asj/y/bCMrRSy8Xne3rbUJpNptoMG
XETfc3Ja9FzHjuDlUmk+zULI7vBrf4uMCuiRFR2U4q0=
`protect END_PROTECTED
