`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tDSce8edF5vnOLrHKkaDCLxD8f9hfvkW+jUOtsJhzhslW+9nQCZCJs7Z2UTtmcmQ
asTM5CaMRGBnfWV+ibMKvzLodjNufdhf1xkl5WjgmpbR8Dq15YEAw8XhGE4AMCkv
d/y7gSiEBijkoD2qPL6IyzL7iNqBA/Vs/A2L3f7d+9GuetVQXBICdEtnqS/m148j
I94wE/V7cMvc1zCy4vN+803zXr7BUleKtJQHC4GcNRy4MtQ+9QnwizHQt7TX4mH4
p2VdWE9/HyeuLFw2LNap/42ttUUMTdYJslukLSZbMIKOR8UHUcv4mW7IIwaPzZ+b
xXHDmotdBHzbYzKE53G9GHpK4IYvhnuQ3J23z8kEdks5ZDqbGLFT0Yib7/uj+aue
2wMslJ/aUlZ9xQ5Gqe3xE7eNSAW5HD+eSzWD2eqmGHo=
`protect END_PROTECTED
