`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
giyTvE6YO8GK/LSFtsFRLLyR+igPIIzagTIesnryjJKHrjj89nIbbmzDfpC198cM
ejkY5bEffmqstPeqEmXne0yK2YEcp7ioMjTuebOgL0YqmU8/bhDMyv9oaN3HmuyS
0gnx393M6+I8fiAzSC6Fe8ABICLknDiLUxIjA56m9uVz0gxetP1gDuPMgHj0Kerd
cPAtbzmU+i+W2T50H475M33v/lfVAHsNe7InoIaFphIZKL+agN8PWE5U1ixT4uef
cQ5l6ioqm+/60I4VXCl9pA==
`protect END_PROTECTED
