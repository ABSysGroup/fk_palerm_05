`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CjKR6oq3vs/GM5MljlYp6OXP915VlTWX7ZCy+65wN2g2pGcZ3EMPsMsSUb30nZ/K
GfOJwqis3IOty0EoYd+wdtzu1XIlB7wYrjrXDlLMTdBVE7F6Tf7fO2eVCVDzCIM1
uLVunZJSKp5h0s7TWVjfm74aaE7CWDFjduT5qyWPt1oRCwC8H1hIoHRJwHj/QjTK
BZ8sykwW9539hmO63APnNJtd31EWrzDeD06qD3KNRkI4BJPVGup+qgd4q6sB8Q00
hxzmgLAB+kxsku38CdwRJMesQjVRA1uomuhOwJoW9Wc=
`protect END_PROTECTED
