`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2MVxn+ry13h1IvBkPqzgHPfjSOvHAF3T2k60/DL0+X6OhFce7ogBCqL2mte/hLpN
3LeH6d7oDoyNsUixPXSn28r7WoNaTlCk1h9y+FXgQWLXoBK0QmwR1ttimKUZ+GjS
DI/rVrnniDN6LMjIjE0USuHK3zauEIXWxbUw1V0Py+qnuxt6nT8Fa39AfjuZmiox
C31a7nUfFM//v0+mSsjdxCwx1JvCsYF1TfhLLjnY4WBuDY6uphWyLI31/uldJtSd
j0X34sClowXi5Sc7IKVKwCSgh47tPKO7ELITOFWcWEZjke1FwJmWbxEbq/0H4Frq
YK028muTNkOWRwIjjBoSZA==
`protect END_PROTECTED
