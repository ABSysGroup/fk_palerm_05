`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wFg3TvNf+k8OhFEVTp2ZkY897d8XYWs8fWjnRnWM4b+tSOvoy0i9q4ucef0aifrg
L3JcJQS5c+XQvcf7kTQNtpYVT3y5dyq6tmDZgyq89IC677s9nC7dwfGiTc5EC+pg
27GeihnZuW6gv6YnsmMRfYs+lkZneFUbCgPGsUDdqOgBX2651UnO1BoyrrCr7HvE
y2ZmkGLlgdMRPN6aGr5VNPZg4xdHZQU92FjlxU0RZo40R+1kSOcrGN9mF/XfKa1Q
MbXXlCUA49XUEW9sv46PCmpeuitbWXz7uhg6axBEliUXyG5y8zvzTLJ3flP1Ikwk
lXi4+8Fw4WByprsJoQK5ljB+07OfjoOjWxpQbPQ3Bg+6iR1qkiCzShxLz+2wPfrp
FaD8NTP5DGX8/U0hFzHgqA==
`protect END_PROTECTED
