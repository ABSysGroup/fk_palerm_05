`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hePMMmFJlwVXi6ztmLEY+IaMMB6/DiRcvcTKz4dTCxz+UYI/1n1qL/zLADArdvro
NzYAlfvj9wv+2q/J2KQ57FahOAQVqknN4CfU6Dw86d+mKOnhEWMsbF6Ht+ZjFmn0
zjY7kGeIOgnRxeVreJqU/ssoqIr/5qX5IEL2IPpJpZZRUISA5D3t2LI1wG/Se4Ya
MPKwzLuEYazsIIRT9+SnHStUi4OYcJb890tuUWOOo1a7BsOXw2DAX//vIK6UZcsm
b5tEv4JFpOhGinVUDwAGNI1mSMJZvvX0k9/bmYwmCuEcLVb3X9zxL3+pXEK8Fuv+
a21RN3E8o8A0QU+1B4+PUdCZ8Z0sqe+JrPcTK73eLwWBs4GHBQkJOMuJh2jzVwzQ
L7q68Z0V6Opi7PccGDOpwxpxR4UEypqoxqbLRhc7CMRDY4GqzLLr8eaf1AGetaYn
3waHzK4edic9++0qELW0YHFHclt2v+DVQbOoQBMPYfNjfCIC20oTGSUTuHg1qmgj
12Nf1oswCI1AWRNck8x+XNFQNLCdp/wb+09X8XZPFWTLUQkdTQWBzoa/farZ6vPb
GRVBiRiiz8hH7ava0VeZddfMPEwYujZFklxHxAWQ44QbFbf5OWSdcO7G6MGFuNci
EXdSHNrZ8LAVHKZmrNJ0SzOYDOMG8jbqNzAmJlJRjdAqop6jImqK+wd9yMdyT0zs
uCXEKN+0ycLAJztuqWwESWK54zkZ5BIqMTy3rSOhiIMBK+k2tQ01AYNVpt5iR3zY
6pnZHRxg7nkH/rAAupmwhxJVaIwx5YRDXWHQK3ZPFrKDGONtkBuww+xKNqKOj20h
h3vpuFbZ8/rjL5l+dmFZaTMXsznEWTPzhFRoMknnzR3+Hnsi5a50fd2kvWv99/Oz
I4rgcPsNmTVZOZZPVSMUrRfzHdBC3kRdWXcGz6f5l93D8dQn3NS2hk64idZenmDU
`protect END_PROTECTED
