`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ghlcbpQ8bhhLyUwrz4+AL2lSAD5g9qdWe3f4q99EdEH5K6tguAfzMRDggE36iZJV
vBsC85420WVkKZyC++was04hgvR4pmnOVSW0Vvy6LyPyrU9AC2kk+Eb3XUMJUF5y
YEl437/B19ChsWIwkLrWhr8OMWwsdgHg76ooT8Q2h9OaTZ3VhIV+AozYpOR/j0B1
VCYXVmtENZj4Kv0nG1WZQaiyNCEdDz+UTYi7paCRgqk6ZfJc7+i6fWdoQA4IhlxL
Hz+HtXc1lSQ/tyczkiiKH8qUMFymLSNVB+kZxuRdix0al9fex21+NZfjBnmdJRwn
wEcywaDanFXpxWqAy7dd2PVBQL0gN43x8+R8hOjkbhwsvurQZtWFJjwFFX0NcF+w
mAimp7oXjpex3CmIGbJVnZui0ROi0r2LEgSlCjP1XnjKn34yjQi1gEFHApEg1skb
H0pmbrZgUA3LLlPMZ5ck2WcfdMLu1oAc2ycPRHKPRxt56M1/g06SX0kx6aO2fJ/G
5MXl9qb19xL2A68p2VL11RA6EDYq1v/MtiQyCEBERVLSjWGbfRCwlDyHPgrFeXDL
0os4RRErvWlllhtnU01vzWQp1JTgULrbmgxzg9USOeR1qoOxbDk8FLk4TUC9IJmi
dTze0hss5eN7bsUU1AlNGw==
`protect END_PROTECTED
