`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GeWHcJl6JtAP+Nyfnucb8fYvvP9+ZRKMRMLeUGCW3xMHLkYl7AkMVtkxwx6H5HG8
eE21EnHMlh2xgGCoCiYd+ZfebvqiY2aFyz1GpBs7cUVfuhsBwpjQXeZJB6j2/EHl
2OK36Gtpavva9Vc0cYl6/M7qqFqsgpyBuhVk97qWBifbpZWfEFM6sWLG3jlBIqHu
HN8cqBdq2RgXbd+ZKBhot/Qz3Ad73BObTMrP4LVjwSTU5jORhnD4T/Eo0IpRDzcl
Ih8jRFsBIbKR3rOWHpH2LBuJwur6pKhQVMuwffmrx3Aut9nN8n3mLMx+FZ9BFnd0
opq+C+8CfE2huOqWFkAkDf9C4lFFslLNcHas7FRpkVE53VeEQ1C2Z+RHvu+UJwsm
SS1IhcT9xvpfWJLd2ziugXxVVhWLUc8FLV8jLM3WTzzgWaEFe/r1HAyZcBxRFxV/
ILy9WLw/w395+tmrRy78VQ==
`protect END_PROTECTED
