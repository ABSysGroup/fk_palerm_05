`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hPDtdqu56rofd5qftDZoufHYK/jS90RodG755Tep+eSfhtpc/hwR+I+fF+z0qo2L
wxUtvKWLfLfI48Rr+DUxJkcXgVIHXQNGLSsbyxuO88fihYjM3ccsxuxPzuloZj/M
mcfHcnpW+YI1Qh7iwZ6XlrNCp9aRwsdxJEzu7UzuaUcs94SaJQaxm2kpO1+2SvuP
bTOOjTJnKaxG5F2IKjmclC7OoWiTA27WU8du+mIuLlsm3FgDGxeBKQrk7aEb6pBm
/T72/V4JbgkRaX2xkLqTQqfa82f28Bs/PUSEA4YlabCEDfk5FsZZ0HjvwdX8BIyx
uc0ACS2ZKvoMMY8+4MI9iK8ZxQ/T2Bm+ErX4qGfsMQTiV5LOc/ntKmSlrkCQJSwu
WKzt22vZs36YD4cZ/pWmSg0sEzOZIuWW1ezVqq0ap3WPRZIkwLmkQ9GIIj4tCWH7
AKY8HOObc/W4Q1goABba4NwvGRZ5VZH5NeDtrN7/DGkkEghp4CpeTAXOdq6MMRX+
id9e3gdocZ4nk51Y6MYJv2kXa2oL+cEGLKbDLdQQk8aiBA7JvChbtgjTdRYh+UP2
`protect END_PROTECTED
