`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sgqyf4c2ZPZh1QKTViXSoLbd4MVbTXJNFqmMLblm9jOGg6wbtAZG42XKFiNf7d9s
gAZs8mIewe8tjKwMJbBP/EEWQE5ZHljZa3W/rotdyjQMhYSdgLgPsuhh+gtfwOzC
H01lyPnQz4DJuRjI9lj5pYpSsZzijp/P5KGeNxjzGQX2QS42uWoXTI57gyvWOff3
puToqBWbFq01Zpg64lJkPB9E825OP6ZuID4wVT5V57CZ07kGcbDfPbL2w2hD2nh2
gwqLBkRNf2fz5bEq1TT5+GrNbWL7EJrHkLxBe2otzshMftX1TrAEFk8yP9u0y4IE
NTpsiD6S2bM6Fw00gQJ+WRRaXEUZWqWX6J6Qjww8yy8DtUJ0lCeAsC79a9DV67PZ
1/yLDSQqLBXSsQJnphzcFxrhSDnuD1x9CINFkIezPVFDv0asEVuoymkmsi9jcD6e
3jrE2Vtu/wrxLPkxM13ZMcChn6PRqQfWrtcmAGemZPqQ5V9/cGGXfJwxBUSBMD+W
3O0UJsk+nrrAzC/+ti5cj6nSQIwW07iUQMk4+ugw3eEIzJqgPxwjPH/euFZnzBkX
hIdhObqJ8HlFYuRqTKqBCxHS62DNmDPK2x8rgThUkdYg3DQLRPwLyFeV+wZI3cRY
vEzstTk2oTJJGr+ihkLFkVmszJ53UjAayeE9s1CRowDzOcB3vWQP4E0wns+WQKi8
wqU4P53JPttH1KKSymlPVnPsesRnQgUEtskNog6AS5EEsdh12HYbzMgF3bNelGBc
eb5SUiN4hbs6IUxdP8ie8LPgdQFOP1uLt8n/FQZxWJMGCJd+z+5dJcA5f63t7b/i
VzUg0PNGCu5OGupyNOeOx9VcoXYMLUavpVvJXueStN+iisixrBcs6W3bbN+6kDB+
CqHPwEuyw0ZSyrs7rVhKo4L0pcmPZk0KmLCF8RNWWl4FG2TCBtZWZbqzpdTzdNga
PHvqeBnSmUpTFqgnkxRGpdff+yOI7vMuTHyiRMwvQaALyouaNy4bY8gDp3nhbN2s
FMLlzqpIw+J6zUKe5rXyQRqGo8D8vt9UcBsvDS7T+Jn5ySc9fHeYGt4sSwsOGZGS
YhUTmxKrCfdI1uvYoqHwdv2dShQPmAbIL26WBd9+q6d1QL3l3bQrShUJK4dJSVwu
prp+C5w6f3O7ty0/H28ECYjUjgObVjCpQgWYOwhu9ID4q5RSRZFYubOXzrm/LW1f
BV3a4dMyY/xeB03Twz+psuZTWssJS2g4Xode2KDuDJxQq3rzq2Ouoow11GwIsT42
SLWn2JORhIAPKz5F5g9fp3FMGPby3xYbxD2JCUhPYYFOlPk4i3zvLRP4Igp9cmcm
+pfg7nMOeUJN5I+ERJ03wlhnJkcY7sE1yrEOIfdgkVXynLRWCX6OANBSi2fCNwPr
6elZ+2HzDx+0maW5Swq/CqGZqhzP54BxhKpYuQ+U72VFyKeIPpOLKaZNqugnrCVv
NRSUxDT1W+Xy6MXvRnQJdDcJbPvTXsqB6Jngf6hcbtfsUb75YlxfIjJDYTU6KqWj
KvGYG1VESdGPlv22B4lSBxXAGBHrbDlpraiA0dRo+dr/6fHc96jOCrJv3uVJyRS+
O/2FVVdrT20QyPdP5Ctn7CZD2dxaLUVAfltKyo2DnyAWLeURrbLMfxZA6EbEFwF9
vm53wSiJfEH0PjMgmyAvnQ4ULWMvhtA1OC8SpiNJe1WhEfuZsSP0TezmULWylX6x
+AB6mekGStBYRWg7jbCNpfTaqUpQ55TQuEmbUcjdtN9Mx+gKJOwzh/v6jva0lsc0
0fxMM4kMMnsSOb1JZZRM3V/h95eVad53Q6egQP2WYnqsNpNDEyghc7Q4EEqaK0iZ
aPJbzC7CR3XIluVZntANSJFF6mcCz5wE7Cx5R6sWFAxEvaEC1qj3Gk6xsosjPvHW
ld6uIe5ECZL7DsAk5X6Zo+LtXZaBiXKR4+x3RpbbrSS/xFIrlFxRr9enmKuikTyR
/vYMhOvTx+bCuqKkglyKDQ97WxmzchxnR29T4JtR5OeHxy0RuqVO+P5YV9/QOOAO
ZiaAHAvqa69vIBHgiDv8qlrDzmrU+YOmBA7lWmLcPAbcLSa+G+jSzfmYQgoH5QOp
XziQ3gyBqV7OfOLlsSICVoGJiC2IJ57/PTq2RigclwmsKKzBWPc7SEPfGIfZ/tVh
deLdy/LmaD4nbuhWIUXQeQOy5XZonG+lKjbbh+WyTXTfHlowU4y7hRA4EevkLEFU
lt6/BVSZAB2NMbR5WvgYTyEPtIiLCuxIihP3otd+EPOYRJP5/vcG8P+jjxdUjlM0
ZwazkqmEUkR4R2b788bS4D0V2wBhPUX0gblJTkKERDC21wAuK7z2YYjUSA69YyeL
B/XUu8PCYCAlu4XD8LuDBG4itBUEVXvAKas0/aIOQcyDiR1LxnpVS7vFZTrJDh92
gURM9cFYraQ1T/yb1bR/RxqbymJDeYC+Lpf0IkCaCSCUFdM4ebKJGnPkq4Kkls3I
sWK0jXkG7Jwr40YY7LXdrf+5aSlxwEIPGNZzWezrVOygq9AcoMePFeY2C8/Q+JIE
Ef0y4Br6fGyUZsG8JEKWTr9Sw2IQVk0sHE0H2AVcx+5XDawVtJCDxeAwKQlESs+p
3bo7rbe8I7ZdWbwOAZKw9jwaZpu7fxDDNlbfxucyWSt4YvVpY9jhxMR60ydAXmPt
GgpzLApbt7TLHvSufHJRdO9f4ivijOotsgOfIIWME9yojH3yidogAY9MM/VTZXbv
6yYIEu6Oei3Zp4k39SJ+87piAKmu7VNyC9vRIty12G6K/OSQMUXuFrXmVsk+LCSr
N/wXOJQUsw/oeeeM/LUngb/Ez/fcYOeoK7ybgI5XdGu0MKis+bMoL0aJ5P1XR2jN
YtGl1vkfKKLJilT1pkXzBIxrjNPCUXXiNsk+OSM8TIu4hlvU3YOTmBPopX8ZZvfh
zSY8EH/qviPAmc/dqWsKKoQ6XJF/qgTO9B3sYHl+AVvAJObWg4iGCLCRe+/t88By
KHohOzPrwT3O9QvyGp4cuPKVHPZKfVHIpP6cofOo/kSL0j2VUv9nJ+v4MTFu6/8a
nSTfVRJ4SVAfDWTz/jSnYnt9s213ThoAwUXXgGDhLGRSkinD9bWbjJoJmLRQS8R0
ZGYnXDpJrAT6euU40goQ5Luh9+0dzIVMioXuJ1uadGWsjKnyipwqFyCQaRRNXP8q
FhcziryCj3OkRuH7f6FTeVWi2jvc16Rbej5YPC63VFFXDtCjDfY+xrpP+XMQWwCf
XCIBkCZXhIM3FpCRVIxlfayyqu0iqpNf8LkzplrZH2C6qvJQ12sycLufLt+jsMkG
nJPHRVyyFtuGw6G54EMtElsBCabwwOfcUU2jyAweE6hKcICeS2RCl/daCB56fzJr
ldTH9qZSxwtzPkk05T3TCuXRg38dw9kFVMsRTeeJX1maTtwQwYmzRwTpcueDDw6b
PPJZe/ipOY7OvYLfQkoS/U5tNJKay9K4g3T9d5U+nIenYh90m1pVeVt2uc/G2Xo8
WRRDOllnJlTERBj2c130S0EHzyIvfXXHkUueVZ2ooyzpRVgde0lg7C1cFEv0DUQz
gxWxlpnnveflCelnBSO3qUCMaaHf7612Ye0QbYYp9rtYtrlvbSiXsTAezWno22g8
vluQy+/5I3qWy71KPMmfc0q6t25d+yvclEUXR8PJNSYZf2ALTrB6w9mvW8CW3yw/
GhGeDL2v4dJ/seitCEW7ZspRfQ5SbfAh97fhNaK+H8z2fhNfosr2N2PPf/ZcgqHQ
+RBWLykgrA5Z4Ig1tHI8P4zGH6euFH1OLiXxOxAZllu1+jpNZhORotNfh4+u/3/4
s/6T96yGv1nsZjJ+oTW/SWAnzKgSb3aG8I4GnqZ5PEtDUw4H6NDAVeT6YPIkVfLE
gpEoRDonk7+uLpUJ9GDyDk8zLt+OMf9NvkBN5MgPDqPIclwTYlZ9i4U/ZlsnAbC8
6KngmeXJW0ZN3WM9S3ocnQpeaJ8v83SZC310s5BE/yoCMnR9tg4aXpwyebV+D6AW
B/kCEgv+djbH3q53uVWsX5pqmfX7fCuCOKdBBACXiXBiPtT0yR5wSYtTdZYaAbJK
eojjW4DDN/NvuzRs1RM+q9DFM+/HCssEc7HHX0qSJKNiGnnm8uo4UuAwC+srE7OY
qdTovnPamqbESxkUGkds3ZjmksFBhIsTutfCK5lVyyo75KyBmmy3l2GhKN8hBMFI
2IZ8CWU48nf3fhAuvxUURZZ2nDKWdSma5pg7LvcZdYnYvbqJRSNu0hlgVBaG7iy9
4tGm6auk7Uy9+f4FRkmriq0eDCEMI5Ij1Nf2dmtDNEw6JpjHTKdKrfLBVnwp0UiJ
zZ/m6uXE1BzhBouQQ9gMhonao68oNyjacZggVvsCwsjS2KcYmHXHwDgTSGSKiqpW
MB5DVOH8jLZ4zbJ7wuIZQL0OyQQ87vDKJ5KlkfW/qRNeq0XU0VKheaI/Ik4YWPqx
xrPfDxtBsRRTQcCeXse43mgK/22WhSwV5hWaixp7yhzWYybpIIxnJe4nYFXQ1QHe
NjABmyCtqkfFHhrfXSn3Baj95Cx0dHEZrjNcva97b6pKqnIuxfu4c0OOzSF2aDYM
qcioYvuwFs8RcwV13NQqXau+cN1/Bpv+u6couo52W1Rc8ZL5wLNI64slhX/Q1T9+
0X+Khu4IaFIOlLQHm9mF1Wz6AHHyTRpcvHh58ZIK4YGelkx4EGLlL5Xsyh2g5oPI
yXRdahQIWjVm+1mtZIXA+MrT4HJ19NWYAoUx84zmJ6aYKU+3iAxs15qL1hr03GgU
xJ9zT2TCJnilx0XTJclSp9LAqflgVg1BY9WSGi+ex6E=
`protect END_PROTECTED
