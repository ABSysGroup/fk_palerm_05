`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rwf+r7wy86U8qwhSUMCEM//f+O3maPhkOHizGc2gZezm1zXl+pOiICFVLxFMTY/B
mQYjdMS9SUAUaT10BxsqZwx6uqQuk2htAfuAXRG5FZsBJN8uAII4iNFeHFpQdhuO
CvwMGEROh4I6aCv7Yy/Q7j/DCRRNE1UreLdQ9WFQZbDz0vvlrsafaP04SKPpVq6+
5g1gq3xu9k4GDyDt+hnmtG2eTdSrL88CjDqUh4Ro01B3UZ0CdfBuHM6UcgtW2Rkz
crCPDMMrqUp40GBIA2cfI+BKD0EbHVr1fM63bF1zv/Ni5zqHXSq6IlcYAjB05yxK
Um8b/gxghpYSymJ7HcoMUlRUQ07FdZOTO7Nv1821HXMTLp/4SGGzdp/ugfpTfzHg
Q4zzZomkHjBls9g33AZqFSiqqy5cEcRqmICFDo9V2kYnJHuxCnLNmgE46BCk3VYK
fH/BvHqrylzD/rQ5v2hjLK8fTrtpS0EbDU1BOsnpA3o9HVyLBGmsp9cE5eocBYcv
KuQp9kRA40Vv33pt4Lks/y2fmz5XBl8awbgIjLqOB36eTjEIWdAQ+FAwuJGDzYXM
5RgSbhmT6bRtpOTJyikj12FU1vNzxCxwux7Zkz+U0Lupb0m+TASI0Q4DiCr3e+1V
nr8VfTB7WsG5lTIjgOpsRA==
`protect END_PROTECTED
