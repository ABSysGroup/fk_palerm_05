`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gUd4Hl8mplZ0E0RFFzFQ0qmvE6ksBY2UzzlRsqQ0BdjF48fotvZG1+f4YuHb9iKy
wn9rba/iBt1Zin2ZUxuElydmY8erW3XQZOWgUTHkme2/gQQSNLEX+ZEv+sXIKXkj
x8JFsTU+Aw9o1dME9HWR6nozCaO4ivhMasy4LM9MH5Du++iU2QoOA7a/WPtHsZNC
wMPrzvvBH5lzQU13LVaheUxb4/2Qkl2Vvrj88OhkB2ta/pQmOk5wCVJNQX3s+hkG
LTlcwcopDNK3eeQ2ZCKC9IdTXfSa6wYFGcdoy4aHdYQkLDOH+IkPvjtV9aQTmYBL
M7zNXWbKw+q22mtlNwKJAS9kdSxWTioXGpzYUrX1cVOe9wbD5tOUIh0j3W8p9QV9
FDQOC+sjliRyiTtR8np8l32tPvXwiws+4BC4Oq4bXKGiXHxfPVcSc61VGk6SNw3L
GTSOIBAZIUJLfD2nXbUFyCzKxz8Cxm5NEzQoxNZG2fstgqinV+3Ei9UW7H7hMwv1
EGVRQ6H3hHgR6EYYrped6y+nwC3aGcQwUNqYR1KO8+I=
`protect END_PROTECTED
