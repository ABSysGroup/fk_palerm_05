`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iaFBb+u1vcB7/Si+FFH1/bw/muhqgyJAJ6XeENCAlqE6zKygL41brW5dj3dVhExy
eXuPW8jJkLIX7rOfzJCx9Y37y6DMEF2J/q/wpSVfprY4CdPRY4/gk4w3Ys4F5DtJ
c+2+7ZfuxqcatLtYT/yzqhgzhNU0tltYjZ4+IhXPdSeRBCPWPqirI2OyyCb2RK+m
ToNwAYBg2tkoY+3l2Zf0Oj8kqXyTuFK9vcu+44F8V2JlMAPatzOK14Y1PGqWKmWV
HnOU77Zkbm/Ww9VdunAk/C7vXRHmBjUio5tg+K7v/8rH4xzPb+GegmqweemoDgTE
F39CEebLzMTDdlCrB204BlsY7bHR0nvgScgfGp4tvXIB78lT6gYUFGdaNCL15+pu
SKoad9A3XAZKq4QGICxqeTAdQnbyjC6mFyp+zn8FY2Xyzw8gJmp3Vcv5naYEcwJ6
frmZC9CKvvHM34zksBAwBFa4gVRF2NkNZXUFm2zheiyaGquTt/KYmn6ubq+/oDkS
h5elVSkd+Es29Jv79c1EvWgbd6k25SmLGtYZvpw9rBj9D6rME4HXV+k25at0djT8
l59AZKK07yc1cag+/cXpJXAyrBV5Su+PWZBovv2Et1SYEsnCMfPhzkQhKkKHrndJ
`protect END_PROTECTED
