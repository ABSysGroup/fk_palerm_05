`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3K3nEOkdP6KRechiyuBPg49PV6EOgoApVqROkijOwVEOna0P0F4u+b90XgDRlIzq
x7KsOoBbuxOoVu8VwgIrr/N5y3mVjAWdjHKY2L7Px46uUVQTqHgU89+EffI/U2BX
EUn+401aWBciRSmeSxluM38FmZYwT3ASYsKYznNwVuNaH63iq8dg+5d7MzthyTXU
FyHiAZeDfm7ojNUhnU4y+vS/tIV7Zi65Go2TQ0fYvmIaHF8rXLFr9i0hsB8JHv0G
Pt/A7BIOkXT7L+koDmSlleu8o6j+Uj94KHAkRDTSl4dkkFqeizPz5HlTqhuwS2j9
sJOvOzUFIxhRnYB5CE/BiVQsfObS6l+RbZFH0jj69pqkfptxR0JKqeBu0nQ7dlAW
NwHbZ12GDvYuNFleGxrJtxM4MMBr+B26j3iTrY/RMyL0/nLxHXg0SWZpwlWhRJJR
VRgmmCLEEqCbKxYVhp0P/BvRsCMG64+vw2+doSWpThcaCQcDt6m8psNQdYFQxr+O
WtFF0I8svf7NKbetm12CP3SGv+sMaT5jksVTnTznGEFyhp8L2OAkqcDQzvD1RNhI
7NUxpcRDfWOhEx3TGk5RxrvZpmtWz+x1FS7jXWAU4+HBZDDFVUiZ/Gz6ZJjAdHzj
pM4RF5+92yKAeILLNzs7JWh4gUq4JOZMbJ25C9JqYhEeQ3zoGdVyJxe/Eq6xrFws
fDmvcxjPijXRL3wE2rq4xwgktm7aWn52zbVgh+G8vXZRtMq1GF/9CiS0hF/AgUzV
kZoPo7QtHgkNyQIRbn6mrFegrqkhGI17cbkI6sSFrqp+f9O000jVdxuZDHGCz9nY
9I4jez+0Ge+/6cb7XknoBz4ylXCfcmVFQKpxwD68Qp5JzR+o0qFLj6Fb1pWHIGoF
ZIK0E/hgWoc7E/Hy0iKd2f9eozEeRFJYfzcvA3bVToNtumW+RqQG1zwVyW26M1pT
d1M0poYH/BpQ08ityOKhjiN+94PO8xXkQFjyJQj9rtC7kpx3sxlalnseQzJUErsr
3wODvLf34X9Hvegxf8CdDiIaOVPXHVYBgFqUw5zelhGjyb+5H9IowJjns0k58u0C
kVVvMUSVZgE4k00vUUbfKxLTgg9/i/SWTgCvqdiFbGsNIDozQcPcFG2Lz9Fgujsy
xJs5Jj5IEDaxR2sKQfaWodGU0vtIokG6aUPvbFSOTs/WPq+YG1ROyqaOcr6+7wil
68t46VnJV80OgrxEZhIooZ7w9paR04S9sWQMpg0Di2GyCBqY8EpmDBp2YqTlJXtW
EosJG/J3Hu0IJumrtvyZsH7k+3hUYj4ugBBfxedz11HS5rwaNq7SYDE4jd8Fqe5C
Zeflable2l6vBJgQGv0tMlZliZSkTwel/ys7veG2X0fKdEZ6RS5KMf1ZEJUctJWg
QegkABcu5qoFIloJTmNxeVkDEU6BDv8FXh9P6wG0wyhOCimt6sr9CKm8kEB94y3/
kKLvvWzFL30BdVR+vaOMg2rJZEtQubDnyEiM3exuB1c/R2eYtP5UThCrvIF4COw5
IXXCBht1a9FDP4sOy/h/l3wqaPFV2uhGGAQigWSJQe0iQzBR3mdFtXr0nCzfNUSi
MkfaIPnmJaZ273+GaxFXxzI1aqHV0oGmcjgkenWTvFT0Xztwv63zfzOB29haRgs2
/mv21XC87uS4HpQlr4r0yw==
`protect END_PROTECTED
