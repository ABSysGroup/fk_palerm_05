`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AYmqz54EfTKyunHLJWFkgCOMlWWuNN+X+IZHhDwm3sgrIZtCS1irVMjQzkIO7Ppw
Zk+JmsOkKxvuHJXzCQRpSqQSEUyo31Vt35pCjY0Y+HwToQIaTTg5NtTfZACQB0fe
lRxZMfyw6Nr3KsJTAkxDmJDnrdrZ8WSJQtQFDvEeNkEUmNnCs04lL/hjHDT7esd4
aY0AWNdSAOSUR8i6Gu40xEuQRQrvSdmAfAE7Fos2G6pIiKBa1yoXy2daUF18aS6D
6cV9wJOHxNA2jfQZlEbrqo4TXV+J16mfSBSkS4o3ULPEX6VL2eZTaeKeI5vJ6t2C
tYQXqjBpxhVK+86EiouPT4jJtH94tS2Dd+0dxM2V9HTgxHD5wYdvEZGOeC23WsNe
eOdWtJAS141P/cI0sHVlCWPVvjsxZ0H7utMsrmgcCAhDdU1Nl6rQdktZ5aVTfJd6
NIFyZX99XSrekG4meirStfhyKhdDSrioOEX3p+Xvil4mDIl07P7wbDFNIftLpZ36
6CwMlDLgUQIcQiIr3sJh1d8HS4+ye34oflrPm2W495GBMsZqXN+ovGR/GO3uEuMT
i3OlktR4eSxkMPT8R0cV6tTOZw3plRu8pBZMqaMaZwefRBbCHvmGeXcFzdQN1aGF
Edmz4iiDK0+8Ikbn2UwOaCwcwBwDCQZZUDTsCh4b1eWHL7/q/Ao2/5NcsZ4OLG+y
V5J9qcgg6CBF7oStGp9d6gZkhiZFeOeaJTf8u6aL1qBcSEuXCYlArE0PgkLfAAZn
1z5YB1Kld0aG9W7zbQCMVc0FiTSNJ17zbKBgVnFALEcimXbq8lPAvOf8plui9Y+z
cwfD4cMGUbpRZzACL8m4STqhTUaOHsnrfstrxUzJscKoKwbvCxjH7sqFfE8QErGV
TEDV5Neh+C7De8FbSJTurkdhILwW4DOMOU7ep65BjuKQxCcq3OB8lc+ORFjLBuZZ
`protect END_PROTECTED
