`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vDgU4wtv+nu3fWwzsDYqI1EjjxcZ9A4sNm8BQq0BBuRr4ceZ1VaHWJUqNck02/vS
GofvVqj9npDM0EypWJdi41zLjiaVlC8gnOCF8kZv09dbaPhJkt7HQvDmYlxu5gBw
X9AH3UtuTP5JZi/00A1Dlw8fIQG/mWLgVL+dB7BeQoXlwV0MuwZ6yDc9+sX/LtEz
imIJDBGXpcJn7MwhDHVD6VSDyr7/1/NrBo3yasrH8zOyYclWhPthkHpJIe97/KxG
LA27VNru0hpmzzqAjy8MGkXkL4m4Ry1JJ4hKt8fisbGo8n2ae/BjHMRapMP0BYSl
z00+sdCvf6P3mKbd09dj6AGHpNMF0Kh7AxoKqoYd+OJw7h7D0OTk8wuo8rbHGvCM
`protect END_PROTECTED
