`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0PL0pIMes+4ljOwu8IZJBor+kXEA2ZUe81F9dfugiCaStM8zF4sLd/MwjWjdWL18
zsibsqiXnh9Hsa1vDFwkqZcXM1gZM8UlLBf5oc+0rdPCL5oEybTxwDmKc6icD6hy
G2QniADLk/KNMdKyfEL/nXSQedL7+/g0jM1o7R09mucbj7nQrsL/oClLoLnwGSZQ
ZyaEvlIV0dAM/Y7RVMg7EeshvTrd0o801y01rPii6rJlvqIH+VI6GoVz4YKpjBFa
LSpWwdJX9ZXNRvTCdY82aXMbwhxKBLGjqFusoMWtXVa3bRlJGhvq3ysunUmbowu0
DqFx+80ojkdg7AcsXu9T3iIgoIf4U7tS6OFW57mDTZrSdq838r4fAcC9vDgeMgVe
9dqRv5zgUc5nPEsAX+/RQA==
`protect END_PROTECTED
