`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I2peAcaIrKPEdf2JpUA8nhYzpxhWmyQ0aAlWvktWKhIAEqUk5sW/8FplAfT5/267
jDr61BTlmvKbBppn2VJ6/j2KPzloo6z6qOPtBjHhzLzk5RHinErXzfl5a+/6EyZC
UJXcXW3j19pEPXOqzV6TgAI89CzWZ3jeElGb2BQj+Z2Lsgpd3YTVeWHh9btncYD2
COGANT4ZsHakECri+CMKk3+LJ+n3qDGJ4t4aAFaL5WTW1MidI1lWnRck8DTzTglx
ndHrACCmtQoW+DMnYc0eEQhsl/08D3CywCtxHY6pRSrNojdzxdT9xaazmjbNW+67
V8sKCEfMuFZKIeBQCB8kKwmMhdahCsV9YVR+/rzadjzTjA/ZaAbncVeFIaj7kbwb
ljfLXo5OZDIqASSo7HG+Of0KZj8lQ7Sp0I76MpKJd7CiUiBgppUZZunIxzaml6Ll
rWTIuQVtZx8PuP0r8E5iIbpWdw6JaEbM/3s0wHYiWh6VQ7W8CmFo+ksycY0cdb9v
0OnEl78ouNL7WutOBV4OjjUg4birB+2eT5hVUPox8y+bgawJNClF6wVP/tTY9CG3
jlK5yhl8OEpl2xcGahkW770Yh6ccszV9TnfukEH55p2NOCaB++ogUp5Ovgc8k/KC
1L8njTgyE0/qwFF6BkLy6B1bF+Qe4XKOpj5/vRLnOGnCNSsPE2uL+po7PfS8jpdD
uVgnX2R+iWoJrP/RcThH+vBGL9z6nRJYDDBXceECJthHg7oq2Eo970BDj9VJIsQT
zReqL2YyGqZd8LkbsNm6/SNikorVQXoK3+MbEzQ1SDsrcky7NqIoz18Dh2jCqkCX
sME/5SCJ2XkKH11Bw1NVsnUMkZ/tgyIyqLvaLLUnCN/nCdh/mUixDBs5eg9qXPNt
Wb5fpuJSa/PKU0UvjZ543rjax36ZUAs+MEtH4V4wk6+lNW4j1lPZkjplevX1Wvac
liHi8k0BkTZiAlTXaqPGhcaEcMCXsN9HQm7387K0+/6waQIP6vusTKCOS+z+V8V9
j8jlXO3rcM+FZw5bsa7snA/pWWm6mvrK1txL0JQKgMjHQ7udJt+/7XMB8JLErVOY
9fN821dmBS+CJNBBsgc3vbKiSMl6QDhsSueu+99lsD4MuSHIPrdqY7sMv2RF0qWn
`protect END_PROTECTED
