`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FWRv1IFtKucjdfk7u63eUcbEYd6F4QydbUboMt8C04r0aKxsOLQPdpYqtB1YderO
vEEFa8TUNppB2rO4HfyUnfHxWGvdRVOC9nm+FVZVGMF5ysFCUzBErODeRHx3LsIl
wKWPugSxCsqNqOOe2n1McNAFsARjkvtsxUXkpMGYEIe0siQsHdcmizLgY5nsajML
loWT1jgkciOjjwE8WNAv8dOhjUd9uulgem+aT/Sm6FpoCML2m31ZuB1ESNpOmGGE
qvBsZaPP+8nBZXMCyligXZ9aNQrGLfEQJzjIw/m1N2f6i2+T4YbrkX+GWwY7kGfv
2QLRy4ZIlmMwUY4A1+6UyOx2355bex6AXtouVuR8c83ktdHTvlTT7f5KnNL8Zbr1
XYhYleWnyUwS6LsqY0lo9vtwXDnc5wWM0WGf5BuP+K+0Vqh/vInq5UEXd0R8KxPH
xv8KqKx9Prwh4o1TQfZT09ElPcDOrWnBTtRezfS/SiyNJsQ0bxBGgf+VRDJvjzO6
JOeVH2E/b4zGxdNJFWUg7fH9+KDzflXk0cpV7qNKAEF5X1D8QIntM/Quu/uYIxgK
L0hSOJjf6g5me/z+1pM1W3o+5iRobFiFwvsWXrPajSIftW/BKBnmX5a770BvdQb1
a9RPNE/rErSrvFr7Wy7+T5LoeEDMX8elB5A5ptqP8r1BsamJm7S/ska1KoFQ/522
`protect END_PROTECTED
