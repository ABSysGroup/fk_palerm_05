`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/4ihVMAXa0Hh1bD3VaDRenGTIb3EaXBoBX0n5e1LjCC4KlQo1hvpqInN9R6SMI3Z
jqnui52s7ZthaMrKSX9Sx2F9Yis6PMNMvWQ/jGRDS02p+21ygh8691P8H20d/9Du
0ofgeoRsuPXpOdLL6Q6pd/zG0rdWiohHtL4bedFr7uHpPrJWS6h26Vlen90KCHB1
qJtgSkWMSbtcu6EOPlFK3GGOs57y7uE3zCvHQevdtBMXrcH3RMdPrLXNblurcfE5
gZQpUEd352DtmvkvmB0Uv7SNcpnK/Oyt7EOrDkgjoIPMlMX5hHu7XVPekcck49uK
h2800vElwlM3c9USVEQWyNYUyvauSCgkn96K4Amac+kFmk5QWJvGC0NLnP2XKoKK
wuN3Q62z+g3nxSi2ZA2rzkNG5yefjtNuOOHlWlwGxFt3zFUB40uCix9mk7SdoxYr
djEa39If0d0LuX7WeeerPvasOy3ZZoP+dpp+Zc+gTEqloZ31qFOUfMDW1S6JNY0M
xeUIyTjJE+odLaB21UTiMPpBF5a2URqmDy9LEdxJl6tTKQmmHrwWdNvZx4ziBvlK
bwyGFmPBZTQVuoWcUIonjJm1RRISCEkKHFtVNWDE3oNknnU3suZhG4dtiLTQF3F8
c2zZDD2N0GNVAEWiNrRJ0D6fGpbnhOFQ4bt8migyw6poxoDYV/EX4LnEx6o2Bq91
EtaSJZNXnBKkgrK8xXoqEh+X4DI5HcwqDLzA7pGkOhADRO77iUPhl9nb5+uYUOU1
VxUkiSbK/9WXl/7mEyYvRy1JSiUmzlkn/31eAmnDbXJSQDzgnviPBH3GrKqO58UJ
alvyCElBuHSezySp3x/sFn2rPUYONberIw4QtfK2X3nBJ5kCpwCHFV8/wod+lMBZ
navmWMro+7hCNpQcSSa4ssQo19p0Qw1pWB4P77bFE9o6vSlw8Fm3A+WNKJV1H7rX
IZrRUPHVBudVHrguxL6TFwlYnlFUQ8uAOitiLofunCFZAqpMBR0uDlUoxrqs7vjN
QG74r/wXCzNhfIa7vI7HCPrpJt/C8YAoVbn0VGj5M90GI6gK8HW6Au23yQQEmQHg
hhqjcIp/dI49io4/cvB2f7P3iJFac4PU/x+9dAoIj3etwIQfiCLGK5BN6ZVH71cs
tXIOzcZu6SzJzehzNXIQj5qxgNMtuaBQMYmL36Gr53wLcooq2oXqgo+WRoRiVuLT
S7i/ATHOWcZ6DJv6OwyPiwGofSVLWHc7i7y4Ym8vSFMvac8xHj9UZf0t80Sqa00+
3Uq34zxXgaHfrMSw3uTP+q0GGuCRxJWGpSD8qSaZXq6KTVtFcQsBVgeVOAk7Nv0O
0RFEkInhp+jrDOU8BjjCOd5V1Ni2XWUYUGx3Esdmw/F7O2AQIy7xHAk2AA++GkuY
wny0L2bS4jOoIoE53i2ywbVAuYh3yFRq9QRPrF9fThSBhrpjw8y2k1Xj61zOCMrC
0lXKsYkMi4vTSpWKfmvOsx1eBOnFNJBAqZ+vGajRxTlliBLsXpLt09xpRcmYLTd4
F1rkpUXqku9yVahYf6TKuTH5aveUfFGezX5P1v4XnMZ87qyFFceO/RdaptTb9O2c
`protect END_PROTECTED
