`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wqzi84zzNYYXM4yGA5GR2zERjt7nIfJ5M9mGxTHz3eECsgajGEz7/6crQOY39ZFg
n9gDUKGH6pdv7Xo1j71FfTR36e/mFMAVc8t/nUT/CPvH3nncQXO43XkTC6pPtfRw
3/gbxCsvwnYR+dPe0axh1x/Y5Efu8NFV6JBvywNrT8HRlL6bJ++cWAxrErvkQ0Y9
dGDWvgaoSP6p4XDJaZhEqYfqEYhqW1KW20LEye/cFybajjAF4G/3eF5BTRdbVSkG
aR1X0i7DLsdAlp4N/e63TS6KsC5wNQeS0BefMy0fGmqdFqMrIuzoynlOFbUZl/jp
`protect END_PROTECTED
