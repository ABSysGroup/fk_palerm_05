`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l+bY+g920+meIc6rZKEOrFPkd10MXIRoCDedYKvVqkhVai4VhOfw3R+UGFnii1Yw
CLGfVCiC1pgzhchOOFvgyXTMydyAlGzXjKXJZ8EljqzZAkNujAG74XsFxI37vDQm
1P1Jx/beUeewQfYHLf+7QtVXBXp+qgEtdh/cN3vy1rStBlkq9BMASOPFsh7i8F+U
a8t/ewl/O3adFH9f+ZiKlCjGhM+J68zJS4pNT26fWfI9X8O9jfom+dwd3nNaBv3/
pLmp4trS/C7iLTHXgtgM4Vbct+sPnMaS2nK4nvne49nuETH90Ojw7yY7HIfOc8zr
uIdI9+PasF4p9xndlpWKurZAIUrMw8coQRgobDAWyBEQSz7MQbq3CF3fYdbU/aet
fmUkcT8moQdPayELylCcpR69eQ64p3YYhAjWcGIu8Zybl1+i58a5Bv/R1VQn/vE2
5dZG0U1e13k/SHgHbc3G6wBBpTzz+f+7INNVvdcZLtsx0wXloDrTIqBXnAgW5KME
f1lc81X/BoR7kVqbDJ6H07PSRzFUOiFMt7W5isa/Tna1fGB03Vt4KCxCxyQXrRzc
N/vvJVYnhdIT46vxsLJ9UDzQEHkgDEGlQ5yUWcw1xk3SlbTGrF7ug10dza1ZKb1N
dQUWcPXs80tLpNeGjsE9xdQRdaJidVcnHU/xDnzsjUqfnNu3FDM/o2boqizL0q6G
WMWNNoaFyWcuQl4QtX7Q4PfF7Ofy/WP9860w5GiaeGTkRCUnONUsJOyU5gniQ+MH
lcQRhQV7W88b8DnIpt4CItwOBWUS10ulbhHQYaEWyiO/zdGI4c46+EsyqOzwaN1Z
XuATlb8//u9uLA8lmxtl4lPfIQsD2d0PKKRgFfbmCt0saZGObtuT2ZdGrYTmq7nx
GdgQcmSW8h9aPegnNkclS2Ej5sK5QJ+I4OCyyjdHB5bkhn/WLiUcMcYMUIDEssnZ
9OCix++otZ/1GDabpRrJH7wxxbx9RPgg3ZNvyrgDYB2eRVftx1PJwExBg3xT3rJI
QgsuHCt8kx1MOQ9nfjZTFrFunpuJhfEyGbwivfw6hR5miVbFBFZRDPUUpoqudmRn
565ZVZKikfvnkOAN3y+3m+dBUvGA4AqWCXEBLErqhPl9lXLWR3Ougq++653jh9L+
IzOFxiI3jbtJSpnwQsJJKQ==
`protect END_PROTECTED
