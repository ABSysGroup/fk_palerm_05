`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t/E41c8Bq/H5HA4k2OGAPfWfvxEtGtf1nq6AlPr6Ngu9weWsRVthUwVpF42eRrEe
0SLYQRifls5jmi9MBZpSLhJzXHXvGi4GFhnrcmW/ANYkzjfF27N89jIrXj6IW2Oa
aj5ON6aXS5X69QWQjvq5B1ySxOmMpNo9slbBikWoumIar5vK2dtlYXfVVVIZuarI
cm/RpNeIwivgwDXvFx2Wcn18WL74aJYfswskNKK4NQZPm0Gwow3DSnUxoMgeT9U4
Bl/oiL/s27wTBVHynA/XKta78nmMT2/EJmlNYjfoDL2H49qUGrCN3qK2XTnHArOh
tAkacXpEY4H4CsxoOxYDaKMnnm/9ntpWuPJqpqjfLhF2f9Cbz76OZ9I5iVN798kn
A7z+LzOMBuIeTM3CleanPGRgZDoNxxsNMIB0wIJfR4Cs6wDO8DGckrc2DJaaFun7
A4IBl/SZyVF3JAHPfS9rmNeOpc5SQ1f3K9AYarKP7hXAB2ZonxlvwhAv6zsf0ABi
JE3CCZLBihVPXsJcuTIEer8FhuZruUjETYeEBzvi7B3z6M1Fcj9RVJw7e0Vi8cpg
/oIXuTv7RHhMHgN1Upo6U2wfT4vCiHt5A3sncFGEH8lhms9y5w9lnNpI9wY2f1AL
AWTsfE8ozckUwlLIMUiY2D7QMf2w4U/JYbT2x9IWmyeryAHSNzgK1fj8nsJ+cm/J
ivmdW7JedGxXn8viZYCswE6E+O0CJpvPGUtUYUvldr06K3fHQtzfdGyhr4HqoNcA
AO3vHJLNFaCwTeqP6Wh1dl9L3euVAGd7AQx68v+hO+gDTqfK8vChNW/tUs2muTTU
InsKbWo9uo2DlgPsr43PGXHW7vIHd+KSt2GkWr5LaIboWKj+lKjFol/HIhFOSRjG
n3X7ncWFLpzh30NLCcAE5l3AyURAfWl5A4k0AcxwAg7n13BeseC5Y5c31tqzpZa8
aph9N6mHlanudLAPN8owGtzGQ8ZUAgJzjlqDFxYRM9uzjffqtdbKQTte7/N1v3WY
RZf+QYkQh+jHw7XON8h0oZe7JrbqMfoin5NTQjKpCLzyNq4z6ui9LCi3ROoLddeV
XwCJY0uhigC2GSfunkuuOvyvizjw4hRthZn0czkb4JOnnZMK1FkL9AMw+878gPFT
QbdYQ33HiiWhXAh1hCkJMLSnIgTNcPeKuP4A0aVZOXQLCZZxo1Wvwt4AN3oDMojM
UQVkLKRfjgE5iZEsIb0O10gVtgrocidlzyB31y3UWWagBbI8mpqloaHmvEhTxHgP
fLMl6l3RXNuGkhFz/6N2rF0idTpoPlckOv6BnZ0p2O31TGGiqFiIXI7Qea8mt01d
xhwMAMRRx9QlAvgBCgPrfW8+PRQiUDkwLUBkycIsLQQQQcNEEPj4SC8sX6fBB1Rt
9Wl+IVEfIAV+LmQG5YE1HcgnA7GPKLW+9d+JTvUYXtaUJDqPMRd++2/HXvq0fwBD
GtNk2kHb7nsBcLdfT6B12aTNJqyL1ucMgIjwFBuBhRr8Gp78wYjB5Y/Jl+fEv47u
eO2yWjIsZ0GPxIc0qqv52L/JXNvbcMjPe4mwtrBoINuBMWqgauMz5F9RPd2MtHI+
epT0FapScBSMierbReObOq5rwsUu5RZ9yEBOBcMsExtH4CT+n1CGwJ0/P07FE4CS
79r5+aaEHZ01Ie9rwResj5cCVCIBXvZHTzu8TOiVfGq3RoXtATm3Gfc+l/HgD0cH
kWXAfrcOqCBHyYdux03LkQYdeaCIUpMzP7uDqOPkHv/pUJyOj5pT9ZcrzTEQU2Ug
S/si3L5dMqrr77MTiDoF2dd9DfSEV4r+GTnzVmaTz8b/Xgq0Bk/x0/esiqZeEuQx
h7CwGh2/yveI1HJ9HD1Qmp4BaENbR1whRbI73zMLD0FfRm5WGM6eFPlQzU8h6ymh
qZ+KUXKaxXc96BwGHyj8Kp5zl4UNfFp2ss82QxS3t8Jekdr+c1KHAlebvktp/5TC
dl1EIIzXCXhCzFHKW5pJob5ed/laKc0iCazmKxBCFUcNXahmBVfKRZS5YSUkKdmL
2P6L/1dxbLFIHmCVc1Lqpqu/KXGB/F2j+tWWFa6PdlGNrI3vNjSPfByaGq4SbP2k
laZo39bJnASTNguzjDjUls9yZ8xclwaqgs3J6NOc63wRVVuYdyE3D5tuLvFs/0rw
IEotZwqT1AlRnns7SFKUHu4X66SWGxQXVVdEsajqkRmWN4g3d+1hpW1TNgX1W1Hj
7glYW4stecy36EVisUbGKp/b8L55nsCMztx+AQjEs4hp5FnwYXjlXnpYz152pha0
`protect END_PROTECTED
