`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q0Ju9EJHUY32piFc49aaRJDcTyPI8ljCYY0HG8nlt0Ej7WFI0FhgJSnA5LjUfFJO
2poVE+P9iQYsUoHk9Zo4UQJNjIxMwEAmkisQTlXuObSl5IoXvgKMggIN9smL/0bI
fuvcmpRSaXTvkVRrlBkKkKym4QbckXY499ZHq6fzSoOM3/wb4X6ixnJzAeg8dkFt
liwxFKsw5OLoHobSqzd08sIJdQqMmDt/x+4Y5AFbx666O6sc43PR79Y1pGKdZ5O+
E5pGZ0/p4bX+tjMgNm4LV75/3uNqVvIwCZ9WH+30avSy1KuNnu4opRvYVcNj/4L0
24Wz5DdOp8CVtDdt0WnE4w==
`protect END_PROTECTED
