`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gvNoFTEZIUE7eAmIGdLUv/hetPUR3XjRAJsNcysGfaQ4M8PLfNjYSzMSFJOq4LOx
Amci9Btof9LHpdzzp6+VwdPlkonHKQisH3Mmx4yall5Um3cp9PGD5cRzbE9BdZyE
q8W8UDyZ4UBAZdy8cA0iUXO+f7w9pk/SihaBJINnsA/IiikN8L80kqVbTGO+p0rL
5in8K597Y4oDZQuTzuALjIRMtmTbiUxvjXewYeYywaKVSq457DO6MfP+QuuwZQlC
ZcP94UVm6rEvBxkJfqimtj8VTjRWuavNEPI27/k0J5fefLDh3y1VibM9ZlfhaE3X
fheiMoiHTxkrAhfKSkafNNRKatyxe+LS3tw0pauAVpIhYWE26EDcZdF4oxCmSEiy
LShznP9/ZVRMpdh36xJUl3I4jnCFmhaer43ddvgpq9Zhg9Ug5rYHmuwYpD+DwOw8
tuj5gcvw6UZnV/tY4p4NQw+6NOuDxusWQQLKuGe0WUzwmY0X1TybcqwUW5VA0kQ0
naBsn3QsfpdyP39KZg0SavL2U+y5ewRiQxcCXhT6McYFGncDyjwMm24eLLWyUSJ0
qnbRWbweCKyZjNRyz0INM+yhS92e+2UWbGovcRUr7vTVsB44kzf6zukU3ZPb2MTh
xIe6L3kdJ3dyUEmf2MQaEtK/WZQ3d7QanbbCTlNVJzcO1qf3GFwQxbRWcD9jZVfW
td/D3TUKJ8HyRbQyYhbH2P88O/6oTuhvR+l3m644lm5A/Mp5YFvVKdBL1jaiMFIx
vuKaa7mfBy8UMTzDyF1xqhFwiQE1bcIFn8Ca5zGY+1yHbNgbjttWNxXWDFPOXHZf
uvGLLXMlY3RbrpZnxaoGJzyYTfVWHxYpBsvFyKgrZEVjtwVXpGcht5gII+0te7wY
aoHj08PIAgvyHHbNlafbeI+8EEjZIKb4XSXLDoMLviRXgrVPzhNiTuzG7dN2AlGJ
jOADYJGQDEC7nwLO7tkJo4jMooi0U1vjPCXKMN+/rNrIYZdRlMjrx+tui0TfuCyb
oFHYcncOVxCoMyJ2/gQTJeJ9GZqugXAzHI/Vqn2SgwpvyoMLp4IJxHpzyXKChPIa
7uEMjR5PhpjDHNqzwSckCcbquQIGMVeBX53GIdHNO967Pk9PUljBtbaRt3HFqpJK
KFp5skUhyD2aQtUlEoolLcZhPmkht/gvwI/HS6D1PeMzezt8LB6FlPvq7Lp8aCFt
Wite3wmwLIs9mK3ipOgvot+M7Lbb0FKBcVFex4mkDSHkzrxfO2J2Sad6cKoUJ7J0
jS3LFzZyD3CXoPi6ZMJWcJvNvGXPbPWCKuWhx1ovbu4WiLbuifsk+Uj5updxnH/O
ibgzWxrF6e5LpH88aowIpxqwoEcuftBd8JdnFUwdcCmwIWdq5ZdDowLFpwowWMZs
DSJu7FPs3ABcF8qu5APp2d7igSC4EqmRm2VKmWafGU4pC+PMJUEtXyUiThYuqWT0
OADnppPiHYaQMDLql0GyIwBGAszHMQwXyVR/RiqB57I7k/K59csjcQgBQtJdmNCy
63LtK3hZb9BXyeg8EkcJDH02AHFhyHRGzkb8dZ1JXYlmftzzNyQTbBwLuVr0EM4T
ZYFMwYjZFnOAA+SDVjHGxleFXQr6a3vQueaffH6q4PFmgHm1FoPec5vfoDAB803v
bbSF9Ci9sigR8OKA0kokj2OFp+JsgL/jkanB5tH9q/j9TTSchMKyxh6qM5zsIu3x
0Y+rbomzKiflzsDNvX+I+GJqkMOqZBLpFMKzsGD0phdvIvunQ9Yb2uHTV6XOd3yE
T31DT4BMtA3dC6QrE02A+sAysoubmRGmty+Q/p4CK/WQlATc77RswE5k12TXNEe4
D4tYY3Pgwjlj+Xp01l7mLqIIP/FVQM2DPT3Q0f2OkWNzCKaMR9J+b3h/sOov3BGW
P01aicpTx2PFFmoaFu6z5/PQVZpDv/1loRPyQ6YVg9D5Trev8Ybe3qAYZwYU5Jxw
mzOZlb9udPrQhS1NMEN9iQyRhzy8/kSHRWyaaEDzDljFXgUKaDF1N9JMWUao4aQK
pHSNNmW7acC/rO/pV1kKCpa3kDjE9CZ9dfzdvIQ4MaJJzchcz0sGpjmdlnv9LyYf
FBSLmyZUK2op7TOJ59l0eGctZ7kTQcW7k7J+81MngjWaSq78zPNDiSf9fNDo8VmV
sww7wGSxCebkJ4UNN3MG8TrvgWl6YYVm+KgV38B8S/3SmJH11KlwUsHMpFqhrtSO
MalqSb9m+K2PIITSE6WIUWE9PA4YOiuizFOMAftsvHy/cSSeX5FGDqLFEkCuKRch
hEdB4XMiSMtWPfQ0IZmPBhCzmzfh7iQcww+oto82nqMHu/WqyqCDNvKtbMhfaScz
`protect END_PROTECTED
