`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GywSR0HwGbblmN2KeSybnzlPIyG3Da+F+Q27N3LM4dCCzV8xdWaML6s62Fb9d6U/
bMGGqN5zgiJexUfMUe3CXfdbXjD5TEpfcFbpiKjpX9eGngXPTp07fXENIqzaAlH9
ZJauJ0Q1i+/QYDhhft1HhrXF/e0PjHvSCYO/XaNA0D/GyKC8dgGdPxhyJgg4TCQU
qnSkhv/zRNsQDj/fxsmakx1YW93pMjhwma1bk2U3chJGTWbRTnN972MM2i6DhaYq
3mHdpsB75Pdntz5M5etmcg2ika41uu8L0ToVqWSUOtLLEEaqpYxToDWBFEGYPUI0
e/n+THpOEJrr4LSVffxHlA==
`protect END_PROTECTED
