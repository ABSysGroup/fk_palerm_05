`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VqHLgXPlvOLufVLap326jgSmqcEV15f/5vmzsfK5XhOqIcYDTzfeXb51mbP9LGff
aiauYzM+CSILiIUl4ps/4Y3doBYhB9bZDogzvDtoZoA8tXhVQca4vlPKKUkq7cJz
oqZ8EsuJFwNS4gLNmwfobhnqQR7u9UPHjkYixE+s2e0CI4KJ6YTbO4a9PiLHDAZ5
pazCtEs1cdmP34ZR3M5PdApQDmAHpFGjB7YyS1YT5jh2uQ+wF5HqrvZZOYn4znih
1cnLAQYx0xAgpj4Huj8xWKTrE5GVAGzssp67n5x5GHGvYlV4AUdzXttlpKjHDu+d
uuVMuDmsQNCRqp6u2Gx5DkYmbRtkhUypSmi7mco5QwPkSVDX1uQj/A9Mpuj8Jf7i
5FXY20szVk5Ynn34NS1VBoua28G88V+LxkqEd4kcHaCwM+9VKisNAPbEEQ2ZKmAi
Zic96vjqshY0HCroGlOwx5Yjp4+O59Nc0502nvrxE176zt3E6QWYgp+YEHJSO+1B
/mrMLFXJSf0UHh02r2qITR9Dit2p1DzvYqL163XF4UwweX9smn3VEgjkV3JSGs1y
thyW9OsyLq28IDWcpbY7UW9QWCAptMlIhPBshGPNTmhCxqR0Zwbv4tnEyRmYQcK0
DXwavCnL2Is9S/oW+yozVbtWHtDtuS2xYnat/Mx2ZQ2j+4LJ9IS8xY64YQkWMZbG
93DAn6hsTnraboUnvWPRz47Ydy6Q7uoFtD5/S/kxUaN9D3ErXKdVkLZ7fR8ne6VH
xzCLVlEFZLf23OQiJm1snUWINrdLS9/UXiuP2HGFyVF31khRoL5u7uxG6qfSbvlR
VtmKrs1CfbzTINLoWld9yhPwaf+H3k21AYCQExXvKVi5gBF0QS1KWPFW8exdtlFn
CeATbeInNe4LS7Esvs7cZnG99WBVCFDTy8/FJ6zqMJfAt/dfUx8P9oC4szYdMF/n
bsL4UXM7FVB6v8SP4s2PVo/j3e9Hh8Ti7NFZB6aJS/2aqg0uk7qVzzI0OcUe1+xO
bMAwB54trOg7Lvf5qf3KuGQTAxm47MkqdRGjF5MQsd7YDQdwGf1j04u6HwAm3KQC
clqAFuLAzHT44tk/QU7442wqs5NYH2F9uV2eVW+nt67MXlJo23fKNGyTrVKKlnLX
S+ubQ7FPejAOxa7az8PRWBmdI6u9UrMzeBbtAfN7GSYgSSt2OHB1j0p+foSEwt3T
U4TfpRLXthbWs9EKkWG2qYWWF+0+/poDQ0Rlogktm5Vz5kya+9eQUqI6YT4RVYvI
soe9EZp/oMIej3l6u/zIZnz8zvDgVowgKhrxV1YeWJWDFzQc6DlY+v+OifmtHJ4d
NPv/4kQc2D8hJP3ecMGHOqEC6/8CNe9M4/qgd4OUQIp6yOGJOE5G3BnrLOqDd0QG
0St0C6gLRFrY42Uc9xdKiKThIyU9zBjwUnWTU6oYZW0v6kWuEqmpuwVnSggk73ox
OOFGellKbFMpJwENIsIX3ytnV5oSRWnTqiuJVaCLcHY16Zicf0q5rOTDabg1jwQ3
kGWzWc4CbrqqLWQIaHu6DAAxy+7VISJzYKlwjHzVOipRagfcXxX/YtR3bqAZP+J6
1lnMscdRcD+It/AOTVPzXmIcHJ3Cb36JVVljckdShTIP16Fqn141ogvUiBpivqYf
jZVSIr986vxIUTrceuzia6AUIP3bBB5FCvCBanAUsHx3gnIajTBuP89bztC8myNI
oIpkJgbMP7YeEzd4HBI1DXLjXBdnEG1KthzTixX5fPI=
`protect END_PROTECTED
