`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RsrWr9ttIO8kCsiQklsPZZEuXRbx7czWG0PM4gv1T29rHNs07SLSm9Ve4ic3Y+Zu
0inroYT1sM03bBdwF8nlQsAFpjSQ30qcJMdAdoygG0MrqutvHSTOLKkk/COqCvzf
b3qpEzW2Xeik1v5busIbD6ChSY5Bf5AxwSYqqvMPjloBTI3Hf0nvLduU1bMamRQ0
94RjE/S24k4pre/pNbVAEXVkTfUim4DeMC/TtTUG3LveKO88R69qa7yU6Bl/UlEW
i6htlALwajyK20ND2bPxJGjQmFLgpIQ0UZF//v6MjUGkGzCLGNL6VqVvgSKn/j/X
ZN3D4XE10yaDC5bSkbMzVclJbEiC6Jbmj2YnGmQ+ZFo/RHzKbwugSOUKLq5q6YnN
7RcVcPEXxhzkiN6BuHV4LZ0FGcfCYefKB+yddYIQtmtfUPBNlTFlfpn6Ij7/cUxi
QGZ5xq2mx35I9oD2VFJvKRsknyoK3hV6NSpQPFvvLt9bXIfcpeWJJDWBPTKFimbr
Fm0s6CXw2RLL7+kWLQfEmdv5IhOM8ls/F8urrQ12PhIZvCYIiDYnGmvrxkDcvauh
JuvLqo5IgR4/VhjSgff9dLIniIUcmALUxNDmdyo1VZo41SuPyF6OaH/AKgvb3J2N
rKHnJDYRJ+P6qoNp4PCYvUQp7nZcM9GcAfk4AO1cz973B3IF573OnFXW4gzYfFsG
c+hQJIfRbO+g1nCwTht0jc4I/jcjGL9NHH92d82nxTQG2Cc7AEbpqQrRChFuE7kC
`protect END_PROTECTED
