`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
alkc53Xwf6LoioBlGp6VLg6tutU4uZYKHUifaA72z7wA3JNEWvNhp7ma/YWzL+BA
5IL68Gcsor65EcAY48bcynYtWcAnrvi2jRXboJ+lSlQwUWG8h1MoUvaJO1yE/qLd
qCP3Rz6pO1lmHzghMNxmqm9LmtC47tLlfxGHpxcuxrnmd/R1DppgvuNaMouZdp/w
hRxv0dgw+4z3f8hbU0pfZVU/MDs91VQXmIcssis8e+l+whmBD1nebIMCNBbQvx1u
h+yRkWWlyOiql/zmOxBVAbWlX7rM5ysBeTC5FnjGMlm0E3gjApJ+cI8RdLce2gte
peu+laqWVr2ljkIEDols+Llv1J5twhVeYr1SQG1gGiEbkk+/mnuch8MVHEe56Z3e
NOkILwkT0xPqlM04n0ElGVd6GrRuQHvv/xkvkf4T1Z9UJMUt8hPnKT4OIvaRXvYq
wpL093IAlATREBJ37uOfaOlppXyli7BjiEQ0EyLBahWOViWFihabXL07Rj4Mz2uS
gtq9/xhVtDq2kVg1Z7F6aLymq3TUxKYs1y616v7oPmilvlOEFaEPyeyYU3HeEbb1
7Aakl95DjPSCQgoriyJrog7Bkt6qCyFgVIzXw4cjN/iDouJp6FNoV1rDtILsOx0/
b1S+8g2SHBQ3bVS/6bvGEdVob21IWgOgbwXiafpQ+U4r5IFU23vW5NngCxSwrpF0
S5Ih8yHbZOWLwcK/zhI5pG9iUrvNYsZnKagDP4vvF/ATa+PPy6J4tklRPNhTUaSV
+knefe0yq8OlnlSV+9bphvN1IzoJYTcAqPqYnLoqSRfhwV99t1+FGwvPw9a5FbGA
E1WOZqvW3jnftU53v+vrWtd3PwCqCGJ5sFXbDBXmDZCIlt3WUFQKTSsLaCPbYIvZ
ESmsLnpzTyVQsbMJ5H3fWMG3bTeWELmesOwo0ki8tK5aFPpkSfVY02+UaU4FSbnu
Yd2VxGAesIsxncDmzxKTSM+PjfSTzhEa73CZsgGtfOCEvb1tbBssYjMADi6iFQA6
W1aVt9liLsk1Ci9pYe4indD+O6aUqm4gWSfg4LSSSimWGAhnxn2PiFs82gDr7IqZ
hcK1d9f1Au2YFo4vgGAfpujVwwSRGpt5kALhHGjW7Ku0aYy5rR1Fcz1ZsERH/pGV
7zyuZWkikUKZW2fSmJ/YJH6jqidJ18bj6OuVH0nUEdGqLx+j1TzBYOSnzK/bhI69
sl3cgaB4R2hNZSRLVAuu3RaCXKOVrMfSvwh2wDWwwXmZ2dcIXjDphE6xrnnjl8eh
XDoow5yk33oOOa7zjGHq2WJqL9WC25L9WIoq3usFjmqNN846KSrl+5BMkJihJFJc
KG6BfTMb31kNGMuMDlY02ZwPJ0fyK/l1HeiWLbJKeacs4lHwFvRrSC/sPEQ7U8gy
t1MLK7uli3PLxiTBcQS5R0oIZxZM60JvSBjKEEtQSeZk5PfxTsY2It4opOybKxe+
ZB6jvhL/KIZCM1ShHvdNJl9+DJa1HqEI1pjbR7OVRM67Mtj+C47Tpgh1uRUADeKR
hY2c18SjUTIFTDWzucsFynzXLAfqYwBpFm7tSQt5UbX9vlfnIRbZqJFZcuTR4gyb
RRaPhSRbI16gvOjdZmcO9soViE+EKtQimraF1HlCmgyJiqkGXb5b/d+wF1vW9g4o
DJKpzDrsdE2ita1A5jT8bDlppJdPULJzqY0YwfO+ilaOCMZ6vEDJHMgsLQ3+B2Wc
tjPY9vxRBVtKEovQM4Hxh7qciMzn8CHiiqsFQylVTcvTFbBymLiMIAZFpPlwD66T
mdcU2zhqFW2j/Ubf+06s8q0DKM1VP13OLNEJZUp5L5k+u8NMYh9SIhxXambwQLYD
u5yYOpwhcv3qivmR6WJ/Pd34sS/NRXPW5wqLJ9QBY5jyahvCSuavqYWZUJtkErSl
1Rk6uBoPff5mkvBb+DRuk2JDLsTYzz2Udt5N8S3uh5EDKFlnoUwo350dXdTp/Tuv
+JDgcW2BXFgIHVjusXeqkLPapLtUSSTIfQ3Fz2Ek3eJ7fOnDR3r0JrFqxRk35Glz
9eUkxvTvJ5uv4MGtwGrKJQIDhjF9yRmWOtBMRx//GZ7gTJeGBcMDNFAvxyZMlfK7
7XMxLgKKs9bm8OaovZPDdWRow3BqU5ehleoHWJZ+EqHDjFU2cpGcls1csPqFUrUf
lkx8iC28xViGLeEsi1OaGj+uHEQHyS1JHKUM+wGIsJ5fisstZWPi2xWosb4NkyyZ
Kk1hxPbdL3KpbjUpNebwJSnqQUUYVU8u1zoOf8DER5XmQYr8RnxAZD7ARtjoW4uL
pO/TAkHhRCwu1AsssEGItysR07JlN8hF62FMDQ3SnuIGVXoYtJe0as5jPgR5uRLY
/d3FhFrZ36wdrz88yjfKsE2rqmpHAtwNIYUFiTKq7U1YBWoMyt10YJ/zUfGOUceO
OEPinoG1TF5jEdELjH6+hnAP1xJ8E6nTsX/coyntCJQSOhe/qSVWvShztRVfocMZ
+lLJH/kk4rmLVtCjRw4eYMOXKphd8KqGNiI9RhzY0WsM4jveME7DusR2fg50+VAU
unPnt+0tx8EqkHH4FaFsCHlKzRIZxGMApNKPjqziSMys6QXLVmFjtxswzuho4JHj
FsaurGzUt1kYp8MExz8hB4AFj3GEcs/YagnhOiRL3GI=
`protect END_PROTECTED
