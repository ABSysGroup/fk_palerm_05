`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gH+B+FK7+FrqrGM1rxChKMvIPACUifxjGi1XTUwuX+ecNalW5qQEEC7lNyx8bPDc
kXomJCrDNxEDpImi4752zOFDOh2QG6j0ZJrJgMPOxe0huhdAKKOso499U8TPtedt
YcnScCpugxrGVjW071Fn4QhG+gUbyduMnZtu0CtAmQttqvbVDcFlQIlY6vp5UEs4
RnEoSEdnTg6g2VjUUyJRQV2ZMoW5q6nNg8XQPWxc0O0f0kptw4xXouiFqVpzlywD
J564rEqmkhNG0JL6UpaQK4nGlNCSFc5ebb5VTNYlO6HS9AUS6JGA/326zWBLPQqI
Qh33cvPcpNn/uz3fb44c+5mQfdE19tYUt85vkWcIgH7cdmnCmojYWY5tBLN+LX8I
JgYla/cRtXsMZrSSfGWYcfQWZXWwLkLW57UH9HmhrQE0l7rvZ1a/F9sXiLKxQQaV
YiUHRC0GHLQbTWrCJqyuej8Upsa08ZRrEE0REcyLfDLQSG4bYrQd4a/QMoWuAhm0
`protect END_PROTECTED
