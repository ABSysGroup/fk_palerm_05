`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WUTcsIh7PuHq6Dg5jUCjmPnHCxptg3A2BYGO/gOIFg+QoUvzFfe/Td/S5/WCLkds
ffOIbDrpp1A6+XtMH18zCz8Lylsz4dCVloe8hywcZPQoSLWXhcFXH9c+xEdk0MIz
SJG/dsqDzfZ9sUnEsFr9NBbL7dPbG6qc/G2yIRrFEAkmFWNLoSd6WfNRiTB4G6C9
/JDohGeDjgnfOpFQxOV1QGWK9r2CdyepNBwMZf3XA0FvTvCmf1r1Eow2V3/MpPyC
6zLX8RXe5dlcqF7RKiQ87bGUsrWKLPZhBhY5Vnx8xR9CAs6+fQ5wt2SU4cjXXYjJ
+37MqGskUeQmMzK9gwmgbmuz4Xrz9smsa/jHyt4GPh88ZsUhamUt0vyORnRxqe2a
v1r1bGNGV5dtZO0gZ0k00787oP/TrEz5hS1eGg/ha4kwTW2LRT7b2b0E26WJoJ4k
Xppay4a2Fo5e+WlssEH6b+R+GPXqcid0bM7FuVOmVuYqo2p3rRLDSVo9JJlfJ7F/
gIejDbg8dKNWvTDQP6f0uT4ya+oTOjxTvM1Nx40EBVX+VxaNsTWASnjoOo1Z/PRA
sdN2KldavNP+2dG5NEU5UNiIQ0QbrZwRZHFDr/LLrgeLk+72VYk7Tm59a6zi2nlF
IMFs/lItbjK6Aqeyj8iW5Q==
`protect END_PROTECTED
