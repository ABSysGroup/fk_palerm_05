`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ym6K30j2NnRNwjQEW93rmGzKZW7uJGuY9E7NnldznS2EFxUvcfCxehc/vvaCczJU
PqWz1NjKc2qUvFXVauRPP61gqs1sUyCOwQyNY7gChBVWHDPs3uMs9oMGtniiAAKU
ektPh65zJXm6FDFElcOEBh/hpSSXkkNrWV9QqfHlh7r2GxvM2PQ3/fGDUUzFNzOT
6aa9QdtIkh2MGUiUuiIr+Jpj3J3Oy8hDMA3NZLz9M6jAQdEt2vC8JfmbhuysF8l/
usO76mNyvwqqBAoqP+dL7+JU0Rx1Nm5pAhvyeeLXxIu0bpgSunAYq1bLVEdmUol0
u62OxGWhWzCvh524hpofeCdYp8aT6CFq6eGw8gkQA4ds3foWmeQ0xFrz2vvZkH2Y
iSQNeaiIW43RYLMy6WjVnHCzL9vxaeWuraHSHxHm3iUxeMEtCrVDr8xY/LUbqAoc
8Bj+Psd+gpXihA1tfLWdIEGZs9P+tZylLHoiw9AEIcODaZd+zHu8wA1ABaKMqX5E
dE/Zefbin0hSu1ATRu+8j/N/jzA3TCAuMIX+KZKG/xzewevydzgGeXbqpQoDFiYt
eJ56BcUZg2G97lqxhyIAedD/5l0ajW1TK/payVXRKau6XOulW9D9LiuZOwU7q0eP
tvNrehyNLmSAMr3SlOlOrRZv3BEbivcPxTCMbcGlgvVnxy2bbM6VQzh2t3pZqniL
W8HCuix0/cWlrcN+raSqFv9Kl+3rpMKVAUcdf+WrNcrIZxumJvTrbaK0SJuKENkT
4iBiLPp1D4cxSKs5b2w7ALNfv/Rk4rvtAM14JWgGXvu8f305C21A891Z9Z1FMDgr
7hVRF+qePb6gm8vgxX7ClBiPIFOeZZviLGiHbSWotwKkQ7yab5fYvZNxPPKQDagb
FaO62FQBh6MMwmL4CWglYzg0VYwZqsR4Q06P9NqGAnKhQJh1qvXw4X4fUOGM0Fv9
`protect END_PROTECTED
