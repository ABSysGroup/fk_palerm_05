`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l6g/qQ7ra/rVnkS4bWdECzNZ2Ah8UbCMn2HqlSPeP32itlbxfooFb0OiBNAxJF2+
uusSLWpEmpSuEGgjG+2hRLFF6f3tN353Y9csLHZx4NvKHgfHQ12eNvvv4KTQreMQ
9+d/bifv+l1r3gx34CNv/FP1+V6NGSfeG1M18SDx9BeKOAWkU3BIu7yOFhPsztgF
h6cONYRziMAvbbGkF/r6ewZRIGt/x2sB+vWPUziGRiza7lTZv3iAdDyb3ne1mtR3
GH4zVqWXqcP8GUgD7xSsk7KrE27PLvTMk25YhIQclutKqV29GUMOE5HzcYDNjKOg
qND3Ail8OpRN+DM/QoEQt3VAKzfQQiBABq9riSWjuE30NZgM6aV9/adX3dVxHpXf
pNOz46O+dRgo/HSt6eCD7CHko/pr1/gLSQSNtQQ9HZj/nPPbuZsFsfpkabZ2ygVC
HBFhnHX8XGWVwDCb7em/MQNg1bZ9tr/3zXJPCuPXtxXm7d7frMq4kyCP9BM7R76K
+9PoQfhO10KjLO7eMfiYGNXzMF51INmXhfj0+ffmArUaP27+/TTfsqUsxYZlVjwe
42jOxVc2UHbWvrRdgJyDcgAPs5MuZBeWTQ+IocaezgElfi+L7F/peDqPuFXWQ4qr
cjKdPD4Ovce4e8FEqkApcSYx38bIKrG4AaVGu8Xax2xo4dJ7WmX6SNzPZsEIyZhK
L9gmSXbefb9sVeqI05vFtRXdOoY8HQv1liamK4iEGmpXb7xFGIVDNsNlATluOBtd
DsT720CVLAXuq5dufPWsuVJ2HH4PhmoNgJonhay7Rg+pEtpu2+cngMvLfpEDXeH1
JfTCoVYZs4H+fybYlxDHJ2PgLIMlXPQ389vRY7srk5e/6vzd/+VoGg3QJpCfaIHq
5FydvtsJTLLkO9NVvia0q38fbPWdDapprzzmZ3ZH6nV8WR5IiPnCNGc/USV4r5+0
xQE5T7mXJmlBtE6eHpOtZ8b2cTmDKxfJfZp/zQg8LDVkHA0yb6MUJNyqkNIm07vz
BFm5MGnd/4WaB0kRCMM+tZLz9SpWgikxpxlPGGIgi3GxmbiBySiC7cmPWJVSpTrP
n+hcfTb65mCRYkDb2GkVQ0ALEHbEyJ6yhXwBl2wpGaKbvK2XhzhMPLh4Vi2zHAqu
BHosNLxAIlkDqhbLdYjsaRt4+dL7jGH/oHTziIWgsNeKHLucjBb1DZsQcX6FVIxL
z6yfWLyO3QAVH9X66cIkHbDexaI1rTjc0XoHpRgNur/vztqZFM3igXoHrLXO8kRc
Q3y5V9aATQo3ecKbEctM8f5FjPLpmIH4Biv6XQ49y/sVrHgwHExk3aPRuC6IEmsC
5hIqFzF5MgUYX2p77vEVssATufCtmBZhWTWWonkA+/Pb4CmzHtgTpJ+qvrSh4NFZ
fE+h2ffMFcNajBgP8n2/2Z+214pj+3i+JHbnhi2TKPP9c7T16Tr3d4hWLfurmfP1
QAt9IZPrS9T2CxcIfxlh4BSiAEkVGb9W5lmBfvKT7fB1GtqPhpKN4izJqtf0ZlJc
nu5e0jl4gpVAG5eIHjRwhQHle7bp2k4AQbLokbMzhA7EytLjPnBCuTONbrEBBu/n
97nQ663zC8VNT+WzRJityXpwXgJkI38amjO6ZtWgfq8vneQgqnsUR30awHl+gUEX
CNZ7jqFQySER5l4oBk9HbiZY+Xx0RkWJfJ/EcrJiOBKaS6H8qC1VibbPln2loJqV
s/eWCY1X0CL3hKVoaYaXOrlFIHeV/sdjtSR/0HJbJ3rwahZ8K0CthQr4p7F1UQ47
jqZsLNrqdUSZZ/sCBOOCB6TN/DcNEovKWMaOfniippdHMJxU6rBwKq6ftKon6sYz
bz/w1LZSft/xcqWk0BSVMxiLz8rNEXl0VTzZSf4leJImPCTCccNa4C7K8shefBsl
WSa5JFGf4eA17xgUKuR9Gw2WMYR4k5Mfiu1cDzOjQhRUpiUIqfqgkPssKJnnFuYw
AenmSgT6YNXh4QGnEovFTc/BOFdvoCqiu6mSPG/wIhpv3JWCvxeApjZWOiVul0Nn
04Qj1ZnpsIwmmCdyeB5/yID8JvwvVJly2j6Qmf705VJEIedoEZwpX+smyIPmR2n6
m7H3ueXVpDfvaGOB/j0O4Tw8F78uHQPxuatvul76s6jNBzx6d19L3z4JFVuY2dv0
uB65krp0k4QALUxle313kyvwcmwEsjb7V/Uvk4L9+9kIdn6VkmYXHRQKOlHPHrun
aRF0Z1w44ueyFHC193qzWoi1cmqS8Oj6RqvGNcnFKdH3T25+Kz5StV04TooNvYrW
ze1p0My/zUQ3smBDPuGI9IXzLKfg3cOzgkpMU2/tGiTBRwaFW2rDPcQ1BS/8tLOv
wa7FVM6+5cFn+zVNts4lQKPgLimGI3xjZ47mYIwmQtT8uBuyXZfgrxDfBcK9aKKu
Q6Nbu3ioHdbA3qYs94n0fmf+TZqk8YHB2+td0nHelJLIfq70aPapwl+vVqr1i2hO
ywNB3Hz/oOOyS7DQbojOx/pXDFm7quFjpNkhcqow8TftpB7eV8JQSZwzavE3CyAT
QyhGHAY33XqQwhQKrhwAVDbE/Hj1ps1pN1A4Lf99XAZ0r1IRorSkPoyZDw/7dLDM
H2kmwSWnf6LG4sKpZ82GWocnVC662aFlBv9OiFqIIoDrtMkP2zFJa6j45T1BcYxk
kMhtT0lKSqHj0YFJ0RWzBx7BqyXURtu2sTkiVaV0BufS/RqRQPj0mO9UMBZHNQJ3
nafdOMYfBoN98lN2pbi7tC2gaBI/NZmv9fTDNQWoYiLB/UUkpjpo2ypycq7IoBjH
p+l8P7dCA36C01kuC9g/VyNDiGRjK2OICUJm7PCCpqJBmyWoJcB6smEwMV18Zr59
BFlZIhO8KR3lE114l82ysXyV72psb8Tl0tqg5MFinpuq95ia11TLNblDoF498H3f
TXGcfigODzoBQDP1vDIWmcMPKkEdGmsVbVhBObIgFZPzEI/zCXjRCkGU8UzwuQhO
0gqoFehjO2nCQco+xmtEoFRHb/LT86fom+RH2On/TpnPeXDcqSdgCCOA1QhyRC3L
QMXmia4T09haLsLo4E6Ausz3grwxpkvp5JTlETapPvGFtkKdEotvVO50BSbd8NUE
DnyJTZ38KjvSHRSPoXreYgrdfVdkVrdoTx4qepuUJqHsYFLmzTc3vh73mVE3IwjK
INhiTFP374ILvZfQzkp5wW87hDVdQfwKcZnoIPAwe9FxYSjyURWNy32AqffjKwns
DeI5dKCp48KN+4Zot5ScZyCpaceNbaPiSmZjBKX7wbWs/i/gbGLQUPSExeQ26vz8
TbOUE4Dy7YAbkwqiVY/7WPY8Fi1Dsd7siXQScr+abLStZ4cDt26DGRJfw4noOgXs
jbbgbK//wh5hr6T+qF71RzpmO7pLkdTlfU7QUS1Y88kpLJSOXvVB/8PLJkycmOsZ
RrNIFRt1VTda+ScggCLR0Y+HMOFiJ+mCaS6vI9jasactAitnHIbUASOIS87EjH5l
ry6NUVTN0qN64iV7ceOGQITDm7Yv7DzlFnuZTXK6QhMdrrUmDmMlyfSUaXKwMdNy
XnroqezvCU5XJ+RQYdd++4Nd64tfel359SDZloWZ7lZvcr3AKh9VOYSdSQ0hsEeC
9yQplyaIbmD+kzk1luOxp2mG9PDAWT8v1L076GHA8eGsFhayPxSMOvo4Yb2FORfp
HA/kz5degx1uARnMexdg93KC4+z+G/Ff8HTezZALeQnP3tTwB0anIvDZ53/hnwz8
E4NzuANVnq219q6CnyWxPM9OZZLiNNu62YFd4zUgsOfBZrcUl2qAiO/AkXvI/YGm
WiKPZwU33UkLtRAQs4REjr/eQPWU/+qAdQpGN1tFnGBZgh+6Khcvd7RiXGy8+uJU
45m+AL4frPf2mdtR0Ydhk3xzNZOHgZzhUHn1gOGoqsVFNBTWSVrUIlZ/BCubiwIb
S04xVT+U3kQ2HNWDVBUBCcRQiaOYv3GzL854pPYzfiieMhhLlrgY1Tz8otXAZW23
VoLcqgSKi44ZjQ2Tricwi51nO6YC7Fkf9/T99dy6Hz/moY7L+NhFkNKUK8pHSJ+Z
LDhUObMyWGhbthmcm/L+M1TasYsCEs9E8WX5J6hUfw6Xd5s3sFLKdDWFudw2JTGL
bUituRRLf1ATusilAgC2LafwRiPkKvfzOGLVUqBNBYCF2LDBTWBgL0qiZN5YQjGO
DWOP/8AFS3rKwfCw+gZGj0aUFhjXojGl+2fDo4uvUVdLvVtwf5Z+51DuNCZRWDkD
`protect END_PROTECTED
