`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J/EY6ufCflUY5cou1ZkyU7npsV1kS3eXBuXkPGm19wZLiQb5IFl8HdKYcudfC8En
qgLjR0cDAB9buXAniR7D10ugH1pre2UIJw7L10JYAB+sXqZ0ZWngrfUZw2JoxdUQ
/PnPT61w1e3GOqqkVVyZj/pkQ+eKM1RsPYtOeAvWRDF04K7OCFreK/XeMZYIcNDE
qs3Dey3url9y06ocEWJQUfghT1bENPzk08Tli26zL0MAvJi5HVKm71zklr604WKn
ZVkYqY8Ws19krisR662+9vnBr7bm0Zg+CVyHAi/8AD9MSDt8aXsbMds5DmRcQ8hu
XxrDrG4wNEF8YE0ektv+zfseYDlSS2rrJ3eO+Qgtnf30wJ9IGjmGQuAT1qEnagIJ
FvsiA/z0M32eE5MwhdSvvU+yAdVIucz4cebTLT90daM6IiVBt8kBb3Y5q7vXLP5u
VqXzOccWTa89YVaHif1IfnbZsHNbeSoXMFD0v1qP5zsiVQhTplC2W238EKyzYfX6
wQEgOoFzbA7aUR5rS1xbH4+njgiOXW9Gq49rLm8b7fJlAgYHmECDh1LftJs+Umy/
LgjOCYoWsl5GNIwbH6NFAsmlz7skeCNRP5K5hg6r+N9D2Jyxt1FWkfvGEeHOTi5E
abW70Hd8zgIF5uwFJa+qtOLAGpYZuC4H0evPpagndkWlSSKTcCfbrIryR0zoTs3x
Q2Zed6RHDw2bGdL7NN52Ae7p3JKtlm5WlIcVsBVMTKNJC7OAE/HFS+hcw/0nFlyX
z3z2vTXxZWNltL6adp/z2A==
`protect END_PROTECTED
