`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pRPg5cv4ERUePeCbVTlFcs6XUxWfNmsbb6HLUOy5x1U8w9P9/c8FcNo+LNQIl0Pn
bWhjK5IDLI/s6ZvlsPVFXpFDUdpjK2DrFreBWXDrICWtts/JGqHdtgBblpNPsmte
YeLVfPtaPPTcQK3SCWQFC8uj8Aee8DYY3ADnOqlygWmOfwFfTrE1llLy2Q8L5uZr
EM2b6TlVf7MPXIyGmcvYtvUmfYS4xhOQf/gXpzeeAXIDEo3KSnC5JloJZEReSDnd
6Std3RmG5Sr1VRVhAP8dPcBUfdeBWaP7zZDQl/uKyHfoNAvqN2QDF4NoJ1TW5VoY
`protect END_PROTECTED
