`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5+0qS2quXXqOl9145CtYidLOiEOudSNlkR4FwgPVUWJHXIeJxc5nEUVVLm0jE/zf
GRwJnG8CinBTQ/o09WT1skxJO9OknBgZW4igvFWeIBztY8IN8JFB5cckONjbwG16
wDPsND/O70ZpR2ACy+AeEktXTUChcdWcAZpk/2aEIAu5RYj8AHx8XrWZqwYFrzpQ
VlUz8oiw+lhWFd44t2VWAkiJ5PXxlh7bKrzs9OghZ0tUSG1eGiLV/Ba5I2+x46yI
7ejKY8fVZv2NwZspHLhYkGoqcrKgpwTFeQWZSFvzrz9HC5W6sIbA9YKXUO0AqI1a
aQuIDNxQcuuPCsG/i831dqyISIlmHv5ErOFTbN0B+EvtOWrkXeA0A88NPV5z10fK
bIWExDKjeJsgtolFIopM9ZFzOJTvF2qwT/qUvTiANmCK+Nfk+qmVdCiarEGfHBf1
1gz6WJc3NTY1RxbwzP1mklpJB0VG076JyY2ESOUNRsEv0j/kV6Scyd3FpbW4cQSb
XDYYX9glYuRvl7Lwbk6aPtAKBSpilqsT+8nEjKaSPVatgpyILWsm42zjrEpbin23
JoaBMA6FcBR1gTpfI1PCfynwSm1+FrC6XFHgP9Oa3K3JcttLB+yjILJ0GvJdj0Hk
EGQpegVIRR2Dn7PeaLeBDua/qf370jwnrZNIt4OQXdiekJThiC5+QZ+woOKGCiOy
/J5TmvDqMXF8UT9ct4OZfmp1jlvrNwZPgwhwR/zdLjilnhTcp6d1XvFKgwr9oACo
Fy0x92gtC8HuT12QbT6zCxNAR1YAnOpXUsEIfNvAitT0IotAAnQC3z3vNjvMvMmu
bJAgpL9G6kGHOrPV5uGH+0JUifXLd/2K///GO0CzdVBVXpViIljglSssJzMTH23j
YcXIcxXgkCXBLs6feaXyICp7xiNcU7g90wzGLZMG0r95EeB63rl8qE1aI26a2tQc
CtBhHQWPZlFrUyukAgJGlwajZ3tpjpnBFxrlR7kNC7Loz764LoeaNy1rjOoQHjPP
FmmRGFoMBgldGIrFjjyuS9QeV74zCjIYTqikxcXosql0EpulMKV3higghI7jFr9x
Fy7ioS90zeLmNB2RUHcsCfv7M3xTrOsj/wME3A79A1P1nSxQUZjxp1agwuSFq0Pr
Md06zryZrK+Rb4OqfAIaEc8+usxxESDDd7d0u2sqmDoEv0G+e5UUi6+nZJ8kyDhH
Ch4lA7ntqPQvACcw6CoO+KmcxHc1lrfQCWLGFPwlDw9BCskfJKRGW/dz8F7o8IuW
lUaLjyBHmsbZnFYaD9Nv1FgB8BVZx5Jy+5inME+jAep9mby7Bs7rNP+Axc1GqaSB
s3nN5jvayDRll6LaAFfNRFqCyYxUaPHjS5nOyy+NDeyL9ps6tpGaRUOEtX3KbSHj
904DqIEK7IL5S0Wfg3fY7FJ/klmABfwwgo/L0fll/Zsr84c51naromaIdXg0mUzx
xll7n4d43NbLvmoX2kx2ZrqIq7C++V6ZymxogSP9CQvzhku73J5dyg7re/zVQtdJ
yZWD0nKJV9vJxxIr9fyM1Wc3VQTCoXQJnHQwHPpemEKwhOqf2BgNFgmCKvhKzVJw
wyUi/COeTaOTLafBEiNi47tPIuVDv3ZOiFo4yZthSNK0y+8WaQGv7aHII8k1WsEH
lkZzDzZ5r6kqxlH0KDGrSdXVHE5B7A5jsjOb302Rp9v6ZuCfvG9EFqshd6EacKjf
O7BYszI+qxnhcJ2gJLi8nfSYkeJMXeQP4m0OoXLs1NVUVmMNLwG3x2rysZGu/655
3sHEkoZete/pCRQJd4Qjo9NXD36dgC4JulbrhN9voBDhUkrLnFzx+1ZpGLA27m1t
k7c1GOwLRReBONZ0zAmlAUNPFujqE8jWa0VonVRFHgyxqkpKdwxGmuyG1ZqoT8I7
0msqDlWrOpJWHe0AFn1UQfibN7vSGG1lnd11mW0MP6DZqwrDGWxyqAkn6BHPfpsN
WD6RF9xj/qm0MCnM0Gw5IOe4aNo1rjofx9ab/wyVoQlZohT+LZaNKlb1FkmZIdh8
Lv26lLbyhVU4y25mfaekG9KAwaAnVgATylT3OlzJg7ew/vKnLteqk+3/izWJ2Xzw
xEwx68OqBQEmTZC35VYdn4ehaIICawwT324qzdJz92R8wrnYYIFFVed3EWKj1F4E
brVwecmjDgBj8DXsVDWxApeXsdHLGZNk3vXKzQPgzNsktaDZZS3RSNzRv8W0kiF1
jirwiNf8ENK2yOJrBrtoT+EbBZzOIqXtFtLpRhil0VtpTTqQJ+vCxRWxfCIWMhZD
veBzjv8oIoU+Nsng5MeZ7a6M/TIXCRRTj9hQ/1urXzhZQ7bIRZLgWMHWNVAnbPHO
3VkHPVOp03kIvNev4weMB70nSAu4tzH6ZHOy+l7L4v2/gij3giHsiaEvmAt8zgsj
PPq2hfUGj///xYS6w8pni4B5QSbQhLLlUKD2tYA/0PTBIAoeOYd6/Frxdg95R44b
5+mEhjF3qy9Uw8PH3EvorOqLrsys3ejVkfRiE42PnDyeoMhylYyx+wE/bycOdbZY
95WXbcpf/Np9EF0boda+NcJnYCzDiDisGm/YAQGrWtySOwMxGIQvJ8elUePad6el
7w2mDCrd1Hm0nhJjeUj62AU+7hm7FApB6sEdtNslXwv9Z3u7t66hpep4VUmZLGWD
yBhpCYLBEmD6oJSVutnF7pw2ME35kzTGAzESWf7lee7Edi/oSOKcs5URvmBq/4S+
`protect END_PROTECTED
