`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PazZ7PcC/6rKEVJzzkVJdeiVJFv3ih9wk7qRhEyMKyovG23gDXIYKbY2sGLoub/3
ktUN/IdOAcnuRuWYYp8CmAU/T1uVQETL109ZkFd/lf4O1wxXUdS60X7PetiJ3GEI
tEuWHnxHKhM0XM1GqZp80u2l0wVncDpdwPxosAfyR382dfSpTAlF/WvaOQm20PXI
fx3hT0ivln/7KiA+j1eVfILxCQZGPWyaSR44Iq8vjIc7cDJON5ndOSE2fhG/MqEJ
dXLa9rXbWTEDFsmw9c9IZKHENWTEYt1Ly6gsGSzqjgaat8XuGCTAu1aCWuVxuQZJ
bbq/FC+syVkoYfjTbVaPYVY+0zPNCrPYLbl8+JFXRlfUrwFeKcsteDmjzOUj6uqR
qqHf22y3lpET1bvAg3VbaMegxYnSIuh7Zu0ozL0p+YnYjWRFeDdRpTCkrk/POYxQ
FhrPPyCTQombDAv5Aqd4h+J7OY/JVWdxliz8xWkCBo/Ep7qI4aOpi/CJAjvX6H10
Iw4X7kBfhE+7GbXIwh4xg1D6RrvJxN6LjK6z8QMNt4VFoG2QbdocCGzyNnajUama
sRsWav0Rdsr94/DOkjLp1r1LZmQ47wsdlgZSMx8/sGcPle2G7npctgPq5dJkvqFj
R7rYb3ze/12rQjSQcDTqdsNxjL1BF2Bu591H5YLox4oJe4hqKqcrnqDGxXJp3DRk
45do0zxnxa1mPppCv/1DuOQpQ6WCTHaE5UhheOn2/VPQZzFKEct9nbUMv3uLNfk2
jF84gUb7HpJmi6NwjRGZQp6AzlgXRRPGxuqFyrKr2bfcZPUXi8XKJgD+Qhphy/1i
ZPN3bntB+8S6z/nA5ozjs2Pl/LGmyrR1uIZhyT9h/p4xmgyHZt57aKtr8Zb4u7WK
Yjg95xeNmebvIb+z2l12PSBMJjdGr243N1E+Nfpo+YT9MfX9tWChyYrtVB+MJk6o
/gIMLIbAJjLybqFK4WGbi2aD95mR1nEXNyg/BnUtgKr2BM9UJ+/M7MOUhQRXBy/I
DEUo5dKPVAzTCAoLxc/pwbOPwI8lkiuHbiNvitg+IIBy/0GGGjx/Ut4RWthRpsV7
x/BxEbp4Y0qBJLqAVjNy8gDAmJhURwKGBXsNhbJZCjBNa/GeqD2fGdRLZSylxWL0
z4aWsS8CUU+sqJU7G9PjsUFYBrhivTmprb+QVnQ8dEM+tROMv0nnYo9l0KsWNoSX
u8+xgooMnuGvw443YWNhOMwWD6TYHqRgVmXxzPd0uYdEeGfbieCEL+Z/GNjms2cz
t/29B6QdL91LNjAhJrploUaPCWvMznB3NC1ltoU8aTbcEufDm+0L9IUhgYxepfzs
tn1Aq5JxWnx3ENzSPoM/J4IGcsVxV6WWsBUhKwdW04+yP+mNEzETwaU6vSuzdACJ
hxutykyUMVL3IvrsOSNHTJB7//n0BQjK7J1k4rhXtMd2Fr5m+5ANG8P5FCjdBvtU
sgCH89H70qnt7N+Ox+Kv+NIIDMNIFp+f6RQqTdX/iCKGaQkNjSuJsVu8uR8zqwLF
PogYwQyTawMITwd7G4prmrf6n9hBIuBaZETZIVq7+NNWZG+W3+/ntWwACWFG7N3I
VPxfyh5sNw507Zq4r6fQ6GrRfIw+RlMuF73+k7TEJS37HsxkWlzkA2AlWLO8Bfad
dAB8EoM7bDaz6XFOOIDk4WwkRoDHFjQvDgrwwxdNPvo/v6kaoNKtQ2DsiFK2YRw5
1TD5RbCo6DPUmEvYc7kvTXWeO8xcX3tu3IaDJ/3wbExFxE5LxEJ3Dpxe7hA/bkXx
P1P/I66zLL1mlbKqAjWTft61qquwF3lS259Jb+dutDTpg0Ugfwh2aSbGkTYkIqIs
OwTeRL9DmozKTzzQcXIc+7xYw/jBMFYT+sFcMvPSK0MmdOayaJb9dHsYCHxAmSKd
D3zmnSk4nYC5B3jX30OOVi50DDX/5pV4HkPmmtSu5LoMr908FKZ7siMHiy1+MYJq
1TPq+matn1F2Qsnbf5ZOSYMd4Yh2dfJwGD2PVIRV94bcs+UUQkFnNksLS15uj/9B
nIATH1C3XquEcaT7UxiFXImqChmFLojyD0qhenZoLGwUBh9BtX9p6VgbOUxbAiPW
pQoi5S6MbTZj6SNyMfjdiTzu1qspS+sZj796C7n6lrfTIz55fVUP/dn3OCA4NjO+
ZnVlXMPmO8M7V2Oi0XzLOH2gGbutPd7xo5PqTI37pE6H4UBcQSwZpGWbxixfCSeJ
spyK/p6QhkfWLqsBQWrSOlgrEHmPRbRpB4ApozOrM776mDZA3iHwTE7DpyNc1RV5
zvIVPG0b5u9jrzQ97n/rl3e8SmbCjmsZuamW5QWssHL/rrezfD+2H7SOmToEcBya
ZQK1cthDjec22rsBduGgnmsh/9Tsccmgn+yynHMCl/jp7YIeXpOjMQIHGWLJE+9R
S5c4IEZ3Cx0siO0dUzj/xSMQldZFj+sP8U7otCHEQfRJo7NoueHu5QiQ7uzcTPeE
bzPeNfGcHpCLRQlzCVqdvzw9o+coHdd3gqDk8uEwqck0KdXjUoaz4x1UJM8pPbpd
WyC/ybP14Lm351aB9+Ky5MzVFtYHNLg3NfpIkm5h4+YBiTkU3P6KCzgV7/sNFNUq
e2YOavdF9dJTe+shjUHn+1a0mECm1sdIyy8X7CdsMWAIobe7WFF/pBTfQxLeUJsi
vpk4gIvR95Xtyyw0lzr+w7XgzuLEpzhteNK93/thg2+rJexVMhtsG0fELRTAniyM
KAoiaFhD1XpDrV44lAnhrHJgJvKBqvqySRQiFi5d+U7D4755VCkIn2ysaeMmTxfu
NHB37TlsOmkOf+W3p6s6bGHbX1ZRfuqiVZ4mTqTf5ybUmD8AZnJyzNf/2eDoTWhp
0LRnAfED9+pJ4Wqr4LmIJqjSB8cfpWpUQ6iil4d2syPis85Qc24jhMJuB96c1SIr
RxUUySDZU+h4zRzaFKbmsLYo1XRcna6uBvZjK4P9XmarC3Gl/okFLCACKSjQvQip
xevHIXc2NciwParOUnUtqgiLHk7wvil7zNOsZ49CdXy6kujBRf80lEPLsNuiu6yL
b6cMkOQyix04eVC3NYGCQcb5dR0C52pCU4Q08QJDZqmJxs/HKzLIhRHbjlxbQr/f
jcc0T+EPsECQ3LHkdg2QA8Z9zSE/hTXHE9dq34eim2yP+44N2Ft+6a3tt7/p6pVS
hZWZbnNHiGJ66LDalFqN9149QIasCNyAqIRr7aldl/F34YdLtXTHRzbXHxXx8Dfn
Kwvs56CkQPBq6Da2nOQX998tpAGRj1oMAcF03h9fluGY1P8MJzt5mR0v3l+Q79lD
FtkJxBw/cvxXMAexNXeJ1lBWlTy+/jeTj5SLM2qWIeDqRPhtRdUeYjdopNWLZG5j
EqWnHYyeLfL6Tm0eM5hihl7GtEz6o2D1bVHxl7XcSg2IoYyF6BSpq/FX24dsUhdi
Yfzeb+8CisIPW429QDIgkEgc2Vn3xwTcHl0DELX4aT278X705+8GSKlfgxwSiWWr
2/FZ6Ok9ofQoB1ziYAPO3+v+n57uUKSA/umXmTfwNsNxBF/CZpmfi/6bMx7AQxws
OXSfQy1DMXC6DMYvWCRMfkztv3AypRPUXIZQbmZoHStNvLbVtMawMkBEG21Fzv7O
50tqZozEEEqnrp+HYJQRDzBgTl4nvrKT52coyyo9p7DO17IrcenPSs1aCqWqQHmk
gLdgw7wVYSVkUElxFIiZ0duK1Cyz7FHiUG9euAGiLsW6NrMwpVJJIeLL31ajAfR+
dV/BYktMPf+ZhqNo8j0wg/2Dbpp2TtTZrnaKQPSfK94Ld5Fd0Kzf14uuxzpC1etQ
HDA+PO3CuGggcZHZ/bhU67Fb4an/gWSMBU0ilMSN2yv0XdjeBJJfiarJWk9TrHM9
glE6SfTJUCvCqfg8k11zK4yfrTRo1p0gBFXCSFzk3UWQdAFar431w1AJbcREINan
T6A4bzfR2/KWAQ5LMuidVYjYcoKfMPc55xoZfaHbXSyyeurMzTyGmJo2Nwo/i3VP
FX2yRjABjfRkmXgnhmWF0SazEvX9qDu/XBDou+8A7zCVfW5QH95xcGkNLGPM/GiG
Edl1pQFJqlI46/lLpz7hXA7z56ZRYZuVfvkqK+hOsiIdxMjJwR4Ho9KoXfEVPhG6
LLMbT1KwOgOpkH1/zeleH7G8wbsRD4RCFsd575eh5fq8b5XaIG6GGAr9wzSCxNYm
tI/wb4nmjzzZdPLP9FFDNCpF/RwD9Wq8gZ69RSISOUGIn3zCUNvhBoPL03FOc4ZG
0URj6xhrd1oDuU1GA8z/olPAt7IrcM7EWwBbkj27N3ABrXy7QgZs8ZfkMIZuZBqf
xO88ZzlCKvE2rZ9feP8cqmJ+wdwl/FhPKb3LF1J4JWSCstHG6CVwe1JmvdG5mW9f
PGE2ujn5iT1g0ca9IP3fa5/U/WpOczwxXixk4goJalSJ374Uv9dg3hY0jMhK1kPh
DzdG8cVld/xgUx8k6cWe9NjD+KsW4dDY3Tzmw6sIeWwmGaU6g/TUDiGKgB2cCSqN
wf/wBsNGuHkSNKE+REdq0ExT+EDx21TxDbLCFEHiajo/jy+chI/kA8wR528+8ij+
thfsJlyfKawlGOGojjPCncaIR2Iu7pLGQ0P9wrUNyPlZlvRYehbhJnWdkPIjriRQ
3n7sfzWqTorJ1RQqCGYqyEO31/L/lYqxpDYBlMQiVy4SMYNZfzh3fHAzyazuQEB2
hesqDqxLwGQz8w4kkJA2uIgDBLftPzfqInYO3J3Z9J6eiYhFcNj3X9bJLrKtiAIo
QEUvvs1jeoLVa1EDBcRRHBZkrbQjlKQqWdJp5cMdLcum9v3PBSpaXbjsmssXy7HG
HaPKZr7nV1b3orcy8qF6lh1fRRIzhDAhvzlnxroYO6cF4fXyBjf+WaEyTEWiCQfH
xU5zW8ce4h1RdrsoYchpnetBF8iTSmo6OAtfYWxtEwEytt8qy6cva8M8oa1vyIuw
8NzGUns4eoTw+FR7E3h7Sw==
`protect END_PROTECTED
