`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kcby4jHxaHaFJ/M19hZ4aivK3sfPX+uoCtCKrQiamJu2+VD/LjF7ZuNq+w4e5A8Y
4m0zG+Qp1Ksv8j6wfsFSSs7ahQ6pCmcM9VS2zRb4tOikUndcl5TS5FRTPj5dMjno
XnO6jVwmL3Nf7AzVjZTnXu/mkmrHF0EAAbUNj7ryUn3q1D8TCbkW0cCgJ5h0n98K
ZZ2PCtaPw0O5uHsuV8XdZ+ASDBJ/pMsN8NFYp1XSVfN0KcypT8nWGnXivdQjDLUM
mGC5FWkIIwYMXwGBDR6Mxipk5gueO161Agg9TvX6NnI2+afE/VvsOZiaYxXBpPY4
wjAJxVGrdubxuahmeyYtpKkqlGhgEmEUXBmu9dKT82MCkTfLdLbsxlaLLMzmedC2
eHLdMNxtTjhNbsm0FEVNIxl/1Zo/K+JNSHwKmQAmE84Q4862s4ORF/Q6e8sHICNf
GXf+5ndQrYV4yWYlvHrvjfEHvwV9gd3OEL1lxbM+AF62XlJItSsTZ/QBK/SGdoS4
FZhUURsgpzqFXtlpfP73kp2glLalklZADUJFFClzWwZwU1wKL1NhuFrRrdMwyjPL
tioa4AW0QEm40+/St8tz+ebUQTieArwmDkj4u2dv3JiNrjHowL0usrL9JHuJdlU3
z8t7Q1F5gDbOqx7nnnXyt+JMjkZATqeQwThou9ltFgp6mkb2FrZa/wr2Yi4cQK92
7vVrTeiJMKPLLtf11q5hqfL6lux2CXgXlQrAwNdbBDr3/ASjrly+3TlXTooORE7Y
F2TuE1BnKYO4qhAhOizFwu5E0+z/BsTefWYm7tWF7MltFe3h4VQEKJ16LPy5CjXT
/LwylRZLsvQmWAUOX2Pr9L/IsuCzJYHtG1x2f+7Ufo1nXwgUOxj3dbawum2E1XpX
/h/YqvTYSgO9xMfLXgW/fiTr+gD/OfxCP4jq00y1dh9dsdu44lQ/KHnwinJtb0lu
eHkPXeTeds8b8F0vkzS8l4ON4E7K1WJv+7NBvEzRd0+AD2uX22IJntboZLfw4tfP
eADyAOOlVEM5uiqOzuY/p2IC212VMNgWSM0YDFOUBmf6dVeivt5v35RxbU9476CI
xTdVF7CIlowzSwjUdXMHyR8RqiC9cRyyzatuS5vd4tF4lxBiTNCzfSC3A8u2vboI
XISuf9frwcb0pKGsYyIFGbtFW8s1niwim684P07wrqA4fQzwkvKkQbHEZgQXRlUY
PfHUWlO45FaeKBBkMkzKmIKObFSJ6MrxVmQA9qEW8KrXEHNCIt9nhSXOmr+FgAVh
ZOqfAt8v0NNSElqP7PWusM0awPO6HAJ7V1O3HvJjnM901G0BX7x1J7U9JooPHQTc
61E2c5uBYzEroSx+gq9XhmbnwCdIugfof7zhhB5CNC/Ck5M1Sx46kaiCUINZbAYf
wZM6mv6kXAleOtc0o4QNkSBDLYgM1ydZ5P1K8IMmRwQyAJXpW5bpUThVtL/lQUPP
bPbkKuHPHQs6Sqnq5RA+vWdrYIVt/saYNhVLhQqfeAUbFVEY/u3oLNG4Ap5I/H4P
+91XH8ufdGswu7Oz8YZ6QZbRC7JxrHwkImv9pcyFsgJ0n0UFlpfKR8ndYjV1qjDk
VJxs3fMOidBlFvOt6DAtngyXr7BmqbtG1D2A5DiakvEzj8d2QI3V9g11SLNEK6EA
UwmBCoL85M+eYGWcynb5SIEd1skFbC6Vb3Gc0OOwgH0NDZ+MSev2SQB66zWF1LXY
IxDOnveT6271vk62IspUxFSzukw0ZyB4TzcRXjCCMdXaM+88z1FFIyTpITaAoY/d
Q8OCwnntMjerSzoKCNrbvj50GaAytCp7+FiDtekHsC3SQ0YleT/WyoQOCepTS9EW
XFVNc1ef7iXrH9xLFnrl1XF/KZjD0WdzKF/33yZZeIcDDAMz5Lg0G7AvYmBXgFFG
2aUYQJNu1BCVa7UICmOHI7+FW0BVgKTakKtg7QFfnudVGsn1eu9hF/u9HYSPgzj+
mKywGD3V2c//R5jeNZ2yWRRoSkGHZ+7ABD+MMZLwEkg5SoZMQ6tL/bnMY6ryogOx
ldrAoRi7FnSmM3MUEfM5k+5LX7XQtoWEqo4QVhGIXwRqP4fr0wvl/mm0X759KAUo
u9bG9O2CKvFRo/VDcJOCgwUs3utI84mEGz/eSLIJzEE0IE2W8cF47mjP6vDFLVkr
kHsILDsMqcU+IXgNOwPZk6HRPWXcXuT3vgRPbxOrUT8VmNHk4tTyg8ligiA8FY62
mthzhkmg0xT1i91iLQCNJZmdtmWkEeHQtApyA3XsSQEwMKUtt5ZkoVU9grMNzXsR
AjWERx2ixrd7VUgsOldelIe3Jt6ajyHi5Pr58/sBoUbUMHiYfH2A9baqXKT5Kh/W
wuO39/zR6omsDgmhiVB1h9jGrL038Xx8B/RQy93clGkzr585p+yLcuPbmGuyZqGz
Y6Mh75bsdB/qF35Tu56evYVscKYo/EvTUU8JxKCKLTcRAt0QD9lDRX65L67XMUyw
0VfZzAVVUvGKEiPhyiTSoj4RL8QKjcuPn71fKwmSdJ76Y+ihbWQaELND+6/rxCTl
0hjCyXzdPZYXGqfYfuMgHGS+3VhOSRGlct7a7NdoP6c979ZZcnL1jzMb3rUnNBpp
BRd/P/9hBHie43SShwlUHSCZItjE3DTYQgPWcpUMRp1x+TVjWyulvYNH/gjyckh1
TyWuCCKgQhLRniEYq+prN+lAzlWf3/h/VcwjOvM0HRM7+jdeqYOCHpGkWEXzoeRh
LKN4PJTchhysrme90Twu/kAng1c3DproSzrTyGsoIFFIrJH0AOp4Z1NDvBf+Ngva
U3jRHTE69FQyfQQ0+btWpxA/H3Y9Juzeo9YgKXJYiwXv/URIuf/6Lip2Vmd9tWUJ
Tfol3adgy5VM/N4slblL8LZj4OIVb/QCGXgfF4scw72fn5vhugKSutvv8Hbq2Z6P
f/4IBvOcdxDIxxVGBv+2J9frKv9RpYWq65NZk7RHTdrb9ioVf5ylhpQKHzqSzh2W
OxLw7/HIYc6wccOBTbDS4snresTi8EW0LHx4aPjgsDCScPu3GTUaJy6pUfb//RUI
HQxwSIVLwuQlz/TRDa1leQGm7rxuiRXdC+f6FnR3HXEvSQP2kBOF2P0aic2Z6C/j
9JlK1ZASri1Uv00/tmvvD/ggaSi3SGe1dCmDAQVdaZYaL6VxZ8Esdum9z1Bruu5G
aew+oJHKssFC8XE+bWtXcWdQ7Upq+Zcz5co70EcbOJkvZz4JbBArERt6gSsRyNrk
LyOD3ML0yKKRyYlObcrOfnP2SX0hKR47I369RwFeNVa7M34pFaPqbLKbMR2PuUqE
s6nAhIlpE3Fvq/A0bjnEjmwSPEZklt1/y4E2O2BRFcQOVl3neKs5pln2Go5M7emz
522Ju80ts64sxZo2VJOaQ7tf5bv43QHlhnKoX52XE9YB7hHfzkbv8OCZ53VUx9WQ
IIyxkUvGV2QKUo4qV5Vm2kc0V9O8ESrbJl6C1NaMANN32Qc8yMv9yjpbBWHo5a8s
AX1rd1U3S+kGi0kDjF/U+w==
`protect END_PROTECTED
