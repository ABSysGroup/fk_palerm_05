`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U00GrSTv9c5niKZ7J+qcvFmp8eVe40cql4RGevX/wm8frgqH6/fss3QnYYZUE+ZE
T7zHCQZoOrpuGnxbDkX07H59mt4+YrRVbHbT4GdUiYfr5B3hqoHVYc1+OzcndnJb
hXtKQr0zL84fRMQTJWPZsAUJRn7IGHN/sDAV7VZ+nNy8zw6APMf4djKoLx+Jyd8k
jQyfxfXTjjWGHoe1d9h2fHxLDWS1E4jPCXIIuphRCYiZhP9vyhnFw393QhgV+9kL
M5f0Ty4n8tu7XzPSWkjl4FgNO41/lIkP0LX1z+3vtW8=
`protect END_PROTECTED
