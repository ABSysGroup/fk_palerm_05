`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hmtvx346YMK8AgEFRJbKkHodpxZvrsAmKu+O5fpn+xSQWp+3W2r/EEnLCDz9BLI4
nuc//emWsObx+kuz/cMyVOtizkU3fQ7GDjgnsz1VNlxrdgEM6GTlBqhJyAk6b4FQ
wz530QTmoJMoVKhvrtPAlloqK1JPoO7O9qPTIChwaaXlZNqGYnXpf5A/OkpAfu5r
R00FOTwT9J2vY/jv6X/LvaIWzyiAKdjxVfYcoKsfmYSSGM+QBNCEpmBe1Slr5rZv
3m0EaHYMaifmpLEsEL/6Gw==
`protect END_PROTECTED
