`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3FYrgx4TYv9pRALdYgYPwgEhEVVUFxtQHNzKerwSrezpZrFKdUlb/oTzzir/QTJW
rgUvONdURXEe6hkpaE59z71HG2Auf+s88jJV/w64LvFoxUn5vvY8bQm9cCAhR2v9
ebAzbmtF+E+c3anDCZf+ChUHofQUcuIXUhPq9oyQaHAnmLft6OV845yfhNTPNZGT
bFA/6nGWSjHKp19xv1QnTz0sdORlEfxAKRkyo+khng5m69FJGclrkqWlaMotbmyH
tKOQvPQEyIQoY+KtVsXF3+t0YHwmmke2L6T0HllcxYEje/1FPCWeinlVgc7+2Y0f
NiuNP1FpdEENX2fS7EsEZK1z9ASS1jdrSHeCwBmvZNyeSGPQkBn4TuPrytEYS/RG
rMFUE1zC4f3xHBDpJConWnGUc8I4QILvsY1yZECUukYfy3WMK8TOn2SJKrY0vL4i
WbVyeyLnFtFoFE9uqhGHYvWWxuB1F8mETFlO2u8hGuMHYhSIcYTYO/3cOl4FU7zY
yhDjQwKE6mWJrUlBvLT3u0rQbVLLkx55/f+gLSb0OEBUK84eOw5Qf1cxQpuGbop2
W3YTIjbRGAFjuGo0EooR5DOa2xAi5zMLCA6W7BucFpJxVMFjsRvCd7iARU+jqf6F
rxClvpHCGnBLIBoelTEm1r/ZToALSNHYnwsGlbzi4Gl12RTt35klpBUnTCHkScX+
c0gytxYq3q8EIbHg+5L/jIiTrP2LmY7af1/qxlle4FVhQQo08alZtXdg4e7cB6X4
mnHTVe+KaPOmv1WuumCJ2dlnV+Rw9dEtfWJH1mCc2KTjQAfBCSsIm24l4Dhd6zO/
84cQ9wRjWs0WSG8u0S48dURV8Ps7xovIKplrpStQSGfimMV+lNMSJ2rufIUnzodl
XclTFKIgm+Y83D3bXVcuKjfeJN2HYIL8KMf/M5tdI3ikNK1DqwzP0v36bUhkj107
7DasmTSzwdxwPSRRite3nYb9piqOHN1AxaQDxuaUg4TkSyOVTxfGnQCip247YlTY
5ZqPWaoHmliibC2HPtPFk9K8Few3mAz4PaZ1+JT2vkfo800/RfweIM3BYR7acSxK
NoF8boaKrrd2b0ONxbqMZyaACpUBJWuoh4j082AoRhmIoGhCm36goNP1CZ6uO8CA
mNWG4uMuAcLRzKSZragAtxwVnFSN/Rmvq+xWt5zzy2EffkL2oIGNYhlINIi987Ct
evVDvNrfc55+Fmsxz8D/m3A79BxKWRm/3FrFhp3jBYA7eEBL63FZXcV0VcEJjpDy
d+j4+uvrz3OAZdOxkQb+SbluvfH5FCIKXNXFdKSQo8/Exnx4iSBzRDGa+1Un4qtH
h77TSi0S16QVmoz4kr3W0lGqNZ1ShMM1Re5LmJv6OIOXvvqPIJNZUrGVpKkNftqg
lSqK8QAjvZX0ZfoS+q5+ME41NEp3Q436yh+ercybweBJOhoeoDQ/FlN8fVIm2lO8
D/00pMEItzlug6YfeDrD87JoTvuU5P+xMycjWKOJH4M5R92YzWny/q//tDGy24ll
Atmbl8jDpHnUbz2/JA/75SyEDe0XeJnmAE78C23RmLEBSmu6zunFpFU2SETud5Eq
NxZLok2/1F1WC1DrvxRtBc3nPQqrrAfswI5dIYTX7gZ6ZkiHN3jkjt1wlLId7yK+
MmUv8E2L2+7GMZTm75VHfb3JGGsWKxCLzPfsC7Z75sn+oL4CgvwZlzoEnm6b4+W+
hzWZOFAaRitsFE0N9VOKXG5eBdIjusatPSvCYwZWMSOYRUvKXGlUChQ//rPZsYG8
J8I+gij7ZIU84Dw9RXlg9SyTbqhGXH84bRBWnQacTYxkkrAydtwq3Yrlek7iFr2s
ThXP6NGsgLaWURbHLOUirVDL38iHAwukxgaCH6PgaHk=
`protect END_PROTECTED
