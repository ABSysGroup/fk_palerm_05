`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZRYYMLOlpUg0Akh+0DGlekRZmEBypWi5PGcL+5iPXUG/k1oDvKPAcelNuTDKAcO9
jgu3VZU9TnA8BCBA+9RGKgc5/K9/KEN8XwAwF/NkqA7os59STS6EDWHuNTx6RxZ4
MZXAGnwggO2NX20h+Kq6Z0zqNTdRhV/ell9+9Yt97ekgA+rDCxLWuREpp/UeKVRu
36JMfx0OPWww0k9tlG09AF4eGBauIAm5TUIghYe6fUGgwWKFvdMkDHMQfkvy/2/E
ldcr/HEC+AWItRIX3+lyDhAGNdheVObTTnlMNhiW40khJ224aM5HLTI58S8wUEQ/
3J/d1HUjCVaMO0bQTqA3LG4HIU2lb4syAFFv5iQgG/OVzvZXxZEVcNuOv4GFOaQT
zKTCO/HH5S6FIc2mD+2JrJ9rIv6gmbLyTOc+iHJWhfhO5HWvC18c4kDhZVRfrUSm
OYn1Xv3SDNAyPUwGZFcIe5t40jqJ4S4jzSwP1a+ewMGafqDaqhzXDFbXGZzSNk9K
zFhMERHWbnAKYpqnzVLF9uPNxGQHaQY2hHgEar+DytgKYSy6FDqCkzEWS9PaEl/1
`protect END_PROTECTED
