`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tnO6ZK50Rf1Gb3X8KBRt0mD0xxS60llDbpnniQHHcdCShDu1H8xbXXtd9i5J53nk
V+mXcA2fTfLXERsPNywntqAqiNckBqz3BogRJmk1yJtm9w72CwSrjk7PMRZS3ABe
tMWRs3mv6DYnW821Hk112MTBVUM76tJuV4H9T9ETeJVsWk0z7Rh1ETm1po1xNY+D
7kQjRznehxhcuXB47644gUz1uQYGUlQPSGFdwSq5UHF4eEjkd5P3LcpBzDzasmeX
bDJCZZhzeTEhSFaZ6tinKWocHLFiRC2pwMi/G7bBLO+l4neBdyt1+2PWQkR2GXda
7rodFqBpnVE1wRFui3tixpPQRFZaX4eJXzZ8D83551zKRitqQll/oBMgfbdWfRLd
vZLOAkphk+8c1SI70rvqBIPn0pPSiYh8oJdXTmGRlJCpMniWgUR5kBFyy1Drs5iJ
g+yqkhilLdNs8/GCkpcTD2AHX+pjnCsOD+Qd6mjJRiI8PQNn3rWONxU0hafePTNr
daOxHOr3rvKP0n9axtQl/ZsFLjgU/qL4wP0TKbSyyNYzxePia9XrxXHaR3PFS+oc
9leGTdEVNpYnPucKAx+faXOoplAjJ4XduuWuSXYBk/IgQNORbPg1ySdW08GSBMHW
C8pacocHrSSSc4ed6FZgqKosGFtKrlCI+1d/Q+/ExqMfmjphsWcPn0jNcWrEV3sP
BwyaLULF7AYp7Th1mh5tkQfcZDrnE/fnWoqVCgGdCt5oLZoOEJTIK6mrZBYfb5+i
aolDNa5iyMndv7L88kTIL/qfMOFO5SIHljafcCK077SzcOCm1verPXD1jhko2YxH
qepbbwiOG+YKb6rYdxqhBlWUJKQcEpW0MT1MeVefwFGCOPPLP5jiK9y9K38mgXOl
jMIThdb5kykXVZrEWc6NAu03goTQ+YqZNE9vFGqaWL6P4vDQYQ+OlqwwpmBqKAhk
8Lev8tB+ERaigvfZVGDBBgwhPgqRZsAlmgMybklwWqsdPbzzcMFjC1iiOZJpboEm
V4Ks8Jb98yn1niVP6AcJ6C/jLZVYweMyVU0lIuZLFoyIzMFlzs7XNTy9qqUvry8n
ewq69FWIB9sBhUL3rvjhyz3+zbhcbfiYtJjk0sP+F/MDcBnhzbBO090xBL5kjD1z
T/9fr2ohp2mf0BlPaIKMPEN+wmqr77zithGNZIAr1OIwweBezJ5cgcWcc7LQTOyF
91rZmLdGR/mlt+sPqiCIjZNTOu/PytTIHSKM8mghMIKaU+v5sbpesv79b3T0ZlA+
su0xYcaLEMchGqeCMfqUJ+Q6F/7FNotEkRqfXMp7fM+4Ds4vT/4rsDl3xzjRpxJ1
XLyCFsU/3thf4qsef9VTCaUCAIlJ5++aMh3uXkwH11mYGBwUEIR29DygwOHgJAi1
3m7KS5utXmWaVmR0vXuykDAm82GuGDbqNVgm4QzQU2phCJ9IDmku0wAgRfEaP7Yp
JLyAY04Zp7VOfQrAYc6WWD6/eSbCtV7KvMw4RUg4w7qSUZ7sDkDYf4naG4isGae3
Z2o55AfiliQdAY9rM+UIZVdaMhgmfASTW3cBcfpduzO//cPV1KpGvD534GhWInJZ
J54QFFyUdTpOcPdpR5bAQ6BXEfhW0KIFtQC/ZuNhaITqmGvDLfJuX+fvIINtUVAQ
JOYO3DKdzepjNEakUfJ6XnMLmRZb3HbbGPccAIBdwwI63+CPdKvKG68k0tXBq3z3
KkkbK7orkWqj4CzwBtXioHmJRh6t4NVZwuWhppbT5NsUIz12ZT2T08mtMnUAkrp1
zV8FRoy7HVS+JkZdlSBLTvi5R2wv4HvBSWkoC2kKapzGPq9Pl5G5dSkYcMDLIz9J
Cl9thpc81C1SOegundbv+YkhuwRnzc72kUzNf1a3Z7fWyn8EF5wmufE7xQpO7HQ2
KqlnoQ0bN/AMz99wWAQXRmkA3TFWCEb/05DBrw+1SEQUz1FenEOGOun+KeZ5SGl6
Cq7ulK14in5JO64CuGIKtDGuSLX0lhPzMbGndVI6z6cL9c7RqFBndDI5oTZoNjSR
L3weLB15U08nOhppoZ+Bi+yQEbf+cucD6rxSDiIYve5N6E+GnLfWhRVDzsH30qgp
5hQfVWv3q4cU4cD0zSosfOsIpbshYnnR8ecrjzHb668LKuyBT7LtmS22UDxNZHyq
fS0TbwI4RUixVZhaVLfcVe8lOW8fFVcqKYD/PerEvYlJx9h77XnVp5FhDBfC5dGW
g6Ggxy2iggfFMJo2ZwkvA9KOiY26MtDiReFiYZXgd02bz4j5fW/WWC9V50ul0jQR
auz3z9oZnMofHfCR9TlF1kiPnOugL6NOWGAVT6DzbOztFEVbNWSwH2I704jeteoa
IMcy2uRRVFSSIJThcIfRjYftky2Q7GVT+GpQetphuRPSJLorO0n/dmnnFxM7tyOY
sfLBpDRUof88CCt8pC4/POOzOnVUR3r1KA9ac+I3zQ7gJNauac9Ev/r2NJa5yOsW
74O6VMqQxqwq9xEbSKH638sRZL7kcvnqOaVPWe9xtHzxKVDhvUkkK7z/3i1CIOtS
OHHl1tpkSVCcBPE1WZ/IDId3zsZPpxD2JXPN+7hO9ctoeyTSDPE42RSqrSsStXb6
4NwVIQ+RK6Aqadgi/527LaOY6XsoN6ed1gwf2ZNCfZkqketDI+gHwSHBHY9NUw0h
DBqLPc9C0K5DeFf3PJlWfk2BkZkoBbuIy9kfTbb/lsqlUW2waw/DQGg9/q9VtIMD
Tvrm2Ber+4z+LXyxxhOzPcJaMvlCG/m6rfm8m/nVch+V6Xs/NUFHD5yajM0PKAld
SIYXNoOVdX2UzviAlly5iQpmlGQCk14tl04q5clHjwBGKRc6jbWb/nChYYXuADan
PVDCEIdeRtC05tdEHXDGYREOUKZiB0pftcrX5ccEj38ZBtSwQNFKCG+VwH0ZDfeE
ANfzi4WARQt5ZDPZ+rvhvWTdbBGiRomkNiLHeLkHkaMYt3bBwmmYVezXuhstaOHY
a3OWrGaym3sqPl5R8Y4faIx4qUHHMSb0QmY/Fz/4iLs3o2uMO2neMS5+TdF+X+nc
OV/iIJCggRtTBK+WuAPgOvzvcZUYry3f9j/UyuJ4wy4+gMxK4PcYyjs+rnJ/hgjk
xTLC6EN0NwdKbv0PXg6jZNbEOX1fcLBiKZhh87irkFX25K0DyS8Mh4CHM6FYchPs
UypvSWUyRxXTtqLVzQyl6nJ2MAKvXWjGR5WfvQQ7IOCChI48QCv4XOOPCpyyVL1n
10nL6Eqr4KWPO4gOk/G62+EpWMN+PeU1jllIGBFabhh2GACFnjfCeHBs+mvSyd8u
eyoAWvEwo2dElWuCCh4E8tI51ZNLFN8z0zyov/qMqxuTEdqqh0nKDV9hmGq6pyEm
fUay5FiSOp7nPZMzBkxXFz5MoCSRpsnvmKK6CCylMAP0f2Vz5hMLn9DUBhgjwmbD
EFap1xvcLegYdWesemvho3HAcgSV7EqyN5upDgk7ChQcTze9V7mNpSALHhWukW//
17cCIa93NRRnV1M2n0a+bTURmlm7PodCHKtOp8QvBk+sX14Roj1MfNjmyfZ8DZgg
1AIS+dw3xhVObqhoJUEwtMQIS5pwCLKJkSiUhGcW5UfwapSj7ItW4N4XXTGlS/Bu
w1C2TzizU+Kfk+6DOxRSiPtqqfAEZkaGMxx+ZHCdD/oUygvYXXIsBpYVKd1BvgUG
CrU86pNow8fx6HYOXyMRpSTPw+w+BvsB5ngKarUWbzDO9CSe8az+nBb/2PBaY+EW
f+I0ARr/GxmWTYBM2RfBemH5nH9jV2BvbU6rXO3poUmsMbrpyiaW3NXC7Ax51HnC
MpBt9bft7DnEK6RhjF3EKq0232sH7g8q0RqwKJ08oAesDIPQeR3PjGZ+lJDYvGyz
qS2T1gcmbpmugm3YOQraTQoPdA/A0TgvH1gFfCBR8FTexAyEMmiHu15DBsELm+lZ
nD55IfZWUs6U+FOKn1+mHC3VJlFf1sx4l5BOH6sex1jD5JkSOrl5vw1wYMMd+bEM
m3ITrqHYY3ARt4MP8AUcm2OlzmT1YKXM3qU0Xmp1m3S0tGVazWgzWpQk4kXRqmfq
jtHIZ8J3J3XXeU3iNzsmnB01+FWbyw5zXOMfNgL+Z5C6VFPn0vtjNZENdctNfVtp
m7dbAnrkEX0Q+0Xo9orCMxetlMCEJijdbtZbJC3thx77iuRvRmJ9wBOUemqb0P9A
ZvVVw72dZPRtPNTIWL6ALMShqCG0UVqQZR/QaYD3CF0rTalO1lc5Z9N0NQ75zVeP
ZsInrfFztNXEyKKYxv15spbeXqycnS+GZ+9NYIzg7ngxpI8B1jMMQLsoHMXKVNoG
1VfUn8YnCtqKNpCedu/grqwmHqAaiI52MO33yOFaRojmzKhyMzmK4Yl/pGCo9x+Y
RxeYLry3vgUjHh4fD4H9ucSd/IvusF548CKCSphJ6CaZVeQVQMHlU7PlcpCvBUV7
5x+6SPnacHD1MBGMuIOqxgdsIt8/78Ao1Oyvs+PS4ctlgXjKXQxqEOqZuUZhcP56
XSKg7C4IzuTX2la+dXbFFt/IUVlxdzU8mW2u0cDVQAj3dfltWPAUNvML/Yf3PStD
LxhG4tUZk4FuaA1xodL+NqO+edh6hdRyr4NvwRs2PkywD9lK9NRS9n7yotG19VWc
/S6WUo22MT5lxbtMIQ/LxtJvBEwvVB6pLe2kYqjWTkMtSGkOAKy1Yn14Ht1oGVBs
xJqbgU3+Y3/eMkVxIjLm3qF1bGe7XNMKjLMo6xuacYLuTkKBrzJ8vLdMWWHTsSna
tfO5D/ZySw8Z1xXKa5m+e5QW0jKBvOe+WtrjjdNmMxZwVGJ6Wf2eZFolcmBiUf9o
h6BgdyJrgmoxMmspLAZmd7qD0GUGg9YuXfLt/D3QE5rRLICO+EK9ClsDiNrK8UXx
JJGP5XQWnv0AeibG3YtIIqVftvCcrc5tyEss9WWguBwp0eWOVyZj7tAdmcTaq7AI
cq4BJmaWn88CObKrQvycHvbRsMxFUNNapU7HC/I7mZfZoiIC0BGVo6fxj1qz6HQo
2kbm9zvZeyxEJX3sKw1/osZfmTs+1Yeht/jEQf6grLuVp2N1QNKmPcjXfq0G+YQs
FvpeLlLivG3+zQ5WiURJ+1VoEjcPMP/43enuhCStuLdDhANtPLcd/OZx3kw4P7Qt
lhv0CoU4WzV7vt/z4ZfLA7HzqZsQa8P/P70nCOBpuT340LL+AgOyI74YF9PYBO8j
GWqhJjhcIf1y3t0u+j1f7wYl6e/jsnk2zxZ4KxuNbVqPfUAvbSWFzKmoBK10Z5LC
kzzObdOjuQC+YAudL+dZiMFzYYNCHzoazdoXgAjMb76Qvd1eApfHPwkLWxxCgCF2
C94FPAK6mZ5QH1lps+g48zzCZePneQemZfmk+JCit1k2efDs1BFSPTeEeFWx1eBA
D8AEg/+GVWVdqLomWEVjvpIn/U5WWzIc7PZJQpPvWaGxixRUdH9wEk3n8c5fAULA
a6rbd6tMiE8gxTM81ji8hOGyM95GIqRDKL1SsxWkcyakasIg2OeQklDhpmW3ujGM
/IaZbclfVExbp+F1aAmC4kPXfFn2Wbj03EsKrnU6C6iFzDHi2mIe9FEtW7anZe4a
laoz8A9KL782sb4qUDsx1Dndw+q0amJk8IBlRH+d/EMdyaE4BUw6WXtjQaB9Wd23
PzIX5ux3ElH2k7byIfa52Nv41nkQgFut2+weQz5AWYOvFYqLl2Na5atr+SDnzH9u
sLZAnXu4xpFEeOvERkRWIcFwJS386L3OB2yauaqKfqZ9DjS1M0qgjdRQJSZwASft
PMceGThx6RnhXopzWOKJTF1ycelnV51yg6OX8YQismqhvv/qmC8iXb02rKgusYgU
6kiI/+c/mdV9sQSMlKxMSyXvRn3IFpDoWSToKlQUdtunpK61yFalcTZbBlMPVqON
MGMBvQTotLRZ/4QN+srX9kdKpHuNoeQMj6hKhIAFHSXFjz8m03bK8GgMCi8hjfRv
/t5PDqrN0yhT9ZJKdyNUybSCTIL2Fx2oshHxQzb9IhjLkGiGoguFR2mekkQ2Fn+I
R/M7RUxk/rd0tpEUJppn7a8yfJ5pZgJwZ10vZjze6tp8IP1idjGcf3tVGGKKeiZk
CA3Eq8tAG/pSHz5ZX91ClGvrt9YenwBPIR9HIcnwd9DIpmiCOBiX6Ete07x5Qqk5
lWW/n2ziM5vW47QjJegu/IDvx+oQS5tfSXbvCRHkbu4wUw4JK5ujwxcRzWeXwkFY
XAguqhX0xCQAUkj7v2aEErU6aPZLbrZCyGWyXJ0H/kNUQZBZBYVr1uDjpQEwtsPy
pgBqhZD6CawrgGQiRutaqwG9QdpA8oycvZO/tYU6tuWe+KHOmshWQOd/ob9lYAR5
WoqhToD5HkFwF3bNNpqq+/Tg/0JyMw7m0448HW4iY1g0m8iIj9D7ciO5dsoX6wH1
JxcdU4j+/1gGQb68tHni5qFhk7FmzJ1Bu1Dwu/rSgVv6v2rI4AuY9lhUgC9wNJ1h
VpBni0N7Dml4x6+TxnyZCnlSFc6Dg/9BJ0lp4ZRn3TUsoFCsdC0dpX8pAmpIjitb
mj8PzOIf4HX9zzmEmK1P0TgGaofJvh5aUDA2NWaXRI6khfzVPqbvCm/Zi64OszjA
nAapuuzVEeoCh1pddIa2UOBLuxdxCdZfjWxq0aqXGOsZt+W7FUdGkFyLfOk84M6O
klv6cN2LTQrWCF9jIA3dQqXimKtteMBVkCYf2MHFKjaHL8qGWoBAbbKis45WbOA/
6n1kq2zwTXVbhrIOGlDecv5Ru2ttTCJQxIMFNzrlIpItVGT6oOGAuGicDUElegd8
zOEeXh57FNTQWDynm9K/QZKt2UhRX6CTaOw58dnDYp7IXqUElvtuFXPFUIjQBJ3C
08jlwi5alXrduxINRrAwQyd08tWt9n/zb6NFytzsklpNWpuVpDhC/WssBdJJlus5
rqV7Ht5KLxmJWavhMSDnzMQPUfH5Kx7C3nbPjxsu9B9LG9lpZGI+ZP9siNbh40FW
fViBslPnuAQNj0sq3muklmx6NJ8pl95T8VYcLMX5KBNnCqKAsmnn/+K2MCcmqF9g
ZG/PT9hKCMiITSNtSGeFApqDIXsBM35I1smfle2/8+HXAhPEywXplsYclwfh80zJ
+NtsbhiRTo7aceSejduVG82+qFfMkVny4SePUyA6439Tk2WgGW+46hpUjtJrzC+/
+EasKbZ1xoZltIBgzqghWN5EclRRPs0rAbiIiJ9YjaA3xS+Gpf2dYeN4XvGp7rwl
YV6n2bGiLjki6U9UVP2D3wT6SC7GiWXE6aCyyTTDPKexTFvJVuPM4l7uyeJfwgL4
QuppXBiEgrHrTQc6yylOcfM6ZKd6jrJV1fHanobizVckCmB2Hmxvtcmp9IBvNqQ5
xeeKu96vdFCJ7zg9NxgGnTIKNDYhSR8+hFS1NLHTf8xiqaigOLF2l+R06teFMjx9
DyzxTFTlLbcR9OdYbivNtIPUGkq+5k/Nae/Pqco6++/dGNAqyNN9YWr4dlsYpXmd
oyPffRwtFk/zXdYeuUvxsig1w43dXQ09GYqBTRWASA/wgLyuSBZtt+j4yZm1zJy6
ni4GYDJq9CMG3R84x4Nuso+cBgN+bS6Ggqe2QDMgIMu0Y5xFumyqMxM06UcabW9m
U54Up8Q/KNUt9z7ozYHcwJi7DvoTG8L7lKoXtDP1n1AhELBkGZJHrkGY6rHVM8oV
3FwDzUx7huEPH9qMYdCP6VWCbTy7wtqRsDag2o+eYmSWXVVLv7ls58g2PYA+0zmb
rl9HXz/gPkwsBp+ccOs2fgSD8ezKEtbNZhZQ2PDxzvBweNYFM5v/wDK1QW8bn+iY
eGArWfGdntTNJbdYWRKWijjvkKPjXcVV2sRxVlibKZbTz25X2nPd2ihSgoLoSPby
K7w3x5SqXP3ASFQDH/cgLExZgcCnnVEpx2rwPZlsGX+yfDkBYLYBqpZ/HHg5s8ZW
dW2zP7DdzQTxVYPNh0KpVC91F/T39NjgRzuSyr7uIaSiBDyHxmq8fSjpUNQ4UrVF
5GLy8IifU/UYccuLE/PuVDvc5Tt0uU3woiwKyNqrTUPj3BDaOoPGfPyWzGtEsvU+
Ni9bJ30OXa36l+nazLe9GzYTJkDU4A4olI28g2CteNl+AXHy3+Wdke7DzS8SePra
by2Obep/+opyN1SsBl0h6F38YIkeVnlwNGNh0AzWMaydlag3PIDPXB/4ertQcCKo
gc7zVjzkLIjEdFj4ScuxKBiAPqeLtG8G3tNMdBpZ5fCW2kwbfYFplpX9146PrZL0
Ihem/zWBhEywtWd98U6SKD8ct0bB4bYeGUyLic+MyoH71k9yYzmGUl+mzgjSBCbk
R20PlVMLQaUiiJjCC4Iz0BQ1EpWNC7u0q9XD3ug8Lone4FGVRWfJULsid/XO5rpN
7T2oPLeiqV5WZkjGCzw+lZ57n/MMz8e7YsUdjMlJaJf9Vbxv7VV05zAkTfWruxNE
0NdmzM0MSO6RjMISh75vOLwetZhWc196Og3+jRpiM9AR0qBoYZ5pYOYldwpYze4D
SpppL6sVv1E0RVPRnzYa9dwDt+zS9XxUhVm8HSVisrQRDyC8RdRvQDzYbcBOo9/a
YSaSHii7tMH/HoUzlWTE7Mqf4JWhSSYpEanFQnfE9c3uGAqshPDB8Cx4GevfX6pW
KdkZ7TiSRGfRzlwvUi1sIKR3SMsofbfRqAlAGRL8kOXwnKbhBzYZPgLoYd/ezyHu
zdqKU7umBmQydpqCOO09hhMtk6lVo1mNo4TyNe3WsJPjEH6z51iTJFR1Qd4eLpqH
Gpx2Ivtif2NYNwXw+U6nZy+Le6xFM4/9CD7NBJGtrqE2NR0iyZ4XP7eLx/0gvY5y
fvg2xYZfs63DAvIN7EQwT/mFrFQ5vcFRuDkOG7fI99AKUIaGhrQUi7R2I7a4+syS
tNqwIQEG2nfrm4HR8WVGnO/1xibKZI+9+tIQpo2c5B9P3ouItUfeT3uo2jFwTfCd
8RuMblsZqfgmVPyQxnl3bqsfpROE7avCKhGFRmJxNuagKR7JZTBQMU1zXOHnATD0
KXTy1piaufB8fWTya2N6JdhA73Ikg+OBLCVGZ5k8MacknYo9fgHGleyAIWfOKdMI
3Y0wM7+4gFZkN07/7r2oRctuZ1PcjUAMJzaU2auDTlOdm9n4speKwBDVV/QFdDeE
9C6a+kBfU+rUczQuocz8qHFrQE2cOYoFBccB0DU5763kJ6bgf7CCAS5DhAt4lgY3
E9brffYtyV6sESHYoqJK8QKt/JA4AiqNP+mE+7IiGulw32egRYhwm5Xs1qVVkd1c
YMtrrySEbNHdqwHKQ6w6J6vm7Y1d5qzj/GuaCkBP+VJPPuDwOz0T0KCeoR2fcz9n
+HQmjMJe+VIIWn0CeTktrrhpocZqeBwrnkKqhfEB+HfLa3UV2b0jC4z04FjevoB+
TJ6JQt2u4rhZH8u6ZYdZdQy2qpy/cy5l5Bd1ZH9FL29FTEFt7HBt16a3OYk8aMlY
ucHDVCi/vtE+BHUCXq4sfF4xixAMsOl9UmqePiwEka1sijqR7gt8KuFgcJpaUJSW
0FeBxwMYtlV87iExQZshCYgNtbs2wrDBZyKqlSKdq2qOtugW//CyaIHTogKGnTf9
ZWcimTPMrMnZzmlBErT42fM4x9noYOy1t2bEtpqcpq8/14AG/t4ffPUl4bOQ3uZS
ayQtsDgNqhwFb1Wo7ZXq4OfVIXzrIEBE3pB5jzmdNZ//LmjjoIrTRMZfSXPuH6i4
`protect END_PROTECTED
