`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xpNlpxVfdCRcy81QB3YeCz3M6jdY6TivTE0DtMa9rWUr5/pmt1BbDiVf7LpqOKUd
WNjZwyOZC0gNwrHYCe+OmeBue/EmopklbJ3XpgxE4JePZKcZPR+DzWSCytJpllaF
T6MmcEveO0QAMBoQhOXzYrkVgQD9TTYsGMio9yRtlBlyWHkehBgloIkuxVQhZ57z
0khDyNabCjo+UfcOfXkt1lvvCHGNkIYO/LzMxyuo89sKE1zxuugcvtqDDF2nFXB2
SklgSf9Sat+ZmItTBYpfApQGyE4bXNF4UgTRYqK1bsHODIkSWgOhIAIt7lmlF8z8
NGwh7IGFEjV92LT78mJCVqshGFagsaAq4i8wpgpywnFLs/rlz2ylKLgHhWep+JRu
Purg89+Cmq+Pj+ZGb26NiUp6iyQyxtdwZ3kCjku2vHJvhdb/NbmsJohWpoZeyWnc
SBZQz4qLGVPK9Z/kW4XM/x4VVT4T5iu5oGTx9QJtX+4=
`protect END_PROTECTED
