`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
12u3dsCbV22D/Kte5KOD7eLUbKapGGUIrX6jcYTjAu36oLalDNHCyhNA63Qr9jEd
I/w9Py2I/wrTcZDBFyIluPZmZwrLvOAJbaae6/CabqKPXB8MfW3gKs47tmWKrre4
GnSvIIQgVD1ZwGwfng/OHmQQt2dztpnEgaZdvVkChaiQEm7h28qlX4tLRDAImLDa
YnVTkjoV16iXHm63PjKeGpwwycVD+dFXvIA3YjeRRl7PfO22Jm0QlHymz/hRjo6L
D6VqifLt1PWgenLIT6D8gRf4S9vjIIS4+vO0bmqCAWt7Qkm1E6/3peXwU2KGa8j8
qEXBSjr0iBA8S1kwqbrjLZO3kQGdmA2BJNOySwIkHlJM+pbK5t0PAE+heYbF8wQp
tK4mBSQafvP69yI7Mrw8xBy6O4mmz045+CwicgGcwBM=
`protect END_PROTECTED
