`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pRQklv+hUh27EwkkN3BKLNkytCIwM+uGrRIQP2q8Q0qCLIhzFIZFMW+jyckpJnus
I6aENDYSeCtJD1Kun4CvawzPZAEOzG6MNQirzCcdkTTC+8A7Xvaq/qpGVh45V5Kl
d2v3PW4uxOuimAJrjk51EpYMXM/7Pv4mlSQdwmAtsKqMNtyXTGtsWopyGp1KMOMD
zkSU0/gy3CI8XEydwVEH+wffjx/ljiQYS5XSafXr7UwsNaGGBA2SagfNMSZShbnf
Vc5TJ/HCQUgRqell1f4mJIviA7HAN3UvnIUFXakxFdtzJasVub0SgKDgSYMKNcaQ
AQ929TlQFS6rQ5cehCrdM6WRl0V/p4HvIwKdPJaP7JxZaeg9zcSktdIoN4gdkI3E
W29eBeJd/Hsq+yzfC0MU/O6N2Y+95hLB7ivwbuZ+YrR5Q4D5f+b5Mmw0UuXihwKa
WXDqDm4ru96ufForDAJHmTB0lb3UWpkRVVHAMAyo+iLXkOrZS2bWNpYI4WSDXl+U
18cI096qlzwFVSVDJUhPg9lk/nKaE7gTNAxaTW3Zu0VOju3gYCV+8JlERU4Nc2VU
PYMxnlX9LT3iQ+C4HYYil7JUQ0F3SO6JZP9uoeqnFRrFqCH5mD3R6LfRpQAgOlNR
sGUmAygZVCr5otyuBsNaRA==
`protect END_PROTECTED
