`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wf/N/2MzfimoLDhSynODq0tqZxUar/2Yo+ORJhf9ofB+lQuFfHsf2tMn9CBo9vqE
P0EYdBQyYFRG7IfOWuQMPExNJ+EkXcKagAX7+NTgo9mc24fCW6MuA6RHZXFKpx59
J4CNJ2kGzsiR2U6v4uosqqwbjEqi1D0eez3g4hS1en6elRuzn9va7jtXtOw+oqud
kMovm6wVhi79s0mD5lkJJcYVAXTy/HHoboWGdIyeyF0JaM4p0KnKajn4a3Aw8NxR
`protect END_PROTECTED
