`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qFBL71s1FcaOAPyGVwOFsOjGbcWqOSLyItIczY2LaLLdRZopOU4qyynHjES8Unf8
GD9gf8zcN7uweJEhclSDsD2y92Vx7AzKJrrw3dVQd4IlB2Cw7seQ1xM0Yyn9aa77
ZSQgHaPcQezxaIuo2jKSgnvSjpgJFgSHB5SPRLPE3GA9SlZOiuBMGfggjpEOsdAt
th/PXQZYNHce0cHJdsMGCG/FUUXyezQdoi6mXhECRkCOwVf845nNv7o+VpEcadiu
G7VhS4aiqxYaRSI+j98oq8kjwZ04cxkiZkRzoHMDdks/cCbErJdD6gfLrqCdsM4w
608nfrQjFVGhiKqhEFr33NM7wanE7uWGrg9vF6udEJe31fc5B04oJzQXun17l38x
CO/Idv7dm0DBcbNUH+M0KCpZCzy5hD9Lm/VpMVUP0C+QCZ4iDFNR1sjhgXEcEw9l
vHpW4W7I5J+XmDoQajio9ZL1AH6GdhxWYVTtPFf0/ThgbsPOVJNh6899TtCqkT53
FPe7XPIRTQ1Vi69AFCSP2/Ci4Brwv4iHiYsK3TP688Xmf0pan2bsiZISq2Z8u1Bj
S7I3ovnsJZ2LL4pj02IzMuNUTfpdJlL6bYjKeSrSyogsLGOoJL8T5LdpI7iO+ZmT
v91Fq8qzmvQZ7gCR64g7z9je4tipjN7Hi6VYphR8Iz+3tbvaLGZUTfXF4Lwny9Nj
DxvqX5CxIyd1pvd7svhR/NGV1T/4i9TCYmNrcVExbdjE0p1cIFguk1NZEVS7CFtp
8djbEkmohqGCCxWZhS6XkgJ21HNiH46whDFd0+P1oI6qM29r0RFmp6YHg9AHneYN
6hStt584R9sdZaPMrHaveG/H7lHeTDiIDjhxpl/bEKpASQBYffTpwWuPdMvWNRVN
9AkMdSlvGkBxEYKR0NynDqqS+CEz0rQicXRtkA37e7CBzBVg2lwDUxjQnNlh714s
TXfHeVrOwCxFNXIz03MY713Hb/KjMSDIPoVsuugGrXpC2G9ztRSimzX20aPHeAaY
G02WJx/+xKQu9SsQ57RYMnv7Tf628526DiHDDs5jeilVfwUFQLfel/K7DhVqhpRA
QgIxvcR9aSLwWQRcIU7acpGmeSVE91A5lO47HFQgFJiracTSPp2EqvHsWNq/zwGJ
E7CmwmMz7CXhEQauAnZ45nRBB1lUNLbO5EdxYDXQeFSLoDODUop6494sWDeYbe+m
v8j31jpHZy0x6O0Oabxdrm7DXmC9fBKcu0lMZqUqoiRZwwLMqYP8iUM01ZgKAVYu
N3e+yAlR8cLg8aRJ12fbPjGCgIsxS3sA+7vZfFHaF0s8NBswB64rkXatxmCDIBVj
mbeOzSuPQvFnHlFx/msvA+LKVORYbRDYlM0SNTFGGwnhD21R0UL3+sRjB9paZcag
RMEaQuoUy/ym0w4HlVVqQxcsD7e8QZlD2cg9PNIvQsLGX1WRn0RpvQM1O8x747q8
+IPttsWf6sN8escZeQaxB6w+/Q/8GlkoynXc1okYzbWOT0xRxoQnV0e8uee0BqNi
yd+9UGqmYQKv8/q+yO9GKnSnzdkyw4uMU4MS64BLEiE=
`protect END_PROTECTED
