`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zkGHcIutvJ0SiGeAn9mMZ+iPG0cHTlhtxV75biK1OTGoLcH+vM4NPCAzwXNlxK9K
2CtVuncGTAS1rZE+P9mZnW/MLa28c94RPQN8bYDKdXucSBuWJ3KGjCLkUq8BUwp2
DWwXUVJGLnA3pYWjvrWusuXpoUoKkbjJIGtS+v+UIJWgciyT6G66rdgQSQ8OSwvk
M9hVMCNm6WG8f8jiUjthwQ==
`protect END_PROTECTED
