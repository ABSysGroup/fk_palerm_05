`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QMKlJ5DvvgqmLIODsar7msBYlgDWhXSGfGi4RIB+qOwNVpGgog29koitT3xib1eH
JCdE7lbhj07oH83KmzK4OCNT86tlKhB5WG4n5jVbInUOk5GtCz+DA9vfMhM0cOR4
S5MYBM50oovO0zn21Rb7I6bJNP6+mf09jeoJGP/jlGvfX//U9rnB1+WxVezHTnAG
hRNy7md9//qhNJRqbtGFYnzpMaoASbPk04M5DpFa1MtldnnO+5Ix1GPgASKJexTC
kLDy/XJs2A8AGq2y3q+G1G4Ndu9FE74QZgV5WGYklggCD1WK3HCy+B/H3NV8hG8l
0pDZADJ4CjLygU5OdL1KrA==
`protect END_PROTECTED
