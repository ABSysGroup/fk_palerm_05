`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b+z/h2cbQk6nFVBXz6Ua5gxoIdKZQbfjv8VMk9qiW1NXKKbDfK3HxbdnVvK0WM3X
hRbx/qItA+ec6DvP8/cKKJbmtxyV+uXDyhcaEzWGNJA7hkJ7VwAK2SJkfRwM3NnT
bJ/FtxDMFfie3GaHpUBkW0stqUd31r+nbA2JUIpZCReDW7e34e/bGuTQ59IQKJBv
mzXlSYu+lM7mXoBmKFs825nlXpwnM4j9itctNslIQig=
`protect END_PROTECTED
