`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NEsruB6dLa2IgNFknhHGZtHBkhGUM2gPJKehBEyZPjHPScuJcM8CPL0yjvgbDt1o
dVxOIDHTu0ZkBeb3wBsOG+fdgMWp2Tr0p83YjQBZUoQOtXb6J354H+WLCpNDj1HI
/FLDdSrehw8ZvaWuZD0Xza1uAyvzbxRBJuOqDGyHHvjaLwb46zD0o0DgQjaBm7v3
/jQJUNLU5wlVjHVGxbj0m2+gAOs2y0hZitKx9gbg9iKIUwsLvafWG5i9Q4gUMWb8
+SzG+0JVFAVFmpheri/qop5H+Lmoowtxvw9OimmWEwHPLIzZW2r8uTt/xJRQpwlv
6f2VEqzDoA2MVJyjJpgLLw==
`protect END_PROTECTED
