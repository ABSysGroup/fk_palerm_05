`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rl8HOIMd/oe6IxK7mDtEGvdGTTYptNyP6S/LvLalMQtqElUFamTERvfDytEzBPrp
r5IIxU7TDI3qOl6IVRloDOahCaaUEWFkf0GY/d+7hGlRRrmO2xs8TWbiu7uZFGDk
1rElu/BnqIEbuTlJs8lXKk6msfjMrpmsrM1PmwmOIa9fCqUhRHLVBZ3eutnz6mXe
aT6so3sZ9tHEWEphdBuI+bP7MPVXmwZVgyFpgU8tmjsrtX/tlZTpibXKUaZkqG/O
sTS4suphFTc1JrSFAKhbm59Z41UvXxskulgdJkR4RA87UZblCmmpKa6fM58nhWem
`protect END_PROTECTED
