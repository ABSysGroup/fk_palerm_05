`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gMaT7sH/PCMSL5+jyj/pENc9ndbriS0nXW0rGQd6kxm7d0lU19eh5hFAEiywXaMV
o2YtCBVVxjEZiGZ0+1F50Y7fsxhIAqImmpWd6hC/CXLFTsaMaQmIuHv+//Cqqn45
lhK98K25LhNlmDOWUJBFJqytvM7xD517lqqeVD88teA7SF4sb54OtN3mdo8oeiiG
Cnc/L8blwdSLTBqPh4odEjHIXikjdeA7gYDr8IqTrcKDd/PGWtTdFTiI/ZJbBZrP
y4l1/R812SIDkTaSv/0e32PTqvoLES5uF/3Tv1E6c6WHANubLScBOo9p7u5Ow2+z
0kq+3td1Ht0c4oNHAzwIq17twxiO6fYYG/JAwuCbGnC+4/IyY3I2tUh0NpjEA5+d
GN4dsFL10g8K2fKYL99EDwnlehAbyAXtNKDFmWpIqojvYAtGkIg4eFnLsoDjhvp7
TgTuUHjCpOc+Yp/ofl1R6iMfDNoTLXW1sqre2VUZYyOHXMneEJW5PwxBvjVUZ8Lm
8Wb+kuo26MvbnSEWO/eEBm/MdH4MpxGZ3AHHS7m9FuKcuS1Pt9QWVOaj1jBkVYIs
5yhvHbKYVQUYVnHdovovsgs2iz9xJzmDRuFGL7TUQIRux1FVn5Pjbbf/D7xPlJwU
4Vp89cJsfpkCaBfrjoGdiipCfpkFYzffFdyQa7k4ZetVjWBXw+UAny1mP2vAg4Xf
ovq9CYZAf+emT605cSxhQPc8p8IzlSkNYpxYDbW5n/u+8+psIr6eKHNrdYHW26q6
HZkHphpk/0YbPEby3lQXOyzuk3QHrkI/regbscGpOMRXVfTCJtBc/+668Gc6lnQq
g65n4Y6xRGSLBCwfD3aXOigePIxGOgn/FHBfSgBvHioAA03zeVtbX1HDS/U5H2rM
DIuE8HKt3dHnr0vA0pVC4uBa02UoCtZvDzvQ39tve+6zCokU/4AA/KG4RSr65Aew
`protect END_PROTECTED
