`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jZ7rbiHboOG1DdfeecCxPXX9xP+HdEaM4C5pAif1XhEFlHHDvPkt2rjf6sL7hvI5
aJoblO0Z0ADe/9Gc9f7Xarz6qhyxXVxWTHUezhR02vOTPj/wKjWCJ9EX5Ogi5g0n
9uo6RuzHACavlLWZuj5LXl32nleUNIZC48Vb+NDFz2oUJUxefTMzXDnMXbE9rteM
HwljqRFpCVw/URKeYcT4Ih3x2XegW+h4/21PzKFNcBw07ST1Y8rnceWcsdnm6kVw
kaACZENGCxHhfEfWWSBSFTtwt/zKvBnTYLpjkPL9JYm30ymqBgTouiKSdJ8JHgwa
jUQ/o7iURu+f1SaecxFcDdb91jgSa0FlgD4/JD2KBap3ZrJpFt4Ue0m/bdG8uMhl
dQVLGZnt/41K+6rRbaHE3y+SSEHJArzXpFi8YXhK9O9WIFPA3ViIy8+Ny4k9VczB
HwkHuof+hoAZ58E1g2+ezQFxiBDSSDDozFkY28sj8dPiXDUUE3mF5II9p9a+qyPU
fX0r9DU9z5oson3jliyvPR4qE+m8d32TJDoRt+6W1lnxvLtS5xHHWeDo1a1zAR5P
`protect END_PROTECTED
