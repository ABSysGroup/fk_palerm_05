`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ONg3fojG9bzcMT6O0MGovXHNa0i6uoo7088CQdClgrQVs6Yqr4sfhdCmWcCK9/wT
DH2qscNupy/kqYEK4atE918pG39Tic4XO75g7vgwnogg2nt6I6ABR0jwqB3BFZ34
YHtiNIQQQAYvfln1+yAKwfZAREcVMeJn/zJJgLuoOI4pfpNQxv+l+RU4C2FovYmN
395KecLUGgdfJJNl8sBxWBA6VlmWD3mxnopwEZEG0SQy4LaEINl+lk3pVWvFZ6dU
+LkJPszufWv0DyTfawqBaoACFpSTIt0rDxwevWeaCJA=
`protect END_PROTECTED
