`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X2cau1AZBHjuEhIqBVLsIPavWtO7osFpHcmxUbX2Y7L9ncvnZkKrOq9LLcSz/BO9
cx2o+rEqF2kWnkdIi3vl/xJWJxNUOTX3KQ72//jCly6VzuA1sY0FCaYJpIeALD0R
ZqLB13++HkYcxhpEQN92YUHpVBFI/Iq+dxrMs4ykWG3BDVG7joU6E4fn8z8s6TUZ
V1aRTBSBZNoFI4QonPT97vYDzMlrKCGPcVF9lNYE/h0C8dWf88NItTLWAC6VS8Ro
PPbVxPwP6ys64Yf0/mlsPzG9Xeia4B1/SnkyrmMrsSQckP8xvf8svx3fM5TaLOUz
ZMn1nxXE9iPOapxVsY9YNDVOciyrfQ8T5JY358HhyKaF9vjRNSr4R0w6uG5PYiwc
L2fZyQdwlAM0CqXZBAxTEx9Kj8k39rI0iQ2FjycjSIw4NPEwCT6jCtQEHod+tzeC
Vo4ffRN02AWeUgTFBBfvmJSEzvwSeZxkSmG4Ka7yvSVdxI6vHJ+mSgkGUlKOOxU0
1/kHs28P7190mJz3G0rIXfFgZOk2mQGhyjs2V1xvdLLjdX0V+AvxBloNAGa1LZeb
eS1KJMrDdJenG+RgXRmEUzneDeSIcu2phsp3TSNd1I0Je2Bm36ooyCkVB8BKzTQA
Xr+2lTSnVSLNJYGJuHT54jVXqFbyKNviwUAuC510/yD2Q89kw7mZfvu0t89jiqo4
0pOvLLnaElzHA0LUwSwrf0maFTO8uA8xn5tRTZMDDm4L82vsEOSGQU6qtF5eMenL
R9fkx0N9l5+9sbe+inEmhN7aa5xNygmhR1ML3raRZRauGIjcAweQj5PKzE7qFFQS
e3pkzowtbxpbWdt+ikAiJOU/o+BnBd9jUNkU1mnbAQywrll3DIIwIQXZxnS8j2jF
4hKWaZc6t3039/oek2UNiVEMdl2UxO8glOMaYrZQUSplAWZSBnjj7N6zRSvi5DOQ
G58G+SoKL1RcpPlnkDLwvYakVZ79hH+SMVVkd03aG73DJdFgqS4okOUYzaw5zpFr
HKYFJDZCk+FsAztRdp/LkW+J/OvLXnAga/nJ8Jw6P+/YJbT5cLqzP50Ggaf9TAtL
b13UA0k+aLc5tuich5gfEbzSeTqWbHlVoo+6D/oolqkMFW2Jredl42tz+kc8wkMa
kxg19AF/Bj+Gmt98ONpkWZJxS0NV+BE9BwpLqt7DDHuerStfG6OP9sCWCX1rV6Lq
B8ozyCuaoVkVj4rZiJC2CfNOJi27B/rZRZmkZi7gktaefWuup1uvaBgHaMXMjC3x
/vSSir1rP2rRV+ei4csQcclj5fuivqGqtv34+ZZJI/qXtpGShgBSfOTYfKEhBTvv
v1v3tjPGcgRIAg44ShvKilQXwC0jt8DBuYI+DvRpTRGB/EQXeg5gFbbFNYkIxO6T
QoBOEDuW14GBmHtGa11EIg==
`protect END_PROTECTED
