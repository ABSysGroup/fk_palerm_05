`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HLQn00z+vyKs5e9m5/Udk0ao6keAftHYfllWBicUWA/YAiWR4q6wiarZtLfILYYn
5zwRdZvr/roQn+xDU6RT8SHWpduWZjGyc+TycaGvzJ9jyVw7zdVSSN/SVRp2J6Rt
HIXfR4bsIeA7wP5PUb9w1j8tDg4l7m5icaGztkpElFMqPok9Njhbg50eic+8IvA9
mfhg0fBx0lYe004YZoT0CwrL0xtGUO0Udq9gZxNx+469ab3Hzeinb3sOKp2DEBx1
pinzJwFbeTYs5UobNtpmpXmqhWj4e/k/orjMlk1jDdCFK27MJy9lzleKBTrd0zWq
5dnhf+HpzUPAr3fFkO+fqLeGB1QbLEaoztL1gyU/6uhf6774SEmU/73sA0RjDW1Z
13JUG+n4+Ooqt+PSA0+UT/Pj2Hvm5oClWkstmMgZ3g4WEuWieZh1naVDiJx7d36h
MjrfEZI0bkpOu3YqvHyLUyowKc2IcdDKkV/dzptIlnkQ1NLSdOHNLyEzM+C3MW1A
BVDQ1PfSojWZAo1psnpt5/bYTt52qRy1L4ANjYMgaLL/NMWwCTCTcIDOcUBmGpcd
nutFeSD0tANSPFvZBTixVyB/m8kbjuTjhZAlNi1GHAK9DeJs7gPaaveVoc9yvQ4C
6z+08ERVAAWsPtD/bXkGWV1c7YmJMXvMpkcDPnIpIMvS2TtcM88s0QWYl7Dx748F
eQpu7MeoNi9TCChs7XyX6kFyOZlxK2LJM9yrVOqf5M9ccts49oiGWHWV3CC61NqV
UqS6yDxgjYhfZimIiA107UiOU1GfW71PsoBXPeZcMLyu305iWHKxrydB8NHoXi6H
6EzxKxPh/D/KOV3DLMc0/tNNxWVq6UXYONY6cIQ0HaW1ZTjP29O1f4i1V2GGFRhU
L3ykayyA9NC8dbzEaBbMgz9Aq8L19rNFMaCzbCA3xNHiCtrzHSnaLm8ZPIk7qTgk
ZBX51me2GuicQqobMYuM6dvoIVahe8/LDijDzLgVJy7y57rTvN+EoeSAkJrlZx1C
qVtgqhrXsaF2D5k3dNMBzO21KWlQn8YCnnFpXTptguuV032rWI4wqQ6dcZzl5Blv
QulvosTzrHDwel5MasqNC76ZnWWiBbJCa92sTMKUtN6yslQ9GYvxuv4kgt5kLSoH
ay6I+kurtXjTfw57we1q+pvr0W9mQTz5gH8U+VVjrBJ6L956UuCrAUrlEb3h+Nb2
O0SOU42M/2g2c5QNrzBZO+cs/GfH1l73ktMkUVCTPbTbeknhVRwU672A8rgeMOWW
6otluIpN3/qWHrKo/dzbtX3JFptFTEtvXKacNOStUPhfvqwbp8e8+82G2DglWorr
hm8LDr2yPyXJAM4dfmCJeNvgNJpKtg2p24heR6LFRyksAm+at7Fv4oskUEwY5quz
`protect END_PROTECTED
