`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dfs7JCuPZKWWBTcBjnhft76dxOyIs7Y/59DjPk0VvXNrWcwrQNjKVZEsHbj/bZXC
hM9HOlJBgmyQGnYAJCNiebAwHBm5m8ork2ZLZfpd/MLh34xcz1JMoirNnVmy4xfs
vnvWYQrObkYfPWQI6LyzJ97Qw1EtldzjHGgMd/qGnnspC93pe1d0QZY4yWxqNiwF
2OEw/8O0TQ5QJSiHIea5nA9AqJtu/gOajlRmuZjJlC3m31bXe1aiEMDyPciNIPg1
f7043vYF1/vbtaJOieVXIlLo+41FEW1fb9UwzKGYF714O8NxQarYPUjwS8fJWylM
Sw6MQBTxwLBjYJK8Be2iS+xj0jYJZJCNKWLI9mDnC6wAyr4DOM18K4rY23LKyU6D
fbC8FNYuTh49kJnNLgnn3fGq4Y3c3nA1MxYqsRxbstKAMGK1/Xk49bJ7uTS9wqun
PxSkXnYfdDJyjT1ABM8jQZKxWVSQE12qZjJKF9EIA8n1kgidQ1Yw920DL7ykKaYv
1CVZ1hajym6/dVDG1pO/jywki4Dz63QTw+2G95jSMu97NZ7TGkKLnmrFJ1LGICrS
zXnnIpFxYmZtaNaJrDIX4gGG255ipD01yTQPO3Mn1EVQmijK6qRjqqLY914lA4JH
DaItf+Cf3KukMFCinvMqJEcu5+uLePdJqA/pNFGNYTZzZ/BZGXCuJcDAVkajsx1R
YjiEkYgoQpwpR2JEC7Qi4u1ba3e9JZFAsBdrc5/JCiQdtfQyg2CZkt/tjU9Sjmal
mglwr8OQsgsHC3MCkWOPE++9U1rqhYio3lr78oPV6JHMrc/xLVezhx1QZX2Jy09G
D+NXIKeZf9aH1VitlPLxhUwoTk8KrKhUKrIOhytjYgjB1+1rjZ4eZHcKA03N1Y1I
vyi9JiL5kFDWd5clt0aakEUQxB+tZqYdWSradHkIYZ0oIkyi/IeWXSwfmr7Odv4z
BsRCMGR0BLP+Ct6rMuJzENDP8a+iAVZBT19nqAdL13A=
`protect END_PROTECTED
