`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uJsUVV6vQNjwxuf7OR0N7WUYfPR1yU3iDAyRxWLujjGvh3xqxVPMDpKUp08Z56qj
f8br34FXcSxPBd6TynNSViGonlNqbrcE8QW2gXdwI3SUq9Xq7GYykIPDEg1gTKYv
sw/L53sSiI69I0b8YlOv2ZlVD6P9ViRR1f0ctvEq+EOi0FFhl9d40FI1Q42hsR0V
YYHxWCRuvA+qB6Iu+WWkUo+LEUnSyPBUfQNbIrjCVO+ZnKqCezuz0NOGFOd6tpIW
9gIu2iHD6Q2VV1QjpaJjWOkuPvIiZpMIbieshWqIBPvpL2jzp9OJ/KzXICUPVU0C
Dw0hpGLIlRAltg/YCxrVTtkqytLqpdFxJbHQDNdTnqS1kmjheeN9rt+ehX2DCKE9
mPlz3h1OsCOI1r5vkWBnzDu1nO5oIegN/zfGQDCJxjYH+Ynd01blWmWrozk3H6gJ
BBMKIQe9J5sZBh3iMe7w7juouN5g6NuZx2//it8a3pWDek6YoRHjlONjyHLFOlMX
kAP5/DEUpUCUoa4WhdyqxwhMCEsvpXCQDXYYh2ywMNZXzVjV6TxG31KRtkyLKrXN
KJknr8jKv+l8RURNa25zwVMXAYnHoG5YFA4gVkA9vGIOAq/QbhnoXGco8l/vkYTt
oVGsPTAhzc7HO8NrqZlNh8IeJrVoyKUAFG/jkNlmZJTuNyrDTqw+ICmg5nw3Vm/v
K8Vu5O2rtZuuW5qDdIeTqzPGKKCNBnoUOxxz/LlJNcM8V784aX6mvt6bmxJAkgbU
hgv8xhLGwVlBYRPA8b/u6IfbYLYNLZkiCB2vwx9XChSv3k6tLcJe8v0FltFq4lhq
t/yqYBSXYMqxL1dZORCDNIVxqDO6zzSA0XDYyRLawoigPgl5Sp9DaoRO6b64RO7d
j0sFEsRBnKw1TiaxvcoAwSrCsTt5dqaK55mK/jAFWVc8vfisBZexTQJcn4lGaUUa
FhF6oAlW2x0grhkJVvCGARnp1n7jMx0h4g+8NYqHZL6QPGgA2gJlbChPEIRGqdzo
8dqer1LHFDOXuUgeGYCxnkRAYZdGu+qEzb8YlBrn5AkowTSlGa4htkBS4edcY7+2
dOB6ePS7CsrGMuXyjUznFHRUBoDfwwnDlOIOMyknqRxdjtBoKuERVP06PGV7+aP/
e4fAylt+mqgrE7hUi5SSCCHKglcARDOe5EgfPyUH8zY=
`protect END_PROTECTED
