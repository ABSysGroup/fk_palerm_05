`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pYKdWvCDS2RJBZmFKvEHA1U7i0f1RBmCuOkbefzL67eOU7y6KWTV/H9GFvcNKENS
nkMgogJs0XQBbR6IBNo0h36SU4ccMb9oAZWEpS6HCTXHYslT/z+O2X8ZXPNHbN4f
wup8NkumK99wFCyOKQmqWcdibzF0V/illDMItViEckXGCcPDiFPJpzMBNxXhsiXt
iYnvzIsqqVSod3VrKbKylHXZcED1BMQugkiyE48ENHU9kxtxv7fYhP9KVC4PZ7aJ
`protect END_PROTECTED
