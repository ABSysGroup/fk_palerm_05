`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IZbAEoHj23ohBHpfK7wQEAMBSdUBcdwYaLsZkAM5DLlBWA4/fFGq5ZX2q7OwZFdA
NPNTL+t5JyQK3id+bRxBTNbJ3hcO+Ie8Jzxjam7MUKfk5m7goFQsOUb8Vi/hugKZ
WCpdXCGwxcKZJO5aXJZFFU0Vk/1SVkIkgzPwuaatU/MxBVGuZkfDqz7PeuCCOaHx
vnuYJ8PM0bfbitqBwWP+S4voJCM4Dd6GxG0++VUVT85PO530wZ29XmxUArdIsmi5
zoRHDVyc3RB1aa7aqsAC8NzHWFWKP5JpchZbPzbgtqgpFtXaNsy4HioViiwY2G6b
rQtwCcEgubMNMgdWBmElqPFygNiv24aA0LzmJgimEvW42sqjZvkCRi3muUyHvLKA
taYlO9WX3R5JL8BjiTqn0QffZ3XXZb6Of1APD/lEkwSTTg2uj6xX6JgH0tMEJdg9
`protect END_PROTECTED
