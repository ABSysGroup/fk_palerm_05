`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LODhHY7k9Dzw3lMhGEoeY7hFK1HG3AwVX+OhpmpHl25ugtrv5o4PH8vtzVRlVSiR
yGi9lSCk7+tD9MlMfO4d2r+EMIGd58QQTYOFyVOVyrcHsrKlX5l/Kec1KGzUhZgv
WfB3SeGklq+zosUD/5wGuSmvdg0r0Jl0w2SI+EwXpeuHzeozDSgo4IGA1QFEkWMc
/VszDJrfUoauDafjtBLmG9a8HUOfEtLO7yezUSrXG1T+qrz5TBWvmS/SMto5dquA
0nq6d64DMnWbeLjxXfkV1YSAcgkB0Yo4ld3lby5UR0/IbQ9dt/zjF2iGoUfiqCFq
UaHivwDJ9WXnaoHYfiejtAFBXy93JX972mTXTIV9SH5NHQBSxjjaKi5pQHhD6dmV
siofDoCeAbMmmmVkZPJBZ7EQXcnY6QXeWw++5D1/ecRT120hNCZ2sqpg1Ix+qDwP
IDK5SXXUb/Tj9gnKBJ70iHzhZoGvA1nmB2MwuhlYBXT7crFM1OjSG19ScAM2LsP/
2x8XCs9Y7MbqffVxpJXBLuAjinITgPmCrCrM800PTfuQxofUE/38o0z9SokYYxGY
2ftqCrnKH1a1PXgusOkJTtC7xtGVyyvQiqG460/D+HlniwmC6R2B5nr166gYYcc3
P5PpExgegUD5sRatJ62dLDl4sypIhLB6O9N6WaYXaep+iVvjHEKSexy7ZjGoIGx+
oBmITclLrEqOURrk0SpUwK8sKM7YnLPhA2wmf+xX/RJ6hdHBXRKjZkaQqFbbvtEL
9M0V3eWM1FFob8vzMJcMtL+W1DvOiizFXXtwip8qBmyvGx8OAKe4pLsNdkX5pTBU
`protect END_PROTECTED
