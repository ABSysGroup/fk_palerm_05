`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KScehmW3XL9bS/zabCvK9bunnioVPwXUrMVB1LF+kPDFQAIDWWWLf7X0b8Omnzbl
bPPPkB4In20gKjejQoDFgwrG9aSNGErzQCYMYgSsrBtqLKb8Fp3BqvkERfNfI7P8
lgeBr6Zf2dgwJDO/70uJQD63sCGzHOKdzgmhfGx6b3uWc/dIpQoVsQoTRm7wYBNP
6xNwk9AQlZyY4GDDiNhkjWBVgrz15qEC8err3ysxs6GB5YCWbGqJ7r46+CPZHlR1
33t5ldEq0GdGyBn9kDh4nRAJjwYuWxCMQibO/sL10GNhMBkt0Yih1tdxgcBnFBg4
`protect END_PROTECTED
