`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q+ctEVKg/kUTTwhaIAT4v4Lpkg+0tDE3+dRSxiMkmr0ZR8INgbDVjIDyAds3+/sw
zQIJIXm+pWokS7dcgRyqOPJ+3cdppslzcQnKrLXrAxlxtfJdbX3+AlgGsokWRl+G
ht9pskrv+hy0NikzgcSB4P0ugLzqBkQg+pLvCUjSUpalgClyBgtcuWMq3NsIGMcO
BBFDv7yNwE9+ZJHW6zw/qcxvV5HFmDhk9Dc+QyP2jArb/hqzqHinDGXX4moUJece
ZMeRMv/3oVfUUznnN/VqPStwuLz/r3nh1hBT7QG3hshhZzuNFGgLQ/dVT3T+wa4G
RAAa7YMjeyupUqzcaE+jog==
`protect END_PROTECTED
