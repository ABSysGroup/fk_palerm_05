`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
evYrbx6L6xGxCuV44rDz4hlyOR1flUn/M1g0dkivbCX16pFl++5/G9rbSVZ6uGBx
/VIopx/B0wLCiaQ2RkyQZ9TT1NMd/wQosoLDcou6k1yt65LEjaVvz26oUsrizaLM
WpUWsdu5FJezvcmdlJeYF8zy3fQWZmk24m2c57Nj17hMRiqA1IHKz/HqmSbGoH9O
+1FayqhTOB5h3+VmvOcNVAUF/XOvofB1hdCKGvm6dWV8mn2Efj+DXeSLw3SLok7a
mnDf62eACn7AB02CcUsX4CfYYovf642Y8/dbBN4HF9FipNl9MdcZU9/aEfQkTZMq
fAYA95qVUqSVgTQEhxZ7JlDfJ2oCjJIEBLg1x598FFJ1HVshuh3Vma87eZOz4kOH
CROjQFtq6R4ZGXzDAx6oajjWb+mCCEzEIZnC8dOEWkUNMQaSVQuHj1EMgF36UUUM
lbzFcg9eTUCCFpRalmhv4Hj5E9+69cj1iRPuvBOzWTAi5uvCFReehcPaM03YQM1r
Lig0JLHbsEpS2QY3J8gaLLqQaMpSb0CV7DxJlt4OkAqGEFTAOMOLy85QfTOdRuMB
`protect END_PROTECTED
