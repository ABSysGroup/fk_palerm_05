`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6NR4FAqZVKyasQ/jcWyFK04lOzd6QEAHVvlRq4gIWUMytSrXyXdL23IGdIYrXoDX
/1zt8HHCpvXCmOiB9yHmpEiOczmiupcnhsbvZHDpu2WNzyECHr73D2sPpuUo1pLi
0Yhapc8r3DxaYWBumhNwvA6AFYktL8pUI4CeXT2hxfZ0RArqXuVPkJrvu5uFPvJS
krZImF5Xth2ezH28gS7UpjzBPnrxGxQh/WR+de7REecvvO/5UQ6a2WHSPkNB8jZm
V1hxaabNJLcbo6PtI5cCzXa9U2bLanJhJ5cJUabwKQfdLRlG3Jr1IP1m/oqRVgOM
D5QiY7y98SZnhQpC/j0FrQs+z5sznTzfUjJ9b3DvSj2aR8z0rug18cVvYLd0qNiD
F4p+0jC+jCcX2s8Me4N1VUdyYLgPhlOneuZLXutgo8xYW4lfOZe9YDxLf0q8oiHn
ra+j58KEFgcpJwirsa6HTZFr4o7v25Mj5b7JZ1vih5W1P3QPaXkuZCXY8TtE+PYs
SUpBCHqPE4X4n5gzB/iAf7I76oGtI2db0KRJj5MjI8/WZA29dpFbA/IZncvVKtaQ
dIsh958sYMfKA6sb4rsVxDiFH9VPui2DkUgRXAu8NlptKsciJBpHDHjgrcCJkA8K
DyOXMMlkIOM9ReMOtson5eRft67N0sv+QOHODPlF99a60mbTb5KGfMI+xE9DNzIF
9aSJMxidk6FzblacCohve+o7prvYm6qYmlejzoyiiB16F6Ex/UkNdOuOeJaX3auz
hLrhReCQykHn/WNPdYpoYPWOKHAoBrhm+7h+6PQ/OAR6ntn2yU4SsKKegl+Be+ps
JS3Z5eYCM9ie8nWLOVgIDeGDrQUo2bLWMpjFWb+k1WZIwPoD6VgfuBKPHxr6w6r8
2rVkhegPuGWS3hS56nGH7d0/lX+EpZTYRgJ0wWuibAtGfrl/Idb+gv7fBiy/En9G
ITG8npD/WK7xJXt8WTFCTFqBzWT/D149Iuhpv/FbOR7GbGOA5T7S3dblvkkcXkwb
9swsJAsOZ6qe2whQPGux/8ioRBpByQ4jfDNru8tnvV9CuYonAR4pikIqBjag5lZ6
4+iBJofUUkxYcUScOFbdaj8uRIJR3bGnzL4YP+0YSMpiSa8ho0vSVcDC6k4LCdg+
SV4HHzz4SiYaFMHQ0Ybvxq24kmPfq0izRjShJElqbcXWSPXqQlKmqkbyVDBDZRfn
vvzks3BvXK+ZQZCT5O+BYLin0kEGr8N3kcDggU+Br6sGY5RpR26eMCw3zzO03CEx
m/4JY7k540RGV4GGuhq981gqoqpmuYAAkzgsdmzMPbJekhME2rwWKezVE55t1xB/
s6ERJmF5MzN2EyYIfaD9IVRvZIRo5uSYuBDRit/2+0lCuS117TZD7dtlgewxRKjH
P9V4r1bH1OdeB9XXCA2L0IxqUi0H9luNQa8NDNGe6mPIHgSJ5sQeXqxyLDqTyNpD
Qd0xGSEI/+WiSNUbJ7rN3DyG3JmpxDN0h/LCN11d1A4ARUVI0qZ/Jc8xetALSpFg
cq6n4fcAo5Da4VRAETNCZ2MmAjJQtbxlSPNfdaqH5s7O1zhrJJ8ONvVbjKpt85Ns
uAjYUM/U6rVnhuklVRu5nqT2iaCE2G/Js7G6Z9w2reMAf4gS56qL6GCSA+W4Iq/L
EJ02RZ0oNnO/Gh/MZLPZBo8DpOxlFbbdRj4zwfWubwjgsYF7vWB5Geisr1WKf2vD
XQY8/Rjxg3fsY8Gi/6lSUkldRC42rZYyEplB7B6pehZKwH41j0SjiGJmVaqp5z8V
JAua+sqEO5Aq7zgg0DkA98iN9N+efTtnvBMI1QWrPxWSFJvdCTDH6vS5T9RFHLZB
TmBjjMDzFxIud/c/BeoNKe0minnQLzat+CLEFHc3E7jsRhLJ2odKT3YplmP2wXRd
rqckaF1x8gb9v4C6fYZBHWF5WX35xHp0xqITeS+diSTqpQypS4dCeNtdoz7DuTGJ
KjA6E6+Xdw06NXjVbcLhE/4fS7sELB7x6IqAxGI0QN+YkO1mOCB9kB5npInQjrK0
PntkpnGjBQsJvIXmVJeZ+JFQ2+B85NoHCHfb8MZpFYycLeu9mR6aAuu4kLmK0L+k
bnkAvxieQkgOJDToma0LH9PCK3h0XTf6oTU1DrcT7PBEWSIEgRV/6gBGIFnNi/+j
8yjIY84sgj0vCt+50uXFaHw14JBZGE3bBppEjLKOSxph12UR5Wr0qjgZ5h7bFtHo
qa8CLxdGP5SX6lcb14gKZuL/p01tuRewCXXt+T4PcBq2+D6GwID9iyMeCaIJk3rw
bf2q4dIduHo89+P2C97w/+DkodE5w/lTJmQuMZ2zdcnEw71jlLrWJmbfXkalXHFV
PzF8mhbOPvdqbG6nueDT65qOi87jIonV8omx0dtIZ0vDdgJ/4zuv3LnM+lEL5MrZ
XAjIewy49MPTWXZJMUwITy2IcHTNG/P6Dst+QyqSZRKb4oVAnPbzwW9j8FzC7orH
+n5o4HiUh80bj5TdCl6OwaU5S3s4ugZOF1P1gUQrGUXENsRZaVSZidZCFdcuIzWm
Mi+wsISaiAA1DmEkswKhA3C1NmTt1UdPbWCrokj8OInvrlwvCv2291kmmiSgkr+N
9SIudI2WpR7A0b6FRy3MLDFDpbExIiapqXRGH6zDLq0DM+cYwBt2sptedqj/5Oef
sMeiOcm18vXljdL6mGYTRlTMy0O/zgWPTqI5YHcpA77EdUmGUVlBJb4TnP1YikHn
SYS98LQ2Qv0bI8Y0qszhk+Q/8vqCl+rcGYl49l9So3WWYlxHGJ5tF3BHOsSg9Rbs
gS9dCB0fESPW7lA2K1XM328HES4c64TJMuwnQAMq3HerefdiMq8sBgviZGMn6nRY
Ry8FaRGWuZkhbEOMf2omCj5PVVn7OyEolOYotAKhK39L1kYE3sKDbxU1E4EPIjcv
oO+TbvQdcFNegHo/wbVVHTzoKtHtC3tWR3fwH4BzQgv91S+l+KMCCVsHFszJmwoy
nAShWZguBxo0zvbTCOEWcMHhJrLw/GGyjeikIP1/CYpARzdmaGibMVSry9tk+qSf
QEjtcUa44pWwx7x71XWy+QwxQK1e8CHfXoh9NFwW67KaSZPWXFAnvOA8K+pkxhx9
MAvhBsvKJl9XtqQXmTpKsdaATymMxUbnC/NBZYv9g2Doz6VsaEE+qQf2k0JScq6G
mltB8H85C7aL6M87RoECo2wpsZwvGS7vB0fRcp/jYTmfuU8Qt+a4PXKcM6rlsOed
83xtT1HtPB0DyH3zHI6/BXSiOyeaR6rUZyVMf/Ca+Xvl1cvivkiryV+R68v0cYJo
XxZUl4QMYVpBodYq9n5HYCuQyXbn/+eQlKxpsyMZUEsP1oO1JlSB/Vgs4oPm5ORm
RnE8N2AEQnfr93CEnMGrJs6RjyIP0FjZG5K1YWLc9Bnr5nFY5mv8W0PS5LaBcJhB
dMUkupLjttcunlS1BgzGlF4wb5foAp5IggOD0nTGYuca08I3Z7UzWFqL61UsGM4K
n7UbSgfF9FvXfzH9txSQDRrDtDczobrFF1vNshlT86rAxNRb8gSsLyo9HSDsXcfw
m+OwipkJ8hgjJ8rKvYkZVPNhoRrFuQhCh3ACL9MAUWUHsPz87PZQCdh0tH/RJKzj
SJAacn1oYcUP9haJDW3HJtPrtMB4OTI4RoHPmwH6VAHYlB5CI+PDz5653dfzn3YX
gyqxc8RtIG6nEM7xgcJjje18XmffIMDa1yE+HYzS4GZdx0MPXI7MvMSMZei3AWS5
3+RtEbJskEYt4NCGJKhQOAxpkxVCglcFKk1bHzlT4pM1cCXbwmky3Wm9kqgjCzUn
2tmFV7N2MNc6K2LgTi4QIb/lVwCh/mhtb49Ft14jXTFxIyxs8xPlnc5dmFqag9h4
yfuD6jwp/M/Cfe24YCxxgfMnOVZgG+h1NsuIYqUFis0=
`protect END_PROTECTED
