`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BLNse7cN6uIoKWIzMP7BSc0U0fzbvZjJO2haPKGc7xUsQmm6AVF3DkH2/G311PQy
eOgSDnP+nhHQnL4xquGakPubJ1G0IcKkeAdo85ej/64KgIQctgq3cbq+v7UA72C3
MpImPUpPUvXrBCyDyfN6y3SO1D/Q1lo+ZShat9JjRfHxrf1pLHzaeaO95bSpBULr
saq7ylkQWh9AXGyFbEBf3cbyRtcMNq9rgHC6vQa6ADHuDx9ETtdqgZPTiqN90C2h
48DBZMfQ/RU+XzJf57bHAZq2HmQ8DooX6lWcovBLuwm2m/ThPGOhchT+p7yfdKAP
Ai8se/qi+d22ujNSNTcuAi67J+mZEInRQI2pFGSH7kK6349yJ0J+lNBncCA3XMvA
UAykHrd3cBObibTy+4Oa8iiCIDVpSYPHnIfRP2QIsbVJIAD9Av0wzFMKRNFcwfhA
tsphBS23pFNAph/Vgq07KmQgItQx11BrwXBc32Xs3F53WA8DxlZQjmSgFsoSM4i1
rraxGTtbaphWVxb40iwAq6luoU/+4mmjbZaiMqZeLyS7fj3CM9C+dsMMaSb5FnC3
OHgriXAd84/R2buw6VvcMt1tRFib8sOkpAeNZUH+MZvwcoaHTCvJ3QkXcQBmPZhc
mqNjbdrbnuki4Sb1Lof+Svt87J3QT6p8IBQrJqZ2Ffkwb9Za4Fb1hCdLUmOOe7aS
tHT3+Y/5SpuFMUZVPQNYyO2OjzgtVh5+Czk3RFyWh5LvtsuMvHb41aU6agR1ZlB8
N858s9yc6I+ba3Z+uV1QG3omfSCX7mn/MVwx2aYHS4N75+rkxdUggFAsB2a6Om5o
ZYSP0lwaKf/oWAS9+ZI3SZNHfdK8S3u0MoIkXCAZ/MluDn7zeFNq2Ri9fjs/hF9e
PqBSuq9ZdU4vV9fR5t9QBCDnGe0PWlFkOcXsVeFdRgT398dMbVQlmJ6aB+ifeRMx
ZDYbxsJTeq4583+eW9f8wB8erSqZfONO/6HQ/M785r1rOp3zvWKRM40MVG/LTEqu
hfcnis2Bd8HCjmpoc/DvRSB2/Y6aeeqaOcBKi7Hdk9HCjkL55ZirhvG/ffM+bMX2
lk3mWlbNRjqQtwC1RmCKRgZX1+jw9aj2Dpr+bvQjrkYEKBnY72l5ZMrVYv6RXTTS
GZsmxfa0Ph3M6mjP/PltvE9I+Fd4ABAUX56MiiQAj47yca5Qa8lIy4usXgXRglGS
D2KupeXzAPZC6zAFmdXAfmK0iWZ4Cuzyir8FTVqBVujadnFEflykYbZ+di6I/BZE
s0GY7K4niRvo+ATolB+Cy8Bq/9pyXqrbBxAwP07gizy0M6F/bBI5SN08AadVbd8H
MbVuHPKAYCfNKibiVORh+oWIvHMBKBSnDyG8o6rhWislV366LOzQ8lbmI84Du6Ic
WIT7DU6FIS3hsoT+NwZrfjtHg58dNr2GJg4vsUI2k2EQXcL0rPtCDWAvrGGF60ZT
KV4eshtb3GRF7vKvaYamv8ZE6vzNjBD1K1xjmf0uyCxHgLvC0l+bjQqTcNDYgwiE
hdAoz49JdBGE2raq/k9tjmFRSefxVIHiE1zaPfP6S3vlBldZYSIJkjpw/d0VwJOX
/Q7awj+kBNWxNAxRvtKYd6mtYJujaHvydfw14lg8TXhM2g9Z0bLf8dgXdxP7g9Ng
JLxDWjJS1b2l+ejIArYUfk+ID/Ve6yGMUzVuzXN9IuCaZdq2GFgmEFk6JEO1ausY
IXvk7VsRCWnmYEkjbBPNXsqGdo0NRu1LzDBN8aBIzZb5MEJoXzobua23Ymk/UuWF
+kSdXohs1YmcHVuc022a3F8x0jUGABlk87vN/AdsHYuuwGjdt6pQncOeNegVHTSi
TjzkDvFgI55JTR1JlMDmYSxSaAM98WfhN4sS8w4T8KrivtSB4dwHvWFZLjFbus/X
0vpdhCFu3g+52SqRvEDV3WG95Nx2lK+ta19GiJLqSpAAlKcY7KB7TSF5IONacsnb
U5cRgn2tKlqb9eMvqJgqAPeILUp8lC1uU42qkzOpO/xjc38lUIQv2Hd1Ms06htNZ
azyxgXtyNm4D9TuwAstXZmWN8pmZLsihIo8SzoU4U0SsnK3irAzfSmb/YiBa47oQ
N1U+SJmx+9IIsvSA6kyke5oex7X5CCSkjCe1FoVEpgjPXgnqOLKpL0SdvHirjMTI
rHSzqcXOtt42R0NGdV21U/Z/GnBV9sY/V1ePmFNUFIAYbzexh4PiJbZK3L47UCHJ
Dp9cpUBkc7ROTdIs7D+DIToh7Idzsd4yMJLyT4JZrluVJmCkKjy4d3IN0KRBKtXh
eKv1nB7BMCZ+yELOk7Kwu8SeDrxxMONeGhfie++kMwewe5J3Y9VSCqm6+G+oV8zX
VLgV3yoMy1lEwqwgvTTFkXiI7wlweIcfib2ts8IL0kXi8JVvPN/bDZb6tI9GhW9+
tF7GSfY7nQddnlN/A9ITP6KndGvlpySPzgKg/lvG1lxQCzUJ2v0to+r8ITT031aK
ZyvmFiCa4gTE/Xwx5Bb8KEzxGp2E1J8aG755LXpO+8gzKAQppQkUS+i50V9mnKrF
O65ADHwjirgUrYG6a8Ed8dX5c1XqRYf2xDeA66jcZTBpDAfQF0K+pagMAH7eoaz3
G7E0dpYsbuewmQqGnGme77aR8U5VKm7Vao6isp76UTNoM8LpH34/B5fbq/gzy7Ev
zLcA5+X+NH08HscYLCGV6dlZThLLLd0D6ezwmXhoG2jR0aDrFhSmI0msHnsUyFe1
uqqx1mPuIEBR9Cwhehx9PTZCL0/6GcRP2sHdJtQyDCacuZobMGOHiLVg7b2I8A4I
Vu+zcrbo72cWGPGwSBBFofjIX7WOuitjncFx2eMN3u20Aw4YAdnqs/Td+hcPFMNZ
QN9qWt18zIijbGAHdS3c2itacbRRVjunDoVUKlmTe5BVCg95D12ViUvJtr59hnOC
jldfLwOtBuBisJnVi4EngBH7/vQC64TlItRxCrS7TLugqhJtQr2+46BhrkW9mVK3
WuLCzvpbw3iI48k75fqfEkhogjFUutOds2eJTSFm0RQz9gEW5xGEwvjdavXkhAxs
3gO/LgVP2qO6F9sbXTgPKxPhhaoCuB2f7OfK4l9ohBx+KP3++oOrXZoL7rY5xstj
8NAGkBEiKuig7Jl3CF3wgu2/xfJYxK2Wik5P5eYw3r8MUgNT0brpeVDzvPYiPdBL
ZPZggErfyrE3fl72T4K5gaP0fZG57Kskyab6a7jYfbyjclCPvaPJ76NMyChAowV5
8tFn3uK9T1XF96na/taOhvLy5Kji9NBVHgK8rCGGi0zbRALnCkZLf1AZyJzKzFK7
`protect END_PROTECTED
