`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tb/5ppurfqyGcFpBX5Z5zsawSTGAlZUyjXLUeI82QQ1cp0SakOwsRyV6OG6vphxN
kKCV7wc8dANeHG8SC7yPD7WTKshqOjvM91k6ACFKqM5aFWGyiA3ett8EbTGGRzW8
owtRrKdOiCzOz5Gl1q3oP9lvUjNFbwh/88r2Vlq1ozn4/h3bzP8cJmocD8hyA2Td
MVElBfDUOeYvm4Pzy2NM45r78DCqbwtUx82RGYX4UCni4d4I0L8u0P0rxuPtaNud
DxBs0C88bK4jIdp1meNGRDNa7VLYUNq+Hk8r0ikx/wHYzBw79mf4FOvUWL6UQYdV
QaCLxOr5J9DaTX/yB55gpe34L9ywf1EfjfgHhk+j9Gue+0GDivGLVdq7s3EPT8dc
6tb9y1fV/XjhPW78BHZVxonM85dyle1zpdY+IjYY3Z3huQCr2QJYsf8Z+q9H7vSx
`protect END_PROTECTED
