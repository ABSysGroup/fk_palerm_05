`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GBYNTUQE03sYfSaI4SYcKsrn4rZmyaaLTSoTr1mFDV7JO8X4Wx4H5U/msdiaHxzJ
1GhuUYei9YTXn41KoEnP6K0XZinRWoDylL5tUkJfae2LEj8HDK4DJjU5xIcTmbY4
tv+251b2njTwukxQ5Gtc7EP1dMcyPQE/yvqaHcxdVXe9ycoVTIH87PErxf7GuuSF
0FpOC8cyBuX6cMiTzOBPBrl+kf5gK2wfQFVhaBoTcH0RROt0f9ix6ea+hGNLn+Il
3FE/9PXp8QC5qa41nLv5CGVOTgCvvrSe0Y4qopAIr69uOYMZsWVMfeXE/O4kaf7N
JqkLH0nIau4/8cdRWKFS53rbDVAKHqsAT3vHMzJsi8wjPi5TBqUzcNjkPcN8Uds8
/Yzo0Ovp9Txv4KD1XIQN/EMoDHkqLX+ZBpoKiXHTPWAJCYrgdEzJ6jqbojRMFUbv
6Z0aiFa0tn8FY/GLgwM2kNbgP0XfpLDDF6rVpxwXS6GxlJ+V3gMZGdf3IvMF0D25
iIx3+YZXoYZ60gaFFVozZvzjG1Xdq/UwjSqkoUqXfusFUN2j8yK7t/qHQeIxCoih
3+QdcZGV90DWlqxzuiPMLPD91ojT7DoVdVTGSxLVK2Q=
`protect END_PROTECTED
