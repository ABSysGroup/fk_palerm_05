`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kGXdzhuadnnP27ILSgxSoHI/r6ecSDp9p5rMShrUj78sa4lJl9e5BO/EB0SOKhqo
kOLQ24af6+nYpmHFWNZ9ThJxWHauekmv1LcChv17NTduLIJnEQNpjRxMRHirBH9X
bLDb/9urzq0tlgsJwU1M8KVwoLLc9tWjRKbpnguuM1MDLVJhj4PZd024OryDAua9
6uyGGj9frZkC0+kfQ0YLKbtqxn7h0ziWPLR3fMJC8dQzie0Fvq+pNw8Kam0fvjBQ
P3IIWB6RhselRTsX8sCsd9HvDw8RKK3rIScY1OXwbYKgwln4oFJsotkARVkmBn91
QV/jY+9aI8D9k1vNkQqtpfuQGWfghujcn42pbJH5TsK6mNo9uTQL/RbZ4IrJp1qQ
1da7RTaew/8qPnbS1BD5F2HqW9nJkLBRzIrTW1yKxfLQUiMk+Wv1CKiwZYt282Ma
hZxN0VDw25JNGy+3MEJsO617Ty/5bhUMG9GQ2k4KPmkLRu9CKDjJ/kdVhABEUCd/
TNDr9rnV12PODUOCEztxK3y/By3qpkUQPMqNIpE6KnI86OYT5XYEUiPIGk7vDj8k
wPIlOMRZsI1yrli9nMrA+TUpJPgNW2yiuZ4qiC0GMCHkAkZ0hdgJL0g/sZqcvlG/
672zMEbIwcaWjgDVa2HJNrupGs5GSh5VHnOIKmPtZ35miOVYeAGLKH0dinf/v7cg
Rpeuk8huSXmFj53AZCl0ZVe7FobLDKYSUkTe7uWdYs5qcyIOd/N6VWsbvrm6QEeG
J+qmEzgpyxYL28gqciKzR7gK5/o0qqKPwHMsUFw7Jua4OYrd0jRBEqe6X8aopgqF
riY+UTmOtN+BMD+n+Lnrs8kibv4xVwUgK+eXiwBCzCfcuXJFrkhscmBCcVAE1Q5X
bhYD0nmKjw6aij0fFxZZ9aAQ/AanQ/Ws0Fc7a2x29V5EB7QqKva8F/TSvnBFeuc5
OgJvliYpLthdmwkqeCPvGLQfSvT1uvYPxOxHfjfRQnKrZwL0J0yNGZKCKtrfNiwE
Hn94OjLXfD1R7N+uTbEDOM8ZpMQ+8zzCkRW1Yfbe9rtLJ84ahtjlxLsufdVDB7AG
3mKY+0wMrTYjGoT/DTSW/ueuA8VUa+d3E4zoXWfoJFRfdbbO4EU5A6KQhjJOlCVj
RON3gVQb8bM85AT1J0qdqIXdU+ng5EPlntLXnI6/JSrctTmnx7JkKPVOyuFJ4F2x
7eOT6vPQ6amxe2L75DQRgdvmURc3AI3za4yw88Y/L+hZbM5AmKs1sdlw4gNLfQdv
k48MtVGebkPK+X1FA/SndpBRDe8Z3kCFiEl+O2kzkhfB+K+iIMlk6jNOe41sckci
ghXS/os0X1RHQOKLmaZB7lhaCDtGMFpFj7edyzsUI1cQ9VJaTzaBT1VGakpZWDX+
rzW0QKMw1N7UFzJP4/oi4m5LWF1MSn9jsSQDEUFdXagP1+aAmrNlZxiWnGFIRbml
0j+X760KeKNJaEbB/IqZ+B7X/tRq8ROomG+PW50H5NmnrRu2FEE68BPNVW1VaFGL
lEc0rQEdzdGkd1FQHbMo1TUucyodcp7L2lo9GCfIGyQWikAt2Ij9Pj9AbqtodAU4
qyS5eQ4RX2ART606TjZ+LkL9EXCSMeliNb6vkl5twjHTEI8lljTdeQzRTG8aUViX
XoIRmds6kQM+ZF+Ce4TSEtgQDDnNBQXZH2ROPLfeaF4zoO8ivSK9NaYhMYvBYgJN
FYewC/IJovaCUFwNLFZh9tv1K1lGOEGX7GTtMBGIqowhGRo3oo6x9FrLDM4a5Ozd
oGd4iQVo7bMMjVpngpCfjaUn0enaK1trWSOj3Hv7gzDcq945GrMWUhYqYZslMrA9
a4gYLpZMbyJUGgE4nAicHEaQJnaD9IlqrBLlh3N88e5KHPSu56FKkuPrxJ708/ue
GI1Wg4iGCVtrGDV6s5jHWM2k3MD5FzSBpHZKmkk21UQGc+mDriG9c7kiX1OL2lUD
0bnBifkYl66HKb4kjp4uGP2t2/3niFdzcdsAS0o3/GGGS0IEqv0gYsI/104f7MtO
sKbMTF+FwyPmSHVJtm2WYoaz08jWuGxvpl+a14JYGUPu7J832JJo38AZV0TWptTu
DO5fBJv4OXZKgANPQz1ymtD4r4ak93nW6G0G8jOqEpqjFW4/GDd2aXvTHOFQPSnG
nbeK2j1J6rWD36y4o6LOX0Xhwv373tMR0zmflj+vAQPyBpGz/xqa0EFpv3oKzYBR
FAJ2WuZoBddzSS54UjYArrPQiwh/RGVx5gcfKUxvM0yX8vP9zI9ouxZlMVegaQxY
c0vK4+swgq7SBV12QhMF36xvZ8Upbdu9RYfxj4tc8pPGMxdIQt74CE4Sv73okgAU
HaEtPBwDUP1rHsKckhdnJzNxswilJ8v9O/lfX2tv7QY2PgpB35uPtEA2uQHNq7j5
vnfOFsQG2t++km8hQ4LvEP13Pv2bT6vyTF9LUYZPlhziw4AmeA85d1HW1lb4F5xs
cz7ltUH8w2vrEjkvohyoZWNb8/8nPuyNX0rqq2BwlSSDJuBeFF4LP89RPEPLnJgt
6//v1sMeM4TRvbxJbXR2cIcdVxBB56Tk/AoAx6oO/N01j9uCbU1Eau/vNiFt1572
sj+KY9mKuOo1Cl+NPmnzhrGh/G01PkDnHgY6yaC5XqYOFIM6TdGDpeA7C/gRcr9a
hLbfgBPY/9Zm9sFHoeu24oAY1Ckw+G68eGHmMyejHZQ3G8EuTdLF84LxyII9Pkdx
UcP30fOqbWIgHVbJfl2rFpHsLt/MNiY8SAcbkZnTznQXQgzTQEPJb37Qr+jk2jHV
p1rpQBr5g+Nh9yoZ1YneDAD/Vk4Q4x+ygaHmTq9H8CBpXjSBtpvfWqiqWZ160UNR
xwclsP5raIEEShjPZsWM81uK1XxQ9xGtaXmXb4ibS2/u2gNqSniFu/tcutyqYi8D
T+cZ+5BrwCD1DnHs1hXA3o2Yg/wzmyyZ4vAbTYvy+mrQfgDbkY7WlkNZAasRe0e/
iaoEhH2grIadK8XL8Z4+Z6wWpPwthYjQN60AoBi+RyvsDm2/chHRDKfcYX896wia
lcIBii9Mw5FASjMAK+LKp/TAT5VAYQNS1Eg+Erq9khOkvJgChbaL4WsVuplIfhcv
72+ERGjSh9F998x47cmWyWIiiylfico76PxAFzWay+Nma6sb63OQ4OVCvq8o/rgE
pmaLyO1aDQWqWXYsiKBWmy+4/7bVRDI0QgZNhnqxKUQ6RxbCgMDfOm0lPBUufzqQ
c9jhEegJsilPyrGAkBJYViXd+ETC4h305ESP3evFdSV0tEcI2v0hGhMndTotZAij
JHAGKuZbKKNzmXJ8tFs0vSDjOPkwp6x+fWcwn2iNL59mV19yx9UyPDwEvFISLirU
SHxorogrC6YAoIVDX4WRcWFqkO2DZvXLe7H9H1Oc52F8Xdqp+aOD1ce8UqcNlxKp
s/qIL+KooAq2TKlg9rKryz2ETJqxkPxjhxQ4ILQMrPjEO0Y4hsvUGYkTH9qenQ1p
TdRlnjZWHVMvJDcZhsCBN8RhwqHtNsSQOu6M2WsdU3zomGlIZmkMwaK5qH3E9XLi
I+u859a2Ymm7oimGJoqNHY/KqNX139FPq5XU3pc7OV6IEeaI3FmLd8LZBDFJ7WTy
7d1HiriXFxC68rXsqnHlQhLHSsbbwaok2UjaRJVi2frzu9Xa7fYNHPfc7TFomXSz
5cc4w9m3Zl40L2/2qwcGGuKSiwqOwgFszawWuWDn3STPFMv6bXtGgC+XLZmmokZv
aKxSF3m4QaTzzJx68xLqOCbe1aMoUbacuEehsitOCUL3KGTYsa/ttmJ+rw1RKUVL
2QmATBKW49YMicykplHS8KmRXwJX/fD83s5qqzvbJuv64eCQ/zasEjoGKtkMdIoZ
GZ4Kkjm6mDvhWubErrk3MleZ01W/2+0svB6yfn9oen3AIW+H1GgYDsFDoGEV5VhN
GgO/hl0HZvqoBgq0m77zpdwtc3rpj9n9QWrSBx962fs1tgIGeQPoFbl1DSl9mNNh
izo0z6wDqieKQhPwlYWFovqvxTbWk2cqr9GFzZz9iBG2UmObXiMZiwEM5PQzcrJ7
mMQcMmzXV1eYGXf/bvjudTTSRokLKPogE6cqbxqQnFxy0hB8O/BI8otz4w6JX6Ui
zkSs+R6c3Mz1vfwNvLclIhhPuCHhY2sCpEcnQeN7vqimwfQEH6/1Be5IRvW60sP2
LtQjwfrsD4MCgJbAHBoQfRia9SPneXJwgbjcwdBUf8VO0W9O20rZFww3H47KdNQW
wyDzXVgIEMRdlHJxxXfL4FQtVBhkbe1yWz84E0NtoSKQgzxeZbIjoWXyszERSAFY
w3QmKzfYf1NlDjkAvQu1UOovzB8CwP/siQnBsYvou2Tr/2X6qG0mzg+Ph0TV1rzw
qU33t81kshh2iw0B1GJiqwk2SJPbFm9sLLsgkT5gekCadbvlfKgzeN92d3c5wijh
0twQpc7YXr4lBfOA/qFhrWJ3LlPSPHOSKg0iQo62EaOHuYWRQNKDLSwLE9wtQ1H9
qhBBdjHEekmk+EVX/AyB0EAaXjrSfWwz4f1h576e6wOatSqtgtiRMb90TzvVJcs8
5Gl0/aloTLUk1MeEn0PbHZEFNkCCUqoMvPkxOAVrqiiqUW7iU6VPieq3zS00RZzl
/GA0hJ/aGcpf6LiCL/NNyRwdg4scGZt0iZgQ8P8StPWip3eVt3oPzibgzIhoSbiF
bsGWnzcZuLftNwseJULBhkWDKBMLfaUKfKjd5EKXdzyswTUGg/Uu2d5KvT4lP8Ng
FKW7LSCPsk2Rw8GVPVBz33+OPEdQveH/SXlUSg9W4KnBcFoBwHqMn39+QKN2+GJU
2JTj2+6ttn9S2gSw8Q0LH/zzi/GjdewbNPpzfaQSqVdxgTbtsGILuuwYeyh3R8HT
WgW6ppFdoRSBUtjxlWUwEnk1IBooS+kNV0J3laywh6zbFLEWcjdNfMkS52p7ssXt
K98fkT0eWQ0AVjE/wcQ5E/oy8ZwfgpIcDTdRloaDN0YFqklSZ/kfsXfsn1GhuACh
VvhUN045nkjvgiWJ/vlQ7CVdbfU7nKJBSIOK8fOqTAHLVMw0A79VKtZuTec2jArv
eUKzLKxv6XHBFSxFvJAumeupey2JCX+Gvqk6ghlEZ9Ih1JE693Y5o+HBVkVaxsf9
6/6wOnX9ogZiwMInYmIE8Nd6UXqjbU0GHIY/vas0IBpj0REHDER+36YJpbvPRU7Z
RK7p4YQjyG6jppMAjyBIfr0VN+aAcrArVPQmkOPe667xgLCp5TM43GDKokowf7jB
5zxIipNk2W3QIRfoErDN8a6FoOIywh30qPxz3rtOk++iM3UrdutDVGlRpu9uc7qM
pm7x4kRUtBgVnn45s3i4XPbiZEHN5/6o/14LOUi/EeHgonqSe87Eg9ztfGZDsoXJ
fcCOxuRxMTVAy80YP/YDJNwggDp19HxVpsUfIh15+UZbMscn/aeu5M3Pg7kFVUsi
vdtAeToZqMINIep+qB3026EOXyFPALGNiV1OGk3EZlLX24svMhM6TC101vs+dnFS
hrJ45t0ctKz2LE8wXt1eezuYqb1DwubGGa+iRYijw8O41RMGUGd5lP6q2MOq/5Cx
CLVqbKlIPgaGwuq9ndCtLw8PHUEc9Kf2hE3fNAl/tk33J/fyLlstl9d0IVsc391w
owzfRoMiFvtoHQWP+3JcWA+s6EaInE797leQjeBggbPSEZ11J7HiDPv1+WoPpjx+
pHEcv6BOk3Znw5C/aA5HOEorr3fnP2Waj4WbFODznHt4f//FsnvPWX0b9Ys6f6qU
5LoWBmlU47CGZJKvpj/2kkjaoCbaeLboyc0dS6ieTUssa/E/rVNA0ZcmH89xv2n7
OFB3IPHQNho66QNyNUNjq6DPhFxdOLUTofY3tlUhqKX/vi5nBWXE/OMDQJDcWlnQ
8g/TY+djGWWLYKNOR4lZLoAbPwo5IARVOfaqhQtE5KH68RNf2nEItXcvXkbET2tQ
9RsG1uQf5DSYl7aw0Fb2DZoeVGyNXR1Kr63jMfOw31oCZl4blkziQd/W8e4Zszzt
ch4FC4YAVIXxJx8TRmk9orRo7QeZTJJU2oGGNoEw8730s+5zJtCCrokpP4jFgNrw
JFviukw3nL2H/4l7WD6hu9UrMQuZ+rol044Nc4R7J4OfLYsos1WNj/5OGAP5eFBU
wexVXDxmlvxSWoGAWXn0jzlj2U32GHalY9Oz+A4ASnTh5BBU2jADNa6LZWMtMQ0P
ipMNyBgzcnZW+qNRg5Z0fUHPDW1KwKzmel3smHRh3Re4xb22gbSx+p8Ex31V7qCX
ghLQmDNMdrcRsalnRDdGxns8UkncUQ4C1z8b5ntICbOesTbBuHkf2UqhSUjJqU7f
BCkXiOfGmM2lTkm0/a7N09ekikDq/n3xIzzK4ehzfoZMKXCrPzdgRo5KfriQQ8uV
IXjtqsVTYh2ZTB6gEeUcDoGupKUYg/C7nbwOPBhfyfQrlpQAz1nHI7NqPOf/copd
y496Y35Fn93hwMaXqeyzTpgUQc8xhjCDoAoSn2Z4Ab/Hgw03ZrjDf2IeDJLmHDK9
IpKkVmUs2biv1azUEo4kVfjZ2WEZkk5AcCxKfJnjbBkTKFDdaLABzeGyJCyROwZF
do6VVV0kbHplQvqbozxDqQQmYwz5OGfJnsRCkXMSW0ETmQPa2TcK12LIEWn3YFgT
TDNKs3eRzVVjVJKXpbdEjhNKAzxhLbZuAwQOxs1WGToe5bDPifTkplIx8JRvTP46
nFPWoQFib7gqfb61CJ2AnJ6K+xc8WGywFxskTDj3RZCIEmoCEnTEAFvkjoIXm/Cg
4N8md+cf9mG+pt8Pep5RnAcVhhcawwUG7HnGuUMY8GujGOmELx/YS0HNUS5aKTHp
DUejcYYcePisVzi4czCxdc+eswVq9ciiTV9+0+JrLtXCyAA+VyXWAgaWVGc0m5lG
9Wr0JharbqvSAxFf2dWDiWvIGYK3f1dqKp5f4yS9lj4hsl5AOtVgZu4SNzmzCSDA
7G/jfAZBdKDnxHNyt8taa7F9nRwVmj+1QpiXamWUV72DASOs5ij22z86m93LFmZA
s1MWVUMFraPAXqhACd50xeKaHIo6/ib4pMILrgqkWHdnghYxyo/z1tYSVeHBIqrA
+jEFoNoBE7lk0do6MzZdINsbK3UGRZspOD2bj2crl7iqlumcuIpOypRC21F50d5e
YLms3od/Q0mq8ZpL+sRixQwRrrR1/ERBoy/ydiUaLtgMSBocTvPJNzFfKpLyZzlz
p6ulOTUM0inyA7eJQ423VG0+haukeOJoiUsElvcHDRC0Ozskhy1RBBX+8+snUgiS
VWyB9Ys23z77rdpIKtQbY8fhSNUOiFmOnMRO9dUorCaJfOM+iEsrGp5vhv9GhIT0
h2ceOQTYJSlm1m1SuqY/ieaR7G8FUojnax8y71lBcfT5wFMOyh0PvpKe8cBbj3lX
WrgLJP/it5a9LkRtzws8HVZvAiDjMdf3xQI6Lw/lpFFd5J//qG/4GW+ET+X6nfes
GA/DiQBltQPUUCAp/D8ot9U4sx83vPk4k8/I09J5JLwTNWiSd8dlXap4BdsStYZ8
Oamp+iiW7EP9pHC+maiYaOGjtSBNZQF4IS8HJd/6xIIWH4NlYWIoNwcL3Sbke8Sv
VqI1bqeYjF6+Rkst1+uFt9KCtCl5uA44ctdNtMprw8MEs/HwbLRKpyafXPIRuU0F
vPFYS091sesUEEgmndAkH9BFXstsoD9npNYcMhkh6PS/qd3n8L+16jth2BpQmvZf
JUx+a+uQTIbWGV1v0byiGzMXRu41sXbyeO2epcQu2SO7IoLWKBYiKy54A4j0wSmf
Rs4HS41fMeKhfij73Q6ULFQBU6xefZi+tXNM18kTuBftxCVUZVDTmMVB85uhl+7R
KxCGg/imueEV9a3qRCU4dvtthqOXW5GQPqHoJaJRASYcTxHEc0x3YBxg24tWBVgJ
Ws47iIqH5xbjLYTLpiI2Noene3YtmkmtkrEkVSR935siZF7SVDuCxzxSaz83aNok
VSQ+FMbx9tcFxveDBIDFz0bP5aCveqVfDeJI8LbbJYbRZMSgm+9bov640f9Vsm7f
z24osjv7NXZtspbS04VCu7/TFnZ1iJ2BU5wfvQAeI7WODLOZ03+Jp/hqBYaOPpb7
laCMk8Ory6iTDr6S6Pkkt3hG7En5EoqEC/SFGlbDxXX0x45ZhHawbK5lW1IQE3YL
0M1kUeq6Tw8Aofb2vCUkgh6QvF9wHhzf3aYy1XDd9zLhlba60r50zcjS6+Kt7+Vf
SKGRx7FO3fmLylNmrqnmVVAkTGEMhwDwasF/kl5TNSOhpXmVNV9I6bsGCNbHgC86
sZF5VEROmURAGxmGHlWB8kpg0MV4z9tZZypQKONWSpn4qJHE2v4ndsaZMYmGXE5l
GIs9YsggGEadd+JG1wZuwM11MiP9xucNxLqtviPWS9T2O2FlOz7+lX3n8XXkJhAX
bo5ySO+yZFNgoUGCx9gDg0PoBMGJJAdMS0oNL5ZhA7u16ygDLtuvCUcRcs8SSTFH
HlpVqjT3ikkOXTBgoK9d4Xb2A1HUeHgule24PD+50Bv1PfqUMUuIs5kHtakEvrFI
IKOdfgkVbQ8IBUnqe5qmTceVJvPH/4+JH8zcQupClLS22aTbHeAZXuJur4Jw3kZx
8B7xqpNmSjwB2E5PcycbI1E2rSCCqNAae2FME6wn0s/u5DbyVKV7+u3j94oSpCtX
Dn5v6IC2D0/4O0AHPb0mFFtmEUfmzbYMQvIPTSY4zfZ8VlFU2j89bZ8bu7PQxpg/
6gjiQOyGG2yQ1wY1D8yylDLwT7aW3lzrBd2kkl5vSyUi2LiXqFLxO1g1ozZLN4kY
VBynmSgsYbXO7Tn8Cj2/+GtCD+MsNxC57nctsyl8gkOsBIWIjFkT8ChdafkX6REs
AYiK3XeTxI2TqVm+in3/cg15PcNgWVlpB3AnLHqtj29zm4uo99s3l55Z8WJoLORa
AOfNNoj+6iZ8S67gcbM0JisNjEc9lXAm5CBFuwAMW7dFp8BUV0/iBH0MqSNNo/He
tRN5Q0ybrGG+mkhY1w6iQD/D9AulOxZMjUrwQNPsGrqtk5/Q60DR6zOZZk4Iuw9m
I5Fl5l3FOMa4Zr8YOiCXCpQ7I8QgMiuFOnvilGWb0u9oF8v8j7HKDL6SaIXPcE8h
XPpZtHhyqATgfWqsHZkaE3l5miJT2UMWJUVYPGSTvu/T+jsdYHJfWR13Fq6jayBy
B74ad3npxhxGVaI8JKZldMK1e2/Tgff3m80uANX0MLUXfksRZbvmnafE2BGOhSQP
uKMlboAd6uSnOhuytVYGKZ+53cLTvKQp38ssl6BLYpg1uYUAdF24Af8DC0QIBRmZ
zw+bCDDBNXcHC+ejHTqMcKD0enWXvWxY3JRft6LV8fVGlM55yJ5n+t6YINbJuOvC
lBdCwE7PIKaP471DtSP6aO4J7ZkkvJ9ET7Snf2419wFH7DDus9W4LVTr5sBK94bi
CK5SX+dBJVWCIM4q2tdQrgBoHd27VLYuxFmS9CLLVhsRF7JNOYXX/4S6uq+Nlhun
XJbYZTS1Uh8nP7GDzS4RMbfRxtTqZnSk205kH0auheublveDzPEJgwwMflffYaHa
0CByd/VSwKL+unhPbJpzYmSuRfYk7h15luqQFimY29h85WAd3AZwztXoh5fhFiV4
uRNKQ4D/TAemuvfOnbxoPxJTgvF95trZAgmZz+v+gHI7IAmAtCwtF9hTsFLBa0T1
kXKdG4oh3ZsYY+Yq5HtwT6ZJbP3bKY07EYnTYUMhZbVvICDE3y5SdJLvT2Bvm7M3
ppjqDjUrUBvkemyJd0mUDlzMIn7TBv/cQUEmAPOXTX8LDFp4QXihh/A/QoEiWGVI
h4IqtbIKedHcP2qH7EWhkitlh6/sjXaJ9eK+g2xOn03uS54pJGux4xp7AoLWHIPf
tqQK8tpipA09oZzL0dQeTD+uM6spgddU2CEnXFfbbKCurGz4BQ1Ec6vPJLkQv8ii
ZdUcc+AEJ/IEUmYjyoOaJlvtZqkAbPeVG7LVAVIgufkGnqcRtWMivblMB5AdmF/+
Gq8bMNndiAdV3k2WiusvK8YPNkxGYBpIKU9TOQI6A0pKw6vIRTXtWeh9zqSHJFBn
R+gjDGIS5Kc+fPatrlJvkQQfoE2w+jI/6an9dnvKJknbUovoQ7BcOLbWnIwGS0TX
QPAOdioAEuGk4pcKrnxGKaMcAwnWOWvr09Vtvh2MNOrlCpycxFiAb2tL2CNP3TgJ
DA6Y3mtBWATEt23WVK+McV7fRHdIl5lUCBwOw7nOIMhKsHvXh4ANPEwkQmAuD846
dwTsSCtoeeya/ACVhe7/iOjjbDnoQYG4Cx9jS6KWDnzSKW/g3drEYlQyWmK+6wtp
RpVZwUzwLSXpw3CfjFwKcRc8mTBEG1tLrRLmU9mRLUUaA22L5xD94Za1PgGA/Ml2
AqW1izLBrSFkB4GcFiQdqTqsX/GYRwFWcx8AeIZTJlhng5oJKZCtADh1u8mdsFdz
2TGcx00qBsdwf/wEniPRMXtW0PX9gSqA5hjxUTWz/QnNI3jPR//CU6fe/i+4sTx3
Y9WQY+Oqj5ygbYtPsnO6xeoViLLBUe6w1hOwjpVhZiLH9eLX8fE4as6AA+DCACud
4+PdkJLugmIXZBfhS6VFR62UvLcitqtmnV0ewjBv9ha9jm4BQMRwfXnzv6/7PVLT
q/JLZjJoi7bC7QuVklXXuYw4+1S5DRZt5SbfvdyV72xmGP1UTmu0d8rWcuqGdDO9
tXWqe0xa5ORURXjnatAb4DDbhjQlXkPCAjXz6LgC4T7z+g/enkRqbX/ELlv+0ETT
evX+860q0qCuNEAxaWPimjyQA5Xxh8YHRR3K6c9nft3O7aV6Koj+V/fpKzejkF5w
PTAcbFP12oGwIlVLVMgnAjoHD4koYf/SOY/gJzQfyATspcblJ95DnoZ+pM0Wvuw/
TSF9dF2T3JDmQA3xaDIqLfcY8SrUeL5hcTLiKYVmSLPOABj/CX8JMSEyfqE5rclJ
FbBsChwuB/ytvc5mVVsChhP0vNoPXSQccpN+qrI3OagxW+bClRetujeXmZuNBpOy
TwuA7wOm+zzj2jcr6f4rOjt1SI1m9dDmggvtfNzvU1hH27QIpN7P6n45RBVSdoic
SxpE7+7K7cJ8wNkuHSp0QlXqzWDlg/LH4m1FAfzcdAoLVs/WyTe8J7IVuArJnpLu
52SEA/CdcU8zGJ64aMe8IkLLXa0FY7CIlzFDrFdvHIlgVRU+ujdtwdLf/wSHfXc1
f/+KDljB0x/Ip/cM7hCpz9X5T9u0I7vtCOxGal/Msd3UCpV8kP7SeChoQZavSxRS
gokCJUBKhLYCgFewL7fgnKUf+6+zBXuGY99INM3biJchpTv3F3r9hGRQYIko8Zsy
kav+Nej5FLajY6QbxVDpd5cOLpzNgIUP029crwy49ZXS+aQbmrshz/uahwKAIVu9
vjFok1sTvbEudkQBy4TFuLcXdxEj8UOk3n3VEkFNVAjblPA1nHviRhe+3sYbVYuZ
gTsIuIX/3Y2PdIirswfsURy/j8PoTzEU0wgaFyQIUyR23Kx9OoHviRRtFTPHxS6D
j2Xg2/XL++e2oElTlwPWKmToW7UhDMu2QDhdjZTzX/8bUvoqaip3owVYn6xVG3vg
gaJbKCnyS0MM3OJvM9A9FoT5+q2ckteQ3yZtUKNUK8C9RLt3qIs/3CzJlk0mejvP
j8f1U7DSAqNnOBZxkuBBKXE2h7F50eeFF2DEWeEdZnMSheJCBZ+A/U6jv3rkyy9j
c5jA/LHBklB5dnQF4kuMKoWkFkZ0xp6vGKwG9V/VdFPdPDtaQweN9R3ucs7e+ZAe
XcNZT+ACY+yIkEa2mnkkpf3gikQ5Hsq/JvIeWEeJdPNNlghkO5B7ASvuJ/lgu506
AYD+GOZqDcytHwYN+huHMXqsz2mGLJ207SrJQ0NWclMP0BdDRVpkc9GSm9/A5yqf
SOT260uVftA/+JM5IJIy2nKTZ0WHMS2yPT3PUnmEiSFUIgUfzYJcLUJ6/aRcbjpz
5XEcWQZ0gXWt5SVzyea6G6YRYaEJAvP5bcK0/f/HwMBopuAgiRvm0MKI2/0/TQrE
0NMy6/yQve0ogjIXST6alH+CEqrai6IXZLx7XsHCIPsJCA6chYVUo2oWf5DbtAen
lzhe6DIgN7zlz8vnVW7JOcVOxkAa28H2B1WWXaDK20qDCvHJqxYZJSR6dJ6ampGH
qzgCcT5xDvvOKFoo3q9lllsT4ncCk2YZMBf3x6SNlFhqpoi3KWcG3kcWHrdVIFB6
UbS8L/i1bMZnDAe2I2dpKae0jV7GVy3QSD/J7MT6c0JF0zdORn+jWc/DVacX/quS
+7kH5sZ6JZaCKVRVGKq4My7slkdMWYX+S69nVk8BOj0Gj+xnO1jkR2VCkYKVDTo8
zpGJBF36iBwEfjUmpRLq7oJA8cKlyNMCrQQ5dlM1RpnDuYqkdVg3BGX43+3feHO2
2cMoMK8mMwkwiqU6aOS28XLPGK/zEWsS1JSR1Od2DoN/Ae0qHOqyFFQs7r/pJoPa
jTakjYjD3x+4/CwhyowZeYUe9bRXAzaC91hA66c3420qxRvBTH2RvSx2ADl4AxJP
LJO5ymREzLeNXstEZO2b2D2rvvgGBabaQN+PxUQwir2YQ17ovtjWSyT2FpGrkPfN
3KId82JR01eO0xwFb/zOMpcBsV2pEHBPYobC9suC2E6AIr3hYssEKFtajCy+RKmx
+u2cS8Nc0QfbDA8z/z7AKQE/lFUgqBvHD52gOMITsmts7qZ/vOlDhxJ+4ehAyU9U
/Ai3tfUwxI5P2tTSeV0w2K0rIDowUkPQLR9HmuHikAX897gxsPCI8FMvTlwzLgb0
5ow+eAlkYCb02dTDZi08j7Pp737IM8vvzcThKLa35h+x+5nqHZysZDrtjjkoKKg4
zfouDgSeONp6pf4IIegU4oCaw3wKEQWPcEyAyGPIHYw34ocnCPLF4mW/+kAdvXIv
i2cKlmPxKBsj6/OmeI4UH0ndUzbtSfzOHsFKFCrbVU2MDDm664VDv9NeO5ma0Npl
2nF4u2shf0GhB/X64mDs9ceHnAf+D5pP6vxtyjhMHjC7IQjxlnHkfiiof6u8OXAG
umB/dRtboiLBtNaccEQur095HelwyMfsYoiMj9Qa9/gN3vzQTL7IDKO4LTwdgnZK
SZGMWsV/XGxT6pGVL8ZDhNx4kV3fDoFiYjJIMpZVmGTCZvU2+jFHA157mO+5Wl1e
wqOdgPnTNWB8ZEJFEtOuEeK8SbvPPO1fPAGUeqLAM+Wq95l0qIY7alxO/tJXIjQZ
3fhtpbqvM3mRdF7i9VOLgoLniH32W1Io8lTlfWwg1g1UubHu6RcLoYYkCSmJ1Xc1
Vhs9vN3VCcwYKdy8UWbruqSpkd6LPn+rXyjIvC8fu2rs0j7y0YtwjBcVTqY3iToN
vQHFwL9M9PfeN/Gs5gHIFtSnVo9kyfAQ0wW3FiHQdK8KL2OxIDQWPWtT/97Ep3/h
pyKFs+jELqay35cldrKtym1GXaPy91+TgbuXN7NUtbsIJIB1/SBFNTzM9esphP9D
E8BVCAYnESG3nSPN3sy+9NBgOSR7rUBKzSpag5suRDo8LzIdoH/xPbduRSA8j0Fb
wUfvfdtK4+XdZUNhw++4ui4mKUMqXCLVbizl5R6zSnZ4gAczint/2nW+atM6H6gI
QK5fi/0PPWAXUJEegrq+bu5QXOLsjegWTNHf+VYSuPIR5v1dEsK2Rme84+E9K4qp
mYPsQJqq3MIRYH0NWNXmNalGVdhXw7/kRQEtCqfS5WsP1iJKcaVEHOJZVVc/JWh9
XVT+Nv+RWrzG8OXyLrCurxjjdTcTW0VFNh72ofKbBn3gvvrxCb2XGaGtmsfjbW6R
dcAAvtirwAjA4DzL0DAyRjqp7dgS4ulUNBXP4TfUapjV6B4ZCGjCcxiDuTLcY/sB
fmJZYWUZhaDYHEz07f4IH8so+cNTeNnJETM88H2egY+gTZb6L0AJLn1QS9MNM6Xm
hPAfL+vyioC3b2weCAr5NNnE3XNIPJp8UxxOB0GUmU9LsDX/fvT4V6+9n9Bq4PP7
hVBR/9qjmi1JqIyYk8GRx134Ses5bkV0acyT4jSKULa1q1CSFfQr6xnfy4Xm+Zqc
DowSn6DxGOnEO+pikAKBbpt4iwDuim9BYrtcTAxeI9AzuSpijup5jaKFUcWMVnTQ
jN8ZZmjdYLUAR4Qj1+RDDQOq2L4fryKlnMq68vHt89KUsBytNuCCl4S2liEA+kUJ
QBE9yD6qBCWQNg8LPtxJOanoTrnPXwfJu8sJ7K3C8V4blVes3CFty1s20MB0xY8v
87nq7xfK80quNVyHvsXmNoMwkcnWSCvSz1dzix+IbCHoKaWFDgJR3VnqkZgjSMvL
Yzc0IvedFbCKW08ERLLQak5t9uCOVSUisiNn7HVevmMUn8g8zhFe76/9j57XoGnV
M020R5wWaHnvnHlBv8At/l4TGJMjA7ZzoMW2qohh4IZWDj7V1EHypbYeF2ewIpXC
Vu6fjISYosWu3tvm2DS6sxsikbKhEVR/kCjoi+NpxellgpHxiKEUI7/ZdQBedTk2
20oLk6MkM/x5mOKsD9DuLqtma9gUXTjIC3y6qeEEGF7p0pXlCGYpyqr0xn1hML4y
DNBroreYkHDc1Rrrfz5ELodtgt7K0/44E9CYuH8iyc6n4tLJL/XXCujX1n2RkczS
Ql+wDPwXEZSmlOT9NUd6imJqKmrWPuQJgX2Y0bBr5NDq6KonYwaTU8Tqve21ntjX
tNZqZzmWu2ypV/XRgaTq9+o7FsxDWhxwduvFNLTrWKIFkTiz8hUn6o1FPwuBO9XK
vF+zrAd7GJNXzwwTy1jSMyg6n00xH1KOzqqHe2T7S1ghx6xr7sZpE736wevWHm3b
FJKXsiSbi/vrcsQ4Md8F9ODB4FzPErXv/luD16ANDYvl6ouv3EDOfxklThSeGYw1
UzhrDP5wNB+arMz8u/x0V5YigoeXzOfxaBQjJHspNVuHbJ8/la/wNVTwaWTpQ5zX
rXJt1YKjZnfeO7GEPaBoBDTXahlc56L0rdqKEZge6KTFyH8f5NlTTUqkDVXpp5ox
495EL3UfEtr8eiSggiSVMs5Duyv6FhyfdRvORfARHKeO01JJ2kUyeWY2K/VKiSzi
HU+A5dr1zgt2lQdUEY4BiXjWWO7REkIX3H8+Z2c3NGZofLzaXSzmnvlkmQ0p4/7q
JMh425ityKafaJQJi9/7+cO7weahd/mGJmZDbQhZ3xJGCmnbylMa9ojTMHSiCD1X
RDPcmXkxjxaZCBeIHvmmISoXzYT/4hAh7s6r8i9bze/2YO6oIfuXR60y4a7h6bWS
vDSsEJfLc4dW8y88FXDn/p9FQuMxjG4VQBiTtf8hQDFlkgk18Y2HyNqtiIbGw3TJ
zjGJbRlKQquWqnI3ikCzTAUE03WuUaJeMTdlT/f967cZbJe3Y8ujBbAp+0wc8e7U
OuQPEGgSGl/AFXGVdEG59rjzhJQA6I9Trhwr4IxbhaqZLT3aKCk3m9FYxvC+gwqI
I2q61eaTkKrA/i1flqME8WxWE3JhRgWuB5Z/kxpMPGAmBqBAi4PTmKCkS2eS3355
ez5ueQAy75tr/9sVShGc9BbZh5mlrucfqKFABkOD40z0kCeMSFTtm9UyufxkIOzH
x4DmIKqcBtaNt2Cd6RnM708375USWt+pqrf8hmZPEs8LScTTU0O0+YqzmAUPVFaR
sx4cPGBMfwt+1Alp1tjv8DhxP/KzMVWfaD/SAyqSqo7ILATl6ywEASreTEOmf7BZ
xHFsIbY9/5jG7+RzNBvchzpNMDTME5fmYmzPHghsHmdcM5WpLPXXADNHZLGx5XS/
cPGj46zEd3yj0ILaW2Pe1++yLP0ott3yYD1R2TFx2FJh99CPLuq79+duNAqR8pX/
blALj1B8U3miUuWvbw+MHHk7cj5BHusHVMSQ8Csp9DOIqusfodYrhgZ1mMahx6JB
M2xrhGAkWvtgaXluFPq9Bio0yXWmw0PG5GDeN7XB3tusEDQqFI5hPga2bcEIAzM6
g5QZZEpJg2KgsqCFWFhnGPKqALTn/nur85ahnZVzynyzFtz1HswKJ5Z4tU2riLvW
ulWPbI7o9minGBZbvgS2/Vd9e76MOrVZP8tQzYekBSrJLuAGpASmHSP5Z2WV5r25
vwhzh0S3+SMAXVRPzWbYq/2IfxNCAngNyVoZpz0pHs/IwBo5JRgbLXS0msYjNcYz
lLCdw4qpgaRZ1BVw0ylska9yzhgMYpS92WeKiLKmTzJzrHIGYnttSgmWVMUBo9lM
UezMDKRp01h8jzt4MS2VdaWR+2mHDCn3Yc3BmBh9ZALIYo2RS0AWCqtpz0cq0n1k
p29LFV3gfquHE7WPpulKLloAvI52y77N+jF76N2iKFkd++g0LaUHzBPwy9REnGxJ
QVnVAm2jfXZLLH4+qxmiBgVSASxQwaOWTNzJSiCtwI5Iks6Nq/UlmW3GrBl7S2Iz
bCvbeJ3iLMAESPx0VK0WpA+AHGz2MHFy0rlYWGY9GIm7g5lN1DEMI2XJsVxYxHQP
Oa6uDwK4mlZS7r8RZq8+OUJZzD969gXZ8VL4Ohz3gVJEXPLrc0HPVCx0qIrMcW4H
b4ECvTmF0OXOYevEYJTTMjFtwIRv8cf86vnNCR0rLYy4nK98gOuv4Cc3z/B63Piz
4nP2pnnF2JYhRFvROWmFJynYQ+K4+VAgs7uTBlFt4gxVV0fuTmBsRlkhW1BXB6LI
LejVTm6sccEbDud2/HOQp2W1RUetBRWiHJDm39iVuSO5CJRY63OjIeMjnxDNiFZZ
mTlBcHu8rZW8n3OEy6pEeY3hi+i057gK3HQCB7+73q9tVmmNxSMCOkCgEhkErXgT
KntNAHxSHWMbt0f3Px3TRf7buOUjhBOLaOPZ1helM136/XSqIpnvaodEblykOUGK
sTXMz7/TCyKF3JTpBCQpoCq7n6kx/WGeHxARM/7ZoPjDxDjXNs4lkkWuw6EPeZ7I
8Yt4eBZVieQqMCfcKwlvPambtDfWed+HFlhY4YKpKuAArm9bHEeHd+4juxQs3Z1q
rRqhiqQzXysz8DCnWZwfCGNsrTQ2RsG5HUyS+bYrKmtgszR3OIB+HhDbrZLfVuZR
ZkYmh3XN6fZTNaIzMlY9Rn5m6hlXJ1jyL3jRlXqza7evjjxoaLGoXNvilhEmV1qi
B0UacvPtQmoEdnObyOIiKXDuqCAex8l/RvBviW/Duj/S2wJm1h39nhyyM2ChT4AN
04U9hmEJAjEy9jHVKj4yp3FHXu5jQCKcyBgSGxQku6b43xPYYtRzK70qBfIyxQA1
0M6wR23b4cQZqZYDB/fAGozmgYMrqYFq2J4NZyI12psnnHMM1meW7npKXeNxNF+B
gNS6DaSGcT7S92KeFU6eYTnsxELPrrTzpAsDOmc3bWfSxbmDFfD7kdWHsak3g4Mx
lT8EAhhA9pGvA0qizRkj/AAmR1fotSQHJQcA7CxEp9iE4uwy9J42YJjy64x5CWS+
7XImPkcv8op8l1cnZLk1BzjHhZDwStlXsRr2EjeR3LFFtLrBzhGpvNUMnm8FqDCb
AKSt7S71wjSVDBBwCT0LNfsTbRS5E6ob7IlvfDhqutk0BPVzgH+o0i62mYmK/q+w
n0JkolVGixUiyq93VANWiNpNc0sd9YwWhbwb8IOhlX2UK5OtdiiPxGdN5LbYVD/j
3yG3A686LpBbYLxAzkv1Emtvr8RVptpi75zq4mrId6HmcN//U5Ub4Le08d7QTFBE
sgex7/fmomE+HwpodF3yqFbzd+XpZvgiSKQjo6ce+Zmaf8s2gy617Efpm/wtQqgS
9iWjTPg+Jvy2jRe225PIXqi919VYLzmEYrNlOTIw/dQuxHu8YFb3SyfSiZrQ7AQl
hLgKOpxJgM3IqM6MqQ0xftkwR7nGvpyxbdwZaO8tEqDT9kl4b68qo2Y8Uu0EysVI
Ox451lPu2kSO3vtQAYSKbEhingpCCX5Ve8th4ac+sqN4/q66t3Xvx7p0xJ7Y5y7c
Oz+mk99QQoanBeIj1+18sgrUx5zS1sKyIpkwRSitQ06YbBA9HS80Me3RV3uIqHwp
/+ZKYklO2iYw4rUYeZnu9chcLqRDi6AYNRWEaE+DFeTS02+gon20hXWHbLo4a4MZ
2ZbG8grnTIMEkfoz6/v3dvrCSHXg52zZOPaABO664KywBsSGpP8EdIMUNhmhWlxR
35Z4HyFKKiji07FhkthxAhuI8mRcnKBWDw9sCcIb19hFkIQt49L5ECQ0PqFuAje7
ZUxSgPNm9Na+/r/RwwThdg9ShBrA43Bkaxq3sxaHJWdi/Bcrm35f+YE+9HPBXc+n
OEy1e2FW8qb7uYTm2EXbGMaRR3rhdxdUc5u12oz78uSNgeEyLP0HjIth54RwjEpF
IoHecwk46Qh2qckknUFRT+D/tX1W/SmyZECUQpzQre4A29SIUQt1UCD04dEp7ky7
AljtuYxBY+FJP3yv9o3UCANLUlZJ3bpGAVhTT1vRU5DhH8KsFJz14iz98fM7EKnb
xhrPZgoT/C3w1MR37HDHFuXxcJH54XrGF7pnyxP9urYj65TTfNw2MAO9Ur92dexj
9XcHbYnsNSotS6YiWlhBdFTDkYo52j+tMQm+2Bik2HcB47FQdQ82gW+AkE4BZofP
IMOx9wKjEgJ//VzUpyCYScxVyXEBdvIwhWedKm29xhNV1NsCOK0Ifbvr+mLG281Z
ikqMV64tvxyT2vJ/uNhoKZYbfEDtvaF/5irgSKzQXmxixAoTDvL8s1js3aM24r0s
FLWWtY9MUa+7x/wknxMi/bA91qZEPTVVxM2UpiziLmD5uj6x+dECmXBPaCaccoPr
TqH0h3DDu6OnWTgFtKM1ZnrxZDmCkLSqjRT2lqwlm+I7x2qfLJYX/4T0uyNOOYR6
2HAGZPfOulWHoqoBfxqGwonrtmPFC/7iU4umSurIwgANANtMAwYk5lXLRwWmI/nv
Ie/ukJcV8rKFoRxhC4y/uHlb+irk6+pVo3aUVG5drE62Bg/T/2mKyFEgf8fXpcfG
dMn9EoxFsVCatzKdJKf4Zb2ARHYiihb06hnP1TKWlEpuf2T/WjPeQ+667k9sNRPG
ew58bm6pQenUkePFNOU6WaY71g/yJpzgNSiWiB0lyiMTC9WNrxKZhZBUx89Gdb8O
zyoO+VByt4Qgnp8DdDX/KVA6QQkuvi3kajp2sQOItFW0eXJrhpDF4huGmpLelh4j
pC4nVvP8ZFdoStib4b0aebHaJdEl9AdJAqXA6Il1is5F6HJfQDa0B1MF4K3PRsJf
Z/TluXfXqzHTRhlMquHU7CAx0pdFOiwoLrPBUUwA2W4P1PKYVeaf0vbxpAe4gmE9
1LAIS1B0S/4QcZhZKbBsjEhtKGiDr+/MUPLOLtvzvAp9Xvn+j8ML39KjtLFlHtWW
E8weej9LbMNP9Pl8Kcasn00iQcZzMfMzlE9z8utz9v0MwYHhV9WqR7klB4kinEhl
hwdu+B6F70hs15g1ulG9+GBbLanOs6sk3CeSeMkiYtUBSw8jF+wE3Bc8GgrQy7Q2
ZumBNgCOJdFzIdwG/y81TEZePOHR4MfW+BI77reE/e8rFE3vThammvBtp/RAb8cg
AuBO8VFz12t/d+Grz/APW0fUG09hda6xTTx/KoldJV1DFgnaPDUBJr+WjOH+1eS+
dJaLe09PaIRFH7kRR+lBFwFN0pDW9d5ACQz6Kgw8XAroHQC4V0s7RcQF9J0Jm3me
POzNmpQte+fB7ptIM6kU9p+/7Hm2L25b5C0NV2Hur7i7HhWOtFl7x1/MqECRYH7z
+7ehCLI613x5GEEf0EpzBGAygpLZ6Ldpk2N1aBo0jchiVDCxC7v8GiVM3A6vIwhw
HmfQukIfCODh0SyIZzwFJBekuT3n/bwuDK0CpMMBKkB9MGiuvaZlZudvz8WF9S3Y
dNceaq4NwHU2L1I3az1jRZQst7sDcYORWhzimNvowetCOktVYT3MgMl2o/4/Lsmy
TxcXI4pTqa+DKsoalkjX8iHNKKHimvG9y1UfYBGV3WxBnGaj3klOA8eacJHvUA9v
yXmaWrP1G6g3YkqtsF/UlMOiAgB5r740c/AaaN3Lqc3Hj4+I0cxLpII2kQ6Nd9pM
c3xUFZMmsi8KkBbvp+WAYhGuZ6x7GzoxlnVxGuitAAxYzUkhTjPBFefXxpp378o4
i9ZsvO8hoHciFAbT7R2yB22gKkhjr4gPts4WcjRTIYA6zIQj2HUNXtfUSQdvTfxc
9qoCEz8FDs9WOFmQ7AmE4ckSKOpJLQLyRvGcMiGdsOJkDX+98hxnG+uYVFJz4fqx
QchPbkSgQTK15UeHXkWAkXG7iYPmWgM7PIiD+vCDbgzOkIG8o8RsNstpZDXSIGzy
Yr6calfDWWW0hfaZwyzSZnaHtii+bdxH9pcbEzCTqxZKhjeyqMRQI3G77yKkbmom
zha9rbZ+c9HrqqPlLRMFAyGDAfCwV9EseNYUmLXVddoUyFCwLnixV+NCs+RC/PHO
IkyxJq9U9rv0m2KZeeOpC7u/mxffMs3leynoOql8KhX0zfdP5c/rh5U3SglqMA0O
zNRFJyQD96SU/dEKiYRSGQnZ6RSq+dKrD/2GIP/lwwf5wABLgo4elSQ4XKcScsty
uUmBEStAO5LnxIutH7VfTOG9JFVtq2ggB95NQ7AZtAKbIJz+FiwXGxDSiVUsIhiH
OOswqUR6El7XztWuw7P/F8pm/EzTfAs6rntP4GKUfck6s8QiHeLZ9phauRXNBCMX
4GnNt7ubMK2rmMM67UEqe/MvCiR1q2YgBzEAHel+Kuzz7StyHfTmzAaRc5Ina8EK
8Jgumy704wmMdiHF+oGdib4ayOJUZHuv/jnmpvJIKMXuvu0M2OmKy6M/j6AXRIO3
WkWB/pR2TRprfUVk3WnjFdv6ft86JemJNtNG5j5uE8bwzO/ulNH+4M6f8fYRiS3L
/x0UGH9fuGdTHuXGYWpytK1qA3WHD9eJI+bAgM22+SqrpKFzwGUOMRCVII0+/x4g
srtcan8dmn6i6XlNZer3miW9zYGm4GUKv3lCzotzR+cxgmC8c/YyASuN/WK9EWNc
eBUTltOgW+GfL32mpld4WF/RQvBFipDaITzxQly8AHrk6EdLSwXTUyA5WlL2T+Zu
/IqeLro3lFfGDugw/dA8yBT2RPYOVSHJIHhn2srQfbkBdsuup1fO8wJERlq4tUfG
ZY7WGwvnJyiwGpkk+xq9hhP7ufdBl4rJLVSTujaCipiRsBsbP2x9UV3/BbwRygX/
Xmv3/lmwJdiTZ6loyoKMo0WdhNJPDI3Cffjjrf8zb5U9ZHomwyHcrZqMEoHwhneK
nfQd17hPuVL7RKgpiIegp5bUHg+y7Q4O+3WLqBo3QXpI3LVLE2/AZhiweojnTV+4
9RXaeEDai3B6+JTom6F/YT+73afJpUJ9xM4Nw1TtoOkpESVlnfACSsLACI5qD+WZ
6IbROc+mx4FXf9jorcW86KnKyUymPcKvgVDhzwDezopbZyY2U/cqgIKb4/0twPDw
um+TvC7hzuvWIYKx3ByxkzwjS+IaIMRqQpO6nQetKU/06PEQXyvzpVq3syVRlgia
xrN1X6F0qAEOhwBzGcSbrJyfgzFck4EDqWYVPbtbubfr6ovc1JI99tBaxJ+P1/DI
FEk62GiMU16zjRBMoiAOyaye8nERgJbgIGDNd0YZL47ls5Hy/YYhOdpRnCcv64Ai
PG2DxV0lZJ3+OGzOGQ021PbXZkWF0bkZpnjbJtehKAFe9ozrthUu8qJ9U5fUPYoF
JTop/Uc5YVMzqvI7nr8fCwDwF/UC6rAOGAmeE3c+D8AVmMxyEKQegq2Yj45K0bBV
ZC85hYMdmVXmGurvVlVAB+F11utDmpPEuAcOlmEkUp8tYLoSx6Vbpnvxa89GbbJY
VdYwdba34FJKbKuMc3YaCG02DJKJcZYWguZKf1eAyPIybLi+49aAGoGUsAZ1KkHy
CRN/rGGxladmX4ju2jBdm3lcy2WCJPIGw0mGJ7r+bkV91r1NFz0JDXQ4/u8WmI68
LbJKsI2vXMbUvfry8NYVc/6vSUG6207HDfu5g3XF9Lg0fNNwArXO5k2Dp5gb6v/4
aOgkidQei0rHrctOHngr4cGkL4Jl/0Q/NaQFeWTuhu3IFVNBOg0mWrk4MNgQOXIQ
clVkyh1bV/SNVrQKnqysvubzbmSmAVEFobwI7WNj+MNsoabb2xRuWUaNE+lps/At
atRgzNXhiMoMF3MqtlfWQQyCHaGgToBjJridtd44ebfzrbegDe+ZqRyaO6a/A40Z
nw9jdlTgE01mCHqhlhMfJMxJxJYh5PSGEuTfrY3UkmH7PyuwWR9bqLgwVslr/7Lu
LV5togq/IWQMhd20/S9Tz62Vyt/08eYEff+CnFGOLNfYL2ath8DGPXrNGzt5sj7L
SH+rNfWoQtgv+R8lwQ4TEqIMLPONgjOdp/heqlzOuGgraj5rreqgMDa8LOzDgoMc
5riYWz60/rloVcHrjANZHxe2v2PUruu3MrX36lmqy5DvywMKPqBuve08+XpgizLY
79udrqVmOzi9bTbb9AM2Qiw+MUt6lp4uHR5/0PBsgl74kIl65zqBtLq2rypTM6Lp
JL3vYNB8jGCCF9s5eLyUk7DhWhdRsWf0aR1GKJR1HBXi8wgDWUaL8BY4RhWvomly
prPFOJpmqXq1NSHVvb4pGNu39WHEvfavpaRr2LxnrKGIy+uxcqRIu2WHKpXHEUHG
9b3rYSN8vkVJf3JWlSm9UTC0pWkUOUuPA/A9OQ1aPjBbn3OWIARdmbrOROil7dsX
Pa3swl8QTe32vntbqK5pJ3G+aA7k2NwLa7BAOyxxZ+3YFvSmYPQcdNvF15smnf/+
R3Zdf7psNmpJQstFm8vbbaED8uXwkvYVNwuKGGhzKAnz/VIatlcZr5fVQ3BSSQ2i
P5+tcvOxAxIN2FFfoweSMZ+MPalisijihf3s3Yd8TlBrqspbX90BDEjtxv9sSEKg
6TQIZKmmSNDoa0G0DgXAy6h8d9RcffKKDUQ2qw1UFGNgDJ9f6E4sZGtbHvA2vrGi
Xn7Z9ro1qeh4Yi20wzrzCb17HZdAJBL0jmfE4AQAdpYnaadVPwHaFOu7BWGv/SmB
Uihpg7ehMZhZ0IOox7hBLZfHFGP9BBr2znfidTbyl0ORpSx8SXjo7DujYchbNtdI
oKHAo4/mxxx9hDmLqtztyW63stcvhWiT3aB0csFHTEdlwwt4g6z1IexgQCYHBOzp
lgrswYnrmintftK30gkAo9PzD2cNzP7ZioTXJaFzOIknDzsyXwR15I1elH9mPvmh
MOSdYfnRwwyQx2MTZ22FL7Y39lpfyF1cBHAyA5EuGgbPluJPiHVmCFQsyKSCgGf9
RzT9+GYP9gPcxT7TJMOmqHSNSof7iIh2pdg0HCFFYhgUHnvJ+E7FM8XMknCkpjFa
P3i+O2iYNOTl8q4KnKDoBN75ZO/I+cG1+FhZqKbYHbbM8NJ1ORAtNxD9av5n5VtQ
JjMauT8PzdGrs49lpjbQpRD9cEA00p0RdZR5BKra0hHqviVgTq2F/D8k81l2Bg15
9SHefzBkvUb0MoEvM3MoRlVZsuegy1lQBVniC4s3B4mqyPFtkQ53xhDNBSOk1DQt
gJqFRc8IlPExqyPTx5HwjyrGxz/h9iCva23mTgibdfKwRaE52DeZ0+kcZ1w9inCa
TKaEPRS2s4BMbAjIp1sKOFC1d5B6EwnyeJ+90pnKY+hmSz10OQNVSuKa/SgWfzlo
5ag5N9lHQOpmTVw7teP5VAMDPCQRuA3pjFt2V2AbUM2peTwQ4Nl2Nixmmb3OIV/9
gyiBV/HCec1HbGPKYS5L43tWJB+dt/WpYgNlZec3/J5GjXdlomL8Dc7VqvbtdmIJ
xwSHaMQ6G4u3Nitlky55EQ7rAdQx5qGnkIJkTCZ8BbGoptYvyXxXDKhAQ3LVELpz
UXW7R8VSy0QGwHiJJqOM3ckypJ26cqN+aqpLvGjY3cFCzgSHTzJiRvOqo0i0SKlO
CY1G5sOP7ALuROHH6dI31WSMCsc5exz8Etstg4s78A+goV0XDqSTjSJbHdFZqMB+
2G9kGsULR0okjzyUVd+bWTGUdBkMpi5hlDxU6Bmt+YtpbxhQ1e5NXK6PLaQKFCwv
pDec/8jYoS7oBjwhiOBbn3feRDxDdoavAkFdnOe84xXiYPpfpq4SBBrxeld1LJ8O
IF2wI7q+tj6e8+H1hxCbBune3IPp8q3PqD1hiDc5FIni2fbSPBHI4KltiqQp9enY
x7pS4n2h0K8DRjGfIff7oYVVBwy0z/1Nkdmb85FiPo3mRMF0f+dthpfHVh0FWGb9
8gcmB0BZEKbnssnRERfNqVhWFpd6/HtxWM9VEfOb3ZZ7UHTA8FPhqEDzK8bY25Bp
wzwJULTNF8/IKKpGExhZCc1HV2wDKfPaPWjJfHsC9009cIj+eM44l2dlicn40mHN
jqEjCgkKpbjF06ddYdXROueUAD35A/ba7zpizPk4kAcS4QK6HqRmEVaEl5oFpTFd
flYcmY7UuV4txDeu5iRKQkX0JJW9nwsxD6QO91jAGku7E+kw/WfE0tX8heDLWuyE
/4v+C/H/mCbjS42WdrJBJNGn48HXli5o8A6vdg24BHwi/OkHCJiON+BCG37epJRk
i8yDhnHpaoPxE+1IC0KHq25I+avDy8SXnPV5ZeYqNs4vov/b0TYU14WSqLVj1dEp
IezaM9B2fTWGzHoSr0gmC0EvQUA4DEMAI4f6ovGnC/G3ZKg0YFuyoyVfmP9fhItI
VoyN2BMw0Da8hWrMrfNjwFyFc6hsvhFJYoiTx0nABVTGRtGZKww8uJ2iUjglVwo7
6hztQ3sWBUuo2bIth2NRha7WDVFXY0YNNGIyxB8f17SKYIbLS6yyRa9cOku1MgTr
cIZ+icWgh0Xw4ziBJT+g8lXXm0Qu51/pksNlYCaRZTSgsxAmxMJTV0yjKxwrTupm
Cz/7FtZ8WjPNBSm1X/MbmqdAOJkqW7jtAvb6YYMA2idCnA8JkNjyY/uWzusBuMKu
Xn0Ok7w+gQ4x5ROBAstoZmZKL8CYQiW3DZRa+IAFW00L2DUBgM2H5/qRdE60TQ+d
dpL2Ly7pLp6OD7lsAy28u4G4QUsphzbQTFqNOKF8Fo9SUvHaBCn4A/p9MgJLNNiC
D8cTg6nWVR8MJhqN8nNY+gKciAaiUOx7yqj2YEiYcq8bfK35FjlVnFUki8t+ECej
z9OyNnwDN3q+BZkXoLTyP83q1vzmERE9tai1kY7DbxynvKMNqBmgeznfyIDzOSbj
5dGGUuxo3A4cA5tpwXJfnLI9cNOHg+EhYMpPEy5noAStU/DKBVE9+nse4Q5c8Zx4
rKTvc2M8PX998+TjnlCvSAuuc1x2unkDqEF8pXAXAqrcPMxTeSRgzC2OwwRoaBGv
Ysd711eScSQmnYmPJW1TIioxNmt+ao9YeMfR1F2MAU2tWYGIAkEwEKzzkWMNmnuO
ZDxWNP0m5Khb6DWKBjhVEixyyOXXMDF66f3du0LVWQELKzpr9ONxmalwYPVKS8MG
K3tEdCDMAWdbP5Y4EtBhBApVA2eyPAKqaty+GcD83NBQEyPb+YXciubIidi6d8pP
Y6PvJNARE6qnyOo6uv67Hvml4SYL4VQ7FHBMdjLOLasvzjVQvjZo08LZaUkNIRdh
eIgmmywGy97oktNEhUYs3KSmHA+uimbn+T1IM+xX3KS3jdzbMcouqmxEJKliRDmH
anhcDvlToGI0Pw9yycBiVLmmuy+DnDJivPpbusJtSZkzvtDdxzizXvSU1aWE6R9k
llACxXK7EDjHe1trw5uZTYJD1U2XgGxggQg+J0BFOUBTNfaSeoDMqUzCLZuVb0v9
Em3EyigOtnS+E+NNrfNSYJnmzhvSK/PJ+Y87WAweN+MNYYif6uKCSkrllo17s8+M
HRm3FrOdhpWNIHyny+G0FPa/sViip8q2uIt7gCn32xtWvxQUoPohT1qkTNOFbq91
IlAsSusLGJUyTnZsHeG/qHpJRsTZp4CJHTDJKq/ssTMZiBNhukrb+9mlz+Nv24tF
x3EXrQiBeXQsot8UI8Es2cdNQSOsEjNYX8Bajsy0QF3Hh6doYrYp/gG4EoV6nDgQ
EqpsaMiAHfO50vmy2NoHjEw9uGhPBmc1/t2kALrf+kds/EtfiuDoatSfPYudKv5+
dwvwkjtBOTgPRCQLBaDVzHoooRv6gM9Cv0oHeZGQftkvqmuGZeCbZbgDbRK2DRC3
cy30rGQ/MnYh1OJWOnFSjqD0iFzzgYkOHKVmOcA1RbtpbTDO1vWy62g3K/zAS//Z
XxPz1U7se14wL1OytWQeaxWC/pVvEVQC9AGnm09lY9rhXNzI7xIADgAWmd4bfY3c
6sfVIRXBc2t9lMlc04pFZL6/GYcKOU81GWsUumzpLcWQWT0LMnodP+nXm4nCltsb
wS82wrTRjPYwKihK7PEN9iQoK3C8C9AqT4GTJns1epOgNUltOXswTCw/0AiPtsHh
YBu/NHm/aGtlohL+I2w9qxEMZ3dvEVI5ovh+KkdYxCJQ0J8uzODAmcvb9iNHL5js
DGjqM/fg/9G+lJn11y4BidGW1lakJ8GLGk+F87qKYbI5L3763zdXEloKQh+RgX5J
Gx07KR567lJ3Ml/U2xkxIhUANa7mvt/l8r/bfJm1I3iIlCTB7Cia97F+6sj2vEAs
xDlmVz6wXPpE9p8gb3pwM/8fERdIF3A+ZIKAumwAIIE5oJDpWHjLJAKZHKU5I0Jp
owmSfldX+jaDaiI3RTMqNbroagoiDspxnl52J8obuGp3Q1u0DGi6vEUXSd9GCCri
zYrLnpS/ZsQSzqOw7nvOOVvanjWBc6biIBJ0dBuh87l2KIslpI1zX0t8TkgVii4G
siVeChwwNVQMmF2bKjLPH4EKbHZzM/BHGU+y+dJceSf9aKwvMYQvhfZTcWyxw3Sw
hPTpVUueckqVEd7VcbSvbnZ6CYhPiDt5pTdaIlor6TrH11wLwgV+Z+RF+Q1vM3Iy
EtFipE90k7TGZ3WGTTqjh7Q7vHJi85bjYL1BNull5VZn40X5EPZ5XDExKZL7Qk77
EB0bJjOOK+27m47sYFHDwP1+pmapHn1ihcKoyObskqwfdaONc5QhBKOkfCq/ghy1
+xKFW6dTX9GW+tPdYSLXGuhUREZcUPKgFuvXofKGCrK0+Q2/1+cSR6SmY7ymnYZl
hlD1yeUPM6BDsdmeHLzK/qEylfjiRKnp8SBm7NfTFQchL4N1aTO340ny1gHaRTjE
osnjfJPQb4MRJqdQeIZLxlQ19mXAUJllIrICe3Q7YSYoVLFrgIgs+6zUUtQKIEZE
ceNoqCEIvWtrcNrxT2kzAPtJ6InFQgcOoRyuKzRbt8VZyzonCiMbmm2STeOopFh5
nMFxc7vcf4QZ5ilgELXmv0fFr8ckmx/o+11yvup13jFdnvVkCVQ0gV1N4M8wgA+t
xFW8fvGTfYMplbA6cT+8t5jenKVYBoBXlkFwZ7YfWXe5R2tdIrl8IDpcSqoDJlpc
ngnQHrmQwQIZ4RFSvbFgXn0nXSSesbx5bGaoYnffOy0TtTas4YdR9/91wyEfNTgo
cbt5flbc12Osn7LEzCjalqkg3EByHMm+F3ZAdEBWSUP3vII/zgfAVk+xYj3xexu5
ttjV6yrF9SDbvzSAEBStJ4jUdvij+1CF6q71ZquZhPxnkYXtqdyv5hDrlRo/+tIM
XeuFr9guhVFhapwFod8V/fUhcgFBDrQnwJwx5EzOBw6nXcynKuwDvUtxH8kRmrJO
yoPj/FTcVv2C+bCF/ixJDVHxtm7UWc+mqG3dAGoRDCwdyNqKSGQaaijInhHrvNF5
SuC+mH/kd0Wlgor2nymbVhkmuJ8aIFbbypaDgRqmtZixR7BCqivfqVyb4gLrna64
VbAzalDuknhdMflFL8ikwDw8F16IJdQjwme7EHGv8ZB0LlwCCnrH4SplRMk8eFOY
bZsq1OP+jlTn+tUya/mGp4iDa1iOUfd4ZtPZKd0Zf3DKZNdiUKuHyXhVy5GVP2uj
5v+BZXbzaXzihR/BCx8kV78OYzafWvsxPCCTeLyUFNmdJK4yhm0NFlrvv4nRDuVo
YitaCUDtmDltdvgPjgBUKFMrHGoSJBaFpjGS/BmLEF01AE+iAcdT4kyn1w+rHQCO
SO3oP34DzTJ3y8AG3blw00c3oKxGtxubPfHFawmeOeRcxCljx7I2yWb7Z7Lbkr4l
3QFg23+t7MESdBSO+9hzogBxh5qKdzK8n4+Lp0y2dbldSsqsBl4lOsMIq/ebcFm4
GNYxw7Tn1DuqIBGBgoL8X2+MlABYkACArXeflTs00Ac=
`protect END_PROTECTED
