`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iuWq9/GXV/KMDkFGTGJ2/jGVW3Tps9j+uhX1ZisNi+LJgeslmRTtyz3xAJCD15fs
b9vT0czVYHRkQsFCWmRQl5z8lp0SwIxTWGTmCiNoNwjGQnT4XK2reT0gqXsUIy5j
o06uhqdg5r3uMsVR8HpMayOH3RFZ3zVjqrs2SryQcXyLbqX7EghIz5LT6Wq1CRdN
S6Luu3xzOcgAp+ZsbmeAsuoRimcxBrYaz1FyB9Qj6gnFWoOX6UBrP5nhWPZj1yzq
KfDNk4EraPB8KK2Fe+YdIU8LIdCI3hJJSiVeYnJgya477qEY3iaCPYsPaSeIyflX
`protect END_PROTECTED
