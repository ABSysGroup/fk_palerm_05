`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xTwqGDF6RzWZZOtC0s4JRoyZ+7muMykIVaxjTO1HMCUxESMGkbnpeAgBySjzpi04
VgvYUW9aD7Lj2gwx5AktNMv0hPYnnWCkhLaN9x7r5OrHP4wcd5F8jyNJ7whistXW
U0946dh6aHV7STEJ2jIjn4a2lthyPWuCVvCviSzfxUVcdO4iwd6NFkNN6QTwk71W
E6sMwLOLFIg7C6omYgbBWJUYu4OdAXLRxHIHHWwnVUqPufLh+ufeEw3JSbL/nVGh
xx2vBRcF+VtAlfHOZ6KqmaxZN6ZE2P/BDs6CaFf2sHMQHt3u1TWrNslnM5y5XVR5
ZlxqFh3s0v3PE4N/d684t0Geo+1Osy4XFDCdLsUEaL23n+6peFvZSwgJW/A7unjo
2ZdGPrlq6afU6JXqg6qgA9QRpMUmFM/6uBwZdnCBRws=
`protect END_PROTECTED
