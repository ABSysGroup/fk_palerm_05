`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QwpKnXstV7YA4p4QETBUgfCoxayp9/TROPArg0hqP6sHO+vx3vTaTfRH4OcSfvwL
xslmy966AZxGjsJ7xlyQPQ1+l/z2FAozE0n/jwEPjxugaTA/k0Z3yF13AWXKPVrY
GaerG/ugm7WdcZJqGWOe4lqCCK/pTp/OhQCfjtIZYeJZ0OJdoc8h5RKObFfgImbe
5bPzlj2UXx7joWj1h1r5nQ==
`protect END_PROTECTED
