`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hJwVeYjqJfxq4BLpLeUG7C9aHO3s8ULKrIGdMEVuDvcqxdPPfbw24wDYg/bdqHg6
EahTOMVvIcaPyOjxaZDWvvyYzpjih12XNELK85iQe4Uumv9b9vQbTu5egg0CnhX8
D4aASr3XuDVK+S7GNOoGEuuZU2bDiSskQtjEWTIPsb4jrDIZygn9y//VOB8GE8Mq
IfnInI8U7L/u4nsnyeckUi9MXmh7MN0qi+9OV4M+1YV3BgkId69W3b2OstMnuu/O
n32x0OQofZDs3fHr3UDXdr5ZdZyozwr6WGLEaj6CKd7LL7LZIaDQmRogoky2I8v/
cBc6Y9O/PijiTVjKb6/qwKjFsj0PImDtLvO+n1ZNLs0=
`protect END_PROTECTED
