`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HcKtKun8yDYVoipk+/toHZ8/C4v51AIS443MBcvvG9Gpi2j8TBgN0WLMbxtjLHZW
aG4h/HBZYArk3K6isC0XjrMJQyyDjem+uVLuwAQe/EDeDxVjc280Jwi2+aaE2nez
MjtEjsLzctyGHSoPAh9wbE9OTMOEzuCjE5biT7/5N1ua1AiYcKbqvRniMUmzWjx5
Q50FwMU+zoNZ/W/tA3sDf7JRVADBPFsqIN1H79DltIpAKxXVbHYaRn1UtQu3gEMZ
1jZ6ihMAT0YcB8EEczR8o7tnUc1KwtK395RcrgDDDSTZHE+t/hC4WEXbis2f0ByY
XrBVnOsSigvNkgyukkCoikG6EeDLd1b/vOvXJXAU/utxULKQVnu+gtLD+A8r3CFZ
AhoK9Lam+yneClia4STJ5aATTYpZpFcORT/s38ooZytTVH3BFiVRb/PzIdy8Pz7p
/RPOO9hxpsAUol7b0SGYcW7XUo+GBY+JPAZ5owcgFC11eGfK4U6GhvTM6s8fUufG
+D6aQCImt6eYi07tDya96YS/kJ3WfFkigp+wKUh4mELYhcXeH+n43dCi+d1uiTJ3
DEBIkfKlnMNNn9rfZeY75NzwP0VEZeYgmG1drnQULMeeISw78I7L7iXxWxgpgkAE
mZgj/xADPRknd76ebdG1okYofBRmAKXRz4VQFr8wuCmYx0d/iKoFiXWtYTlsB6PX
VM13pvcZPZINvKm5ME12E3mei0+yaASgEZI0HBhnepWqXhid0cM/pjYQ/hF6akIg
DxPNBcF3YsQei+yBGcHq+3D3wgREY5bSCutEyhwvb373IvfYY6k7OnmCjMqHm8Wv
hd4q5S5aRV/0gePBZaGASFLNNEByYzF7cFXILI/AjHf+5Y0vJNZBZJh/NVNKJ6SC
ROevlf1Lv3eJbf0x0XHJ5EBdMH+DKSLA6dkjQGDKZ5jhawawKGZAt+pDeIZSYCqw
joEyQnvRTRbGHJgu7JpFBBS9/59OxRUfoQIe9MEgldRQans0SLXZaKdOW0cS1ud7
v5Sn055jXyI+LJieWLwqCf5j7Av9gm/1YD1SdumkfiRQwm6AzvfxnDQVKMBuc2ey
j8ULStfjYtbvaqNfD/Rg6FUkXfucPDXWvH2sqpb2dzU96S4vXmNtpAnSrBCkEq80
6jt8yRhgUI1oeua/vxPB0/Nr0bIPsfGOwUcFAnfSXikWJ2SWf4wOFA2tTi0FKaZR
mGKJA4tvr3NfHYI21I3i1JtRyJcuGVZZJFAYAI+bFL0QgTF4zc9pZqzOQ44gPapv
q65rLLvcSRnyox+iZre6nPq2xx6/yxVyrZ3X/ocPu0d4AYxSTK+HaWCJ2gZGdUbj
f37yh6MBuZM+keYFZ4crbpnu2qM0L0h/RtLBJzxKGtojPTDdHgb7ShAYWtoc8LV0
OncWRDmWJzV/K7nf+etqksJyoYVdhOY3GeFmPKkmTol4LKtd6gRaAhojYqYz+x8Z
YMTjHzy6BVJ3VK9bckMt+T48LImy5e+GNN0bdvh2/BbH96Q78xUp/5mU/XrLL2nc
GJ9GXJpNFqAEMJ22BgZbqi+5J8ZnNPtCSnncK+F1Rr8XeqLl6nv1B5vl73pxZuGE
`protect END_PROTECTED
