`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pHulX2VgoaLHWfrTqfVMLO9tHUem+GxQ30PYmfGg3Qpt21/IYfH2aXYc0EDpYNqk
rxuX7owNQBkQ2kERG0kbZhSUCc+nI00SShw+vKw8Pg3mFcMNDuP7VM93J/JJqGJB
N628oOTX1HdcLsu8Kv/9w32eBqBH2uq2avjL2ppQEVKYMYm3WqRu8NMbCLNr3Wb0
Uvf71msV1XDCW/rZPVa+b2yg+8hnP7ZhkKojJKOabzZfalLbdnjDa4AJsRp+SOi0
3uNE0Fs1iglM7/HMBlpSZxHCaiH0/FOf1Q3DFr93HF3cAqQg/FBMmuZY4d6YCUQZ
p9qAu1A7TMcH587J9SaLZTezHXXpgnuwxLYlF8StCn5npytdC8qrBpQnjXC3AQwU
Sy7hA288w/0qbV09IoU+KTlWfQ9YCw5ceDhcJ+zDY+jcxxaaDW5WJOfndsKGvRvR
cLayGxVfxToo3zEX/g2UR0TxY4yrqeJguIiZzb0UhIob3g84mKDiEenjFdxl9BYA
yPjYMAjQb3hf5vJmLjwpEkQPcAG7X3JnTJ9UaWpd4w+Y1iojO4XBChjKQ9ynTM48
Ezu76OPQRz6fR7ivr6mM+xEwcv9Xr/YXTJmPXABjQ52t2HGLMtuXOP657h7ytUUZ
4L0kj7tCr+dfaI7FCxJQdA==
`protect END_PROTECTED
