`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bl1RK3NsnfQvdF+jaC8wRHkK4lQtGpeytFzJzCgKsnYTt8rZALaDIYgtDyNvwFXm
J2P/V8/WgPT5d92dxc2PKHKWrJ2JGuxfhV63oymtpS8TmqDHR04/4FMze3YvcZk6
IZn3tb0EY9trsdSl+AY9YA8TsV8bcnp9uoxsXZS4PuQwHKLnaMiAOmDwj+PSwyLf
swWAKFA3+xPoMOf0NjI6qKFl44Npt0W4xm01aw3atYbMFWop+JR6FIQVF7pvGiqB
svzNmYCShOwdMhE5ssniAUC1TQ0vC6cZOfDOQIH+bHPc9ABMnxoJQIZYJg+YI2cX
f3wKfgY+JQg0ihsRtfijgQ==
`protect END_PROTECTED
