`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6/vMS54umAQxJu+dITQfL2gSV763Q1/KEfZut/uK+aPFmmDEnX6cSyPaNmKOp2wD
aawzUDaex9zRr2qnpii6CCEv+cVuoMPuIiOzsgpu6X5P829JaykxP4cjKwp64YcF
Sz0Ge/EZ5l29/0R5NEvMv1Urww4pY42pVdnqQo9j4XE4eY0P8y/KDifdTmVqodjz
OjmHWPuUU1IB4ElO+66ku2swA9ULLkzCrJR1SjisLDykXVkRc2Tc9dqa2hRtHGDG
XWKt1lFGaNKfLYDWfmElsNA3VHR+Le+5+/5MWuq5zD4bubMOnooA4G8tLlb8UqZK
mwTSpzcJTiYBY8UHXccx4VqZPR/GTEp3D9UXgli6VfyL0YyP8jsWeAuUf7L409+c
qZ38IkulaYRVljLy5P7mQG6bJedtF//c+5Y10qAP3r2FcptEU8iXgaXPSywEG4bX
cEnO4uiixleT4Azje+0eA9NgwD2+csCwUgvmrrjgNAO+VuS/nmX5OaSO1g7qy6uo
Jg7N2syyMImoBCVtHJGSQw==
`protect END_PROTECTED
