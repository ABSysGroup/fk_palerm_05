`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2SYAR8hFUNCdkxCj+MBwdyKp2Bjk5DYCqvyK/wq/6BInyfLrk3y7j2pyfF7m5VIc
Ly97neP4D7UoyoLUDcvbnrjXJb9rbu6VTyioqXEH8ZCb0v+QSD0G93R8zKLWF+UJ
HWpESMk+anIScN0JlS5XhyIvkpqLkUC0EbIc9wkDflV3lm5DtUeTARdYnAUjPUSn
+6oUxQZ5pZm4DVezQ9Bkl7lNa1lk5G42MeyNA9I8hFeiKdiVHVjwPHLO/KdcF6Fu
w8hipcXBBTBjTaB9Qx4z1g==
`protect END_PROTECTED
