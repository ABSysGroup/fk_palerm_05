`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NgELhhdbrpK+kJHrYKppFm02ePNah430kfmUOSDWyRGbKNrMRo4kVblOLjeIihvB
2n3qXKs1c+7YknN8O9PgOfDSubJhuYZEOtXvD6Zg1LhFxSPvqhHzk8AoI9VPIDdy
YG/NwdnjTfDPOOXHUELmaRG6E2QZjgn9GIO8teNHPhdkSaZogMOloV38wauGeUQh
PKWre/KPlmn1md55wFNAGCAfMxIPqaRrHKvMB7y+MhCfP/bSJYvbAuJTkattR56x
9GzK9JW5JxK8nH5v7wCSCoX1dLr6RhB0cpPKwaNah3x2FnJgnJslki0rSXFUd4R9
XQ2yxESzPCdDvzabuY6d65qeGZoZrAnWZWSN0yzV2CJTfHqlFgZN8H9KzwOrrQfG
fZJGNw/5/eBOJMYocnnUbr7QMp49U1W0b7AQ+kdQw8KEx1+nKbMguMjpZlxbgyYr
9kB3XzVMFYpNaylAX6+jrreoakCB9jEIKS/lJYgD9P3LLqdp3/JgFrd9E60LFg9c
`protect END_PROTECTED
