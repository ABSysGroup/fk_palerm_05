`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2oWVRyRsnQqm92t/vN9KR/XAuG5CV+3Zhs7vJfwyjm0Pts7HndwEB9oq5BIcbsCI
/F77WwoQ5vFbRFX+q46W8KCBbllX1JPD533jSIMWYMMmkT5yw8lv+DiVre5gEdTm
3Qo4ZcGF4/cOME1CxJzISd1r6RXMcrwbucMjJ/nuTa5RXl63D/0kiI51tcXj070/
276GuMwZ5gkKAqixdmQfbocN2H9o4rq/2N2hgBHslya79cpiBmTTA1vDjyYu6o1Q
gJfO+qTzRY4x1waJsXrnGHRYmuUV45CQQYyHOVKe1j1H6PuBSU9GfwKJeqMlHl88
uJZ3/hWpRfcybXJe1sNtzgCjBPVQK5PzH8zgRwdnEz48aGliQxC+5qmJiSm3/IbZ
ssOVlPCpM/Imk7HsgWVrIlzouKsdSuWTVAEfiuwKQKlL+mULIWz+Mbha2bhPTC2a
RgZA35WW0IgnC51b2tNb3nDxXoskCfT0UWFeYxq1dYpL6GXrY4Jzs+rFxvdK3VAC
id8vQEkKuIXyy7LA5UMGtMQUEmlTa8tQOe8+3VX4iBXQRE9chiON9VoqeWUH6FjC
CFfeNPykishv7SAV76Y9ahNfOx0Ynt3rHZOwvK3tILU1eDwGeOdBxmYOSle/mzit
XlJ0hqBNyIE9GRn4hNof57PO66nX3Tf/Jeg9P3Tf+cbf5OrWemGhFmHJ+Fyg/xts
ZMU8rloQqo1+0K64GXbMJQV8rfKZMNdIS6zWxsYv9NWazXIyOmNth+cmJ4qsE4/P
Ubupl1GXqFyDAYe1hKCLMgYeUVJkjAP8OAV1voHHojuhW8Uv+gxAYugWgcYK3svS
WRpblQI2wRZGhkBYlzHwYNPw9cRY2yOEVYxWxEyloJXzECgyalloPmXoD8FrZpWT
a/gAGDC6A96oHRUA6a6vS9oRse5DFbPSxIFLcpEUgGroLTeGLyxczSt6IpujkLbz
qr8HKIBfhSGUUuyaOIXbs23qYAdGh1tV4uOBCLYRE0h0EmZLBscUKCeP9OaBuZ9C
JstdIThrI/Fx0RkDSUYRTDCH9D2IzDXTMoI8WZ4FMQh69nhGVdaH7Y4UKn3D6psx
H3OpDTO+dHdDiRkYZZNHHLeQwQNGnn6AlMsVgTC9yZwjce8dQ+CekPRXFWRiM/nf
r1PB0iDjgJIZqJBqqAeW0/lT6Y8Z0SP5YfDQX3xsnmu5Ey/Lb7/gj/5jDnjOtw1K
2q1KPfoLOyv7uvxTQfSGWGtMffNXxTPnNd7cG4Nm1O1OjfEhBCZJIMb9H/vNZh0J
qGJT/FVgOIpWPvRTovDI0HHWwT9lca9b9fzBL4SJJNS5NhCIlG9Q0LjhVmkoNBNc
aqAHGBFSiLnO6Rs6j/veiX6tVpd0pcBhzYChQlUI4DtPbf6JMZkdj0/czmtKVKL9
PJ1C10st4KiBKTATrShiUx7XVUqSx/EDQhBDak2fWHOqPl6FPcGuilsYPAOCMZ0o
L2mIxalL5iDJRgH1U0yJcCSubheV9llrl4u28PszzlJ3NGQPM2Spg58wyZpoVQha
T77suciqy7oYkyK5TQbH9vQ6tVlGcfDODDFFf8BlvaHGKoXcqxUlGELYNJW0Wbof
OBTBlrfU3DUAlyPTG4aE2tGZ+/zwwZe7Z/dNXvtgfaciyyjlZ97Ft6om65CiVXhI
Ua9frwhyKVvgyMQlWeRR9XWNegYdRsP9vZOKpwL2vJcdimbuWcYS4XUxc8bI5JKH
3M5dx7NAvQ48+sSdv23knCpW6ayGLxgbje6oM2at5QpNPq7Z47tkR80Bq3Jb3TK/
gVO+O3H70UiPlh3Wjrq3PUiP7yhgLwfAVpB30Ze1QT2/dpnuWwIlYz/JNrCKwB0L
L0JAGLoHPz7aH+b0f85aFsr6gMBkxZw4LijF0ZkU7XSwMcuLkTDIXa55Sq1ztm/R
Nvv52ZoZ+eeeuCTD5t72Pyx2kLn2CowfjwUbnhWzkJh2hIe0kd72BdS0cc/OEoMO
9u70OvdQHeB77Cu3nhDucF/mipGrxIqTd1YgERVZMtZxGjl+30SBQBslYBz0XHdm
2uOVRpDnk0PtsDnigw9mKkixxf+0AuWKsv8P6EJW8/1EkE+01TXBQawQxroURVCs
Bf0bakeK1e1TkhNklNQRhvoMhs8ypVJE4ZGfzUTaztoO7fauFJmjzVZhFTsK6Hby
8guA/eHVKV8JxTsM+dRqFl12C0AIU4z4iFD/VxqyYMh57rzgosYsESK8YZarvgzh
sn5Kt3x8E3fUWiRnpX/OBEIWRNDoyk3Kqi9IAf90sMuBgupyvvIB8Wo6A/yzZXGJ
femnWpfO/JNYZLk5E3mn1cwKTrbkpJMR8wbHu4A1/ejGtVqRkeNqGPpxQVcSsFya
eFmWe3WLyGbUvf4hrxO4zyj3d5Zs7smpJlO2sXbzy0oSM/dBqhazKOfH0JxsDUDV
I0u22xiF8VQejuHdhat2SmQjC6J3DO7I1ItNKmWSzBZHEmbIUYBfp2k/AEHmMQ4K
wnSD86sDw33r0xW4dWZ8M1hpPzTAlmWQUpBM6K8XBswVbrlkAt48uhAQYNROhHCz
47ACsrrzWjRGuRVFI+UaoE20uWZZIVuvlcXp8PomBmxT1Skny0m7oqg7/6FJ3g78
xOnlNymnmPatC48J0RhezcNqmNve39vwS8OkHY4rixZH2quJg54Lw4BckrzwlDD8
/64gTIh2DS4/iXWsKVNa5otiezLQQPDo9g2eydnFdX1qfYJWddgiIdG8hAPuqnLr
fclRFTBT5Se9sQOhaiyX4pHvRYmGpD901BllE5/BIEK+1cZfaNmRx8X+tgVe54dR
cLeo/ddW04i0cjoD78PmnE6caQ/wU7AKuO7r5kcy5MPXJC7VF6g2vek+UEmOi3V+
PYZ0UslNQPuUrTznLkT1jfpRQPcw4zOuODUf3t5x76qWFo3RbnYGH0LPjlwjddSX
/7ROswdB0NwC0LQKXIH7nDLtlHuuAPo6s769JA8Zzcv/5azwAhGAoDRl0c0KJ2Es
+71NSFs8tqBekZHvyhDq2EDgcJ5NIxiiV5tz4y3zMM8LJhJxyZpgSbbroyB8Fldn
FnGtwAnrXgxZhwzvMkbUG2yVNTi9SXVBcPVEWxXtDdNXBioNjuDRSOYjGrzI6I7j
OuDKBohRRT/4HlYs/0Dr0IaTVAxhqXg2tgQGdqMfVe+SRJy2E1iMrkKTWV5cNPOP
sD2LQzaRubltCj77BPNpA0EMTolrWvQYXfH4JP1aMojjUdL26PKMaBAg20nypdSS
srU2GKHQvoq6HlDfQrlTOQ37FVcDMB9LWBuLmM0kVgjArH3wCQPnvTJ6oxrJYulB
ABey3ukYYKMZjrZkA+5PSCtYqb9jUHmL9FC280N6NHmcw+935zBobFChR/xhK+C2
cskkvWO4zeMmBdwRV8kn0/ijKwpi3IGnKM1/so6+3JP2uKAGiH35qpiR2oWdgT+D
VSeRP8dHg04pE5SPUQK0VdpgTIMXiC8/9RJXa0ayemudmPJVLGHRxgz5gBdu4CUa
BPKiFeg1+3taNbs9rtQpjMA79qfev8xb8nLbOSvEZf3LlVUb4kZ69Ke/zUmTn2j8
9z4LA0R3tyM6LqPn/r+p1tvNB88+DfnyTTAHxyYmQYwxDLOBTirrnI1RQvCdIa0a
jGOQT+9LLhfR2tu9KIxrR+IXbzeCHNKAPhu2y7bvMmPgIl5b1FXFl4vJvVtzeGrY
eNDWbzVtdK8UzJvcgLTFNQ3FKrGI0JBdgG+CD1PaIVbNDaQEl735quodqUVcCzCs
LT3QEgRMiivDCCB1yi9DA7yzP4f7lbRzJwAgVq/z+9C8pGrAmq3IyzoRet2ErG7K
WnYtJuc9LgL8y3kkbk98GkyfYPTLjHlyEuLcskoEBg5HS5CqsdqgToJm19oS/WHR
FtwM5cIOKvFCBZBn2Pfc/ogJnEVJ57xmXuSoSj0VdqKou7z27+9ETIv0MmbSEVAt
pA1ch6ArnLXi2MXPgBCI5IwKIE+M19MSSHwnfhb+0TkUo0wxkeD5Xvts/mhpBt8F
++DYt9KWWBew5On7fZs49Y0dIV8khvNK12xDXcnG/C7EyGw2YVoJbj0cAw+LMzAL
J6FIsz6MFGQS3qzaRVMlFKT2xI4KDOqcQMiZbuBiqtAZvRKHrq/CcpWEOxcGL6Kh
W7k+J8QEDbjsHlN9LbUl5P/+71rznFqgA3diwGVkApYAwgZ8UCXtAjkEzrpzxERU
qhYseGR+p14Fpc4wy+XPKAAu15TcqtgQ3HSKc1GPq33x3gPSuZL4n+yHdpPCgGJM
DOjcOOa37jfz2EXvd52n/Z5Tpn7BJyXpDAeekgaooG9epIoWIO/RhlXdSoezLH52
UAAdOU+CUM5gpY0xvyl/UK24rTCiPslvW3174RzEywNQ4nBRKuEdCL/mx102v5i7
iUTyTpy4pYedteL5E6v8FplEN9YfDK5tEJRkKvjNnHtAi4jDBWSoExKuZIbRg979
XmBq6KQkfVjGMvb/ykQBX5YS22HlJSYXqtCemuhOQ36POwKyRLj7y4NJCzBvxbad
IP9+BLveik0lXFp3GzT62+AQ117fvH8YeHPqYDFMqlupA4ynkQzKZzS8+WZ6ORtE
2ssmbxhIDez5uG9y1FJlRgr5PRrPTauJKL1qldnhj+oDg2t2Ctvt3COolOqT4Ynj
QdhM5Oj4WRQgWVRPk3DjzVMcGbqKzk3xnoLbo1+EwDa2GeQCkfPkn0TXzskCH9Ek
IAcGwtzd0W84+CzgggUmLfdcdWHjAW6G2b1WS/PBZSX9K+Ky2Jca5/b3AFip53C7
QkMlgI9otTowL1pxmGGn582Fofuy3rLEKQ/A9imcXkA4HKPZ5kGajyFGREGfA+BH
IINkek7nT2kcT+OSovGxB6z1uSOPj5Whcc9W5HMFHYqMfVQ/wC3ychbH12NvHAL4
CAFyiBWmJ2mvyTgZxgTJTlaOH99VJoa5SfXmX1Zj5FaEel5xQvyI8Q/94WVmju3P
Ld0RFYSGPDM6lSt7cuV/gqMaxtCT1arAeC4ZNMQ5v7jlQutMIY8y300IEG/jFi/n
s2FmmYvF6Ag4vdn0z041LRLPisDIisfc4ZbYB0QAPfs9/xcDpdSKuPbcCsc4FgCK
VIHVqs3NutRuz+xV2ui/TnRLp9nT1G/+FyAVmnZgSwd5I3+puVN5NOqte7G5MVOn
ln4lDMtGt/JRoRoZ1ejRb1tMahq1DGdoEpEPf61g4RaBa83t2TDZMLA1rY60KrHs
84UpK84p3O9ZfXyOjAtebB1Gks+XWO/vL2d/Ne3meKUBvB/G93Re8XZXMd/6DlDK
/bEsTjMHH3hX40cuF43VRj1yW4R1XszKg4GBmhiQpB1pfolmd1TTMuaE/CTjj3YI
72Tl3TycVv7jct9qkIUggY8SM5saSCOv4SYVukFm+tYWsR8cb6sI+bXA8J7I5fXc
ouC99BFM7jYV9RfqmyJ/zNvY+fk4bjqTWqntSmd5day+xVCZsHg7OnsTzcVhziHT
qTv+cudj21ZA58RTgnXNeDYSV9d2GY+i58dA5VClN5/cTSGKXCf/Vs3St99hCa9w
D0U4gaTCEK0fTnn5i85EDG3gwHCX0q2SsOD2VtxWOdo/xPZxD/3Eft/2MFQia0bW
+utYeS9BugbStWnPm4ZiOPXRTB2yvFYYZ0BJhMMRe9IRUvyyJtc+JNZ3a2UmvKAg
EaDN3JhT6WG1sg/ox3KSbElaSpga3PMHtNfsz4jWVXg40m6Ys/8w0ROFQc9/72Op
KTabNrMHC1czCwN2Tu7I+Q1ZtsgRTrYVgi+uvZjrq0lCLx+O5h3JLb2pU2qN5aq2
5ojqKBfs5fw2phFIWpj7CZ3mpAl6iPI4sxhp/xPy2FCEIGSgX9rwOxlNU6BEaY0x
EiJ+vbdBifxikTTW5nxWJsxKdfLI19L6GUrUfjS7AfLjBZOH8XSAWHg1pmoCpkeM
umMVkwzyj/VezXU0ED1iyIcpHvYVOfV+TKQjqi7iEkM+uH5V3TCgljfs9XTOMVXL
pduT9HqIiHRLm9QeWFx0LvwfeFmhS7ay1DvWbGpHz4nO8c4sy0PwViifHgpCUkBZ
EB5A61mb4pUDLg+uT5IboLKC3FQKSkRvG1RHO5UF5XPW7M0iggU7P4p4Oqimm3Vy
L6gqBLZtU093j1lWiwVCQRc/QU/kP5peNDKTS+4pP+Jsm4bn8Cp3vTyple9ABQkD
fOq5ee5iHhFVMRCyJ8cPJYBIIep+gwST7GqQ4Da1udp3yEePg6Wi/nQRzC5ao9z1
6NcGv0IviNQEhhsTkJADeE6w8A0A1GdeAecndjBwZUKquN8LOESA3LVUbu6sfzW8
HtWD84WA61aS0BT6qjcKonQ8kVCYxHleMzIbLaYYqlfS6j/ThfGv6rvODM5XlLdw
/5ZCbxerdYN9E6qh5M1HNCQ2LR+a24iY6BMMrUs91qgineGHC8mCupvMmB4Jv9oy
VyBLxGlvSeUiLuEQjP+iptAqoEMFGsNs0UrShnB8ofcp2xqjg4oK18OtZxYEv4YP
HIpkL38OfJUZOl+1pkSQHegjTYk7Tvlbk1ewRNikaob4Eer7MJNQJvxDaKSZNNjm
+k/FQsQ2jdfIJWXXlXb0MARH32pxKdV5uXuZAllCQ6lQoCaMnT7Te9ZExCt9zA2u
yZy3SgdPRcUCEaiPpIWkLwa7pfQLyqXt06h9WSy27s/j+wbY8+PQoUOoKdet7DsY
wtlfLL2BjYB6vdzPBP+1CKAmwzkzpVX8WWeb2hkfJJlL/tXz3HF2BcYOLoRlXYXW
41fWtHqBhGy9ZiqCl9t2SfnW8rHB6fmie2D0u60VjACcFyeFppkCifbnlCb+YZBA
aaYMoeSRBJ3UPXBnZjcDEbJud+hsjXb7oa87xyxvFKiiQj31sJAWdjQkz1+KUvWc
az07u/e/jf9iCdUD8C2auduWMw0K3/C2SB3G3yJJv3hWwwRNvcZTCAOnC4EEh6rg
LxcVqCGtyRqpNVBUewRiL3st9FfexAFWXfwekxP36OlCgmfuRCMWdmL8mdRV4gJ5
MV2XB0iqHbVepnjgI1b2gFMb0DxygJDSaLeIhOtKuGkAytngMmlmsw/L2y7rygYL
FwYfb18bmLWXZtNR5xwfj1M93bCFR7JKOeeJAyxtSqrvSxocu19TW/U3wzFoSVOm
1njgyFGt3JCH9ootkyaq+l4P8GwZNEWSdBB1IJop3cLUFWQoY9fjbJdqNZZvwZRn
o+1/QI3ATs01Ol9QMg2kQN8DPHmtNp9vdRFDPmkQsoiezfu7y79WNARmLPutiDn7
S00Bx4gZUxLLap5K+zoZefQpSyjw2VK5RTmZnldLqgLjnsXU0PgNWExqAPVIXhMw
lGvwIAZBLaLeLBT9dRhAawCIpSiejjYdpy9QebMT/tqWTrpIht4MNpp+mmsieTlt
AXZsEBl+LuILibAUUk9pZ5tMPAteSLJuUQ5Yd6eX/vOIDoBuNxjzK5DRFk08tMP8
HRidowprZQQdB3EDpGWb0jFTThCe+trmR91COX4+FyI1LZyH46z/33R7UiZRKixc
LGyU2M5bjm5QUdj63TZmOjpIpOxDnUFtWNmNFiDpQGDfWcY05s9Z4HowgmF5Wlwh
aRxMXPXWBdT2pRi7ooDbbkXKfa0/Zdlk2qgqkWtpxPXsqhrStgrABQczzh+MpzMa
F33cVQUe7Qkx3jvL9tNaspZrUxFPnGmUiDOwxRbAJ4Gpop5m7dQGP470xg0hQe9D
L+soO7hrK2pKkVapSqJK+7dCLh0QlrViwBuxq3d08GX9K5FqFOeQNHQHSZeddor8
hnUCytOBYhPQX1gOm89tuDfqou1lxY79JPDKZ/3KBetDHYE+YFyuT/uWpFxHmuE1
uC5vP0h+nuBsdYxb2TlObg8xzF0bGJQEy0h3vOMg4I0daWRLWn2JpNyS+QF0kt3o
3slAxudDdyYYpW338IwrFI1+nQmoe7x59I/gAbGsvGskrCseP7EoSu9jHk9auuMi
72LTwxCT4B/h+UjAcJSTHtCEkkQllu9hXaasfvPME0U/lBD4u5CNFd2xGpFNv1zH
O6XQZO9Yd7Fn7Vhf+JJUm0uKelbyBwW4zQRSq+haDDPRfaPh+hKaZDLpR2ukwgG4
KJLcOE9sgenJCO0YodvnUDhv6XHOOWaT81k/+EfifvjT/CKVPRTiWC58FA/1cIcp
Ba0cfSRR3E4xsXHkmV91c1QNZbruiVUxreBzSG1aqu2oVeSGJlx6qkuI4+U1YFfr
3ru+QLNizUi/AaMtigncXOqZ0ktoD0u856SSfdxTsFXHrj4ih42IPtr+PKSu2OSC
dN/GyOuveKEYZQO4O0bZ32P2bKBu1IiLT1V09BWuuwt37+4FRUM2mwVbslRtf2DO
+Rup01Mm9aTek2c24KRO7sDXAdeNc9UN/Zn4YUfNt2KLdD0fnt1AAouYNKXsKB5U
ZDVW9MzQGOszUIbu8V53ttZLw9CEqp8L40zjyGPKqExo6yjSNn/4zepJkfMWkBw4
5AILd7c0nAbyYi9QeaLPf+LZTdgtqFlbprkleuFoyKT+7ZxD/8x2f2656kzeQfsn
5VKs+m3UU6XgjsvZ1bk19GUOicuHQHm/srlElbkFs2Rc/swvi24xmH4hj45OrGOl
rpIXHRGsrDKog83TsU7TvFPuf1IaEMppkOiHesxp0hQxduhbdEnxhDQYyohu5P4f
Q4yLE7BLX5c3AgRnnWsOg1yCtd88zzyrTZeMcmDAHiTiVxMMxpvTcwQv64JRXfIl
otMYZrUQo2Dw9deiyGCvpf03PzIzbqrVWENUb9wOPwtFretEwJzHbL5jU1dAMTwo
KkbxCOf+gxWBsM+lOIKW2bb71xa2it7f5PbV9qZmwx+c6YchRd49+YYINC4DagBt
qb4E5JGxFDrPeb1OY+BcZslHHHc++MNbG/4uVdKuzCRvBfUzjwVd9LKxZfqZP5Qx
taSBAsbkTLVUV3QH6bHUPL3eRL2wxWWFEYFQMBGwtZ4cR+iSj63aSGqpDWaZRvJi
KZOOKJw/r26WTvywKLDOvog7fYEGj6EGZWCyoOUORF/aNB+gHndNwEMzGrNppxBf
KKw+2x06zY8l6yL0428+8qtMUO7MY32aepxw0QOEQ9fsOMTZ+sNp1Ugw2GD6Hh6a
eufn8KwhKN5pV2PSCaWeXhnnQPCcgWwotFQ4sVoBisfbtRv64TfGa8Mi6jhVFVBc
g7eIMwjH+TEOjDzSXjrm+ViHSkc7N4lHxj9np9OZhaVPunH2GOJ8jewsgEY4G8qa
OQ1Ju8WV+hYIHjSwAQSibi5Ry7Gb7fsoCtHcGF81cv7mIz7R0nI5PrCRVWpI0DCQ
6jmeVeRFfN+r5o8ODURBkYIa/uG5sw/gO+ze6HyQPyn5G3jEuU9GrJ4bTwjwofg9
fFAnpZxpvIHFRxRG/hwf5g0wfx4tNFREy0DgkZjVFC6NbP70CdtxZSF9yviu3Q7F
V65QsA4KvFQnLrcXBUNkYpOVK18R3T140fe72Ye1O0V1UFvnPEf5kx2ycg0yCSpn
QUMELRgDz/39+bsAgbBrOflGr+dSptSMFpzgHKr+rdIWzcxYbEGHOF4Dp8fG6bCj
qjC0SOcKfZ/2soS7Ix0MrqQWY9HLcV531ncA/x6C8l8TI9s91xrz6yj/9M7NLLLP
m1FBypN5z6j/AEQM2eVXBBCjk8GqWaCYMMMNmv7A9O5CV/9WpD31BAIdP+SBT+KO
bP28Jy2o7oMCNDuxld8bmYA/l83RZ7K9KmN/6tkLgaucr+h4NgDfkyfycfSXwYh3
IBmHVfJeV5iCdTZGFdHqYfPepetTPOlp7eW+yyMyzarvHmrK5VpkRG1zadBBYDLI
3YuB6p8DKs5J/cocvVpAuEjLWhGoeABVO9D9DhibLBDst0qzZraJJHJJfFnJ5iZx
KuA4staiOZTFvrLvrDaMRpxQlYXDhaYrXXfbVABZbQZ5sR0OeJ+YlGqk2OpljNfy
P6OyN86gzLJYSmhRf7SqoZplJHe6FElXyN4k3wwYoklpV7qF58SB/wJRc6B78Fd2
7ccwCZWWkzQB6uvK4nCCsM+qLu0js6RcODtFDcHvQkimKTyXy7M709Av2gl1lppE
ea0kdqe5Vzv8xqsgEX6O/VX7kMWPh1wDMQJ7Gsj3+oL1omWhIOQXc8RweXYSTeKy
YB8bmKM611VORzO/GbFuewb1KmenKAWhm7rrjOXUjCNy96ONjU7b4Lvtt/y9LxQ4
ea/eg0CNGoAid2hk8Oe+i/AXIPF4pD82ky1wrwACmdN7EPA5knxd+yu4AOl2bNQz
6XqD0PtmS386VjtitjNW/s045WaZO4stCsRgd+au+g5cOiTCf1thQK6z5th3a90R
rR7PMjLsXFmq+OJU0AOHreL9iiVnZkDUQvpbvNcrM+6VOEnD0w7XWtI6a2gx3+0s
QcNivcPqU6rTXMROOdSJQjYF5iMmLxT/t4CxGhyxr353nAYIVB6sWipDqVsTqKce
5Kv4wpKKTa8KskFuRs2GIeHj/W4oAKiJEFWqZUSIE3yYUp7c2RtO+w75zgwt0X0t
2A3ZQJH2eHEgOPKc4f0FsTcpj3bmkWmz+/6BX9LEgoX/t/HNs2w8cyVFmhdcU+7f
Q2MT8RRMH4+DiY0mmpHDJA3q+9q9HDAqAuFl5lG5FurRoOriQ4yMOCDgmg3dytMI
oWTYwB8fUOG9vep6cB/lfn1uOSfPGNwPNpwBRrMhyQrNmKoxgg6o65h/sLQn/i9w
IvTpEHuM+N144Qj4nPZuvgPTy96rjMiYB/swg6UCqgG6BZxzW84TP9YNAbY+wCYZ
ZkhZhOAr70XVo1+C0KiIQO49lVs3rYxXU2/M9eZeer5r/gQRbaBypgfDU4vFM0+Y
hx3FTfT4THrOKSKhakaLnt9ZTf6lAogQSqpjfVBhVWN7lB25HKM3/6M/DMvklXvf
x/3FFaHNmogGiA7q6iJg0gGVhpE4AR6vf9buImUX5twXzKQB0MFzqZ4ArKFhMSe6
fTlMqNxwX/La2BnhISI1f8qV/1E85+cedJdKtsvwNOQzGm+5y2z09pv+djLFRq8g
JKiTlv2e3BKVUch+nV22+cKNfdMy29If6Xjn0C0duOgn1sMp9JipEifIi2v9ArZq
th1Ne/jKcaG+r7vqDV5nODXiKlm8ijx46DqfWYvXmofHnNuDQCE3zER+flXhA4Xs
jBtcP5f2mDrNuDJzyysQCmwrQ4Y4ZVJXpspY3NVWBkp8TX7cllRUEnmOtmfere3B
nSIvNavPYEiyoJuZdXd+KX4N0Nb8sptCRM3hxgAIQTQ8mgXs9N3o9Na5snU/x05k
mSiEnvLwWG5lj7tS4+y+0/+DRmwKSywpOFxH+JkYOVYV/hgDpi24uJpv/OncUCA+
A9lnp+B9fIj9vq40oUxv4Gkai4AwU06iP4LFrpPgd/Tzceh3qZ6T6VKyoUJZGGeo
I6JkQbaHT7USat89AN6vEF6W4e8hwS4gzvcIyTlODCbuiMv7Xk3brRXv3eI/HsLr
NZFKxSXZR2kvRU2+uHraCZ3QhwYbDGeEk2yX+AE4mDJng7dr1vBFQEZA/xNz70QT
2D6PhznNmosMWtyCEECOZadFy72CB1JnMlJmRZMDadimcmbRF6Bkz4X+Sx/09Zwq
ZIEKNbmKcDnTXOJJbEVjhFy2uGXL4ueH/5qTF69tCM3GfUhHQw6lda3In9lNjuM+
V9LpFPAe3uOBQg8BUx+jZdsjQTM/LKVolkXA40iN1P4RTqf9xQpyvpg9E77RfR66
lZnbuuHYLULA01Udt9F1acpDuKfAfkuqBb6cVw24EaRJVUhqcA4U01fa68Z7ZFp+
dUnCC1lhFaqdOukK1FeA1Ym7UpqWqTMA+/p6IkxMoQX7tNjOleENOyFy1gVaU73U
nIfiBXc43OSTTvCYZi0vK3g1jbu9yg2uuNQpZOxEta2mJiNtD4G+EosGUPhRhHNP
dF2VFmuL7ZIic48p5KY5WVC/RLdAqRGEPVd6tuo07Bx8wtCVPlduG+cHxD/AwSGB
aryR0YYd3tK4UbHzus4wSQroLaMCYH7HHtnoWRgWqHsyzS4zngw1Uu+oqE9RPtIb
bHYjWc+3HEtR2ZZUhzjvctF+UmM4IJYGghTmD1zgyrB9cVCKJ9bf80wmGLKZwgOD
ohuWbTOkEqaYqwkEOP+Er0ZgMg2JQ4SKSYnUkH4rayOVxlW1g6I0p4UzG0f6zfcI
amTFP/1hoAVxkh622GQ9aSKIakGsrZmVNL3KnETfEE06jFcfHWfOGXxXVNbklz8z
5xx181TFNQAowPjGciyyoPrYnmI5pt9gWGMqAea+aGgBsAI7T/UGu7v2+geHvAin
GBXXrLA3QHsaFSaF2DQJckD/SNCweTJB5rp/2O4/KY9ARs/lvvLdq4rZ5LNBCutc
s9F27N4ny3CqWCDzOFe/gnUqOY0FEGOhcDtOmvbfwkmdAUtx2sLhBRMV8YkKYMIa
SSAbKNuCKgtBKtejqPkFEN0jS+ISC60OBgH1pnBgqWjguUwBSXYPN7BVvgGPGHcH
XUobEcBIgBoSyDKmwwToAVvYL0fO3UpmbY5OBY/9TXht6+QDoa530nwRnXQgS2HG
9qW+zCfRy3OBIpOBh2IZ4oS0ryQIDJiGK3t/zBFjO1hcAGddAclTPYdl6+dfZ9/z
Q8CXf+qtXv+NnFIvJjpAK/7h+N91lLlSMzGl34/pCmODuG0eVooJsLvxpovo/z9c
`protect END_PROTECTED
