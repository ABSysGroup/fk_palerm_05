`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yoHXhhMVdEcj5cjoIoFkbos8t5RaUpqOyDWo5C1j0QiLJ5nJFNIySifMIsKzjc/I
oN/l6v327Qj5tFsObom4m/PbMxfwLfj5Q6tfmC7gMUN4raARZKbtyh73mTdP9pOl
rxofqOYSYPic1PtI3bG0pvJl4+/9UPmwT7P1aROsjIEZ9E9Qe+3iAj+6nGbM9Zp8
9AyjHuTELhgwbLk5lZ/bbAf8m4nP00svkoGLMzlayaELhNVdSVlBJdF65FJrkRYs
y9SvHSXygnCSAMFYUaaOn9JecEnMbtynDo/w0NR+0vCLgu4H+DmxDjOXLDo1rlrg
E1Li5dphAmRy8N0VLcX2IVf12WGAVmMVL6qAjgS0ZrT9/VmdeYsF9ncMEiRVfhBh
ijahmIkZqkt36Kif6gWni3q7HaDJqd6hwMbZhrAx8AUsRyzTzOOloMxNGHEcBAH6
QUNK9AXHtrkgm5HvCoXg6vRk+u3brpqkFzP9aY/00vYSQ+Pp4/nfM67qktUGcOOO
KoxxHpKtJBtChRzWfRcR4CXh0+fgL5QTkVL0VU9jzXGbB1JdngNveEBAuOCK2nxn
zMgAhGpPnky0C8lDGoi5TbgcegdN4/THUGpxPBK9GjdTQPCs8LiCY53b5bPQfxOr
qLzp8ndHdufuZepsKvF/KqUk/xDo/2YGDAux04nFX/IT00SNYzmNO0umnFMck1mS
IXXnjYwaGUfiptyecHVmjJZ0OzlIAg+CF9UZlg7I3wcyvZzu+Ksn1m+k6AIjnYag
Ha03G2NdreJ1jlb655BkyRVZo1CR6hjmtI98/+rTO1q0MyAxugw8YWmTOLKd31vy
20uB1udmfkNG4klZbJKS8u6bhLPJYdxDzlf4Wy2SOL9o5cZjfTMmpe5PkK+t6fgX
LeW1NMKmWpJKFiNQuFJ0uC4VUPpb5CeUXJEq3/LTbPk9UibDxSF6w9Hb4mRPkHBL
`protect END_PROTECTED
