`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dbhlfvx5HyqG0zhp3Q11MyHSgvcTs21JVYqk0h3pgmeTVNdTC/zGNfKm6AmeD+ie
5DCNgVXzK6VaxuZO1JPm1FTAIo/OTwhkNSspnNdRMnWYFrJDQCgIekPFS77pI7kF
rMOaWAPxwOqN0naSlU1uA/U5sq3Gx5IREFqsw/Ie1reqF9udtUaLORkXl26h+LOq
22Emd6K11fSqp3PMFnJXy03JF52I64jFgm1N1TGYc69sLwKdfaX31tIVqcEVq2kS
Log7kUymgc9TjYBJ6zy/srVS0YvQmB1OLfAWnbzum1DsZYgzMTq+11ngIMB7v7fn
JmIW6MF6cwkh0a9di1hzfkYAYf0GyiSIGQla2f9R0pdjPH2jI7P7mA8wHPBf9aY4
bFQmaMU/I3Scp7s8h5YsFJHKVuiKZ1tIHgNSdzue3bmH7oTaZ4Zf1Gb5tTPdUHfn
PwRJIIUvX8XB6/+UFYJKqOsiaoC3cjtkc9ZGBencO/PwXU+XBU+xZs1buoYAfi+Y
1WaGKrnFsLMxQrPDW3TSYFD42ygR6JL4uyBLZv/TqnF9Lm4Uzr0dIklSFBIECa0R
r0ScWRS4jSJCzuJZnOTZRMkGaUISJXEEJTYoODw3aX6wB7Ov7CSwPZThV011ubGS
myjtQ36nTX8YJ6Zl3njGsD0bBwjcq7+MGAEvYBBiaNp6j3DzVw1rJBdel7CNx6/f
ZVzHSW9Ospomr5Eyl4j12uWLUlmmhp6LF+pTayFfJ/YqbboUw+5rLLcc1kJTsZIn
UQJWXGA1MFDMoPd+NjZuav3Ulythk4n6L0e+gLmaOmsOR/4KWreccqkhB6NS31Zy
46hvKfpUbbF7PUayq8Dbo0D0h8Ku0NA5xCdkXrL8ZozuM9qQsQ1QI4yuZgsFXie9
ZbHgCQcZaPxMuDzDsjYHDG2SwCboRC0xn1e6qEHNowBtSDuuAbdZGGVIaAwcH93D
YJeR9cpZp/+yFp778okCTKtcSllitHGB5U4m/9Z25L5yF/fWyd98W/RlzLWK/446
RRTs+moSiuKn3bZhmyG540ckd870ZjM3pf5mJJyZ0xz8ZZcrP5ZFb0kKTqiWw34l
gztk/iQ9B3xDocR7Jnisv40dJpPUD7ZsS6u2w5gR4yf1av2imjiRMQBfmD8lArrq
bIojhD7HaxRvumgbpqnFd4ZXToLN57OpJSvuaE1GrxwNSREgIFnOUwodmQsOAUhB
JDIh6D+5wW+QHzAuLPCJpGA/THZkqPCSQnDZmMzth7hwn9I94hAZrE2+XCAbq+3/
tmZYePycEmSD0VijEDh2ONhKDdLl83Tyu5HjW6dX2CHNJiGRnizmyyQa47Nz9xFt
IXGSjAdfnN3rQRl7XB5IDYjTnBgN6krwF6LCmPdb6JePe0FBWU97TvxJNuUFDA4f
WEDMxcHHoLrJQbgA2R5NYgDcd4jcq/dc/Gq2d2tlTtrFUw2/9qBL4J200263cpli
zziyJOsMVBPCmKjirY5tUFK2LiUApwYaWRhxNwv4QIacIZPedsxsfKaBjRsZU+OV
9VbrxnLXZEfnWRTEMi7EbJ7+ZpC3P5Em5Ndtuf+pwYGafTKV1z8Vichd6Qs8QL8g
G6sDkQQrrZdWR6MImluNyjQH55qy1uOaS++sdN10hX5ZGV3Zv4Q/fPYINcbjm/Qa
XpKm8aOkrGBHtn+Dw4GmL5JlKvZ7rSLZjjdYRwqlntnocaZdwm4tQDD/IK4Y1yW1
vuKR31R/w9sp7OFfY78KrGt3cXwelIaNL2p3+dRhFvbIyaQ4aIln8f4MMwDsjvoD
autZ+RdaKenfu4sY0GzyG+9WhZ0eSgRW5ep35+p+qenQRglwWKMo+wnOpHi3MDGb
JpuLIrOq++6DcDCZ6RvzpoHF6CJq+5nzJ/MQQCUOEFoZFgSQ1AXfaX1En/mFaPcJ
ay49Y1OyAeC9MGaUpUXU6LzM/rGsZB5eHG8APxvrzSpdYCydILMk/qh/pNP54jry
JjOYsXvhb6gf7fe+w4XIiTpuYGgydHXWTzazHbGvigmz66yhocucOnLluucoyhFn
qAXbLiMbSdkC1nu1evScn8YN/YUWINO3xdIT6aHbAFpgXa0s+fjqyS0Lj8xmxyec
maV8yImZLN/z+9+otsq4cGp00WHB3OPwBmWJs9VezXmq5oMBgGJ2eIrciyKpVQWB
sVfieAtIftd2oykAMwg8yuphECIhg96CUjCVSH/WNrh55kR0eX8TjCMrb5VLOG6X
xB8Gd7NvyK/2ZkCbuLh7LZfwp47QjUVksDL+vfJdVbCZXDSgF9JSS4nc7agBrWMi
i8V/oyWNAK6p36uik6JNJ7G3abFDZZxZqhA9YUOqtC2c50Of5AeHrxiX0SAluY65
mRwMk578ysJtp9ND3vHT+3km2xMllfwXPCgA5qfDBkRaG+ufpzmOVoRTfWljZ+xf
dNMuMo/uHxSf6mc6pUQ6cKZUQ+RoJawokR3yXa1tkNbZBOB4YcXlXStj+EdrJW2L
tV1pofuYQJVHECxcJvSN7//RuOS/lhjp3b3jouqJcoayTYgRpaEdwlh80w0Kcq/O
PmgCWQ5HKlQUEand25T8OrYX3PcM9Wao6EJbhJW80X2S3vpRmo4IpuUn256OMKca
vYU7aJbDXuC4T3IxaEKdE73VEbwc2b84MqcLrN39RmDxkJX6uhDqCcOct7+lNDU+
L7v+QJjRkhKKo/N078T8tcr1RGNSzwY645lYd/bIdbypPioHx4AHoIxAkLKnyKld
RHr3vUH8tJT9550xOKWtN9kQCg/Cu/RKhBjiRky+wGGEh/ftViXZb128Amqq01Fd
UTWhK+ktnwYxLf9U90U6PnhxY74/pjnWMy4xjEaOFA+Mlp1E6thGKFtJBI8/f3ik
gB4sJLA9JYsm81qOYJTv7Z+2g342UK/zDL25lY1bsRt7Yk174v5Kly6YAoiGlAPJ
ELSbnjla3zuuDnVZVfRD28TAiHPa3hjcLgvypHJp2n3OS5LBU+dijNiYZMmp2DKE
ZFSSHgezRTmV91OIAiPc+ockbz8GlxbZP6/Rnw2GLGuwzFlK+6tPf32b9M8SKA3l
DT9d3LidFnM+6GrcifTzSvx8noTMalIbxT3eKEo2/lRDUnkik8JVTyy7zd9tRfMh
tyZIBRwWBTlBST6hlrYkImStDCpody4tK5tbSMxzot+FsCYDK/KdyT65bZXrDjmT
lGv8OMEOeluMEgnEBnnkl5Z8JFYgObB+OS5qejnWIYDOOKSXJfm6b1JYGEszN3z9
sTmd00fHaDUu2qAGYpa+ZxZ/IB3nIMZY0SzgUKO7gociN2MpKU6KFSjV+OmiGRs5
/iN7ogZePSHRVHbaF0b0ySd7D7EWo2obZdpeYv8FOB+1ST8ROGTbEdJ0dIkzRo+u
HefJK7H/gp9Nmp20gipcje3ANvp+UJvNJxqw+MXjIqwkSLzUXXub2wesqOowiVoV
Pg+FwT2RqTeytFEUB8TzmpmV0xVcCSGBBVN5q4hu9+tDXImjhEJrelX+UD24danP
7w0CUkaCz3e4Dsq5vKjt2U2VZNcaYiNJ7LWwo6e7TO9Q38isA7FvJ73PkK7svgz6
t25CKXl31ydHxiYBP26IoK++d95MGDzlDH3TiJZ/LxUUYFEk8tfotsdurO+e3Uiu
KU4XwbjHiDDmrkCh/uLjh1jcX597RmPuSyoFVejlSnb/VACjy0191REwUS8qj+Ys
C0lvV7GCoWXT1gOkFq2s7fHWFIRPOeQoBD5OwMIV2CEk/JsPzOS6mofkF1g52WoP
BnxvzsRIap+Gk9/4EzndmTFjPTWjozViBmAmaD1FTujvm5t5QOJfi3N6hJVd54CF
RBQOPYgiehpQTchKqO81JXegcUJQk2xp0D8fzG6TrilUEPQRuUqiCvOBrVRX5QnT
Hv9FFpD23E7mnHyiNcK7bQwegp4+cr/rZWOSniY1qVUW23OlLvU4TbtD6niZXrhN
dBAvmm3c+i6cerBxcgzsgV2NBIMHMcSe+01LReziRenE+lSDeLhq3PyESfeHtviq
zD+UOnLLTbuj3+usg4wGj/eOhCB+5WGnysIoQ9UuGt1Soui21WxxQzPHrJAMHKcy
Gd4o12QJlnHmepka9fhmvw6I+KEuOjEIppnCazF2YASN/rgVxu5enCt0isbuQubV
SDw48WmhUMp4XJExMzjJa8bANfrT7q55/7aJ5T9huTiNQXVmPEGL9dhlx4miA9ZH
T4aat2QxmDVAc0znbNRKHEgQrILQr/y7o1nBu2PYj2bSYmiawKOrfAo2hpvYIjgb
tV329ATqObKp8QIOyE8xuIHxZb1NRN3ZuIa8NCClKscs1sYWJxsnlBHSmX9/DOBt
40mXnB8Vg/hcScdzQ6HRSFk69nOUK3Qq0lC1OqBxM3ixIfYndkwq4SlX8IpYmYhj
dhkdbwQYUBY2duh1siqPf44NjyTfdTGIJDVX5QnC+SnYCJyk3dfVFwcRYygLNRa7
N45GRH+HxfLDdhy5zRsNTPoVDQeW64DCVpC0XN+IWWEfBOAOK79M3AFP4aeU0brK
ygefoiF0IyFRVrGlLW3xsocD5GIrNZ3eV4/havUw5VEeB4iRsDX6PeJIFDpIcLlj
YOg/AfDf6fmfWrvcP/Kw1UPqZ6GGysvz1HZ/cHHD0I2sBA2CmqWbDo1+q/MjsEfR
/Qkvm9/grwK7pHEhgVftK52+AOxuBaOonuNYhCr1zPjE8THA8EnD5WcvabMf0C8q
1tBN+FNXPpMdQVynZI4i1YGYBj6jf+TDVD6J3xbwKzFXA5vlpIw3ueSVis2lG07r
Q9bjLk9EgJ9SfctG93gFYUd88C1csEaqi7f/mpdK0TO3eFDqOT85z74rljp9h4Bw
UNKLL7PbT3y4lv99zuskJ/r5sGXWFBSbw9w05eIy+zKdWoyndiUP73DvpPN50bs7
HCWI4nKrtIZpJ/KIfwrk23TVVuC9+CCGio5X5MMYwFhuqXl8ExFj2FKRiNl1WBmV
c59VKhAK0Q9y25zvER+Q5LxtSt3f5S0jdRYBniksHRC7c8AIbHciTRbl357ymRfe
58oPGRK9RtOHJX729uQg7asYEpkkrMRcC7/Ucw43w0ETywBrNSHwyrzt+nltwgJG
eD64YBYaklY2odwHu7XhSaEWiKc9Pt+DEYiuura5ovGNdyscWnjZyAIWAGlH6L0N
qpRo/C0KQLL8HfrRJ4ZRUhR2NrAAlRnFKyaXB4JyzuPB+OUD+wyKcJW5AFqx/1w/
+AEOoZMP4tTxPcN5dgzuobnJURTsCa20ZrYtqJ/4HW2bz1eWkmXmZNLi4Q71/y8f
sXxOKzMuTN9Aj4jsXUXuNRmca94fPvZXrQiw1eM1IMKZQ10SFJJp6fC5oUd/fBYu
VtKHHzypLpwJ981yaJf8K/Yi+luVU2OllJ/8FNW/Fql1sCWvMNQAjCcMsram7F4F
CQO1R+fSS0UhYFnNLEVskw8cyBlXRTQf+NlBmSIXBGBlDMLHVAAoU/R5qa5tH6Ku
lcXVfnM+lJFZVT2/6Jfl4+6s+FjLhx9Q6G1N1Yr35Zx3fQQyDZ1QYAr2Ma/qf+Zu
6Npva0kFSG/tbzDM91X81p3gzFf4r9zruIstANXc03BzQiOxAu8GZVfQImOG9Hio
TLQ91eRhMYYtY64N+m7yptPc6jrhzam3C+YkOEBgxmkNooihmx5jYjlsqnF89rlz
8uQDOLN4IUeaB7nfRk5x9LWUA7eQKMBOdAu2LEO4GLSasogILRdaYcSUbFwK4ESV
fuhh9xf4RRinj/gKrk8PbZ9x0EqjocpQgwbU8KmdbRo7JzDF2hQ81qgyzk4RDttL
9dAfw5hNLWRud/CYgW9nS68xMj+JfhqXlVgsPtHTYvv5cjKQrchkum5r18QvLvcL
CI+zal7US04lm8stAA7o/TdIfFAiGwZWkrlIucl9zmq+YfYd9OkVGi0D9XB26OzW
mObpTiPLT1pX9ZVhI62b1pFsI1WHWD+APAtd7JbldginyzREJ9eLvTSWkaKS7+zr
Kzqg0Dx/C6Mfmw33SxakPPwpaQp0LVSuW6uxzHBwPzHGEvsQK2Cnus5t18akTJmC
9Ha4pTzGT+TqWQkJz+ViwCHOa3Xw9w6esTptWDYi22//W5iTjBlgy4tqGFXjMu94
cNZCeF4q3ELHlFd9FBNGfI/TyMsnC2B+cwQDj6aFjn1h8lEjdnaDJZgEqBFKqvJS
ojD/x5oLIBmi0TjBMDaxRVhRSiFccBHPnblSxnAYLzG8kzQOped3FHgYV/tNhu96
sT5RvnOUKsPHHJBe/TXhJdUlPGdBrbVJea7j5sKfhL6u430Kl/0NuYlzoUDXJbqm
x6RWklpVF27Z57ESP+B8wiiSu5dGEuYueztiz4X+8kyR7xEBs0dxvQ40aCCojRAa
JW7ifQhOWzsQJGFFG2tMbmQdScC7PaGYjTqmaf8kUqc/vbSZeKLqOVAYYcAKcTSK
mJtVaWcAW7d+DhJSpL5tMYZy8iDvt7J55Mk+yvZNz9eHWHgGzCwy0rN/XYn/OtI8
iQzi5GTwbPE+Jk5W0FsgLHLTvUDBF58iD9xvczwEFDoWXNtjOlrIBjUdly11BGrV
UVelxOfXNL8H2jntk+agGbAsJUhU0hFnyU2Doc6dJj2H7rExXlVrPlCHHqDMZc4W
SlIVgEA2KwnZZi3sVGcEujU9QBIgVYF1k7m9T4ARgAg0qYKbHn4x7JFCdNaLmBv6
oMPNe45jPHHhSAhEPzkhMDauc5mE9jbWWEQyBwhlF4uWvPkUrzadPUAf8EKbGVpa
0Y2R03QgW9JG0luFNaCdMq4FCySBvH2JKcQ2IiC1Pz2d9nLymg69uC6KoP0duKdt
2vwcHu4Od5b+N3qXR387hJQV+bBp2zQHaRjIAP9TxjvLjTqvc1rDwEFUeQVQ1rOn
JcOh1Dd4orfNNR5wZOUkfLh/IG/ZWrmISzaAiD5MYrDwP8IUk3QgC3C+16PLbE7O
8JfyGWCZYu0I2sS4e3ga3yy01dD3zm0jeXt0jGwMBX65b7sW9kBBlnn3nPoatQiu
dQt0520QLbFI1twYA2BvU18Gqf225Da/fs4wWIQuZjZt72bWHPwZpw/D2cJi6+g+
4N9sGjbMPw8ubVdupYdf4WI1AdpbU38Or7j1bNKsbknNtR0NTtDnAfx9DbSMBrvf
OnQ75F3eK0kJhMdkuJL/hB8HtvGnZCo/T5YXK0hqHGbimXRy/wnSPcBtK/JPxAmZ
TOx+atEy5OqO4CHIuchB3BQcJ7VApMWQ6wGsEmLitid87g6/zyM6+vu07sRK9+Sh
vQWvyUWh3sWHa/pkKJhjDRWyP3sXc5jkftf7wnumZOAuJvSDfikhvCRSkeA5Hj4Q
75tskprvR7IcpSjERGKozaBhOIMPmUvFnsTt1Z48nly9lBd3FXRH+6iUhDifPSv+
Mr2rMG6S3LK+JFK24XcAgEUVNXTN9wRWnWqxUKGZFk3LtXOapvu0WKawpxHNutPH
DcylDePHVQquQaHd0iEFRvMcG7hhv1iKOI5jGmUWMXVmfDLevd6UxegZlpYDQPdY
pVCvCjuHWU4w1nqnq2JE66Mp21N1qEP5AYyAVxt9W6b02j2TcVPzOB4lEPuFi7QS
OKesuo0uXQBUb3PonBCKdiOwKkiI7Zzn4x/nqF9aSAmd8b1OKUiYb+UTPvkL7md8
SGup2j23OYcpFuRximIIqU9SssXQmKpZLN84mgmeg9oXB0Umil6XX6PHVnJ4FQys
k9PUX12EVSDQ4btKgq2b2JjZC63qCO/PoDM3Q9gBXG4FcM23QslArY+Ni4HEZ04R
7fkhX+P+aQmj1fvsrvwq4Gwe3y0KWCLUIsPtjerE775BjrdZ7XxmP2ythqp51oVV
/9+jl0eLxxk0zinRjJHOduAFu6lXxByzdy7mbvgoKwPVhKXfgVdXps03S9TcE5UF
JUkziFOxC/TnpOHjvMc94JjgfAQnqaVvsr1N2hORuvtiMHoOV3FOfyujKmqo3awM
lGrEYqwnX7gDdbcI37n/Wp6x5n4bcQbbSCrvCOn/5Onc9NbSXzDK7ICjtB0Mqr2k
xY2QMacQfRN5HFBivtj0TFhsxFelwdszoA2RZZyrl15TsoJ5ub3VIS5iZY++hkKi
dKRjuETHLmuO3mm5eKpiYqF6jnmyMlH3QmX02tyrTvGKC4qcxqxNobEtKMsXM/0T
OhTG15gLHpPCzfptEuuodRW4CnZBjuYVrwa22q/a5C/g/YrO+c0zxJTUIQYkaACM
xCBUAtN0OS9lz5LwWPsyTEtHM7TtpHcx6tNo+C1U75SgNUsz6Bi9KgXgwls5dYIL
kA+AwQbTKvPbHthEfxCC3gzPZu3v4AstGd342bqR0aIMq1Xri9JkCuKwYUvxKwNg
Hs0bVYt689ZB5ZdiZ3d4yJPDFJ1+aC3FhLDE9eUyciWu+B9kvANp088PAr0qJLsL
wEtwU6tZQMLJtgAKwEtu4UtR4GqLFONqGsToIbE9fvbxiOkesM7M6FnjaX0cpytO
QSYb3/+Iu0vbTNCPWBRUCoYEYTwg8NbAjtDnN2KWZ5x1XZ0pJ2obMnllXHBw6RFb
1oMM6UMbt7B0tfw77yE3PH5EuBb15dsKcp/o7rE9ykc0rllqPLZ2kfw6YeZ9yyry
QEDQKYQdLilN3500ReU37+8kFKWx51F1+5sXSpGp874okbuYNNYX7ONzqhOoElMe
OYkQ5IJX5+bUsH4aT4lAP5EKoDaWokAkUImP3zWEKmVuodE3+lMxOsQkZpKePcg6
y0uV+PMMyY/phQ4Y1EDpFrApbNfbIw1mZyYgsSdoIX4GbdaB8mLK450HxnCSpc7p
Y5rd/BSTUOSJ7lclGdq9HjkbUkRfvwi+Y7g9mvIeA32CwAjoP1uEku/iZL1FTvzT
ISm1BabGWeHskGMC7qfMBvH87y++/qMx+QoP7zdJvNdZmOyDHz6rwQy1w6YOaCjT
E89f1UydDS16RC+8SGeqvZhV5Ut3BPP8ShlesnN5gaWmahEpzhx70qJHyq+1+NVF
eYTXPpz6wzsA6H1gXCUFf6mXw8tIxARsX9AxTOqJze/CJ6Y6Vs0IzVB4WmeBAqoX
1YudIucSB2iAeBr+8EFDpVzNrbEmHqjYV+l7AgSEBfGG9oq1dww82EHEfhwtG2tZ
Y0tblW11mlxxhlAE7RI8P5ejW0gfYBix6kc72hrNIL88G3KCNhqMSnHWekiLxh52
AVNMQADcEhO+cOMO417kAJ60enPaYWwawbl9QotbisMes+DNQfuhJ4J22QsC+igv
LXCeDS5rdgFAQMOLwRctrbg49JQCFLKJYA+8krK2t3h3bVhMaeWKkoOmf7U/fzRs
eLUA/lmn/PK2+89wpUXePfty6AUIVJz5RIuBiR/qFasl9Z2xcpGAYiUOiBkikXX+
4kLd8mGmVR20VxB8LM5YRYtszoHFJ0lYWK41HB3G1SKZ+t+NTH8ROigOLuN2g8FN
EIE5Ttpj+QGcgGCLjhImoxHCOAXnbHx6ineKi+64LEVOgOlZot5TSB+5lft7mt+V
Pw4XFZV8loakTdkoZ6a4iqgCaYlGPFrMF1u+U7S/Ig6UoCYx1RICXPUAXlEISLJS
aXSea2R89pVIvy7HfiZIHHnLbt233nCkhmWJ/f8fD5UJg0jJhMPx33muBA7dfoLD
ox9x5kXLvWY7ayA2FyckiIalLNGj396AFQHHf18DD4ivwrzmR8sU/ClSrS0k71GR
VRyTsXEANikvoKmrYOLKqEvBUMHxiExsMUU2J7C4Znb/oLM64iEhLyyVXbJhBgHy
06k+S+4Hx7Preiv4BMk9DTDVCRivKMRzU+Bn84WkwmlaXRueZGQJTBQxVm/oF0L0
5lXVxpjucGPI7WRtlx2PQAqNLN4uFyiKK2Q3tPsjxQWNYLKQzggEkFBZRVXYI0pX
v87HGgLA6xQu6gPGvpzhZ+k/lBQzA3dA+RPqtfH17oO679f7u/Le7gD4N6UU8uSe
62Q/+2p5KM4KFjKgFFfpZUNhN9FkSJLE5m+1qehRYBuwreoDmxSa3upCifNjC4Pp
MG0LdicbpxuJAgRqh6gnMuR2lgYfMxX+5bAw1hk5ODSRFNEtNoGBQlq6Z/FkV62r
wouDhdcPswLkvZUqXiZqGkQQNh/ui5ZHbO/88DJ4jWs8e9zdmA+pruOuZFiEC7AT
OTy2Sn2EWZxGURqrCp9SDFbzg/pQnCJ9/aT5O3HbewJ+ysRRc774ShpvVf4yt/pQ
lQaBj1PDOfy/8zrrq9UWALQvA/uvzs6QzkTENdL0a8sRqsMX3mbNVV/0M5OAMROq
uVWTXkmeFePPyevBueZB5b4qbKHAk3kUFXN8Nm5+/0SQZMT4u/FjRixAMf6/SV/V
KB0k4xm0rywwSdHfmOdnPdJJEmP8BYpxV4myamr+4Dm7g/xuza6B2T8fm8PGuqir
+l1CReO0z2jjHT700N6R1VUX3sag+neJcj1Aq9FkEld78nMo7bqxpGKO3LQCFPcp
qKH7nEMAt9RgDhInMZ+R56g8Tj4TXOpuPvkpgK/Mmgs3aFK9FmB5w0oIBmmfGNAy
4HD6DqDOOg/lTHhc4sZMFAChcdBWiuakzFzzh3tC6Xf1nYL9HVSPAEbg7AZbW247
qewI0zPhW4v7rzZoluROOeU245SPYrG1xImyQs72XDD1WOtXYN2zFLB3jJKuDidG
1JqXwAFYRYPQKlZnr3aJddn59NY+fZF4XxAl3xqGjXF4y9fTbvMgfRo8eY5Y/H0M
03aEfJ7m4qWRUTa7wrzrXYT6MR674reIYvWL6QDGl77e7JFS9dHG3rvrbWKJOXjS
bhVntpGdvq65/G21ahaW7oPmCZm8N967vfMesm/Z98ulnT9yDy/0JUmoGgbdI014
GfaHdhdY27kFYcXJt5ruJmROQexr1fIAwpAYAnEEpAeJCt+b4jTslAe3FPAdhRYK
4InQ/7L6+TiOhMxJ1ikVday7FmzTjcCTofm3O6PgBwIUlKkDfIAYGS7VebZD25cQ
1WosOtf85ddWmx3TTRfHQVxBVWcI1MxnvByXCC9bARAZ7P70RMqYzO/GsZ6H9Qzz
r6gUs/syREF+mPzb5SBOu4jyiAgSyUqB8qEhieAp7r7mLmFUFQHRrAt9koErOMnJ
7GfGdb3D7GZgwyN0NxgZdTcW3F551ZVYIbMZ7WCM7gcYtgfrMwpVqsrrWGGrl5q+
x4xjV64QvTrK+6U4n2xQ8LR2RVJDq2KHK0LP8JpaSeL9jHhLvFkXtZgjC27xKTMd
eBn0CNbUZTujTsUcfa8NvF+Oyl8v5Jt6MpOBGl4M+bXX6m2eMaAbjSSU9noZiTMx
8QXoRD1kHntjylnqESEaVtroZICuHMZNly+WQixKJX7LGUJlevgfBnGmmWsXR+iI
BoV+aY7KGfUyr9vJFOAjhyTmI872PX+P2Sd8XPuvhiFq3frPOOQ7/h4vAOJ499I8
pcH1KmmkUam61TYTpV1ckRu07l6q8gujA6dq/XG70rbrXjoW6MxgEtBV7BXI6d5+
1k7xUFKlXDnuOF55xoufX1xl73dta/OrdURibhxEUb9cJUeIGqO2xCzZ/WJbFjiw
BTPpTab2nOWBKe/AsqKEbNU7+UD9B+XWWL7tfpy6SANx2gg7gaew0k8U6rNfxn9U
JqJSkCRQI0ZT/iUAw3ZGHoPnUDCj8sMl4EC0thZxlW4PH2A3A5UWPbb85DlE8asY
EyPqmE8rvvMURXqwNoGHEu74WqWJ1W2K/oUXHK1qziWFLFV/ZIpdF11BmAjy4b/N
7AwhxhoI9RUrK7gofZal5hFO+c3sHTD8EnbWZLSmXlufwIm1BN8qOnsI4iZVuMc2
GBTF3yhVkWq3XLeX7pGCQRQ8LBTrfJRptYXlhQGwJjZx+4WVO5AhO6SoroEHR64A
JFhr47VaM/wRZBIywNCbbPu92im5p5JCGrJ3AD+GpnEQxCwoe2SWp5he8DftkkEG
R6LUz2mvV8NLzOBRzBR56EJwjigEfyt3KbRe23rZyzBrIGcPjhODgK3YQi+MHBSx
g77a7TQcUuIJzOm9DBXOFglHfSJivoyxq4TQeow31LPNZNCcq5HBp0/tXDa6CoYb
Ex+w6zM/T8WZvt/+Xp9Ydv9psBHB9Iqhh/qOWXWg9bQmdN2Xq9rX2RgMwKGRSWJd
vT6r7YvKY/xQV2YeODsapIJYkv7dIdBQvUcoiTGLhckipB97Y4L6rZtf5sRjQc+R
vDbbKuHd9cUDUj3GZvJbgEMFPsqEi6ahAZsVjc/+NpI+93ujm8e1S047g8YLH+KY
mSAZipP9+WkIW4Yzff+kLXhrDWPENv2oph/stB+kOU1ObXcd5/SngCAH0rXzqgfT
tcY244CdFdP5vxuHEh+4BEIzAXrPJ4+4j3oNP+Noqcrnw9nnszpJdt3P0XIFVykZ
ov7Yz6J4pjGYqpzFRZC/zFmt6dJ7YUNJHdLW7nmlLKPUeRvKmrl6pEiteKrKV8SL
cUFS34lTocZpArrdOEjmovZ34dKQjZ7YQsfHe2JeFsnWeKH7p71W6ZlxiYZZZSIS
btzuL/AR471Ib3JhNZjBRjuUcFjiMOvBeRsG9K3fJQPJnKabTiNRxyDif+CqFEXW
vzwFoxh76uaXYfN4WFL2HojT9Mf3s+9hJF4UyIwUIAxZ+V1Uz2OraPLSSbiPM7Tq
RupDcqCm2TDUBaXjFix5aA4tpM2fc6xisfnc4ojiRu3wb+4VEanZOllwTiJgyzDr
QMabev+UgrdexyMd43D85T+Jnl6O9VvoF8y5XP75o9k6SiFvmUs9MT8rBE91vA2e
v+A8UaXozzCu0V4mGK2f34H8U54O48Mwk93dtYxGIln89a8VNB/KrPjUDvLZXK+9
zUij/bpXjth85FuaGYIoTc2TJH+ZF/qUFkAqJxRwdqcuBdT73LiEnQo0om314AxZ
BKASM9y0Qv/IaizamV3nWLK0J4HseTvXVndP8T9p8qRjDdfKOJ2WqzMypaFIs4tN
Pyi9X+/axTJxOFKKKgqt9EDOue4kLim8S5QiOYAf/kyK4ev927BUQ6arm0I8HiL9
YDNmie5ASTTTdkjXeEuVVMfNnC8+s1gPUOr7MceLIOODTwzjXN57XfBCV8NRb2rl
/5CnHqXX+LAiFdw7csZYP7FirfpDnHP7yUHhQ+TxoJleiSb3o7wx1SVjV8Pl5FDm
AdRy1ow5TOn3Xv85N6Z18D8qzInljCAnZMTpXR4UL/MPovJTAwniXt8XmJV+rbD9
wy2LEw67J9u636zAeszSNABEK4PDoVqmjCVjxSK4CNsCl7hhV1ZaYZ//oHyP9Fp+
+azH0XyXznW+4+EH1T35bIMMVLiSGGuQGLZBCBaTA0l7dctArpdBBLXK25nOqT2H
8Mi69hNF/GBCz089Tei9+wI+qRoPRixBLXrSLCSWrLtmRzsC+kUicuWfaW0Ef9hl
n85Mjlk92bgVmr03jEGmQ5KiYpxl9+Zfg0rRkmwuBXrkXjMzi1219Z51Pantn0CR
pz0hiDuYY39PU8jEEsiD2SHI+d54Wte280BVnInY7qqvyMCQ928q6L02G/54otjb
DG8jbNSg7q4/hGbLaaeZBa/fEdsZoGiHorzH48okFnu/M96cQzwuUeNaw8IKD5JL
xzdz/HbJ7nA0WTUdbCBBgyq5WNs2rzwgwzU8kdICI7nJVX1KaalvY9yllKhFzagD
2ZN5tz9xoNFg2Kdz5IZg7vT8wxzMrAUb36S70vRBIV7uX/zbjSJoUPZm1YmTUf5G
wkTVTIhX7MmaWpwkvPPBMtE99so1d1l5FZXJEqwwua3ordr6S1r+I3LglYVWCfMI
S2PNrbw0cm3hETW8Nw8ZOSEx/6mL+5MyUB+SSw3H9TZiZf/LOpkTcJgV7hZwmwOT
UOO3zTMehJPb0+KhNIEJvECeFs0Ks8VR8sWKF0xh/MxHyM+PqoI8ska1bjHdvvkR
OJaeHnFOIlk44WRnRXw+nTC6/JeeXPBcdZ6yoloMw28uuRy/SA9x+3F2C315HsxA
9f573hXX/fa6810PJXHk4ccpy3hPCkQLT7adtrmXOtw/WJKQgKWMnhVAGHBSvGyd
0sHxG68cixAjnrjCoO1enVYpXuTqTgd9EIh3d4Od6Y4LkEy85elUHkzjbG/VvfHp
+o88G6cfwvE5FEFG1/sNyhx5yXEgfV9WKKb6L08siUZw8LGIUwHzYREMM0IwZDA7
wzmiK8gQAciduGDBk7ZWfWAXKidxhpFT4heqrPO/OUah+UsV2yfmAfMM4Ab1I2Hw
urk3pVaQo/hTFiEUnWk7UDs978ou14qaUnZr7iq1aq1vdjy3V6FsGKp6GyJYmkoL
n8bhj2k+VGpa0TrXUkPY5/vlRrCAuqs8ogwbMVEVNl9mD856C+6P+jTWFNg3d2+p
AN/KMtFQBTTi0u3jrloEoR4+YCI+dYWuU9GLZ/Gal7jBJCrv1RqUqS2bD6Ad1kc/
QimIR+iYQgAr+O0CCeq14AzRiaNvj/Tab493zRUWCW665GAYFrfR6mRJHSRzuwpU
36C2zdj7adVYSN/VUUrtcr/IwxTIdms+9VpU6LpTeD6Cq8RYqu4vOWGFW0C0xwRH
l3M5z2P7y48XjMg2ENYJZM0ecn2C9w90sIayiHGGlrHNlsQ8fW2zACzE1zLOSoro
PEzaUcQ85n34bCUKAkxSPgkrmGmeYBpR8Ye/t9X72ey0e7tU+XeocFxDXX41s7LX
x0uqa/5FQoCoz726FzN7jC//au4QrT7tOe4pg4ZrQgO4UgZq3Fys5Cj7cT93Zibi
fVJHIklUW2x7l2axucYkiuYXOpiRAEKj8RagYAsnOUEtnu9uivibWltwcl6P/v6U
/+KP5dyTbCOyzBocLl2VKUVUARXFJj4ZPm0kGa3Pg/ZTSm939CduRl/VuFhSFJ0p
4E05gRxWEddxzqb92VlaDYNIsWydMM29w+RC2TfOjAdB09UqpuawsVICRdPBAZzp
SUJnPtbOZLxHOh3/hNqYLrG1sD2G6hVjw5C13jOmK55ClgHC/SLyN+vES+Hl8o05
szuWMJBa6BDF6jddObOMqDKxdnCeK7ntQW59gi0OXzdZ1dD88xlhPI5gg2gIaNnn
DeUmvZnPwpdRDTUpwUJOXLvhz4d8uN3yHrzgj5oQWzIrIH6lOqO5pG9CWpJhITQQ
fzSb5GghzzBL2iQIvztX+HIXZ2/4b8pc7G1HbMRSrPsVe36mlFUdlA2Qc2kxG00e
FcoVPBDk68PW5CJJBMDfswA98f38dOeGiOabMtRFJr5Q9xeEb+ERjKKuL1ZpXH7M
J9ogskaFVKaP6mUE1eCMbwm+jPK5+WAq8xWsRpQ/dXCB2FhpPNHQtRU49PBX9NSN
mbN56Kaan9cYa7qtatL3EcxszRQNLrIOW7RkNM8Q1FI2iaDgt9Y8X+dUJpG/Zp1Y
ttvYD7rl2C9b7Je0G6BaAFqCpcKdMpd2Vg2P3jZMH7jONGo/1mFTsL87opGj5B5x
kO1GSjOYWI7Hy9/45mQwBDb99wg7mAqM+tWehIbv2ILXm3xgamPBoW1luA89/z2N
upwLzkRJLeBxoI8RjqrUaHpGfNZ96OciIPvgbGP+VBSlQKdTVMH6u2Jd7i3MwykB
Z9sh35Nk9W90Ii8mtE8PEhLkwc/8rHFCsQ5J1rFG/hNKLfblPQTSkVw+90CFgleC
hHUEe2kMqrTvCpoWFcnn/Jo6nC70NQm4CURAuVNuaR6iBlPhX82dm1PSPxRfW4f7
8AgNLqk5Odsj+fI5Ipu1KV6GRYWfAjX36aVs515Gp2a20049UTSqeIlYE19yYmN/
5ZsI/XzRe5e4Wt++RYd+7fGc99ZXHK/LIFf1ZlxuCnt9qYa4f7c4ZGYOvkRkbURX
kkuKhRcoSQGO1m9Q5lp62EOmbwXLEwoNi1S6fJyQUQOHeAwUVfI99ozr3I9X/JXR
w4RNIiI9UC5F8pEhKmKCAwv13nuYPTNIJh1wL0vXZkey96pFriOzG7q8QMVLKVJs
5a8O0kiHEJunCjiJPQD9i5O+9pRrZNfPDp0s/XbFrwqw5OL0MnHk0414RbM3wfdv
SfPcGvd3dK66MTZ3Z1otW2osXajZZxV77yIqnEvMEhJVWyc9N+Oi3XPoTc3Y9++7
OlyPX7sr4cB7S1YIZFq51VChNU2c8fBmblG4/zpLYUo8u+vMwQL6r12aJGcUnd8P
Eet6ZZD7JSEoAO/XSdd6X60sm5ntUC4amIh89uuRhwmEAO9TWUXsjtb5+z5SPZmP
MlzuVtB9FHHaGpUz4D3b3nvt/cd+PGhOf5PsVZJJ8KOY9Rxt/FrdHgtdXX093h65
/BZhLc9AlkrgdWTPoyRS+SN1MQWD8eNHubtVVwqoy1ax4ImEtvQ0mK7V8B8PePAh
58+Mb7jleapvsa0m+acSG5e8uKHJXMi+pJM6It2WWc6sTINhZ4ol4u7t4qtivIls
AoJrV6ilhokaHztL9UPIc4VVKqAQTEHMB7juTHEuyTDJ2FI0QYXNBZGiqJOe+EWJ
IMsrXYbIPlOhkgxOUQMrJSSJPAfM3jxCifI7iqdmKGpDmtUSqaTqetHqojef71G8
PlpvlvSqXFbr785JG/4/4uWwS/NRxmIOC2cKzMD8eADqduVaKxPZu9XRG9V1o/g1
kjsouai0rclKoA1crQHOZBlrW3T6J/0ccXRiidELpFZmDzWBxEYw/Cv5Ol4rwB3P
Fz0LScGrBoOE3pSVhMj1Pia7+iV8e+sFsHR6bCod3MMMycG/S14j4zENOu5vMEu0
4NkMPyv42pI3Bjj5o5Nn2MK+/HsLqjNtWGo7tcW8y25iM3UB7gB6riqpLTI6vYPL
KnV7mLdU+o2aXqqKJoE9nc7RAAkUkijopNp3qGXU0V1kAXLMkkHyOUVcxYkHi/hS
/+o1A2PZZHjDnG/L45v70uH0sMbQ3qZfQ+6UqwZH5cuxDd3725W7iz2/FO5hHxdl
cdVmQ0YEUfVPcS43zkosxsamKDtO0HLzazY0I/qrv4XijuS2atj7om7nLRCiNLCG
Qk5ed+fKNYZDDVhXVtNHpvahDvtuNLHlm6TPAt94Ylyq/Cg6OE2J6PW5wtUUv93I
0o8nU0ZjPC3AVns2by+8q8DxlTafldYVsVSwIbFpLv2Pqx95dXYiwCg6GEhIUenS
67V/8fqhkAp/cjW5UMM7yjpBg62jdsp++O+Ipyblg5dfGXaq3pi2EdJWaxDzTrBP
8j933vRV6S+AATKFjXu5hLFC5zdiTU0tetETNyVWwBMtoYfnf2SIRzv0yIxuBZpd
Vfpkh77uzjy2uY63RUpKphuW9UQwDFCkrnClRYQyYIhYhcbQEsj9ahh0Ck11DJLx
DS5aJZTf8EGqcuYEQejbR9V2xLyZi5fyEPWARw1VRYDXO+Gcf/W8i78cSJYA+4wn
XpuCX+E316jYTO3kMmq7+1h4nWrhaUQYY7juR0UUzA3nJU21lDFtB+ATuYUlopw1
CKPF1Q0YAdsNqyQw7wiSwgdzCmF6xG4+Ie6P2MZr98cEDb+HuB9fqPFWfdJCbpBK
KdJ4CHRdY3NykmyEqGN5aDbJE9XgD8pZ8oJ18Z4DqXooC5KacT2Z2ulF/Eak4wpy
peuNNXQO09e8zc7JK9sboL+CCJptpEK9gXZm1JHRCm7zp8vq4hXpsyFLdm5dIjVQ
zTjOkjJfhwOIHAj0d1yK3ERdFfxtpFC9d/yiq7afnPib5KtvpX1g9F9aGWHUzY8X
v0N5yN6aLXftimH12WkdpBrcl1OBZbYdT0Mk10u9EeiHXXoDFBJTm4oGQLbegsC3
jNe+cuRJ02QQxz6TbqqA3a8COntcfw+V9rmONaMqUmqd8ERFYAPsRfNDFx+TiXo+
0Xb7g4ggDR9/+CkgUS4XxBbYGIIcTJW5IGfg6vtnfJnvgNW8+bnqucIjITtPDff5
rZDlnR1bUZMnqmqGmjnJnA97b4FKAbRYTG0wYMK6o+MgY3hp0Tf6J5ubtiwEuub/
BN2rpUZvyhPYA2E2WI8IYA9l7AdRgfkpE0E4NQVYfbCHp4vRNQKpCOwf+ypmz3V2
1buR8DJhVmx3YtKikw0jng==
`protect END_PROTECTED
