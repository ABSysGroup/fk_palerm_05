`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zZ4mnQUnnAUv+UDG2VlE1rTuQDWuDd/N2t7zpFgaHAG90b06azs92LQlntswACyT
odJJf2Fx2Vwui6snF9yO6DRWa7dgueUZ8DyliTwrZB5CDhAzZ9f0Rhulk/MAIOhW
xOTei+XMUquYabD9eTnGQGJD05Gb5T0zSwUOxVGiOI65IEMEXk7eFLBbz6k22tl9
aH6qaiF1zR5mxJ0ckzJ5Fv7yuwbEB9uoD+hTJrwPVEUGuWC86FtUNhYv6tBtUDBs
aa1vhkBFAyo2YG/9awtCnfkfgQQRCVGmnvwujocVTtx876J27z+LFtww7WLVCZfU
4BozzT9RfmnxtEMEuRDpF/R/fMHumKQZAEwHYHEkXjITvOD40XrjjpK2XzW64pfH
eH5FY1Puu3XGlX8NsnhVYVNgQgnfHser76j+TWZMKwHRHzWvj6F+ddrGy1KYCGNC
ztkPnVHjXmmOboerwdEBLjHJCX0kEJ4sfEJRkXwVBwPgPDGWEi4Aoxi9sYdWXPCf
mS33jwyi6lJhUkThrdLADwG3iLKzeOIzmxD6+DjxtAFOH2DgHIG7Au1u4FqngMS6
yfRdT/Ho6FMvqjtxvkFV0VlUZyXcICyDY8uLrng+sJbCwuvKsyMW9NXAuyyXh/x4
SHsrFamJ1FhAsrRZeSlKv22Z37fC8qZQ0J8MMYmigJY=
`protect END_PROTECTED
