`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dHAX6NR8LfgedPB7nFXKEEmcOVFaCEI94OLodCWLypOVZCYo3NV2dJtOe86XgBiD
djWN7XbfEoZMctOhuY5yWSZ35kXCOl03mYfnhQHBED5jBlhAuL1Gl0ujzwXQSBHl
IvaY/4F9Fz/jUZgvZnUpLpjHm4U8zffBtiVVb/oj8Bu1HT6A8SONoMWf/UDBdEyV
rYZVNbo9UyRLuDebGJBI7ZNyP4GAXbwDjHa//sWxOc0Ih55bctEi9r+EAPhtxm85
nE2ArZBSQexPNbW7Skk16+6Ai5Yp2jOPxCtXl0PyEvnP9E4Y1vskKRe98HYEexAV
o1AZ1c6SlmNsncdIXAQcWgGVmx/FYdNWeuqJiRyIP8bOnUJeU0dTzbfVfovUZlSQ
cGLjnvcZODLJTiD6kVdfapYJl1p8NE5XvI8ZWowdlpFWzPSOjB1p9BB0Lpm4/gUa
lOQaUtmUC038gpdECEootw==
`protect END_PROTECTED
