`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VJY6wdsLLHvxcvFSPP6xlfsmJdDxaV0w1CT8KHVbPyz9lSTCDON40RW4J0676Zck
WxMKCo1MQqSQhEwMkwn/m4j0kHBpPkSHDA0Ew6V+w5z6I49qinmRxggiQSzmSq2d
Eo8zNduo6cG4dLRH5ZtRtq3ieW9Q1M4c8fcjGa7HLY0dlEL/3e0iKUqX6sKuFOZu
dq8ep6udv/vrdmJkSqE7ZHIwlwVEaVDl+ZQJ1bXDp8POZGaDPvj3J4H2GeQbRtYA
hUumpyEBfO57AMqPg105W7k1FnSawsoNhyPRFkEg4WLbHIh9rVgFeVJ9OfP+q1zr
MXtvoHsCj4r0w00i7BnxYkgyYBNTXMSHRQIYIlX9kBjDHHK4Df2juLlPwJ6NfB4Y
fC9GoEv3wDFlLS1CJWYQxP9kl2v6/wP3FW0N2EoMb7vIounAKEdyjpwG7Rk6TPar
bkwrNoXlCp8QzCe+Hm6P089heUHeHigjF4qJmTgNcQ/6HDgxMIyrRi8+0m77crQN
1XUgbqQ4XYyjZbTHI+79LOizuawmiXlmd6ZOG+WxXupvROH3DXQyOMEwmFO1duLu
Ud5Zqrqpxi51qO6EsKDBp7TEneQcQJxC6BcnmavxMBCEo2stkj2OxJ1AXpqJ2KAf
qReaW/knso3p9QNJKEcv5w==
`protect END_PROTECTED
