`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uEsQ62qj4jKhpAdZJmCysuLwnVYU/lDlc0EcEZYP5KJnkgjO0Sz8lEOGGuhptmBv
VYfpFGov8Fz3UpU4jft2kqezjl8cJkpM58u1aa9vwYTPLe7+5gKw0na9p0lxHVow
kxQXwCQNmRMr6RKMnkeMpko+EDq5POloBEvLZpvfMFGsG/m+2ETW5waG1BqxLJEm
4ANQcYaLo+vttq+Xg9xxfVWm0ffb2AFpoAndxs6n4Y5xKdDR60v6BBKcRqkjXkb+
EWbmIidc/4YhaJXZfJYeSgQlWs19IISFWzEG2yfWqjceud0NU5RSh3GefUJShKXn
KS+E6aLiyZqXubDFXs/mZctpkqOeDXcKJozpqrXc26sZRKUxQhutCCR+Nq6zXMIv
lL5sOwqBVNhblTQhDSahU+/u0s+TvouQsNvF0gPYbjalBe2gDyLv0M7npq2oE2VL
dyUr1ma5AchSQuxRis/SRoF3eTQRMtoF5LA5krC0dURgHqXl9dJEj/JecGS21fss
IXzqfW9mQhRQmazo8Uud0467/0GIhUl4dexQ4kLFVPiquKR1JPG+1knnmP26SoDg
7HJtxDgxRSqUvpQJkWnlqG7veuaqtWg9ZjRlsCbZAk6vQ0Q6O4voCUKHW9NlkT6T
ZiDuE2tSxsPybVMeOGxo7QtCRe90s8pmFDUytfA4LIsCF3TK7QBfhgJEy4pJ+75A
2TF2jUt20AC2iJb41QM5WbplbzVMpa9tuJkL11CNTCoBwM4QKK/ao855yMzknGrD
vcNOyHOjtd//G5400TR8EqBmyAbVs1eHc5yRfmtC8y8CIdgCH/jtf64yLlVbVUlu
uqtMUzxZVwXbtItbviT9PBlDrIFeVS7G5+Wczz4qpkO6Fn7iNVE8oWC8KPKu42lZ
cHqUJPGU1z9/QTx3AZr9k6jkhAqymjFzvQeeJR9plBGsD6yA6m3ZyEW06PQYyoEq
AONTxH632eWycXyLugiqsrdq24xA/4ZWlPo/l/AyAXtz3grPWLqHj10GTj1R/XaP
KyNwOK8qi8PhuNNSR2aR2gOpdIYhvlZDm//KkIxWZr8idI8AozCUHQx8qmeM9Uck
LLXI2o12SADaMOx8d3oGXEc6VsVp1wCM2WD5Ii6m9s/4eKTBn/sywSsdCA5KyMlV
X2AcNw+SfWFyKz4gWicja4XeGHAb7j3cFW3UGMS58x7E8YrryoRZ83Df7fCMuDAI
zLWfLlH2zYHn35DBevSz7AZkjLTcqKiWBMOkJS8mmtlFr3aNXR3avuaY0Ky3vM6u
/2MkoEkOvuQdWui2gP7lKzg0TS5aJmvOtQ+2qZ1laM5LsCgf2rl9OWEXagnipJbV
MaAbxq8+gM/Thj2tCMcNMovQeMRI5wEwStykJfo/qzGEZpzIbV7wBrLCU70CWkp0
EuYw/eckMLq3Tdum9WpCRydAFR0YBtleN7mPL8g7XnXsrd9i6p6XLfVR4RdQFI+I
dOW3NGPCVu36Eet4yxy46mG6n/T+LzpxvgUf/BdOFU1K3F0jNoVegXUVchilNAe9
cAEb5Oggitl0G5pXbUkZ0/kvM5RZAXzl975R/OGssdkB+vw6tLGEdGTs5lTRUUA5
USt17McA5KFr4R6pwdGF63k9iWtqFrvxdICd90gVv5bJj10Fehw2w0aG6DlhxIMn
b3axNqv1hGBZQFwl8a2wyx2bZfK42Hbj11tRdsdDeMmYUmYKPY2DWRBvepHFrhAz
YVRRE6X5t6OOtAUoz6+XuL7gOqhnRJkfiEsy9XK1uZy5lq8ubockcJQK63pq1z+K
8c1fEU6xT15ANEA9HoOk1Uy8dX/CN8Bu/7+vzD3LkA16socUjGiVA7JGIx6VLwP1
Xb2VJ140MEQzh83A8WZSXu3JjKe92vU2luAuXAbligy4xsx6gY2gnfOi5P7uZBkV
j7V4+0ppYBaQ1pKQ1xO8AImLvMC8+UpD26zdNEqxFpHQX0CWsnzGz1RiwBqyQk14
XTVNBjhJo+SaX4Pr9+7LfGHRtLfsZMj1oAFjs/4iweLkrU+JK/OQauaHOnydD/7+
pSb72gyBGe4L9QhIXiPnEzUX1NVRVMoAMHZdqzSjKOvgBGuh3DdpF+8i3pod1C96
4FzBybDepAThwwq+7TTcQGbfinf0/1lbO3nTbflhYP6hIl2AlpT7gqhCCzQPz8MK
DcfbdfA8AokZd8EdN9i9B79neVy4Otb5P7deZSjCuXXkhaPBykiL7HtPEWEwgcf+
Y2AuggeDPAl5gpyl7SRKup3S/ZZ7p3JGudkGBykeFTbzIfiyqXNUlWnw5Pn3xA1v
bx4xxeZ/J3E7nMw4R6N1oYCBY/xSXN5rw58WS+mtiXcYgxOXbp7fzi2TMUYcDbRY
fSrOyMR1bGD7KbpvDpGvHIkaXfbyh2YvHoXbOncayVcVRBl003OdYFLS43rM09I6
jK3kOZlMf70aTokQnTx5Y58Iz2tn8X2Oy7BDjMu/4hHQ/4XfXhTMmIre7VcsU1nN
1wenBUv9tBfzuUj6oiCevuk5LmNR3WJNbJZfeApi0Mb2vGQN6OfbBh9r9seeYu8T
t7ygjKAseC63b0ZPIJTIcdj122f4f7LuXjrOPJ17Wcmx9T1lEYUp6ELtPch8fMAO
QfAPlw2/zSteMka3q3AzwmYDUgFZFhE3HPgybGf63y0Gs8ZRiny7Co35Q1VAuzbS
NuhUGEI30TbXOncZAoLP/BEgv1z0aUv446oJOE5mZ9QfOuSSO0vVhoXVhPYeU+Pk
mwM1NQraafl3FVBuHg83tOWGowjP8zFTY1Uoza7f3uaYTh1F+6Hg1bC75sAGOkQg
kKDElZ1bhQWjyhZzwFiymC+lQdeqfjRDBK2ftT+ldmds66ZRJgZNg+/HMoO8E2Ks
1ZrR0DUERz+EsFVoU57n1dtkODZrvzUc03f9UJwmCZfqFwzLB7Lgs/ipMNUwuT9L
JAcYe/kV/QvpUyFbK+hJ0Zjzz2erjEz0syRHE23ubUoyiaN6jJKIxiz9o4XRq2X5
GZDpJtiTYJuWqnuckACxoo4xO58tQyXY3G0mSCw9pJyeunVnypVRC8FH83g8NPMA
ggsXKZk/13vSFg49+epc1Ma++lti4nZgIAjU+M4p/N+mmhMr3lmRzzu4t+o5iK4I
wG/QTDtUyzK1OsvCpMvqPNTjiY0waCUFg1wmPiQpIJweKKGJDme1j1PZD/kVo1jf
8GDEbB6HHGrv3UBauD9rFJx6PtY/gYAIIaFX8SK5Jk/g6EmbL4Y1bxkatzKKvdVJ
jEGe+IIBxcIJIFL9Ei7rW7lgBJ3BTLRnnWyseHEwBPaJk6VaOvj3TP894e752m39
kbd++BJlqdaDX4OBUtUuVa2Zbg19+h07SDEH/PPBH0paeCpzkTVnt/DE+gNx/eSR
KONVY6OXNEK3YGNX6DRRkpuBVc8fHyoejTIMJgZNkKXsHNYmuArr9eiv1V+7JzhT
974B6a54yLStP11iiVas3HZ28xyrx5RiRVounxa2yijair+UGAFuteFpwkMcYg1m
0tWaqyqA/VMTadZJSfWY3LpnJe8Df+bLxoLDfFczs5KT6bXJXolsWS3L9CxJ+3DQ
A4lwUxwYUsvyrqcyjmGwoElRk3aVTiZOjn9zrQT6FC8F45Be3hj4xu4+5L5L0C0w
lgi+zvMiQSIAYz9YRmfkveWDgOEdO9I1PQSPNTjbdvf207O4Nv77SN4hFgcyIFXw
sJCv5Vi268mNgQ4WM9sUGBLj0pbGirxm5ZLF8OB/VSXgNkH6Q894wNDpwIe/cKXl
RTVLaXYXvx1oYTMdoUZIOxURGTpb8yTQ+j5iKMidkekZTLT9EvGIGqid2mitYHJQ
Tyn35MAPy+2XzB849g3oPTjqTGQgFPrTOrdXRhp7o+o8JtJhlaVcUXShI6AAWvxg
/Ih2P6SIV2dbMrjLQwVDYi3qcx+g6f43iB3ZsvxiMZMAYbMYSP9iqSCKtpW/93ha
DMs8K+13Y57R1y/gN4r/f9mclLN7TsCQO6BZ4aIpdXfe9c39wcULFRP5F6SvsjXU
PQ0nuOcfbEzALFBuKAfYZH1UiSC0T3fIL2MnfGrgDsO9vnkb3J2BUnNTKOKis73Z
31c2Tm5vSulFgNC85iwkwsNpbhYhYAgwOqx15/tHoOuOhsthp0kXzRPR0XUuhiQf
tUVnKuEtTt6lAOCirKnjNgQttVQsEmmEd4LHR8a3/ufsvK32DBoATvJzmMtkS6o+
VfxbZaSlQ+EbC/O7ZzVJAXjs/mBFbSqEuERp467M0R9cPwPDoiJ4hzk+w3KQQdv7
1KgGywfwENo7+eoLTClOAq+7rI7zSXGuHgGjVPkBDzL2BYCkGwVkwXjsPFRkOu7w
wjOALRZgYnJn6thiFBbiLRInJcz2qMafC9pPXStIgtNcuGR4gVFIN/qVNChO1UEP
9wv/O4XyN3UMTAl7tvlo1u1qRPRvvdFE61R8JzC6jkfJVyMzewEmyuB0Ir1o5SV5
E6MfzccVN3uGV8tCLyR7/Ibka1nZlXYKO8+P55mJTUi82PDtti2TQtNk5nm7g2yJ
OQGTde3ljA+sJp3LvDnV1utdzFkK5APAHxXi/pXUC1Lf1+RYAlfvmv2FLqzXVEMD
vQ9PIvRud1r72QGr6DI6hrZ7EDaXF9WBEAq24srzHr5/BTFQPu4Z376ja6M3c2vt
yZFM8JqKgiaz6Xw9n1fL8wrOrQOjsvPrQ14bDyLJIlSBj/oGwx5hDEpbaiASMOqc
CGUBukSw11w0zwfq85y0MNhlpTSYveUu1GOVX16WqGvfl+2+M793Ky9RwXtjoo6k
ilmWX3633okwiQoROxs3omhuwhkRvi3OwD0Ak2YocykUcVI0ClEICTThSsI8tS6F
jd7A6D+ArvDKlT++RycmauUIFYV9oHq64chF6WGE2d8GofkyY226MvjfAmMQwTDR
2+EqpbpqIVhqYbUpwSTYxBeTlYoy2f/rcBlCipJim25e4GRGJU8wGOZ3izgnVw3B
4XRpxfjgu5YNO2LtUdrb8cdvoW+bJhuLWgWg3HqxjZfu12A8IDliRXWZgGNj4VOX
OIFpcaGzdOPm8g/Ux8P1AUHzdArizwW5dS9gAjUT5PMncoSjavKwqTIoGU2aFfwB
r86YSuhymRQFNqGO1o6HzwgEk3MOnrslbN8ABdB9KXC4lj/oIkp3tE6GJQUM5KRv
o3UdNLLXOrvBlCUF0td4Qw4XM8W1j6gmqYQLoKLctjf//LnlWWTKdT6Z/oI0G4UP
mnzpRKe07i2vcYGmWDYpRV3Lj4X3JPxBGjcDnnnYtMY6UR3uWvrl9wqzGhc/veUm
mpxkJKxnR6Y4LY37wAh9SyWZ9qYVwtWq8t8BNGZv3tAQdGiuzNt9VIK5EB8DE0wX
qPbWsmT1jcqcYHTlqb1kLyfSKMh2IZDue8K9SOL6BqZNl8QsaKPUn/vL8xUE+Qo+
wN45LcE0QSYMbJnDd96XTclsLNyi+0obvpk+PsXOY77F3Qb8UXiPKunVSagyebKi
3e+pCBzZkTsfYpA4nDSBdlTsYqCNaU4c9tdlcF1uNmWYR5E4m2/3BUO+Kw0tgC1x
gKtR/orCCrenvDZIjIAQ84kuSfOrAUBs0HEcIM9AFqWby1se6uWxwSeGRkJPl70M
FVAMfv9RGFLqPr6s3TstYWh9NefUA6EEDag9f85kzFEUNMg4jT1fpoF8YmgFGtBA
mPCK35Ooy4InoFNZFVavVH0QEuHfJgfr93y8Q8Ie0b5XviuaekuZkl10wlM64rzL
MvoFOLt5hbbTuhOJCaS0VIMArid5geTqrM4Z48pfznUdTKDqiAUdJzPvwm5SHKBd
R7nyyrj93nBEKDJmZB4ZVY8/WI69T3Rw0IYy+D7XE2ZQeehlCf4BFaawsksEeXXP
J5mYpkNO/d8RjuMqiGbOMumHhDl+z/BL2vbz/a2L+qsErHkUSDyZvLEABnK8Bajq
lPYQnuwz2HmV/VLbZu4CcXfj+xMUyssHIIifYj2aBcH0pbRqa8I3JKIy2EkF+RZv
/r527evbfcBFLMPal1IeqgTzsX8DBiDtcpot3RS2uJYUF9DLJAvdERGCmi7DeaAx
emqYvyjCXtdpmN59MnAeCNtSnSWrGzzHEACt8bUVugokzJ3t2aQ9hpfrcgJgeC7W
fXoeT0XOxOB6l9hEfhC90BdUaqJ5TPCAXAM0GYaMssdc1aDEphTETvm661KDsgBz
6G7Vpwv0mJpslVfMv80iEQCM1T++xer6rmA4yPjgmEBZDnR5iJwOCuX2TYxPYa4a
NeChiSKIaeqEpHn+QfnuddlesYdsZ9u/8Jcko/0qncpJvQWjf6YU4L5CE4RpciSl
Qft5m9Nc+GMqGeOil0jak6AP+qbj+IDL9rispLSxWRSFOCwkc9f6y+GCvEWsW5oP
cfPmHk++sdq8XnATlpIj2ZTQSXDZFVTFpl2zWYPLnimyySFJWeC57f3Nw7F7i5kg
RszlE9Ouspd9kJXuBohzVR4+DDiFI3QY2TKOFH8gZLGEfBHas+LVwVQYGwF60eYH
HJ7EyqNh/JSirg1gIq7wUxGlZJQJwI+S+CS7qz41MzKpILU8U1wakvCXIcw+a/mJ
bkXQ25r5gc/WJcSvl8OpP4SvDf6b+WH6MwdFd5bdYsZG8nnzizRAwJzKbpHW7uaD
itgnYQQy+qA86nYIt/tyFsRNevF2LS1CTpIIe8+Bs8382MtEFX/yRn3Fy6YyT9C2
NxqcdfyMJz/kKnrvxfNHhzn7uD4gR3Q5m/FHSl+76xLrrWgXR7BNrY4YyP6g+Zzs
CcnqP05Odl6dGmnvkyhf7BCXrrzlOZM8TRVn7QcX1wWakk4ugW+SIll5Z4QC7vZB
+CKmfJps7D3o9lkgCciROwJ5HVu1papVI3e0gbgolMiFOQzh2x7H17FPaUMNjGLP
0RzcfOKbtczLH2rcEzUD3t4DP/rH0AWyu3MI0/CrTHsscDwNWB/phDuY4Nl4tNOW
YIUik0EYoiPK7sSWfYgJm3ay5QvUUgdfhp0oaKMGsoniMJ4zXvqWdjPGHvue8/7Q
gTTLX98f+gMWJwD9uUXRdpv/0p9bkI5W7TZL+PG0HXWlyRvNIUSQtXBF/VsStvcr
4GNhwEb18dVcgtVTQylV3gkjRKBZ8vr99oLNMVyTiZr1NmbBxxjymLvEyWWW/nXB
tWon1mnawv2HDop4BCxNIhasZahMECK6RM9lkssiPbFBc9G1xNeWI+iWKNx+IeQL
LneaQplU/i1O/d37QmrGwTtke1gd/1lmMtYfjCujeEPoP+9CQj1MxT7eHPZMqkhP
IIJ5dBgFieF7JZ0MwSOC1SUdrVvAqupivpD/ljCZZe2zTVHKdJdul1Z3+OcGSn2w
fucMoirAbXJYKLj9ZTIQkKIZpUJVZwp2zph/1MRgRv/vLUxCvGCS8CWEYJqbh0Hf
skBiYr63Zq+fX73w0Q4SRMBUNKunoJCvhZOUA/ejMnceyiDXGAYWRp99mnesM32y
5h3xWW81lLLE4gDGGSKvSvIjEcfKXp3XDjDYwBzRPEUtluHv8KXUQ8wUfMUPv7sa
1/T1pXLlfs35u2Yu54fj6nQPx3yBdW8qE08pChJPMAiXesud0cL68lovo2nr1rU/
BxQDT4C4KrH7qkTP9QoUqwbAILNMGl04CMQ9WMLLY0rHjVix8TLkpnMAIgb9ml4B
PLdsSnehbgzQUpTBhLMpSfrPT7Fsox47JfW5r3zFQWhFgs6f6s4Mm/1BiqN3xsZT
i/oM8StI/IRXryhAff2geHhkGpU0HJs6Vwdw1D39qdAgNtys2xliQpWwt3RB/1wU
AcylsXk5jRFeM+DPeVEoE6S3P7m/zaoXnmPLTYGsV81i9iqUnQAatrm2tCI2zoJR
T4FnMOcCFW6c58XLe11hBqiD5G47RxbinL6xIhmhHJ3l0aNoSQobZH/BAzZjAb+U
gwVlfhyGNHB+8FO3H5MHfXZ+u9legMJdyEoS6S8W9T12yL5EwctQVk5I3gIMqHpm
lMmvAun98Z/xJY0OWYi4s4AGCrIGVVJE7zRwEtk7d4xxBijd2PpLtYKNY1iBod/1
8DGCPr4UT0RbY0BRwullZIkd3Mp2W02eN0glAA0p/VaKcK8TeKxvxoJC1Yu51zUo
8MqOypLecNJQgfcd+AhaQM2TSGoAtaIXGBb9reea0iGHe17io636lkA6XVBUZV6P
lBDtYCHxcGDqtgDElPGBY0tFYF84DprDk9BGGG2CzzCb5+EPb5NBIQmltA/4+7sr
tcUkvDOEqLRFec2MCH6rsBJacc565BqqdOdva/uiGBDpEvg5J5qQ/Jaxwbb2o5PX
4FToFbuWW+r0Qa3tCPIoP1BnUT2Jv0WRNmIpOPwEh5dEj8hUdpBiydOqN9B133bG
pwFBHqLh/Zk+soZOJ35xoCLQdhHaop93HFcjlx6IWulLgF5ozWZNFXM21NF85W3i
m5kInC0vdNf3EVo8fdCTdenACYT/nCV22iTACue44ZvxX5gFXOrvQJktQzJouTWA
6ICkSoDuDloR4JqUYGCZAhmme6ZP1TqTTFyPmQSLjpzqOUP8TMQraR3fEAK13iGP
sjpUXpW0N+J5kr51ha8NGZU1rPh48Oky3XQrzev76bUg0ypVWMyQ+qXbKxt2CjjW
QZlBNCDgX2cCFjrt6CkbL6uAbQIgh1TNxmNbpvE1McyqC87C4uoNvApw8iVzfac2
uAiZ2aZ/ACe27hhl5zqJ8UjCs1Bs3sG9rzWqG0xGcLv+RsB4oced0ghzvIQvwGco
gY7YOB0qnOky5UYjgNsqSmyvoHbjWr/LcvW247NRAXGu7i7ZY132CYKjgYnFsXs2
jFRFTQAf9ogZFBgoroNT9awUfRIgf6efQdiuJPSSoMGigF7jq2cTlgl/NYJAFHdQ
A0qu8A0dRxiyHNvL6eKYJvaiLEMiPn1F6/aBpA7b9pMJsv7dN3Gzl9kB3Fxom2MO
OWu23SPbQY7mLrJ97+XImTKkbC5m7d4DjVYrYg7qLfnfTZRSbwddgY9aidkEvwVh
Mgiot55EzvgFPr5Xf+Oni63+YUkpWBUyx6ZLItIkIxfZ70h9yZj5FC28HQ6gdDIY
prqOJQcmakmod6K7/7/+bfOWbWaJNXl50gW6XY3rBvaEGvz8+pv8vXhBAfdi5UAb
z4C9K1JkfGqBtvk8F32VpFaZcVkEDlOfDdOfEUHhNVqlZx4nAH2ZrN9Q98ofTDl4
glr8hkTx3cj0Opl8VLqcFpK7RDJC0aKXZyEs3/jnaAMUDfiGLKcZhXCTypwAiMqP
123TsLd/xHELS5ktuvEgUCrYomBg4PiYXt0OBrlgbXrjzB7W68BJCZPfQFZf/s/j
ttrWSqttabshBEBq4jrwzFKxM/R2ZaA2kBXVXRHyVXaC/ZXmLVz7PoMAzLHymQyV
+hnc4bfiTUnTEMzOF2EMbLjV77JHHLcXKA51mDdkhreanTMGhUps+h5o1YBT//Rx
o2y/G6pilASdaP98EFZecCBIWAckZZXRlb90VJoo2ZxP8t7BVBTNbXv4qmdHnSDQ
NXoKRm8ddMt5tgiebUwlFPgf+5kMiYeFGnpoOx0Y4AscF1DDKk+tp6nwxW7LZuyf
kibcJJTYcIR+e2/u4SV7XTG/OO8BJyyrSShwkhcCQPOBe60MS2FgBdwjeUo9dD6i
XKsWQ9IXvBSU1rHY7XUJLQL31ePmp+LtBtQz0nhQrmrIV7lRHzLGmr+vFg27Vyr0
P/tPUzPqfn60pg9YC+32hp3u6250T/7HHmttZVTr2Nn47Y3U2RvzxiYGxd4JZgmU
E8Tv5NRh1vD0Ziuoi81rOFB/SPUCCxrpyCKYMC6f3r8JsY1IXGejHNODvJL5+3RV
k9HmODLbGROcVwvKA+tbdoQ++s7rjqPVd5rZxcRS68wbq5cQT8ZObx5UETFJNDtM
tNXBKXPDgEUvbDNS02+BvuWpLUWhoBfr0UjY/bmAdpsgdryTQaXhSdsBu6NBFSYw
oDBvp42F2pxwKuxAr1tzBpL+Sc+l3r+QET1F2lftNEY7JPTuSwmIEt0U6EUWjW8x
cLC4LepvKm/2DNDsG1A3t5EFi2Nw9du2LkkLhnTE2GHCJYodumvEfLXkYLtC+/s3
zIfGqSaaiA6MvTjZdLmNFCX3Pf2rgiQGe/IDJImCtyoldtjS5+Y7g52C0UEd7tci
CnXED7zOCEtMG0xL2K7O4knR6s53Fijl8MS+bcX3GOIv3/IN1tseeBZWeyB86ytC
X7tIRgCahNmbjgRjs15DQK9KgmMYdGs6lNEek80vyoHe50cG9kX7tyl3quDr5TKM
2gMsigY5by+hHNGFZUa7vmxY5rw3GHAGmm1NqSxCKldyEF64W6nfM1on5HmZJMcl
cKJ4SvjkSZREdo1vZWzz+bZcVh+A+UCf2K+RR6irpDj23pdU30uSzgwSbaigNev3
U5YsY5uelkc4b+lsd85idwYNVxJNoHXM63mtS71lCb3bLulRpxzwN/YGCvtbYIBZ
Ma8OX2FJsfrz1GGqG2HhjHa5cn9J8X6mOLOURA4xyYquJt8OgVHexKoAV9dmCTUu
VcKwnQntQzG5so/1q7beG1OyxFciolhchVsuQX5TZuNafHprSe1AtBLuzWYcGTdz
qlSD8oWZ4NskD0/UUaeWpO2KqAM0JzRMuVlL47R3y2wQ5GnAt1UDcHcdGhe69JQe
ABKOEacLNYySQR6jfeB7iTVuRx2//8v/YQTHsSBhHlw+P7U8OHziu29tBlJDRPQ0
QVzLh5ujQMjVjjD4svrIuqgOYTYN5LqH2bKLr80blkL/WgMKtHVpo0GZmaO0dIeX
Acx76QuzG0m7nlDs0x8FCgg8lYMeqUJpzbCDocad48D6gaOGm2pGZ3/c6SQCyAKI
L25d/XBx9xmtBPFOADDPLLDyGNeI050heLiPcQlyoafMVgNNQq2UUk1pP5VLZMZ9
2n4MqcqvjkXwxta8JxX+J6+apte/6p9q7R/yOSTQiOuJCCCsEIVQ+HyReESJfEi9
L+je0oydg4m+26j4mS3Fj3OIUnTM0YJ8c2EjeUx0ZbBYFDRdXST4PXKmrB4cSszQ
U6oVwRkxQwvm2j79qGGYnbe25qEZXzp1MtALdNvbfb+WlxMx+VEleGHv+3AwjObx
sHJJNQbfRdLPIFP5cbiJyknfOtssmizLzeUa5XK8emMp5hNEtGwUCqH+xWi2xD/w
VG6hKI9Qare1yGTPcXm5D+4+Z0SZHWYOouFZAQYKIJNBjAjQN/jMLMRDdZPVSIuO
G3DKgGvYY4/ehhPnw7j8D5lXSXDYz4xX0lFhL52AYh1f69v3y6v7bUMvTauFyJnO
FnhS/A2oT+A7KASVR1lEbD+0R51C/XtBfAkep2Bd4rlhz/8IW71Hc19B2pDY3Mzo
1wYDPU5+MmzhcY+ez+iUGnUFEi1cqr/L2wEg7tbQGj2HDjAvwlEbtqN/VL8+Z4BU
ql1KtI8fKTbIFZOAPhrSYL0d4qumjJI7mEcTvXdsjZsYlcBWq40vda9rBV5d5tXt
QabcdFO0hqLTM970puEua93gz5b9cBQBleOtymbSfY7NwPH5K8ZKG/6xIOv06ZcC
Mk5Jw963K7JaIcMrGJmxweCZehCIfmcasafmSSnEEgdnWYpFf7t2rDzqcANvTqSD
OSl0djzG+ZY/UdSvh2wrjdSubmYq6xZIdzVKsR2TFzTrwF/yywaj9cCuqlLt0fBn
cLpgRh48tPMJeym9RhEh2+6gmWB5/I1DpkiAnKYkskR2TmIRjxAtIDEuHLq5O2j8
BMgemoZ95Qs/GlRreq+w6KIENSe3JDjFUg2USz4yrY2zitP9H20wYiLnxaPek7BH
5/kPvfNcsZoPadEiGDlEXIkUrmg0IHplECvMvi1LwZBlTgHCOkF6VpiXnVHz7ijm
BuzojOlTJ3mSirHp7SuXjuDNaEE1QcJVAP82k9jMKT591GriTYZlFXGQh46ybKkn
RgCEfqdEob7jlIMmtrwXEYp9RAx4w1JKWPUT1ANbiPFX26D/PnTSX0EqNltk7W6f
Q+4qLVkTP4Mrrs9hrg7vmBh22wNfGeamhBZOU4H4zWIDoiyXB7jHKao7VGIhIbdR
aGgjz/4K6juBTTQYYpLqQ66M4ikZ8Ob74Lu2R2HRB3PZvW0XndTHNITjfECCzEqu
RY3h6kD00oLQcXtNc1Zkv+44ATPWF7pXBsOQqVUG2pQVSnQTxoWXHlHWuoPhz3ta
n6aE3lQW8INSwTCS1dJDtu1WUv5HfSGBvDK+SiM1i2uYUgxft1PxoegyyEs3INjl
Ht8MuyN4NJxSApksRf02xE73H8oooZicY2BhqYr2sQ/nDlZBZROhBWD7uWXS5itY
H3FrywNAJSY8Tftqc8alJuehh7zpmFjcMQbZE4SZEmkCqeH3ESZ7zNXTX/CkNUT3
ymuruq2rdyoVxFNcxpRcxivwf+pwx4rTzOG7ZZD2kY3UQb4wgsd7fNvKXbvxcnrN
CRFU9sPSeVMVu1G8bQ7vOdc/1WFsf3NLLaZLqHaQ7UqZR8tVqyjp5d6fka499qsZ
BtwYeFefmCAi9k8ah3+YvIr4edQ+VK0NR5LA8fz2qGmS3P/FwuH2CQG7QK6LNFTo
3XErhn+5/n1rp5erlwRmVFUPQPDcIgGAMNSFGCnqBHaES5WjOCPj/bELxVvHimgG
CQkKk+axfHyZHPr0O4yBPxE67/TbIvCJxAv3paf8aBCTEWkzz6igpWq1vjrtme80
Fxm00cTEKx0SvoNU5pOY6r+rqf6Yy0L6gQ4VJycktXXgiBdo1HJFcfitY6es6aBs
sJwKc0Q+bwG4lyjHvvOFyi5uBll17v8z8owWoytVjTnQ2s+pWygKJ9BygbL8RUji
R54LKkE8Z8/PtIlj/wmxh0SCTGBg9AKECiQ+9VjiEnpptB9zafVISxO4DV0u4Kc6
g5764nJgNz+UYA25AGmlRAN5wQYnbnIL4ARR7/J0TE24pCL8celI6XZGvzM1YQ5f
RBNIvpOYfjkBwzn32MfzR11e7ofXOELLYhWr5vtCvWkbx+FLEAROWf94li4otEFE
Igax/++NufoGHED8XDHN99LuGH+qeDStbQPGwrEZFPfkYe+VfcBxRERnffVtzm03
wYy/dciRzAImsXSrnelaV19iRlj7e8vtqhE9bz4+6XR/Otm2h4jEj2O62NCt+vRl
WtqTgNqo/2Lazi06Jm3aUFF/tDq7KYyyRsvYK7I46rqa1PgFFHE3MbnOcoQ42i9a
ROlDU9hD08n9nmGzr3lLqIKotw1zkx4UurcHGmS6xvA4FFnQ2ZDKyX/ob6ZqLF56
m13i8DPFPhdTE905aFy3dJDWb+IxaP8FvohnTm/uQTWcPcvGv+hFWmWUqGH+nEp8
rLzZkGkwvoa20GPNlA54h2HlFRxunrk011jPW3Xrw+/BEaE+zNLYmzGF6qHVg5Y5
ZziODCOGB9s8XjGb0h+xVi8xBWX5gOBxdrQgbnIkgCnbDWt5IMbzaE5aM7Xpes62
5XUMVKQqFOIDS4QYFWt6IAmFjYbjC+lbMJfkFoj3oZaWt7ZaC8jJBa7FAUTiKrES
TDkh5roqM7MGwe/KX+ySeRz5hTVT1QrkTFFGWMSByHxuTlM29jsMd+NTEjVRQ+8A
v6Ij8poulnuD8F3LAy3w4cM67KoIiWoIjnigrXMRc9F5xT6wrR/HuXrCI6g7zpFq
SCJt2HBbvCL/0h4O57UHBXorQouTEfNjI9YmMS78xauVVGxSInIJZgVWhuYCsghU
rbk9hVER+9XkJmpPZ1H6lQDKN4UeDI/HIoCIVg8MP4q1oIReESOpqk4G+mmcBEn4
XCjRv/Io+X1+5NMjn94TXMaom6Z77yJPYDvN8zusKIPMYj+4Zi8gAtBZLx6nj9ay
EvW2tjTJEjleSgw1sRei7qerdr2xR1IY0uCvIjmVE33FO6sWpBQtW2gKY14ZiU4b
YZxsb8Tw3G5huxrrpvj13D3gaRluUb/8VsY9jjOVKv9nAZQDP0WlLFTFi03Avex4
wvPjXvCUuJl0DTYuz0M85z/Yh7U/nlJaG4gfi13TBfeqiCYrb/EUpj9P8wAspma5
8W61yCEu1b6nktb/YGtpyBo2vLMUARE+gs+izdjQqRZWQ/8dC76+WjZrMQiyzmdF
ALOiGGLzMomoEoJSSg88pklOrMy75kl3cGLDrvaiLQUu2eko1iaBhD61VfR1KS1+
9uLlEsqS3Kua3J1/V4UyZY8+NIV6Q5Ro5gcNGV83MURWO8uF8y20p9jbgKGfvu/e
86PlKWOoDXi7vBrIYtpsvUwvac2iaLeGZMzNOfAwcwnAlmWAt17ki7rKl0ZdDQ0t
tXbWWSZGY0qF/zS7y/CperTAsVSOZzk1gpjulvauN071vMHA0+KuA/Jtrdoc3+O6
3AIpSoDb68OMRU/FWRkqXe71zNA0qHaI0x5v4sl3j4yg5xKlGZ7ZIcQOukGBi4Rh
D4FJ7wC4qcz/snbbMt9MV+Ekk3bRLDXm3Zv49yrY4Q5Nl/QmjrcSLeUPFp6oLE2G
OmmRfVuQleO1899T/qde2KRR2kGQTkH22U9EO1DU3mx+Y9LrN4GeuRg2gAIt2B6v
fLfXivPMaB45wxnF6m26xc/gDhmNKKAuOcqpK+CWesnhjC9YqVL7tBrV5+1kisXm
3yseqvbuPhdhGXQjbib/wMTLXmqM0qoeW6JnLo5FqMlt9Hu6g2fsnHESUdjzKzwH
n5AWa5gmN0xYEXSKr6Spv6Ce4tuY7jvuHe8kYaRrnyRScBkDniWBgeyhNqPeMRKC
y4pA1c689BIgc9svasO+xC+TZaQSg8p60693JnTPMbqeK4tmaPMeFs0ydLcz9LW1
NdsTGIzj05LAFt3khLU2swZL8TpkzeGOUPq/3+S5Zsfzt6plxVqHGI/bwUMp4nXO
lNiE6Xez9sVAGYMYxcS4htgSob3V6ponhNGfCdqs3IDKdIFN/w8a37lQvg9w+Fx2
RKYlUvUjeGG8UlUympWWrrMMxsTtZ5TsRL/TnBb/l+DRu9qm7SF7nG9pqeSMoc3C
9roQVIJ98EKF8rcAwrIB7FavyeTpxEbbZ6Fjo12KaOIV767ozFyV6KZ0Lrbh69FV
tRg57jNshlZIZZ+HXYO+9JK1St2j7YXATQXgfsYTVDgvW8QST165rZj5c6RSixBf
x+49E1PKIlU75p6Py9PXLrgmv/tMhs6BgS7Tv52795AXEtdkfMJiBL0IdCLpc5OX
3QuOAd1iu5xGGdefX4m2xmKf/DmxUZ9snPXqpIbyzL1OA3sFKH32p2EVkiszu3R8
srRhIT210Jugan7gt9XN9j6zx3zCtH2/hXgbaRPtP2uxEhk9Jy2l0XEIgX04/Nqc
pqs712DDeYWdqiqH7xdCr2cw3/8sePhjN8LjA5oL8yQlnkAkfKRDZIQTUAzjSMxZ
KaKjcrz6kfVup9uI4dW/n2mcQbUGbF7rvRrAk+De1Fli4v8E7pmeA3U7EvZFeOGP
+aj9/pIX4c8KjGBP6QDw97ec09RnEg1UBy0Xj2HuhZshMcqY67jU9yz6T4SDrCK3
aHzXXzys3e5J5JED+g7+AZqXbvXf6MA3osokGE/7LqNdVBwbnfVIRukjNjx1QipP
hKvz+A814Oa44QDNO5MdDBgAT4OPPNwULP+fEfu1WAVAZN9XjSxui4xWBc+Ug8e8
QcJG+DjqGagb1MbIuwgewwtGvatzWhI+pCJctLJzRyN/RApv9SGpdjT9iqx9xaWY
ygGrL+05NY6Q7sBH8GN67vs9aPremtWoT0NsxqDI4h8RgXxyGo7AoeYKJTbSE00i
0g0c9ypbgopotsO042+uV4BCE220XT7VUmQLOFFxA1RekRa5WqfwsCsRzylRm1ax
cVYGNmZg8VF1ERzlhGmWxZygh1v6QBlDp3qQU/27xnreed2XUiUr1mS0TQYTxuj2
RdWGzSQ/vE47eJbgktEEhGWktvJdn0ajgWek4/E5Z9QWz/wmryetOWgZEV2I14tl
aPAxvUACvFR48P4mzO/fRfHoif4HQ/JCmhRoSPRK64YAxbNGywDyxJ0BSb5CUNd2
K5bwGuDOhCbj5n49sUsgaA+xDUpfAJ8x8s0nBQVyiacV+zs1pqi/gnex/kvFYoB2
SMGQZfoMi/FOhiGBikJu5s7kNuJpUan5icwZVOA8O52jMxUv4rQv0/PFmWWNj9y4
yUz2hJnNJmKu8ub7BjlHV17c8XOIv+gurLLDyoOD2nTTsqBZDr/l6tHKvM7alrxB
IVsjXYMIbVDwZ1mGvn1fpCvxg9/OTXgsmTKnh9BR0pknc7SXtpilWF90BDqmxPki
ooeBfgRe9xwQmenjabChKJcw/odoJ0OGlcsmsZo9p7deumImtm2dGUuB673pDW4e
v3Jy+0Y6JQ6O+zJtDD65GY+9HQXVl+qmdOYfywQr7VYS3sm/YwNw4kbVG6845pmU
sW7OEZ17kcV/GKA2/itJ9YsWIgkys6Url4s7Ls0agFuOy1bNka/ejLxypK9aBZBJ
naBT+8aaH0wfqdlleFDCnL7k57AF7HxFv0TfahHT0iPEVMppckKoetKeA7C61pFe
UVajPgnGVwYXwNRFvBurswwWuazcoXKIFhB6NhCOojHImASScPOPQ3NkI74agr7K
PRZX5AOhtfbk340yTWW4XN7AfnEnkEVTW4xyrRmkyKKiJCOYs/zOX4+8ZzZpA00X
yefw+nLNn4Sz4FNkuxNEvHzCS5NU2K/Ws/L/RO5H2ma9ZmsT1MjpZTeVuS+kqifv
N/y5GbF2cHBToFaVv9gSdrNNXKZwRtTVaWwa2szAIbcfUHAN6JwM9qLUPYj635lc
AckaR+J0yYOdkNoSskdCvYH/48vjzpZmH0IRTtj+pIejf7spdCOU++kIrECHrcgN
t2Dzv4o+rmYQgyWNzVnWasAS3IpDYHyz53Uqzwt/ER4ZhWwm7Zof2IfgaHVWB9uB
Yow6tcyJ0Xl/QqS2qxOO1nt/yKSlJZVqVyoba8O/znf1k6T7NdYCAOo6Cvwpn2Ka
qeEBn5xYpDGTAV6W1NGQu9G1b14/PACAuo115t2EGv9zsavhph4Daimer2fwtZN6
/QDN87X8hDUZYmqEfYP0KiIFvh/CMpoc+93SEQXKgFBl0C8pI3r5KOc2MksUw1zF
mPxgPm7KJkb6DGPIK7qiqIAyqw9gDW9HZXigzayZj7j41HxtI7h6u06TJuwK3RAb
n0OMYnBLto5OFFxJi2QqCB+jQC5k4j07SPqxhIg+z71/tRIJGdvENbUsy8VTB8rc
kIwVk7Lb1EksqoKgG9dQtejirLBvvN3nUVrINVZzecyO9Q8pEuNqAUbV4u4kJcWt
bxxpSV7xbTaBBjS8yoi5OQu9btA5oj20EEhFaeiVuRg3FeTPZ2sZKW6hdeADwkGk
NE2m7Ksw0nBxSy9+jxQLqBu4zOb/CFRVDl5tjRjDsNjRq8TVDyHZgGgAwqC8S7kY
F0xsMV7pjKWPIC5w+sOJiqU0lK/WExNRtTpGZ/SfxPyaGecB6PpGkBrFcUybBwRZ
Jwsywaf2TIIZ/gXDPbbmCQlK9MOoPy9jlSgqx3b4YJvZQt1dL0xI/qohta27WqOO
Xu0GIjAa7LmJGLhVyi4k8hoPJf1dhVUiTpQR/8bX+Zmxzt1cCA0003q6x9M9S02g
afBRtP27aNlyU02yGfgNFY+hB3kwzF1MYmepBoIVhxYaq0VEhtanWkE5gHIsm07f
IkTihdU57jIsqx/HM8Jy/qoDNRcLH32ZT//MYyVz2wWejdsXJ/BBZRTcZxx/Qmr8
uRPk0gcczciMjlSx4o1QiIuuV4NlxJ5pZsSqkjNMqoLV2mwjz8YVFveYKpLAR6Ux
bS0kxZsds5NJtBc/luj+84WL/UfRWBFNxqubGPBAsGrYTbh9fnyvsC/fgB2dufJ9
392+0CzpDCRtCMOm6q8mJiapUeeN0Y3FH4zziZRh/VWZ1rSbmVsqfOWw8NtU4eIr
kI+Inu/S7wCRZEKb0wanGOzM5/pNa1SR33bWZGgyt2FP8tyR/MN3qTmRpcDjBH4S
0hu0jxKDIH7RQWth2yL3wTbna4oMbgC2C8y9xfT20BAjXcvaoshp+lPwFd4Pgx0h
PT82jLLrtDGBUht3ZAA62hlIsyI5h2erhuCz9Eaa0tmDFKCWn8i0Ers0IvPhrvNn
Mqj0+SO7a/yMUauWlVYs2zP6gXWjcQtu48dYCkoO5iWKz10PYMLVSxbOUrZdiQKF
7OBDWMrTsgp3ZE988zcdmlQX5NDDEo92CzhbDu+VAO94PW1DiPs8MRcI+01ER3rl
e3ce1k8YwGUu+lKzyIpFbsP8vVBHCcXgPzCTKUmyb8LNQWQS/VjVtRRsyv2WlhmH
MonMt1oCgpT5zGs4zp6Uixtqs0JfB9Us2gmgCt0j2sGp2zl46n0ZKU+XsSvZEdJA
vBFoFG7KyqODRVUZc5T2KVPN8jRaRqTgbsybfDJ8S8YsId7ChVvyafaPg2mTh+/T
/9o50DDE+qW7VvWEFSGClxzMwauwauBFXIyffXoP1+Tsl54oOOpf1CTfEKhUaZqk
8ILrs8FNBDAEsiMHLIMVzFLRefa0cVuLwNsqGvA7HNGsWac9d5XXe5xZrxX3eyHr
vABSvrzahmMOaNCqv6iFTwmSh7SKqldi4SBJDyb8JDY+NCwVaz/DJa87xtj4G/1T
QKWeEjKHoSQniugT4dFiCKF0Q3O0Kz2MKLnGthj/zAMHJUzG3cBN2jKf9XLbmjMH
C7Yy9yVYm+WIpMXxw9l2z+RrgKAvfcEWDhaCEoQni33KaC1c1bgemjZcM1BuyHOJ
ozKyeP6Euj7+1OzpTp1036PmOfEHb3qVgm4gKqgjpRGaWBCJN8h/OhllvsThkav1
+HKotYhTZQ21xQ7Jn9V6cKAFbNBJzkmrx4A/8J9yOlexN2Qrco5y8DgJdRheDN80
0SABUpqq90VK/J7SOg3PXF7/3w7/l3XU/jgNcWztQ1hcgWSQYhUuSFTg9es6YbDi
LebJ5Yzv9zwahAftCkP77REdGgLaHtt7P3uT/NIVt0o3C1BPU45JeKuGdpm+6j5h
hMly0pusMnIvyOEcShy5NPJuD0k4Cd7RnBqdKlKIuHqGTfl9dMjodYQJmuCRWF1v
zfZ8gf/5fThAcseW+q0CvrQxVl4CaJFTVDHSIZ7Mdo2mpiTgSYGUS5xLxYUsBL19
36hP9EWixHwdZFZ1j/UKhhC2n0V7CR5g8GM2Pkw+1R4FSWsJDIhVGEn/XkV7WKlf
u4/YEzLT94IyBSNixnoTTMOC9gWT197eeFcsqgP884Y4Y2OShgFhI8J2LZEIuO7o
MaHomwUHJ7SVzTb9cZtYpc2tUugLmeiwv1RXj3Sc3pPxcs/t6SmC0KU+t+wnRD8V
KDRwDE1johej7ct95RVHTJq512hVARjkR6Y01eoxA4NH2zez7qylw3c3T3/i/sdG
my5oEC+S8ABFmw55N1grZElFrvupxKKrcQlr5vd3gAhWXawGdcB2JZ3me5IJygjl
JO81O0nRk3VdQNyGNpOgtdSg9HcNB5JS2AsXMYUM2Qof0mZZdn3MiKF6jNFC9MoW
WMPcy6NBS4lNb/YEU1HNwaJeoCl0R6Hq9oksze5jsT4g1IRjebMhltbw6sjNM0Qf
xHtkCvYu6xBwDYxjo1nR+Rv2g8EyKbJ1HCgU/zh7FS4qgkq3+nWR/Et7KjAZvblY
r+mneV0G3rWzPLN/Q5IhhM1/IlEOvd1lfj/Lo5SDtTMd+LODBOAP+HOG1DJ2Lxuz
Nc6eHh7cmVWlVrg6eLNXnsZRt6I4sxK193p9hyxKxjKlENAyAeULYJK/YeYmk9MN
dPDSfL1lftN2DELOKRbO2EHC1lOwd0CY/ThUScNkZUzSuYpSt7ve8xWi2kYdqN+B
9ikHRvVgchD8cfljkdT+4Elmtsjkg4cYyDTuM3DLBYP10dfSmoWNb+I69Kzvnf+I
CGetj8a4JFwMWasIE2eGQb2lQxvmbMApCclZoOnVqkOuKvJ3JhOxipP6j7aKfeQ3
UPqwaGaSVymkXIPMxFWxQCG4s3tUZxIk1q4YyzrsiScAcNAuqso211boa+AmS9a8
xxM8sjxlp1TiYCGBd8FZpl8g77Iukz6gykfy3EfJN1WxEePyGelD1aWtqMMUnN9E
xflEMa3C/2Xp9p6yNEPYAUyVYWzSevKKvQtf35nSz5tLWKF8KvysElBWgZFyTTsP
P6m/f6yAzeyL76onA67jJptOGFkzHl4k08I/qC0ys5U305D4TItVoe/Vz+paaicW
Y30n/27aciVqomRo45vpd0OuhTiTXE7PO9pkMnlNCYJlkHb7qdnw5KFmiAD5QIDG
rUgIQKzpyB7XLb6EtFe1SoOoKD0U+HQziCb2WFrRBbKoM2pqSX6S4DWcwBwrmSzf
VMcl3dQOSaYXsRJs7Ul7kZFNShqkP97VdZhiRQXto479v0GdnG3xYg9dxJo/ZA2g
0HNI6jqUj0ms++NCqBcJIi5CO5Dt0zIFibKjDcNmuQrjQmoACldGzCDW2miKI/+T
DaBrVJ+tzg95+GFWeD/2GG7DvrFfoS5TssmgeRC/3HoFbu/N6wTH9gAfVhk2zm2a
QunNuJUjdhmsLJ7zptEe/Oa27RQk/tw0O15cyaNGH5KVW/7CA7hsUlgUArHrLlzk
AQV2f+4PVPmjNlGcTZ9e9AGMAajFCMuwbbx7P2c20MvPhPBDwUMwTTet/0mJaRnT
xFYrCa59RcZHJlNNZqq6UAPa+bIjX1eN2uAV9++4seBUVti029eR/iOPzB/7EssE
J2Z9ocUPMh723l3c+f2oFI4n5gPPJCY1m68aTDBF+G+MCpKJoE5JCHLypCBybAun
rUnC614fgX4kkNA1aVbbUNFh6deU2q4zqfayR2vGPA9e/uKm4MRI3L1MVepyh27l
Fwgj0mTtLKJUk2U43ZAi1vXmeX291RLj1gs1haXkCXRiHYhyOHVrk0a4Kxmdo+z2
uH3aXCrphnL6ijNbx4AoO+xyKR3QFbg1wTnqPX+h/mQGov3N/0g8uQz8AT1jfHao
3RmpVKrh9tFDIga+YEy/RIGcFb28Lqk8L4HFf+5Lk7CugB61gs1E3PnAtAuYtidk
j+PdwrsbRvVsl1yu9jVthzpQrKXM0uhtzmdTS2B6fcQxPCSXMJZLV+miOx++gkLX
m1xpBrRlL5pvKv8atvVB3g4k1CSHVoE93/lKJLcVrCusy1yZBY49TxsMj3THqE/w
kltbuRpdeeMKOApMPdqsrXG5EsU+OFTBe8xOdoHYZ+RPbS42uaZInXCfIiqbIgbG
84zO2AkLYvMA9gNldSjCl5cO3Jw1vTCrnGDsWXnvDeBbgPrmov+sOXUABRc4x9m/
KRB8atuYP2iqj2Ef5BeW7azUNAzl8AOqoMVcPQ4cavpCuiciKRrVQZtVkPo/gqWL
iPqgybRzSNn5uCKP7h1kyrFKDigAircD4JC/xBA0GE2ttgUK8Q53OmQQGzQakh6q
Z8nq4O3FX6NnaSoLq3dfG/eGhlo+EARslEalPuNhKFq9oGRRaae0sjBEiEZnJ/1K
svad1V36HFdzZvl0NcvLAkyhhOn8j+g4m887jUA5UCWsbznHdjrUHCCJ1Q9xFZ+o
8YEe6RKymEw94787pxIkjUhByI+/83ooKbegHqkPcd6eoOWjP25cBMn56N05Gkbu
e2dehsg4mXR74bZPHceag1J4FV+V9wUoJtAfFIPiTVFNXiblPzcZIyRFtZ0g5KSe
6dn9AdUTZI4iqT28QkHMY/BLlqwC45A0xuueT/NAkm5SMejWbEkLQpxyXfQoRjSv
iXcYRLZOnEmMEf2mlZdb91S+YSbvdvGreGiLVtu8C/i/b+CRAX3Vz0m+7TD/qg5e
QTTMsZlMdbX05JRWmtws+8/Mp4O1JSPPQqa6Z4DGg4QfNUOTPOQS601v8/YDWL3j
PZizao3Ge4HPsXn5AXtaOYyLSHKf9qJy2SvRHn7TFRS6ws6jbc7lmjv9JVPl4r0z
+3TLqVS6PCs0RKdJVfpcY9+XQbb3nZIGyzvjgHz7zNKLxO2nBtJ39wItQc6GBrxY
9jdrJdtSxwLovyfNfaJf4F6AOb1ItBh33qel4d9fmSx6VSDJzg46WG+poPmQMSha
RbiJMXMqEPpCjMG1dthP5j7MajOhCLAVugneTLKJ2cDKA5V5UOGC+ux5O7SfzAOc
JI1eK9qgiAjOtzq1pmJs7uiEOkPXe7HzdVjup+c9ahlqOQgYgIXeRG21NtMYdBhz
vcla+PinsgdZf+2ZYzYD7iiWdEqbTD2RYMgPDTtXmcmMUgH45EfKAJdKG2UdU8S4
hPmRXg4zjMkqCvUIvlTMffp1dKlOi2a7lQotpv2w8HprOSXIMoMCsp37O5vvoWe5
5Sak6dwhZdls+FIHM3yPcL6keBMrGRDuSUFvKUAbKrM7lrAbIC5crVgV33MChGr0
1e1F/GDBwwLWEzTlWmiQWBLi2lG7uBodZh+c7dpACMcK0/9eyHcRXSIElRQ9nEiE
7zrWSyQTGnbEGOm1fKsLqgryYySImVlLzErXjlW9wX/noRpQSTBn7oJaLcuYR/fo
jQtZb12W1x5sF7rZClJMBf3IZflf/qv6v48J0Bye+OUIcrasTCFw7XVIbPSx51Vl
jP1HFPz0O8cfycJSvzUMLnreGrifdg7ysxJObCfjq3rN3iBxufeJabIz9Kg3BeMx
QuZwOfK6P7HAkSicPXYMOebSYzEFCCZtAYpAPPs8YWtnUpri0PPYC6Qi0Zb0B6Lr
mq0ad+jZIyvLPkF1d2EvbuPvTvycoiEYmVWYCxRHlAeL2YkQ7KPZp637E7/p5lIs
bz1AXKKNJ15nd6Xw9QuT3IQ0VK2w5RnnJLN7WR3jlyy8IpNDsWdikAUetbdQZYdG
AnqDU2b3Wc33u0NxpPe7ohZKpgD82nVBjGnBG6h74tYt6JTFDcbkUex7OO2e+FPc
QwwBei6JsB1+kA29SqP7+MQiGRpr4LbxF7YZ5Gt/89Vo+ms72itBL2T6yvqlcbP9
pYYzo4T5yOcBPOgNm+IiN/oZql419LBjqaepaFJY3whFZrS2af1C8SI/obGXaeo8
j1hq+O6zeaiKuL3HZADgILXltZZycCvDftf2HykqNr72l2TzT6lgBHY2Jhgn5UTF
O+/A8MlBCBtSRSvVHSFv8Bh0EfAvP1dmdKvfef8wl3K7q1ASBTBUtBvCEcec41xH
GHA6gw1AWzv6+VkQl19OqDTydM39slguzvriJScKDhBBLlNUMa8C9861Gmaqx6P3
lxDdQSRyu3r7aJvYGwzt/xpuyYRhC1PbWAhvncTaD4pLbccjni4ZHxPGkkezjooy
Ac1hGkrBpnr7u2e/PRLURZetXa7FiQXFt/RL8gRJrFnAnWoBqyH1UWzoxd/QbHuE
k7FIBsLNMeZoLltboDJfBlNmN0oUKJCT84Ph2cakh7FTdE6V9xraVaePvjG4SYAM
wQYR0rEqxTDr+DqLSaa59AJGTr3phZTvV27eCP/kYEHHzQNG9c4D0QI/ORjtrDsB
EEiHUfLi2UzP0OcpnMxi9zXKz0b+YDBovsqgaucTeSHSbf57BTkxWYFO0MP592+v
uuFwXAyXMjb0/ATSoDjqUP+W4+Uce/TelfJ6XAK2ojJUlEhcQVpgDCIMs7sVxffz
ix2VBc3EPgZ1+Q67A0LfzYTyBW25SZSZg28l1G8hNLbpmYG0Xt7VZVOg+zEPwSvC
5jND3lFDpw1bEnKw46q7e91/u8iX25bu0myOEkVrE4uA4+hZk6RFLNzkTxL6dpYi
Kz6PuK7GPaoNYADG8QUBv0BOWz9ihi7qfIKSeBn6s8mZvVQpw7ABZMA18JxQ+8cq
bFVdBLX7aoq3XWoj+Khsac7BCiLwspQcTApTE/Kgj6mP2DWdgedy2yq8ombdjuAQ
6Jp3Td1fW0wtX+AoEzg2Pg9BtCFypL6kmUpG9n8fLRSncTJI5NiM2L6Xr5o3BgGT
XXvrfMC5gqFJLqnND8auOgRB3Wy5y5KXVaRjpEC+eODFk6iHqbwv1k9JmWM4/3+z
UwGodrWc+kwaBdeBoFrGSFSJ+kJsB5HR9teTGEB1CEhdd4YRroDC0EZxhu1sRt7E
ngdEp2CfFv+64fhAMn81Vof1Y0+0GHg+csPDfrffwmyV7MABQ1XDz3YGZz/v9aIA
FWCDggO14LcdYZ2AkqixiBdNlpM/kcFxVaW6/vcN7oYZ8SHWTQfQF8VzhQ2bupGJ
1H8sLvoV91x34mc21+OXhKjT1uGlG+1e2vV8u1mARYdDmWSVOQKFWPvvcNP7znFr
iJ/BO1p65gX+R1eoTF7m/3ufhJ2UdKF9xaJ58gYD7W7vGqVRK3QL1mPqSuuSmKTB
0PTPfDhFHruvx6+hIJ5EOhZTGr7L1XjXtzUMidHUlEuBSOoqrOnFwk6hlLtLjotC
QqCkScaIbVmIfOKllHi2K9buZJDREaFTtQLv9lxhowaIYSkVtD3c+OBsiagUD1Hd
7UNTQC9pcP2fpSTmSLlfbYQg/HRVSxA+ypS7L2M86p0sFs+zGEIRSdnXHlUXpLa1
NFViznptEJxP4IaKbwyffvv1JKchJT/asmwFhWf14dMw+xygQSyFUtY1bsZ4gQQx
/OrwFIJpw7s2IXq/ZopSOz7RXcDKPNXu3QeZ4t+Zk1DQ4Ki8pwvuuGbmOsqaAQcK
39VYUplIEUkd+nDGL/poirrLUuGHxOqY8ogPE98xlkho/NNAypcbFL/3vriivVmn
65F78Jt0w2lPN1GoNjyAe+AWBJZQ/S5Orx0biqNWGsiuMr/KiY/NRYpVsJOvk3Jz
Bq5nbbu6O6xHya85iv8wxB639qfzvcvqUeYdGX3BwZ2tZovJLN3UHNgtgJoyUNv6
pvIF3wxksIGdGyKvMiIB5ME6Z4V1Xa5tm0GU80RF9nfBKXEXr/5TtYN9450/xllA
1m/Lw+YwY35Kk8UrSqkQ+/x/MAU8eBRsirUvOB30Y7jWz6e2vRbcU0XtOYvBEMDr
uKkbitUKq5lnR8e/wy6OB5kPLMpOHYZZjaFFkofpqP22DLDoMj/tJGzMpBi2+4BR
opRMB/wh3HFtPScIJwV1CFS4ULqoSjvC7pNgo3HVZMAtlbQVmi+Dp8sDdTXu4VJ4
TG4FRCFh+XgX1UPnvC5g9BleExMLj3GJ0xztX9SKo7XAH1aD5rvnWdm9GNp2QKu5
5VQPlTUR5dx7Hb8bvxZFJ8HGV/gaoQs9WJ+p0/BMMPy10GevhrJsSqYhhSQqF1s0
2zJ0P4v6491OO7p6AbCviS8hT7fgIxu/JCO4wRtH4LEJZFGnxIJlP4N9lYnfWj56
sudIcO3GcwcFLxdP4mnWF4R4sUg54nLjz5d+1+NI6lBI6vQV3EbFLTzIwAuQzlrW
/hCSbWEtK34aVO2w2LsyOR7PVP7tYedQ6cSkA3rZDsRYjIlI5GUTaEjHTZelJtb8
HFf6qrVtBxo6Gu+tLpybyFT4MH0MCF+qnaEHX8qx5W1UMbJYeF6kut/pQFdqmbHK
fVpZhruls8X60440eOXSjTWhpBgwT0Kqz1cQ2tyy3TChh/4ZVBOTQsWlc2Ua8kVy
8pLIrHNhivvfwzVAEghrm0gw54q8OZ31zVyaa/ilB2Dk+y+ZclZ/yaPs7PtfHNi3
1XJvgdF7oIJuNCrRmaNADSKJuPpdqLBhFgN/NOIQEiZ03kcBGQC/6HZ6r1OEfKYH
JKM1HJozY1GmPJHc7+2S+mDgOatB/sh0yXCS2QayKm7ET8GBQSR/83LsbLnFA8QL
AXrFFzs3S5rwTz1sOWwz9W5BnSY+ecEgJ1qvRixY2mbTikHnptt3GR7nl4/R7Db/
k7nuwyjFIyHGh1+Pm9h9QFL9vSt0RG80vZxroWUw7EdYtb48Kdu9XnBjAy4gKjCY
oBDXb8vBH5Gm23nGi8NS0BH2YTPKoSLJwhkw9StyPkgatAzYTH8gFPYOsyOYQzNu
P6bJQ4W5vq+I7bDZHz4jRRMRXsz23c4iukQP7s+PFvP0NA2mJKvNZ0UDeude5ubP
iK2PEN84YwPNw9U8xVNLa7VtiJj9Mi5TfiSe307RcywsqjTMU1kEYyAFwSKqYTe7
4xxke7ZOW/qZlcPwpoeW42fO5tJjzXWzy0/uht+WRfkIL89k/YhtJ5JGHxbKon8D
NYBNQsT03gfeouXFtPzPZPLJo0557189OfMe/+lG49EARucPUlllGHPW78I3eq9h
zPjmGY5pMCzz4y49CFk3Vt5A+4XmyrN7v9Gaenl2K+5MBcKJ01RFzO3wq1HZH/O7
ieQiT/vT+d7Q6+DIRzVROhpSLufaipga4iXu7WR76GiCUOfPSEVk5r6+ftrtM1Cx
3hrvLDWN3JRLhztB4+0up7wlCRhJQlptRnUGicjUbZ7V/mIp+JKDjfp8kDYRlVe/
H0vQ5FaP8ZvO9L5ZyxACLIepthjX8+VBLmud0PRn9rJBKmey761CYEM7WA92jVP7
G0Nmb4s0VI/UXKnlaVckWluuiIAgcgQZP1X888Ow1PZT3fyC7R8G9LvaRXSF7fAc
VU1U5LgrqSp221uwm1WIVrNBZ1pkBEIPjs3xNWUy3ofwttigx+peQReJsnbISQn5
00m9UcxfYNv6wtbJz90y9TicW13tNEhCrpWWvcf9t8lanIUdsTYrgODWSbvt/Ffr
VMlfdwnwbkDbchUuOb2PuuWNH1Gt6LvATAMjdeaNglulCiK74NqqAgnspkQsa8TA
eEaWiaYAAA668UbkekTKOjTdgaCzfXaSMBInW+RQbfsBxWTYxN7UaOtJI9WxRb9D
XTVzYojFmgX2Hi44jVczTqn4n6gvCNSNcHxCK1KL8K+X+AkbJafQtAbLQzJpvTax
2SRDCr9j6Szu7hfozEOuG3bEqOvmPDDrU/9Q3rB7hhBLKcD5QMeIxYGgRWHM/syq
HBC3UAXVKzC6TJfmx2LjhHG8RHyGoMWfAZqS8207xmvZdATantAiQtppNxDWA5Am
cx5aLWDt3BU0T/I7UamiEGnpPnrp/Ffwrom7fqGb5ufqPR8S6erS6cJ1TyvJMHn9
tXxMQWPO2gm/WgXpVFPwU1OzIfP0hKnjbazuIcBhFPGdnITT1AwQeqfrSS9WuJHM
esiP23NFTqDvrsJc/SVHjdvUXLKHbnBBH12eEr3bn/FGb68rydy+ubbEbK5XFwXK
jourVM+UKuI0M0t3VndXggYI/sxLoTh9hB9ygEEPLZDxz8yJFWEavBepZXWzBxDF
EIKDqDd/rgSd6FEoYKAUyBMdH9/fFhu9DSRLV7qdtHSDLQhr86u8krlV9hywaYiJ
CyUNrMMyEbmJSRnR8smSPrk2JGghZRIbrPpI3UuE5Qy4V3wgUE8PBlJGeWIWns1y
sBTv/u0396wSXi5TJFVYjWDLRKQxUFe0BJtGQhldZ8j2UZ03apTibIpLZQAqUuG8
lcbDlRdC8vrkDs7o8XaPaKaP1WNXIJSifjremqo50Ril5k9Xar0vk1lqdR9yPFCT
OY5UfxkgShCSL/86+iuujYn7nUDbT/LJRn/vj8exky3ivk1In9xw/VZAlM4yHo0E
9ylBTj3ZrkWPNjpZl9n3hg==
`protect END_PROTECTED
