`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EWQjYdOJQMP75k/FnI13RkeIZA+hLKiyrUDuBcm5tvNG6ME1VkP9Zep4O4MbBX2e
j3FjrXG9MdHVpdlr8bPUaQTWCDZRpldyQPAyI0oTZyxel2lmlaZCpUcS5tTWDYVY
29N0SeiTSBD8gFgPhUJDmyg0dc/HcHz+fIqLP0Ei2TrSBK6d87TjwzHo3ODfv/Mi
UAxAxId8gQV587sFMI+7Sg==
`protect END_PROTECTED
