`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TsLdR1gX6qvtolsT6QPzZhUjp4f0VgIhiWzmf4WofXGWddr97so/WFX5fdA4VhXp
+nuyzYde8XSWNTKPoz7IM1hvQJg+ldxglcjhEaQ/RgRxEHEiacrPK3Yu+hNRxcw7
4JM7vW0ZoGy77S2nQw+6YwW9f6dnvLYVnUuln/qoDncAC8W8UNpPjG9kxOw9XcMA
YhF1QukZMHD3R6SeyMzx2Ijt+ye2C04pESkFgEl9P3foPc1nz025Goiv21oDbDt3
IYMWwvRQTwbC9FwQ610PEU4bkwncMuVWoOrMn/uMPtGqr3gqb6I5Og3NMeACwIj5
xiIfB85w/Gf9CBeBPYA4ZBxewJ9Ep6/OyzNdXX8cJGK1IIMDm+H8Mc0o/Y5n/TJc
h8HZ6vqbe24QhqBy8NKT8btTBDF+W27KTVGO1y9TLv0qRAtArIhSec3AnvPFsPnZ
QGTIbYeygwOa/hMFwAtIp3j5WC7+cW/XRCIBRo2hJb6FI8Zug6+NW8PSetLrjOQZ
oLs1kHtNeSwepXqC9e0y9nLDxpUXVWl2n5+LB158gdmPgaa89OYl3CCrmPnZc3X9
fJdbQJSDzdmmqyTuhDoCrsxIrI4HD0f2NMZXBbntqul3250Km4n4yLR9NBiR3WTh
l75zccGKhIkMVDBxKgd6kcccg4ppqn/MkPd3+S/QEpGBYjVmlZYJmYx58q+F2Myf
fapPVWW7PJqXVibtzVtq/Jaa0HB9kS+NBQ7oEyjjWtMQSGHmciMvQkgQgfUx0ZXW
Raktvbdvk+I1rEVNVH3nbjOl9vaKqx1Dik1C8/83TKr778Fom0pIfVNgODqk56Cj
54NXLujB8+1RaDl5j4VeUPRcQ88/3/eSQ6p3hL9l89zl2yJ2hEGqWFIZdnfeHQUV
oQw8p4b8fe/k/98abWi+JpwKrcdbFjy6xFWCBQtl/TkISYI20+xmtWdEWHa1TtE4
R3N17W4JEU1uuc/eehWTnL1VEyyVDizmPbeE/DnC7oWxdzvXpZOya1XWiZeN4xf8
mhdFbp3UIwaCzJ7DnZH47fFITMxI23gbfxdoO7/5HlpK5QE/1dfWuI09uXayK5R8
L45uoyUlcR10csGipXA7lk/S5X0mtwMbHW1R/7t/2G+7wFJKA08lJL4/9ogtmDeC
qp4ASKnypsMqkJe9v1ORWJxFBpTBtuaXXHmUtVMwywU0J2TOmJBCT+hwCJ/ctQtF
nINQhYmwe6sZD+fUdE7GnSG1+0eMeSRalQAcFkPMVNbvqywEE4bV4/K4tdAT7iac
AHITJLa7y+tDedZAW/wIv37Y1C14tcu8LkpkpPND7FqP89fVXdSgrrXTIsVN4tnl
ia2dbvhprbfwUcUkNtzISYfSm4ZwYE7mJf9TTFKJZhaj0fSv9IcpoHhLZWkZJg8E
tp5wF0XmARwg2sW33VJv05EzjpJbr0zy/w+l4lPadQs2RG7FlDOHZ86eqUjxMtAz
4D+3mAOxNPuebB3/rTYLPB4dQaSzyqMsXI7LOSJ8WPQrs6I/FFcPF92es71LvkzA
JtGKiyxLI2ZgW0Liz5NziF07CSvj886jRrjECeih7/jh6bxMnHgGtFORvZ3mmgmp
0Hai+vy6ziUxjUgtdYgIKBUUuBmGjeQP9TJg0s0tPm8VrjPVzLqXPTKORNjjTrL3
2znf9kglgaDxRNQudA8x6BhF3BdvQMtxxc44/twCCxfnySeQiilFain45siR4yJx
y5k/wcpiOAvTQEi8svEaKcLJ80QLw3q5wcTYytmHvm2OMurSHZcpIhDR1Zvmvhsh
kU9EpMvZbU6I43+h01lIinog450XQxFNHOljYUskYQHoNuszR6ytKyYNRn9kLB24
ZcRwOqveMpU54pYBgofzVFKjPIAF5J3iY8XJOnHwQA3kafiyLDuCVncMmHM5Ch1z
R4eSk86ru9VHeBz1lWHhQu6Pt4U8MJ73kJLCCuZs+QyuBhISWRM4gVcTRi3sC+qS
8OaxC/NP4/NFBHRtkZ9dfT/fH264nG+bn2EK3VSMLisMY2fbA31/JLD5Uf3NPOHk
6kNG542Iu61wENgHbStODpfUObiFam83qyESUCVENURLMMnoIXZUAX0hU1T89VWQ
JoG3PKgFbH0cKEJduUr2oqWEHQlbrjZ21I12WLP6infbko1DjGOKYPywF8s6x/mf
`protect END_PROTECTED
