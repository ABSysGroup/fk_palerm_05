`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dWS1/udk7YxCylfFKQffTwNAOjwDweJim+7J2WoianFvNNEMPjyhcivFG4mDv+4E
16PnicLNatOefbKIR8rI1Zx6RAGkbkjIcAk0wN0HthmuC+EUgougTsXvJkX+CxGp
FLYjxg/H2s+n6d8/cm4gg6x96bc7+BZcdt+KkvamU/iFD/K10LaqahKHVsR4rxxx
80nLJZBx4nmjEQPpYxZsrARIrN7Hb8c/+91K4DCTx7TTIDD/FmzhsePlw9q7IlSM
aGauze4St6ho/nefYqSXvW7wjNqgn0JvfIZIecjsIMacI+6zGy3sHYxC4hROlx9X
Gfu8Igln5+PvkvucnPVMINgwYppRJNNJgp9y6x2vqyfRdlheoaO34e+WSg/RMUFj
NDGvnTpFRpAtdT5G3sAMaWRrcCwgWKsbc48ukko6dAzXroq3b3zH4O8YJJQJx0hp
`protect END_PROTECTED
