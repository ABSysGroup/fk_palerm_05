`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TtN2d3dFXcxOa0xnVM1Xe4P13sQ4XA5MpJX1NxAK1nD2XkApo526CC9cm6WM729+
fxbgD54Pul2J3u/P1IwKgq259HgFS/UylzQuc2FmeBL35BYT4Hijyq3RNgZJ5ZEJ
ufnj+EBIvbHI4pJg82M39cwXIEaLVhe30mdhJgVpPMvc45QTQi3P3yhDLP+CVWbz
QfNPaAHh38vv/OO9e5KjtrB9i7GQi0GvsqO4ktKpGPF78CD/c++1pMnd9ifwgSza
UKPaPFFuSRgMAv0byr47ACNtuBTfiH/IG5c6jQWcudgp3cnp8BbsRbRueUW4xN8n
Gh4aFqgE6Q1LzXySJ20F2rgZ74VTxCv82D5X+1wJzKHO2aUsuZnuXxQpBEiQU4PW
HFvpFvGLciUbrTL+I3IcmtpZDQl1l9AUO6qwdsXfxbv0Oabv24G3GoGbmamcceZE
SNFhfX11j227ycU36Y1/FTuSDPVbVqo9KTdAl5B95En0BDiK1Ci/lKAZO8otpqDV
ze5KlTs3EoCCmDTHQHze9872QZrcFnSATlhawCEeQBcsSakui74Nhz69FRBrFFEn
KcR3cHe8lPOntymhY0+ozvL6vapZXjprr1qlSWd+bOmEYxetprdJbrqicKxPokfS
PqM7KlmLZ1WKAHQoj+MJc5P1kcNTGVk7opT7LpCk2L5Nj+yuz6b4Efq88yt69BBY
bcg0PmpjDeri83kw1KXRvvVi7x1z0/m0oPlmt48WB79/WsFsvscmgF9m0KAu2Vpq
3GvUgLYa2R2v8ho3iPtiHIYOvkEwHzrLpW/T9LCx9aanGBUrlTRmlbuDvIqeiX6F
EiaBcQPccU9/0RhJFJN3GyocMuUODq1hmyl1ijtwIa6j0cqGmmAE7/w8ri6SG/DV
9SZw/+mLY/gG4m5ctJlSSB9YEQTy1syeFhzm+bejPQYynmacnKRQbyK2sqicm80Y
FI9yoNCXjYWWFfwgdMds/mVZnG2DgydCr3AySZWcyzIaCPBvhBWvV14XpjbbSDIC
HDsC9h14lxpeMfq3Jjp2Mllew19N0n81HoN52EJPoC/E20gR9vVmxV84SEd7b/Z8
EdvWMV3g4smkqTsC12U6bJnVCjpgJ5sPI7JOe83Fr7dF3wGCsnneIfunw6LuYD5z
mSGJmFTt76xn0bhWlcNoq7lxO7q3HNcq1ga1RAV9d7H4VHYoNLEp2QIQX9ffQ8GY
bz5OB9ZR8if5UA6qwGFa0xoIu/nP6+PBMbro/X255EfoL3BUYeB2+IbQ/W21n8fT
6Iah1AEqK56HUxVQkyaDbti9Jb2u0uStmfa0oiNc+pIhEGMkLn6mHRPjkEPyDJSH
GUIY6RyZpGl30cKFODrn4uOilau6zoloUjd07fu5SrJ4FzRUREmTLutAr1fmcoBr
Jr6PtmYtrGyr7HXHbd5g1aYsW1XFrpoCboJY/uvH7H5TY+Qayc7YdBNNkxdKa5GR
gIm+Ebj41FfvKqzOb63VvgHF7RN4xVHvO/n0Ul13UkiPNDSMQIeHTSzcLtVBvXvo
yIi0m7SRz63GA9xHUQltpN7Iy3D1FlFxAmZ6h0uG99H+cOOByheD12m8SjVbeEN2
OLWgNo6dzRPJfRbBhgyl3h1/DbCPZbiWbsL8g0C4e8yWgJ63Ix/THio6A4sf6Ll9
6Pl4JxGmCKM0Q2yLyumieOlo7+cLy0d6n+xKu2GTaMchGbQu7eTjmSYjf3KQTDuf
3UvweM7pAOEJjJdaFePZFO6aY92ix6/1vMXDjoYKIDTqoH7j4kJ/ooBPMg1GWL9t
PkMZ1Vr+2RBbSl3Fs5PhTmt0eDfTiCMb6CeWLzOZSKKOEPmcmn/1/ABqirAEXDe4
xp62m4IMh24IYpm+g/SNoX+lEoMNSVBxXN5iun8XK1/GoFSFBvQxFP5Nkdp9zy1Q
m45R6YJpKVIPZ+sBFzzetoeHrkLBPvpRkBWRzhCrOdupbCuqyRwhY8GWZDbmqvHD
iPMtZxAgbhWfdKPzFE6ZAXhTatbewQzypn91YzdU3ihgHmr96/yuEMtBa+i+lQnO
MXbQ0hxUgEcgR3vny9qsrdjOuo54cxZ4xoMMSMtQoSSyzdMwQdKIotNnX+yfKEF4
4aDBGX89MjTBWGEoWebKpehs+izPRBMWDC0EUmxvf0GP4O2WpLgQBSHbjabJhfE9
qfmRYVantb4wJPMlQdFskVXXbRVoHZS1Jp+62MlealQN0k3HdLLKFMVwwS4dVWkF
f+kLk8EQCXihV8FIfJ0UkzUOPP56+zVaU14aXzbXhyErNLJAB+ljbpxImIJSSwhb
i8FotszThniiizIU1UuW0VCpmdYxIGWQDkpUwdgDS8KtC73XOuXHShouIqLFcQoy
5kIv2SaM9pvWKLidKAyqSa2VHbFguIrYeb27opXFxPoaHrE7UMDXiEyCUwQ2jsH2
2fb6pQ/EShkjtAxzIGQyQJkep6CXayTUkWPfe1NbmgNFhcmrHUddrfoauoC3MJG8
C18Y7izmyfyuaMDA9m49N/oIEmH4YnQD16R2iZxPKd8FpG1QzNXqYWN7VsXAUAq4
DlQUOl7bOZqPsGbBwUk8GN2aFDlrPR5ZwG3EQau4KMztv+kTVHRVMBUjcA19JEK1
l17DW16zt1uWgTSrjCNdBdagKaWZyhR5BqfsHXMWqz7tZqqp3aHnTgH4VPB+1EDV
al/Hx1N7VJ/xWsETOxUIaZxCh+/xCs7XuZaWMdIltUIRXYovJ/x3DrjHjjVvYuJq
ccEluPT9P86nCgk+dHJ5Hr/fefOKKoQKtCdCRoC/wvSn7S0e3bmBqOEUKbdTzG9F
tHSYeVCS/isA1uv4o311g/L/YyEO6UeQW664o5O3/D9DQkablx3nUeqLqndj0SPa
PecxkAowAf06wb8IVJa/LVIfzhpTF9ljoBYFdWzsE6/R3Ol1KySxljn7gIpOAidj
FvWJ+8qyMSHK6+c1l7k/H0rdzZKv8BlQOSYBJSMBSH3bsvmWl5F0aaEHSJo4/5OS
4YzLMEvKnkHx2uh2I94w9aEIqxkFFdtdEmUJtGqVqz2Lm0yCnIB1r/QhRomIgYzD
ovsH0Escxl5hkEU8mvaIgT9U0dDb6FvAmmEDCxE40nExFH0h+dwJZIwwITO/FBtN
ZiizdPhgkv39Ok9UHvA+DuVpHeRmoQ2VAGkcNo8ER/usEd9XmjV8/iomBZ8Mb/6+
37F6INM11Xyy9DkRJpt3+4kMQ2nmnudSbUeH+vf+fYUHALRgZFd2TGcoOdvPGwo1
Y5JF9xVO7UjmP6xv09pPJC7J/Y6RTVpMoxseDmc7pV17bh14LxrDyOGUko0LIojS
hrcaODcnSrd5wY8/VbdKpOikIIui0iYrQvdt42Qgww9NRAPOfBnaTaygXRxeE/Ni
bgkzV9cqmu+qcCFS4vvJXvz8uj3Iq+MYgkP+N9kcuSSBtEK7rPC8vVwuFZV31yi3
DiJ+5CAPio771K8YUAM5vsbJTfZpokra8fnRezJEgDtmi2IGsF9Zi1GgJaUOeV1j
XqtbxsfGRn7dGpmi9dPD6ZKBhfjs6h1Dd38uw+XytZre0S8xoRB3hDh3WYyhsM9N
EZNAONIKzF+jGV/bzLgPW5EZ3GjZV9+4X1GeMfBpElql/BZvGSjNkcMkVOkZkzZI
y7vKFA/YJEEetJumxui9mNt4FYNXuZ+bldHry9Xlhkb/EJB7ymgntCVirVhTOJnR
xqBxpk6S1sXe5XSHdgzVIIfRA2igGHAcs2LBipIyLWDo3sEGEpjxsTn6EbgOruNr
8KGsWXRplNwX9WirtCS5yZWsLz/8NKgr68HLea+8TC2Oqzci0w63SeLFEV2L0Y7E
dkeNL9D6m/Rx3CB1bL9GoZCXaVwGIFlpWQ2NL4bbhYFs7nu+9Ekg3grMEpDRxzsc
+SivmtMGumJbXlJxbljJQY3U2mJGcrwEX8liplan5zBcyAQi/I3O4/Y2P4EJvnNs
5X6hCwf3uCUVjZAUXlREMznbiWrF1wE0DT+Nr2h2JEfM2r+2ghSkuHW7dG7gc31a
wD0Tm422EQqnzXoNTJBNeiLr0FN1wGef3xa7L7vGXznMFxjFt+Fb6+ElCTmAb72T
bTZXr5BeHXkmOY7hmoJfwmOUN9cYG42OU9TsmO8gCBMn25eTljsqqs9rVcLKFSop
QLx1PWemIIrMpybmQFxXRWisYopMpim56ZiHmeIHgHH3RyFSOeJstPSgd4r2lIba
PSy4rQ4rBuA91ZVEjsDq0HRG7V7NSGiIavuWqaO6Lu+uaX7zVYY1Ecv+ltm1mCmu
N9XzecpVZzVydyj2+iO3vuG64MiRmg7yvpakJn3hub019+7IKbQx/crT7fnHgSpl
OnleJvMTuMoGZs9LRMLG/4XAwm/oiyGOvjWlh7nziH/NkqvFKOeJdtgx5WN557QM
FVuKAssyeU8eh/2JKmIWLXnWF9T5ej7O8RLyUI/1GIVUaEyZX/PtInIXVxSuVp4I
DxMgU4sRvdqdO0AvuU6+aoKLI+B81XJMu95BLrANgU2Ox5Hmq0E1yy57jgMweBuK
IPlgIBdu7sOfwqtuz6Eidffy9OlDrz3Vxzd2NNBOu87EmGeYlyfo2Cnvjl/XUs5b
jhnp9OhjkUBl7NcwqA1zo5UkgOOaAxP1ezdLTyUFbJ1MgWO6u2SJ6j0TD82Qftdb
L/VjaqdbA6p6a7lbQ1kcb16H4Ahw/SkqoPd3xcLMeP/xgJBHOVQKuOQw+Tt1XebV
2Kv7luLHf+ltpR/MK9hDxlSxGlm6c1Ypkigy1Y2/+quIApy07MMJHxHY3Eg+wwiF
OrSXs5eIo5Di2AAeRhkkx03F2z+m1YlgtZGNd4XFT13BBjGNTKC+ZPJXuqiiI8H+
AMyS3uRK8Mjk7tKZqZ54TvF6RxMx3VgDc/kokePNQ78X73i/GcmSE7innCqJ8Kda
VTZRhaO7ds3JSkKmhTp9XA5mJs/FzO9umcrT5dQhgmY9iFWOHv6riqeL9siuwI2Z
RKUYdjZkAMG+MVfknuLLGiQ0SAYXbQTPoJwMomNsDSIjsS0OTZzrEORRCDFOG+tO
u9ph31u8snsIjqYUNHlWZvRGg3zYoTtlSjJ+wUMdzKoZzTxT1R7ZMbnoK+D9GiRk
P0E6en6JTjRN2J/LfPcopIOlZINUU7eXYh7OHoTKdQVqerIfLu/CTOmTisE5cCKF
NNgPJC3FA71RIvxHAMF4AfE8fw9wsxqhCRmKUi7KQEvm4CsSgLdN+xnIzt9rQQBb
Ek4/XWailwUPX9MierLYy5kGxubsfaA8OKLLYt5QgeNFnC/MPaSASFgrKQIOJOaA
oi6e5NRJwOIHScj/RfBRbyNEloRSMZgteA9aIHTD5uL65lkgvw6/jdV15/h671+s
NEdhPh+LBJFfs9dJJGmBQscjtV8472SpVBZdK6SkgupGmvdv71gAKG2drq6Df9PU
pJ31Lz9/MNDIDh87GNdxB6boO7VGhGb8Txd1cWffLtsQX7HKegG2l7KQ0dXTDqNh
NtIFydJAzTnGiLsawmxdm2QmQakf+7UGQ/CB0jf4BuH4fHpjoS8AfZ9uFIEEXPXl
BI8RXoz8AD0h/GIYC6D75/W9XMZvJNag4Ffa+UIWxqmp7b9Wv6Z+1Anu7s0Car8t
7L+biErxu4qrGRDqu/iNpWRxcqDVPNcSbnynn6l+jTK0HlwsKLgd2PwxC15iLyYI
4n2xF5vLd+4okfp/amc71RfKfVSVb1JZcxZCfYPK3qkyHir1jwncf8zKnETIbF+U
WfMmIIv5lVCv5ncO0n+FuqaQkBzp3hf53SWlZ3Bjj8R14VSVDJ66TMYfuRXTzaYp
XJjUuZUGPp7ggedAymuH0/uurCmnQGhpayqmfviHKIIh0cyUjL4kQ04ssThjm0rS
zgJ44tb1cWDD2m0vqiMK5d6Ms7SqyEQMtkSPoBjPLqZkc5MgExwG/Hvj417+pDsf
WX9PKW3NIhFJ+K7RwYdSCLGhOTgUcn/cIeCSh4041ZT2i+fNQhalr6Bwka8avo/n
1b7s1STWrjjhWwHiEni4ql6Zs5H0g5azSK2aVnOzbOmb2ZmseiZgiXp6Fk4f5oo2
HWHz7oC9+ro5eXNZ/NicZVj1fxn2GgRc9F/K35wl6oatYD7MedD0ILxX33I0H2HK
OIVhziKQngAcGqlZ1oNqwu6X97Hnl/lAMjmRBROv3KRPbdBhDfXgRJQ6J4nZtJgX
6XfiUf/K2HigppJwn20hCd2mCf+XQWl1EP0OLELnDJOOAq0JNVGO+GHqg7eHs2+g
G/A8LOc1dzmW1+qqc6y5bIbVtpnOPmI/y4Hp2YkSL8iy2ByAGz1mPl3j/p8ZhZLN
sdSO+evQJom2SPqQBM9VGoNvJpghQO0nO6eHJSScfIy09p0D6NwCjsW1lh9DW2oc
3a4jwbTo+96u2pyDEZutpBlF9CZUrPPHtIQtobfQ1aNiNIuhB86tkurcqGAyfm0l
f5yN1UezEEZBdTq0YA/lyMBClHt6gG2vkV5gAXWWC0C42qpVgy7sYvPFRTtiCS1j
zWEoIItuPcPmPcytAg3mpxhrjm4VuhbUCJOxfrkPbhzZHzvUHo6WnqmBy3vIuL4s
726bpvOo5Fqnfl4jW3zqasD5CN5Sr9j8/PSCRi0LhNSfca8epmSLXYVzUUeu2XJv
MJZ/ywKERZSJAysq7lisnwgJkDSH1qazJGBeV8+9Ku1UpHnGI/xY8EF38P8MgMBF
5QFgzWtI/+mwRbNPebqUDa0s4e7TJ162+tgK7/vMDuaID1sajkeWO5rPnbYLTwbh
oXiMdb6qFsqfPVWkX+p7pT2ym5NOihdSNVH83JXaG+GEIn9zHSCEdCi9E8rtwbnG
2rFoUxrqqehjuM6h4KKO6DjwT/owv3YFkbJ6hrOQukMXRQpATbT3k3+tH9O8MPWf
KIJj1zwVDN1igpSzwfzLzmantXZB5f8CBg2NEqJThuJI877wF3pwYfubKbDgJfhs
NsQ0A2kKVoOScihvnJYDDdEi3/snMIsLecAKOTF+UFJQBkDZsMm8UX/VUNABZaP6
RxbIxTygAq+kS2eP+UK7u58+P+Zuzxz/jDlKTiWF8MPvXvDAOhUOaII0DCrySMP7
nA/li8a1kpV8s23X2+fGwaupmxMgPd0GYWNhArOebdxB7cYmPh/WF4XUm8phf9IB
1bo4Cd/UGTYE+6hwKlv+T8gVKVbhmxAp52H1PwxGPpxlBI2MIUJIBA4oZKGJ+9QI
8YMxTjrbY/DEQMSL9+pjVhPhLr8OSAN0ZZSqWyR+CvugTX9cDFBvY5uwfsRYVDcQ
pohEFRGE/nelBcYiuqQWXcBp/nHfuFl9EjP8OkjCsPszb+NuHCXVq4wkHHwh/LVc
N+P7iCINJfHNVymEc1yW0zQsNeZK85lE49IddIJkZWMCKps7LGULDD9EdU6cj4df
t3b2z3nB61TBt8lWp9SbpsaN04+njHYnG3/w9l3stDNiaalSV+6fBEM8SmTZyj3N
IaRWsbHJvZqNtpCDaed6pQchZFLvyFjT+w8rKxtmhBc/FbLnpeZCkGgfZ2Ovw3ou
gx9uBVrFuFgzQ0sHJN40zIKaIyQIIt0T6LRJdfW/TASDMhxnZBG6yyNOmceWASX8
yXwQd+0xgEO2XBn8nUyxy5NYuAQDM9SIVOX6THpE1xNULmrRUbom4EVwrkz8/Suv
6vhb6OX51X7al1LJspfDQ2cN9/SAZ4aQKVSnr2FEcvHn44x8X1A1gg+uyOAr/f/a
6Lp+e57oz4m5rU/nZpn4y4KbmsfiRfjQ9SadzmqE2I+viKyFmtgwHILr3m0Qz2qb
/DW/1u+jemmVlyrrjyVLdiUjuQRXJxFixsP6tfWIDI3Ml+o4VNn+DdqmFacxonOG
D3R2dny+6d7eE4VdHzowcJ7qe123Bwk+V5Vq+f9NnxxlTZTntpiiQgcjdqL07Hw9
uIH4FUq2yf1vKOAbcE0jBFyXmBK1o/57tTet0lGisZMrjpRMgxAnKsbfJggU2t/P
kaWMYmfP+G6yzSY4iNzMiBp5iRSCaCw2Qw0i03WzZbT6COJYc8MMKU3zBBQfc8k3
emxodH8tLhgQ5smMfSVvIOmbICYr3zUjRuWCNsc8s60o7pdOYx0Vz/uvsKU41y1Z
NL8n3T+Tlz/Rbt1fh8RrF9OfeJ9/LCJD87Vqq9eipUb2IaW0oWi/V+omCcSorCad
L5Lh5zpZ9BT/6skC7VvNmNeYose6SKgZ/Y8Iw/o6gMUn6ZYdJO6YnWi875uB2BYo
ESd1aqjjHXYQEFaFDpwTT0wCC+NpfZOxNizRdsb0aTZ21ogXls46rDb+KA4PG4Jb
hYdJqCNJ+Y0TJhWuswQijcyeh4xso1kfqnoG5qwej5E0rB1ek6WsBUsZWsLk88WU
3FK+rMN88w3NuD2Po+6s2O2U/jfwIK5u9syJkXN5wTQ8SwfmNy9UHptSX2vrBvAj
Dgl8zHfQS63YxHSU5qEk0dHIub1zQaAhaEetDPb0+9MPmHB3ZQsNOUQV0oyOYvn4
77uxOWVtqcMWrb5PVNRZrF2srdK8ynHrfMrIMbfXRHFs2YAGQdz4CazE/pydu6g4
VYOnxVIru/eQDCPudfGsPgmHZ0vpqp6MMsypOOxo3llGbS88eNl7uGkdu+yvPk/X
m8cpQtPJIZAJQbGojcEmINBMYX02Oyiwh76zKuDZv4ousx+9DqC+qHmAneYX3q6/
APuB4YUdNmy5dL9LyV00Kuk2n4WhBDvc2W24TVpKpEYoRKIX+12n6bW4PAWm4plB
sySdZhMkP37Lk/MqMWNATwFi9NbZWWczSYfLcE8K6jAmW+UaqIB2pJxZuhG0qOlp
DifgrT0x0qKYyEtksC9ecI5Cauw/oUt1GhmIVrSCP0vjaqU+12aLfoJWCvf3HgMh
aC4YjrAG/3r/ZsN/FErO9cOxAbMffBgzNeEm7wrmKXVxipOBiW86sfhOMjC5JHXq
1mHZtJif5PYeuqa1JKoCN3AwaQyJH0MZ2B7M43ZPYZXTrRoIVeMeOJprQzo4o8uI
1GM/seD1o1R9BJWMjvW1qHAT6ERvbfYxEPHA3UEu5OENLpFUI+QQoh0MHaaUx1uN
g/0f5nofwH+teEk0TcvqWDWHW2H+3JMuA0WbGKqrQzMLMSiKROpJfIR5JFYndG6x
0hG/0AX8/g/Pe2lTW+6GNbN9HwGgY1G5Nztq/eUnbIjqfs9C/8Vnqt8oSkdjsyct
9R2I0y3lWJggWVULVrJYpt4l2Da1JnC53AEPpu7NVHKx+dxAkGwdEHlwgkWrx6d/
1N1myQ/3P+yTaCtxT8TEmqu1tk+VasiJe+HIkd2V8LoFSYTkG5qqjwteKcvND4Cg
KQd0yJP2kWJBmADauxCgHYbJj9+BJuTNgH2ThyJsWli6R3PyIhPg6vJ4PFmqEUu8
cgBp3hsGD7NmSs90Rkc2XtbDyaHJlPXz1QbuYzGdqyQi0j/UjTEtZcoUnD73OHO4
ur7l/iBJoQUmRV11cJiWveEDDL9HY8ZjaRuw3l9ba4iK18DaGPbCGmciZLVoX4+b
FdcWbr6+eHbUIZhvAv0NhLDHLMST1ImxvlwuZvT2Vb011gxNLz+GiRd8EyaWYRaL
JhlswccMegf411gST75jK8fh8ee9C87uII0kSdb0bbWIXo/VI2/4NG8JrYEdrACr
7KA1tKpCZ5IqUDZn2kVoxU9JVWQx57Tveljdl3IO1i/CklRd9D8KH8H1aZdZ33xo
2oM3GkZRnUpcy+jWKxwmXlvbqU5F02vLHHFZ/e9tdygj4OPUetcupQhxv6SLyFXe
1kFHFYyHNLa0kgoUybbIdoFw8cvJB+cC2lQtGZhD+P9uAn5zlSZVC+xlG8nkSCv3
tbT5abnxpcw5pRlZNIFCm6Lxu4uJ7hlNkaLqyY+3xQl/nXamsRsQuuDjJP0Bd++R
/udRtnQVJvuxPEhXa1xaFFab8KB5cOhcKgU/weK0uA2F5m7pgrDlocu+2CgLY4lU
0yaLG+uXAONc4NiuiT5MVtnUx9tFhFl1SNJX5gVvz1CYA4bx7F0OYQQE1WrtQG1N
4gjoWpTCDvA+s3DX/ma0D8/WeA/DnfybbabK+gHrppwim7yS/j3HA69WD/IMxTAp
K2OWNik0/98ewvk6FmjGzXGhziaY98tsIo2nWCngTqIJ2D+2EBpUy9TfGad5bGQU
PRNI454GPE1mtGt2pCQVw9T8Zist7FdMh1Dt++vq0reCrCvVZqqUDSvqt8N1dA68
pmC1BrZ2FZg0BI3NgKKObyvqgXbZSSEJfmKJDnnyK21iNSRYrFO38UIIC5L8rjER
zEqVWLdT60mc+lbFtjoFB9o5SuoXR22AlND9zSYUdyHEkOpLtQuhsKZd6M+UFezU
oRjwbhFS4JXo2IVi4AAv4Ey2Wfap/KAMvm37hrFm4y3JyRe/KTUAbK1+Dw8BqCey
RTpD13MOs+p49VfFdyZhEbFrFQKjDRnW/MQARifgL3Gp698MAohLmWYjrN3Fw6sw
10IjPW8aCC7+2AUQ06Ty6+wiVjxUd2reZKjgE9lnnnCIYzi0o6B4MraPgTRH05c5
4mDRXdb4nlNgx/AtrjpyoWCdkowUwh/CLvl8/xcWBfPXYkJHmZS3E70sKktLkrJq
XGpmcwsOTQmE5ifPtmzd1Kohd2k/zGUJIRnU5NJ7cCCOGZdHc3NXgag3cIHKZgXZ
Cp04eTWZ4YOcrof9HdQnayxz9xo3p1P63y9jq4ayVXW6GDbzZeAFsgRiHNrLua3M
+UVkZzONFsE1F6+o/Il4OJKaaPYXVDkkx+LIWEw1/SM85owYvYkNhVi1P2T1plhb
ms9T/qpYk3GFHvF7PNFe0k0kZfXp/t9zJi7oxZrvpkW7+Lr2/98HJEIYTY+Jp4Fv
Ooj3VflOiccN60/UstconP93K1yPw6fEhzfCjIpeKJkXKLA2DqaYesG77UXlB0wY
fwkUCf5mapeLxJzY3wCTNKsuF09BbDhCrj1FSezRgoUtgOWnLd/orXS0Asv132Pb
57A/VoaO3AuMNU6RvTlaXWMOHQfaVr+f/hOOBC6U431/LkA2pRLp86ri03pUL9B6
urgZwY69hAYCME4FW/I0vAed/8epc3l+2gxespspfxuLbd7d4qhVUGezHsWtKIny
8xloYw3lNKJvJaZx5NUop29ASjynm/h4Xu1PplPBlytBstraRlJgjBn9FMysQb1j
NtFHUU8VYnd67H7Tz+Zs6skUQyiu1MveKG5zqoOhrVdbcXCIyXo85I67N1wSSn5Y
vaddGlN6ijs5q0ntwlO9KOJcEWzqx36xlyszbPUjZ9DECtfrHLJVoh/nYU6ulT7y
M7BNHl8qT6RQrBHtHvsDfxAWtzOaktEHBObjyuTE5kTyYC4a2SLpjoDze22QmKeK
9tHlzEMIFcWeiDxlQ8iOK9w7GrrPOFfBOmMu77RalsVmPZ3D14mAH0x2ToZkQabX
/skPC7eP1WMiXp6AroWCwHPyUQMJYqYeRlXAjRLPzEJHq2cNeSkx+PauZYuROuB1
7/VaoWKqNmz2jO+59/kQ5s0BivP5u5Uo/Qs2QbMPgn1PVUlBgme6cs74UUdrlFA9
4ZbfnnXyurhcZRltZpEuDlv3EWNycJETz5CYwlMBCisOHS1u1OImD98vb8q/k+wx
HLkcm56GQxTsfEW5gWwy9y7SD8ycp3dIwQ6qnR3dWbLjVw/4o7YJHoPpZX0NPyrg
doK/QF1VRDuaqbTqBGknNwAUhVtxkemzo1nZgUrJIgdutJeMdyTWD3eU21BlfTEs
fGFeQWBxh+tVbFvR+PfnGDe3Rz+tOWlADXBbe9IgqRp1ToW0ajy/YiyiMhqtcZC/
O9cSJybLjqnoA+GSaBhXPO8JmXJ71R729tdpbY+2mlq4HLUZ0CQosqSO7p3B27SY
B3y1CCU5xre4T7vkMtbk+4Xgr553miNqeoqo8ONb47ibLr+C5EI+4l1woKDpc0iS
+IzPSxq6CFC5Cjrr60sr0KB35gFFaQGW+mk2RicvfIOuGWtyyIT1n0eK93auSmCy
tzGYQWVtY0KIDO0yoJRtVRnJNZVuoKw50Njg72dNJ64RPkNHoj/VMhRxCPeVapDS
csZ+m0BE6Zy69Sn90SctpbINWNM2WXpx6OQ246C3+9stxEWK6cmKsn4Fj79ayaki
aUufmLOLvblDraff0VeWjAFZdBQPy3fBc1oS9sbNrJ0YWBvMqz83wGwG6JvIybxP
cxlUdKB7MVsKt9iU86iNFLQd1cbdPgnimxjyPi1VTQhxBaL7vKICk+XbnStc/aBo
9uQPM9z88pem9LVAstuVWkWVG8Dn5QEx+vC0T+vEgOAdTpWiDtxFdOKSz/TQQWpP
sRJ2gv+1Huu1V12+8SCs2rJ3tgdlBV+HKL/xBo1tDIUN6Xllc7cEKGlon7MF52xr
MsDsoVo6Wbq9AyREMay4zVBHwmW2lml4pViFAS1aIz6lgkrBt5yVrHH/hLywIC9G
fJ6XiCFk5XgBQhr6A7FRAtjpQ2bufLpRXjAGxEFSvMbVDK3M9wfuerTcZjgXydx0
fbK8Y0aPhnvzqyCu15G4ZL1Ucih/ZwLxdLiA7NCKd48oxrkvBv0B56HYoV+MPaP7
MSTmXX8X4SolZVPQOkPuQc6gBAJV0t9tOEenqni2CLr4PtgnBS18yL3+BYTfyAGV
KrlGbFzdDndiqs8bqSl4CFoHA6PdaWJBwsjgaKsrfmAHrImClJ6D+i5qEg/N5mp6
rtjaNCCGOyFEUXFkaNkbmjcKSbvx16WI51W3uufSlFqmGlNgAjHHzCfDamsq+DsV
V/zCANDDhqAy14funkwoZnIY0BkrDDFdrYA2BtudoX2GK5sih7UFdxhjPLXrHYpJ
R1sOTPRqsyoauKP4Lp/vk/qh6r2cbavQCIBgesK1q7lM0gd63bkhrLJ1Vgs7sQ7z
N7+Yn0hg4U6v3FC3ZXtC/NFYErkJ6zeERA+bK1zZe23qCOdb5bG61RYkVymdg3zo
y+oSgfxU/JSfnqeQrPQO6dxvUaRTqVd+DQTuhDJYiHTu7wdHknYcCC2iLMYOU9Uo
Y8ekFDzM+DVYdg/wiL9w/D5HIsu596Cpz0t82re51G1kWgsC9v6ytnxnCKkRDwZ1
bj0SxZbHhoZS6zi5sbNWRFKmUyKcxZBMVJMJJfh/y1kuJGySnhmSUC2WHEzH/qmI
3+6M581hUMDCT26GXQwmIHOl2lmeSSMHsYbeeSeQleK0IVyb4Z1T88/32bGOmaF0
t23XjsyT1fHr7gPQzKamvQ60O18GrjWNZabKEXrx5wWTtzRdAxQ2dcGlj5ppNV1L
glXPYHbtLkYmlAkh8Q8VszVfiw3ZdlLwxYJ31cxUhA0xdqkm0KzEzKb7vvXXqlWV
ELAp9oUG9HkIBK1WdP+gBiGCSBhEMYHsKz67+w2t4NuWaM+Hun4NDXs9YpV34Meo
2Udi14o974ZBfr3mBILBNvwiOp1GFvZ+gpVsmdthymNdBMgzqWnY1OThYdczWFNM
QoOtF85/HmAf5/SieeLz0ap6xB9utCkY08fO9TI6BC67yOZRKi+jI+XAKpYPCj8g
q+EwqmaoaXwdjbW4jp5Pz31hMumxSZUlyZBfkdyiWModd8uJ6Ty+zDDCYfAQTvay
T2Gs8JPYk7zXBjLLnmV9ePK0vi99nswphxNF0dA1L4CEQZLSEh6gX7b22cLEyJTg
CxMkcuesO4/VB1NoBvFrFc8MCoLG0vHKL0ZGreyRXPvSNrkmNN7w07zpOg0MC31t
aynSM0nlL61jEDZ4525M6gZ1J5EO1YcIjwBNmZ3lWMTF8wTwiFozdXVXeWiGkXCi
F+vdhjDnHzUfrONEWxDzXMFHD7+YkXRPiVLhXVtxPtk3nzwgcXVThjuL0Tl5XV5M
b9ruvrrtPtReXZZ1+ADNX7D4u4bif05TXsWQ0joWGMD1mt7GtM9jOjPYI+AH2P/+
FA5vfv+/3bOR9MjacuTl0K/cz1tGD6/ggSUWgcMATpq+n3dZ9s5knxrLO/9QQ5As
W9AGLVm9WFKEx/QHRZiTTsJNwzIj77Mn6GRccQ8WuRlt9GKZcx1xcO/DAEV9OwqJ
kFGqz1fOXJTeDaL182+gtCtXsoHqNcChYh7FfNzPkGnZm0A2kmUVKDyVQ3Q8Kc7l
JSHHvo2w30F9v7DZvNszknDmR57va7aa16G3wyLSSP6MBxFSdrWT/xh8nOUcPyFA
n7/AUpryvw6KDC/v/JKHGU+LahvMVTXyroAbq4Y5sSnX/suXr4BNYPRoI7YDR3OT
AXNkVuHG9jLs4nArgNYQOj6a0Ue0cPSOFIMqG/SF1qrVnjf0kic9ca2oNWj/Y5i1
AD90uNTsDsHLgk5lnLWRCPWNaz6UQSIfBcim6WVfTjLjDjW11CvTCyy5e5AykGVQ
ExvpkUQJhgxLNXhyx31YtsSYuOOjaPQa5ziU+vqnnCqDrPFpIHdf/ZrVbyMZCf4g
50dr04EBzFMlKITEBuZDF35kngumEajWbHoiFyMdnsgJubSpvUaZDWMVFmUZMgwH
B/zeetVyTqje9G0YL7DKdZSITGWiAkUEah1zRSrakxYtdg6lLPJvvTAbxXo4kGVV
SEWsHWR7F3uFQ239xsVCyHNQ0KQi6uDCNdzRx8iYM/ttiSVJ/oPPGJGvVcdD9qQH
gwkqXBVH7DGh3e7bsk6+Y0jlD9gJ0suhhl5hOlDts+kgiw7yBnBXVnn8G+VQCoFk
F0iOAq5N8tWObKncCvPPR/uP55h3l2hUX4xUazP3Kt5EG+imDomwii1at2uFgD2r
cm/MiNJkMWA0rIeuAVaA8gj1mAdWLygLiHMHmhg++EU//eg43EZai0QSVjbuLt+Z
vi2SQ7tEVmvEgmQ4ucw71GEq21ghqvEjmwX/g4OB5xj3bMU1cHn8sGty2sxY6xM1
I02qd6fdNJG3ph2JG6/FHQJD86ihu35ALUgzbvFWiYsmlA2916z8sOk65ZkTf9gQ
QbkVAac7Mmk3qg5g82kSKIxjtPVQMS0NmJOfVfBvOMu++/mZiVMNffet+3lsEsN1
nXf1XmTDNg8CjmzHlftn8fFxLr58aXVCtjLNi/SorPKNjUluzE72N5arV8xoszb6
pHBm/JcttHunCTw6TQXdMrM96/C2fjMQqscZFisaZigVl+NhKX3Tc6ZKI2WSa6Py
7LdbtYDPA/owyaG1eh10eZOWDUM6X1Q8tKnfWdFGkbzkMKwjnVVebPfnmFBk/5gK
yz4HBwa1g256I0VNESG/LMCUkyEZ7hGb3vIAaUdWbM3bkfSAVFM9nDzpxbk/sQ31
BRUS09EGmDHkYiWcM3mYjYtTYS7TRiw7W2KFFOdr4QbnJkjRIuFSsTYfQIEGzC+X
lSDpzyJXq1Jj9A2XuXcjXoR0/umbNAfSHRgxB6S3A8Ljmp4SXvNB5j+85QcWJpQj
Vzn3S+OoL6OVDQTWxer2p8nkcDkUdsN0kPUsVaoChbxuESEzmvPurFPb+vnhxDt+
NxSvvXQeVdjjCAJinlfX5q3fq0+ueU6fyOIxExvh+guibI3Zs9sbzfdM0pqqTPqk
dvmvyicTNSf5js0CXSBNhBlLzeu+mPy0ucyPLvEToiSEVVGyb4FPtcugAE2YKdfU
05Ja6rRSua39Uch4/1xz40okqa1T58+BdeijeXRyjrNcR+Z4eqGDUT4ZW5ni1uXL
omzc+wUTAZjBREGAmL2jtmSyUCx3sSoSkLQYGONyNfodfp6wlUy55XNbxnBo+MXT
3hvwzL0vZqKdzMMMjq5p4XDpQFdi2Or2H1+4jv7hF8TOr9higQSQhIqOMvyEP2ir
7VXQd+X/2FLEMoqu8OJn94jcADTT7/JmG4zZre85wpGpS0SphUe/8/sVx8TYXVpu
17COah/jGfZVeoBDy7jqk0GEBIx+7CEH/VzzDQjR0xBWErrgo8PYDHvg1pyPWqTf
fDAaDr8iIO8hIWowiJBMwOTFehHhJGAXfbrRkFXFax2cUGzI4TcarZ6vU8bBeICQ
tZ/cgxYCT8d4+HSdhcEVfqM5UUXeYqTmeX1f6DZCfBIOwEgNk8Sxygh6d1ieti1m
X8mROxWoSBWzjXdM+aR70HJJxXvOXsguIldeIA/oLT7GH06MNZ0CpdPCtkI013Pi
RfGFw2YqaQGmkHBZBbTRDhJe35htmYn7szJ721bLxcmsYMZKDQBNifL2xJuMVoiC
XSuy21GOFLv6OhXKSWhuy8F5yRe4ivoCvCzh9e65JiQaMqNxmDEIVSWAaXgi02R7
cQmiG/YUDZ0i8kFEYzjSXwpUbqffRh48fnf8cFk40HR5l2z365CEI6rY/tyep+os
tnTwtjBLBBZU6mwCtyuhdEhlqMlxZg9Jt5qmotwK/Nb/QV8BypnqKZ04p6kZDOKX
t8qBOmSqIlLConk5M2NZ+PFE4RjfeR049hsKJ2+4FIlukw7RN6jOGZbjTlJp6uke
eNEnMunSS9W1F8NYiNvo8h8B078Br3YMJNGfkq1EmPZlnOTjlxulqTgqadEzQAUa
D9ViRBhN6ttd7s181VyrwEX2HtWmux7MO35O6YNxo1WHBvgCmUnoO7VDU5x/XDf6
W8zliiAf4uetbo13zcIzq7s1QePjZtDDOAckFGvPlH8CkR3LqXGCLgrf8dFd6/aF
KM9L2cibP+7ee6akNknu2wuU3V7vN8vAZ9Go6NgA9sFghux+XkIwqD1mY/0zc4vo
/56UI5Yzxm2cDo8fh4E1mjLg+mwOhzF1AjdHAmKPL2K3JOeTQsmWJ4RFUs8DkDGi
39d19niVCHVeBYZhBwVFaRMPIjKu6EpHSypV4AAGCcR3fx+K2ojP4uxoqw387cke
CGEIWraDEDnywlbVKRMLV+viGFZxLZOl+9xjVVmYBYg4mi2gxgkPGjxG0qeETxUD
NY/hT2Lpja8R+uhavK93YroGCHKVKyTPWPof1gLoseJ0MkbBH+bAePat5+Q7PgsD
rdQj4VwzQR9EhqcL11MD3px+bA3/trrwqvW/a/QgdHP88BpIZ2mHONp7Z83lTjbQ
iof8xQitHIlldSfsnaC2R3S2uZYzPGN8fxEzlhVae1wywte7QXb3yQkVZa1ARE3F
aChdvKPYNBL/c2ChsIAnkbh927JJCRAdlH7PhHIIfYLthVjXp2kai900Xs5PdYQm
dYL1kv5sUIULU81HmvxSNRr/Jhd/xpQTdmtM3CKMQuY6oIk6OJsi20mTkc4BRYqb
XdR8JQh1ZpMJBzhzJPMgu+iU9nKgE0foUqy6iwLZm5sIe638rwEfZwqap3aZEAOm
cRjylcP9S2/HMg6vQ3OEZOn3rmnqzUUFlzUgcVnwOIxYAfX1MAPXCJ/m3J/VcQpA
YVczQTPsQHjWI7a1CQfPd+bg9V+P2GOoc+FScwD9wgRcg7YzgfxwQf3Ab5drHK7x
wzXyMtTJg+43/kOjCnFfFR7iPKVuKn59sKhK2WLTvA6PiMaxGteS0/fslrs1VUDA
UT/hFXcPtPnB20XIlqfiASWrR8VQkM0ouzC7MBanJbg34nCAFit4tVBMJ2vxDprX
kT3JmBdtjz3s8oBMf+85YZBG0bIssdA1YyiHggDRvAA3mMGP02sOvIq503v6BKjE
YnPE3iCmyC13OpoxLaY/+YmhXzgdogLrdsl58vPOqzr8VdkWKKI04vKt4uZ9ew/D
Wj8NsO9nqfMmfGb2LrZW4heOQbetDC2yOOJ6A4WyWK9JJMn2YlCy+Hcbv3MJGxv+
o46CpfEQypVVM5vVyfaJJU44wtgag98lf47QcZAPDLXeRdYDVYhQdA6jahNrh8Ud
HV8VKga0E3hOZjKo6XSTGspjxVcJ/3nrm99lGxLRliqh6w05YRG4GMKu9CEqqZL7
bws5fCQcmEfM7MeNqlkaOy1W9xB9JEhokC+cAiHGdW8H6MzWhSJR5jr0sHQZLTL0
bJpNRk0ZOFs3PG/NsmB+w5srwvTTeYuRrIeOEYOBBzosMCczjIm29elabV3U5uAA
u7VbsXQGP2wGyIG/RvcurSow7HlOHWy6LhDI83iAJS/UDL54XNKNLLWsmiEEgNZH
e/3nKu1/0uEqj8+05kna8AxWb5xHNNBrscRiS849MS5GbGBHnOBPsF/RzcOOsmun
d49FcDlbKLEBfdudlmfHU0r1mT7VcFDzNmLDoD0bWRbP7Ad0uT6n12zUoE4Gy1b5
SA3PEglQpgz/fqxjtaFt63M7opbdwWRBqTMCjOUhSC+5kev7JvlytnDwuF+stnHz
58hTYL6xz4uXofYepIqQtvczTCCSiKa9QM4rb6J02QEFIxHk4yXo2srhnPkXDgwE
pIT6o8ikNl6FDhsBgmB/zeOgnK9SMofiVASsrxYaqp5PWIDZKtEuMj17lSfdMsCk
QiMaRGLKTYRpQoWlzl9BOyk4UTjzbOVgfT+eqtbIWDJJHWFYUZtw/Gtx+ECTejLW
yGxzA9pE3xxaC4YS1dDJ+u3kyG1UzF7F8bgdIlB8en1hCZRmzdgEyyx5j/V6QCgH
iFDNoft3yhrQ25FGL2YdEIdEkGo6L2IGItJ4se2L9NpZdx2KfIy4shD8RhMN+43y
Hl0Yk3ddgY+zvFgBp4nxaQaIxmGqsvTndRSEKqm60G1OqlX+4Jpkak5UI5Znkny/
ux3k6d6lSPurBWyR4IX72u/TkX3MzGecEUu7VL54W1uVWB78CR4jAF2cmBoAoe+D
PJDCk/qS8fp37EfO++I7edMXq+CicyqjDnclIomHW6zAcGAmGabjCKI2nSUB2f2w
ZD1SW+nyzJDf5Mmr9IioIJmZ9RypL2yKgij7y3j0KNp9wGtM6/YpIRstQ4q6DKas
MttJG78yCRrGPLCK36HLjrUbzk6AxYCtK4wLpuSdYVfazF1kTunmh1rQgXQuMgJG
z6sIS4zcWC3BRvC5rJkYP/ra+cuWi7YvKhMDcYlsinob3NBU12N6RREie2oQZyeK
3QeSNkcRcAN4L8+qpCl8lEPWdqRjo2hJaVrVXW9Lcg5Nl65Y6hEP/7RuMP414Ifu
QLe8TF8Vg7THx4vnJkz5OUMuPJGtXqN6mIkGN+/PxEB7OteMXty8LKh8fYo6P5Zd
2t1+oA6skaVJ0Yg8jffeo6prUJgBeL3C0wrtP8bSiNBr1vw8tA+2PscmBQlQ9FLe
C5OYEwlvOf0rbeMlZokr+mKBouUIN9NMxcEApt50znK7peXP4jIf3z0neZ8ypfdF
Zj98hQuklFyLjaTQB0PYZL6XkislGp0i9xkEo81iD05m5MT6TA3RcO/DzMQIFH7d
LsIICldPIcoarnXkJioVuLmRmBQeGONgOCv/Yrg41QwkeWouk+yQ442GaIurcknR
GzMcnkiZeqUW8SsZ6qC8dj2wHUi7V+Wpkt9uY1ttrRCtA7MDiUJ0OLBi0PojYu+W
Dmk0wj5Sr91z+4AfeZvDqQI1YTa/r33yuxKiMJgO9XaHaF/XInqT0kScmjtnb9pO
PPrzoG5zEqxhJFq17t9g2UhRQOLdHfrNB7+8Rc+bmk7ALs7LwUrYTPIG0CciWwKE
2kHUlUvU7aOhIMvMnp/vqWRvg8yVqGsTcXKz04Yk2gYm0TtVmJ0+/TEu3PWWJCq8
8vFEywN2jKdHwP7ll4Xa0H7znYNrktwCt1iAWsf5DQewwhsHdFt0t3ploPQJr0p6
IHFA1uBd34BmEK+QqlWTXB9IYoguDdyZ1sUgk7OB/84SBvJXiEqBzJSCEV94SP+0
ybBS7ZcBO+PprZr1Ly/cgHQd8cF5anFt5b5O5uWE9MzEHz4WGu2ayWaTRipuy45P
KW1Y24AR6/ROCczo6Yviuiw7w6tqBLYtHaxJkVoV9QCyKtZdokM4VTReeuU1ovC+
SLp+9zWZgldLbYiYOzjwvTGRvEEzzMPgZ0nRfUK+n31HFvfapLkJnT3zFbuicVpk
iK/MG5NarFG+qOCb9Y3zpylw4Hlsmb3CjP8fk05Wf6J3otxkVKwuOPTmSNXiMY4l
nKCG+jP10dfnljeMbr1rqWWwqltZikRH1zB1Q3Yta4SkB6s5yrUzSbvp99CtN7Q7
VnHcT4nfKNWKIO5xkXOu9OraFDnWwi47cl2FYA0vlItg9S+ka/PaYovUIQogaU7r
5iCnAzMcsCsMxDyqoKwnq/kHQj6FzfYZvI+OgXy55n/DV0PFm8vjOES5h+j5yKB2
t4uL62EDHnnla/dpHEoogpU70xVFrb278ntNwm7Wib27s/SEtaHkUxL54R8JFef2
7u12YjI2CkylGjPGhKZpuKugVdAQgOtR3BpiA07t4htOuoD3Zq66xNaN7EcwiqLp
gQMP7EW8PZDX5BouYXeDZAoGzIC7aUURJ8/Rdt/Gg5tfX+LO/cszQ8YGDOtXcsLc
5Ffgm/yGl74R6FLZpcFuIMyVbi/9mA0nqNdS5bb9CA3M19z+MJn0GrHux3DpVkeY
2eupUQoEYR07CkCAbxL0RJWMJLtqXUkZ2UDrK+UrWE38F4gXs5NWSGRzvz9VnfDa
uZneIOdBpI3VMD5ezphCFIPqxiYx2wXb2MLocCZaQG1HncKDZHHVCZ9t/t3I0qGT
KJp5Tx+zkBzmfrBbVTBnzvPN1MO86h/1wzR3TwxQwk4NEvmmqSldOb1ua2oyiygK
dE9ssOZU3AWAAvwfPvyUp+v4YVQe4f/vXrQuGafstMKB17ShRDPpiEMVPTIbIr/j
jNJayO15ePCLXUwfzy6AloF8JXaB6nkJZs/gCq10SwpvetM0JFMVHJOuq83IC/W5
ZDEczaMYx5gJUaY2ADWmyqPsSFltP831FwNa79Wb7/ROPsi1XQZ+H1OrKqgH6ppu
xBsOre4j1Fx4XkYLlRqyWZkEIW8n3Zh8cl6YU98cUkSU1DyqxjFDn6JHTX04uEIx
LpofxIr84xkRwXAeEAIo8lwd3c0o0d5lxTVV8U2BlmDg2iCQNNGe212KHNe9Jslt
VM4VlfO9tuGeBvfEi/67+62qHTIuwQGuwSV+eUGzvGxVWwzyK+CwC3tfHfw4j8It
97XsiIRS0AxsNsmMpN8MHZ6tcyh14vXBZ1oyT8fHunVyJ7c1d8vbd2AhImrtKTmL
44zOCwfTw/vT/05wRn+jjqNIBCWXcJ7R6f/UDL1wE901ruE2CTdzMtdiyaY4SsHw
zW2N86kCZGZyr2K84rvHbZfXaNK+3bHrl99CwxkphsScwX6A0cXXXGQ4xiZrt2y5
hP98ffJoSDDkw9N/0c4JHzgIUkw8/lJEumr2qGOzDnyGn5iw+43C4CEiAZCRCtAc
NdCRiDRCwPUvF3bb6IJPp2twMcq/x4h5bjeV5FV06kbh2fR0i0aMRevLt3btOAi0
pgVuyXCoi0X1YOzjjiLecCDcA+bMymXr6egYOKjIgwmR8uNZaGUbtfNuP5i9U/fS
EwgDNhZxEmbxp2Gp01f2hhRBRw+M2E+Lcu3dHljTq6QaD76JYVIYLsXo5nv21V8e
hO2u9jytwye8a2GJLhbBqRitPrPzPcKGnWUj+5qDnObzc78qnaGrbwSs92NpeuXq
oMHI/ul0f1buJQFAID2FPShMc1qVXggt8BIVfCAGl0Y4ARxOvHLJK6rvsG0INN4E
DIGllL0jQh8SbJv6T3e6vOElIl2SxQy8xGMTZsAOTIPEVy+aFl/iUcrpdEkgpOdm
GX3lU14ZnOAhIMxeKyElNq5+dOws+vX5iM/iasze2KyECKNWSyBLpou03evE3Rwe
cXejrKm4Ne7VpN7trnG3BUpYyS7nxlTivTRsNZJ7vBfPmYVa5pvxHGkEDzqeU/wN
LUKi4EDR0yi6TF9Qa8JHqgCOsaj5xos9PKB6vtq5aY6AKrFSkI/in3rA5v+dUKyE
omfPWEo+5dpXjjqqvIlYt1l4sYNoB7kT48hFs0zOnjhs1fRxboGGLbirXLz1HVHI
5x9DUrhlRoDLYbg06OyhlVupMwCXPh3qKkWACoaNgj8xAvdVdUs60oIn7aBnpDfw
9QPCemMWpKVIUCjXG7n58pJRgblNChVkvnWg9BDKRWXNAG8cvK3j47+y808EC0nm
opmmT0FKWsTT+xj23k39Olu5E5aeyV21sdub4c3AnhZJYXi/HecyU1hKpkI4DjiC
tLZTYLzDSSQdVUwFUATPjccOGBbKtXAH1UvRUx3aYVLKUMl9n6hXAI5bYRVrwndz
OVsC3V212fCMidlct58GJ0gsmmGmNtcsXJZgkkXEb6T74t4N9xLR4BWmZyuDb1Mf
EnZhJpeV4D06Pni8hoWzaGQk8O+9ZWdWzVOy1qlGvBY3OgU0KJq5nG5L4m5JXqyp
61eZcsOJGYpuS4zi3RJB9ESMqZZY+BlTEnQQ0xffP42EZn5wo4eMmIEwd5CmougE
jfar6n1i7C5o1rEVUyHr1x6azLNaAkSfYRUqSbDPHjvydB40CopV2wjqRj7U7FcK
dTfpwV6fs51O3FElw5rDNARCYuIqoswVqbo+xWNrEFeTF38yaK428UNNjn+PJ9T2
aJlpJH98mgvwXGzYwN6cJ1gOzLm5fgcHK4G3cPEzPuBArUAY7pmQ897g3gfwI9K7
OpUbBjmj4+bmd+hOJDdefHb3W5qLRgnVmc5tGtdJDFBzLts0YGtwlk+AOnOx+8dK
hCLMqsKlvqDcLGxXFa1Wra86iYdyfAfJwXWZtaot5W/Dhxcv0WPh6DQZHSLY55RF
PkkLRipSAVgU84hzB5apgwgjOuTI0+ind2sI77TT6gMEAb6w9eLTUtJMYVKK/1sF
fREgBSZICQoW/ppU04avetO2UMMbuR00BvPQqRBMVHm6z+Nx+JiIujg7T9daX3WG
1T1AcEhv7UxIPaZBVz+FqdlaUuFav34TlwZtAkXdQHOHqgUGzHzZPsfAUmzq2MDH
JrBtzMtQorAJnfkAVoCHMXIogN/fpWbeTtQWYz84rL+tiYiXi9jt1say2s015WL7
7fKI3O9DwZZouLCop/KSMmtmmwfKLw+bCef0xlcy5m33di//ddRxP0CaqqLTapYQ
YS3kw9IpMBb1cLaJrHvHMAxSEvdQD+v4w2HdawHu5dbHJY8gQcJLoW1VEpJm0KJ4
WdiHv7HXMLQtHGoN0WkRs91CoZy5yKLY38l2bGw8qgV3xuvP4T9luYoOwg9lMMrt
bD6g2FDDB6Z+Env7T7Ho69b+V/boQZ09+iO2RQfNBjq/norbRX/gaOKFp+j4aFnG
z7bO+DeTVRu1F/ttncRqrL2Ez+9OcYJsggpQixqj+mWtrpZ4w8q9D1g89528wiuP
Pn6q4RB25YoeRLyNyWoBcFXPNHkJCV3eUuPPt5uPsd+Mg11hmT5bAUnEcImGBhBT
0eUYayfVlTvMPESUhJmrw359TanjK/ke8ZEPVJckGURzB6lYyxUUirmKm3jycSM+
Dg2dKPSldMpSu+fLlgHDhGiG2l2k1leYCGKttlGecdHArcBw12P778SnX7JEozmI
813FAnIkwUHRvMMbHHm1gjSFb3s6gbUcbHT8W81gIehIuWwhad9xLEj0ZNJ+FbUE
bLfyU5Xz+U1q4QsJCRnWInCGFnRlRnCJP0i21Hf9sbkQ3tlrBxNDl+NbVc7A5xzj
tdsVxJR+bX+Aa7S6qDj+RZhxuhotEItrZpENj3iM/i4rIQgt54WDxYfHfR//iVsd
JoCilf49GilO8UPyu9tQw6HvBDsACgPYl2hrmbbFRlvMqrstH2PCJmh4bPpX6Djq
S1MgFECIsoqkY8Q8HcbRqlScXt+vQ4bjhdAUx8fPe2bbb1aeexEKn9SUwSDCj+iL
Ax9RxsUbYtuYU8vntO35D+OYz0H6X5iCt+JwweN1+gKscDzLOB8HmJLINYJc9jn9
THBVw+rHS1xRBWs12tw3zgRr7DYHIPi6JISR55V149lj3WvaeWcqlWvmlrAX25Wc
H92yVd4/8TWq3+2+VjcwG2/EbtYXVMs3QrMnOy/Z9FDv2C/ig7PrZddcbzrFXQt3
2myXaGFity/DqZErLVVarWsc4Uile+HC8VMFUUj8roiwSOKMfIDt5fFsPtISmaeV
ijH4f+sTMz5M4J4D66dyPsfEtwmV9egim+FdqxO2OzVgdMM4vvx4ZV+2uj9i6kQE
iPKuqUfARBf5XF9YOv5jl7aDQfOq0yiT+4bZpkihIm4MYbtvAWcQN7nv12uM6C4B
qvQNbxgC+BJDJdS69DcjrOsa785YUtC4XGkOnv0OIjsNGpN61GTD9a2eRqAHwZ94
2IabrKt8bnN2z/JtqFWWJciXXUSLYQ1e/lCBC3ASF+uxUrwUO4pZuSwszviHvlb9
wXf8dmpwQQsyWQIL4ky+euCte0doBfFIfrqbahrae6NS4WAHkZpw/rK0HnLPNS75
ZFL+rFQpFKOEIx7PF0Q2FWf6r8juGXjPVYDoAUZbWUKG7ZCar/UEzbjbOg8xS6m2
CNqxihKyxqZD6+hM59VVqPu7ptBqYbwphWgL54QD0DCvqbbxHdoq4FQQ9dbg2TsL
KgeqxC/ANTVm52YoP5egyjkzH6uAZiQ1K/oh9U4rfUYsjXbvzsoKf3YfPv3Vmsmx
oz34trY1nTNyxw72lbtTRAudA2p3PCUNRjTbqRVxd7E4g7IArF3ZEsimHyaAKfeT
X57hHx8NOz32p2PToqK4ZLfW8VZvH6/6FOpEqyZQ89oeTxygOYZ6UnGVwn5x8+D5
VnJ/7kT86g/YZ34LBzuIlv7QG9QfjmxDd/B5Tp0OSOsV3zRSizfLrY/wxijEiyAZ
9029PcDBj5tMAIBXIwWMNwjiRk4rSagPFXfHRCebYYJDNlPGjHz5+I3//kGwed5/
uWx2P7HWzXZ9dcHUUAfQoITQ7Wu9TGfQti4HXByCFsWCAySFW2tO9R6e/5DzAzvD
4UoGtfTH6tf2usRuW44cJdrhsKu0XXbewGpsE0DNlBGAtA42FjX+hPTvxzhmTuEj
TE7KQWdxSY2px+sKXN2qAlSEqJ8HmEk+tC/sPjs7qlQZ+MeoDkXa4x+mX+wNNfky
NHdCKytM7OyRKn92+2kornGeUSUCGaAbbxtbna+nKhG0FacoliYMDBvzcrqreRTs
a6AyiFoeCB/1kNwIOy4b/dkdKlZrLmQIyPYAcunayU1QbIDYW5LsBmwrV5qCTFnU
N9hb2lWEIu6wmnBJgEPWkLIOdicRRULKLLoV6CnG7OityFrX1NITZue6XH+4kxnz
mTSLFwv5cH0iIsMXS12HbfakjQpnCHMsaWnxhG93/MSdgj8JKmnegnVsuE/4uJJZ
a06FTjUVLnecdOJfkGecIKe+9sDcWSNXUvp7gthOUx5oKua8UsK2ANpOgYfbaDfQ
CYbSCwy2WcB+zRKWp52CsBzn+8ZhuYRr6kM5LXOUKt0TPVA48+cijrkt/3IWU64l
xgvyG0NG9ojjewLVg79i8qQGI85HHCK30AuObwzbJgShf+2CjSSEZDQLqRh6MPY7
V/VnM/zsnfil0V0XRsAU7gW6EFWs5hfBDZK8pu+og9P/GM4fwiMDX+nN7bimpC25
5i+ASrRsMB58UFvTqstlfMktHb3rnlPoSTAEsc85YZdkUe+7GwFdi9TGwar2izEV
SXz7q36vaJxb7JMOlxJzlc9HbQQWClxHmes+LWD4GFP2FGRXDoImDfE8eUByJjAx
K8S/yKu2etDP6glhGQBJmCZIvLU6fAzYj60X1o3dsJw1FK2l9glItjQchCT5AB+L
9JmMFEXAFgwnrcOsP7wqWOHccy8HqzRKirZWbEuT3HfHXaxoJodam9xWip7m+zjP
kyWn6pOTp/zCwATSTT2wC3NhIFYH+UuqviigrEJeUqX2n6VksZztJwPpQmIyVbLl
AuuoLWnlfYUOCsgv+OOLfST8RzLAxVxpCDX2nJRv9baIqsLhuBpiwcWi5FFqiOFt
hVS8g0fpqdOiZYSjqQAtK0HgmxDBFjYW6p4dK/aWoJv51Jz9xZLVY1m8qRXiqjbh
pdZjMcmGyNJWDd1ojky1woIU3FGyuCAN2P5b4QWqaO5yqpEbkz0JVMNMH/MIJDYo
xsn6HYzBTKlO/Ijf36hENVu8e4cHAfcgE4P8m0gVu99+ENIk9lAIswiw2dQpHzoZ
5yRk+Lgwl8Tk/sVF53vSZ2QBfi2/5dviw9uoJRH1hWD3VnugkwripNQGVQ6/7KSw
QqXKPjsoURHTtronAuGrxqfqNvVnw0qZpBq++7pZjNei552+cmsCm2lkC4uQpTVc
jykPkl9MDvhCNGx0AxtYPiK8OdOC3IUz8Hf1TGbnEjQB9geaCLopFx8S10V/csYA
ycJVD3Exg+cMW4V9Kp4AIFbw4dcGS/pirwiFenIa1JZzDwwMOmEVA49N17S5ymPj
KvQ2KVyOk4wiXNRGi1z3msg7IUNZR7TL2z+UaAVT8On5nnBazXZt9vSssos7wTei
yJM4aGuazdr+GJN4YNccC3VzHebmJMj5v5ewisTxtC9etoiN1yK0EMfDEgHidrkt
nZt7njlIZ/5HjDsc3aQOrNt1dnURsAUnZ84Gq6bPzdkf5cUCbHBPSAAg4vhYIM99
9TGWPzQvqRo5pJ7FKw66SbRv9tFTMiXiddA+4UgPCpkvvJJws3zUvFyawVSP5bFW
G1HQ78A2SHquff+Ni44iJXXc8y77A2ziWTuo/8pVAJfGh8kUi9ajEk4Mq2o8sy/s
Ajz0fMmTfHLaD+6cziVR2CnuRiWMbFqNDymsJzqjkF7ArJbvOKwtw4jXbKIlVKuP
OuYtJMZ2RBDQSX6hcSfiwDC/dE8yc8g0S4XdGgN5dIrofw+U1vPXfN2Z+SNwxtUz
0XbbVBq32lLSQFFHKdXUiOitZh6LCRCpT6Iancc9zPuwnezNHfhJw4ZQLihNYXz6
r+V3cfErUVXOC9vEqCDvhSt+0YxmN9lIAo6H9mRqdx61CJniqOx38ZRrt0/Q55FN
DEG6i1+OXMTHYPFs9DwuiPR/rcXPUjLW61q/HVWZTMFcJWQiP39XFwKatnFetdoN
8ovkaK2kuCc3zjLMhxtA/kHbGydLy0y7sMHW8jsY6DPoi19dsY6TGtsLqBJtENy2
511Jhmx7VZvNLCZ2o6k2ZTLvGz1tPfjohIii5B/KuMUPboFokK4R8C337iPuvskE
wfvN6XFjyij0hXpCzYOTGPhhsCvBb53j2pFj+YoEtRXnNwi8kAiy7X4PnWT8UjZH
cF5Is3a9H3Yee3BEHR2OfMTHhw/jZPe3quiHMKMonVv4Mb6L5CAUAoM4Jzs/2Agn
qVurA+EyFhC/EkYSiZp7lWLm6Q2nG513YLZo3xrHkrzyaGI2VpvqHayM+JLPV4bf
bc4lBN5KP9HtPV8jbhxWX0FF4U7JUFeKrRIAYa2qXzg742okvuCd0zdsDeuAR6JK
06d8iQx7GqkQUXGGZuyJZ6DbNq25R2UNXjTBGIQsVKT353T8yePGFcnpxUPSOQgT
kxgzdon8ajEShoO/YSPI/Lr4M5KjhCwsBlQ79Kp6Ha+IO/PJLdA6v6w3NrhIrmlP
8D7O8cVUqoKHj12vWLdRW/3QYOpvSUkEIG57dUnvzUGOtvPg9poviPgn0KDWF8W/
uw6UNIKROYACkN8r8gKemc5Ni8wMOKWsW1jNCS9sOXXvVeOTlCcoftEOwcOLdfkW
AznTIlwGugrZU+3FAVtM6jZDPNwgN2qHgYnfsKt2k5AgDDlvHZikwxweYBft67/+
WjG5GBHXsdV2H6U1nksyzrLp0KcnHPP3mJq9d3kT5lmwOgRBicvlEBCmz2809IeP
asjDwnCD6FwSCIie5wQ0hCs3/A1iVfwTBoEpZM6TTk3hRt0QwBpp9TrdkRnI6Vi5
B2sTEirOlFLscEqeNgBuHQM+J37e9lSmq1q3PJEw6F2h1XS0hY/N7PFaIVV/wwKV
Nse4uFL368UP89ft5kWC4jdQKtD4ts3810Jbo/lnYusuzS9GMgLB7fZQOWE2MDrz
pI9IL2gnJ3YRxckj5MP/zjFTJ+ucpjUdpfjr8eo6juolyC2HWNKh0a+ZnqLzeIeL
24XQHgumw9ikUnD3k7iVOn9UUQjcfnISRB79V6i4h133iSDaafxd4ZyRgAJNWFRx
/nLd5QtNU3l2n8YfzL6pz2h8xspJZdKkmjvEoeXIiyD/1397eE1CH+KZUsdMSeNa
i6k5rL0C+NEn0yN0sl0/oUPq7w1iQDXJaYYigJQeHwTq7hkSTS/2jriJNMSZuTeJ
gWiQF/owjthwADJDk4Z/1ex/zDPnbn2W+Sx22Z4i0XH3tHestuq7ZapHE4vhsQo5
jPRl7KDQmH9hh8P4dGicJz8alfUCJYRq6mX1qJ1SfZ5B4INYbzxfYp2SnqR682iC
LS/wVKX4gA6+4VI5H0kWw48hg7JtmC4b9LcKsiEENonrOaTC8dTCuuFxKW1FPrSj
szKJbX9BAQenZcFY8KbqcnXYpjZJL8s5fsOZmwbUAFVoZx7r5I/haFpmTFOl36zH
cuFwuUr80aclg8KPElnZDV3WZ2KgCFX9KtnA21ldM2Zf/JdeKaQzVBkecZjWyEQt
bpZ14LSzebBwI6W/LgFeUj0jnl7F10otaJO9MDvm+uiPq7doRKQlwUvilzWO9K7R
82+14gWgkWREWMmi6FxPAT2YjgDHjU2OrZgGwT9TXHucR2YUc7s9i4XOCcCo7teF
S9WdtCJ1MG2l8mQKoMMhGtcIh8AU/TpWANCgBc5RxOzMKLuDdi9FAW58fufdFdAl
KqSlJAGFcYapQzBlKnlJ16hAX8ZSatgxXZA+aXUZrl1d8NiFbKLbxNKGQ4FkqXki
NNgehUrHrLc6V5zqiQsrQo4rem/oR5o1TkqtC8cI0c6eNuUjw3beCZOmnf/i2LOJ
D4ch7tSeDZKsqSwd8inG/S22at5BZvvg/s8IdfOglZdw287wll5MvFq8zYsZuwpJ
bMEXDRAovt7kOUqGFj0y19HJRM57YsUcaR6Q+VacvlhFVo4W0uBz/phSEJmgc8Wo
7SQacLZLJEYJb0u2av2zI7Q7Mft59jKJpYJT991JLgh5JS2ta3wKug7j5goWFwfV
Jz8FOXhvr6tmeqjUHC8lZhqGDHr9dabJUcQ9O+eCgcEdQDjdBTt5UJ2Xyyii6dPW
Ft2UmNCHwV+Lo6D4C0blFl/XvECZ9sJpmjysliKvYEYaYiV0cC4juF8XlT2NlROn
kpjcQajEbNEEklXsgn10P80ccNv5VaRalueo0O5fPy26d5fgOOIIQZn9xBe3AgGC
xxD+tkwsu99kegihrMCAuvAzvkKvALn9ODmBYUFrdAfZUVYu16eMLUSYEUeOohDD
T0Tg1ZUs8KiKPMsLqCp1rmTVcbt+j1ZqkCI4CnTfyN5kBPwHrOtTP3/9xAjtQhzD
5ZAycbljudxaz9Woeh2CHYfacYMmoxzzjAqnIRjGG/4VZGvNPxTTQVPzmsE8DtnQ
S7iUScn/rhVVgbHyw1ulnJ79HJr4qtgxGvD+qhtVH2M1Y887hCFk5ullEvUuAP6H
Xj04qoOljoJxW1te171oRpApZSvZdSbCvw3B5Ho2AnskOLeBZ19ePE5Qgr0Dnlr5
M7chVsmhEDMNvXJ9otjDYKJx7VqEAbCB9hPYq9G4QAflhW+ZcX3e2Hu9jyGzm7Av
i6Chkj9hEbYQHy1HhVtRaIC268QZcdZVfmAdiwrGEB45lqXH6vCUTYs7maT6cBTN
cNCEoqs5wX1aGHpu7AlbdaxFxCvUcc8cXjvU/Zufa3oKsQy3FUF83MY5o+nl2au1
UDsOCxWor6QHwjO6CMLHh0gXSl1R83hjLzMcE/C5vDXRGp7P9bGTDcf1CbPFDDdI
ZspJBDsVZcxih/GcTIAT1lKc2u9RV6mWeNAAq96kkUOHDrPwfyC003OyVCYtbU/u
/BlHlgyQIcnr4b+ZijlB741yeT6Nj9DgHm2J1nK8LSma6QnAJBHJfJ9MKR5H5Z9m
Hfm8z9sL2EhWDN5i9jsjang0Y3Y4eKYmQ2pn3TRy+aLsBx4cQoVVXLHKA648N9Dq
OFgWXueVvITEnemDkW9N9XkST0j7fhB78Xo9+GR0/s/tQU8ica/uhxaoyL6Q0+XQ
1QmAMiMOBSdOr1+dc+F00degVvHVVu3/LbALwbfw471QLl+FhLu6+KVuakDgTGtL
PNi/FhzXm58+59PeLKybJuXvslYYBgD80V/4KAvf16HJB1t8xTvOBe+DWQGosaHL
UUZBITinA8FKaIAlvpr2MSZqUAt/fnJhNllfBtU4oQ1OoV8JFZlYihf0PqHoQm32
sxX3X65B/npN+nmaSOS2kOX3ZVjvbE1/v1s36ZjXAA7EoVxYJ+EJpAEJLQB7+r19
i8++UpMJPEtplJmNb1Iu0cH71LrahZFvhd/tMQYgev2sBMPLTI+Uj95uWFHKAho3
ivBfINwOW2oNEYTu8XRuw6b3Dcb06DhbCsipMT796W7krmiWiJia2oCHyEtyS+Vt
xLV9VmyoUp06QwYj/h2ZofkCV+SLIdpHRn6CsiiPoJ8V1NysFRgbfKJtt2geqa04
aZqMsn7TXpUdksP4+CBeClJ/YJ2QqqXFUs++R2QeWcS7FcQdKv5sOY6TLgTf91zP
9md6SWSPUaxn8CyzfJJrEXi5HYdeQOBXn+JuHMSeAoz+q9eAobX3hbneTMQqT44S
AlHnvN1AheutDg6fiiKH9o8pdyjG6hLY+DuCVYHkXzVlLEJ7Dw6zVg7rZOOJS/c9
eFk6O9zfkB22u5IgzUygvR3k+9yezcWSyT0zlTRjh9sM39JWdnrfGbTLTwILQO9n
xTfALDxHyESEWNoY6uqRN7Sk76QK0zV8/7JjU3Mi4nt15vufcZueJu1l13Wn0Vc5
u3Bx2ldSehqLXACrfCuTZlZAfn5UhzWsW3y+u6GFW0RJzQckN9mHeX+iUpubct9R
jW68qdF/tNHZrn2iaULrzsiNDLf8nnx7clZMM/Kuui5dCpvOICfNcYRtoCcxVuws
B5gEIsySuIV60kDHsbDH3Q6hA+aNjPZo3K/fSN62Yez4BOUkdrEPUQCqbwNk64dS
YfLKUJ/YKZXe5o1cFDO6GahVQRVO4K1AL4PHy9iWzQw4Zn/hj+6Pm9aGRBChvG39
oVV/5OhModEw++2EVa3685pagJcOfm9F5frRUuZgoG2ng6zWrJgFS/DLtPRrT3fs
5HXpZ9tRnzmJEpYzzAbGcWxu9Bb1UX+BXXbkoPAZmeI3XwLIGuBfrLMwMJfW3R+w
78Vs1URTBAbaM/MXQ8Tk8MU01BvItih3o4I596IVw+Qw8ZWbbdBHZblblKIQBl8r
OywDaAFVBdoYs17m2vZX+ad33qiGslhY/ubZTvZJR9MUMMgAN6CUFw/zlS8/am6q
mFfjNu5bg1KAd2qn2oolpTSFXq6TXuem2venuxcSEnHtgfq6PHCwNEJkJ2KOQTzf
F0BXqX9cJmmTvevWhdIi3mgF4ZdAuMliUBMxN82QF9Jl0NhQZVnMryZnb70DK2Bc
kFqGJut+vRqU5OOv7kDRmSuko+BKVcOICTFRQrvHRuukbCxO+hear2caxRTlAMA3
iYlbs0GkStoQrpu4xBYwltpgTuHk5sO6eFfPD8Fkjef0YWjLrNj6URk/n1ZkNnrw
6wtF1z9TUnhBh2Zueg0Du/8G8BgRqhf4b1v3sY+Bv2znk52Eyorhm/bGpvx28SQh
w6TZdDm7S71GTIbu2C0RmN6W9KtDV5eF9FYL9ykKlVnJqM28U6yefV9hP1Pbw7lt
HMlaIvnTt184V95LiYZRqqWOjqOljs7PtLdZMJx+c/MIRilU987ZkMCocsUf46iQ
5A2N8Fwtr8pbLpDRvPalXVK7Qg7Y+jNPvxORITKLME2eTEhiXgeGx3DkEVG0R14s
bhxUzKPrVU9YjMpJrcv+gr6ar4mk2oRb3dqnfYuXy3BGfUsyNPgRFnc2XRBSsa2a
ME7G3zmstAfLIF7OrI65Ohf2atI7vLgwP8CmTVlV7SpmmhIxtCXrThE1PEs98mTj
4LipOIqX7nCY++zd9wGO0HwEN3YvX+OAc2A+EqE4W+SYzegMfNnGudRA142zrCk1
mnTfsJ+wErt9v++0WQA7iNn35zmv9JZu2uq+KAT577plNcFhixpLD/AZPa8M3hoJ
kA3l9+tB1dsOuhxqfZIMdXQHYqaSyG9gvtzh1xJ9EFESA5hMSPSeSryjGGoUun0F
x78/lhfCCxIuL77MGa0+aiOGgay/lV0JFHtKmObNYsmyqqFWo+ERP2Yr6vwZJVON
L+0ItBMq1iodNkkqu1Q5FgcT103pUIzLCzbkOnrXo0GWckF9gnXg1Nt9407HU63P
ym500GyD4tdSn1EHoEFtEMuc0gcaxGapR12ZZOgRFW1B0AimJqb+SBFmm8KerBHb
IR/Jz5DAKG9+W/fcWt8Mjx8Y8GnmlUw7JZpvMcjxuBS95dt828B5t3M5gIY/MRy6
SX+XMSMHEh+fJ4GYKvx+XrFURp4q+R3lgi81UDRs3nfuwD1JN/OZ6CuZnYuxdN3t
WXVd/qLUIKLviXlIsrE6vISqbN+heyzAKPd/+O+Qjq6Nq2AHT2iHriBZRek/2i0l
Vy2hQLlnx4kMbwr9vRkXZA73QqIKm9eREnxNWaEnpCuNkAUPNK1dOn2bxxzCWlRf
jtgTZIu4g+b2kSlcDTHiETv4fvpCI1UdU55QitQbKxpNioeuNN9hk5F93/ZO2Vs5
DbgxV+5HudMV7NOosayxuIisySpMfeQ45ua+eKMfId2BOAHHhH88ZfTxPGHpuXce
EbVfoQhqVsouhg1dCbtumUhGH+pInil/t9wFCfQmWETVYh+LWAOWPOdAP5W0gcoA
syIsxhknGi8UNs0XD87onyLf1Y3S7tM0YoheMupC/6TDhLuGuHIFl5uznW/tolCb
3wmNpyqM5jcGWaGWk1E8lM7Djl4K3muVwxPE+IaZDeRamvDb/1VnYxomlCATFIiI
RsaCD+d6QxEasxW53pZlk6gqZ9V1CmHi/60f07phjYM+lW/VS8Xu5OCYbwuC91+M
p7vSxy343vzOeD2bKmigrp4gIMOURjy/+VDlpNI4kFw53cnfL7KTLXAMYGpgcUjW
H6HvI1B0/WSpQJ7R1/ygEEQ4zCQkMGTSvXGoWWr2bvjmu7z9KIvhD6JGXIGL+eIp
ON286zVUgIcwtQZA7UMEvczhwsCpbM72aL8lFD4C079AagQLzoxy1+EDxIvZw1IJ
x1RmSlSjj8TSS7bgET073Jha/Lex0MXZFTjxH0BHy1PG4u4mlnzE+xlXlYBBnPwn
+WwjH0Jpi5zcoO6XR4cmhBvht893fZZ+VSdGUGBnkVZ03S1rIYxmw2tfuwhI1cGb
ZNOoCJ1JbW7FmRFHupfP99UnU32rEktpp2+8YL2F0W85cEtDlja0NKtsu84T7GyL
9RuHREaTNz3vOUqGZh4iggX4MBpMguNj2bEEUINkvJop4LhAc5GyyUHOKJNAq92U
IxbQ94WKQUdrv5gZa22TXxme15HOEI+omi5tZGvyMba+oQSjeDXed98DwvV2F7bq
Hlk+xkPTSIHIpCV1zzQrov0Yi6m9arEubEun6yxu9jJlr3naG+/ALLQ2+apFU73K
8rGvWY+35eoJ+jkxFCDX03EKW2UuauSivrKu/Vxl7+WeSHQUG4GQKYiLNxrvVPUD
mA8muGkm7INr4OIOrsWtpqSAUTL3O9iC/iY0aUDmMN/8a69o4N1V/iZf5n5Or7rm
FFa0iF4CGrAZTGPE1WS+fCFlMfkl9io1+NRn5fWWkU6eIZqUkHX0kMymFBf4uYb0
0cds/27b8Bv3v//APbkrt3pWJgsnNU+spmIsyJMflLf1g872DP1srzZJzpsQiMZw
XBeTyle8iosX0xA3nWtt3MYWIrhnR9qCYiA27nQd117mMNAY4AOD8qDepxb5D7WO
fdZk5j5RJvIieEvTfx641rPeejtZWpKScwyH0zsFKDB5gpCQcUl2GYG8LQrURY9R
GrDGftGicGyx/cZRnTQqBxCmW3W8RtPXTAnV2NMa6ymK3K+d83ayHyezJWHxwU/Z
GrnN48zx++bccbJkgASxp8XVAlmgw23k0HvJ3Jc1fkS3HC2bILfgtUTRajkULTlL
kqHmJCN7M8eoC6aQbmb86vJLG3Fv85fyoGzM+1bbViaUVnMIaYxXBXtBE2e2qLXq
twVEUXBL2zGLWv2SS0fxibnEc+g8NmTU82lmB4XmsoPbqu5jRZ+d18LT50byfKVx
IC9WYRjPlPfgOs/lxfbLIkH62EiRfthaemllFKd9L2X0NqcCxX+uzHW2ZRg0t8cK
ShrdLVv45IXUNJYbFrBofiHlOWAMaWzqkEojtxndaJtg2PfJi2DNj77tDWUai68h
sv0g6Dj5XWDXDLu6MgRxHH2LYvRfkA6MK4sH+RGv2etETPhtw5NI6FdxbtFAzcXi
retQUANJgp+2SOK3Fx7Eppk/GGTKvnzv8gz0BKfpfsQO98+u+KFyz42sxrBqgXmK
jCj9I3UcDPkyWU7FflT9zMvA3zoluhshOKRy5bWeI63GkO8LaX70In9zdtduWAmG
JiwPcD0tK/MKjAz763FLepM42e9n8CyWpKndhy+v8ETFxfpGlarGqqB6Twzg8Kpk
BW3jC9LlhUUO7xXvrwCgHl5BYvW1K6QFi6k4IqU2MNhXhGk7AbfhZHPS7J4U5UBm
yqWLdHAjm1mysvESuSTjiZS+2Bvps9N7yhQH+XfJBThc/E2TpVx68YJhCqXJx4Ti
6LOKMAnsjCGzvUO4P8TUIMBfFaLXE0Puwpsu4tYX39GvidfjX4zelYXu3MOEYwZK
dmfVmCDVeBdmnN8XP7qR0QI9nSpPrZlwyCYGTlmRMA4o5X47PsYv/jNkeSbhZ1Wb
32cx4g4xQpYT90aC+It1+hckSgVHuVn1+2FpPDChgsCMpWkxpRBDkOpISf211ts3
l5QpmyPNVB7C8yjmhG+dNjidd4WIJCPgNh9HHNR7G3YPLvd7hA5X83hexe0721De
YwHDtZF9YyZtZU1SekBnpnu3D63A/RhsDDwNLLkRxHAXJck7DOB9NsNGjs1H112C
QngPtcjIraWka1fl/i8iHTkwIG96FNKlxJ2zZccK7uuHxzOFkU+ZxLZNuEyQWkn9
y6Z5IxCOVh8JjLbB7MvqeZ9cmR4GEGJX8UrkbOcQCYJDFnZgNgZSkek3VHK0dr1f
y+RaVK2k7VN8hraXTfmFdNlC7eKagu1jrHBp0sEHPH2prc9QwiISBMv0+F4nrz4p
dEWD4Lgt+T3SymWSiu2wt3xnycA2Br1zqqvXtC0BadwdYbVtzBm8pNf9bluxRfVG
YPo1PiTvWU8klbh+PEMU2OYAebzP7lG36J3neMKX9eVTWM4eFuTrYOMj/KfgnDNc
J3JvYaZGe9yhn4BXokf/rrFjN2mKFhiRZPm/jeyuRe5CudvJkAhCYYlxeIMDUpt6
E72BsPvfaRSbv5nk30gVoJVoKzzk81yGBLwLuPiufKIzc2+zgw9g62LnYCjb8iEU
jjzwe/zYEMkJYX3LjSu73BckZRpR0Zge17Kbsnm1sMxnUiw0Xlv3V3jWaAoVi3Ky
dSLLs1fMxvEf9zwgaMXsKttQjIC3+JFaENcx/A0QsLZ1ztPm01NEpqO9k2HfqndS
aja+eij2SWlGtN3AyHTApuiNqaA09q7b63QnAhqzfvHGsv3bCMtkp4noWS6vSfKz
DyYfDHEWjDJxazSybP10xdmfXHI5ZQIjxHg/5aMonOMBtsxKXXi984mfKY4pjL70
5chwjcqZiYNf4SuXrExEYO2fD2EoL1fmEnwo4OArzzMIgQkmuvmf89pZSbmzKFCk
3ukX3JyeWKNA7mRndpONa8MBm03EnPWFAKO8goWFSV5siPzkJSrL7HulYFWT3MqD
QY03F8VAkQOtk/OsiMATLEIcbJlQqD3xD4MtHMjBrzi9/6mav0e0Wug1mYwOUzLG
3t00KwULSIFZ7ApS7RYXR05htkiZHu0AKyANdCo9pdIXQYpYhpaRM66gBVMGy84z
LBEvrb1ySIyZI4bOa+fod5gxL0sFn+Qc5NcR/N5vhx/uSn6bCxbBzfrwUbVqu0gO
M1yh61ZD8j4c0lhyR85NXmNQ/K7sheXLUO/s72JDjXBh+V+lmWPT5+vuKU5SCNUH
b7PjPf5G1lNI8H1OfxmtDPI3xHe5gIKh6t1e3eMnB4+3SL/hw1zaPwNucQU6Ypw9
FQ/uxD0vkR7p5AcxEPcP2KdPmZ3RY3lQuUmrQoMvxi2AuEo718MIDvOdGknmmqxL
oWz98+KNYtQ+QB1wp9NUxNIoQSA9Y2PDGgQrjaHy/DwK4SrKqdQDA5u/3dFxTuoI
lnBPCJBf7NynwXuED1+eRFNue27zDzpcaeuWSuJ2i0oCiyL54U3w2cmKMtALnydW
zBGKjwv/cwh4FAMO7LMR2dY15wlTYzbabzoojYH3F6f8OlpJbP7QKp+Qfb2TjOsQ
g3QQ4yzvpcgQpiTDDeYZ9zzYt5SKrRv7rw/1zewz+iqluns5uceI2XTv0KhlaRAS
NQFKy1OcLqT1Xzuv439gLsLxXHXZxepyKhV0jSwJJIJK9BQ9yk5IC53noSNPIuQV
Bc9iK/C2R1N0D4tZ+MFXbcHGM9l7BFYm9LnqxRvvjitwOj3zGY8JHgv3zllNB7YW
MeoK8wvVovFtXqrzB2eYEGzexYLftGy458kMQO2EoUEcbntAuFJxO9U3kkfJIo6w
Skwd/wPNDIyqgmUGgsecQ4XtL+eBMaa6kA97MdXnoS+5Vgfl4i5lf3RZi7bGXtD2
9FtuUvnkcQRXY5bSKB4O9vJh0PG82msFtKbaMxtKT5n9Ql4Az8YnX8ySp0CMwt1N
Vb84JZeqhPAftNlrmwv6plbzn0ugctIg3AobanPP40Ia93AR5qfRpJIgThZCmiWX
nTZt4442sTinugCiu5fQ+OmUWv6gDUTFqOGGzaILEf8nos/bp6E623qBClD1M9Uz
rl7t6bYV+FSRYuaN7GYJJpVkKv/jbQs9z+tet5oaVP/n4ln12CSQSMBevNnKpxrH
UbkeHYsCJaK/GuYVLxwQoNCmjT2VsBqNE0vzW+Zu5PQm/roIUeWfsmHyBvEgVume
UB1O36HRC8Y/Nrz5K2OWv9kqCxW+X2r5yVxuX7iI8ro/f2IkABYO/7tvtmD2vFTE
AfaZYwGIz5YXQNdh4cbkxbCSkPjnCfwh3/qtiisKBOsCIGx4EEYw+VuYbRgRn8f0
KC6P7St0Zr/ylxoarTvLFNIBZIIeXMTtql/2+V9Ajlj7gBuAiVMmcy5FXJShqsE3
DNBvykb7whVKcFQDR50X8z/b5zViPxNFmLftyxa5HuSqWtnRmHtUYGeJ9wv7VbqS
Pa+D5eQNx0VOa2gFaKTrF2CUrPjbkIUiQZXPE0pnD6/aCua5hMJd47yEbIqEtmCa
/wSHdsdYgt/YQb+OO6KLZj4InND5zc8ViBsD2iKTSy/Z31Jr2dFcJOqW8YDemFP3
b/T5R6zB1iqQEjDYggLST54htu6n0g5puS7d3+1CCgQa7kIPy4Bjlc/UKrXz7V8e
r9DpzvCzFMdIsHz1aVwFIb+CxqKIkJ1JnOY6au9X987fx5QMT1t1VJJgIeyiDEmA
Gq7lwqKAjmk+BJdDNs8K6vUxcgszO/FcPKTYjO/alk1hRNQwaoxFwRsGmMPbPc8a
ij2W19s3GwIMiZ045vA2VaVlmYGZpa8oUxMnIuyDloRrqlo2KdGnFyAmECvvN+Ak
cMAGqkdhQ+QhZrvCNouuIfPOqjkaFAy/JEKPQ6CU2aDtG1KsM4P1diPdpkelEafp
PeahAjqZ4NAgkOUZVxs45zjHJZiGENmoY4oxVF9sqN9KLnOFzE1Ak9UrMHlCLDVp
tlo8CLi6sSKIl2gGN9yedVDbu0OfHKvHGVy2oAYqEOHj9GOheoh0XW0nWCyYq11z
VdsaRcNXpXresW0zxDi4AMisvXwGhGE2YJ668AC8Hswm9x91scX7jZNntegB7ivb
I+VX8oxtu4DzgEO8r1kdaNAVPrkytzo1BTC7iV0ZTbJdfEaFF9+aScqsRN1ZZF7a
IR4HbEKILIaqmjmyGcJ4aRjgm73u2pP4to5QGbes7vXg00SqJtfgRGnYGKbOwqzW
FPG2Dn70019oh9Y0SiOxnWdqwlMkE/dUqx9sDaomLELnhf8gohjdzBBYDT3vivMQ
6u7KuDSRY1C+xSdSRVLONDX7Xm0xxJTkvs5Wk7yqg/mYmr8Bk6wUFFqF6OSfLPtc
T/MM6YqGJearAp2uThTVcKJ9yB+Ku9azHl20bkAJv+rqe45vFAurGghCsf+k3bKu
64YHcFJzlGL7X+0niUkTbHU0YZv17RFEULgT6VSP8TTHrAlSj2G/FR0/wDzGJyUV
dYAjTgL5JS9afpRMRDnKHQQVIBbHr9UJcGw6mZF8skwpOFuOEq8LiRi5yeJ2lHIh
IYmMW0TcnlpxIP0Z6ry42Yd5t9521TidOQD77zSIOVUvwTo4kx8CTfjtY9Vk5CyC
Px0w4tpAispitwwSial22ipp63nOm99dSFGJco8dGv+iwCZPn4RZb/CggUPksXY9
QJpKTV07oPG6qVvPCZkkkBh4joox6am29RfZnQ/4R4Yz34PIMA9d1yU0P+PfgNOT
kzH0h/CfNtFqDNW/Y+WyV3pU5t3iqHa5Gm89l2mvuqvv7VVG/0+T9i0n4efoNM8I
yxBzOIz7lhIZZNXejDXIzd8GMfXmDGJyjXfaLseGT1oD02QQSazKb7xwmJjQUSnW
aiS2w4ol5EV3eofmY7gMZf2qPGkyzIbuNAK/+sJoU3uJcDoEfpMRyCmUI1J+tQwe
98m4AcQDig4p8cRAYtCQviGkzDC8O2SxdT/FIIayipHVzdvzmp5IEQSb/vaXy5DZ
yiCWVhz5VtyUNyMo4c2tMuzChlyEN0MJcQeEsT+ZFXpx3pcCmU0MDJ9qn7vmCYUD
iAYoU00NfWnbmjHu9fjL0l2L/HLzESbGR+jWm9bxekYrsOlIY32kPLKFyLSPtiy0
zD4Ds+4oBVfRNp6rta5yInKfnkEmhl0pe1XAALfGTJOMsAlAkIRrVNU13TdKZ3aW
Hg9F9XYuLOlIKsY4Fk6n5dY3ltGKkKS3DGfbYp3rsNkOhEa26xHb1JrvUi+U046T
cL4//dj+JxUt2uroHisPQugD7jHLFtuhvmbfQGXzEDiqvIzuxWXHilxTGrM2Yra7
kcOdiFRPjJZKqbNOfNrAdviXuiKj8ljbVG+emo1rO4Hy4IjUbZNF50m4/PG0J8qt
/ZIVJw2425iMnowxUsQ5O3RaIVWlUQzYGf51j0YfMK4QboERNJXnNO32AN2m/Uuw
1Ajnm+xEHNfTwBHZrcIRdLQwy+sLUIv3/vCw8Sz5N10og/gUTUEi+TC8Zki/exZm
fLqDlYJDgYy5BXmjyjYu07VYLpRyOZNlApdgEPGaa5aYVRmmIh1t7NMy7Z4D+kfi
Up1NxFlC8u47rz/PbEr5noIE5vJZgLg3EzxdOYBanE36Ko2ofNEJeEJMOJpE5bWZ
xrVJNKxFlQl0+pj36xNY6f+8oYGA5g02gap5tw1qsIYdYXkNOnG9oDpcuV+sRwrh
86wVZi5+X+mS9IPvWJKOZUuzQVJy/DUy/cU/Bqt3+C0zrAjVqm2RxE5TKRwS+B8z
TWQZ+e7pbzuFHClvaiEiYz8zjBq/quIpd9bimoZvonWSN8QIb1/Q6l/IZn5EYjT4
EEWOElaJ3slTalKTneSndWJ0ZcNac8OX7zgfTe2L8G7nBj1olMdkDaTDckANZAgy
cp++o/Lkgp0JtbkxF0Qcc+2Hfrkm8jCCzu6lqxzfRx+b725C7m0lZieSsI0VVhkf
5ETm5n0ZwvB6Rt3XYWjFmGKKvcx4E4kp3MnNoIcTxAKR2+X2Ox2BKZPCmBmgiDYm
/zsb76qS39BvvPsDBgFOPfqVhN6SRpABKJV/Los+1P87rEVbe1GFoF07Na1g/r/E
xW9/cH6AeQZjdY7lsyJmF2DcbCwutJBM95qz4/GhcASsQuAA0q2TCXylKbLNlUpL
h2ZybPibqgHM90GpEKbA9J1Qs0DQJ0z7YV7wm6zqsU6vJ+0L/wJf7IhqyoEdjRAy
HC/AsIrqWcWMBrr0jiNP3cqf3K4NL2MgkijuNCA2fRqooshATr9pYJ1eNsA/ZBoQ
tORt3spFDowpHbKpx5VD7ucZoMKHjtr3c1SRjaUy45dlvc5ojcDY9vsTlK1DgJQ3
88rIOzJAxabFkZIuuU8uWoTI8v09QjI0o4VTWBAj4axuxA6Y887YJf+S7Km8A0JN
gOubHzpYNoO8hwHoR08C73XAe6IIrkPQnVXTxbagP+mpH5gEEi6eHiPML1rVzgzm
wqJz9iQxddwPoSwBZfI1LzROvfWB41ERw1OuIjQAmHyXC8L8wWhqPcbDMWjcOFca
r7Q/8sG1b8Ka2dwnU+1dLuz3eURwoXTsBBgghh6m6W/qMKsLXRtIf8mZWUkZCQs7
Z568ASpgAoQkSZwT5X/e6nPuXCdqKhibFeBBlppbEACFhNe47HNz2GTWBH4s5PVX
tcI6s+Pd4Mp+BqF9ZE5k8/TokMzA7hPOGmxxxOo8YmYoygD48LRR6ovM3gIL9hQf
fZ25jbJYaU6gQsj9T0TJwroLAYDAf5SsapyQpUW0reKeO0SFJ7RvtQ8CNfu71S0+
jzt5AQqnKKrQgHTorVjG0Ia1H3hklVUj5jQ66k/K2NFpCVY9pHdZILiQmyoUCFlv
RDi1NrCwGUchZtSUqttFwJEW0lMVEEQvn1JNB5zIQCicBGrNw+WXVLhqpiDNec8x
I44BmR/Auu6xd8wPCDR6XW17PdtQduUtXJokNoiv7dPnA9bp/YiRWNk9iZ7K3j7z
/+CmmZhMSQDB7PrpzocdpJagSO5MGa7SWVM1eRqrC0K6Gts5E1crIaOlCXvOzY0p
K060f88yhJFUFJsY5MHiZ6VHNlcsYyN5HZjuQ7SvMP6/Ixv4sEVVrMl+yqgUmwl0
bmNZKTsZAbavEmy+qaVYSgpWSnIQXe9wcTO/+ftn1pyr8r53Al7wVMmughUbPKQP
KKAdPmHiEz5Y0PMDbEishzDDI9z5bAkzL2a2IRQmJKpYul4Z1DPW95CTT9VM8+KD
Kn7eh5I7GKpVjV2nAVcY+TX+XB2GS2LSxurCBj2GJdZ86Ak8NMLKl2IaGuSR04A3
gjYymkw4ZhaGs/OY5EOXKexZpV361RJTAWjSlEju3FqdPcccNb0FhSdnskabf2eH
/IMuzFC4CDpVYtbQlB/0lzpd/9eKYEU2AJgUreC76cuFJummeuMR2P/f2T44gp++
S+zF/HjJ4DwzUMXX0zi04S6UsmcdgJVAUx1gdZcvYGSZCR7fbw/YSI1ajLKyf2rU
AzM6CEzXFwZHn0nyi1Y3xpVoTftHU28zDISPtTB3paj3v8WQPMa/Fwb0SvxeNVgA
c94YKRfKPGiX6UGgJLshYZ6pJfCApLSH1T1qD/8ia+Ahi115LMY1hQ8NLpwzNNBo
f9hDaODMCWT3+G5AtW6jqDt8ZVtzJNcYboQ2Tl4AltOT06nyOpdJDsiOkzy8posj
ESPcTQF6Kkqb1ukZEOcopPxPS8k/f8IgoWaYq8tHkOY2eG0x8oC9A862lyvo9G4r
sR27hCzGidKYeAjDoP19nxu4nkc+lBNGz3K/1Vj+HyBZETN6Lsz6xqrFEf55HE5P
O5ccQ4EjTSatH2Qy2+vXAAZbtg9Wx/Ml0IS/DlizYHHZv5P6aUprVGovkRJzYMfS
+cofIMVBOJnVwm12bVGQQg7tlUC4zWK9EXX50/LCsBCDuOujSov/CUw42AKiD7Li
gX8pTa3HDhmABbFCBFOam2i2BML6C26s/jp34fmx/HbJTRs5iDBdsVPzB3WpDt5x
F2HeMoqFeWcsmuzqvaelJF4axVXtLfXvs3bDyWaxm5f4Go8T8fY3GrEFtNd04tx/
9DyMyVi5KMRAfpEytugnAq3wOTM7UjWGjq5vxAI2sfzuNnRvtoWgKUGS1j1FaJ43
zPGCCv0fh1esMOjAtJvdy3g07j3xbgdacjTy7SPsbtMGgMI132a8gEqdkqzEJRdt
GPzRBQDhxIMB0o5U6mOPks6f0T5EWFBr+i7504K3fgR3o2Cg5LGcldGtijpoXoR+
h7jxcrxgByWEsyrmSKdC/ZnfQOEP1PgVFCQBzawg89aad/b5EUUqozLnnideRpRd
ediYBb214u83Q5HhLQdEVjyTglGXU3fU/L+xy0by8oSuVWiSJW9CS6Bf39gPo43U
CZH0y46S2TRdCJteW8iPddwEKzIA7bpiYJ0KkFH6ed1xgZShSED+uT6VkWwCEDmD
QXil+YL4BLkt3Xm1U4oKGQ4igLJswKUW4F1uRei+pX7RXYIVmDRgexS+Xf1HMby+
TotRxTqdv4enjTUK+0QPLfCBQfNBUyJvIRACd38VYtY8J9M3R3duzXF0O17yFzud
bTX1FSpj5fsCmzJFJpmrCWtaoBwFihbGrCLBVp1fck0ZRL0PjkaUpyqhPANUzPXy
Zbi76YRh584HfrsWgcd/qE7G/ljqb5vmra/OX/+49sReof+vK279JFNtqIk1ywq3
aAKnm0pfOovsRzDDQ5LoXyMOkYjAekeL8kb/oEQeiI5E6xtTE/D2BIe1/Z5OZING
alXiWIfOu5lFE8gd0SjlbfZdcOEdEbx1grQHGj4EaYLg238hofEv7rQc6rojgvvr
i578sb6ZoaoeD5tLUgmw/+91qfebLJ7svK0q3EIim60GX1+mRX0aHlqIoq3FeHw5
+iO5t4wjqCX96Qqp/dHxZ+IpMmyfGerPOVwfM+RgiWVdxgu4odl766i2iRH8xEOX
dNAwGKJtKFQ9obuqiZv8VCB+Q5w9JNC5DPetuunn+kQ0pPBOplhi1TpHUAbgAqi1
V327Ir3X7CvlcWcED+XEpbjkv3RCrc10FayHPYeOaQr5hutx2KIvD83jJ05KNWVq
VOGQp1miK4vyYsi5AioYiCPhhMm2E+YWFXMEWK74hT5juq6uAJgyNAPxo6h4AyHc
pFhvXKvSOdvMYMJX1Zq6VvS/VAPsVCNkuDyCYunMg3YLpZDA7O1iFvl17JvJTrfM
TZ6V9aVc4AQR0S/hiL8q+tk/7BEpg4RsE1guo3mUihKU9nH+wuc6k8n1UNvMz6WA
qkvPFgmAIZ9PXo+lZKP0Cm44zv+YAtT60F4E97e8EXRYofMSeFwsLohgy9I4tasT
zyl5Jcp32HV/8J7+yMc7dhKrXqltXNDmpGxDmt0KOGUYSN4a3DbmXLrfMEPBbkVV
WYQIQsUeVOPzhb24LfsNBiQ9vUZGckx/d5EnkJ6cqqAqBAMnyIH2ZA/hYsJ3bhs5
NpnWAW2yOitq4rk4uoZfa5oC96wfYyErwbpOsKHep6dExxSwZBQVlvNdE8wMwI9N
adVPZvQp3lx1zN55ws7IaZxVx9JwbD8KCwZVxYlZGZjkFZeEdpiUbOkia3ZSpSpr
ttXCPWFH7/Lx6uSue9CDobKq0lNlr3VX68gJe+7ilPTJvi+SgKvE9bocV8Je+ZoG
pNzi2M+YtWidUkNDXUWxhyPAych67+wVLR1z2O9qxFOt/GHYqDglXQ3sn8Rct+ia
yxtunSNgRk/9isQLuejZKdtQbGavICX9HaecAkC4H/+Q/d7CTPGOZ27jFhbdV407
dmSPF1ZEp7u2Ymx90pmCA7Up4a6QmfC2eSBp9WpyzY1ai1eRV+TBu/zPyoz4IYIX
5FUUwi9dx3YfV8HDZTrvpcauOQY4KCATTHi+3FrDQB/VzgQCY25ZkrNlAnv5ZPzc
LbvSpKPj0t8AVDZvkWEDC89QIPYAH3AMemU2jJVN/a+eBsP0AXGhno5dzJNOsLph
sVJReEmF3KVh5wRjNSylYdOeju09cLD7afiiGaAKybnf1Gnr0BID5EpE531CSZqZ
rf2z+QCZ8/I5fL/iayzOhoIQjMkifKCuxEvwMAuyK1NY+GVfL7Dyt6Tz3Mj2qUpB
gPz0FxZXBcY7A8awD08Nj0yH0Vno9fWKtCLgCc65qxT0M6RdbaXUn5C4Dp0uyH6G
Dr6RxnjoTkBVuXz6jnW0Xw1NzpgK9JYn60nBcHgiUhXlQ0/W7M02xpjP3mQSktWq
u6ExhPONx6Pj0lQcaidElrAeRlUqF+CX502GA2WPjZGoS99SOu9FKGfkrh6bQcNa
uWpUbey1b2v9tWqW11Ws22Oqk9TlEM8CeTMWBBNx5+CwdLgyGA4mgNyfb8QpOn/4
F+qFh6etrlmlLgjk7WNpPmQXazbxgzryxzKTDWAc7o3A1BQNg2KeYAa5eB4GeSWa
8AQgjaJq84/dKf/yzjr90AiqCc3DKrPvrkeW2qmBQk+P0aWHqyine3gd377Stkzb
l0m3TbFBVdg1OhO/91pqneZjQEV0E405cEviRWCZJ3CXRk0M/7LlyrPCRqYY9HhA
VUBfvFMb69CT+oaQyJoGsKnmKvk+s8niI/pSudtfzSj9MnKbJ7hM72Rs8RbWOAEZ
r5MObC1DAEgTPU1mPwft612YJKmDWI4ibnO7A66ArfeLGqHGnoQcV1oAEOzvYQas
F2usyiOwZEwRtnStdcKIEUA1mwYo2JESrLq8wHqdv9pQKXViYLz7QDeeU8dO7eCR
QKzcud3ev9cJE33qeb74MFkZDzSLbGPmjGfIrQDknY9EHvMsNjya/67RM2PCp8zz
9EXnBO+F4CwOkAzxsJ6Yse0132EgWymOF08WtmnNC6l/lkUKeuholtox82xjegL0
r49ub/LTQZyXaK9ib6oPDp8Pg8Xg0IhJMkywWgE0NP6GPP7qh2EW/k515u1Rx7iW
x3hUvtM10G7S7ZX8aLHDk6OktyfYnQGip57ewg+NA9fR+mZJChY5hHf8TdphNvdS
9n3q/mQyEu3BCaWjzJ+konbrR4rsjthR6NYab9qYcF/MAYAbNWus7QcrrCgLIUuF
W94FmbxdHOnRM9205k679Et2oS63a/FhtwaJd/X4r8X6IxfeYXgJFzQDPtrk7HAK
k8N2rMzCyWjRLgbrMeG7aiFO4sA61pISBAVXWyPt1CCjPHcaKrE1LXQ1wQ2I89o3
fttEQN36QCY+O9Up+Tmz2rAFv2yzfJviPp0mqHbSSTYO0kW1iffigyKAPsKxTSMq
Tsn0r2PC2vPlTVgboOBr0IxeXB7Rcl3MkQmYpC6A1ej2peCj74mqjiAxkoh9o7xN
6+1lm5z4L09nCYaTmYb8dnl44L2lsv5pqotMIAdVxqYoM5OASHs9wjkIaE6ZWkdK
NuHWfQxXtCajvy3AB7cP7VumYkBE8HBlJCkamfATtRzZeNIvcJ43jCCP1xltVPZb
tJ6kCZylTDSil8R6GTTsRh3LzdhPbLuONofttG0EZImrXEpmNJACxIG5j6SA1mvK
r4pYy5iu4bbcvcUaq2VkHtxlKtPJ8uUg2FaCHA7ovytRTkUKiL/CMY9/WWtrAZij
oUO28yj3vHSZlpqYqPGGgF6b0Ip18RlUwb9zGNRz7V4PTaJeTsfNWlzyvVR7o93j
7rTZEcXJAqyRPaIfLz4x3n2ueL71rJdGNSnZp/h1IUveigf7WLza4RsI+x7/VkWb
P+Zyd6IK9JVth4Yv7ic7gMyj7sPlrQw1qHWTwBT0B6bwO6GASFO338IR+wOzgdpY
Mkw0xWV45TgXXjytsQWxprSuSTI0QOnfhj+rHlU0iecGdYUJk8YNwaQtHQ+2ozxW
OSJgfFt+/iKgqQs7lP9zn06hbGfMR07g0fhU8INuEJlFCRnomWACBndjbNWPsNSb
w0UwISc/wGCxJiyJVeULLz7kO8d/n0tfiQB1qhqM68DzNfMQh1HXGptpyZNUUCzk
OwV9NZmTuxOw7PqsRJ5ARy7c+KKaEb9y0uIslpoMd+iDsepLfhz/PC+GmMw/osf+
VR9YW5i/mVfzBHAtSliMm6yE8rLDsPZSK/7EdkZLc51mumkHG8D3cJj3cGG80eNz
Jitlbr3NdNIIATvpxCoBVSGyq+hpVr14Xd4H0kCsqlUmG3CTNF5G2vIBCChhAyzS
PmW9GjnmTIUq4yqAGLyX+nS0371yUbLy3EN0I7pzDrd6b7yLPcDKfukNQXMyCsB9
1DvT0z2pCEC9DrILRrWKhEykcA7eTqjFq0xpnOEfRbu/lswReqUrpHUYw1ZmUUvc
IkXHQhTUaMZSn/u5z/ZYT/jYsqz5vXgBpCTNkTQV1Ai3RvA6sZuZ6CZ5/C3fCwV8
+mzaBHT1KjZyDVpvU8ujXJ1suFgamgx4Z+4OlDhPJwWT0zuT4eJNGEcJnRHEJGL5
hACi3hjzpBNnkJznXZ6l4yd0wX+nGy9YiYl3yXXKxhQDs8KK7qPARiTLRSHZNbKV
aRpyWcV7CsZzbRX4J8z5P3SSWKPSdjw8SnzqrfoA5lXi1ldDjglFhONXAOswu4xP
wOGze0sYtGlqFQzwHo5eXQDZObbqycCdZad9ugoGN7HtZo8iCp3DFoIQuUkMcHk1
wVsCHMDjJffFkAMw5crf369TO+LOO+5Yy+YbjRGDe+imR2M8LiA+KO7vwQ7DYIEH
0akkoviRsCvd/NZdaHlHQ5yC18EYjh7nCohPfBgGDdiKeJP7CH3YplkQsXI+IMyC
8A9myCgegcYmWI1YPEPE7UZXftzsCHdBmYVGHWVdfUVaphFwpuvJjMBmmudJ7Iha
DygAlFyodCfhZA8GExNiY5vZv15f0XZ4WKO3tfihRRj2taO9/YQNaP7h7kEf8o8C
5F8rm9J2zR4MoKRAQZV78UveF54KCUTQSg7hP3RbxVtqgxPfWAd/uVUbSF9N5WfF
oLPpK8nt2+tZeG3zGHCHVXywvXPrrCixjdwptxx7iw0rJGW2hwUYAPEgLvwHnyae
9pykOyGPl459iQHHub24Ev9GFXJvaJfuUIB2mI+6dZpO2imvKuWVdwqjVQmkmNv6
2B5n8ksG5ekVooN5dBHBDi4/W4e1M8lXjdc3Ypmlz963y2FtQYv0jfsBX2hxxrne
+yvIDTk986saGIFm1TUcB/CoZdfgBQPGqj3nUA1kU0ns9KD4Sb4KUtE5OoqgT/Tq
lH71KlMyyvYUJ6AUd+agZlJePbExD8TYexCXhY3AbyeSB+nJWl7wLRIo1HqY2KGw
NZsfdoCPba2UQGu66gb7oSZqW3ZVJAB6RH4nF7g6a/tz0MIrI37soUpsFVXt0Tdc
SUak9ivXagg6kBOuEJJxqXkEQs1BpFa9gB7TlJYimAyHYnsPdVgjpNMGCl4vM73W
aCtDefWpC0Xatfq4xejYjbykcrMbym4jC+nD2lEGW9KvU06MA90n+GMaEOSzRDi5
Jo1+0pRfXZ6FQGpKbElzsuD0WKeskBSjYOVVV9KVlaMhaJ4/jgOpJGsqILDffVx9
0axUAshJ92KiqFlsqmmufVBAYiqctFfO3LLkz4x6JxkyQN7pp1jIgeqPlW9vdnbp
AqadFiQ6kV+/plunrgy+SDDQKjdjbC0OFXjLLFaLVZxMh+O6jqdPdXLPX0Arh+w6
8EGyP6hVDhO1e3zj+xCB7feCPFpGBSzmWrW1/u+shRsyScNNiST9BXrfYTCEsvPk
lkb7IcHpqKN50OXEq+UbSD+Vqv1O9FN6nTE8u3LdJB4bOWbaHE1CYgoEsimYXe/v
rkU7Pe3Bjm5v8XuDgq1/aw54J1FJBLebSruZVJ7AHp8cpkHfPCOS8+oor23+WXHR
K3jkX9QB2ERAjBSMJFufNZqOiWWwFI8jqQvv+QhzM3egUDoHmxhiiWIDrZGkCcbz
PCR23YZ1pHHKYvtun5VgWSYB9XNdPvVm248guqii5+0vLjsX9/E/mp3IjcJEHnce
rh/l02qeyR+5pv2wYJ9zq9E2nEfdCekk73LRIxlpJ1yXaI++9aGLltAbRxoBrSaz
+AS8/NWgumYcrvg0Jk56SpGDX7OiQgskmKNFlQhR1Ddr9MkcygNAq+5Xm4gy3jFw
t/pog7qUnAXPownlvdl+awfSluHlcR+VUfW1OzFCaaig4/Lu35lovZCaSXRfhw9V
RZ1IBqobL6qq4feq8vXRg5HLSFDUA4oRFyrPNBs/bJCLULy1s6FMNu61erXPjc0e
04YEvg69nXOTaAn9cuRdumgmSozcs/hnvb7ZkW/fuSUvvykPeJj5xcSSL7a5JOA0
PZY8o4HkEdGWOOanwrx7wVLtzXT42ssSgIW+QhgFmQ/Cjj573qfevHZVVd88n3ZV
mTjGt2h3JwD/0oPt+ksiqLX9LLT0CCk5X6bKuDpjqUBtpMgDNk0XGqbjgAbCE8C+
4TugKCYrvoRFVd1bC/VUwNKTd2OFtVjQpV8N7w3Hb3JZgkyNMcN8OODL6aaG0hMH
XcKcXTdLZrJOQbw1sTOFNw==
`protect END_PROTECTED
