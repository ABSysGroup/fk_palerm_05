`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bDT/SBTszU3/vr2OZr9pXUIyUVO4dXBOzgNVLiO4YSNfxcLQHDb1jkuwi9VUW9GV
2iSPMNViTZVzXEKp6FqtxiPkT6YZD3BYVEoqiGQ6NXtuv32INCBy+j5/2Dsn11h9
X7TYGxb4z6a3kL/HqYE3CIkqTyjuRlzirPdjlWiDQu4zqqvH9kAyNJImpZQC5r15
spxVnNKrnZ1pHV2IH2jGnx4h3EmaGcO063OQvgHokZyRQBc3tlMh0LhMD98oBAJb
V6xYkdLtk/a+SXrbxxI1lVzx7t3IpqWn2dKfelXgww7Fh8eIzYKfRFuapXPqltkS
CsMa7qqR5Xm4enYuMpTD4H5MJG00UBFyqMDGUOYzAOCgNJ1UAwCJ1S1lUObNN8NF
Ej7my5fT067uYk7A/Ru2TbTfe5wjdSCJLLu0CXvn2gAque98v8BRWstowZs8HgAf
bjmCUP3rj181q+3QgUZsFW/csdQkt18RhfaTaAV9nw3V623jOp/gctdudox5uiob
XJWrxmWHITxeE3PwIdt5iMnoBRTJZVxRA1I4TZWk56tqu9WzIM5kIxOKRJncBxWO
KT2dXPyxV3IYXHm5+KCsnQ7pR9VMx736hyJVwuINAadA3bG7/26is1Cf0Z1Mwo0u
VRQ6UyvzXgwXG65lSHg8WEiqwf0c2IUvIx/IcUldHjmylMeNVDvOfuZfI+YCquZA
Q3W0O12SbIi0L+tctgryUQ==
`protect END_PROTECTED
