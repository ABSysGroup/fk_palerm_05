`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aATRyw/HEEb6O0AzdTeQwg+2F69NOZ8tEeEP5V3xheIuKJr1+0U6VoTjdffgmZYa
9dk3HtWuhXwDE1gYX8/B4Z3+IjIFE7zNTPtEMYKoQoRrw+zauOYJATyg+sNVMrzZ
gcJQWI9OmkT5W1ML/+aYtYPBF1oMfNr0HRmHxbRkIhwNKapc67ZHsAonsRag/oiY
0knxxeHOEbbCqLfmXjMXbbUbw9Bl+H8/6Xvegs1mA8/5yZzdjbizJmuhLKiKuvHR
NQtSViFUH61j86oA4/cHm3MMZNyvVnxHRKESpltvj4vlV/qWYYatzxmERJVKyV8/
j0JGHES5KgDxpMzRIGjg6AFM+SI/KNz8SYxJjGZgaDgptAjAiwLoB8irUoh8LYDB
rR2AIlEEmP+rgK837c3i6AolWRFz4rY8R57mRYFeq1awHWQxq6rEf2eQYAZ8XF+a
6sNsIYZl80Y+OimRNMzFnKRYizXP3MilERtDw7wAyiQ=
`protect END_PROTECTED
