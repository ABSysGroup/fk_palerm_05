`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YL3lN0GolwvYqghXmMAh16YgVph7T1qRunt6os7kCwLXWk3O13DeUYfSnq/s/RkT
+9CqFEFaS7aKhbe0i+csnxdiM3R2CawuXo92eOtQaFzkLKh/kFuT6uLm8mpTIS2i
p90979vDeyYKYJD2IW2wimFKg1euCsAj56SG4inGb7k+z8A3O/zrWXFr0RgaKU0k
SKHVWzPaovJhvalkEInrGQHw/6xe1ftDNVJwgclZPSB8CQj7riWAD2mc+8RabdAe
d0RdArvGBP/IqK8pX0YC5IK850WuIt3e/jA76IxjMqH01VJOVC5RpmEoFp4FU0OJ
P9oPa8C9t8EqVAPu+L2hZydpyU36YqOBMqAJlx32x9WbwSgwhzi2sXpAEsNlrZMb
7TFfk6mNDQeJQ1z/rDUZZmis0vGFBADT7ka5yBXnrV3kUoEVAzgBf4/AJ2HcXRK0
`protect END_PROTECTED
