`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xnjO2A8Rm0Sk7ymnoOnaNkYYYwUTC9qupOwMIwECD7eJS3dc672zMNam45dHVUYG
O/0TFtNj3D9a8c7EN3sKDBJJvcRbXQRw6G+K7lsEyCE8WHKS9str1aJckNVTkuXC
j6Yn4cqKBjG0pHBEMj6d4zS2Pik2QRMOIjE3tvzoqfKm0dbKwNtm0ZpjPBHmwjYb
2FOSeXlYwrXQ13cSjVmUlh9aFhaXJrka9F40hcvvTYZEvwYXAE5a4XVNfW3PGoNP
FME6rv77UJmzyqbywqid4fyDkEYAisFm6F7WgrWpRSHqJfrPcXffXMxc97uP8CkL
haAXd+WqmqnmmYb+0Eh4WVerltDyDtOZ6nxX80iRi4lg5Bw3iofQi7eVN93YPAAV
LBNHMNorZrfEYy8wPg1sLKBoFPa5QCjK+6YLYE8t8NwUBzuT3hlec3b90s9AYY4i
hQCFKWYBTrmnhjd1NwY53RnO9Yp+QAJMoi1jlVoCHJatHuhm91dVgx51QA+TlBVe
mQXwZSIlGZNdxlULC/PFdbyGUtn/gwQGWIcIOOaA9Kw7DP10hDh2ElIvqrlXycH1
2Ww2/O7A5TUMRAOjuN/wpN7UMM+Y25vd6rkIW0b1VpuZbU8jRg7AXQCdlV+3v240
beQVRtLwzbd/SNwF96Fl96wlbhL+P4f3iYCCa5/1iIVYUl6UmNld07bta3LGO0jq
bbWTvBDJdgWTcuIfv23b6yOJ3mSRZ+mL/JHdYDDCC9rDONhwxCQQc8RL50nosnWg
oSUOM8If2BRhUukbOYvknW8MbUtu3jd528bmxyTxv/P8kaoITK6EP+yBy6ah/dz5
NesD6rtT4NkxXjMK+2kMl15W8UtaR0gfa0l9U3KzOyThuikJLhlAexwvcMHgvTwS
KWSz5c1uxBphxCsZcMQBpvQrtsql5PrL+Ah36eckgyM5kpKkJLh41CYXThWZX2QG
75Id9Zpud2qqDBRqEk0CogmtqWaniF9HWCo+IyhdJupDqzdVAr58ZW7MWYhT4yyb
M37t7dXBA9OP/ISypzwJAXBtM7yf1fR++0ZljMuCJ8LW5yulexM5/Qy5ocRnq49o
w9QCYhmaISl5yEbjPV114/5M1xv83Fm8gqAs73d5E0UK3USPP/XNw14/+eVkZTmQ
jbsKFWPM7nqFKO4EBeN2x4S1zOf/K9Ib61ZrHNzGimIM8zpX4ZV2gmHnqSsfvj6a
qsfg0jNi/WB4fLj0WS0I32huOe4qKTxq9p5ClLFOxeKAVUVLbISkpI2tJoYOcM+O
`protect END_PROTECTED
