`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a9gKAuqYz6KGHSSpP5w/8GboTvyxhRWgOSUsACjEUae/R9EaB3vR9FkS/D/AqDmY
Ix7mWpTwaLzq6hq/gKnUK5Acr5yB03oD5K0vpXUWh55rF3U9Ew1xw0IRJlR4XhPr
ucRPCNOO3VomzrFfV3g0+UJ3V5RsZB3LRHjxjz2nUwVQYfFsCvtb0/XPwbZD138o
Bgfw2DzhxpkFg9pvGVe5snbiZXBaQcvq0WIC4uB+GhbvGpWJ3sJcDbVld+XbjjZH
AzBpNnbYI1SxJ55bwB4LrfmphWXkZqEPenwbEI3Ey7AuCiFc2ULpf9yDqKELZR6a
4qlsylUIZoo9TxiicUd0+6b85awiBWGab2AGaV5scCJz6v6b006V80WcbhGqYuTR
8y+9Ffw1fEyXrd3GmzpsVSmq0D1E5qfhe69CBUrtX9HssixLjkuhTd8L69XU4HNp
KDd/d/hfSGms2Znp77L9Ut490kuo2R9MFIgDmxg5jqySdnwzJZlP2LA0zpVxtFPt
YnrfWIn5lbITMBW+nrsLdIyJI9oo8lBFf2JbIBHve049jxldrIYug2auHObxYa9r
shChQJtKU7XKifSduNiuWOzrRs7evdK8zB3sPWFZlBEPS/PW9/FGGqX5RQOZh+sw
QV80mHD6Otm+dsqm6CgDdBOoITMqufTwhhsQcnveTOD3Nbe5GSKNPmJITOxtuqrY
VGutrxGChD3wHeJqOs/TPzDNiJ4twiSQjl1R5Vs+Pf5aW7tVOnkn01LlLkUDORpS
Rar8A2w27Da+AvEkqbK/DldsCoUEKpgdT5atzPRm+Ueq/GRxcUKew1rfQMU1shQy
0HTLoPUAgHE9qKFiARAk5fOSCXj5jh7wQdDskGwvVZ3Kw889dx5Z1aYstaCkhi8g
8lnRpyKYBf8j33LK9jxyRaSo8wHaS7uUdil/pBCuwZwuWAl14cvjJvEcFHHHW8Z8
8JZqlPX7Yd6AkZJjDcHl+KYV1KyE9ClEr6f+wOMrPM2ldfYMb5VXY1AQmfzQKWTE
MAk680k/E4j4MYqrA3Z6YGRXVaWEBAxQcj27aXJBGzmkhgxEV81IZFV/BgTQOK/S
SsbeKXNEATYkWXNeP3WfG6HFajKuXR4c3B+cf0Ea3nPF0quYKNVX2FCOZbNjgtRI
RywMYp92UF4KopoGz/nYuwn/IS2UqaLVDHuRjkT34PXdcOx4qMxZTiEFYA065wKj
Ie3HFihjCcMa8GHwKnAudZB8afjQsHc8KUdmqqgEWvM94WQgf8pFdvjHi1/36Nrx
YqIL4Rb8IrHT1z+MHbMg5b3vFfoxnyEpcSWgyeDuzOfCgd1ZxObQ8hf3s0mrxF18
BVC3L0LrdZdEX8OU1CONydu9TsewaPssTvoIz7hmV346/oRjYBhqq76GzjjpJpnh
j+rw/dHkkgZemiJwUVAgHffjnhJ6X1/ov+qfITOgE2YvKHe1wcrqjApX9wDU1YVc
4AfXSTH6yQ8NYdiQF6X4t4CzhAf1UTdY+VNh1XvrTdy5PLhb9AtiuwgRnEkUde6L
qokO/AxQKqEAk649kdl2yQS46fKmTtrf4R7nANL3KcYY2N9vn6Xm3INd4Z+5M59k
BoQFYwHN6nYMjli9Y7TBCGCF2iPiujgHTFTZ+ZVE7WYcMnKqN7MmoxMSYbmhfDTF
XckNPD5+7aGcyjoT70z+G1mG5qsXja+b3Dg5R60rsNX+doa7oNlxFQJ/guv0c+2F
8FwPusqQJObK8HUq0gR8K5y/+ttPHnAwSxL6QY45FIHCTiMIyXvCLzc/7vWb/dUW
4jNWq3GADhflJMUrATkeVSjIkHCer/9swyhxka9srP2mrvJTIKqTFlfTaVm9ZYec
g9jCIwgR69qW6VmwEWfHVJUP6IaRquAW1fVa5RarhjTExP/3qxAfbnDdrkTf5ZOC
4hBloYqcZLUeTE0k1z/U1GCFJ0JDwL4ajMlZgd3zMEXXUcYvauGcKMTYYdRJQtjM
hJt1j4Ud2vPs2XdiDLp+Zfi9K/JDWxqB6h76AaWvwZ14Qi7yJy4Qqk/o6/0jbqQD
ztu7gVavzC6qe4tRpHGczKE1Izyq59QmxX28mYjBUdsAnVtGOmdskIDJdEG5vBMm
YCm/nUApOworS02r9zjwEYb+1jar84ata1g/s2U32suLmRd2pjJOdD0lMkVq1GpR
pkluqnBhzTzYcSKlkCfrirNGpgFFJR39jUrB3yawI8LEBxWwjx7OvUP0ocIJmugS
Y/N2P3OS1ZoJt4SgSCDEKm5X2G2+fmFLqLGsmYvRAUC290WmybbC0Eg2KBMO+RLL
BOK6mNQP7KVJ7A4Q15y7PYF4R0XVS7C2q1k/I7/HWBLf1MTsHvKOO9uf/jaIp8Oz
AxyPqmYSo9bRXXaJtbohpXZwwmjZDEZsSBc65gsfNxW39YRfxiKYx8MzykKPFw2H
gl58hKT20ALF8pc9U8YD+XmBmh0z8y3qtBQ93TTY7KJ8dVq5EG2yjc3p8kodB5O1
IFdTc9FaDiOMGVhOTKuoXcEj6t7Nz8awRNZquZZoCXDrmbCgVyoRjQxXFETmBbzR
Cl0ab6B4R8mYoj9iRrBGW/49HcTAobB0bG+gdR93brbWb7cfCQUeAWXhzaFprXjp
JomCVrK+UVNm8QALChL7e3PyFHnEEGHWVQCUaaR84RzAzTJi9VMmT3cWBI7VfMQs
iuOKF8Ryy3+xHqzKaLsfuWpNuK1x+EwQsGCDpNTu5evTu7w8M2yrmQ4kmWHUiZGW
lbQ+0mx1xLhiilmlIZ51HQJvTdvpO1IwIRkovomL0w6a79Eg+60q90UpGYdMlYK0
bGPyHPEy+By2GocMPsyKDTvESlMRZx6G1LLy7VWeZu4AdwWaFDnpBduHB8czJwkK
ENohgUvGocJ8b0fRBwauFwVtIKLqX0Pl2lO+BgRryAXzp4MD/S+9LYchb4tQlcor
QpL0UKye3k7Fumg6DULNTIT7S7T2TKnNwLcn6HZNv0fuiQTF89mI/0DlQlq/S/Jv
NsLNzqL2fi+PL9PbhoQrRo8eYjxR0hlYDRytYUIFEqVJaGqS2Y6vuXwAi61XHDaV
WvaY7rn5vknq/qa3O4mWVA50lE2TRNUa9aoHGhBdx1L775R4NdhvvFmUqf1C3uK3
7Kdx6NtnoffVmqXSBF/qiAnDnwv/a/vv9CS6o58l1kRA6cwIv40329Bmc6j64gnj
hNZeuPUNjCdIEKDKBTMK4xu/G6cKoD+0H2bDd9QS1OwpswzPcGSFvswcJk/WWl1f
RDMdB5xN4dFxotb1UlV/gsTfQ9lIN6yzR3ibbWHIAE78IJpV4aKGtieeLPPnzf6W
ROyRt1E7FJOntdk6tA5ru6sLtarjLdZoVU48Ltfdb044D18chKBHYoAipYsXFQe9
trI+Zao7RaL28w5U2kBVSKX5TfAUL25Lt1tkiUmbIsVqZ86eM4F4CwKwDgH/RsZN
Jnp/Oz7DZ6fRe3s7FW3MNjwrcYR6vLImMMfq5sAOQ401y8IFB97zLICzZIkEPE6g
qVQcGG2PabYd2LjamEoa8ktSY482pNxMEDIPfi2YtaazBkMS2xuoj5AdyGUKjCbX
Q+XRHm03Qglu97D2DMhD+HjIlXdCC5tOSefA4eXfXQoT3Ec/TKRUrdgMjVRRsNgK
UyWIUUIUeWirmPbHyGHwCWUNa+P26CMC8H1wPrrDJJHV6jxvVTAfa3McEpDGAqW9
0g7kfGQ5rKmFPU9ZLBrnSs035mwV0LEqcp2gPum0R1eqxx4PsFPpV+ymYmrwTInI
txKUv1hSzWlUlQ+B4EOugw==
`protect END_PROTECTED
