`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X91pL9SLU4APRDGn44rQyxpd23I2Hww2kapaIQ3FwMh9wCXHFX0fN1o8sm9PpzgO
5ELkg0wrx5LP80sTa2qfmANONgzyd1H/GiepcbecR+vLDiJYFDp65DGVma8MncIf
pEgFTAdwweOij0RFnWHnwSKjlhLGRJDJjyv8iLbGQ8L6GSvTm4ezwo8GCehJs3Vx
pGsLXfFduOaFA+NcOnZ27YyRb0lGI2kdH5sgFtZJxzWuxFhR9ivNb/Rb+iMtAxnf
HS5XgSLFx+OfeOmbd0DyNb5zDfoM1wnzBOdRCImXaPJ93E2xnO9CpMea1L5fUkAL
NVFOxW+0nWmvpd5SQCLolkaG9qL4w0YE4z065NdD22B4PAmVJ2pL6MKyqnezyhxv
zoPUVPELG47pS42LN6+zdefERoSVe6VIGkoOUlnqGmH0NODE1BDeCnsE6o6M3GIv
Oa+q/l5RFnL+ZZVWKJlBvsF7YHbqQsHeGe8h8nPug7zp4F97RNrWPl/XUBbv/36s
`protect END_PROTECTED
