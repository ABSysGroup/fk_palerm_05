`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WaLsPHEZ32iccs09E9gtVRZ5viMosVNhmyBsYZCk32iOial0ouRCFZmAUa/otucZ
qbkp1BHj8JlktUbvUfyHIgghkqBuU5UcvCy9/jnD5Khn+Q8RSh2yJG0JzxCONWVI
ypIz2opsC37zrh7UVGMqG6fREGXH/5SGkj3njDlMvTLxnQ3NJlDW9bb8VJZT0hZE
fazVo+LMWpPhR20ZVZZlwr2O3Md6tsazCuur+iXpQ+CEVzmNBJlI0B7cjqGp7ctu
/eb6BeqYsp91NTmfg96b3pQQmDBdWVnUCZNAJGEaVZ3QclmwXOEfG9fYI+2PUApN
lkeBhnI1hvTB+h2PTuiKf05rJyEABtjbBsNO9K0qiiTGd3eYOjBj0HDGKf9x3XGv
2ZjQ1AFWf4iDVooJ8Ba/CwcEpy3yFl04U6/VMUCc2zDygB7it1/KNNKQT83TbUul
Tf8W7REe8a5opMf6rQ07AURcNAoQ2iz/JBWzZJhtc21b7bi+am7VQJNEvUVXu2PL
HddBMnezfJPxhn9UV0/HYdcU8kVGFOqdOKSg1v6Goi5eIU2C3CNcWgVmBXEgc6Ly
s987+FR7sPrN3lWaUqPIC4HA5aUefCHb4Lv3OVFvQsF3Bm85QR1zh02JNv6MllA4
BsLghQWpsdxSIz5olR7GMcxHFy12LQRo/qGmeC25B03XVCqRIrNc99w/+NqZaiAv
zxYg0O4RJOAdjFmUR5L53Tdwb3rQjB5nXTowvQGPP66Svw66pwtjOx+UdocEyXku
ElNT8e9v1+t+JVUx6SK5PsUtRQpwi8BzrU/0ExZgCAX8qdhwXqSJC6eutGxSZdiM
JIDehL7t0GzBUTYdki2Q4U2S3GfSeHJqAHCcJiI+mjJYhsXxouqkG65obIdwop9M
lTM8FYcK155bLc0zYxpQmfKQS/+wGWd36/ORUNUhp9QBcFrGtTmQNt6fHpG8x4lr
Pac3JMJEV1KXXb5oiSTL2KrReNsHwl3dkH12lb4TwpIXSQPacjjqQ3T585NJTdJT
+hHvYsQ1m/LQgjXF+pIZzHSijKs06fk1Xas3f5OF/dBr5CvmOmnywaEj2t5PvW48
6jDOPLEwRSOniQJIZQkK97it3LPAlHb8h9yHIjlmZ1+kOxUrawEW1N7xHhzgTzbY
`protect END_PROTECTED
