`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8TRFjVChtMnOd2p1f1j62eRMIqB9LedNjVY6NlM0ZEZAXJcKCgCFo1Yof17rcNr1
TMpfdmLUR3M5bQIchBE1J1UZN98VBzw9KeLJR/nLlkMVR5n3pGIVTshApj7NcWNT
OIjRY4V3N4bSBssFYxDa5NTMLh0k3X5Sa4i5k/g+Hn07MD6L3BOAzpqZh0EVlB/1
Fm7jHMlYiW8ES8r32IaSc6pMjWAkhcKoo56UZ+jyb6Um17yKHEr1LhTQlmLDJTAp
kSmDxd4h6YreVVZh2n/2PZl6xUmoUk62r3MLCcBXjDejYGjfXfWGjH/svy/zaj6s
a2qG8RrM+FQ6MKvkjTKMNg==
`protect END_PROTECTED
