`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
41HTQ50qGu8E8aUCJPKrDfAGVY0WT2CPqkHLPO3XpqRxCCP9Dcjd05i8ytvoTmwv
jFV/73KuSH7dXve008m9M5mOI/CPrnIrfNzYk6PQPuICwRmBCZJZVaMWSnJOn3Jo
tNdP3pSWS86QXKFG2HKXZ0huokdCOUqsSNwcv9nGKXP/ApCIWXnYsCc1pqAUlIQe
jxrrrJJBZJDYiNQp7XtJnEdmjeLO757PRRMFghE2mkZodfI5BWjdPAr7JSAt3HVn
uku7S9zqhfi1ynZldjE3J2JMniOF0mhB41RbGeRkwzLhS3rpj6qC2tgjDs6rgUG5
3IBa3tLCuSr9z1nBSu1ZCVr55PGHN6UbqQI7y+OrcuLPK4lDOIAark28f71Y3UAE
GN4P4+Ne9o3FdolsJK24qfAt3gCA0GO1ADF+ihFpzNNFAmVhqtjGiJTJi1atK7k+
FaJ6o+llh1Yt0hcH34LpMZcHmZWwaRwF4NT+nFk3hLGtJ35BuuDA8GsaHu9fHsb2
488uBshzVI3tmQFvlEznTA3Vtd8xTc41KnwAP9yQNkhemTDk3joHdBrS/agLROgg
pD628k41yz4Apkta9roN/24ejp6Vf7eLEMAUssWYLbzVTYH+chFqyWpB2AZibUd+
IPCp+qYa6iOvtauZV9IMwe0cA60HJskN2f0wvtrFTAtTSwkvuW5qoTG58jnproOJ
Rj0uctJB8KM3gibOm89wAg==
`protect END_PROTECTED
