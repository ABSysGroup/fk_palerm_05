`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pbjHf9hyHPjjTdob/rFC/W/iXmtahJ+aCxll1lSXETbfFn56it9j3Y8bdREs9eP/
bdOdOfJTwCgy3WErhtBHuGHuf5d71vrOseFDKTn/zfWVcvrR5rKA1hhmpfyd4tA/
brMAD4kiqLwlBLwgQMqrY6aoHetILmJ8n4Y5UBslJOuQktHoU1K53a3p+XEW1Lxq
Hc4X/0+FjgS7ya/N1psn6CzzSi9UYAjRxkY5hNABManO2VQQdlbtida2TRF8NGUR
3dXu4B3xcSoMDMBHTPkwKRlgTElT4M2ZcSl1dF143+KdFa+9ODIbHUdLwXm2xyQo
UWGvIzcS6FF0yPJ3DHLgjah4p0R94fgDN1dtRaGASRmll42bqzsa6C7PFUg2jc7x
lgYbYKGxArEJChPTrL7tQs5SUzcHtzQWA62Pq+BUu21aEir0y1EAeyOao1RRLmsY
51fpF5XCVTFR59Wr5wrUku/em+UflFM3nO0Dl1XlsbgfW6MqIfh2rqzx5J6Gvur5
xVpj5an753eIQsCoFF95Q+c2yRrnQkelwmZHV/DAVqcILd6S5YEYkQUrEND1ngG4
iwkbioTQli7kQvCorhpagzJgkGkpzGJwJi/kOrz3F64/kw2J8XwM+u9oidt/g2kK
UYduJB7TAoBV6KSLFET36LaCFpamgCYQWd9cQ3v6vBryU/sIQjdscgiHY+KSeSJ/
wnHWqUjMsGWlzI4D+7AfQzbNuccacIsoe0/ibbcO3zInpz5g4ZvltNLFujzBhuWt
PTLLrHekVL1imNKS8BrLLPmTAC176J/+vhSA9SoepGWPdGf2k/j64vNMljasyPEv
62OyLSbJJxlhb4ex6YQs2FG1SckioU/eJafM6VZwyCp6yTZDFxFKndHXTAmWqjmn
lE888JXVGmNJxwP/ya1Dj0PleM4d+0ZDXklQGA1HzNkhRLe966MeFp6xz0fssZU6
grcI3TGKpS5xuDQ9Koce9MgH1WOXtjdwEuzBYkJYuL8nSI0S/FFOWZoi/uTcL+df
4PmZBOApU/2E+eG4SHDKjU6mZ8AQC1E09+eNQueEWf0HHSFrk/bv5FGI26NsxJfd
2eI35cY8IiUK7OeoiJTGqus4cMaA1Rpl6CMd22hHLsAMkDJpo5Lwauh/nnbPDewm
0HRmEA1MLXzX1NMySCinvFa01etHg8eN9oyJTuaj0+UFnHzqsQavEFyoZ/IdVEtX
S4bma2SApgP36KxTwanWiLWPMI1yrVbsnr+jPuedYCErGspQYw0Yx3V7usvv0bQw
EvvNOzkRDPWRkaRWi8O3wjBTRle6FO7FYzA3FKb4OcIKqy2a3aY5lZbwIPVMMG3T
dsxLxgyCFHli2Ul7faJqbk3HkvhjJ7xZQE4nkCpv8s3U85yJcjatakXKI0XmLin5
my6tH3bguOfWKJOyzPfo0smGTtzXL+iU0ZOQcam5R8GwVaIInMParOOahfdUCCVp
+acvOt4Jb+0vVlSeJIwwRZmPHPK2hn6kQ0q6WijbMj/R5rWJ18mZZDvT5gw+c/1D
fRQOxv8SchYfTPlRgvyJmVsTiI2yDNJdytlRx6ZZN9tX/uh8Pvgj6s6nVCeHk8gm
wi+QjLN3G7ULCUu+Zptc6jM4T63cd7Qm6+Pels9YmPc1sc2P/b3xjLJkU+qoWhmh
kv+yzVIaMRBRzRTPp3uObifpP4Xm9uZTvdM3mMu7JHXQb0SUHa+BofRUVfi3Cahy
x5nAITvHrADF0uKQe7h1cWh/E27LHskhTVMG37uGXx4aWvg/iZlV/cCUSxEpm4Sc
XRxpMJ4rVJ+OHt2an3vXgN0FQTCGj7eaokqEW/ubCgv0xzjTSUoIBfx7uE+elD3I
6pGItxaR7jPVh4GVoR3POtnPxsqd0eipKwCBYLfWxz6YJPNfbxyH4F+EpcuDpUmQ
tBAxYdW2EJZQ6dbO8nZLEg==
`protect END_PROTECTED
