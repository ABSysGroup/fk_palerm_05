`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C8Rz2iVGabPvEkEY8skt30NNelCDmUnyItQmJIj+Cp24THrQfy0gtWiE6DNCGcBv
yDgpcdI/HImswL9/MKl8eqxCbnpElJfuVAEWg+7pU07i2fll6sqT3iw0Mj9RXXvi
7epjdyr+ivjCXD3PRBUMf3hsAnkAOb2burBbc8PGFx6nyxbR1hUxgRIxaLWCE14I
yTdRN2Y5WYA81qqiwPRtxu8hP/r13r9iQie7efFifdXnacTO7/o18j5Iwz2ShPoO
6lZquGo6iy0SPzG5vB/7KLnnq7beNqJHOjs9cXsDec8eAsjFn6mN1JR1qqluMn0/
DkLCa0PsFY5glze7dtgJ7fFxjm0Fbz7BrnzVlf65Xz9hhv6Z8wJufDrWPlzJ4tWY
Eiu38s9UR+LCMYfXMMLPmQ==
`protect END_PROTECTED
