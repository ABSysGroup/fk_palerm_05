`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9bbTNbJBxv822GF5cEafTKR7SSHlmtMhWMjNprVSEC4u5esi7bEJ0W/ItFeE9oFB
B5MSHiGbjgmYwk1TJ75UejWQ1zTSBay1dr7eeokOVpmGcHRlWZ6EnuxmMgQverdt
GlFSGYTS2KzO09JTgO18Y+gyoF0y1w9eblmQBxpoQGkjnPn77ed7abdb22Syh4ut
GbJFQWL45mqQPGAKVjT30PyNNJ6pqah0seLSuym3zxK9lPyS13qYWjucyzxuMTC2
DziZMm8YUIUmrlQqGZlJ8tGf6ulBgS0voOIxvtEmTWvWB4VkD1+roUYbvCTJE6I6
KUjZXHDw2M9R85EDOoGbK35luw2mJoLKLonFHxJxwXx090LRYy/DzWezlft6Nrec
Dce3daYA09EHY3xsLCkNuXQG2f72AsA5wu5CeKLSkr4rxBwgJqaf3kn0K6G4Ubug
7lq+dxukm7JXqL+QR8rFCiQS8OK+3TRHtUL/r9Idb5M3RcRf6CYwaa+F/+N9zkAU
PFqmHJI0R914U3bVcpP0hnDY+OqfeCj7qoI/wCkwKXSS93Th4tcyGEfRYSVvO8n6
`protect END_PROTECTED
