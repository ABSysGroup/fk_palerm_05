`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RxhHgDCy8iBI1vr6CtTxt31O6yXnvvhHWD2dkTJAs2lE13wH0tyh9Onk4+h1vd2f
9H1tKG2Oy2D5ejYMUip+BXhTCrYZKQHsVYrvRHlBlwJYfBDxqJkluq3ATsW8qe/p
vElHAuB4hX/zkbQI8CWVr/5hxqH8N63IUgeLULaDUtHflGSp24pSMSLTgv+5Gm79
Y/7LbXZDlPm1gD/piWBIbT0gWOaaKSCCwVSt1pXW5vZdbV9/Lpdner6iG2cT3qUR
jZR04H77Iy+na6pjyUiUbAb5qK9b2WGFUSzOQzmwGmsipOWAqB18OZeSfooAAJBf
ma74IDSmcuufict59XhZGv3OOTENT9I/titAthi6ZIotMDgVUw2LFmrvzedOELTY
SRMLj03bme+Zmkn6tm7rDSmsOodCYfw3OFFUpbhFYrKFnduFBrlvNvHg0tjagErj
lfT/Yq84/cAQbDqJIWFhSR3mqzDys7MQruU5F3NjgpRPb/jn8+2H+Kwj+76/rI2X
oDQZl0u8ZSygv2u9sJjcrw==
`protect END_PROTECTED
