`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zfbkJsrkhuyYwYnq+JAVSsTEAFVwGhD+4Yz+0jssW4PQul62nrDTn59AQg0EO28s
jBiH270tAr07+2GCk727j0ZgQtDlnMM1yzs3TT6aHvQOVTzshX017/8SFtzkw+1y
HdYcSsdatHHJno7dulaiePDsJF4ei6pFy/SlPRcSNp/j0xefqJGyCDkOJ2BEfEHJ
U0+Ub+Fv8RHouPuzjHWXx+fbrMGlHX0kBCLLWBhlojPgARETBv2Rw1P1n3rQb3cZ
aW3dF9hm4DWwlVblzwlxuvZDKLoIhqBfTRYIPkQ9RCZrMxcNSwy17a+UIceos/9I
Tp7qzTMaoim1Yl3W2ra3/Q==
`protect END_PROTECTED
