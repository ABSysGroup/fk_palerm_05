`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NTckbZsUNazEh+oOps0BD4IHAX6iuFxNZpgisGbGsBokf//qcOu0Lrq81Y8wLiNF
8NIo1SrGOUuXg9KNIi31nGv7s4RXNcG2JqS1LC2vxMpjbqLvq8MIqA+RChKxqKeZ
sV9MrqrAh9QQWtengdlfKfnBbg4suQjU9y5Pa/GwXv0Q67ukz3Yx6/vKw3zKUQYT
q3qktdA55ixSJ1T8FBNMBOIemjVxUhQ16QntsDMT2vD9rmhroo4vgTKj5eelAP5v
/e47Isa0StB17zOOXYObiIVO8acScTE+4pa1Fst6WmJ9FtW1eWxrsyqzKu02bEyv
vOLDjFxMwT/yfceZQ6CZB+dIsu7b4YO9UrEqmPHEqI59C8yriDXIK10M7e9CS5wF
DgZeZ5DiIksUvrp5SD4UlBPBkJgGmOggwFmU2snRw3GfGCIHm13aDc5FVtGz4yc2
5a83qF4BW/B33/+oqLXdV9iHdFwukqFUtWjGaspENf094BtzlYEK50K/d/58O9EP
OGi1xm0/cFzjwI901CrWgvLgobdV01nlUukZb6PEdtUk7uta4Mr+rcgsPitY7JQT
y20cOEj+Wid9rosb1EqlGGZOvzEGuMU/aSV7mA1Rv8dD8zPDIgf9lr0z2Ri/Axmp
LrO0ePsbXHjLvuayJVoAn78ekEwe45RdoeovX9LU77mtPVQ7Ht5vo/hdZxORT7Yq
hvjz5KBgE5ZRH9USr+14vlAVShIrhzpXTuchcPo6siw3aVQM3Br4lYhvbpC8qLAU
57olLyR0yqrASknzXBtaXyxYXxfqLIA+JghvIxlbiv58LUwY7u69pHP2NzmqPBmv
vrRIAQgnVCDwMqz7t7ByzgYCxyeiW1GtHnbQ95yx/SnGx+UevfH4hIwgILHDi1tg
ccztNVYAtURO/vtBISEFHnMcR6Hi0w/9CXxbvdPzet1mf8LNdCUDt46F5CrqQGH+
sm9NSbE0Mcl+OmxeDXC3aXKDPmHsWTaxN8AMh6qOPmJ7wKyBd5laYrgcPuDG1uT8
hkFiC//Xym1E0Ag50ogJhb3ufwYBa/rP9eLfTFjt8AEaGvPeeoP2qA0WOF9c8WJB
CKIlOyCRQC/wkGAiZrtN2JQKtKt86U5w7rsuPNrbiNPghlHFfz/cvMPfE82J+ajX
e4eEkUiPj9dFa7+Ya392OqjlmHTr7MBCJKNox5hE4cQC2JbwfJrap/1RmNoOE8Dj
IKcFWweybUgEiCrqHNyiFL9naKt/diRF23iakCOhx2mh/8uxMTwHK2SWcZz/9k0y
BqX09uurRH2K5igNdN+/cXPr0F9aweBwRpP40E8oQMMlADpR0WRS1mRFZwZI3XYF
4343c+l+ftHGgqdpzv0+P/TMOH6KfOgw5oSzZ3Om7zGnPTkhOd6+A56UnVYwtVcP
zA0NXiqwQGpTqS4Ua6F938TPlhJW378Q3HHXvio3rqC8Yv7S0xliZulp6JjUoGaI
4vmh3F1HUI9IZQ97cPUZeSAkLDFLR86jrRQXGrnHzMVTlooE1jnT8Lzdyf4hAtUu
MqmIkjR9L+sqlk/sTJRpqaItI/kVI5axuNAWeXSTjore+6Tov+HzvP08YlA6t+CQ
lPCnGunrSOLGDaphr+Y+lPCC863igwf/0OT5+GH0waUUdQSmOfi8FdexMicN3fnz
2fj2vyXvqaTIW/tURrrIUyVP+zcPehsXk3+5wh2+6lqZEjyR0CkAQ3yDXUjav7X8
iHgUsLultOZh6fl5+z1rk86uUUUzVpn5/HvZGHqDpxXagGugfUj9L9mqQCmiCuFW
UQy842n+5sBE/90dPgU7AtZNPU/teLka7Ui3kvfFccWQLnYpGxSD2tAyonqRQkiv
UGERNe3pHvE6hKTog0RO5TPDLZujmgyobuzhlyAKaZb6AFZ9Pz6uvly/t3a6ufcb
GJo7C0+HRJetgSqCNMx1dP3IERDXCoulbK7Tr49t951GAOplLHARZF7a3ypj3+vm
AMnS8O4t5f331Fs/zcpV8q2u1jC9whoboObV8khR0b5DIfjNMFicY9SbR/tnnkfb
QRpLVctYQNdHKEGSmDZgQW2rfv00wGq7KcBKpKNUwsDTw9fjeW0AtKNo/k+XqyjO
Mw2TH0Z+nlBtEMsoRX/XUhoOI5iPHmy9Ff+4/vEcpqzGnStTX5s/ptjR/ORB9mXN
O1CQ2aOjKpow8islZGoWML4+GyJs5Ibeqb4mzuqVvJkX58T7jeE1y/u/rQwlOhxa
fr+olTs8qx5uYyjm1H4jLgdEVNq9mflpha9oe6TofZXsu87pc3oIKTSKO5OT0TYV
TTfn2eTL/6TzfOhH29LiwsMJL0S3cv3lFwhsqWPPVLAFg9YfPvFvbFmnT/d6NxKq
R+S3sFQcA99l3aD0B8xmBkQp3AgTdGbXPPnCSO/qAVNrU4yuqlv2brysenTb8Fcr
S4yxh7iL59yF+LACNuwALn93QUXbCr/rY71DggCOx1iBW+vCdZfD7hAhRl2idx+m
CC2qH/FDzzkMDNeGg0OMdoWTrxRA2C4UH/wnIHltxCySTNY/2MMTY+oEkjHtR+mI
CCiOgiIZ1vQCz8MmumLDBqIfQ6OHjeEmEDhNvyGaF+F9jr6C3rWMNAEwoQBVTzr5
xtffbpUdVT2DUya4sIWGXYlkcHs2J5l2BprTkXrKHZt6uE/Ej8eV2N/RTwdmLklL
5Aw/eXk8IeFgMa6tmkTLBg1jL09uj4sDuuYOti1Hp0JAkzWLrRsc6EwfsgwMX5qc
3oqWvwYRnAD7A2fsRLFl+33AUxTnveDcdqqyyX6FMbI=
`protect END_PROTECTED
