`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bt6VOoDf5jE0Kp6EK4HvRy5yvwlEFMSJJ49LYLNKn7t8ea2EzQmh0zqNdVKHru7y
VVIp3TbxZe6zSU1bMei9eenmn7fVV6wDa2ovXvOjk+9FjXixDMv6OrTz+9PUwcAT
kPwQXxu3NHy0sFuBbbmIpP6D1UVy/LHlOIOqOwQNAoUKQRYTBKXe2jKY7uuZDUmU
CF1n9OYUw+iTMiiAPF0G2QdfdYY4655RZRjowFssbrbXO9ez+ssSazEDAkaS9t1Y
iKsui9QgXZonZG7KHiizgA8sJFte8sYsyMdKH9408nA39+lKAdMs8nSP2m1dsKnW
L7BwpUgv8OiekCYAUB++w5HnpzKy7G4wLSUCpByGrCjyGofHsdyxFHtLHA5r2PM4
CVcSgY6bOecR+7rlW6Oe+Am/TKhzYQZpI5QI7Am22jlgVZ037d9vmtfrQWhGm+Xp
HGWiBDNoX6GwOzA9/0pQZ6Op2TOkwcoOHGhtVs88Qc/1LZiDg8m5vSCRILxMNByC
u3HbnjswPc9/fqtBg/+KsXXOlJlqaS3LC0nG5l75by0uGm1a2FRsFCgt+u2xUaEZ
ZjTGY9J2h4h21surpftBbQkXUI136BZYPvkJff3nVbFiRFZisTk6HlJ7zvod4RUR
UVWX5/xok0BahVSoPy1N6KXG13BoCnlgyUMc0/FUr8usNA3oX+uLvD1J5ckxgpJu
mg6PoETYRmwWkK+92ufpz0N/2fnDSJMfhwbYX/9ccmQ=
`protect END_PROTECTED
