`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lefIHJP6Nq2963vfmmgRTsAWufNXGN27dDRhVv9XcMTt8yOgUfoE2VGUe/oYtSvY
2//527HC0mQuEdN//ZUkLh2iqvqU2yqGxmlhUMj04/HuBbmiW/r9Broeb2BgURDW
HIHyCbBmJIVqVX8zGK549l1D2OoSBssruhS51P3C7qWpSV+Tz3Qy8ZpwEtdIIcuY
HX2DH8U+cfHEuXySIcEqCc/RVs5Wg/AUGW1P2sEWibT7OI4IJvQYsmi3wsKYzkIk
qtZw0NN0rH38CXJhXrLWTJS84AcpoRSvVEanKOffp9EHu3uMD2YUu+Qcc+R6lSi+
RQE70RXx//bn6rb85fyj8NjKs1QA/X/SwO9KlSaa/lXFPmuF3jjKnpYPpyR6yo5/
c4ke5PHeAa5S9u9poSc1+7E7S8QCrZEtSuCMJXl83FKaJcSKBCfJzDaC0N3cSqEU
Dnjrf2SLVgKLFntpI7bF7+4eb2WhNlxOqkFLIZ8yGKKfB0rFG5jH8s6WcegsmrZD
`protect END_PROTECTED
