`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cIhkvAC/u+BECRsN/0iiBuKqGR/7AwffCYu++Jly9hkWuBWfr2ofCVsqBvzs/8/I
wCxVP0Q8afYeKmlcLtkjFiMvkzCngP5L5uEWnBJHonXw7/pcFk9qdLYv2+FsJwpO
XcEUECae5sOGlX/DSBc28b/IuyzhfhoLiBM9LO9Lu8B7cQIfK3QLoUjyeisbob4u
5wKZW9m9SFIPCY4FqhyXpgzr9o/KdqA3akDUX6e5/QZEcsbXi4CV/zGmXTosLive
MRdHqV71NGHzBxcMPwq+m0UwfGhs5CHl+RJsKXCd2Y3diYclGMG65eYNZUl6KwVw
yZfl3UhcBTfhtio0nepdYQMGdVLST1PPilmWzstX62venJTp3vM0IpkRKSMN0ISV
jSqa/ZFL0QvUXLatAKU1rNtYCL2c27FD8j3Qqtl1kKBVW8P2qTHyr7vNBNwZiwLQ
vh9NKGe9ONsLdVs6T11Y6yE5az6bT5MztvNejGw1R7UnmRXpDCP/xH7ijp7FMSPy
wrsjqw/N4bu8FtP6ZN/wUrHXeffy49mWctxJd5SiUKkANqEcOMMM0nLQ63t/qsil
DAu85UKZTGHxoG/U2JQKaYYx9ZCWSX0abz9PdL8Djr+H+TPVqbczaXwyNdeWnWnE
JaoWRqEvhwmMXnO23eZ668/aqJtQVI74qXCl9NkOMlZLBg303eAOd1LyBL8d4+Ks
S80QNrK48q9aLBoQbZ/v4E6fkp1pdT/4CI9wrU2sUyePk7pTb9+FSP/WNomNTT+g
W17he9iuvJD6l8zZEFy0iCFoxJzfPkx/IJ5ZcCS13gP3AEIAEYW5QjQHLtBDZGK+
avEVcq1VDwJglvDjOjINa8TvC3WE7yDmmMwUWG/BwNssSBg8WtyiGwWOnO9wmCDI
B3MLl0vSkQLLBzYDSHVXNW7f9K2EyftaRnVXxIZj1DLBn95mbdTuuSnhM2p2WgHV
ugtFahUyfNRcaE+Z9VqvZ70JNvfZ/GJbhZ/u12jZIUoCfJISqu8BARGHtGEkxJ5E
PZ6J+ppo+Y1LllvpEIBaZtt0ObFiRjqOSdqHAIMJtS3A7xJNVWnFXH7F6Dbj+1MH
9SmrN+G/7RuwdCFOGdvuUGQH31mpcBemwc2U95iXV5KYlVCe180I907+tHkcVbvn
EeyrJKvAKIz0ektwlVU2EnOBlpYWVacGvPik5eVY7fvqziefmHNHCzEDyxJ8xFkb
X6cZMQ8rpKHWEktkjSX5EBP3bVPsmdl+kvq/cRkHXVVkCw2lwF5mc7mevgrT/it0
iRwRt5vQOTC8tAPWihCMfolrXMFPb/ot6Rf9YswlQAncZkCnoXNb/uhrWngB6d6F
P7yCeI1kJThD4AG1lpogdUYAr5PGlY9dBNYCYBc9cdSeIAjG3Lc7glvf21v1ZmfG
EhvPOyx5h6RdDrDbXnA8gd9ZTpS0lGHSe62NBNJ7LuU9AVoFSpWd85JrdFJ8OAk+
QPpIFSb0TGWVQPDRkvfuOV1OSjZqtyArRf/S+yoI2vQN8aeYxWrULEOyxq2Zr8aT
n55vmlFAQmKNqhAIuk1W4isypMZr9spBY8hwBugphWGb4dxtNAcHw1PJddlcY6QV
IIrPYMCRXPQuS2jShwlALgElzMqgBLCkN5tlTL3aZ5b5tW9KnB1bl9mVAe/GWqG8
GzBkLAUTKogPzL8roeanBsec4o6C4I72uw7bFrCh9m/xd/S4H1R6brw27tx46tDP
OVdWRKfvBmSYt3MhTlDoN2aAB0CAuh1QAvJTWXNezq0uo94Yb1YUsy3XBP8BK6ik
qfJLCDsw+eraiff3wHrBdpAOFpmwsvBdwJeJ0fzva4kiUzg1nAssm0fDjKGUQHEn
/anWbm/zR0rKYKVIVXiRTDp6NRqo9FSmpedHDPKGYyonMBJTKkrszUie2m4vm8sA
Bm7iJUezw0bEIKJXnIEkZy3T2ptN+9S/ucB8/FW8gTm6m34zJ6YzI6QO/x3mla5z
G9mFZTGKGf/yEisn+ic01mfdP6fzzzQdqdWg84tkfMftIJ1PViNcz4zBu514qWDV
`protect END_PROTECTED
