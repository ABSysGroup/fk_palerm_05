`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mEaVfSof4o9XABeDydqw5PjEyNww9s2t8xfCL4pNXnZ8UeEo+49bsunLsQRmVY1U
AN1b+nsiVnzW4iYBjBkYLbhFeCz21Wvf2xrp5pl5WnDQR2GxWLYEP28aaVPQKCRC
5NEx7Ar4EatioKvyMovD8u+kd+EZQO9FmwASsnJAKzlTMgJFO050FmE1rSTr6trn
pd339/QdvlJwD83sb65kJJyCd/lP5y1EQG16DSfp1u13vJhhRiC5K25QLg6Ipnnf
G631FWObtVZTqvLcp365hiOffAietIje8bwIQYTdZbh1IamHO5cb+A/538pGfA9S
mFPQsIxP0oCX13QFVNu0Dm/lOSmv0S13iqVNDMzUrr5Mv3i/UEQRdLMqMaQIyr5s
GiYb1scjAxrx7102t65JiK77LLE5rtR8sHaHdJ+GWp/KRHy+FhyEB2PRmHC7w+Kn
FOsIi52p5WGgbCSlQo+M3zgXKtovnujDbjAX9UrjWYk=
`protect END_PROTECTED
