`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EQLRO4iFRAYy+hQHyVmqk1VVlC93gNhultzPPL+KW3CYbUcYqjImOVJuPzJEPDJW
+ET2lc1uSCeNYavki1sROXHepGY+VY9sMq2mt37SFC1eYp9mMu44ybZwj3/0T8To
vgZCuRikHF2iI63BIfwBZL1+S0hmM3C/8jJaUArkcuBUytufX9DN8u9YmfWKbNLY
9asZlvsQv5wcGsrIHL9OqeF80Xnp+4iwgE9iF0cCEkARBWo4yCrdZTcja8UfQTdh
mCJQCsuZen9kWmo1cVxzmQ==
`protect END_PROTECTED
