`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GmD9nTk2h3BkkatzZMqahB+efL8woOmc9giM0oTSn/oluYHUmJZTRqmop4ZdtCMN
ntR82McqWh3+UIvOToqOeANGGK+Mxds3J1Qc13ehfM7QyCXSlnFUizIFpfMqBSvL
6WoekYY4pGK1uo5rULA+OwZoDiuMmvxaMxbOlv3HCz5uq4l4fUBZ4jiU8Aicqc5g
RRTD+HmjLa++luV+xmPqlqZtj74qkFs2f52fRKmnp0+gSxoMUKgKT155bW+Bj8Yn
+vyy9FCBKuTrvHTXIvbUpgYA6TfL1aOzFx2l5nosH5/fjttd5UwImOmMl+5bZRgV
S+QezjLZq2ONmeWqdCnpXg==
`protect END_PROTECTED
