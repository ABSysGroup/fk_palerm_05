`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U0ayoWzPiv9bF2+8ufx+JIviwThIb+X2cAJ4iEEWku4XZXEeXqiWmlyQQ3bz5SqP
IIJg5xzrXrEPUhvsNoM7EavH0xoKTdNsEIu8b3ev6SK5k9bUrlm6s/FuuCM5u5xt
zpIeUFEqpDNjkh7BrGBlMpeZDXb3SfT5sbyH8vLavpRDpAKWmopIc24hZUpiITMy
nr5yRzJxgwZ5tahT+dzyi1HiSyQVnBB3No1Fzgt4xVySPWOzcnRriynOwxjoqdDJ
QZiDm1MSRLRb31d1JyFXPlpakO4wSxaFg8LI0+YCBINrXzapYIgtPasyhVFPzJX+
6wxW5AqfI+mqv+hDpBhUSwnp6fdVjN4eyYGaD7qMQbZ0XNM6Jb5Q7vOzcKxlRzUy
JCCxHKNBhg0hyiEnEJFDiEiDXdi9hUCQf/1a8dI4pZmzcbHIPSYzyUGPLKvCieb9
`protect END_PROTECTED
