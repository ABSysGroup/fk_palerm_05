`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fNs7Pb4c3d84X4YUtrrd6t8babKAPMgnsFxsA8jnh6BY5TPQF8J4h3IpFwO7ibiq
3HqJdGKJVucOdpvcBdzc3YOadV2WXJ9c3EcBZD/4LLpXqJy4Km4GbzdPAr85SaJJ
pdAHmH0PKSbZAGpiZ58PlS7XoNWpa1SsigxmVwg5nbD805Zp0s7bKl3kuF2Hp5ua
tSqdbVwCN/yKUOLPKqmH7+NCnBHhA+D0lPkcWhWUUMMtVPlGRgJC9OgaFZtVc6e4
aR/5pfuE4tXOumze1/Ke0rwJL0ehbSvKqjOTbt9bzJR0x6brfIB4ah+hA1EZD8h4
wcfO87gYf7mhHkyZi/eXNSHxaWsuvqmYOoR+zk4QNFW1pzt2Cc5OgyIMElV2Mpmc
lpN2ZnyY7nqy3Qywk8L/0dEkZ4bKbBT3qOJkbRdSUuBEcr+63B1ULfhqjf+S03TK
cZgIlErs3uGIq3ASSGqOaLO/Kv02HpWvyQCZU5Fpu2pLwSa4gWcvs2aXdRqZNwNZ
`protect END_PROTECTED
