`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZSqPCzfzBm/ixikYXHQT/j1sIhPjEYftm4hdQIsYisKBE/IWuBr6RcvT8SmT3jbZ
h/A1RFu1x5nCweChq2HrgAnMyETpRk3HVUrZfUpHfw/AAE8IBfUJgBx8phPHfQQE
FudthK8/1S5xJikuOYqIlwQT5Npq+46lCqGCB8ITLISf2lD2HGqju189NT/ZgTZI
ukEW4aQbyzw7f+rsOFYvy6kHv8oTR+SoMsGwa5ue366KjW0acmj1f8TPRmV7agK6
SUa65kicIJwXPdkDjYlpXcIuf0/7zRLN/fnOYQ9xWXxoVdOdOxzQ1UzKgbNXcyuG
USq7dTH3j4A3uoPNwCh7z2iGnE+R7d0OTetB2GZe7JEwCvwFY40koZS9aYl9J96B
I9GPOB5OinVL8wutxlGnuxC231KyQYuoIn+j5DDDeQzHMtAPsHH9VDeXtNcnzDP0
H6o31kW/hF39g3LT8R20VpHE62RLZtITbuDd892q8TcKHojnx8cNWET3H5UcbSk3
LsRyeYw6QT5YFimYTsfMdFS2EmvjPyqXwUJS1iD4N3Z5Js27jzbkvrgAO0wzTUB6
bNawcMIb6Ll/+FozFnuQAzZcuB5wioa7DTRUiBzZzNLGaGe+e3P3lytaz5cvDtgs
P492IZMqds9XP7CWu3vJ6ebTvEP5eRaqgqcgbcTjRlQp4VloPg2v9Eo0EjyzEzl5
G3ofpbvd1kSIx+g/3mX63HA2xNHEeCDmabIFZZYnML9lXK07R8ZekcKTv6aJr4SO
cjvdf2Y6vfF6sZEeBT3MXFkVs07iLuzwKO+J6oxq6p7WuBfbBoIJgwxxfTvePyJJ
dkkvJs+e+gIPe2kC4PkjoSt4HKp2wtXtpR00wVZfDHM3eDELGkk+k8jXU1IMT8hd
`protect END_PROTECTED
