`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fkrDeNsqqBGuMxNaC+NgNmIhPHD9LJeNOSsOxYBl0QP1qULz0FoOGp6vZFe8qDma
QKuCARkk1xyvsvCrwUIbSNadJlc8TooKeLZARdqWi7dbTMkRWZuK/beNAYe+KjlQ
NrXKHnHSp2rYX4N3lQi6UvzgY3HOcxSdkLmr5vXnZWjBQMP6oneJ3TPevxAA4sWk
vTlClD2weEkkcg/1C1mN1kZlLdMp4jIZBZ/VaLBanc3WZFirsceTuSu+W+AAUWxb
sSY3Ie/KgRdCFDFf+XYL4t56KrhX4GB44AzU7+j/AeO09lCRL8ZfezWoTB5VJnjI
iS4twbRBzZTJ0j2rkk3UwMUq4CO8kHNq5M5b8gMOXtH7AV0OmOi/ShSX+Gm6+tdu
RZdUIQ4AUejM/Xt3amKJcpUECPkxjWAuBheSkoEuA9OgN2fdwYmY8cVRTLW1Ove7
j8a+oWwkseTvgYgipo4VsZ/8u4BitPh7/YZBjcssQXtohk8GpLUK0uPs+0gLMWch
3UhglCnhIJUzsRniNbVAawki55IjbeJWzrLUuC3F/gyeqSg77/qd/broCPTmiIGx
IivE8fx2zJl4RrTPcuIL80Elzec/dlxqb8FvsKQENA9ngPk76SaGvfArSlx4/kkv
92ZUbxgSf4wNGitRJZ0H3wkc9LfJ0jMtXN9T1qIHmvX9SpDnveUHqOMjJXutmRqV
ZOo+NI0eer4u/h5CPFvKLfsoR9zOhTRsSiFxUdD4C4ZrIQ392KlCVNuC4nssTMY4
B+bVtK/XCCp7ctxHyzq4PL5Ou1A58DDHbFECzMjliqfgjDAuJ2Exs3B/qIsbige9
DqU4cXejUpPx9j0n6NalQYPmzrw6xPmoSBI53TBgA/8jWHLFQ7xdSgC3vvTByqf0
GAnkirBoF4vzsYtgrSVa4IBTUGiOcuH06jvJK/aU0/dUguv2mvmfWL6TV7H66ZC2
dLLI3IQTPD4oFVZLb9qfwlmIGJCewSrWtEeWYdgfrCe42JTFm27A4hn+Q9m26EdS
GEsVEdFISoT1YwecNFQZaaDfzAhVP7fzRqnh/FjBl7uag9oLYhP4GVMjCyXsA98g
IaraAGD0WCOkVeW03wF6bpBN2k3G4hsDEDYxVRP/DRQyvHq7PC17GN2kqWEzV+jk
iGcunYJDZutXDZ3sKcwcmhKCNvJvhffVmIpKMc1Kl8E=
`protect END_PROTECTED
