`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c0yGmBxQiYB4LjFN3BC2PRUMqCXyF6JB+SBgEi9tBjzHTKwCbvEAE/WhSrHNVLlM
B8G25qwhkFFvu71udrLFHu07JHcMUebSQujj9ydB+3wm2TRCpPfJZ4fUis7Kf/02
darAJX6mnmJt2QpzzLXJP7uyDQp8A/tp42h/pWqTt/c25e6w7Zz7FtLZrc1gEPPv
yo/mnym6NURh5ZPSrjdjtsDI45iKnj64mx2z/6BedFzZp+ouX2trakjwiUV3hEra
VneXkWN5KdOrDbOJClGYh6hSKWVqFenb+dfn7D3ToRb7iexKWBQbsjebLyILc8Uh
xFrVOVx5pIn5ZwJsLoABvLefmLDSwYTr0eCKpSUbl7L6C8/UV+OhJ5UplbRD9oBj
Bv7QwFxODBpMkfaDPRjRt4NCjN+qLvoQgBpy3Cd2bAa/FSp9Y5JAcXCuOEkM5r4N
LFdL8sT28ua5g8q8mNmx6FUeH4oCxwf4kKDn9G8AX0yjDGaBJyPvAkf+2GoJ5Dk6
iCU6YcMYNNQkceodm/wKuqGXH1E3NYnh8OLrqfmjwpEKRbTCBBVLq/Wk0zNFUKaa
pIFe5Kv5DJWcYCU90u7r6nc3bDOChv8dPqgbfO4g4pbpX7sKhXFMo1pP2oIzPblX
CZ+ADD6TV+41dP14yN08bgATeFrysp6F8XYknSumDt3e04WCUs1TouIMp1FOs6O8
XV1T8Zli3AEHP75Ktvz9TC2HAEARedmDHugqmqLcTpK4rBwenNfGK2h4M2IwRHtY
2IhknHGv7EuGYnUuFPYP4Y5cWMN1Mg2FOlcMk6zTTxAxFGLJr884u/MrbkF+rIl9
OX1wC9RAQjWodf/i3HcBQPdsSF1gsx2e85wxJG0E0I2KEPO9rrsTocReIhAd34gQ
kLG2VDVyH7MWq7mHbg8oRODxpNR4NBLnp0pl2ll8WbWc7gKbx6RsSjsajjSpQYlS
qjyPdrRm87LTKpjM+9NpQEEmchIl3EuzNo4RczwMWsv63WijOl+J1vq7FiwT18h+
RiEFFDGqvtj0IpeqZtRIxUyuPnyWGZwqAf0Ur5igcgnELrtW8DFq4WE5hPhuf5nd
v2bRARj1Y5tnlufP5CKqB9s+7l445qpXpvNq/IOBtZ7Tzng0tO+8Y5h0Cf7UR40C
3PIiXkXFwFI6MuV+GE0EkSxwPQR26cnmvf+0LjZQaPJRAhOsmVXcCPrnX30CwleS
g8AWg9L+gvWoMj9QPCzNXYOWHcSc2x9Ibf23VL1zJzPHMngvXU1udcCWjkAy6H9/
4kc5yyKHJUIEoSlWuCb5spfPXeKuTliGe4TIgOWEb4xk6NDxuUkwGqAudgcSnuxu
UQVSTNO4l/gb8o4C/s2gN5/I74Mq1VnG4BrYYj6MyqHci4VIKLnaY7myyjnJe00y
k0XkgB2234tpqRHzwQwcB72+DFMv6J4M6uaPZm2SVREyg3x3c5hqh0sSz5ZvWIpN
mpUE30WBxbey8OqJbvDCeUoxiYGWk0TX0vCZJSAujCYhoMzZ1quZiikfx+dCWL3f
nSitAr6iF1u/uKNzxqYTG5iiWH4Z80ZVPyTke3lDV/irFxICvAI0+PA1KM9ni4yF
IWgDlxbZJ0xOz9izj4DpTQ==
`protect END_PROTECTED
