`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LjSvtP2xToPexzOyD38stwCO4QEq9GElcrNwHb0rP7TYoge9ZT8kIXsLgQ9gkDhc
VYjzQRSO8q2DuM6w/i3tCivXYPvPSuGOGXYr15AYLGLXZNmMaQrFHorfQzmt5NU+
7nHQwWHcfpzBGXPz3hl3vakuQeP1S8Jwvno0aFuLsnSSuZbficUAYsS2rCGP/cyd
2CNvJE6e4uvHIM5sfCMc3Vjs2xcp4LbLmNCCQLd6lS1Jw/6xPulUWxELUYn2IE8T
aol/KrJjx3A++VxTxK/C8lMxLVjvw5oNjUHeno7siNc=
`protect END_PROTECTED
