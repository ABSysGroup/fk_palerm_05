`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2cYplycSlVhoQz7BSw49K7ZvKGpkU2c9bgmQlKw5U6PatVZnx0UCzZNnAY7wBqKt
Ne61+1jA95T4FoJGHEcI2NZuUvGZf1O8iQxCCRLE/x6LEiDI4yXd2Mp/kB+sFDsF
2DEK1PjfVkrJ654Wnr0fJSFwg84fQfcY3XazPilc5EXImpI59CuJPmMkVsbekEXn
M9QLaQiI+oq7pZiacpfddmT+X7XaoiI902/51HNaTv6BJ4Yb04Ek1qo9RsMiuxS8
oGNPNb/LMQ5hr+JbfEh16xTaqBNhKblGn33KMFl3ckUYwVFK2ruaOC+E0k4yDbjs
ef/wW6JfUnIM5s/te6y0L2Tt6DyTAw+8WvcCsDYDVTgGVIjCVllHFt0dygEquy51
txQh+MpzIy4GDl+I8fbyjufCLXpO545ivF6YC8AwqBQYHPM/bfcKHtIqR8UA39zY
`protect END_PROTECTED
