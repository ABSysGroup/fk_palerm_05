`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hVueciCmV3U41P/wPPVXZ6e6ke9lze+Tr1Keo8RA2313vIMmY4qUdndscE9MS7Mh
tsy1I6bKNZDuty+hc4iB5O1cl2aJdoRt+k8qD1FCKaCaUs/eSWZG9Tw0a7wo/L/L
rxArvsqxSEOFNOp5ri7asEh5OATujvgOp2hGMotOFfwXCs/HH4s2QSsgJk7+/eNm
ZTti9sbbKsRx6SB5+8crW/n3dvdBeQq/PY9MRn8qPT9HFUUoCMNcsNQ9wCO1GvCE
dj7UzkgRv84JPKrlNr2vgVGpA9si8g4dExCywT9Vme+fmnSht+18UFHn1l7tFjHN
nKh3w1OcoKELLrJSiKWwj/hXKRv6ND1fssjLJ0m6yUoz1efXLmO9rMxnN2Fiag9s
Sqm/XnTWlT3j8rzHi0KwWZoRL/eCTJvLHIsRtaLqrG4P990vYFxaDFyCPsNXVwr2
XE4Xzezi3COxzHzsAKpABVm0KRGUIPOT/WEdrTf0GDSvjQQC20mnuazD7Q9Uj3ub
BF1fSeU2JAwTCRHZW7OIE0561/BiHQ5GdiUA6w8J1HJzEA5xSdVvitjERAj8WQ1k
m1fySFXY7dYnvitddJiXlwgfNLeONxZoObkQuvEYX9ygzOF0RDaK3S7tr07YIaGx
+CScQjwD/iXgWCK9Mo/rYFaH7caPNjxqBaNP2GdOpdOHdXoDNFM4xEK1IPLaG7ut
lnY35QDDE+r69I7s2zmlxx8CXVruv1F7WQVxRQN7raUIl3e7cQSuZugHQ2qdGaVt
57r1O8YSdbBwjMJy/AEfaoSBoJrKV7o/BYQ6ZprW6vvBC/ij0xRc++2QyvPrUehK
/aoofGFNO2NJwPk1iYuxd/6kSgD8HNHjxYXGbDqcyDU7ykh2+M7LtpjwvYA0b7f6
V7WsA0Ua3Kk15hVWofpu5wvITOsl1WwfR2FKWQO3UwfckSXXJOLKVgi2XswTPo35
ruVwSVeoi951VrUQzrtDqdieJVeopw8TGrWaigC15+yXQqHNT1jR4dVEsHhFskWP
pEIPvS3e6HntXGvRqdT5drcoljQUT/+7IysKCIaPt5T6YRFkat6EXC7PpuvHEdtS
97bwzXqC2I0nDeIY1nSL8Gn4oK9MK0EI+ZvCpPPJJRPqstGJRHWGyw1gkemzPVky
v983Ng8ggEj8VFRw6R+bd9Qur+/8MVUDJeKXlXhOOBEJHIH4/pfyJ4tr0qyKSqM2
z1hIiX0wamGfw5tWu1wcu3fiPorgUDlcoBjJTIsd3XJvgFHOR9/X5YVsfUZiqufa
8E9jsDeo+T/Mj3/opDfgSAodfiXFYTMOC+Foo2VST3IkEvgG4n4rQEoMezfTfltZ
o/jNdX28ysguO0SICizj2WeRcSegWENmGO9V3AJSM4ZpLF9swCvd7YZMQdD+KrMf
8CM8yeVTczJyf5DaS+yO0+/l7LtHQPe3Jme77lxIW6d7Rjvvkb6KSyE4u/5eX+CL
VmNcwNrthvHXTBa70CLumLlJBlKq6Z5t8Juyuax9PBlMRivkwB1h+sANeyAq61Bl
6ktR86YqM8i7mIuhP/vO6C3eC2FJOI0aGP+go85Y/C8fGLJBJuVev1D3Qck6PJNc
nGplGjyQA/lYShEp7EPcaMgPcxvaP19ruBggWuYYiWUkvEkOd7GPwAtagO5KCeKd
i5SvF36AVemXBJVYM1wyQkQ1twILydQ1IfzaWdisnxAubWIXMaRdsjmIYYF09CTJ
gVojy2JyNtgFK/3lP848KmtJb68fnrWFI2gjcJnxcq/ohPmBLShhClx/RuIKaJUj
imTn5IqhtxfbSuKoLI5CTLZkh4BAQAq/FWCbCLsQWI4ZY/Lj4K9samsMYh4L04TY
qSlbwB+tR0U/6aFoCg2IpeCnnx4/5+Hk0uo9s9kp42+3b0HW4LGyj9OshTzOv75c
sQ40P15rTEuB0+d3kFjTv8p4kv98BOYAB1KWZ6svL7mcBPfvBUnR9ut7UHuOTK9I
Wc9nxqOXBL4vU+BWb+/QssdMg8tjvuakDahQ8RllaTMaMmOHxym23jeUV00mZxPg
xReOcdx6ndzuibWKL3oVjlxrTUVw4r3beRTgh4jtw4aNjdB9BZvH/PxZHERRoRDn
5QSeIjQ0RNZNrnICTEMaPA/XfqRzv8fESBBxbxrgarIKVGl/5Rgz/bS+UAffZkED
+/8MPG2eMrdvwI2EXIkvleNETRPjC7W25qi9WkahdLQto71AqbfR67FxE3U5O104
3op8xV32KImsh/EyeKIHHsL41Tc1uzKTkdjWQ0+TJM4+iRa7imae3MNiVCXKMLrq
kV4BPJ0FAkl5di8+mK70n0BOfd32GTpSlh+JiZsxTpnzJn+AupnKd6DsqKf0SmEL
s/C61NPnm8MLf8zOdl1fbWHtpSZ3ht2JSW8oHLRkMndP8RODZRy0VVTVEmeRNCWH
IcKjpbFDrvJceyeXDjO90rnPNfQCMnYzUB+wZ4oYlp+8U/4mIM2zZ7fyHpGMLgCt
UuFXBpliLwYnFmYmostVbhU1Il3m6xbUOZk+LRo4aKnIvm6xo/viErUaTS6iKa8X
AHoe9Dbvz4ndAsBknIs4jPC3Qnhu+bLbZWgo7pIknwjoKCy8L+i/yzVWCoyOa/K6
KCG47fVMokv0dAM3nr9qBir5F1Qh5Eo2VJvYvBpaX0m5TuniqLNVBHxQEJtBvER9
E8bjRoiSK62nDb88cTpvsmzrzwF9YUXznwDw/x7rTdlwcJs8QK8GJncxi+56sawN
KHcZlQQjXpq1KjZ4izDZS4JpzfiBsMZqfyqmgYOmjoyWWrXxc8/XylT2CYIoDnm+
X0WO8+cNaE8xoNBGiRwti6rqlIZh9VdqIc2+IMg37mG9LBdWJYvR3AhaWHHOo/EL
ptXblVRlboUcprUFWfIElFpHDPU+DcQ3/U0Gq7HZYbQe6aJmqVOrbMfEAqVAQqGx
hohtcrmkzmwsjEouCgZcAy+/mEEUPln01MbUc6HDoB/yfrYH1IUis5WZLqI6WxtN
vJXeJt9Yw6W17PSQ6HL2yjg1nxfM8WcaTGI1Byjn78slu8XgKE0zBkdAqHlh0db8
lEL0BGDQtmfcmC2SGm5mm82bII/JN2k8EIrMehSHl2ZS+9LVwQyvuuUCO87hdftp
C7Q4aWkr5vU8glp+3MwJrkLLURGW6l1grN8acDb3oSTzCNkETUiH/1bTvofkdT2s
YAn6RlODun9pY6Aj5qk2aS7EVO/5CxYf5yB3uPJcDQjHYT6kuyPR3DFRweEnrdxc
o2p4K4DTHlSMG6m6RkGad0BWFNR4q0hsxZsZR5W5HOz7mYu3b6xsuV8pWvg809HY
mx30HX6Dhb7d6cW7qYtX3fg6+aPw7QChyJBEl+1sxqWzYrRH7VrFd2khcUF6JVK8
iVs1Mx+8hPJxcEAnn2iHK+tdRBDRc9u4pLYWnK4nADRtkzLtW8RohMBsB75No/XL
fq36gWtNpdbpHTp0IJNuskfdaVunYMln2AshiFUpLWDGM+A/CoWv1fB8jdMjcPrJ
e1CeCP+v/S3EWrr5B9boA13qlSF0SzO+i2GGGwUCGDcKFbOhoEiY0yLNTYb9QLik
RqES3kd6FpNMf1OCDtd0InH3kL1xbWiUiUQmHX7AhrQnNZYhPh08yyoh/YnO8kGY
4wHRiAcxFqpXzWFRgicc24G4hVIGIZA1XkQBzRmGWkWTDf/6lvgsi4n6NlkgkT/K
qVMDVi3lV7fwyEQAVOyNOPvXailoEayY0G5XcRlQMl4zm+CHAmpeUevLbA4IIjlY
4OOM0BYm1ODlz36cC18VSVpP0XCN2/dB1lGLXyMljvRA/WpdFjPBxV5YCtDF/TIn
puGdoEOL3XZ+/4VS7WkSOriNYrk0KEvA6mxV0zhdzau1S0XaKLjoEXyhPuibBGLz
RR50u5WMXqrfFbiio9+sc+sRh7rp0eErafHZQJSFaHqXRgH6O4pXfyizvNjH9sLJ
wGi3j5dK04xa+AGacFY6OWUgyhTg9N/6pexDnUU2Cv9ztX4rojv09e2hx+K6wG/k
a7xSqwa0IZXme4r3E9vzU/XdvSN9fVV+XCeps3TMCT3K4f6/m9MllxxDC4a2Y+S9
rxwtxFvnyEfQWPcuJwjQhukpjAgY5qmNNhUGYPb/O9+Ubj5XzkAbEQMbNbOWNasH
4Kigzsil3RnA6xoaMAZsWiY9iYyxk9/qXWufViWc1oX7d1PnuH5jUOIrCyaCRYS+
KZSuAj+xlp84QQQSXJjAjVsMhePfQhPvBq224BeF1cmgT/gYKYbQC9hQXid6mZvN
+Q78OEUJ9oF4uXTtxcktaQHqSH/5GaFEVR4ZMLKo7YaFPcb7zSCXvNhhv4zx9PYP
5bfcz6s9kLx4RH/AqXvGT+yDsZaP5T9gabB0vG+HERRpiIGpDXD0WdReSqRBpU1R
EZDSLDz3Kre4AXNoPs4PMSVugGFtC9zgixpASqh6kiUfeRDjjAmtbtw8UAeYQI7H
RdzpM5klnNDDYhFGUd9JwhMph8Q1WwLQ/6a5eWKIBxY2ERnOGuYDDWmM5Rpk5cYY
cXVfSj4gMuvotVfCpUpnD8K6GcgV88RlbfGwvPUvhBPERfL6n10ZN+b++O1x7MAf
fFnZ+/TnIPus1LDFJ4pe/D68ErWjFmQRJ79Ci6ncQbMJTLM6KPk7WUlrrIyEuSVV
qk+Pa3RGCp8OdVmDVld7npHy1fhR56UObhM1VRvjVIlmGtWQW0AHfIyw8ErvC5yZ
1ECfyHO0/cTIMXfsrxPFJJswXv851YCJ3aE7LwUf6tpuv5uXlyxLta14E8KryC+l
cX+OeEu/goet3Trma8SG2r2HecZA4HwoTqfThVF5i/AIr72WjOnRRWsjU6E4eKut
7bhc56phpZ7LEY1TApPOiR6wDfvkoSZ4J74tTBDp5K4sn+0xKiMAv6o/CxR4SP3n
O+aa0l/E8x3sb3XDzN/wMxdzTWfXPUkmG53nNSjJmspbMUUnPS7NJJQtj7dSBkej
QtUFI2kK0I02dtpIMWNU/wR75FESsP6IOjnqozpn/u7sEAWIi6HXOaNTr8N3MqDy
96Ew/AACw/VZ6DVpEkEgopMS+zxCUHn84Y0w+85GxVE=
`protect END_PROTECTED
