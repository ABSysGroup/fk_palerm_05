`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zm+qRT58cHHIkgOm8/yeJRte6kllOrwyFst94PgoInI46H4xn/Y3tcXNjYXmSnhE
GhBo2Gnz4drWGCyJkKR/nBi6zGEURF2Ofpl4gfJzbAujDZQsFK2Jw7GUh0sgDjON
9k0Cw/sc6q6wZlzhQDTwUx6jofAleyr1IpF+ANOynYw6sKrje7O0gCxDSVu9yOxC
tSpQDVUAd3F/ZvSijLIof7A+yN1x9L9lsZHnUO9VWP1alSzYzJHK9GIA6NgofdQ4
Glo0um8VaXYjqqh3YDZjNhliXm3b+8WY6WbMaUtdyhU=
`protect END_PROTECTED
