`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J/jJW1AZPZ9uXeHkyBzjwQhWxBK92Kzu1yUXK2HmWbR9OMlK1TfxRq0M1VIpFE4v
Hk+JRGVhPey+H2g9pnRAL1Fk3CL3phLPO0h8+i0ta4pGDqJFT57xUWkhJI89KjDG
qnCT859RhuD0ep+nSAnS3NB2OtmsYSj2h2HY1iYnVMaRocOwlOfBzDRRFtWX3JFH
EHUbtyBSwI0aI82lYS8XOnqWDKetvQ5qN45VW55VEVXGYnmLZjGEZdLpFZFs6Zm/
`protect END_PROTECTED
