`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sCDVJfekBwSRsykk3xDfVObzicbcYQVdBmfIy3KKAKBujgetCT5457FnkXIvDrdR
+WL3eIxnIVgQ9yRdZHBM4ocH6XZkHZjZ8sA9wjsCHOr7DYXKc4tCiKRzi1SxnF/o
QTqWtSdZPb/O+3sCSRmW9U/jEtVS0lTXEeM07OZZHDmEQn6smYDWEfveverCzp3L
EuQ53LOyCVoGoyFdIFS1dnpiVfU3pzqfLOZouTbd1dr6pOYd0s0JTxned6RwzpUG
e+qWH1YvCsoGepEB2F9g1jX+R1aFkPrCOwFq1dwN8FYkQ0F1J6LYTEMJGokl07cI
NjSGujzamHl/nTlQeakxNoGPG4Y5ikYkj1boCoXDvCXITZkWaZpN6M31nF6rrHAl
Ab8AKcrK77npmgkpbXZxGDyOrcqt8Wm2q/7KWYtjnJ7xaDkrU52CuYjPeMAinsNR
l0+9GiNYBh86Jn3K+xo540l0oa3bECs6RmdwPTGjGBuYBinLJ7vGbyyhzwqx7j+e
I1S2azl/EJ1UGKEYBX3CTlgpx2OOWDhp3/nCKznWzopSaYOAtyXZ7KklKjx9f0hA
UjiKnV4ADKIvW4BBwirFRg==
`protect END_PROTECTED
