`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DIrSSZebjCeMut/GsEOw57k2yJ5gsO+1wsFdQSCfT0348D0z6B4M+6tF9UlsL5M1
fB53d/Gss1aO2l1r7G9DE1WqnCDnyXub8rQK0pyX0D65clCqqrCMZobl6DkaTGwY
HHBEt9U8eQMQx7gIQKecmB0QRbpyWIfV0mmBinKYpi0PkYdimoxu44d1lNAEt1tg
7wRmD3lul1vXqZrRJfffc9s/zQfIFPh7KYJBanjrk7QqD1o9xvqcw5rOuON8GhT2
M7HvUlg4lLhuDtzMK6AsZa/8B2VJuPPDturYPMcQB+H2jvaJlsfAu9E9+Z9PBmBX
s+EaebD3s7t1dHhnqytPz/KGb9JKN7WmAT7p5xoshez+JRhh/Hk8kjJYFo+1KBLj
lyOUnxsEHCUZe418qGa1XVJb8sAXbPMELaiJa/N++27pVvrXQjKbeHl3Ub/TIaAj
3kuPD5Ndt/Zm1bHREebH/aPvQTGEJhLQ4GBT/fbs2v9TvqoxfCckj0RPffoiCmRj
qaHllU+GFUDp9GciQtYc4VgksUPfat7QleGUo2ZdoaYq0RW6UPEE7uc/AJSI2I/H
jeWp3vke3gDau18qlEc6V+jzlulDoNxVPKIUQYoNOZU4LWpb3/eSIM370bDDLYap
aL0noarjULbvalOtbKSTG2lN6XKWSGCaI+QzDEjRiAWOlyKAcCQeB6WCwaKnhiIk
RIrn0iToOxOmvW1uXEvSbA==
`protect END_PROTECTED
