`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OIZ7iIPiGQO9QqN2NTp2/oNvy4vtEAojIO16NM6G3riV1aSVs1PwKy6a1AF3LPbS
HYRUvmU6NSc3Ex38ecaPTtAMrfMmz89dx29GUYT6sAv0CiU1+ybm25N/dxri1gkc
OX3js5XVHj+l+NQmpBtp0mob5TAfkDv/L+1VeIPltthysMVwvyNAX0NXC4vu97f3
jvC7u8cL4Ofy8iVU8CQmG+rNyff9Zy+tER8teyw+eqVxG3wdDI7vI71fSf2gLgp0
sMBi4hEPM+DSedYmMV1A+3zYOmcRVSn3ZjF7pgJYuxLb5osfPR3xXI6OMWoliW7W
W6mAP2GI6zo7XM5AzYrRhmsPusOIs7A5JwWO5//ZXQu+Ju7vbpsfTdBZtXvWYqvJ
bz8lFoz8ZeR73XUXs6slxrW2QXTVBd827TQsOhzYI8y9T6AHqSBJKG32BX4JkBZV
6H38uNwFWm1UQrUkC/wiSk12hElzpgrI4Q4Fm7Q/sFzAPZLYQOxJYzf7xjIEh2su
c30T48fUFWysxSH00iDzAFRK6wyQI9BcP6AoFkSocVWukCh20OQi2eKyKCiOBmCL
ot8Y+Yq4zkaB2E0aWiQlwNY3n1EGqRUo7mMt16sYukLNkzAfYQVyTCGlnInw2+nY
x7vqLoUKSJAvnm3NW5VUkyfqNgoEbL+MxRvslgpb7LFB1yW3xgxdNbMQqlBLoTUI
PQEw9hilqOvTYP0ehN5ChqGGaEyLC8KrG1bGKkBi/p5nWd3B/r6neHDh8KkKF8sS
KQTaj2MaXVrZmba2W8q8eb4cFOioUwwS2u35Rj7uucupuokWdCHy4/D0gb2hhdE6
tY85fm0dD+O4ViN2Fl/JkLrW26d1G1T2PbkeUq58cXX+dh/wKg9gKEJ1562tTqd1
7bwmqiHJRCnqMjJMFxSoaAs0OZW5Zmyp/EM9e7BuNymSn9kNROA0ixXo+3q9oKYR
4GdH0T7MuBJk02osVEZqJ1hr6ZP7emVDsL8s53bRi/9WPgXy16dY9a2UeQs6W1a9
+2l82SgqpiSc4KMPStsZH3T+/llcgkpHnQ7Eqd+RJ851xQLPdsHpfVnUSGaoyqto
+FS8gX1H8ozCJgUgYmpfxdxEmg2jyf8hWpGoFXvvkLU+yirL4fTox0tcnEIYuFEF
V0YBi1KIPRgH2gt8R/XIwHMuDQNR4OGvHgNFPHDVA/afGIwW10OcnUpsLlJmuJzO
BCDGMoszD9C2/RmJ6eMMXTNv3vVjxjdZm9KvAjvKUeWNhKiiwg0XNAFCD2fRERMd
t9hZU+PsSmTMYD0mJUC5DWPSGCMoCCmBLfb2YMhkrf+DGcPM8/6L0/AJ14ate9lT
dC5Zj/n4pJVutqDvMg392V0zjNXAcAkKGGBqHxw8NVnZqeOGkbWjL0GrntcCE/av
ZJr+U3MZc9n99Cd+r3eOzQ==
`protect END_PROTECTED
