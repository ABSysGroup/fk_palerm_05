`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rxwYPqngcKQWaBhYoXH3Kbvg8YbvYECKMWR8HfuMM/Zv2NN9FZvHO0EXwEJLNOg6
LYoeQxnXtnK3R4Wi/nC873gVFTlEBh4n9Y/pqHxdx5bWmr9T9teMfp+lQ6DWjowB
9zQadNlA73Iw+0tBCUHCACJxHhGmpjzs5RlL71Owc0/N6vGiAOPLMvOXkLRm6R3T
ga0VFhN0PpijFWFmjdhN01yU+6tme0ekg8g6629x4ydSVIsHWSVyVH6NviMCR3Oa
U4V7tXuht1+3Wd+F0QHMeYrztyVJ/SURBQOZK5ear6E8KiUBB365lDtPrln+ZOG8
hThp39uzfbUziJGlG7OccTbZArMdBeyHMHocstp2hKTf/IjWLxsC8FCTdj9LBVWk
WpnfDBW5lWAreg35sZgs/swacQhjtFlrJqYRE6I7z9p6TlB3eSjUOUvpGriCZcqW
hXhefgSRYEOZ9ZIDiYgdIhyM29JiY8WPxxmsj/7ngxDNwO6A3QFuCmMxXm8Bm/Ke
nVHN2ajdjP20zap4vsbUJ+l4UZOSCfMnE/cZOxqFJfmPHdXvNl/11CwVuTYounGL
SeKXidghBhS55K0s9OfXoKYmgSTkTotj/TsoXN7IebJXvJ3NziUqdVgDS69SJHB7
oknu2I/Pu03JEm5jheg3gU+RdDPk1kN4gUqq45jTnLYLv17T4WhILuL7jX+B+LB7
W4RMA/nFRz5ZVSuGBhNs2PphdS0eC0lcDRDcnLBSlCeGBuC/ikyb3X97MQavE78G
d9knqYjC+KFwX4Jj/nW8hDSlAoH59GsxLtVlIBT9FTT8Fs0LeYgaea+IfhH8Cf4w
QKOERFWc6alXYvuGpWEPsIQq97BT6tPGwSp4Gc8gtE/1LztPB/g2d66CjS7JGJLo
w/zAayVt1puRE9DoMuTQ/EG1OHn4ze0ym8yFmXQ95hXS5XSVg59yulOAYP9yQ5eQ
rOCQryYpyR0DFFmTWAN15Ls40/fC9+0gWnBb6Rqh6mAzTROUY1xck1jLjAR9csG1
2/a44iOdLOEGJJ8YihimWvUx3e3HCT/Dq/dyBHe6u5/4HJrsRnaXehex2ynuy/Vl
lhw26FGYIe4tgVcDT9D2zngB77po2VfbpjcvYbQq7Lxn4SvXqT//m7emPuAGGJIi
6NVxy2cwuIBrF0BsWHT85Kpnx3/b67tiCdyQT82Ywy0=
`protect END_PROTECTED
