`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q2A6EtgabTBOtPR/QHj7w08tTGgPOG2g5VCl4/yensJDkiDcEuIBJg8wM1/uzVku
IUrCFmAlE4/Pri7RhqzJKqjpIDFoRgizKuSQT/rILq1zCCcwt+qYgZD8LDGrI+X1
3A3JEnehqm0fp3/sCYFWwNWsw3y/buxrkDjNjsqNte6gHu4BTajmbkwYof7pMCps
eWm2cHIz+l1lX4NzZ2d6pSeZT+dENphuVbELbJm9oRY548+WOhCc8BhUipz5e0T5
9vSk7ccXcz5z/Wp+2NoL+uvvul2i2Z6zgroxtZVXXvCmVOj8LjjIVluD1Ua20txu
0WMZV8pmeWuQLoBgkMaxMSF+CBZA79fguBQbV+FmYlNbWvJA+Y/WjxaOdys+8cyd
3vQeRdIs4VgfYegTsh8GZvLPaDwcOcTJkObLUmp6U+gq5iupQFpN9J4fsnD0ZVDe
5PuB+4uDFh5tEo6JMz8e/uVkubv2CHXu5nslMrTVbwlRziaPdkpxWLdb/MfNqAOg
KF5DxqB+GrjFioIapTDRnVOmy9YNvF8vqhNj3nxGs0hiwPEpsnUAHOwIRG41cMyN
rzDQhnpisBuKN1A4Ro8u8dBW+mrfai9N5/kVF/brq25THP1c3KbgZWwK9hBlcTw/
`protect END_PROTECTED
