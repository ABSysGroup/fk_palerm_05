`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UgRj3yv4gaS8gStHoNwLLEPxot3zAYzsrj2nBnUQ+E+6jWD1N2nCBapbUWVOKWih
wF4kHSv1YSYmI+VUSgr73tGRGCSRWxIWO9G4FcKcXEO5+jLfvNgRd7SFClpGPrqq
7odPCGUnweN60Cb8lRuexVdTq/IGikEmJn/dpHoCpOkrfdz/TXLGfuHNu0reozSR
keSkNcgni724f0e8Ihi5YV7vWKPESMedba+UStAd4aNAqQ62uc6lFqNsdd+JIg3v
n8iOhdGqBUAeh5U+AgQJijxKDMa1EZhfO2oXyZdmtktDqK1r7eXr1Jlt4jQtN83j
8UIBLOjqcAaW7PTqCjlXFZ/JB/RnxPv+0nurtMG3njJ4iUy9vwQqUdlZriVMuzYZ
kWG2sglV8UiGRY/h2rq/1CzXCs0nxXTxXFOug8X7G/2MasP2rD3rhpihKoJm7snO
dL697923od6Azzky1+EqKr9W5aFX6XoKwyH7nNRsVFJlfbX0M11umtImYaKGSlOE
mrPTtAuGTxwralx432omyGvwnAUK++ibj4D3WADm0FY=
`protect END_PROTECTED
