`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5+X/6sWA5IQlXcj6XEJV44jTsumkrBHOYVxF70QoTgF4MZ5h7DxQsEaFgACFwdP9
RueI9AYtQL0qHSWGV1blMw+oYvthi7Qbv7adahDHwo1JgBm3yzxEtOn7fWW59er2
2Y0Xx1FdlxVZazY6kSrC96UEOcxIsyuEIGsijsthsTtrBMM2v7ULETUx9MKr179b
G9ZQl+Drz7PxfTSXpdeKxg+vxQOyH3OWqjhAIQVTlyVYGOeTtYo0i9c2wox5wy4E
GsU9Y5vXGaBXT5SegWxDTzTpwCArZ1krngHJwh56u4LoQG29z5QUS7V7DOAa16FY
+T2Z2aQ/rCaBxcR1jlO+0kpKrHCoqRwUN7bCeXRcbE51eWYK3V9oVy3icfJElqA6
f6m2Bt3G0PRFwXRweaPHmwZSu95aLDfp9Jy/lVyIbdv3j8wbMhvH6UgMEXheu7Qw
Mh2cQHgiYZsGOQpXm58gvEMQOUGDESthN7sEZEGQJhPmU68ITMwop8PAwwBwI7+G
dSPl+3/ybv9fMmJ81+quly0C6z5brnRYOZ/CFeOdPKGhbC7yPZyQbYJsiTahSp/h
Zwz+ErmJPMW0O4MEBeAd2nFiIBLOg1wUPU67VvOGiRvm5QYJRzDviBR1vw7dwbmC
GwJZUicwQEhshUijXYAZnM5u5tCmrdL/J+j/GeMiF9U=
`protect END_PROTECTED
