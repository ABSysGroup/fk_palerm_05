`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mBMPZK0guX4+OyxgjqBqh/2uy/sGAk2imbwMCxhfX4wZFugspXmH/ytLWQ9x1H8T
6vJf5cskK0UTwJbccGyAJDoLHOXeWPLOvoGwFqHSZxZYEjUgbKWsS6wivrn1XrEU
zLAivFL5A5U/vavaBvj6VWcUCfOl7jpa/Ob2tPBNXbuez95yjU3eF9l6ScKm9pIE
oazntVvN6Dyik6OR6Sxzd8VEoWcJmyGxtYR2YQT5XLiVpOD8H/OWiUKGwrTLRhb8
LqRqHeORDlEs8h19dCXIr1TML55P6QSVMq3cM9481R0ZlE5NV9JSwlyii08j7Dqj
TgHIjZI+vm4obfjPDHXf7Ugy16ZH0TaxcIdPCHFsO+3gHtp0H2jo2L4qgNg/W4Uw
EJ7ZCbJQE7FtVJpgTKIqu9VlbBF/TGiZ1qrkfPhmJ98iF4dr8reyG8WjNXD95jMv
jLkmCoWfyUHKNeEh94wE9dUVg1vz5gHk7K4fCwjlY7B70lCCYZ6gyN5zdoENCNGx
qjishwhkM5eqe6ss8Pz2cl0ycd+wLI2CclRZMd9iLJkONncY1aCUceveWI3FC148
xzB+WPFdjaLcF1d3CXhYep9Jg9BrTG4UUNVHc1OPY07HkLmr+Rxwa816z44pgv6B
80TnVBuKdlWAA7UPwge0TGvGHgXK/Yh4HVUE+aBQpXSs8zgs8vGohSUV8oARDugO
UxeUqVZBHU3Vp/eReOfudzlJl+oUNn5YFFBzndyg/yT2HbKdVlL+asC6NYyxlCpR
ZXpyFm4L2XYIOIxfHUW9lvrR87DiwpaT4okUWXFgQiNRIrcmgkVP5orVGd7n9bI/
YAejIrzmbCq7vloYRjClyEq4Dhp9Pcz7+fvNhDV+6XLE+RBVgCHEae395O3e16v4
2O+jqdCJFHNkdl5N9Zgelbjl0niw7uW86AKvno2q+kJ4jDpG6F0yLBbdOiZ6rj81
vg15bIfUTTZlloPLMy050h4t86bihd1KvhiwLuAF46+pA/esmNUIsFhCVz0VJxtb
CcgM2Q1BBESThP/H+rsrUaKLESku/aXsNIA3Laz9dQAFtVbcf3+6KLzQBG6YgZy5
CCPWFv75nAb/qnIGdCLLlKtOOikbXlSRPHNXfvPJ6oR3EgvrvuRHGfVtr/i8ga9l
SS5o6WhYrE504UWs2YG5MecotpljCU80Utit3CcT0eLLaqkBgQvZQpFEttYI26Wl
DiWfhuF9UtzjFLpeQnfIgHWNI5MNhM6xOIvlqryB/+/+O2h1If4HNZcWUrt4yHFi
YmiSrlsMfL6HSCaz7HMCIpdxOYtmF35V9X1JU22t898X20Aw2tNuVz6NUWpfYzeo
r9PZ7e1XdOeppkBnx3TFpVv5tUoYYn52ZXCF2Kha6lHg51tF3Qy6MqHuCk/NPMTF
kdC4h5j8AM/yBs1SnzxEAwEENUUkd9wdyzAI1D/G111t5lEp0td11k0OmdNZ1dEZ
N3QovrmLscwNHYKtg6dTM9qfrTbiPWvKy7TbFHsKlF6aBiilMhlTcD3LC64x77RI
l97giuv9FbartauGLyQT5Zn2p70HD3zS5vr3uKkxWfac0jpYXi/A1WJ0eTdujrlj
YyJp2xyTeSOGdsuKtGm8G0Cmx/oNXAq392XRfyAY8i0=
`protect END_PROTECTED
