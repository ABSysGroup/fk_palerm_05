`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yt2vjgoaT9U+uHB94Focq7CDOrDATYZiHwr978esDVr4M6J5l8VisO9VneyBjEX1
yh2QkJ0G02kp0P8jQfhUqMR2TBjan0ySWij6lp9h/vahHAgdfbspWovFNwiF+8WD
p2AnHwq1MBkqB5J6nF4nY0SLOAbqjMaEMJfbyxkD++uDmNZYHff2WVZT0dRDF/mx
xKzhi8MTlea00yc638RFGs1prDyBDydNEZnBKB370RFxVBSRQG6PVQt+5yiPeGux
qBM5AY1NroPOd75sOHYN0GYXW8HAL9VFYWYCRD+WOgQmRFj6rXkRYjFbdjqxCjNQ
L42EYsQWA1WXw6mvnJOKwWslZBNe9I+tx4Y7Rg7BuXkHWJBh0Eqms0SkLcxYKl3G
9LFy1iBQl8OOK51MEVdA+H7ZBnYdsiLyEuktH1keGdJSZTj/z0MvYy2l14Nw/UEo
`protect END_PROTECTED
