`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M0HbZHny7QxrOsK0vu0IzqiydBzoSIeA0eBCczPuToDIh2ahQZBhwfDG9/D25Rij
2CgzLZW0JUZGBk5H6pKqsXD3lmz9aLW7ECiYbtyguZDbfCYLO22mLoVJg2A6Stca
rJ9ygrj7rdRlDgZGvJs90AzIayNL6Ee8bfI2chlK4Nyz7Sm/8F3SDQUEfs7g/y7y
XyRSGt0qNMXhsMGtUjpLrrGCCDsrIgVeEmGZVALWTEkiTtGv8CWqPi2XYxhVqdh5
`protect END_PROTECTED
