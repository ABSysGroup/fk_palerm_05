`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vk1WqmNJA2A11t5p7iSyjQk1lKi4TIV90JTEVA3hXqrwxfnjtfjnJ8OdgtD9cPGH
K84RryDIrqOa/HOm5lxb+PmF8XsJ6EEno+gKxd4SCsr+UDtlq+L2kai3JTaAMEUo
NJoTbc3f/dm/MCHvDTpslVqapXK/P7XkD79Hxg/1hwDEsLE+MQdQvIHxoGZF2iuz
B1oldPjKSSaqz4aiAHqUHjOuaiNA11wpSML7nhWvtmkQ/leMUU/tnccGYSReyWXL
7be4V0m1thTdy11ZDXv4pYQmjFwQwQt+MyQAPPnTYLITcrV5MMWIr9YqjpAdp5md
y6NFGQIFmrK3Qgl5lNrCG6ZUdrAgog5MDbxn0/OIIYRS/+Emt4W4XQABSEVVup3p
Py/Dk1fMy3JqKYrGwpOxUs1FLX1636Ob/N5fp2kI4Iba68iki0zQUOkyJ34R4zp3
I4LCgoTPtw1QkVVgm5fmUSEXD15YeTjVlksuXB7eZkg=
`protect END_PROTECTED
