`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bULPauX8XUnIt5EWM6HyLjg4E+/vm9FawMFoH5RvWw8kKyOQrGiWp5ODNU2kAkPD
Z8bKjmmLwjL3lyl3nGCZv15bqb6tdLpVW1ZrFc4txbtmewymWNli+iSyBZ4qLNt9
ZgdCxVjFTHO4lWKuKEGTIASfmLL6h1wJatZPk8TApZIlJmn3aAV5C/LqYxc2YPIx
E0jV8sRQTQAp/SdOwAhDZJlVzwP07cIdag4DLvBpXltET/quzmBXVrpq3gbHwPSM
eYYAsnPet3HHeOUYeWgjoEpstJHIyjAHtYEVCQ8IrGD+RrFJLgyImx9Q41ew4VVK
ql8CApm46BZbAEmWQWBKZCd3iZ4pm7qfcIQU/MHoE9heqinuZULmIwzkNCnil58V
HJ4di+dGyGugrttUGP5Sqn96krwjFYkcU2s2R3KyO44ErzkgB7Je7wDjSQV6EbkT
55GwL2fXFgKZjL2qijYF8MdkGOAruyl/a3GiD0VGpbzTWm6nrP2QMtedBqXctQdZ
qzIS0OeNAXMosUGh9Esg/uMqRKjXRRThYNBnI+I3NHoYqsLVNkhYelD/wTGhVu4R
F56cXQxxto8MeOOVEvPVv6pCpNh+QZNTqYcl5EuPMkvQGPImUPeipP1xPU4xRrY6
MdWF+VyTq3Y1bHP9Cvya+7DhZCFSm4Y4uohTWEeskuY0q52dvQiFiIlG6xSktY8m
kl9xTrhjEjmdFMo4UGgviiRsu777HjGdYr5CdwnVxF1r+aCfh1/F0iN4e4+NImU7
4/XbH/VB3i9/AUl/OKdLfD4oo94l9TdYGdQda5B0RnmY1D/EQcl+c3JruJR3C6e6
GwnNr9jtqAv0BeI7L8AIdqrfLAwiNVKMxF/9Tz9N9nsK/Y0MWzFlA7q19aV1jEft
xkFL4q9WcGK3RsXnK6qlmt4ZH+l8LJMN02hNQRnutssb57oZdwbhlstZ9PJRUqwB
`protect END_PROTECTED
