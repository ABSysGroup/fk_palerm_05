`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
84atFyMiI7mQ6m3D74AtLk+3iELH9a23u2aJFngPPA3ApD2OBz1guMlytmFK+Xyc
5VSqNtuDnX7FOxDAurxCXA681WKyOflTP2ArBmJNH9N95COgNT2AqaomcLA0cnWl
TqEuL8dHsanaqR5kgabyKY+Jx3YBSVPevRmGHrc+KDAn2ksLC56AL56JxfHF5yKJ
kUhBvvfT2gcNCFtYcx5qPUjKgI7F4AvPhatMButxJQJ7gmTUy4zX8xIDkTL9xR/O
g6gyit6eDR69VpS+J2WdEK7Xk+BchvmCCM4/FFytpFLMNYbvX6or66sqkb7fhJJj
`protect END_PROTECTED
