`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Khr44918C50EYIDFXytv/ivlGGZihdvNNlfs1HGHXR8CxScZrjarQctE6G+Ep33c
A44LjXl0lmXTaZrEn0tQEBYwUZ415QgidqVsg6/ptVje8TuPrIXmTgP/DX2I89jI
INfKk/FeLZwiQMJigqOxHvSNDc9ycNvUxJEzz0m9CJRqLcK4h6xy94DXOzd5VsDL
wW1zbyDYAuImVkb3MK3yfSR7Q4wriOrSMOdNPV4Q55Gd62ETcSPEyD2yGbUxhwMX
PHLd7VFGcq6/f8DJVPAsjZ3ZcSg3WyGwjzydyNnU9+fywp+zTJNdE31ZIn1v2S+X
p+UUtk8htKAVWobN8O4VrEDzanQIbkZXFr/Guib5cb/g2/VuN/2/nuhg2WNRHORn
vJGvSKhLDLWJkLcxMHAphB7V2eyT13/N1cp6+7SCs+67l539XLj5ag92F8L4KKZM
WEZwD6324xF/5BeaPrKHFASXR9N/WYod8a+OPpTCZhC6AK/6dmuSkSdpeg5cv3ur
`protect END_PROTECTED
