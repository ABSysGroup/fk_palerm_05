`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+g5TZTGeBMb00bCu4gEpom7bT+OdAO5YHt+LJxo/6U3NFPLDdJM5L/UF2RKg0L7I
nHJE2kub7iliIJyp/jnjX5mgmMwTadAdaAnHVvRpyF2xL1OVZ4zvygrb5gKnwXJX
TRsJo30cABOR8UwJBWWDmd8n4krtZMNqDAAsB2QWMxdzdNvnu/5MFlABFK0h/kYo
/EOqhzPkIgjAhKueAupy+/Ah8VyOwReF2IDSBJFrzYzT+SGUrqXUWVQieRrnZkd9
2pzBfviu2Q6Eep5oFo8Dq4TcVKCzEQojjmlSCenTBc76cd5f3rERO2HAm3qA20JR
M5crX4lDE0v1x0viHespUBjd9PgpWzzw1ppAXXpf1mHTX1X2GPyLlObv2Uukt/N5
6tUfrAI7DKwD88fOq2TBmH3AtotI2KexnhhIYH0VvRGH6LyLuEdHmsCVFdTkcT5m
X86MYq5BAQuhunM0zvpHPchfRoW1j1bt20N4nAWBf/WWQ1rQdxBjG8PZariDovZe
WzCDIJPcvgPJuvGX2OAJhNrmNCkg/V1pWgTEFpJOf/fbthE8m9w/BHobkD3OgxiM
hWsAGxyul/kuMUyCpkgcdseI84lktSWZIy7voOnM5mwsBCL0JqEqtuC4eBHHhZTN
rT++V/pMzF+H57haz2DSersNR3mrWtxdJmSAb4iiAFtOSDyRwuMRjXGdHsjXiMwq
Ih9nZJAak9YhfB7kS4jVhyActU4nGpkEZ+8un6rAjppJ7UV28KT6AmE50VO1wCHb
WBgGxABTJh7cwf4MjGNJs3iz17+9C9r4bqhpHblNuZAXu4UJSuY1dx80crRIUvXb
u5Eebw7wEqTNRFJJOiJBIKQNIf2wNoi3RbV2NjhDqtzJp9zXAY2YgYLqZdjagaIn
tpLCtR9U6tcj6haJ1QaFyoXP+7OXZ6S0K1QxraME8WzR3jbFvoQZRyTTW7DnqH4Q
508KU8NdV/Yyl8vavBIkDZ1eIcg3V/V2gscV+PKyJJAiBGhCTlOzDxqBHPz7Uzw+
NCNbi3wdEwdIpTZGcJ8q7mCxZtZ0Ccbn8UgoEI+xxn6w0G4Asm7UcxTidkKzUkbY
1Zquv6hmU5WLDLjbPzuz53o9wWRQMpxdxMetV1fe6RW3psXxRA3Y9U/M9Y+tETf4
rb+wHoOOH5UbvgcbN+uY1MRAzUYoBxWQe04coJh0zbZU/oTZgDLwj/0vBal5+bt7
ABM4wbk0lxdtAQcQaEyQWymQeSXgCZ53gzQ0RROGrB9UEwFqfDvekMJyZxUs114y
iD/grmnxKok5laaAV9lwBCugsPV0GK9//oYyjLOVHi0KC0hDZdGXWwbFVXK5YNQ5
wRiX6Q4uSpHpQHGAdT/bcuBdZCb4ZspfuyrA40TTo8NMJEqpqLBVdClNTYXdvVHy
WZs+N6GKXa79yKjzD9qNVM28Psf/3x5djs4sTALhDwfaB2dbX6LT88BrOruVXJLJ
pLSgvF5gWZqw0bpmyfRBwnuAAry/FAxet6ifX04kGygz0tGDV4omlPHk7TI9KG4h
zYExicikuutKP8tkOZx9jA==
`protect END_PROTECTED
