`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DXmoL6WQ0yBz0Q9twuZ1hetelkqnybEbLQDBTQEOc8/al5d6/CtvhaG2n47qFh6z
XU4YlOu0OnwmugbHM/Bd83GpNyf1v5AoAt9oEgvCy/zSaB26R1gaS3LoRHu6/Wrn
o//ZylR2ZQDcuF+aEACOXzVr7TOJTzbjvTNM/vfzPEZOhR0wETJ4ak/Te5ZuAFi4
b5tqkWyi75DFYuRrxZNLjUUCaBEckEXtQ/H5Ws6MUe68QFYmrusRXtzm1Vo2Crnv
4vOEl6kQ9Vri+oIJHfgqc6gPlL3hZ48mQBDGbDWHbmkdfic7rIDI0Rgg6Wcti+fa
Y9TEEX0y3YRlvrnV6Gph6Q==
`protect END_PROTECTED
