`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KlDm8cStpWzz7q5eXwlzIAJigIGb5t+C9gaZPLwXqHA0xPUoykWzKKVK/Sw0AxG5
+/RdA8BDLf2DGiahxmjg51ddnFUYJ0HI8+xaw6A12+vEb7ZT2T574tOzpFc6e3hO
t3WG9JrvQku2NUdmLSQHsIs5wpxEqVE4ZFahWX2/j06pZ27mAY9pvgSFzM66THoC
tzpyCm5FRI6QAo9szaFF6O7rqGYas1/3vRBEo0MjeVmsrUsPU/9R/gR9uPqvHBlZ
IfFEOQO0cL3U40kr6ClrfrmLpZUjM8lg1Mv2yKm6hGr/0us3osQbJABCA1plWLEo
kuxR2eXufXLrDMmqqdHOzyhCl7MIy87BnJGd6sD0Lp8DuAkS/Hg0LmhW9QbRPEGw
519csHx9QMSw0FUKsW0ODELaD97Ew+55cCJSsuYNufZWGNDJOKOSQO0/6MHnW6O0
raz/tKjzxSvcGqC6eCNpvNLlNNaXGhTNur/mWmVX1Z+tm/MLfqmvRlMzb/gHA0Ym
fPaB9vG3IJwiW44x2xkGDMOQ9kk0j0G+LUXgacskrNhQIPKx5bZPs/1x/KPL+t+N
OSTgp++0pZknxvhL9QUPyUMYmQJ065NiGuBkCR02x/55guJJVwNw3qSD3EFp4YKQ
956dcPYEF3BlgCoQ8CKU4tOuquAjiPVn+aDXBVGfkqHbARRa5JNc6ucgABeSlf7t
sBU82lcRkpn1iYE/U701J1CWeictrMoPTQNZsdGTIhljJzTDZ/mGU3fQFY+9nZfq
WfiOtBzgWFhjrUY8FzBWLe53PTM5PJuBRAyDCGEL5dgt5SepGlRsF0ObI2RN4Afy
yR/ZtAYHK7tIe2amdeFzCzbx6ZjeKJkUcPxt5aPzr7ndStClqN1hNUFZZqsuwMS5
1VL1M1XQdQw82ATvql3oibXdvjatTu3xvbRXhfN0bn038G9JHQxC7cvDoYHkaX/k
Fmp/Uuk7YFd8TkBfuIkcAzYvFUOvQUZJA8qv8QHa7mnxD9vbpu7+CmkMnJG4mABw
gHcmAnJ4e6J6tHoTPvWJFSxvVf7v0saCtwSYx15s/k6Tn/Lm/SPiTWspb8dBkVH+
sGtQPNQJYbWYPAhl9Qy0G6GOE2Ou8AjBogaQOfIMxucI+2X8ze3DzeprfAgeKjtS
KZfHQN4XKKVc5wLKvheP5B8r2trsGpNhsmtgMlsZ+y7q0P3veHK1w8RdVXxVnG7y
51+yndG92aLiCaX9pRi8OPVu1gvdDDdfacDEinq22pCjs+GMxlDw2QTiYwr8XTSY
Nt3xUeiZoRa6NgVj/N0Akg0GbJWHNcvhQj4WZpLLePNenpmAS7vL2PXZSbhukZ6U
42g2H0+SS5bEDSbEpr2BEgxYbjrp0FoD/p+dGtsdHMHsEDbAwx3JxzJLwsOySO4L
rUX2JNCHzsYF1COkYo1l3o2DMw8p0Lmqw71t4nWXTA3PaebQrwUjX1hO1FXN0Z3Z
ADQjP3jzWbA9q+iij7MCCss6kmytUGnqjp4mYJhuVYJmT7Vb/gqrjoRLCnh3LsXM
mD9ahI+9FkX4ZY+3FFk1t9z6KrF54cCXBjKrN4E4x09oLU7TyWT+IEU9vc9gnAEr
UrODRJhyGuXyob3Stj7SAJmLLs6AJLd7krp9RYLC1Qz8XPwq+yEKw67+gIl0EPuf
CTbFq8Wjk9UbFD9RaUxeitXNectVk6fuUVUsKF3gOtGUnVxz3MPrRirak0CQ5lPr
wYU7HIIN91zng6UCc2HlWoX4P9UvrwZWbP44OpjZzRZewEPiq9CyghhWciXBpBYW
JCWI0q0euuOcxyDjJ0k8zm30IUItlGrokYJ6BTKZmEwPggrHAmRegS0v017ZYbgy
vv5mjMsf/rUwiiN66GovoIftYjIYJdd2cuIf9aEhc7UFr1dKXtXD812q1Tvq9Xq1
4oV8WPC+DIB/zVsyizSzvgPYy7mIciEcUEl5luFRSaACd1ov0uLWgPQrFKoBz4an
NBfO/exxL5bBdsFL5eN3MmID+vYUl/b9LL51CH0fqbDa6lrB2Xj96AR0aRywhdOZ
UPlhbx8/E6wEO0F9cIqmOiF9VRgvmJcjSjF6fdgr267seOOyEIYlE00q4mGYf66e
TRuKOpgQDIbEku9QBVIv4NFQ47A0VR0nxnWeov7vhI+JP3BsRV9dGyApg3Bdo64J
03n15uIjYdl1m/INsMDJYFoawLYRVSnLpAK2PfDHV5OK0DGjfDz0bp+/d7woR6C5
yP5EPV1wXk31pMzAn7Tx0NnEs6iEMbTEuvvqcsA6i6i65lcKzp1yyzx1JqxTYbOv
lhP0lef+lEhcBoT9Nu4aYd/CE3rsDI6sYooHfA6V5B49IR8xh39xmY06kAGhZskp
Fc5lZbrWY5FFpkXsD06J8n0X2e3jZUsg+9IFTJr3kDrx94XnmrIFqFxZgl86KuKS
+xW/eamg32rD3MTtI7Ak3B0EobNHKnQm06wi4bfytTB67AgtTRKnx+rY1yCpJuqJ
XXbHv4gVydPsfvXOUZC9s7bHBillyuOXrfAZjJJgR0oovwGtMS3feUO7z973LPUk
snCGPxKIZY7ST5EkTj1Z07XGIGmYM1GUFiCmNPCAz12+STJXZSFz+YDPd8JeQX6f
ecCFSdHXfnG9CPnT0T17BK+PAsoi5ZrY2hL99SfAdJSxYFxsqEFNI+rG0UPFo6ol
0zEB35YMaaildAgHf6YIdzCsmOZphwY4VAc6R+6X5r1YnpMqcRnYQd3k9onIcYp7
5m79dRl00y8QTrzNqAX1OMQEHBvY6kVh0Jx8S/1izyccc57F3UDN9MrsDIHxXDix
fQXrRuGuMO/ilrt9+JX7QWP2Z/wmdAk0Zg/TTE6bcz+a76QM0eyeWYotLzrX4oPr
LnbTNkOlXnDA5lNDGyHtkEbzThVnM4G/fpsC9R1+CP8PX5G7c/rY+Zt31W0fYeaF
+ipjqk3LFKlFjcPgalRgL6bS8AwzTdwkzAWSwa4bnTt80Qq55oB3NEK5tqbdZ/vi
obszQFdhd1Fkl4lVu8hXKaqxKGOyO4Hcan9l+FzEfG8ZJ1ForgQYxr4b7y35+mNl
jp6XBBAV4Spkez4YPP2m0ZB19cRADqNIsU6T1kJv9bWw9BdUltNRffA038tUCqxy
aoNnurQYa04hAgR/cz4xdcJ302fCmTqBHvLUm6znG1W40hkRnUkcXblsq/SUKDa0
c6XX5wU5WlhrkLXlxoiLPZkTR6Jn0YaxJrk3j3D5AHIEU4+LUeXhTb6cX4DnnIz1
WljOnuvfZppZdPsneiA0gtFR4GG9P0Z/LHztqDV07B70RBwgBaDJ+jPqHTRzvoOP
v1kYMEaGZYnZm/9g1ny0+uSo+NgIi+3XzYBpKhpsxSyVQeUlPTyroMG3pDauP+fh
jJYhEgj/t6tuuXZDvMDIuXnm6lVjlCauQHjXWEgnOXyILhSVmI1Cv/3sLc1KVZDK
99bAkY3nfEQdnfXMszwVCt+AkrYHKqu+W6OdP2Yd4RI+SLzp9LWrdPmQVmavOr3q
Fp9w/UWrX9J4mWUZtOXKpT14fHFM2IGX6qesF6dd4vuZQwUfzG383Uf60QKgiW4N
5MPakcNfLWnX1E7V2tsx3mRX11ScorAhvqCCzQUBDsTQxabCYQd4BpDaMt/RdbdV
c1DxNHiWPcGLgV/MANdp56Snmo/nuX05o6JczyUTUWhPDCfR7csJF1IfBDcrTluf
FDqjuyksWayPJ+VSt72Pp2G6QuypkGh/uZ51j1hlGs8K+4rEn/DD6MU2dPVENeib
MhPAQHDNm8xNWhjWHuoCRV22hECs+s942uuTnDXpc1adWLfNKcFA120E84lbX1jH
iS3Npr4W9yVBo2WIBFZEhzKitQj3X/bIETFsQGaOSe+erqI3WaZtWRwINHaPwV0d
PmzHhcJv/WaK7HckfckEcIKo3kJ6+i+qpGU4IISeLysNygnuAwwmUg6y+sJLQdgV
TdWoHWB5UVBg7VLFWQ7fo4wqYIjonNTkKv/yLBuyCYeWkwm/p/PQFVeEuwuvoUPY
LrRCkGqZtjyWqws/sn2c3lNmo7PZWrm2bf8IhTiNphF8Izchckfs5AH+6pYYezYV
ZS+itsVhFyckyWmsOZSMczJLsdJd9iMb+Wtbs1O7kO+ZY2gALo2rEBgFdlJtatqb
sdUEa3p6581pzYYLpBl0xEEso/zbPwL3jZeoIdqik+UsaK+IU0KgJ5jerOWTZLhZ
sSBysTYMu1KD/f/8T1L3SImzF7i5tcUZ7EuOt5zJJc7j0pIrzGQgSmfnu9G+gqoK
dw2bQCQwr5XW/ZbpLHnCzz7KBUdNQhRV90GUfw1z4yE7LcRgMx9seSmu27S249BG
quSF6KmorT823W6eGeD5ZGVhrljXJ/rfkjE1LQGOiAqUgoh1YKRog/StkYBt9NZk
Uti7N11QaDiUcL7JvtM5Hxfg7v/TuMPFPvp4kf69/D6Olw1fzvp0aPm2OVammsCS
Ry5YzyrpfCeuzqn4SndbqV67I2ynlWz78HYJIFSuugOYavJZ1oCsSptyLcQN5VtL
0YrrgETKX+lRTZvHxDPmpiyRrZdBCwi8K5glApxDDOIgwqCKBCdSZY3yPbwuCVsN
+2DMoc6Iu3yeu+oBiZqrav4PXTT7WAknL5rRKDwEB7LCFxnyzryqlQMCpqoym7vr
Yp5+gWW5TGcI9xdLApExEekOUyX2JZoZE9zxDvCutjVTNk4zYPb3JpkA5YLu0nJN
l42jWQBGSGLw4q54vSCUq6gRNWbR+jnVokX8Al5V4iccicluHwHoGamMgI9mVnIp
nWw2mLudXZRhW9rgiEEh5O6IcLYiQ10B5mUln2WRrOFBr4gafK+/pE/8kQHIcvp0
jzwo5Tax90oXYeV6QOnuhhM8KNaDKEfWHA45ZFp3qDcpvFyvxPmHWgU3vdyLi4h3
rAwIqKtQDDc8d1FYGrOzd+hdKTd3nnql1FTiO/qPdgh/3F79ieFUjOM5cpL3UWFb
hI7MfL7Or+YmokmKdO/99BuAmrXamYCJHkem2K4F/xztVE7+j5+52h2S8FDYQxcl
M+4h4db1YlkWMEmo7+72shkGnbPTWfeIRl4HO4Yjd6dd/S20Zg7BpdGu5WguiJ8X
Iwp+Od7GyH0XgWK34y9N7FSvcOJpXAgGf5WnUjuppsqxkFHjU/dX8sbi9W/J6HXi
ojKJBVbkWcu5ERWi314EePeCARWMHYmb3Boyspe6esNBW71y7BvWiclbQJ4J6Exi
aRzG85i5W6nmM7WFfsbVNz3jNj1249odECdc4p12IOnt/KDbf+OT/+o4fTY3nQCJ
n9dGmGZCb82A8RV10Q30SI1eQDjPpC66FsFT+YneFVQT79b0S70j/BWwf56TdJxR
8McviJxsiGHJjMOhrbI1x2V2jJM6TuWsTosyoPxLyi/Y9wCxb+ezvPP19g2rNQh/
nB8eOYQn+39CTiR/c/V3Tck+yU1tTptCKqqbJppvrBwTjCezs+a4MHCc4rEmTseN
i78CfUDHsGsEGR4x8WOtZwqpy23GpwqyWwVeUdgmrQwMVR2VbDatnAZtxLpwktjK
HromVnO0yORCssdqHzJjTWNIzyrhdhbgVqSJMLhhSBBmLJWfV488kcZKZLXmIWTG
857BXjANkfWWdsEMQT/WEHHOzD37T0iwvpQaVK/5Di02ltJJkEgUfTfKgvLlVF2c
4U7ORV2fVuNYuJp4ID2/slT4K8s5jFVs/HZZK3bh1GZPbkEc++UeAkeMthZjDkVl
bEeh01atjwq9UCG8ZoHqF2atYuZDm2KJR3yOIBhJYfi+zZu8ijMZ03cbAu1NG8NU
cudV9Uc3Avr3d9RVnlhPrznsDIhQ0DKydAYMe3X0Q5fadImRLrEh4EwcHpmjCLxi
x8uE+h36BgkPl0PRQ+F+X4XEKVUEWUYwan9suKCdTsKAH026izD0PoZIKm+2EL1H
3sU9CGS7t4dqKEdBMr0gTOjrcvKLLe22hQ/HtL3XkAruquJLTqJwjq+/NqIIw3Qk
LXgvUrT4lMvjjVV7lLSQiaN0tveUyVqB7mtYkRxQMkupNdg4aKOCh/2IsMu2KF/r
WCQqv4qmNyHqIY47XiPqzj1Kq1Nbys86fVYzHJ10gWhLSfqv4qT09EFfjbjbN2tD
k+f7ukmRSGnyho40t/ogRrncIZ8BrM+xIMNK1VFTEDyGAe0XUz5G9WYiCpPMlDcH
1yVu9dHX34L8AINOIh15CcLYxwk+fGdXw/FMdMJ7W3U4inHdW8vK4AnvcHcnsn79
F8IwNMQQCC4jaoUmxn1+choFeGaW0a9Mb3jd0nXPnUtxWpTXOfm5T7zud2ODAosY
PAosGRkMwAYpSokzfFuvXYEkpIyF2atmS5TNBL909FvgIuoYm5sG0m8ajC5xBtjY
S0FtOj949NxsawoO4g/lqWqoIaYXF4+Iou3SyAQipNmJLLIxzOyIg4xyyOfhCs/8
gjJZCj0yxDO7P+Mk+Af8ftjUOTXUIZnDoBMsub2Ir2W20S9WAjhMu3MKCtC/czG/
YCJ2PvcH79Lm1mU8vxXI2hQlh5437uE5p5CGy1tLwf+0HQ1uA9a2pCar0GvHtTei
i6H1m7e3Es5jhZfYyBRzL5LGtpvZMDOUTo6oMCuiwecQ3/SjIIVclg9mElgK1tuz
5dKMjm/KbOc8vkx6Gb0XjCmdi46ysMXGVW7extyIkfy0b/EEkg7mEDAqQ85NrC2p
bJiMuMwQk+SCBEXgoXOTIYhKsnNo+ZVma2CxBk//PPtT5JenrPHU0Ej1TRwf4da/
Q+JsLjYKc3+/dIXJ8p/zGwhE/v6YgJtxaZ2I2NWdk5YXbg65pexnHDC2vNDbr07B
ly7L73dgBvnEI3jBY54JOoF5z0pm2MSB76QVyrV/V4CKk6AyZkyO9B/rlcVD+ykL
6mw103OwGcGSMNozkXoqm56cPfmt6rTFqB8WiEDDt16NIzJqR3NKbF7XMbQVw9fs
q4kvhg79g315IBUsATUnYZqDod67yxXBUmS0TkAsCtsyHzBhVYjiooHW72r27/oV
IOPqALHyC4iG6iCbYHbMEgqLKjdesncKZDpvTbbbR2Fuf8JPTJTC7SX8OYwqVFti
ns7Sc7kTxt1S+aCKWSopR1hDsrRRT3+vYdgt86R0G7dD5osxYU9Q3Pnv/BTLe9s0
A5je81dqlz7MVw3FTKii08ZZgCWDZBvz/C6SoinQ0i65D5gfzCbsQFbMN6RmZNHW
7fInFV6sbI/eFPSOXsmLBPsV4AnW+CtrTXG/aarEo8g6OgGSegPIdZYbm35SL/9v
W93D8rTYvdyZcEQPd73T7dE+mWC7wjJ+6npi27MlHt7R3scKU3q1yzv86s9pZfyd
LhRNfPZShNedLYulYdrnYgSkM41wHXmtcu/PQpf60ovPT3JB5DUopeL3e0feAZ+P
Wq2G0qKWwxwiNljqEr+ocRo+ndCBxyjbXojC/3Ptyg/5IE4l5Jx5hZT6ITJOFEFS
cVOYTxvewlOKTnGIyGjnoLj67T06YPB3FVZ701bu/JsEo48E7774MikyixZtA8Qy
dASqhqrIdPGLTuM/D/5ZUcM1w1i046MwKHkMuc2D2hiorxzQuzpy3ole3CKu6zAj
osYnortFauu2MInK/LCGcg6VP3Zbkyq7MfLKz5JPtgq4QrPKmhAZ9z2bnP3VPF1W
luvR7pneg/Sh5VYwzG/fBBK5YrU6kMvzoc2Yk0fGlhAe1j7cPH8UZXuWW/WXj4n4
HH8w7B+UOqUH3TXS44Vbbwyfzg9GoUb5fAhd8CcBPlMutdQbxWNgymC7ZXhdokyZ
5cDhFNdtNmovSDA/cLXQ6meRJFqRXzOZ38DTTyeecXe/Uk4jyBKKXn6ZeDZ9QJyt
Uhvlf2OoFShYExhNK9wkI0FJLOXQMb5SeD3aYJRX/xsBnE50G37bdhQOhbUr0G1n
NUGZsmQrxSF6j5dWFqIQS2+TTQVvBlNSNTAn/LfbuCioirSLcKoyEwMsxfPcwnZp
43pAX77SVc458mwOR0008qrSLENVL44LKCzTTYMRqluMY47R15y2cCcsbviXYOYu
LPXGOO+B+vosVSmFS2i9kv83KXyXGMym09BnKaSP/oIuJRmm7n4LuGlqcyrRjMak
6I0b6Q6eYhEugewS50BnSAG2WtBRo4KVVBZEZhH10e5sxSWA4cGrqU/sxTjdH9R7
2DHvJZcuNwQsWcJ2YxSWpndVkINLZ9aXoJ3FrtMMBthObK7lFYzhD0cSqsdq+6uX
2U4ZZiq+Cqm5lS+bTuOG5RnlAWa6vTvzySY5CGsJ8GTqeQzdzHXnCkI/hQFG6k8g
UfaOl9InyJAheivBwfMK8LRrz62ah289P4PNcNa481zT3lVhGfGhnyMv0V+6ZCcu
oC3GG/Wa6ODbtZTgtQMpxoX7+xf00vijtx3WwzPCcwiuPpQlq1WMRLcouB55X0JD
HXZAuI2EUVMpHxVlZtDw8sx5IqLc0JYm8a4CRtvTyppmshYd06htw4MMe5rXewm8
LyoNJkOHGt/c1ZAr1m4UtCT60MxIJDE2kYmtHuOJbQJX3vezRmVDjzMBrsfLrwiZ
LZCUNFiukkDukp5siEMLVXOV8Rqx/lKvGLknT+nzYu/SFv2sXDEjYxLJmXy+NjnV
1Vw7tYVwXm7QZUPX1FtAqqCTGwxjjToMMVAzga4IKz0fpfxL3q9LHTQ8Xr3UsyWh
aDlnqN92fERxtja6KEZ0xQKG0/YHoavuCCmv9l2hFzadclXV0t5yQSYjf6NaTMcz
apsnoupAvnZU5tEaucrneRqwubEJfnVcKMg6CLKXpkGSsTmEVUuz0qOOPUhDCz5p
uAvGhKEJfBPX4+YWUktKMhY8l0ZTMP2/OPEYDyq+zQQhPHrXTzP5G4x74eI9I8GY
3vmzlja9o1qefLT2xkgjbbKipXVgrykHVJ8YLqfr4jgqIZmkrEBv/YXx648F+GLE
JnBPvH/fYcIyh0PlLp0G2DN4or1WlxQ2qcwdHxgXIGVcfL2+eFJe4GJfW3BVsuFx
DOzJvNeTx3kATyvG9EEIcPqvLzG5oilgUWQ38dRuXAvqGFJYZuYVEXFnk0PEGlmi
ahPyR2cR3nt1GsKPRbqWKk1q/PRxdWbugaftqptEBbXyJ5yDMdLdhU2ktjPSWPeu
GDEFcEJzl7Wb7dAWtDmsVqPq3wyUefKTZu3xBmCaYFcVgeVc4t70sZ1zIIJVevsW
y6xCvrnXr4bQl/PdthT7KYXciJEEQXFRzg1hPBC5JJYE/N4c+ECgc9agMukhm+uN
EjcOcOdeGy+wQEn2s5s5BJefJjH2f1SYQ6aRM/9LpOexrN31nbApWmC0NheyOXQC
GWBb4UMZi/HbwCJzkklxRmtZy2IG8RoFSC50Kn/qiaMWvrFKL6aok2aI2dHs7/Sc
Pm6ORgjqW5exaCLxKzgvy6/EAp/LdeFZMnCJ/nP22vD32p5LnNQOpjg9lD+l78lR
thCo0amab0bkENWu96CntWDoTuS+I4Y3ExVH4TuHyvsGZxokLfofENZdTqFS5gpF
cEExiC9wZJwc1BCPF54yKJt83bfmK1BLvwkXxW1QxffXr6BsyQJHl4Hb3vAXSRHX
GY/wX4QyPZ7VW40UZQai7IY9cKGRkzXq7jZ5/tr+aC1FfnudkWRr6ra0/nNCJaWX
cBrFRt+4nkS7UcS3ECWmOaPhLUo1o9qsCKk06LdAK7/wJTLCJDIe7H1In3GTj8mM
BSCetNWHIA+v/K4JJN3XlP6Cd9xnspF65f2nQAom2/IfgW4xsnFSQsT6L9ojQgS0
oLd0OlzXh0Umi6QPQVaWd+WPsLnXOvzcOhXP3os3WdeSoD05MgaJLzWZP6Kx2uT4
BfOwNJ9NgvwKXOx+oe9qwUUeNh5gKpnTqcGc51PmvXYQuiJMXG3+lOtzm4kBZc1y
eepQ1YqH4ShKgooyjlPZj1ukONuICuyEEi1HQMUAhTJ/wgz5fy0c5ADh1pJ7MjWU
wVAvld8bbF5kKcM1QPO5aPoUypUIAcgC8f0Vf10tXqtZKqQd9eFA7d1c0Zuxq6bN
NuoO3Nx5IuVuHchMnq2NCSz+M/X+l+zQ496k84ZLoqdzUZnXvbISZo0aDSjFV3PK
KKRho9f8q3Rttm0NPPixDW0BAQgzVx/IrhZAxB5UeujiqgMQcoDEpMtMMBkwf1Wq
Sao+iGOfDBLPu5DBzhRa0qGGS1EaCDdwNWTwJkFXBWfmfV3SneIxUy8Xvt5i6h2H
8X8hJwmN9fgAedn0rQQGS/8vT8h4lonJBORmBnueRhza3YxKt7ypJGxWjoa/oxda
UTF6yRzeFSTFl6LQkavis/0af34u8AC4+ujxd+x5JbwWnMLBpPogMWYhQ1DlLKF/
oaxRan2ZoXz9VUOX7IEwcxaf67r99TBHzIAET92F8kLx6UxTrNq9T65GzzSrHOxZ
j5XqH2iHekTyM7XulSPy9aW9noZwpkbvoL9aB9g4ENeYUJ0OJVWEAXv17AD8J64q
7+5sTAUleL0HSvjRQFIMZtrY2duEymdpZ1GMj0pGGuw68eGDy7HtdIat7pZFkNIr
BnyO8Wx+EVlf50NZdd88muFAjuaSR57hFiEgtYj7rVcjq2mtOv2QxlCWTIl0ZZXu
pwE3q7ew4My5m9TxwYM0qCby0in2ShYpsDzmlU97JJZ3t8Ju6dpyz9WgTWwZfdnp
ymUt2Y38JUdCFZRRVKd+Aw8Stey8kPJuPtfQfSKyHjtcJmmSvqeXU7ROLl6pJyRt
opojdurIB7RgJQeb8lv1aVZDZgE1aK60bkvj+x8JQiN0lskeqUptSwFvVKp6d5ad
JDKKcEbtUCwcFxn3XCWnlZF4HX4CowvM8h3yxLAp7o11GDPr+OwDvy7D/D+QUVQM
K5mxOERkg8HJqGpPvvOZeBdCIdA7F/o8KT1P+UfIy4FztGbWd0noER0Kta22378f
O098QsOoAbjzsyLaIxM5VFUgdQPUmP8MDahU/VK9wmEPeNU71+bEjhoC9RmVkAJd
fBZTLc7rKCCG2su9StQ7KKPhseNccLJ73dk+GWJeRfHwA+oDnrFr6XWAfw627C6v
vcnb4KF5lwjVzYd4n/DzEamCsj0EfvWAPyaJti3grr36UmGJunaYqcSBB3A1VLRm
62lvS2cLXpaiZ9OEL2BSXFqS8/t8d/UGPJKXBnnsf4N3YcwcgdxdL7Cdg+I/5BFK
pc2YfShKEk8S5RYOucYokE+kgsXegjvDZTdgxpEfHpc9DiojTDoEdUb78XNkO4Zh
3n6+dibNBQA2ncX34FhTu6NgM2hdyH58iRphzLFijNf5q/cPS6Di3FZttHtVP2x0
1F9Zxpda2QXlMu2LaRZqH1FMrIqUAIJsb4iaYx+k2ccw0uah5Vt5LX5nouEXR6TZ
Urx3FSdiGzNrWs63kCxfyN+wy7p+1mvZB72kE0Sb+CtKdaRyJEM+OLqYLWb8voYE
YCaRM69EputYB3Il2Jz+NZUrLS+bjNlw2odVWOnsM2h/E2ebbSDPV1SAINJ4c6HE
U+FipmTnGNEtA1NH92n8+wt1EVV0nZGKLmCEmToPonP29xfX6t2uVphqhfDM0Ail
UzciK1COkst/pBeQmzpG/6cbktD4wjWUn2wWhl8PwZ8h+YVLLX4PBZiMT45opNcc
fzt7ouhyJPRZq4Gb5blYjDv11oJrb3Zbg6lVuFca3tJq5c8sF6CfzAefeHD5eXuR
YXA4So0RIEnHdqC9bc7svT3kluAmyGxmsdS7sJXkVi8kqRw7sPACzoM5B/oOSTZZ
G2lcv6VQWz/Fu1ZkxlhJzssyyFKknIW8M5Bo29ZMzazGIqINi0g7B1KOF/xKOQcH
efzDjIsy4OlpjVl7pPG/5iy1BX/XGcK68YoVyvKAWhMlmZDq3UMcXnDnDVb+opKS
bmF4yah5b1oaNJDc2GVGh/X8bEMSUtUjFu61d5gehFsV3rIcLmFzWrXE8Wpzw5TT
M5vC++PPmvULsDnpZxRy99dYQpS6jrBOGV/AJU4U9peSGWyj8SbGDi9biqRZot5d
Kq+7lmQq67LOzy+jLiA6hlQt+e1L5otEd/CFG4Hsx4f0BOp3zq49fOjJAsjHRS6w
PqpSq0RRjsc/dSuTUlAVLtl9b5EHI4NrsY0hrUciUgYaNLOiBwNMM06EO2lUcV9J
Y6PFqElKtYn9YKrcrGEwBPZsxBpT6UWSqqpTYCfN0EwMTMsuEQC+Ldx9RiYbnYh6
Lhs+sY/ClrRIucz/CIM743bKUBbh99Gba+gQkL8ayzT2Sc5Z+vjPkK9ILQ0oYj8K
PEGtAzWOw1rOZyXoCIcYgvzbfH2PuU2Sohu5cVQPo5sYqUVxZXkKhzXsP9RT/A+N
qY76SO2S6Xa+gdJWuTbPkuZ+35b6i2WCmgqH0Hzbw9VE3M12n6M8c/wSHZi66kxf
L6S889FOeh0Kf35bmglPD+N7V/jdsrqcFMwWhCRImNBzwAsDQ03IJjzCp3jg/id5
DU8s428Pi09Yv+JWVMLCSDtcf+9uUobHSqSzXKxOuMvKeSXVgXwxuS2fwJ43yDLi
oQBvisd/cjjXJX1w/kJXjj1bssf8rbrONhry+frGsw90b1hcKZPuzvn+tuja501U
MBxrJlT5YY5GWwUpKTdKyNAS7eoOl8mpO7PI3vX1MbsCEoOCTLVgoAl3KIr/YBEZ
trKzwaCoXb/IQxsahPgPyiRZ1F8BXg9U9a9VrHskGPpIyQGRcqAWK4n1yTikgcfy
nk5lPYTlE26MrqqkmVAu6kybGs7wD7fYL8EItL94egJrYrL5hUoZdo4EkPszyCMg
fgJhNzexfm5NtUW0jXK1aByQ/s4PH/1dL53pnAKnvSYHcN5CyXP+/JBh5YFd1DX8
aFnFcilho4AUHs8YvBTBNliBHOIIhC1tCNRq1MKg5jlzo56kWsnXUGhSdRjTARCu
BOONpi+XegSaQr5WvGqXahEqkyH+QEb5x5VXq1fG9ItctTv1gozqnYOfvQoGZt8K
i73fSS4+CQGLFX22aJzYcAvnnZiD34fNfw+zofD7SlTtn77GP7YhreocsGNYSErT
J6JQTB5ES+u0yWcyEckkWrmgIe38ydTZ3VwpNFkEWPFlRlqboy+n/ynXIJBWUTZg
H5ilK+DXBqSuLXRUKB8hKdIWpdUjrPlnqA7pnHMu9+5mGkaoLAqJII11ZvMkcAMI
mvOd55lJqHOjv1V6F3yYEIk5ulDkolKeDAuM7NG7KDAqdBNHbi02KuHMpzUK7G9v
BBbnyrfFOcTqOFDBcg0ZHecr7VzEgtdi2qmNNPe9/2EBNeYnWdkLhaOJi41Z9gGD
e2akMGrrTE8xgUuHfqIQVxBGY1SRd59eARiMN86CVTDTTR4dmol9jeMfv/2Ud6Ux
1mjTjJOhfUR9BTnUCM+dk/keFxJa1eP0pvAjZoDqWoZ9WbLip3b/v6x+QI66qvKB
O3B1R8NU1uuowFqlwyq+u7ah9h/cIJD9QdSLU55MNLhX2uHMgkdiGIb3tVKZRcEp
bZJlekb5Xlg/p4cEyKkhqNTkZK8MX4KG8XmEIY16L7Dhtzoy9la8u8FWSsnGwWxb
qGs9RJIQGMM0O2dbn7wJGrt+Bw4W1kB+UTcdstCrXy6+6NeU+RflBgcLuFC7KK3V
ItYyaaYraTgfK8UNqWs5Vkp8wwS06NNCYnlPrVn6iESIT/Z5daxNG2MJpzYoGdvN
kyiutc94uB5t2N38wf+O/GTrDvhVW63KNkkSK04Ru2t0c+T7IMxfcffLSg6UelnK
T88Hd6QL/tpBMSlhx496rXn1QEEOdnR6QWlV9J7VBzc1/wGDksls8Uf9wD3L/mki
GC6CgiyPTjyCpPkMVGdTBH7o4DQTatDTUKSJcxOXVIOmEHEpmBG7UdjV3rlLsfjQ
TPzXinYHdC+Vk9FGG3+QnNfSq4a+xFc+x2Yea1pcPerqHptH9VQKfWsXNmM+Ogp4
c9MoouGfNyWaCH0UJpMaAC2YTpvA9KWfbdge/KWmHa6h01LgvY++2xkryshoksMn
sTVh0F4QaTmiLIEO2+Xb6BsXUwNSkDG6mwZEuIXkvGTiLDdKB8k9rQPaqCnOVA8i
ZLskXkT63h9Mvg94+pTkUO5wy/7ZoLzhiHBynS3rJTOPg/ulAflVclWG2pBxKByJ
KexlSqRoF4/4Qx+4f7KjKyE/eXhNj/nPxHN4ooZVjzqPILd+eJei70KkpB30IO7n
karSYGt7sRG7glO3Sy6ARlQS6SpY+yg70zMpsRnGn+wgimBvs9VIY1Zp6ZvYqg+g
p2sU+/6Zh01BHWI0w7IkOj1PZKaeZIPpCWVs5ixaK/3yAR94ihXeICEkAFVL58KI
Ldr2mYOiXzmvs7EZVdOaXCZX/PXUnv/+c7zRS+dSOk/gmxWyLn/AoJlvWZcaeWIV
qXNSruY4xugH8NBW33ZjJebtI7LYyziUPwM+0Hp3t/yE4A5q/9QC9mi40JCsytof
9/WHb7elmlaJLKc+v5qCGqLzi6kVOgTiQf/cCs/v7qspNxgZsZzugYF1fIXCSDAm
UTXMZ49fXg4A7esWVf+wwArKwgDD9SKIdXZ58MZ6fqIMgzL4BiCDLywUMO36p39J
M9T2wRPpHLP7f5wtUhLQnSFcIxm43zUA+lhIrbantCsKXiM1ZeGo+f5EGoYxN55k
aTJu1TIxQ8NXQGtCkrqkXoHDIr1mqygXN82vtUCxZk4LoBzyMgunSAe5FmHVLbb8
IskW01PSEsEchrQ+d/Qri1+/bJg1aJoxl3w3Tf0lzlKNR+YtvOGpTdw0QxVTsdFX
8fK4nYPvWs3G6/F1XUiWDkybDdTXr+m9PM0hAqETFh/O077Gx0lWVfGA7JUgmvtY
L2hopHEsBrQUvbjivUuL+WRr9pH9EGh9IfHqsuLIkgnrBu0463zFSBa4MpIhZaj/
Jb/7DmdnOFhObjJew2pxfuR8x4izHUWXOZKHvGFRBxMJWbIKEkPWbJvE4dh+NILh
qzzszbs1HjOLABOZA1jtZfEN+5zzZy6rPdrDz/FUNniZY5a5jW+YVnywx0gBq6z6
+aNAhRY1ppgowcuTAbibTO+vlRsH7f7EFWrT0gc2NDnuCHFLRL3GYGNtWbSBIEn8
LzNV4vhGOdw+JTtAHqA52+CXFR8lRSjGiXUyz4sZRqCN2ACcC8a9WNLhTHaB5Dm7
I5hYlIfrzmw/BTXo0NQG1mJsuQc1pJE/lAHT5XqrFbCbkR1Im2STOExkZaxsBUrO
K/7sJl1vhnWMKO67EnMY3zOOMfBFdFbUvO59LepVwPgcTX5yxx7EsXzFt7I/SslP
XrpkSx4Xn7I4kzgfAefDkON+wV7ZRNjSGWgzRvN06/1eZVe8qJrrrJVvSR/aLFJz
XeXccVBvY+nUEc8oK5VP9JxfOaTS67afWsKgQhLJX8f2J4GV8lPPgZyF59C2yz32
b5xTc4nozfHxB99nIgbJf8nSBTrd2BD6vmT2wQBN7vC8KkfTsGPdPHZiNqzgJ4Ah
YzJD8mLnsM1sp8DsPrx6Bdaj8WZNi7p/stbFEgFpPCAtts8xfA2iaw+Acc50xEYU
MO4/V9dbZer3iShM4arH1O9ZKx3nA7D3lCDh+65ASoGTGlQQFQ69n2U4Lsmvqy6G
b8Kjf4bkjSPT+UqZqz3Ftf/DlsPgSE+xSd9ckHzmQMPlUglUM7s/IIME+AG+QnBs
J3FZsHlAVipIC3VUC1bsp5+gWdtIXEo5XFHjyE2nkfnSjuDvEN+jDl2wic+vsk3N
Y6PGV4Lya9Doxu4DpTgsWU8isUgdP80+b2pNVjHLZePT2nU1Id0YpX0XRUvVsmNQ
XwMsFQMNgVC0klLLe1XHlM3zxY7OA9BioxcoyuQimRJTnetSlSSWwYWIBevDtFk9
xvdo9uFinPnj077PqiTjpxEFg6Ts2hW3aA/HRmTMD3m6E+p3UH8kV5ifr4fbG2Vh
MGuI3s01JWYNK2Z/aA0kX2dZuf4PBSUDGVelcAgxwVwAhxAXUPK8hpdyRNDMLmI0
vwMDLSMIn54r+6PclzevZrdAayaaWH8zcBKdU8XTK07vFY2Kh1GeqzeIfM99jWGB
EvI3Pc8LExhBudIovn1f/VDZbCvi1Pz9cnYnrCMw4Pi0Jqy/k/nVMdakdu0t53xq
GwR+oCLQU45ER9Ng44f1dHzz71QM7yZyHCL6lW2BniV/FM4aGmKXPxPkUKJ339uD
P2xE1jKtc0qApnim5U68vqp7YKlj3w73EHh0rkq3+TpUkgKh4ZeRsEQMV0l7LRhu
paB8s1R44mFzAmiYIw0+ZHExMufXJIX0Vp+DB40HcYtuPAaSSWHyBL/STEmSucyv
dy2SNgwrcmv0TbP2Mjf/KiAue8zoHs9OY0RP8uDeELWUlNHRH/6vSB4hgQfTwKaE
6gbKgvN8bmRZixvKCMoZhKXQV8gNJexvzd5b91eDgDZeSdxvTmiU9dGZFbCWHTZ2
4GxyXdAr6XwU7huYSU2C626N155AxBpqrVx+RqkG92i2hrCEhod3VfEW/8vz39/4
+sS2ousJi+XpsDoy9wSHSw9CYmSPrd+v4Rnv66w65OXRfLNM1gVcJnn691haCQMf
2mKc5Ff5Zo5xVfr/7MfCugr5EDnYgNvh+mvzlljIZmNFUaV+DkXu3RNrlSKt++9m
n+8Q34crVAXQ7Dg1YoXKZFDTUJ2J5v3zS3wDjHo63dlcUSUgPGbUtYtupH22I5Ts
EllkmwhEJDwpYP7Wft/AhrBGTwvqXSahjo+Nl4VfZQ6YfPySHR3hIgBkMD2RrUOA
5TdBXJ+uMt0SGpCYhgjsGyKRK7OmMCRe67hqK9FsCjW2k7Flawq36eCZxUNU3KYs
ma5iCLDdNFYOQ8F10nRDnPW9yJvvKaMDVxCA0U3Dn8vAiODBJZJoNi0x1o96EFeC
uJbvY3u5RLlTsDcoSVNtmHGM0omzHNOoeJKQ5B4DW1MHFudXvidxwHKkXY9ueC9y
eQr9LufBxTIO4iommnJlulKtljmCvThC3ziL4AlDjO+AY36QiK9s0G4joL3VMSOY
X3F9D2yhw9DYNOw9D7NeSVP7rFEn7pdhp69bd8L7TLr55rNgJj5hA059+YbVzmqc
aEe2lD/6AxYqugkUkgdHLUKXkK8RZsYQFcLwaMVCvjVdYEYBcg37mgDpGNGkYuiv
1baJUysrZ/vRRn56KJcXhMN3USY2p31hMqS1pRWQcWlssTI9ZJqdtA92xA7/U7yS
dI3x1bN8KvxEGlwQ02qwsZuKhB/wMTmApzGscSsC7udu6NfyW9K31Kl5fATT/DFI
pKCnyO/JAZ/oM2Kx26hcfP7qBahi5avRMjSl8M2XaDLO/GeubZHHjYpr1x2qX31w
/dpmU1owt37RUVlCTyiZNHMpdcYy585h88r/n5qSdHDOJXiIvwhsh75iGij2h+K7
/gl+FS9P+VRCpcxcTAuzJwobj/UAfJ/jk4P861VPHV+KKQ2Z7nz2b3H0RV/M6dTX
cVBM64F9UWjCrXPMBy/ZByPRqxGWMp01tCJL0BuToQtFBecHud+1SqQg+HYHcfNT
g9GYCuX7HCBBjC8HozAM7JAjt4c2TQ8MAvG9afZE2t0+L188Vt/OKW5fU7iwLkkz
3JddAZFmjiUSUjnXo3duRw+yspc7kFO+Xiym/HI7pSoITRcd9s8ztGnMnVhSSb2m
ED5kdFLTQcdHoZh7siW5hEEJ+qaF70sTimSBuF0/tNNiYz2rxCll5H5FD9x/8kth
NIUOTSM+p8n+/OOTQdI3Gr+YJ36krY4ZImtPX+o8uLo8msn8gfX+NLHs3ctWpUzm
qslDJpT7PfIsC6u0ZWm0t6ib4P5i7hmYaNYcDRcemLYf0b08hmVhhfvbfFoINRes
9aZjsrIQ7hFwOxKCbpPPGn6X1Ppmay/fQCXvrbcO1cp21qYlE1EGvLvPYAfo32yG
eWZM6fgS7w+aWr1fJ6iBehvZJRyu3eNrsgIM+8BTZll6MMqBflRf1ntiSKS0dvHe
yffJYQRByxoTLYHT2Ab80jsWthKn866F1L+TWeXSEt6zs3jJ6Gv3LflzY+vaNYhq
PiN/hhv4UdzsxOUJizMxa2ZyAbH42TrMezAfp9XaDH0Y1uqgEvlDU0ahXAdHr8l5
3oP6OddoMC8WySGSUr7W4jtPRGSez5AM9ayVq3LXINOR3B8MUFvshLSOC6ZXq9Sr
dUwxx269qpnUoeErojJ7QSPdLFRWtcSKr5PpdpWRTnbc4iyuTd6OAI9DE7EY5tZ7
4K/IGUPFdknhnkBvSi3KqkwWZJt4eSa3fGDdoZ8kLQj4c+PO6UCUDElIqx33YLYc
RyzUHG9kEffcUHuDmVxd8hOEambYbxEtmlalIrNHtpTarWWxixCbfL1ArC5agOFy
NhxUXK2ENBXXk+zcsl/GK6lm08d35Z6BoHVkFCwlZR9LczCMeyXJr10H86hdOZRH
pT2JbtUxfc+jt8GqONi5ThIa+fpjq/jqnQiaX2VnMmXwxSTyX037gOAOu+KLxQ4B
KOckXwnGGCkCC2G5N98ytS8STDRjSnyoJ/t/hnYjUhns1io8J0tV7wEBK3koW58G
WZHxX+YuGZG3J8YXmQoCfvB9xQz5o5Me+q3UskxhCmFJ9GDEz5xMMtQxBPWy057l
knI0gXu5FVnOHu1Kvbegwr6U7auCXRyFy5zIzHJAjpAxWEWmp0N03KrAAL7/zo1d
B7XS2w3m5BreSsjRMP9cW+e/+L3kK2oIl7j2RKYuCaAXSOx4mAs8ZOQiOEmsDE9m
iW6t4BENP9Nh1f6rwNKcMpfdSYfRejRmQMMyCzDRWSB/kYs0B6vZH5MRRZEZgvre
PGrmJ5pXHADxhJSupV6toIPLObpKVhjT0o2/znWWxGo/I6SdkfCGTv3xDMe5Nv0U
hzv7nA7D0h79P6E7RwQ5WekBrPWWtP6mn7+GmSpQrEmv5MLAkbQSnw2GNB33SuRp
+hQMVFdfWkWJ4FTEH3DKrmut1MnqvPSuFlAEueL+Q7fpvRpR9r1ED/dcaUZQoHQj
dlDpwh0ab6qliBaIW5A50qW8QlZjEL8OZa/PhqgGAhTmrAIfq8JAba0bSHYAzMdw
reSSibkxOE2lyRDONB6bs7WV2cLbPtsP0sLmxeTudqCgrJiEJw7Q0c3YuT172+b7
YA5pkpXSQVQWtGQjlAm2V9ztMUG9s5WESFLIcIclbaoDzMXDEKgz5lbJ2jaf0ieL
a5D65GNZNLaaT1FqaO/gUpeyPr9I7FsPDaSdrRZ/VQ0h8XqGfOgvm8KKvOpAEbdG
KIIq351UVauBHuLzcmB52glIXqMg4gIhDsZ7hqd56bDz6C6LZEuKUFV7nOpBAv8C
e3tGtYykD52Q3d+N/bSnabTaAmQ2JIN5DOZa/hzuB86MK+pYC/vLmNq9me8nQKm9
v4eYCeH3PFGBjFS/uDr0upUg1akRvZqc9hyNPo7qBqkLC1IkoVrcNnc2mi/VbHKc
OvUqPKLnuZgxUtCFwraXwaKtBfsS2TIvbU+nfmSnMl1kdvfHtKLq/FOB5OPCBzoP
44xP8ZIVNrFPOoUN5Z9BneuWJdRAD/pxiFphBm+9FlTCfguJSNh9eDg8KrmLBdFU
TKaM46f1akkV8s84zj5feIzbpSEvQRclKVf/ASVeTF2zJLEAjxWoMaGaAG7AibIo
sQSK3xIuCglP1c1X9XwD4I6a/J9Bz6BBK+4/6mjNSmSpwUdQEF1c7Ry+B18II5H/
YFvbvAqY2lfnkKyjM7nxxugCLmEGR6sEO+Snzy4ZsJjKfHQz8s36mY4WnlHQPDeS
h6WmdQvm4vWo6Z5KfynAYK0JpAVM3yNH1eUUFCL0Hixhdr44tEhwzQijXkr4s0eF
lZ3mlgHApFe+Z0+VorcTzjbeh6Jjf3p8SEB14MN3h9DfGjxE1qMQJ/dRavtnELfa
1O+TuNng4sFBNtP+AK71jjLHWOvmus0vys6xTlqfq3VQ2guphOFTwNomJ8WMuY+p
K9vJ81A6zBI0bWCEsdIsLWsTGJJfxrPh5dx2RmQrgIHsoZrvV+ms2yDSKdlzE71a
vRuEc2rFy/BrvuZjbk79zEvrVLySSmP/UvcOy0Y+oLmsrvYJ8l/5h1oUB+GToK0k
NwEf42vQ5WgYD7GxPmX+TLIDGNH76Y4m+RwKbl9bJ9x4p0vj+AQtErHhnWcCqAlq
CqaGIVWFU6m5LvzKeVYR9gmPYOgy2TajCQhyCyb68BCrYKJQlK/l4ZQNBFgwNuI5
WtfC6BLubiXyDTSAMuu0j3iuxYHI8gSaEtW1ufK7is/bTAwyo4sLOmZD9OEKMQBn
nWC0Zbc3TJrDtPJ4MnwGqw1b9lmvDZ9xnDa5T3eB233zBzi2OBJhLmhZSgzLNOAj
BkOCYkBKTTLo/sAj9f36gUCMzKOixewToLZMyT3OQHOjE0fHzuT5M6FTJ/7AHAy1
/cK8aTX0iNEVMpw0BFxYYPyk1iXFRICqClgPyZqyuDU7o3kp0GWDcW2zUgDiS9HB
GfHrIahXtwnkFHKfAc2rI9NDLL2nwsgXsmzhs+wYaT7v4Yntulxpc7/uDLVDJ/4W
Ri/e3JiHtBMdUCLyVp4TUBRIv4w/d9+SiCRHxQ0v+C3Edlczdca/1ZQvLQthOtWS
5N7/6LBFAoGYvjLWQhAzQodfphknV2nxPREP40MrhNqiiqj7Y9nSl4s48XvGxpqG
NCXUwSwG9SRAizDSE65rv1gnOkoSoPpuLDcDw5faGiw8mbLluwdtZkSN2Qstv4I7
j6g9iOTYalRlVN7mDYefUzYjfGeDxsFsLG4i/6aNWFzlodnnqafrDiZ9MwjkK1Vf
yNLb53tDkGz3ZYNSUyVL4wMfYuSgILB3FyX9zouVK7chRDo3WwFC7apQjhp3YwJO
NybTHFbdbQssDU41mPfBVedpHwrJRDpufTMWY4ZTF5aL/gUx7N28OWdq/80vY6bm
wJjaIJqFHxOvdasPft6dFC/Iv91+XSgntQN9BsqUDk7f2AydHoV+yAvkdVnuBa96
QWM8Ye+QCI2o0beCci30vTZpaNYO2KlejfhOTw+Lze12CeN3WMvvVIIYjG8Hk2po
2iI+vyjLOv353yV7LiXtI+OfS82UJAWtvw9TPH7onWuPvjhvAlL1zfE+dkghtfTw
3BCLs149y45LVRrsbnAerRXGFqG+J9sgHWvdjYNrTr3UvJeHD+tJ4tBjrp3YdK+i
VIaYKzbCLWsi4zOLCsZMkFQdA19ZwmOy3yWpJCtpS7DIRosMWUWOLsHV+DbyPhsU
iIUj9Wj6TqAFvhW/WQ13guAUQmSjRMxaMlVqAZ4pO1Z0SMsmB0AhiueNdLeVxFqp
uUueWNXVfNIHwrDMrJ79UKEoftc0fLZkfCKTZbPu3hSRJr0oFnwAAnOSSzYpaUcu
5mgkW8Wxjgf+kQJwQSS4MtRtMccWATTSSqXu+KB2rEFOjRQSY8dksSp4CgzQw4w4
Xj9m9DRZDb10MWsfwSKSMl5WReRiwQY9qUttXwoGKXs3er4o/8VUGXJWvVAn6DiT
cr6a1qJDTwGPQskkm5HnGtoPzz0hDB7mjGr3Sep9pOz0uViiKZv2akFbyXE12Wv7
P2UzvDvku3Dwxy1+tNCJvgZObuKv+NDlxzpBeBLmeO9PXM6uG9//ohToVNkpo3mU
feJHeuzvQzp5YxEusbW9k+XbVkqamhccfg2etGuBprH2Y2GdAk6jq1b4GOTXWFvg
pJBwg0bW4s2dscorBSUhMhpOrw/L8JWaJzcBkUIiYYl5qRWf6y+oWupnAT9R/TMX
Idm3XAdli66RAQbK2ydcv3fFMyaTK8rEdLhUgDflEYO5ImbuimsIqrmEFlVjpeGr
j0T9olZOD+2LNpLFGHG2sk/dMiBX5/ZvCgYRVP/3LjATENtrcpVMpjF6+cavVIK3
l3MccaB0eWnTdaNn6jrq/7/iQATrV9ZucBDVyChHjl0eNts4rfoev4qrlCLr0G2I
nMe5Re+EriP/alMlRWPst9ZrPp05waMm+pcA3dtNl3nG1lxhzP5ciJ91wk6yDf7f
WVmBrw7qXDvbf2z9ZAZFl8qJ8X1BZcNJiHEQjBU63LuR+pWfcCjMUwmTQ0BEojjA
YOAvDLOf5XoZJKQ5NRFrwJqIU2nbyrOn05rke2O9y6NHX/uyP40sFEUQfqVyC3eX
vQRC4kCEK3SmaLuL5nV7zi+iRvKwbllzBJcu1nQ0x8AlFNoXzxdGNFGvmr2OPEfd
uWPypP/5vP6BqwcL4UDMBndyLckkRZbzrvb87guhZcQxMpVUO5F9JS1GBVsVdU5X
/3y+EwpHZgMRRsBL3u7s04OqdHpgdHArWmuHirXAaNCc0YXig4wxsmeqCPHYS6x3
fCPyBqsq0WT62Xb/qFJmdL4ZeChXtls3OapLurOLKMrhw9mWJgRC8PkRe7ZXukJ+
qYyAwiwm+rLV8gAU/QSCxvwYeLSRtSZD1honHB8rKN0AqlJ/ZgfqbQTre9pEdmSU
NKOzt+ZQfJLSg6Yp5J2ZioOvuhxYaZwSKL8+G+WaqNqaGlN0QY3wAOK8+N4ZI4nq
wkXC9JBOoBu1SCXoUunt0bdIdBRbl/DYBpDateLByWD2R8gYOUxeUtZhQQhCE3k6
semjAGKsuGW+wig3swhfguYlwfQkVeoGkeFnmXi0YRKjVZ+lybFzWoMoBJ+6wRlS
7qYO+WAbiRKWpCRNtijzAuUTDyeoBZEAGVu/LbgaT0rZfxTOMcEvTFwXuJ5gTJ96
h4KCJCPqzPzgVqjKQr5Ddq8MdZWhrof5bxCOb9auj4Adsz9yN0ZpMSJXkCb98RYb
hR9s+qLhVc3JVZdEKbFexN1XQcl0HB0Wv6BcdGCfpIVa0ppWP3UT7zfEvoLjrDlb
fIDPCgzN5RwOmjHhFmYNKkgMmAi2xLderz98m9VCiWVg1LS6bEJkIF5ZPEnTigCA
CSx61GyH9qiRi79kF07Apkb9V8Xpo569rD060GxtK7WFzF6fUh4m4FPt4bxzBJyq
xzJa3Wc1BUTQ9DPNTKAU2vBViklksv3p4eWbVeNlPSXCvc4fMY0kVB05x1fyflPd
m4FyVIk++OFBXBvWD796NEj4ccaZ2p9TIEpT6bV1lCSPhmLWweeUyIHDTpJHsK+M
J0nLN2IyeCqw3KXyA/PoTgoDaSHgZuAby3f6yR+Y4fGcbHZCjHBJXh/RLQWB6y9Z
7QNSf4/lFWQ8FtoNUbR1cIF/dK3lsVDXn2MaY90fK197n6F5Fp2tn0JtKrY+Jaj1
lzL3w0d7zllR+5eiYSECZOhvYya8Gw70Yo8Qt6lrqIZJwQkccylgWX0JNxA6ZSkt
bbn0neVLX5/exXgVBh28hRWsNTPEEuNyMzqquV+X5XNi06eSWDx4x4y/dlWbSEqF
ONS5mXWLtM6eFwFZrHBKW9nrC7q8onq4ltpy+27Tm4r+lueq2wQTDqQ6Nvp55JBq
5P10Ll6H/+9pPP/pwF5EYg/zVSeWiUpeO+U6qxwXs5Hdhka2b2JtME/BuSLL0+oJ
IHk2xtfz301poG2gXJveZdZIFQPjY7oV0P+KZ0Qvz+Pm8/Lmg/GzUo3IgOyWm4DS
iYlPr3SFw2O2Tf16zCziHO0V6ftzfiA4VJmoSn0gyM9eX6xC2vLV14pudJJtrnlt
ItiW5Vykli+QdZVdM79qe/QtQSxSNmum3an2FuV8zzPJi9TXQyTu7I7XSkmrclRK
kAkjZ1c9Zkgt94bcAko08ssBXwlvlgaHSEeUQXgr/hZmk+kxo9uzK1CH/60JA6VF
XBgqw9nzfh+zpwTnhY7D7x3X4VWCRNot/co/nu21IDxyJqKd/4c1uZnWEJspkP4m
B6LDwu3jsUoMi+re7RXLhiCCbraxg/RThvOas4bEiCgr9R+KHMiptVxwt0a3+hhj
eLg/zx3iwC8LtsIHJ4tRrG4LlGMvHkbM8aMhQKZugeXx2KoE+AcK2AT72B9pWaa2
csVeui/I4dVLtQgwxVyLPs0PgosPc6jq94buM9Q8Ql6WmGcr8TwL/2HWLKWXnbrW
STpTbmHVfZntA3zEzdCvfD4dJO+uRg5Z9WFHZWaSZ0UGYous8MrWv1CZ17fqePrf
b3iqV65G4JzF3Rk7qNZGGnv7d4h/c/3V2c/9uKiJ0BeUIUlSY5tP3nS44zJ3Z4Oc
S+XHXuYWnHwqC7OhQKaVO/upLlKzQmBPXOawZu5j17xYj4C5wim+K29tZlcFk2Rp
gGdzOi4Hhjw4K1r0yvBtVWEP/nJK7VdfBnuWO4i/zJ/M9GCeQ3+VhGkjRv0r1uXu
swsLdAUZjtKWlBYJ5rKptjYiG2NTq2fYLB6xoYZ0tJQ+QsRV2tjW53VaFxQilGKf
N5Nd9Rx7Mn8Ue8C6VSEBhYd8acqrQVAxqWimUR5EL2FeaSq/YKgXTEnN+R6gev9o
SiJ4NGGfvvc9zo+fIo8Gxk3CET2n7+1bWQUthAm0Ap45O+D7xhkbcH9eAsLVrZmo
h+JSfgW7/27o8vrTPALkXggUPUU017MU4yrJoVRGXbpEdKTyh+iIGvN4zPNAMCs9
Ii8Ocvs8fIbioUjyJvgYaExl7q/3YRB4vwpkM0M63ByUFOYUnaI6ZVwwt1SloWOl
c1dakPEgeowHuHH5xJnMkAeakwAsD86gkNll0z+yHvZF93itDH8K7li3Ap3mv3pl
ovDpHlZNW1zd84K5HgcIppCY4TjaOguwlsuNCu+54jveou+eseDacJ4dlb09WPHo
aR1AdnmJ+CPPrjd+rs4+sgGJOLUPOf5jcbOSa4H768f7iXrYciQUAMZekSOwgWIe
kyO7H85bjyNKEtB9UT4aQ4AHU1UYAvF6RdFrzFT2eDaL2BWY0kYsmb+Ge0uaMpXv
2jyTcWxqy1E5fvuUPaKf9oOSnlxagYVwWo62Jh8k3vMxt2a68W50QQ3YxSpCk8Bi
NVnqYYHlLgGbyBzELNJiIkRB58n1sy79dw7JYQmLZcNzAju8IsToD3hAMi0NG3Mr
Ku9L8xvIemmH/kve9uVM0R+4FANnd/2xdOzoH3PT7gHybAe+o729b01IT06peVOq
E3j0L1QgAb/hrw5wyctZkAKCyQKMbSSqynyqPt5A0Ko1Y07sKek/YG1QMJjZpYXf
TNpAwG6FBcH8FX28fkpQcYbcxud1Xrj4BYKiQxjdV3IiRnSRumjfNgdunFIlbkZC
In7ylzpgcij0Gwl34aCfPGG3nBEDjPRGsIGpLAFLjfMF9CAxrWWIQx+fge9Od0h3
QoPfOnuSxozRIi8IGvd79bJk3a+zz1+2JfAuME9LNz0u+FUjZPaTUYjMdP5jYu9o
1Xe6PgbsEm+VTbZ1qQhudKYrLRDCw+BIFjfaErjaF7ZF+a1lYoUjJr5rBftrskXr
zC55YHGpRmZ3HJoPCSH7A2zfJs3achIaPXm6t7/MsJ0XB32C54dC7d8TB2+8hAo+
arpQuHli0ZBmaNq0btEvjWqhd65FQgmjvEEJPpNHYjy4IWP/a9K7rwvjKXwP2iGT
fyqfLU1dYOJ19g/EqAnpsXAYjhTysfo44FlRAl3kn62AqL5p9RspoyFRe5WBW1NS
gdZBynu/liCkctS7vVG7j3b+rJNOqtau6nsLoU5LZUMrx3CqbgIbHzoGC65GTbHB
zAiM5mTGMva47Fe2jU9Kiuw+CZw3xZxXG6EUGUqWg+ttwWIIeafhVcR9iRwytu2n
JbuD8CEevW3bDXT2H0dy4DqpR6usVCMoIJCeVcq4tsALGgMcKuILBkWcFOJrB8UM
Vpn4hXQEgZAazi6X8yWncOFMHDVFCKEubasshLLQkbwS29gdO6GnOhc+pmsH68IM
xiVSsgtyeLETNxEO5kJEq4ndeaXcWedLXfflSVZ9qHDXYIMPifHAEMkBj2hLLtjT
/lPn6LRhd9J62DDZ72fKiFRwMvXg3Gzzv02Yg5zES8dvmMJE25e7nYhhg/Izbrug
7v8fdnuKvIjqU8UR883yePSqVz1OeJrZt91EHp222kAcdSeHwIQhvzpUJ4rmVeAD
eeAfd/WB0/6oX6ip6IlbO8LSXxHzatUc8SYY1cI4ocRTdQ/tUgDJeEmR6N2rr0/K
CHFk2mKFdj+hX3F1sgJJjoCbUa1rG1FWnZb7ku4T8a1POL0JUjailCDOr6cynRn3
8MUK3M7f4camdcUmuLiPP4bGv64bQSB5KOcOp7BOAfYbIjsOVhjPElbZn8TbUxNn
4R67baXxysNZn4n2rl9RAbGHZ/4s10qdPDvo29c7cnH7jsJvpv9mC/1p0/qH+rwK
qx4WDQ9XpCO2ITiAS81Kv9d2tx6my0uPrMyBkfBjdfTAhZ7WMQeydJCEHowiuQ5h
9Sob9Wj0xgorv1Mudrnes5VwMzY7tTyrdOam/j1xp48M8oWc23jI4OK6vDzSILBP
L22bNRAwnewOFfDJUnZdUsN3wSpMa5oQMVKMtiyFrPMNkK63J1Uy3ZSBMqhvYuyU
KcBzSvXYfY0/oHJxv1yPKJv8/3NmZSNod3kznnS5DJNCFOyNnsWSYA1hAe5WK7In
LTEODmYQlzdQNfBy+PWUs+lmxiBKb1Ms6miLLRVnkqzOsCBChx3SvbJS9jeCnhUu
SPG5njM1dY2DeBT+DQtrvkQxavdi/VkJzq7lv1V8Yx7J9daCK0fcClQNoUVAazZc
btCLPzP/HFEzEL5YBMU9P62rSimH37ZFHUPdds8y36YawJu60d+CQkUKRlEZT3fx
UXINsOLjGvc64ke6/3BGFkZSmayrv/FPbNSYn66RS/8KhUX3o868qjOGzJb6Hgcv
HEhfsLrEppp/IgqSlSAtWco+6izE4xCarTi41wDG1JQV2ri/fT+Wwwp8z7xUG8yh
Qo29i4fS1scKeuPynTGxHCV6u4zoV5PeGyeP5c/u/ojeUHmjoU52d7if1oc73uCg
7Ta8E0db3oFQq7SQmekX7hQzjAWURRUchfwhMy/fav+If4LeRX2V5b2Qg2fBpXbV
SDnK03rOP+XO3DkIQH040qBbjvB+4KfDpzEt690R6kS6pM2QYuV2VpPngJ9aFYn9
ekgeOdMc9Vmh3Dk6D7al84uycSlPY9gU0A6QfFl9SkwAqMo8s4LDfyMXkefmV03B
M120QzLWoQZlDIiEwG/dG4b42ec4Wh2jAhE1eJK5NR0O67dLsyVKkymJvTpKhY2l
6c4b4RT0nBdJXBE4oXAQtpo+a2HfGwAChLfc1fH4/nlLCDCm9GuGlAW1SK4pmfY6
ypP5Lsf76gaTEHKxNbLBXUrVmtkvv+9cv1MXDo/8f2/M6yuzDDQgJoykrCB8OTPD
fVa5dIVCTqJen45gBpFdVcve5ZQ3Cigmw01o37ZYzewb69zcojT39n4f3peRNQMX
kTNSaZqHNkpPoX6rcqinFjmNuAVSVL/nQJOnnXfqvFe8mN8feyeu/aXNOeRIc/aE
tqDzjsAEZh6MAfRzqJBKIPwqp30egf2jGm0juyRuoE/ZF565lT5gVqaV+Vvs1Pvz
ST8hJKtbmnyytmxiy32w/Y7ylv5qT2kZVaWybg3NkKDaW+2fc8rZwpfGL6jyntBg
ioHm14wOr20yjkNa/2yNp6OcqpDFZuCZ4kSDcU/ef1zrAiupWdSMxyGR8tYAeTgB
euwF/vnkkhdqJQPSv3QaUjAm8HdUIJINdrP/kKAbHEkS5YOPgNd1/ioSB+5PcMpT
CyLaInFbPMMhsMZzyJcUphXyO5aDSkmvLbMnQ1QsSXaN384fh5DoMyKltJmzj37H
cZrMauG7cXUS8OxvThcSL3TZ1065oQe1YJM9zXaNpkhkHXzmI8jyjuslz3dUMyTM
lMUsv0gxJQVahuZ7PgD/muh1hjxHurcihbKEho10ob0hS4Z3NC/JYPHeccx1M1r6
T8V8YOC14XQTnSwOdsagNx3DKSCMGfjwYvPKikhWqjuHt/gJg1ltxWW5enF2vUgH
1RX9yDtTn0XnXgi9Tqgp7jQ4ufKwEUPrdXMZPIIYY4F9Pw3udbm+RY8bDq8QdQbK
C/K7uhrvdBdM3jbLzToGqzL0zgsL6pwUQnt/2wPzC1N25HiiarhwyQmCtlQBJfTo
esVWrWzszDAVae5OH3Dcf4imaOQIYqYfXXujis9avurtU6hahdEQHWUOQ0aDjQ5B
UTBwzhL0BmcF0zphRJCrOnpoNm9U5wW+Nzxb/T2N04oy3RIDL5milif7FTBMeZ2f
AzFtGXLbbkAnAXibr+wGW+I7XNC9XUMBaf4rIVSuAcYkXO5pNR65IIPrkl/ztYBo
JgOAGrH7hGxeSjGjTTGJnkdL+eAJxSmM66xO/p7GCDEvR94jY6ZemjT11P7Ymltv
plsLyLbXvR+V+5vHVRlcQBKIr+/Yk7SGXPYKRGfTYtlftHSTdgoyZDuhO8cVE4KT
Px/KUPodxm512brBoPSWn7pFMf0HeO8lce01zY6GjQIHUiDhbA+8CpRU471hziG7
curyUweab5hIGN+ZVel44JH8JjwZ3O0B9C4OHktnH9/pNzoDrXE9XbaW5F1savOR
GK18qE0hizJcuuy6oR63+onwoQP0qhxsnD43j6Yb1ZDIa2QpZfYGk/GtjnHvPfNA
sjlIt3Tr3OYaVCMOSZLtg6yK0MKcgCVB3qSG5CXmtVunbIqIRoCw935Qa+zOajbB
nJ+cvTWRDPlg+6QAzen6vEqG9eqsVCrq8zN1Livz9CngEFmTGC0bFZG0JcDn9NMP
TKBwqne7F7FNYmXodVUGlGO6cXr53iNiSv6r5Qa1HaNcD0p34GvAa9NUEyQhFV/J
VC74xHXq72CWye6seDkDmDp1r+bKqRFl92GYZ6TGcqzAjnT3tqAXFyorE8DNcWt2
6DSuLqod1SSJmo23HXuCA/RMRLX86o2PDfjI+8yqQGJgYRnAl/h2kAp6s++epz14
acg7fy/0mfbZ8wJg6Zm+kxTaq/JvPmK19Av5UJkKzivDqsjVN+3LCK76+XbNtgOn
JuBbcK+P/TdWnA+3eHMJwIRjzx7jTshuBrLPtSXKfLMxRQtiRT4YqtpcPWi0mdpB
g1X29Bk3e5/jXXitu782bTJFFyw91NXbF1ayg83cDm5ti0a3jsppnHzXjL5LNiW6
XHO8az/3aLuPZpV4PGMLnz/56wJ+UdlJySisSU/2aEmW6jhN66AfYjL/w+gcSZZi
0Mf6QZ5R7uqX7tuPLxEujFj0BbZiaKv5fmw04eF+cqzVtlO02i6zUs2JYv90Ju3r
f/x1nxn43SucaDpP+cv0zeLh3p1jSoGlnB2yuFrbKGDYmXDDs+rQlAeXHwzozC69
KaQSdC1h/G3jnP4hMq9/iFCBhKZWGd+e6VmHC4dCfQ398d20eGgs7W2wJz7uhCag
YnDS1vpAOWFyBqbiFEodXQ/9NaLShbTwJFAmUTzN2h8pHmcN9rRnLzCFzQCmQnXs
FX6a8QoZHKZzeKdtYC16RToh8xl27wcxbFrxrT4LmTSza3+yhCDtmakPq0pHuVKY
V2/8fbgJpqc8kt2E4FrKhf0NmaLKkEaA/0Ij5k96LUupsP4ZzYjCJ2qaTj0hWcgz
izMrqtGSQk8fYs54dIpSPvoFfZ537JqBPxemEK5KJCxABtEXnLjIPEq3JxZj5d+a
UY8WTIepSfDYuiDyJ4qUACyVY9sJ7n2z800P0EYYgL1NSi6FHqsBI5Xmx/KlMAMI
hckVY0Kn/Fa/yso4/dFl5DiiBr1cKUEOx/TJNdf/zylfbrnkHEHUk+gqbRdCTTkZ
9mlwANV+oIAT0u8h2pi07ykfT8cughVxl295SEsPhilgtlj5kFdRkmmmiIO6U0X6
amzmOY7qo/dYM9QMK5eK0UUlR/UB/cTy+c5fBIV3PBkQn85olj7Cgegx9vPedETZ
SoLH4egJ/9zPlySXMCie6YJznGHeLlf2gJ9zL4dV9RN8YYZ8C8AHzKVtwaUPcNmg
PKD8mgkQblvpjVFQVCid4Gl6f+inHoBcZKJWTy01SXOGoOWx1v4qqABvxeEkR+Rt
BYtm+At9HEAvolNBfO9XLEUCiMP8v0FMAN+7Ytk+AKFrMl8GK8J5j7+bxt5SbobL
urcnyFWqQWCOD79ifeEPZXGxX8HiBPO4UXQ3mMbsYf8udl9EM3DLoIyTzFBvWmwM
EPbbhh5bR5FoZT2CB7Ew/dBY8wwOXCL3BXwdilLrfBWwPdduyXdr9mKaZTAawsZ0
nWa0QJO3p/uvqqPfH82Mk2t6cRKQk0JXup8P6kRCAFbDFaPzCuv7kGq2Emc2Hw30
GNAonZJSvkUirEngeULBTMnXXdd299oyBNATjnye061iPGRK61BlH8qsVMmNscNS
GxPbBtMpakc6WBF4uyAGjrqxmPAkgQGPuLl2WJTFVqGkE6EQ7NzpwI0iBuY6Z6Cu
q5mn8u/b5Dkk2jnwQ8W0yVSrVr1m7QUPDWMgxA1MDZZGKDE5tCQ7pe+Sypx8l02K
hxFuKZ22zyKcuXa20MiQMKxPL5JQQEPD1MNGf65jmGJj69NI+Ndia1lTRv/YAHxy
oZyyJLbDeSTqKzJiYYfNA4bUtedmZAe2uPegTn36h2qxSNpdeoZEw2LnJRkC9QaG
ZgAquwvEjHeBNP1qgg8Az3npng+UfolW5uIFIQtcQkX5VlAvncW0yrIeKXuOt/zY
BufmjsHUcaHg6ZTd1N+6NULdYA+V8R62yRJTUP8NPYRWyKjMCtFUqVJtskdY2rS6
PNn9LVBRhXJhDHunYrnwSja6Q+fgqPjum1F/7jcg6+eMzYOvVnQugeqZ3iD40UCP
B6BoLBOUhbZHS3ef8Nw79A3gA0NWzab77U7GhFdU9xKGAAedIUjlzWaA3NIaZ60Y
nHNfbuzbc1Agj2rV5QodosHScaYZnMMgGFBHBdYIwHqz2p6q7OJlgKkD0ehFuwBX
xV6F6t8MiCi7maGBmNy3/g8tSPdoTvHQ0iPgKHB454JaRogH5zEQaNUiZ1d40yL+
RHysX6BUuIMiAre9EM+ZZr3pJjMMlSlL/oZ4LfXWD6DsuFPm9PLwAiouLDaBxflm
VBWYskB2ze8Zui7FyYctIChdeSonnImFseZ/Srnl8E/P2MS64ILCKEymWPWiKpTh
FGda+sXCpnLOxTwbpy6ZOq+X7XXan2gkLrsREnMUNRCc4g5PTiuX5VYrgRP370Bi
n94GZksxr9N7CFq3zG6jP30RIJS4q4vklYPzmOXqbWzV6AmFM88NH2WlwCd4kVQL
SDAZUMrhYx5U22cv0k/DAXEvXxNyZXf/brkFWFab+PMEZIyI21lqCkIoQiXa6vQO
UlTUrtP6GREH9rbRGtLNsCAqzPuk28ZqgCaYesJs8Ab3jwazsuoL7AtNg80v9387
D/d4mMEGvxPUBBu1CrMQ2mR2mCl8vNL4nI13ZUSR0sqhAf2rH5LCgNYXaAppSaNO
KIrF5KcocOyVwMFXC2qqpB50wtYs2XQDAWLjOhQY4m/WiEjYif+Ou+EUjI96tZwU
rhBQ4ugNK+AS3HkxxWIRZO10FghsfVLl/9tGabJgXtR0VM7LbpbjQZIuiRgeXyLu
rFouVbpJ6hZ2HEpKjhhEuGTod1OlhEs8NFG463GC41ITcBmIYdSRmo3/lPodBc1G
k+oOSvHwi9+Akd2G80FtEeIO8+i0weTn20VCqwBzbjGlRWRtBVNqCZQW29rfVoeD
P3ggkpn2Q0lrd5TR/n7+AMueVfGZK2GfXswribcBpRYYCP2Q9QauYgdgFySUdVVi
gjugr2B9KkeYngFvFCJkNAEuh1XgLYQtIT4m7I6Glq87r0AyrZkJK/8MboTLXVE3
YUsWpzylUWlyvmdzwH4ZcK9ahNa6n9pW9q0+lpZddImbua0jeO1D5YjWixncRE+p
Gq/Fjljgt2yg7ycuLxhrUo/jTJVW7mOtN4wUPTMgqVNRUBLYXT0gYRE/JZZ74X96
mgZt8Gx8d1ihEsmIfTQD1zZ3Yn3mrTILYPw9NsrdDyXYcIWNdBxEhYTLkh5QtVGB
tICkvq/t0a1ucw7F7IGTG3+txvyTSWvmmaTgIZbjp4KKnMeMy7MotsGpG86PgATv
acZjk2PwlTTXMNzyY4pMz7t5Ll8qwVTdD635uPTL/WY4p3gex7v7qFkHebZLF/Jv
E623yf1LGPYxdHCJfv3GzeNPV7w2VWTie4eX3sqZ0/aQFxqSNC2aEQRHsySTRu1z
EC3diYdAhWgW8/TGeZx9xiTguZAicpk3yqC4LKijYkiudcjq90tBDV6pjJo0sutu
KqRz2b9KcZIxf93tMGtN1D+wiFkJ5FjBlVJuypk65EdgG/4Ok30PnRC7PJwgwOdo
mpmd3i3r7VofaK8fDFdq2p91TP1teFiGQw+f28x2BofcczuPnLR18xtlnmgS/lb5
sMkukVYG4b5k+f3WvkxqNX5Ql366Mrq1NmM5YLKcXncXj6leESqdK5gKFYnW+hHV
LNGQCVclXusQ4gHXWSqU1FgMukqOLH7OmyqTYuVRK+lydxn+PNBPyJLPXMrXXD9t
n5iSaRWdYhKO6EIfdN1f6xA5onNC3hUFcGuHNiuu+adQTyfEBLVMLNxV1cpDOKVc
lZh+yqO8UnJyEJ4w5dcnasRMhdjWEQa09t5zOjuqf1rbs4CQDnqn7c4Dz9Kcxz2N
POMPl3TrBvuqxxEUuszKQpZxAFla1cr0O/B+zxNsFON8w+KD4ohtRrldvtbUHDOg
D0+hg3Z+W3n8IPLSllQxj+eEzY7UH9259Qxhns3AI9lARUZu8S+MXfvy6r+3CaeS
HTtbF5aYAadKyJQzbzaftF+SzGeUuAVLATO2rKn39YNbTw4BNNtpzhkbTzX86DpN
G+6SoIJfIqUrA9dbIQeHfZ9RvbD3RhvGzL9M76Y0NqLjxu8Dn+2WJUg1jAJKQmEL
nuVDZzjCFUhWie4ZodzxzKWFZWszru4bCqe/zzZEafE8vj4zfyiNue7Oi2Z19gdG
mXg0U8yMiWUIly7NUm8Ypvxqwvo/xjxEiFrkfDvf996YCipSDIcEuTsnr7XR67b7
GBve8JsIZNMbDM+pcUQ+WtbsZp3f97JwYepelhwOXQA6grV+OCAcjKZ4jimgOAcq
4Sqo1vjGN3ZvxM1oPl1x4MQZx5YLqLoUvk0eI4HEDhYqTT71Ec8ShKq4s7X+Hx7g
bfUN75R5QuE5sC+mgTWL+y54GD4HpJyRv939Oi2P4jbY1bA84ydtSvxhg2BNm0yL
EmVqLjZjwH3CBtlVbQNbKruTdaIgM9w0bQ6+u0S9+k+qjMVuxaVdJLmQm4l4nuTR
olzJ61yL+cgkGCx2de/Lc58Rlw1rFVKGAvOQvrmTHMS8LdB7nMvwt7bP9Yg09p+U
uuZJsevCjO7u6wyfv+q5hwfvoUOqsT6iqb7CRZYZAUKflaWMZcMsD9i59ekJDuDb
fnLDE0PqjB/zFE9lu1ZaSEYE4Wx9YefQWuNREkTsG3/oSe3kbcG0VrRGWATNHL5u
tDDYRiKB0pFPh0/pmwrQ3dYq6nBztqrSss8AlyGvWcXyjGvONkIHuk2vYsFPhWsB
wiesivimjSWfUNcwklwL/NQhWS0PIuTMe3bRbBAfYLh5jyeIUnwF5wMPvFIitqt3
fncfBXfci/hjNWLNKmYM+M4+jjA7gIgbIi4e9Vl+XbzLKnMo9lsgE5oCxdvnEcq3
6NT97baoL4S68AUrkuq2tsaLUpMNGPmxEd5iMIgjow1mnvKkH/m6nmUxiLj8IspP
MSqEXcf2KBRVc1Kl3xXoGSQtD4xH2bakhrANkmv3cRv1/hBpxOWR0dBNS9Fw6gCA
HNw7Mja5Lj2L22SN6z9rZeYwvbC9d3Hl8IiXqAEHUiLW2nfK1iEITFNALWXY4xRV
lf5RW9vHazui8HB/CFZsFYFT5Lqg5Dd+8wlCALzGLP0jWH+7+HSNmE7GbaeRzJgt
AC81APiKnB5eT7ob1jROaeVk1tZ1gZsTz1bn5Tm0lSe6+6KW6GefQ5W8WaXkK3Lq
mG/LqUNT9HOMP75+dFMrdI7BZ4tjderDuaLR2T5p2ywZYIcHQvf6+YkUXUn5rkPQ
U8YAAhGV204OYZd0ABYqLKAsPtcQGmQ/KquCyQ1AEoBrGBHFvYRGNMSM7Wc/j3qF
HK1xYkxl7xnTfKTtsPDj46fwnonoVl0excLewqNVhLBBouye7EJKRpa4YIYQqXb9
j/FXJquXsCjJ2A/zqh1lwJM9xX4I5qX8wCQxYNA0DAD7Hnxjxy692edlh/dKqW3m
jmDvmJBkZWDTmv0e39j41kV+fWXY36JNgaynM2JS99HjRPGYXNBIs+apk7VHPx6i
m7cMZB0jdvlYawMCFvmtGL/rweVaygwEIEvM1dpgyWnBYp5Lt+YxrciGvWK9lAbf
OgCkPCfglzWjYG5ueY9Giw3Cu2O3dogwm4sxuJakWd+2uCCwLKTgrsm9zEcwc29u
E9qKkIhMbPiGn9NjM3WFmSNVHuwxYmapKQveBDr7D6h7eKBMbOJo+Mz2dQxDpiZE
pfaBsIQZK1JYykXZeCpuvgUDVrclPWXRInuX5SS0+w2fnK/LrKRMqldlFQ2nO0jS
1ZlsonLTHtWmMG5QMH8U2Xm1fH5O5T49WE9oqcNTW2hmksIS4A33UJNEdGFEAvks
oooRXF5gGCJPXUCEF6Dh7Vat8WIRasb0BKtWOrYexGcMK6UgjJckBLioljCMy21J
ntB4KRitQVJU5W4N6vUz/h4WCMbycVXyExx2Zb+B+OpCx46gQKDiCI1fQvWVIWmv
el1xbg/Wq0Gjm8nXakszqWAWLRLSycnZgZOLAl5xoS7ouAqZ+tX75ofggHZutbDn
ne1RoYlz9ZNtrESfszXblLySzGGXeGyZHaVS6Y6HAMJyyeZgbQjSqbWvilfIy+7T
1jGjqSY3MUOb//kMHXQ9XJhG1D08SG5W27MD8kbS1Zo1bbrba4dfvCC0OjisS6eV
Jd4Mfy3GyeOZCTgD9I/2brMcqxWIv4ZNuUdkiD4Fk02eRizkKLjW22a+rL8j6dvw
Hr6E/AIRU8J2K4EDjZv2fKfn8q77rG/JbOJNUef3EintKAZhazvTiu13pL6zhflO
of5sljLbT+53sFqYttBM/anl91v+5F5EHfkPgWsJZw4BG1E1u/6b4RiKQoc8RS7m
RbGVoJwdaXlQ6sPHiZJMVplzEUzWOrzlqH/7Zlpl7qMe81YlhBJbScqdh5kwNsj3
vdaCLkaTBsgKVFJmmIow0xFc04Kcvniry4DwM25Xk2R/ehyoKa2nbXurQRYkQxvk
W/oNA7Ua8O/UCqrukAsCJb9UcPHGnKUUu2wo/xSfY0NYxg9RBcpWH+iJiP1R/8f/
bSl5spr1Wd9BR/63Hdl9iiDJBWGB+ZTahBbM8rfRPyAS3mFy10Sw3A+vpJxTyJ6Z
qyi0YGWG67ECdQ49+acoHal+i+3h27SNLJyWd3aKlLNYBS1h+jxyGCZWYIDoSSz5
6q+S+4wbqijEew3iKKYz/eaoAMFLLMNRNJyCf/UBagzBeKIEdSf7JNn9M/JWaCSS
xDfgJ2tO4/3vG6z78ob5yUT5Y4C9ODfO4LLHd0x8HAx9Ux4OMv/aXP4u34KaJQiU
uIQjVJl/N4AJ/RlobVY7mk3Csdg+KyUPflYN2qJ+dH95Laq+N9iHABiAQS3W29x1
TsWW60Sr59Wp/2W4S3eRsm8xtu5ZvvSRzo8STztcwVRckn+C1W0zOpXgYO7XqEBO
r8m4EPs/V8LZOGONe0yfOmhSif46aXmQl/CpufmNML+X0m2rQMvKo5/jwRqGYHam
70QuX/ozAAazJKgFxVW4JAeF3ql3gbFRl2OlVQM1ATlmMjOd3BkKmvXOj71YvZjL
DklDZYIa85O5wf9T/whoGuZtuu2SNvFxRR0pSMyvV1Kb8kFo461V50sRvAYS4rcc
Xw21lz463YexU1H+ixtl+0lf6DOmfbxwh2yldY4syB/ceiGwKcm+OwoPTApC7Thh
wv0mUbLP/EnFoxKs5pX61lnkqr7QywtEvYLNk84WkQ/Z3dpag0Km32Bv1lHC0ThP
xl41FdvZbHpohuI8XKd5SR+1uDgFBMeANT2dpbSipGetAEBTyAwsw7CKA3YqzTfU
BQ5crb9F6GD0sXyO+fkdT3LfM40mftPtoZQOdStDSyyLiPgCZ9SDKdLmbmSLtV+m
8hQcSisK5llDhz6/KlT4Hpr3TNrkKSsnJvfs0Tp4hp/WTxzv67QHXwynfj4Bx7pe
OHqvTjps9UAuSav6x506GX9QFejcRYTes4wyJSNNzRKnS+R3ZX+o4PATLmNt+nKV
uDx9oASAxOG4XzIkJJjqPudBqwdgbQHDOH3D3sa3rW7OKS8pRaFxQvyBGdxjulWB
HYOQNYtZnvMlZlRW+GzBRHKShW5doBACmfJi75JDSudA8tlmBZOXTLkGdl/ltwiC
cBTlOtwrD0FRa9onYJNx5EdUqAitJLcWUtUnnlFETwhJUII5XrHZc2AcWJaDiSLh
r4dXnOD7SnteL7bNZTlbdTEjcibtRv8LPgsFR5gTVNL12e9gBU8P71XckoVb1H96
fNxeK3rEAvuH9bZNq4tB6mTXZn2sIAEx3SIfvH1bpflp2aB+gxE0tp8w/yt8+IP0
AgEw83Oo1wRX2nFmWnvp141M27B6HTQG1g0B26u11oqYs7//JhXsk6VNZSu33xS1
3fcQhgRuQ9vDhMk0FvdUcWjnmqgGJTNPlWRCKfO+scxFhqUm+G0t8X4ekZrt1TPB
EG/JFLWyDUSAfCInYWmyAQP94liVmc7QsCT8q2v38n0QCSND44IQTbQRgj9fpDzd
0boi0Q05NiPHSM6RnQJ1AkOU9w1az1oOwN5uNYG0VnKInPxwW+blPL6a8VmoGA5+
MveZIBk77PmJjUS1lw7iE+hx+cRS1bt9+nxPSJZHve3X/VyLVcMd7FfMwXUXi2sq
Alap2HPhY6QWG/CIihnqN1fzj/hgE1S6lGyRMhGnXl9JkHuvD3zpKB95C9JPm4b1
2wulvr//TdvtdrnaNxGwVmuFSlLv/ZdxA5uC2++L+f3u/UPyq/Ren71jZrU7tMPT
Yb7MwE0Ddc/+ctVunU5kg70M3OFF2Nh4gP0HPaq3xF7CO8RTUd3ENjz68lVe0ewS
/S/cOYEuiCKs0tu8QgVUbdDCPAJcQH8P5dFVybr1vGuxAoKa91+bycJozr8QKoxE
GrsJ+EU7FZi6ATe3HkvSnhakStLui14B1IDKxoxY2S3Ctlw9hSUwpRa33Kr10Gim
MabxEpc6ofWBebzm43HWkR3ZnVRQaITH8U2q0Meitc9aGjwIntLO0IrVhKS5q9Xd
zzfkI2xkAMI6GbVnhZeHv/RgIUbgoB0L3jUIh7KS/Bk5Vc8ZmHTaKM64NPVScSI7
YFEYk6hqKNTSKbiEPkUcMHcjJSDxe6HumhWvDFvI4f6jtJOGHbwYnAhFK6UgtqEx
oMak+6rB/xTb1YFeVuGzAhjmK3TWWsYHkfxuphCXL4IpYkJWV6W++tExSHWCrlVC
l1Oq4AJM0we7KeUsVMMvlwjtZn4+Rpz0vFa0tU5JKz8wbVSdlxMUvh8GOs3oYP02
3li1GlL5hCAWMrpy69BKXTnzEX+9TEY6GIHaXSSzpvfefSazmyvKBQmwz4j7XZAv
cgcX99DUKtR+X6HfUwRSpSP5fm1UJLrn68J4ElUAxju+68PT2GEG/PPBi1Facdrk
G0BZ8ZuoPsnUSqIlxV00fHvlcna3DCMCE6buFrgOTk0XEpLNxTIoeoVufQOF32tH
Fo4+6985HPQFwq/N+hWJSl9kEkFSXLTjfJX9EZ3HnNi5ZFzaNMlCrkTs8TDh/jSy
nOhlpi92xK/rFgktMg2iZ448aMCdhRoqNM8hLQz6jxc=
`protect END_PROTECTED
