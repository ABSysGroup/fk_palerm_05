`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
obk1dSYhwr2ELpFIqVARWCpksJ/qW035H7rkp3O42boVDj8SkKzDW57x02h8ySCH
UlL9F1TmhxT8YaOu8GkUB/lR/LaiiucQCdWyEpZj5EWGX37dEytwbFOlJEdk0I61
2fdxoKWrcDrlGj/xs6G8eeDJ2yaa++u81hAZyJnSWbMsM4eZTo9tXNuz2pO4MfgO
Iv8zxQzq+v2cYvUG1mZoX/lbFsig9bXlc+vUO3f0KFgKG1gOAxugptpc4Z9VSJMu
05tjfjsH2vXxuYkdsXu5brzHCO0320b+tuMrMQRBfnhN6xyRQlL9yC9QpOCXoBOo
JIvq5xfjEZNhIE7GNwnuPI1W3xzbBhU9MFlifJtfoh6XyVU+jk7n55MxDxJk98p/
NZIghN7BQUKJBRxJDpNTJqU39Rj7pHLYV6+j6G1L6hp2WvKn9ECd8FxNgF+OxJEP
GLz+RX1Ov7aFhVQOSHXkPw==
`protect END_PROTECTED
