`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l+4yhIE6RhIf6IrkAhQdsgmf7OWCit40qJWr9ADpWCwfvuPcmAQt9rcbf/1rxptp
uFzlVaXznGcHEy4qik8gKqK6/ZXM8PoY4Qe4aOP/SemUADxeAdoNj1FdJry5Y/lL
LO/+OlcyG6XiCPgJqTcDm2A2B85D9BhjysXTu0YscqHAv5Lb+KN+srT7N+NCinIE
RG0LZwS0bx2pcjvJBaSyu5RBiFN0zV6In7ZBrEYWddJfxWyisDxUlwm7nNgZ8/46
+cQE1nxPHa5KVnoCJz6L4h3ia8D+O0iDv9RRU1k2dVxfxad4xagX5DHY6JbG7wuK
khv3s72CxhmDR/ZZWhgE2M4YWmXS9LIXT4N8NBOVCuey7WipQvAVJHiA5k2W68Or
wyVSijT+Y8RkbnXpPYBcgUNj43cBKwYEmu/AeN4ODDRPebDZAQvRc736oL6yljR8
v2yE2YtjPjvWrMOo7yPu2MBlcipsKNCmD9ROGdgP1y+X6j5rFuTXntwE/D/F7je5
aKw+Sf8+h+4fZzB4mCvF4V9e13srwAKF9oi/1L0AXc9gxlZjzQKDTKiGARGiDzu/
Ja497hkN4AyyLmuGHxkiaZNdPBLy4FSU3m3L1nTK4cF4QyDllvswrccC5OAxwnKU
Pq4a+hbn4XU+6uengtAW9vtj5cpmQfvC+5u0n1oyKkvLBoo/EK35bWKaoUlpmtM4
ebHX5JhwRzByxpfQRVAqq2x8PjOQhyta16y5SL2O0BbAWU2AtTZG+CdX3/gSWbE5
S46i4MY7pyfZfxORaB81R6GzqqERPJQy0S8ZNnr4152tCtCjE04+pjrfaB0uhpGn
aPS7hsfIqatwkCP0YfH1Mky6CA342Uw8MBWe4cnH552ZpT0ThBq5yXCnuYYcvhC7
yc0xraWalPq90PPkUCtdj3w7IEJO92m8E0KZctg+UXtuA3kQIqymArf581FADe5T
zUHkG6HwCNAcwjvKn/cPPbkMzeSjR2zRv5o1i+ErlpenlFWkU2Ff7/f/883dxhLU
of3pxf22IumzvQEDjXHD89fiuzDuW96uSmUSsPIibBtm919m/sl3YAtpKHIdQjkE
qZ8y3R74wh2SSBf4ufsZn5S2H91/Eu3gFxRPhXegb+01ATSNwUCJkYyPgQzpbbpg
YjqvtMBnRkfOyScXpM7R1GY2Idvk4/fg6Ou8HdIAO/BH7Uv3wunVtpOgnshpql7o
p8Sdmo66m9b85WngpWlcD4gqvP5Zgk/bR/N58vz6W1/FUT1QnoxiG+9wKz4b2CmZ
G0LCUgQvx8Qr57lVXDveyN/WuFa3v4jcy1lSWYiL+olXVbLxx1qso1T3J7eTYZgi
nqVZbvpnEzxQf1UqsZmD/8khK08vTAwmHR42P2hwwhvxOvbvGn5LWyRTTFp14o9V
mieJS8MTHKu2iLR+zC0PZkX6g5k3otmJw+7HYIImwPrnJOOoxLf4KMUYOPVsXLQq
PBEYGAUgiaA3yoE1GxCnlh9OmoJMi5kme4Ytcmdg0VS7t/jkRB4ee5e92OI2e5MM
I1KyHyrdXLCMfUkM1T0hZPKvvNy/AzBOfPzAyYqYnRoV6DE0EliCjTRj1lXRIafF
Xsu3uZSe1IAK8uHPPcwaY9rpeWFxZ51PVJ5Gw9T/hTnpcxtHjQSjbdwzDtWE8DSa
zaLhmKHjC+ad/f3tdgjEM7xnYdBalR5H6nvQlGeCUdq616O7HhfKCW6RyGspfIgd
5kS+ehLbF1nsq6P/3PVltm6H7l+NOyQJgF/lJXHoi75jXya/hszDecsDKnq2hjxD
xF9+yN/tSyiFa0dHs/K4zqU2sYBBkrzAcYupEuuIXBZaFmvDeNLyLSP4/lc6WKAI
bOatw/rcBwQ8XaEcdwjNz9WKDhKHK7pcn9Sl1Gg/sAo2obAT1fqjeNpKGVSjBlMY
Yjr+TRw52zxQ0EgfH5RE04B6mfmn+gODDY/GQnT90OEAyp9gSqO336i7h4LYFoMb
3spXYQnerIUVRF1uE68b+aT/ioNFl1R4FlVNoZNRCog1pqsLcRxNHWhEPG26ZiK1
QAQp5xQjsg8YJ0AHJBYGt1cttIHaK/+3pZrlqrDoskk8BVIylHgNFkZzkQ2u0QGq
CuPVrc21KeFGxoqkGRfppXxjYxuFfPEqUwmvVOsAzyc=
`protect END_PROTECTED
