`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cz6WXqYckyXaJ3W2Ll3QF5L2M2q4h2KDvQpzbhrTWu1XfeYB30iNTy0gKkcE7igx
dVwWWVbwtMZUmS1xW/9ybv8Ske5eI8LeF83rQAIkD+18X9m4Iz1yIeRcg7fQXzZQ
34QpV2iuqz84PAWiCKFufm4NOgBd8uOQ18NRg6A3p0R9JBRK2dEkFes0bbBNicNa
1aEX/gGWQ4N1CTX4AMMKtGof7zfwaLsS46pgezchcP+hnt3VFDe7GAcgkxwWubvU
cDFQsFcOiUln91gKHQ7r0cAgYWYRu1tlqcxSaX94/ReGFKtyIH4P2ggS/f9inzd+
JDbwRTikXrSYHnhjni8oELLPW9hqBPYl5aFUf2WsISUEPqL+p/Amss5j+5t6Rc0V
WVDeQPwviH9AlnXEdslNU42/dmjkp7ezshvcATj02biEXMjCyqYp1zzZWJj/fXsJ
i/CfDyYUx885dpifgCk7pmz3R/k3kPirho1ce3qCCT//y8rLirpStXkqQwmDx1Kk
`protect END_PROTECTED
