`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cHAgnIEw7lsKOU5wzAqgs4pO7gq3uanCjxX2CDP4iPuSe6MaK4wTddY++QArMC32
KS3V8OA2DZWGPjlwT1ArhhAkEHRSCcJ3s6q3oakH33OkPsBdzqN5f3xoZY11v6u1
+Ha4kZM4Bd/Yh+1Y16YSviiMeDXmCZETIR0HogeeyKEfdUnnSmxRlKiQHg5NC7nG
cUJ40+s4lvMLIg5eDhAafuGHGrQeW392osVpo1UBNAOQfsFEciqct4m/DCX8jjNs
C/FVh8DTbtHw+rYIQdv4MhSoMJXFtfXIDQoED6CkPxon0VXYRW0r0Za8O6kCJsfb
Nmhq0t664WbpJKFGIblDu0oPDSbm/CFYHOrXZ7fmgNRxSu9yYX6rEkOrL8sGjkRm
t1y/x/HQB4yLIoMNMJXCK3jRJGDWRamRYpFYtImcLM4FB6/kWoileydKHgX79weo
SePtiGbQNjqPzz0RXKD9h21HZzpx019P+j2RpUOlMDcEa+D43L/gpztAD5yHw6TX
7c2JiVuMFHiI7shovw2Lx2q/Oq5SvlXM7h4dBjpcbv5/py7gNTnZZDqz4mqDN20u
3ETEah9fT9LfIhMqKzs8xuzgkMyvEwnyk+Ic4aLdNN4cpeAPTU4Mhb8u3nZt/U9U
6/HzE1otNeWCez6vzrgVnqwCo9+2alifTZ42O8h3ZIzMyEyToQyZCLE98KH1/dRw
crR6J2P9+bCpokW5Oq8kVesx+wLgS5JB1agPuTEZn8uHapPOX5DDCkiX3z4LNK5x
46MLgJc3piUW8iB7TxECJvCulaAIg/WD0+8NzuJpZMJtLWD4RZXhusfsiFw+XdSR
wyw1o4dRHKadXX8HqBiuZtOjbrh8ig4zAAPaw2wdiyHnb0ygiGAinTcuRZfce9zA
SDhdBAPapFFPxREaLXyuf18cEYXUPzz1fN5vKPBzi3zaQU8oNBmUhuAEShtigwqb
b5nst8oH6eygTeAwlFqUNN9dEtuNRn9mZlhwGjGMrEC3Zala9WuGQBZ79cvB3pl/
pWUzJ79Kv2hhaTQqU5Tv/dLC1nCMyCFvgWQ50C1qVnK8zSf9tGII/lX7oQhL4PLG
KfQzLw3tAZzYVZGQhfoETkW8acxzzGKdux+N++nCNjibIvvi0YfugeFeUiz+vbUw
qozpCOVVG0R/LB45a4i6/Ri2bE/wTecmwSb43KQxq9rKnjnnTRKI2Sn7eh915aw6
ied2A1SYVyu/h1NPpsVvumXxnfy7WLBSMYt6bgfTkAwY3rt0QCt84ZNUo3DfbxEC
ZOAFIFAS4ClMDMmnl7o3IwYT84n7Kj/h2/6AwBvPMuSgitudUINV6ml85amc4e8t
eFHouQw3gkpb6Do4LRO8yPOD3YuWeDcAB1YVz1qRng8=
`protect END_PROTECTED
