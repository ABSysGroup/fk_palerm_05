`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kwVlCFYA3XUfkdJADNSi7/5U2TLmngSPoJDzzbAq8FA/ES75PsyzeGv+OGfstdEp
ZtvMUXFEKLuBbSOIgGCrZYDEET2B8Obt45w/DIS4WvneJ53/gMdn9bhndQ5RcpLJ
7LHYnxTfzAiOHb8oZ2LXtjUjKXgzP0rKO40qdg7QiqutM3gDEC7O5wzbgySmQPRa
lzsCns6j4pSBffrh+wp+KO984S5B+Os7B1ai3IKV1BxaaayD6xF2vUUJK3zE7kmq
ScS9Nrejd9+ysKP6N5eEhHuPiacABzKbXGfYNeRWlYlw1tJeZecRUXpx0CbUWDUT
PlxiLK9irEA3/1o/tMv42z1u0tMJkBDwBhuwBR/WAn+m23KFuO6VkcCkJng6+bnX
YlZTvP7ay+/mN3pti6NtvOm5WkfhC/r8vci4In6oZYQ=
`protect END_PROTECTED
