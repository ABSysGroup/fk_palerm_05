`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HjBFs/4RPPqX11mKPHfEpQ92ToKnBCT61zRUQ1+hpLKp0rbFMr+LT6wkOZrLc+Ex
gApPQPTZrkS63ZXEi5BfRDvaOzd/ksDSY0IPvM3lziB3hl8hNJohA8ZZ5YOimGLE
5Om6cU3SIxWtTQY8q55cp+O3nOc/178dKNQ6Fpd6YQqG4OMi4aoGlHsr+3/DGG55
1jfa6l42LUcvr+LHeXINH1L9ZPcqwGkOV1RpoOWsnHBLTD6c7Lru1Oh6W3KEEo3l
IRybom0YDc0IvhOYUYYBpcpEM4Lk59teu+m9RaZ28T39065qR+/7hQjNg96oGZ49
xISDOwE4TtROILRqwbM4wlixOKBYqifNoE5lvkPZk9HOmiNkxie27k4lPfJP1i3v
5uxCgzdhWL7/HtgKRPKKPsJB252/7X9vrW9ATJEC6db4Ru0wG3b7uZaKO5PcSv5r
7UCcC5fd7zBFXW+3m2R77e8DM9JE5+KMPvxdHfat00VdxzXnqXBXPnHhqd2R/9ka
HjGupWDp9/cVGTmZ57QVoAibQ+lEH00ts+oIFgAzAI2e3rN+G3mFA3a0t3Tg5lb4
2JofBhhLP0S/TY/qQ7GUFwZn56qjczJ2pr5XvyBXU60foUr254F8Qrmet66MJ45R
BbgG8WgsaR71GsXnS0M3d7OdSS16451Pu42RpkcP1rYhSTq1Z0gllONSxo9KnHPz
NALsxJvx7oxnkv3QXXwaoWlGs0jvvLCByeKBFYY++bIH2uK7nKMlXbUA3cDWECOG
cpi3JKGex4Xa58qGd5whLNhef8n8I6MzFJrH7BQ0PWY=
`protect END_PROTECTED
