`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XeWCaNf9GYfXCwY6XwAp2ayZOZvZYsRWvaLMNSN2MJwcSkDK0VihKqIfn48IYWIM
8gU2Q9sWSGQj+KHN8noe/bnGXVmavSqenbZrbzYy08CYyRLKbJ6NlaZ313w+ZRwY
OdtdYflsRLTw1D4uwg8lqnfJsAYgRKJxWSjfftOWrbonpxtbLpxemqYjQgyU1nWL
oa04HpfYK+2cCtmOc/4QQEs6ILOhtL/IT+zda7AV2/DnGZLkGLHCpiMQcbD/m2L7
WBY9z0D/kAqfPDpY1bfPMpXhU2cRMKazzL2cNG5FzVoNI5BL5iyiyQCjIVrdK/CZ
OEQPbhssIVkspYtaUjlGGA==
`protect END_PROTECTED
