`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GKferL8+n2SJ7iz2cnk5LSQScjS3ODz3EfyHw6yFC++zpvt2aWIQYax/xgfzw6x0
TL/F2kkvdCZ6k7TahfupGQs+CjJNPzhYsZWX5kL906p8EbvnMpneONuLyDXX3TlK
mxroKHEx0KgmGkzGqpi+ojFARMdbrvZC+K1L2gL6qoE78P0MwU8E98cgTn/ur0IN
p2bxscHnQs0TWNhLj7YIwLJ1ZYB2sIzoiZuCeur/u9ZUMZzjLZ1AZpW7CC8k8WvZ
AON965PEeTDRXrZx4EOehw==
`protect END_PROTECTED
