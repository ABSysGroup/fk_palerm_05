`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ti3MaEZuFs3Vk7Vdh3faUgS/ZsY4Lgx8JXSMoVzzBfHjJHvLSRpD5qKHO+nA0jEv
t6L/GrcuvEcfkZddBuHLWz0iGrCdN8eOieLkOT2gnhGzT8/ZJp7lC5secrP5pvZR
YQKvqfWMyIOhd+rYDkvxaEigYPB3r7+OEj4bvXHmC3YKj76BawDhuaH8rWK/ML8n
S2LJPtdOzCKQ1VxHCaa+Yt8l41AYPk6mhMB77ldZLuiWdLH+Qwc/t5P4a32xQw1Y
5BhMBzzQ6UHf8JrZo590eKp+2VVZHhcLyeQDVQxFLffXbzjhj6VFvFPQOBexK56L
E8fOwec2dCxiAXUZyTrE9p877tQmx95Ca6yV0vWvWWY0ree1pneY6juM1VTVEMpk
zEn/mu8nxmUwb+0+KAbpTptK8oPlDWsLH1I0lkSxKQA=
`protect END_PROTECTED
