`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nXWRwLWJochgNWOhpLoG2INVKlmmk7fnJ+wyTJ3eU57y+XopnDQgDIMlbWHlFx+9
NmSc2U1swjXVSpR85rfky5nfUfE5Chmo73fMF04Ld+GUgGJrSkiEIUVWH0FIFRDv
bYFraFgjK+LPnqNWUIMy9uRzIaa2n6C2fwDeRlGpdiuEiApWAZ3i63OjP66acn2B
LgPiMFwUXdaz+6KJdPmlY2sobxKQgtT3Q77QeYQIujIKv+niLGlO5jRlF4RF+cbR
UkerpVRE352pCJG9yMWbbbIP28JyDzQwcoGlAY4b9Vg=
`protect END_PROTECTED
