`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jqGWThX7nN4+cHiiq/EgRYDLrRMAbeelzBRrUAOJ+9fDhp0yTtcoTxCrDo9wkgmC
wjVOa+q3SfumESqJfZe7VQlEs46ddiXGPGMDMS7aDiYmEmkUyrcJQl5qXecBtg4N
OwfH3zcO2QX4fyR1KWdyIOoAwzCimYJBlN4u9bhfg6oEk4tIqPbNB/iCBco2OoPk
UBXJgKNVcUmAAStQ3MzwPYMYBVyKFUPlGIVVUOMYbSFnc67aQXpcIOvlS0ygGBZJ
IeTjwvGErLNeDCze2P4yXKdfaQ0UvBtF4Ut0B7xIAPSLOWfloHPQ2oOgz697LvH1
Yv5AR3c5XAcZHSNoJYMaODgZIuiUsv93f+I05T/jchh+SimFDRixp93DgLPnE+xW
+CaaWYGdgvvkOrf+KkFUIsHmYMeHoztNP/be+MlgtGZCus+UlIj9mb7wSM7eCYvI
A7qvRqHAntcHK+F66rhsYvo0Iu+cFqT8/BXAY4gp9RbwEzSpf7AEt8LrDOKxo7iG
`protect END_PROTECTED
