`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t6PJYCZLWKRNA13mdQJ2B8WOUmsU4wUdzY2c5PgYQcoG8mTQdFV0sf2rHgxwSfXs
qOgohMnAUZOLRMBTgS8FAsG0BGYit3WKoqQrIFBgTkxlQHIabw0r2wyDXYmrORpZ
13H2orCqIrCYVgo5+ZlF5cQ5LKFZCHBpA5cUxyo18An2ahft3UOPt5bA1g2T7+uG
aicR+hLoHRysbbTau+kLRHO5jgMMk+lXj2mEhS0xY0tka77dq9vXqQ7udjFoBj65
xPknuqf5ziEAO5eQ7MWxqqoId0MSfIppq++eQM2jcBcKxJWN1G4QxxPsfuE5CWzv
szQuCSmp7bV1I5owPmp8/4c1+LrX6aQ2gN2fRsmZVYzOg6vGQwmGB9O7eCCO1YjR
wTJPtF7PwHnqvYWBfu73rmwwkNsv2v4fP0EVOJ225SZAHyMnrn7HTC3yYT5BfTIp
P8fd+J52VXAWDNs/bualof4ka08TOOXhOmywCRuAVuyz9+oQ+Z4DdNOrTs+lbFxe
MsAEa5+Qk7oJH1PylNCC9gNwr3ez3PL/ni+bZdzNxx494x0LhbnfQTTt9vsfDftt
`protect END_PROTECTED
