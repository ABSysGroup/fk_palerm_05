`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HYRgX5FgUp7w3RJWc72wa/ApPHQHj5WU/lCZwrPz1ORr9+QXHFhEN3jGlMByQqaH
1yuc/H3qhB6ff8Z8aUxz4kCps6/mGyuP5aA7LgqHzEu5qAvmBI2/nZuYj0q667jW
Rjv+Vkyr8rXlesNKbRNHqnGAVZjBSTI8LXYok2crYg+J5rHvRJOQMbsJ9OUqKHyG
gEDklhBIN/Qv0pvJvNSRAbwMHp0N5wkfp1mv4Ef4eA3gzrzLyn58yB4DmMx7MRLx
+VYEtC+VD6rtyEDykBJ9BZ3cmSWKJ992lw23W24hSwbSaThovOuv76mov/9kVu0r
jwZtIxsuI48pmtsETadOHX8/D4MkDReQHvu5ReeCXZ+Wnm0/rmxDFSZ5VKta1sHn
3+NiNqF/EBtlUpeecYr2SxIiQLLiBtUBbN7UCB4j04sB/sq7ORYKZ3Iy2zwKeVTv
/33nZCwhVK9ti1U9FCzPktzcKth2oJSnbQCt9yUTjVKTI2+y6s2b8aG6fV5DWpD5
lPcfxP8L3ML9d1Z4mspwqjU7lGHK1U7r69/zUdlP9VABD6V8dfFauQSmQ4mnxuMr
gCclkZ0f+6xb2YjvlaC6aZYrOt25RG9gDfi/ms6BTQ5whNS9fNfPpWp3fbw+uv87
9dYHoKKa/gB40etDWeXrQTwkkjKbkth5g6CUhnmwzbrM1r/cfi5NlwRjDphVUK4X
q9NR96ifd1pHgy5aa1YkoOVAJ++4iZZFLkVxpyFiaF+TcWCUqfslKGZc4vjbLzGP
0E4Tg3WLDkn6U0PX5KQcUZJolt43VBaT81TAltEt9DjqB4rISND4JBmwqmDmDwR5
zeo7y/BgJ8Y7NWbT2ZO0zQN4JGU/3V0WKbW22FJ/q1Zby0ZJwTgTDpJr1vhIkhtx
hqPZFKedf+WixKN/7WYFPIKFJpZl4p5cKZoyDDoZPiol7uu4y+X0Ms3luHZTA88q
Xu4WeagjuvobE7jOIxPMaw==
`protect END_PROTECTED
