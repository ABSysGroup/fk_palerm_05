`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BTyEzlwR77ze7g/lAp1iboo6eqneB541M6YQtNXszlWdiYdN6ZggMEt+k9U8oAs/
WhPlPkU39ilZ2H9NDLX2/d6F8o2eDqLhM/rLyhsXCcyMGrHQE4mFDfA231AqcMSt
WO4pGl/jW1ovuQm45v8SDUP1Mb/QjY9URUWOJYSKjxVvmQY2doVrANltUoT4abug
JrQpckRnJJSD2kOTlU6LLdry6sR1/jzFXQ9RIV/vHju5RGhZbRcs9+GDMKm4N0MR
JJlvw1liP9vT9CjfT/zXRqLwSud84mMQxbkBoo7An7V+ym/Qt39kpne9JjUnHkLu
Zkz/h6p5eUs7EsvNb6UfN8Hyo9wwi9m+f6k8a7eOjWPf9fm7txMmPDrJzILhpzb1
ig/O3wcRc1j2MD0liSw+lgTCwTExTtL3/zfqLmoYvNQc4NULMnyYxdCITYWZpmgU
dCkkwNUxfLp+t6DgSS/htrq1MsNJkcqSGX/s9Xu/xYdbDaiSA+bS0JMJ09Pt59h9
45n8oNxgNipSyji2gN4xJ7UBqx7HXL+Jo9dbYt30I9hE2Fp5bzUBhdLTHWNU3Bix
QWlyHN39QeJx04mvIkOiSA==
`protect END_PROTECTED
