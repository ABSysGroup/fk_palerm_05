`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1G/aRUuR/jzsBVKmS1QzoY6t1zSMpNHlJVvCfo1fCku6LbSWyTA/ef0SBxDAfm+A
4YqaFtyjXP9XlWQl+GWXY8uy5+RcFwytTNYwqrrsQjzukaCZFK9tC7f4CHAPupJ7
nbsPgx9ZDUjA9K75JREKumrVyvmdB7phFD9prUlrln9Rzt8UuApDyYAqLZYY4rht
K9OCTzhbnKggpckBxaFBXRAyIdNdw5cKH4adSBPsOoQC9MBl0hTukZXkCSFbvYhX
D7paxnvi81yrEfuHkoBPO/Gq4mDU9qb8FF1VeqzD3GmCwu0rMRTcPikC3KNZhgru
OGgOVJx1VSiZo3Zq79yKeRelKYrV2J+eDaTHUNUfIwhX9y8BTV4i62BClpGbkZw9
x/0wSPNzIYw00WZ9618gE7QQPyIeOca/kpRUMO3mA0qU/KdeOV+Mvt/lF0iQJEEe
Y/Dg+C66Cud1YIP9d2qXEhUpPvvkahk4DyETWalAe4VGaStqERS/cejX0k6h0KzS
Z2FD4UzD7s2vtNHx8TV8wj7hnOoW8gyRGv0dIcjKz9Byqa8pMb3dKtxHdtb/lbtF
2kAem4EwR2g1pRS/+fb2/98JY9+YWQ7EytEgowvcFBQ=
`protect END_PROTECTED
