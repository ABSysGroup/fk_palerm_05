`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8xYd4eZEz6K1D3ADrdFC30zSQJNx4PlYEnUEj0XyMRoJiZ9PQFjqEWHvu3jIvzNA
wVIiBiqdeyw4+4pD2+fV8xykVFY33F7D9Wr7lOGbb7Zdj+oxAZYmur/N2xvbZ/VL
Ep6MlG7caSumZ2Xy5aJQpu2D+diRWG85yF232Acq7D97z4EH2rwAVzBmknWCWXAe
q0WxA0yY9Jgvi9fG0zhv3NPdsJ+Pjp11pv3sVHwnHSwXALRWLdsmmEby/1OBFIp2
MM+RDlA+dvrXrpAni6/JEqMqh7XIyyuqdr/7ERY7T/Lnw4P7nLy4s1pvr7SgZZ6N
+dqz2kv4t6NwFW2bwXeQ+a1GlblJcIAQ8HYce0+SCVyUsYQe3VeJxxaxzWM2HIfc
`protect END_PROTECTED
