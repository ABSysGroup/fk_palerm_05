`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9KKnpY/E/ovgGgyc34aEKFOMghhGOvi1DCDIX74FZqWKXNGKjF4jMSkvL1EVZAhQ
sh09KV1J/Ei4F15/q0WbinLktTDAlSg6q3gvujI6SJniFkl2ITKtJTb4EbtNJRxy
gFQaNRXK2ZyFe6nvFtHh9m9z0FZ8dmVQRAWCwOktxNl+3GP7aXwZZV15JXwYodfQ
A9H8MXOBwSpYrRrTLqgG/IrU7EkbQ8agtHRUhJMLXsrRHyUMPyvQRt6Xf50rRlrM
OVw3SNKu2vzqVlhgVw6c9LBuOo62eeklC79o7nwaMCIVaL6emAHTIMi3JM982Kwr
+nEKxJfi+NLQF6hoXP+ne6oRgEe3m9hXLh9Mu/JkdvbGjDCuKvzt5NMj2B5Acvn4
0rwYMYznGHKE5GxbF00T4BauL3FbSyZbT85hGkGGLA59dOtdnVQIiBK+oa/RLG/n
Xvy9Q+rOA6CHRh+ViIWQP2KUKxbwxa3GQG+2gR+JTjtckubiU/c+6r9aIy5QPumP
2FthV9a2YcbI1kWmIK5/7rXxFtATOEhqduulvPv9Vs6tv/ULj2bUKFzkZoetGysw
Sd0X4wlH7bpCWa3qHUkp1CBHEhNRevF7IaiRkUG0Mn7klh4q0IiwVfB5omLx805r
vwmaMiA/WBIx7uKIk5ZtABG5wJq6t3MXb6DgSNXDTJAnvcBQKbo7otsuy9xnGd8r
NCsjMEK+vQ6Wm7P8t7NLHbTCrma/ZzQqsYqXbJ4Wru4TnEn9CQmLBw91A1NzgmrJ
9aoGekTerqTU7jgPl/bRhHLnneOMMkt0dXlMPVvmio3uaLTU8oaoLDnKnom5Q4hA
kn2fAKmeDq20GP0w9bLoq5n4hgSBAFO7BgpQNUV6gdcEv8TNQEo3Fb07pXGvrR5l
nGC+8ekzzfRIWmF3M+tVGTzDXIcy+cG/NRcS3asjeNQIzGrnEhyXoOVwvT+eJVbI
x8hpLEEr+Bb3NHFVjAaddjz6Oiw3RXcml5ghccSSzker3cMy+gOhM2pZeW44Ku3s
Ssg9L/gqUuG8HulZXIg658OZgGHI+OVDW8BXCjI88Q/PkBUg2cZ6sbS4/PynesTn
n1DKguuW2zha+O+vUWFnFOYeCtPjnKzMwP5Vbg4CKarjk29HVTJIzs2IaF123stG
O2WTeLkF2wGCZ13F2xhEKNpAXc3QA5kxhP8wsaWXsEGF+6TQs8oonNvoCTMZeVEs
3HrKNcfQF4MDflIdi1jm9t7wsaOds0atg3sjICvZaIaZ7Wk2sY7wRUsfYyIRFk3Q
GOLKqZ4qyxCNJ4pg7z29y0r0liV7CbswkD/ihZmKSiGz+gXeSEg763FvegHGXPGD
3h8uPSTJ/d/ZQiqC8tRWtyMRJeO5PgEDGMAPrTGSi95NsqJ9ns1gyMkgOqWV3Li3
`protect END_PROTECTED
