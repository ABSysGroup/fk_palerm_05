`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TJCMt/6tVMNJKcRDZFg358kdUvQ6TFvl9cByHDrJNw51fg5gnk94O+x8LsartwJc
XOP/0wcYHQql3eW5HKsgPbZG1kKwk8EOoavz7543F/qBJ2Q6UOfHX2riHjZ0awEK
CVHNVz0AJkhQUJ1poonbHulhxxVQFnFHwYSXTupgwZQRpohPNruTYSJoxAUPm7jf
SAcGk2WpnGiT3yH6oX54waApriaGo+KlzxdjxNx1lq28vNLc1INBOP/+EIi6pJ/O
/tMufx4JopwNahDDxWbvG2AUT2yxZ/uQS6VRVT6dfjOErMlfJz9X56iDDL7D7IM4
PUQmBl0EqyWiBe1aZKUq2fvm4Rgdl2QhoCEv5wYYgLzu24KjdoaeqzhR4T5kcTv3
PtnAEt5tPZkxMeSRfgaG6+QgfapFugKAWlmL8aWWpfeM5Lgk26FTZaE1MtuYVc/U
xGut+KviJlaEnt7F+SU1eA==
`protect END_PROTECTED
