`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YzjNL9NkD7nimoBiv2fTIJhA2/o4W6DmM0is8leKCjfBKcWG8bbGiGjvmuBKEVgx
ZZtD6BeF9LkKe7LXC/1iGFv9ZgRvsuTvEUhx32WcMxaF0TknMn8OLvnW/d9+3h9V
tpOCsTnFML5fkDfKXpBLzg74fNdancORcDSgA4+7vtqKbmTcEAwb2mKBv64729OS
27k5xQ5GHQb9t/ClwalKAKKYYuDVaU7IXtYNUDhMi2ZKD0vgmcHH1SJOMgk+b2Hk
sTh7kkrI3uyDnwwAZrqxeMyNA9JuKUSLqRBa8irVOi3QiHNqM0ZDoKdKrGJ0fsny
yiM5kkOLEz1EwfcmAVSS7c3y7haU8+/dg52/bfOygQEviA7PodpGi85N7ewE3SQO
iHLlFU1sa8nJxMIlGNtnbA0j1u1F5cTjANyyEzLBFyV4BCcO+9JzRF8PFMekXQy6
Bgfz1QunSnFCDn4PyvJYvdTKYYRzjWJfzAwmh/UKG2hFKEslXcpXcR1n3sM63ZWo
VaE96dnkv96TMlk8l345vOAgV2L0KdTaEMhU59WHkObWFOG2L4ldgbZMRhNZ6tn3
Mq94VKZFyMVMSWlpHAFx2Kmj2+oDYOY/DR/DxIWqhQp7djus6aIrdKdUJGE0yl04
fbLexqYtRywx5x3EROEXtuFIWyYOJ2gWCLpQ5jize5ehw/FjAeMkmFk7N4fPJwoH
B9Q1/9rqD72ncbdVzYitYYcvVr+a5BWQWkFPJuXONs70WE1/XKw4+qdTSU1xB7WD
1/TgbpaxifBdJxV9pgeXN4MgnjV2Pq5UOx6zNPq0rH85sjid1xp3mj/pUrPUxLkB
8fO6JlJI6u33imAfzwde91dAS2eEbwo62yldDFNFVLi+yQZWsMcmfFtn4YlLqgkn
iHstXwBIrrOehQbJvEF0M89fcdeECdI3EQ2vt4kkr4YaUAPGw/RxGYarWe7ywIVj
5H/Isx/BcnfWaO6i62vHI7BTKi+KxzMTF0FeAEgsW2FyWC/Ab3MBgnDQrG+momHe
1BQb3uchTQSahzjiXwJIzfAT6T2f4eg8ah4skbNbwptIMugiLGFK7C8+FhEnnUob
4JdOA+qV+f83JE4LmmAMRZAZQL5tAoUwiN1zNlCOGuuBbuS9rr4ToOLUaalkatVA
jaNDn8Vad71K22u/o+3vCRTAo81aawAoquTTy0sYx85eFgsGCLhEl1zpYDxh63Xm
FQLtYzYry2c9ZkWr6kRgmgVofcmN4DqOM7+VamEjoocNjL4zlIH7xKorMBY++zpV
CsmXO1bM1LI3nP0XrRboX1nuAhUv7OtbYdnJWKWXDExqXn62Fcb/g0n2CgZ++xfF
3IuzIkf/CSnma02COnTWYCqwwn/lCHpBFkbJKPgtEWkMQWplPBYogSN1/GXd/giy
ksHxM2M2Cfg0MnHCqtqHJuqSt1STOjJfJKY4VD8XXwYekI+74aNmchhF2vEmh/FX
JGzwbGtgcprPkdFxCpw9NgW+l8x2zszREwU8zj9vRNJh6aIAnHJAJepEVwb7f7IE
soXXNZZEaAIxNjwyHKL6isqRkrDZYKrQY1uhKusGEcuFE4g5eTk+rkJUTBDX/+gD
FCiwjNZajAFkSiDdPBqr0mMLSTIJVUhMjUVhm3yqDgzSnLGKe8faKCQhcfABGJoW
Hd/K395Pg2XSkRCT+gC8QnN8fy+peuJofckZEhBQQniqkuyZhOFW+qKJeayJL/X7
sk6WgyW62tlD3x27S4NvdERFT9RWz2lhvkSbit3zvI2YA1oQSruurmi4ObSTgDXZ
i279kgy2flIewZMv/sMdEuOeQ0GrlSxDs5CU0sveF+5cO3ORLUnEEA0gwyq4bPOY
0QbErKAbIhMPlwdbXLyRCtYG09UIWcdZU7f8cGWOxh/FYGiXPV52HOfSxUQrGymV
7iGcIhzXXMHIl8izVxV6+h66N3ox/3NsbfZgmV+NmMp3mGseXhmaoPiS7XdcN1qi
uA0Dt5a1auN6HCK2mfYmzX7yrkRkN4UH3MV5GufH2D3skXgj1Uyo1ebJtxXOr5MD
kDszOJsVO3HMz20KgdGocueiTyr3w7476rorndRealOzU9KqwAAVc4QkKxHugl4m
0bDrV/Q3d3UzitnWo/H86oGyll7myJiDQvuzDn57aQtT1y5U3Io3Azp7K6mjPDD0
ZLE44abNxNvFfXrUaZ2gsBWWeAkXzlFXYjb04kiMWSScKxWYw7qZjP0pLHgTXRgY
2emnbgwL+asgzImo01+438BR1p98ZStm48phocNDi6g1tXfH0CxKjm3bFwFZnctR
WvPFF2LBHuFD7QhDK/U/z6PkEs5/mWgT98/DkpuHkw8gZW+9qcyA//wJnyjWDCrJ
HuC5989Kcb03RT2kzYwYGFHq5l3kDaHiGrRSrZ/aMsW7qcuh1ZGx8yrPlXD48KAs
zrDG/gnKaGeY7YiRh+GGUo8DarKp5/0Wc+7fwE5VumT3/zY+EAK+cCJB7HMD4Q6X
5iXmWsk3c7a51Br41vG3HdRdpU1EimLzqNNstz8zq5FqhPQ7lLaWRIUO7tAm3J8h
yFBUwGauUsH3rYfS/n/zLVTpZlvT6FJqRFeJyltYw77gC95l1RRxays4lRTJsjfY
sC5s5HsixSO76m8Zfpm5cQrr43B0R2506STuGxcquIZc56ABuLfwycFq/5KlcYve
wgdG6al/hidQNahjqsFQhkybUBbQ09h8vJjU5Np+px8UbUxDvWHuGD1K9prNLPPS
haU8sFnpJVLO0+TJuFbRFS/tFDglTlFZXFxHrwpSYW8ETwWbtiEZtrwcAr2t9GjP
Z7ml8cIBqZPHhKhxg6mV47f8r69wNHphP1u+QrvL/pMzjhoC6OPSeEtn5rw0ZDh3
FvF6/bK2s/KQ0x92xKKjyDFVYejGDRssAPogIQvK88//b6/jl0WOkBoVv1Sc7RnN
04pdSrSwlUTiT0BjMQyNGRO9DiL2XdFj0hmQrY0i6PLv5bYGtTnye5CMe7BJP+uv
QMUmEzQDQ03+O/rINTJTHu7mMI39b3wHFveoCOSd9OV9ukOT323cZEHrUXtdwGyl
FHIj9WZMMysQM8XK0KWzHAfyqy2B0BDLnihLZx8AQ2noifoY9hoZOsYtKSQUXqTj
EakS6rTGzTAnQeC18gTTXEcOjjVN3KbuPuJesmc2CqhrC1w7RtJHAdQuGq8YaLCj
E7vCd6TGRNB82f2pRh4kzoaj5P7wdGeXtqc/ep8RXFVwOLYV2YYHnZz0n2ofIqH2
NKc+cxI1+/Wz/A4ObKqNNajsuERMkRf96YL59nvIeBIwbfiBBIhPlnyyJFSoe5Tf
JPpSwMKR8DYFXTbUIz4+UF8dP9uNiNZolLXGmMrWCsBAESCV4kJ4MeXZF9tUAqHm
x4Cao90ScHuxx2QV6+o3UeDQm31Usd1nDgAdf8fkvnFnhru0MzqYWMB9h2WDl6Rd
tgAtjCZQjLrExWKDGGNnw4LW3pgTH8yX6qls227ASjTASR/+qUQipFHV4kUzDwVy
gLHjNmLM7qVyAd/86XVzF5IQjbKCQ9M15decnWv2XizG/89SVqVFHMeWUDtjBaiD
Q7YEGcVx+Z6guHY7jItz0TW1f4vtNV+aWkAy9M4mQ0H4yEJ+3sgZPie6clnFOE+d
erbkKkb1dAXskOMTiovApKBCtCBUraFMV6NeoRhCjXBv6bnwIvzqY63Wh6/vj0V+
EjaGYPkyvel9n40va1w4do/iob2TgReeq9Qz4r8quyP1oo6N/W27acvBlnVtzlvn
Of7bWjxHgqAy8wWxyjwgKsPLTusqQW3XElwyShEgk6l/w5BnweYboP7ZjQvAer2S
326Nwto2hFM8ZbFqAdXwfURxo76m1uN0wOdSJFWRjtfLqWKlqkX+cB+MMeSLYVR3
C26n4e4xCs9uVGaUib1LDsqIAwp1nXPe7NQe5JTSNqzeVFuLwsw1Y8X0MAQHlZCc
dxysoz9Y/g/03ig35hMhnNiXdyZ8+BanqwfuhMpLBGalyboWwtT2k5L+6IlARcVE
JIP0WTdHXsqjvOtTcWVeO4A1KK6aaIuG2k3uTE70rqVmgNaCum3AttEDMWl5V3oa
jjDf+Wvovk+sT90ZpiG0bpRx4vqbMUvewiMxETkmPI3d03zHAcdGBZpEVOdilDFc
Fw2Jo5BDQEqrohSurIj69TZ4OOzSZT0SM3kA/mp6z560t8vPuhCiRv7EoZWmfsNw
D2kM2ShCrLXYUjrS2ha6lHnA+ZhV1GUsHyOLrES2kAw/19vsRMfPPnnAbTxUuQpw
BcAIxbCS8p4aGAOlDMvzNUHA/NhgdofYhraFcsqBCAVXV+qeRA25Uapa2wKMpYYE
HhjQDmN1pFJjZ8Ucgir5zeKY7kEWcCpCczp2iUh2Sj08poQaShcYcugQL4+y5IjM
Bqe+IhWLE9vKKBa9jMTvw/Hesd8FgpP9eYuJChDcFnVhj0VYeI7JNi0g+tClT2DK
MoGlHm6dZomlieU3pdy3QxxyEvmk5bSkglLyykIq0L6SUET29eKKcgVWaoLW+17+
tWSDPigyh/NMEmh4KIiIN/dfl5bv7lz3tDASgYCXGtCzflu3m+htmofhZP5q+AZ+
qgDQQk9WGNgTcozhKm2VrMxVAZ8g5iG6Dp4O4FaJp9qlAwfeXBEIUZY61tSCN8kl
GCyTtVFyhK3Rmr50ffOYlKaHz6JgnlKFT68x6Mi/lKo//sYJRs2Hx9FK+9BFhsj7
A+KviO4s/W5sajlyc6dy3ruB4ZKgT1kP/XwLmzDQI2D7mMe3BDJ4l1dGdEMYpr7J
JnZzArUXbBX0wYnF4qqCNj9SrdaTGFuYTnIYYp0MH44J2WdVLAfeilBD9ITr4ydf
c7KcA84waRNOBBw6lRLvRSqIlnVvP+d1+kM8gfvWnPxCtFVNZooqzIW+RXnGRttr
Ce3kQJdFbVf2tnWHUyRP0gIamxHQ6egWwT0IBalubwI4LEa5Z+oyWGhqbvaoqk4G
YO0WvjANvmSOuRSz4DvKVOBEq1EAwmmZXnVdi+wFf9cpi8Swg/QAyl3Ui+rzcMhg
YZtkV2eDj/vKPZwA/MHLu3GjhYxv76nbUvZ5MHR82VqwH5VKREdHasE+x46vb08N
LibqsVsqWwRe67lY00hhhYToOD0xZlzUrTG8djSzTOE1R5TnbY9ZtR/LPcJvr59r
s5tleOITeQ/z3EThb+au+BE/5tHfzNzZRfGZxUik3CCDsClmCWsxfAJcumYWytWO
WUFXYWIOXxoKUL9EFybKlEL50A11YOY9azLaVvM9PPO/yrq2c0MvMGx5n57HcfI2
AH+HGytMOauCirUZqZXnbg6q78ytNjE4BkD2SbAVwo+ULtXZv1AnNYEv5zS08aSJ
jhndG0s++nnqLHXEgfiSEVpmkpEKloq1or+FQW2BhOY10j7bzXFCmHPIc8Z4Cf1b
F2uTdyuhRgz92xeQqd0i3NNGx/XeGT281zFuo5BlHxHbMZm7CZ9h7yMX+J1LhrXO
Z6Dabp8O/AsJqgSpzcrQZ1tXpStsalnk6z68xPC2bULo08FIqSxoAhB7wQC2AGdX
v3U5nL+IW0Q5EbQmcatkyJnj5eBD6wGD8A6yJFFwE2fP24k2THqBfpD1yURGumKZ
o+ZIMk1WQwsK/fnImIhH7wVqoIc0T0OgsuTfpy0ia/SBxwQvtIuomW7NEa4pYV6O
LSG0sU7IOl5ayJdb0vHljBJFwlfxE/a8zr1ZWtpDuuVuHF2BfWgJMCL41VNx/ger
VAtYR59xB0aiZ1Wf/2TEIr5fU/jA1jgf8WgN6NO9bZGgiucZsW3Qxu/8pCQzFREc
eV1J1Xzxe2JDMnKbu6kkn7KDu4FBKP2aQRA7+PzFsd1tK4yZ2KuzBAy+t/X5BVFM
o0BtnIHHnYbcRWqadXo7VuKjEQsdvYYO3L2HwZbGgp1x2qU2nlUnfvBDsYwwSA/1
LD5b0IBop6Doo2XuXCrFak+8F6fvjabOrWVZeCDQzyJ0wsG15xW+BcDNqliGQKJh
wdMf9mDOfMi5zUJG8qwwkwOsWrSzVaF7bL+9EmUUZIY9b2vF7mf+KJiWb1OG1YNk
b96LTvCTRbi4IGF5+9ay++2O2tGnHpFgqIdx3dyLhUIHTEy0MLE9sLNqoJmiYK+d
3xYemKxMaOVv/oPPoeJH2C3EeQKVCVur0NuGc/CrSYm/aQ9cCqDafy7bsCPzAApL
i9LkXgG/6Ez6lBuDNvj/OC3/wr8cjkWhaeK9H57SDHSxPCrIzAYAnAKaygPrM5gO
jXP+D23PjOfnZTZFA2FzWdfysTLD8yIUZD/uR2rMBlnirDXNklmal84qJR38bJ/j
/06Alfzj5fJYUUhirUMXI8PBzTDW4Z7EUbrMPhyA+maFhAA5Xl2SrfYHnq7zwvRC
WiULIPcGlSOfxFnxFE4G7H7WSiNH+45dWm/XhjRHYakGXT9F3HucEkUjAIJTvzRL
hxtyWPMYtlKtR+64HcZtm+kOW/yeq9bPUJByfp8izIvccGS3CZDjMnxjq5w/QWo0
b3h+EBVq3CkdYb6irogrIjc1d51e4uWROXLAc7gLPCJWdv6YNAWGifKbU0NdopKt
JeO98X2nCxsegmXnFTOFtiqWIOIR6V/PZWRYTIb6VNJ3H8xZAzFff4SyW4z04uKX
FY9TrbPITH1DJLMJSto1tf0eDBNkiX7gYPYBvtBg1nRBNlXWamXPhyUpdIapaMM3
6JopO8RWfk36bjcb7YYC8/7uACAfTKKi3LXrUQcbVi1ijQocgPFHKMcXgnWkJF3K
SPX7Z99Vp/5Ula6FXPniXKpKtcwp5+/G8aoLQRHF1+JLwXd6S5rhrc/pmq1ACOFb
saK2rSAxHKvZOgOgQ+IV6gGH9ggnmTw+bVO1V/tdeWEkW0NFfTZz5GD0evZYqUdt
Ze7oF10qFomWqZQWID6lWjyt6osZm+AuNIB4mveRMUg0KdunLqfyv/hOtDukzfpx
h2feR+hpxBKlr/y8Evg6KXz0GprgNIltFoz6yIVNoOR7uy8Cv8KUDiNysYBlUwvc
W1etZQOLZVmj6aRFyH/wNNtQ6aUFHfgbJUj7KPXi4aXC7QtQC4+1V/70kG44W4TK
+IfJ1zs8XDNTBSSQyg80nnYYQCud/wwGhlynab5IfGZok5/s28WHsR+5nxh3/bc+
J5kQFJyddJ50d+fARumVjpiwdrPoAgSMH+qGgC3qhDP2RxEfqp1x9KVX9wpQSQ3u
tGEqq4br9NBewhIwMQLqoFRPvNI15YKQ+HTzaWKWegP5SGQOUH+JWe1iI4Fj0lkv
tsAKir5D8NKwfurzQ/hSmGXTaylFi7NaTdL9jWLK1zi057RXmF8DqCoLyZMbMMpB
/7s/xfb9nAW804RAhg8xW0oMcoo6seImlwQ7mP2+xKAT6XX2tW65ht+7tb2eqvMk
+VEGXVPoBmlQ6WlMRKy+9HKQbZHMMwweYSTv+hZuzblMnJIGnWDLC7tbCSrs1mHQ
JI7A/K4W79UkB1COHbbEK+Kuja5XcKjS1L08KGsJJdcO7CSOjJ5KAT5Y2MK4NFcg
siJwnV2EGrlWX0yDBw/vKNtfx/OQUIUDKzBi+OVgfIZDFn13xmvcmh3GIm+0xOZF
2gg3+nS51ES8pMZhjcaX6wGXvp01SSHAcvM7TQNKtnWkI1XPgJ2G6/j/U3DFhUHv
epUUAC60mHABm6q/sM4k0VGeGo1XxsvY2nmDgDTV7B0Wtdi2QxVg7vDJ7lTRhpcg
sEZRsNBFt2pevUugTQ1cjCZzLy7rCHFwAXjrS7zzLByg7cwfoM/P1KCz+RihGeSS
KqZMwwAoGUEmhOTmPBrXh0hyoNobK+TClwsO/poM5mYiSNZX1nBkd/p02Uwp8nkt
dPHHYigGDq9htXSYObCitHZLImgPJWyeppdELXPnM9e/R+e3fLbe8SxWCiYUzjMJ
P7qZLY9uMle1SRmnkt8Its89dj5YB6jTmH2HUna0Gs6upTS2LNvhO2LAbVSk5LYX
vYpB2nCwRK0c4APCPSyh+YKgD/CxOlbDctGLpVEOqzasI/859DVQLiecxQoVlOhD
sQ3ThXOt/fH3jh0WEo/oF9x0SGYbPSP4r3jnbstUxBUaghZde7Q7UTotesiB9V28
LcQT6THTlSJb4OhnIe2PKVSTU3UxKR5+oyOzsdvtAGYjWnEthWRIGDVA0D/G/23q
+82FR5ZVdZ/8K9Hkd5xEJsowgDt+u7mQ2lXRfX5bk/jtuUrf1RoVaJ+zw9AWlbYS
Dg0MKr0JytyYbMzzl6wsN7i2/aeiVv8RwP8JH9xomR/ZV9cyv0Dllg7+YkjgGMWE
DBY4zgWV2ojOA6IIM+jskFniZRFISLR7gImxb9WiGWuG4T2x42o/jhTS8xHS/qSt
lxGBiipo+h5GNzPrdUSA4935cpZxGkzqvF2eNllIIpjqze4RO78ntNFxtO989Xgm
eEzMGEmK0nZqbJfzWV67tau2ZAYih9KARrUNxoyVUN01L0iYLEeGziAdb5gXNANR
c5M7iCNZGC5ezb8DoNXV/rQCpN0TnXNfh7/pprId1n4b/a931YxsIFucVPJzR17m
E8oDvp+SBMtRFkMWmzmbHWkXmS/ZDTW71Sr0+Ell/zdiM0tbj55nnq9GKS18EUNu
3k3NtyWlWj9KcY9js1UCJWMylycvkfiGUiZO/S4m+4SwgbixKNSDD+kQjq8MDtGD
GuZzaud8bdmnt5hUpouby57CmQQ/jvYgwHsF24rqlF5uIY5+Yax90u9Yrsp7SBDc
IjxdbdaPQMiBOVkREUeqYjTyvN1IDrcRFuwRnizHCOkpOebajOz84x8FrSnoksC9
cCG8GegQYYmZdL5mA03jExzY1xk0dEO5x2m8J3/eEfnb5nPDzjDqYzmyQfXj+Hq2
PbEjhA34x3QMZLjcoPhASqXJbUZFOgG/kqt3CKJtm5+bEIMoHPkZND600bwQkagf
gm5nSYyS3TZp6i/9WO3WLWJhZ3vDaWzvZYC9JsmUbU1QXX5kqhHtsxDfVZlH+Y8Z
IFrauG6cpvtXu5b/qi3e+UmDLKk2LMwkZyyl3qISfg84BwnCW02eRMl8qITnR8Dy
9/JiYeJSbW82PF1tTNnS04vvT/8INynd5Xz299NGUuWBrt4vilGc13gDhVmPNzLq
lrpRrsLyX7LGXUcMjTRLo3dyweglE5tIGoees13L+CygfhZpHRoDWQp0iIFqJ3VE
N+b8C9T5qPnjKSqT/vvBdAyjmm+iuE15dzq+1KpuvG9UQvttQ8C5P4yVwmrYiitD
gDrOSVUmXEqtGj8i3SBg++03NIW7H1ClYkRfKYyKTZ8/tk17Zr7gMa0CcfRVPaIx
sHDkMoad2LUC7pYyKlIAWHKTPPpcwO7QutDGgvRfMyBH+uLi7RjUehFReCfjXdaw
jRGh1yRNzOZ+IQ6Ibd6m1L/TgPbcQKrX9Rr5ynJz06yBmLhKIr+NcLVHpYNOqUsK
c5mx+bq3EASeAOP7WC0jmD8kL3/9ZO2R8D+5ozrIysNcEFrFW0nAJ5wZ2Tbgt/oT
xPY70E5vsAP5RyfM0fVVHZmC0u2PlfTIS/Akj7BKXTH8EzCfVEW6nqa2wHbF/s7V
3MrSIFj7pT62s7U36XWwogBdYoGApyQtsitHXjWihIGjtxT8l7IQX6ScEoShcNxU
xk4uOmhevppLVQ1NhxMUjDfAon9K1LdeM3Gp+M3bP7NKAWmpJWkNakWEeOjETFSP
/jE89d+xbK114/KP5y+fyUN2m7Nq/d4VP0jNOFq1Hmv3PKXz/6k0SuhzDFS6CUJ/
TF2Q8+e7oXKyGyhSoQF8voQXOo2L1rQSwQwEHnZhmdKX0ENhMSp051GrCoJKrexV
nrHC7YvPnpbYGt3DgjbBt9lwPNrUQHT1xeQdPvzYYuJPZGdaQAguYuJ34SN7p08Q
tdAu1YL8Tw3beGtWCTckPR+RgbTkNsg4tV9NkHEPU6it1iF7H+s9withO0LhEZ6d
80bKys4DxTXSZkgZLkyJ9o/L0vmI2ugJycthr8AKxvweJp11SwJ2lfHfBf35g/oP
qobFJDyfPBn4QbyLGdgTZuykE6IBswxvasPSFfrAwpEdmezq5WOSEeAriXBwANaG
U+Mj6CBD3HHjAKqoXhSx8uVfSDCqsKC6jOm55cwQy6PzsGcchusiEbzSwzTW7Uey
XNbhgHYt2lehJ2DkT8K4h9VkuvRSFOsmPR+6YIQqa/oKE/o87S4QYs4CXVJEs1Zp
UfPyaVZZizdBOUenn6xjO05UU0hywTsak3/dOHPd02uMm8bCdj9iHIiRu7kNXi/x
m+tg0Fves7CWrprP/aLWsLOImViMTFvDH0as/dy6/ruYLWpMha2KVJ3pOX3urH3R
jAOQ9u/9jRRQ7R+rNbkhUNhSdxSFcEr/ZpFhfaDYZ/f96vCnc4njXJBJX10fOych
LJUc+nYZEN6LGE8+UED9pP9psp6Pv+0X+1bMIJ0gQLkvied7q0ukWdPkCJgfNFz/
uIxm+mmhb/Hw/Nq4zHsN4IvyqEd443ipa3g6jGI1/KMI8TAoEiGnpfEixHNCZQsN
5oGcScxWia7fZZi7XOPyOW2f5yGACOe8uU1j/16JEV7O5u4NhOk3SPOVKh+sn2SP
StvpjkUr+YxDDyMh5gzbS+SK2gKxJaqfIhodg81Mao2RzSUFKJ5XPUMUO1PoM/Q+
7WEwIV+YHzvAjE0vVe5DrRA/3Caw5AAMDfs3JSGmOQ9WYaum4ihh/N/nwE2qLtU3
vEAGY2LbPGkZ/kdEGY08zUJ/0I5WQN7g7RR2lnHze7bUhGqmRsC5b6f3zKB4Z7X5
H1nCN5Ojk/WeiksrbbLzUd0ldvsyY8VGPWpzdpRm98golLn7ZturKhqnqFUgEtt3
BSpCvPrsAx7sznr6ptqe3oJ1KTRQN0mvYPULa0bsKHoBhWApjEASTzz+6yzO0nyu
MSBwDGmkzVxrRvXs9NI+1slWIcCtP7Sr9jWp1dNXiXd8nxFteFfjwr777YH1BMyu
gIBAvQ23v6ziYPDQ9+x/DjapN9z8PZ+7CNYR5uQbJUVFgOtuu1/p84u/xdelfDfT
j8K0PCA1IvNL+KrGidAx3NC20/ot3j/x7zDaX0OPuB1wfL+rOeQ6vvOzKAzJKxCM
ZZcAQM7NbXduwv/DXwQbRSGmQ2GG+SHxtz1WKFRBqFr7i8e6cwaXqTF1iCKyYRe1
PE/1Q2PS3S8r5063lnRWe91+mPedeVG+nf6SdX7tYuw4buyDAoFF3KeIGY0f4sF8
dkMgeGBK8f/16e0qk6jEvPOiCbvBTVJ4OishsNvnN1lU+kObDuvy+kS7daLodceW
+T4QOFrKwiZetfAGv0jn/dL6c737z9tH+5BDhJkXYM15We8jzMWGsO3IACt2AjkK
I194Xw04/bqeH4qM5PXvo35wgP/KGxSuzeerD7aexXGmaGTAVstep1+DgPS+EN+s
eofYjXjYzVOM9/xiS233v59MO66WRDmpgIkLuCJThyxbY69jgmFeetwSgJ8+xsnu
Ow0r2tb5MzeIEyXu2CepM4pfjOLmg+y/aJOyJl7DNPhiKcgOKYcpA4tnb+WYU1Vn
/TFL8q3OpsYT5tOgQCB/oozerYIVz6pfKAjZqvzOsFRlpeSXfJIj6QyqjwgydIju
WXizfb9jM19Tbu56N745Oakv7Wd1i5gJIFG81cQXNsdQteIw/vhShwzP2KTMhuvg
n0Kb2g1pkX3IhkduXLYJ06dOtUUnzWCus5YDRUhB64JjQO3UN98kBhgoGPND29Zf
8y7isy+e1Pb01PFTlLmtQhUcf0MkCh2gzzOfm3GT3iw1pj0as8vl5TpF9V2k8mgB
+quY5ctNMihJWHkdpQ05NsECA0xAPp40VCsnVsBZ2Y3ske8nWLnbLx0mbkCRzRH/
9hrQ6FHAjQ0v5uv5KPRQmOtvVqERmXXO5siCYo4s/w/mvYjOibvKbz/v6LyJGRPL
S8WyFRhkt8sYPYLjyskxJ+QtJFbQ22AklDKQKqGF/9hcUw0ThRKW0d26ZfQt1gaS
WQyqIOSYcfVsHE60+b19zXPg+q3EN05P0AtQG+yf7Iv19OGZK8ZiHls62CFv5Y4/
PUzzZlWZyckDiZBtcz2F3Isz9sP23la/5sDrSIEQXjvih6TRHeAHYfpzxB3arYF2
CxjgFjTvQg4+b1eoo0uLd7tv5FDhj9Aiamn2rv0MTN36BYhkXuUO9B0pIF5m/9F4
tTCBs3LiQvNr6FQozY7oFNAcnbR8AK9HG3mUWXqqaSSAVc3DzotIiI+S+lKU4tDY
pGV79+TnbwnUFwZNERJK82Rr6Gfg/atJQsoOSqdTZkZkjipOU8M+2RioJpzSmYKe
ZOKyxxSXl1QqJC6DCpKPqM79rcm0s8tafaJYArw7jeBpdSsgfyFXzMb2EjDAM2SN
1Wt2V+1N4oV9anVvNDZnxACYoYsvYtGZ2770brrFbr9fbVUxU5GMRcKxaGOANHwU
0RMkmstaFoS0qIl5SnQBZXLkN4PJWAI9evzhZqb5c20yMPyKzF464eaWY/j9cdSg
KCG6rPAuUte3TM1twDsLoA/vGkC2pAgklhxp3ntZtR6JkX5S/87zrlVPUepJqLCz
IQ1GIuHnwog5qo/iMijvceTrToKWCKsxvzhASeCPzhcPZJZeLIL6kdKOEMFe3uT3
LiW6dicXnfAn8xaQsQGsvhyQyHr7dX6k4sl9eWLWhwAzCiuOyLUHll/DPqLxZcdv
wY4RKsQIc8SGo7EOeVHop64tGGNc84j6uj/YuQ9qDQzitbO+u2yweO0A0LvUFMF6
vcPIQFUM/NJRzKfnt+Qshe73PLCxbtvOWZ0+l+vy+znwviUrD1Ao4zMYE0URAz0P
QvgLyz5WBfU63KjYyaGB6WFtG/7xpikHoVQYB5MU4kK7FPTXXRzGX51gkKN/mXLc
SmNmKUOYaQHYMmWN+CjuBPvyGggUzYYoxfzzm4zSBGGp6nqqEsD/DZMeWIwyt6m5
LYdXLiuYhI5gOJJtq2mX7Vk+YR7HNMXrB654enS/OuRske+pALjboTJt2AhJyxws
Q9ZH8GFybFJ12DBQ1Ey+/ba5psLtyr/tJfI5rEK9/GW+5Dy+lnh/skeX7ix016On
Rk4FbZk68DZJawA9BYipGMtLMZW63m7bQx1auJP5Q4QqDaLrtKhwS2othZfedYAH
pC9u0VhaeWAlX8cmwB6bUXX5dAA5HnytUUa6G3lEt0mT66DBR4W5zhlajTjnV8XO
r7bWZ+XbAZjusbLvDOshW06NUUS9bIRRCNymZQQnizUzi7GtVqHFfpUbYefOqPfo
eL7YjJQ+Fw8VzfT93hH7XINpWgkOm9LEsOO6WqtUFpLl8kebVCsJDA6c8HidqnQz
bNFnK7wQFEjho6Gq8VlNkov+V1p/912g8zQvFiKnsCoitMZpjR8kygCJRlyCP8Gc
MLQ/6QaiUQBoOEBaKT3CEIuLP1IX5N3DTIGbHqSlRoqKXwm2/uRgWmAiV77RAaoH
9JSaG4K1s88lh8G5INMtRqKHrDes55QbNBsoxwHe4lpx92T3UBZHVcZxwXGfttPR
v2Dq/tLM22mjfeVL6wBI9wVklrYIWZ9Yv4KvlGJQJscdDgFXGJ8CjWF8sWxMap0W
V3qYH9SoZ1aSZ9KWXlQpy/fd0xfTEDbzR01sWyjePvgNR+kC3ok22F7/u6NAjunb
koluoR+dHFKlLXNiFT9VSqxHSZtgyjxNtb44rldd1d2Ly2GTevWHZfqJxJipsO10
c+9cn38zSJyU0+XTQl29LYftowhecPcZDGTMZRAI1KR5uXhJct5s9PDrU60GLoIM
KekGZLn1ZxyCccn1h7WQIJuCGTGs3kI94PzCUBBS6Dg903V9Oe9jLDpfZHgGuGV+
L3V4+EbA6m2tI7LeuvVtozbQXprHd1zJku9NrGdo40tPWaCQHqiRqbNqMpPNQQ0P
WYl1znPYkOqe5urIDj/nR7AuToe2ud4mwVXU7nVeOxOR75nXu3pdQII23EE8EBdT
ZyBTrERRHnMEguBUD54vn53hiM0geaaGE3XD7BgbfWwz1z25ppSVtGCCQrLQoPjW
d0IHMSeZ/JQLZL9aJiQSHvaVIkwujqLPQ5V2zi9rjXCGwZ+fZGq3C+AOgZum/UDO
dEdWhn5/WKGsHI0g5VApEPwPtx9LL35BSwb57D1qJCOWU6X6SmBbxwcjt5hYjbm2
vS26lw1VbeUej4lGwJchCG9qndKEet1MlWqpEIlIxD8C2z+ufRTZ9sMO1lwfvasw
L/38WskwHQ+daOEHUdpbhMwf3oDuWkXhrvrQykjk33M+a/wO2LQrsptzgvAlDrZf
0sdWebrENKsvuEtFzlr9dFmYEfcrhL6IuXg22W/jrAcfWeMLdfrFsMzOmbvRuEsw
HooIkk/WWjGCIO/K1AQhfbqk6kggUxTE3PCSVECKVb3ncCbS4ARD4pULkMdyjiON
gEmpW3FJZMBXCFSP/gUa8leuG7qOHbN6NhCZeGKaihBdNsD7s1DDBtVGTeq3Xys6
XMvbppDSVhtuPTeXhjSB+8lhBfBo5Y63nPdw0TXnECzW6TjJiVJHdfn04NfnyphA
BukteE5ZAT1qI/Gzl+6wDnDr2gQ16pcepjRYWl8yz5Pa8GMXOr8fpZDCk2ZaXDV0
VWaq/LHby+dmZvdXrtLllc7OadoXSnNN3g5xluo0bOlexDXAo8you9SXRnMgLZDb
SWClp5wZBGYm8K9DdXe7aS5GX4qFcwLFBxg2iBimy3+pvbFxlVGiU2mRuiwZeA4X
P1jDRGbLaukO+neL6/3uOg0CKYzdj3augfKcINE29deZelMkLmT5doHxSQtBWtOE
yqMRkrJXPpZQJTMolgNizph8l5ZQUrSc8AHuG8nRdwWUWUo2bRT0Fa6eOrnipl6h
vaYgWJIQTkzxX3NMV+J+dGhFQnLuO5c5vfVSxtLUI159QWhkkmld54KBn5Hkxnor
amqKylHa0vvT70zKuLO+bS9pbFov47DL2Nb989gLW8o2OmhM/ZINVgClPVr/wzgB
vvMXj2Jhzo+77D8bLwdEF5Sl+u4JlP7lUVrmsjwRFXqeMDgzdCvGp4mA71HoKtVn
LbSXbbuUyT+2d+yUiKRMfoD5j6DHTSSSvudYj20SEto59fAJYiNr48ERx9cx2It8
HzSqiSpHYqS5VBekdhcj6ChdBC+7mxVBrdEj6ORc/syMvj7yLrc/VWqs+6DqxrvF
hlwOTVVH8HkTrp6l9FaPwPDxzFQUYwp/FWmSvf+Ky+akNvRdA3rHOWPTUqRDTRSU
inOADO51U89Nv9tLXP50ybfprHXku/B/rJej83ROzw4cn+jT660mqyhyiYROvaYM
uUixbrBlw/CfOUx6KA3FwTMe0KclZaFhf/QtP8rXmZ1VRNFcLkJjF2bowSnJKIDR
FDxOntcX3C1Hgt+AzHKaM2qPjpzAKAGqb7JkfKXNmWUHSrDmKaezLPiqBgL9byH9
UPh4AnRnTfVTUAIZPnVdVvzmsg7lzV08k2BbKANQh06EmwoyQysFTfuIvvHERmQ7
CNiGOykCPJrqdgZIUBzmBT0EZ8FA9QbktebqZ8GhjwgT8Ase3mcZRdvE4XhYhXLS
0kpJiV8fuEwoHolb8O9DuoP/oh+aAoTZm5j0bZOKoRSM4/l7Xf81LvA6AFUPyDc7
T4Zm1GShAAIXGgFVigRgQ6Is47O6ytAS93mXrF9a71TATP2QHIDjYYxy6TLJ9Fa7
ZIjZdm5L67sVcDEStA3H1jE6m3xMFArcEadbABfHgEeS0T46PMca76WGWd3Q+XCT
azY0AIPoOSL/wJaMKLCLzBIR3pHV3K63xz55KJk7qsP58XPTkW6hZ4Ew6zYIY8fQ
DytX8cWKBBoswH43cS7WNWUWQIBb7Bog/JsbytgkxyF01SKDKNQYrq4m1g6E5rcO
sMMdzheoCjJTteGYHrW3HmufTyXLKmVjMfq5xdN+xdCCidkxhdHX0qcbZopu94L3
9+UP4oodUBORJV/+lkL2UKeJ7xkqEFj3u++DGZUh6ref3xp4/sHETzMIBrIvi1/H
T/4qbokx1xJ1xv1eQyju+568L88nVG9KKdGq5tKf/GcWZzGn5YEVbSn8Iw97n4FZ
oftufRtIteG5flT5+uHgAGIgvl3Pak0R9QJlwcxCnqzaoIGExVbDWOTCQwljXpx8
IGF8tpaaIF+QqUm7N003RvmNj+AZyRyZVLxqQjVAnagRPf/hSZUAPnTF096J98UF
1LCbtA11jvxUbxruxMPp+5uV5QR0k20YrZ2UM6qHzo30m60qACBEjpqnjQUv16Pa
g33NL3r/itrBeB+rol/2lwIRSmTxcjgJTVlolJFP73l0jgWjOe3NYksIOvhSWomf
1YDsxjsQznxE0HO0gkXkO4p8oqj5rKaSJDuX3PHspuU8LNg66RbPUUsroXqstcBe
osP+pxxN6qmVdhDNZcE4CX/9a9MQvChaHnBNT70in5B0Q4cA15g1uzm6bPaQRcPz
fcZfWSzhaDrds6VFMK/Ex2yrVAhrR211gj+ZU23ETfgyshBUG/J9HrKj41SLj3tE
cHBYmq9Bi42MxF0rdrqDYPUOPA6RnGIgACVn3xkohKZU7RzyNmorU7X7ZJwe9OxZ
eqM68YrbDfhtFQ3zC5a0MXSUcod5Nnn/qnTepRe1YwG+i14lyiAIv8YP9ufoZ2VJ
VVsjrzL0iNNBqPtIgZayo7/tOqi+YsE6+BZjPkFfpsOq8ZHsf3hZ1JJXCSnjuWYA
NMbKNDUL8eBQ2V7N+MkuS3xeo+QYqqwi9gI7Jz9eAgRJD7JApTqfO3E7Jw0eMjyM
ezBBw+UEIy5m+R7EVpfCaEzRisZ4i3lf1PuI17OQ8+1K+YlWpK8Iuu5Gp8eK8s2X
XHqoKIvySGQTz/uAN4OVCpcJ5oIvsAd7PJvstbuZNEhHFL14ZnG0v6q+GKDui4xo
YRARDM/Q4XahQ/y14ioGTw/BsmfPOfLKL+jX9mH8C0X6w+ALnhZupXzRscM4RSeY
FgFq6TYlLaMiRqUYOA6TRdbIPit/k2wXk0XRGdMYGhfHlzfrkTc5QZbuvTmNXaSl
UNRqGFOY3//PmyRwqRGri4i3amAt43IcX6aAUg7Q+b/yYkXZr6Ij+cFTTtD037Hf
umHNm/ucOK3D2zqNwC6LJW9Dl+pCsnwE47TVi+HTuF1uTfsGs7A6PfjtjS/jiRIB
KMpzUBRQcX8aS1BJdcyKGUWP42fPTFE1CS2NOvzCZzRDVjD/jbvwez6z8gJvb9Jj
otQKXvHkt//tAMjnYv8B1QsNbxBEd+NtjPWrKsICsnYPunwiJtrAUeZLi7KneHxf
hqirGSMz/ODm8sRlKr+dRBErBYF1QjygOLxpf762s8F3BJ3F148H+ZN5cpDK/T2q
AG56XRQK8AxuLWd3TpfLhtWQjjjKmPlSg9Hz64Al0EpMmG27ZKzum4EUUdmRWHRZ
o5UQWC+LBNvT8R/5dUow/By3OQkrMeStDPAT95gmEdhT4R3CExnciX607mBMG/gz
3Gz/IbPtvsITe7hWfegVWlwa/Jk1AzpC1oPEIbVITnhayfNnFrCtBU7ft8RO+4P5
FbmQzb6ilYhYJOMnUiDQH95VXesvTSanPIEyN5aFFUD75HxWB22j58pqWwwFmVka
KFb7K/yd2WkYNvOLpdppbu7ILVg2u2XHAlUSjx1pBVSgCkzVJPdv5k+C4ExUmkL+
lQXfu8i9Hc2znDjOo2CO0fI9DWENxznBi4BPnyt1YyCczO/ah3O/TAX5R5lzOgPn
gOL57uIHemTFGMaxe3Bc2+v39QSuxAmBfabCE6ACFHKeROXluiBKm7vwwfSvjns+
ZexglT5o5nSCTwq/f5p1vV48DCU3SSikQhvmCAXGk6A6MZVd/i6B2/iMklufsVNQ
he/B1LRf8mlCn5nDcIzZOtW+BGPMpImb/Xs2oSsuBruS6IUXAMp5tEJVwlNm1BTo
dCxlGlXJYNQ2H+ljVimleDlE8r3LLKn8umG47N7zjM0XMo34YQnkGHD8yFyM/JgM
mBIlS6eoJHYzLMoOe/JATZJW7LJ6aTzcB5kYR8N3BB38sZbM1+V7FA5pnOlxSEWT
gAlIQSd7NoNHKo6W1nCgQK5t3cXZQEeu5U9XySX7RL5JwuV7ZZWVXG71d2ZQxqs/
ml/ru8tKKy6ZrEGh3bnEQovDAyLGdWkNseDcomm7KkK45Ke4BRlTYioIty3biVIL
Z5wGLe/6VFveQwernBGR6JqPKEqchK3Uj8J6Wk6/EV97GC6lz0FIrxEMoNErJbOM
KJXSXTbzk/rQr9OaQ5iD8Q/4rVvgFcJKrWfDqrccmTHWj60UkWvswI6KT8fOZbRX
WlRa7CYxexKbJ6cIiOOj894RaM6cKZRhNOXBRQYgfY0Q+EKqwI9rn1thDp+zPDEw
vX5LdAvWmBy7M/fDE0gkwOmtUUFUNF0SHpXcEVs0hY6VJbwPlfaPE20eqfBCWE0V
+rJ8v6EZYKpYftDuJc1VMKHzu2N5mBlq3b7+KFKVIDQLF9K92zaMLtoiwqhQoo7W
API8q76YYXd3EPL3v/g1a38u+1ArnyA+ApxO2/EnbxpdSEoP/CcpKLgoS993jDF4
GuKEbE7OGxNMpsJlsh/OqCS10aD6/SZn5FqCGnL0lrwN3Y5EILiASgKn1l5Hr36l
mvXxVhrJDhKkUAbLxYN9wBK+soFIsLgYLcKXP/6xRjN41M/RG54EaHrboYMvRtJB
DsdlPqIX2jBdjbB+1GGZUV/la8yMWKXH+iXcOMXb4SmOYyI9JYUNh6g+D6iX+V5w
om7iPFIKWOPu1i4xUKUIB5NsCQKCHeuDYuo4W2fwz5NlTU8EGTNKKX4PlSPpUcDe
sykP2LAyvhxj0GLGTqMWBg7LfFKmlw6DJVY50UQIgh3U+qsao/c712//7xKGYHGY
d2B+0dhSRFRMeUgqQ8igPk0YXlt+obzaJ+ltWbTjJqiZmrioTVM4WatNXVmc2uzr
RBwrF9ljis8MmEinQVJhvlXozXrAd0g1GZ3r6wW5G9BZnse02zsLIC0cefghawlH
cAZjVD8C8FibynVqgeavyom+sQQoVhowZrq77+f4ftD80YEI375kOTbyfdq+Dz3n
W3Uw4erREg9laJusQ6kWIz81pyu9bn5lKg/QAdD/NYlvPwlI5wFP2iyRkgU3Pv7i
kYn/l4iKu3IofXwU5NauKAM/MMcyiVz4pARBZieNRcn8krEqqXoYbSdA3t2ofRgj
pOZp/77ok6EDANX8L2904QNzrCPnMAs4vEDU9x2fwWytOEbEAzktqvmkPWQ5iKNx
hDaClf7tKuyF+bbjabB9z/FFkz1FaXSf2hxrnCc8DYHmL4NMEt78uDA0P6oA5d9Q
+UmfIoBLWcCY3shpkZCJcxJEBHPNpw6dJzJwEKwfRR0HEMiTu34WjHDMuD38ADza
+ukVzMnsG11bAGupoFarZrYcKPF/ePiIMiBvkWn/PvmCRKeDezwFy0V3I9ga1ZMw
7RU9FqA7OvtMjr51lvSvAu7RiZMl1QMNgcQlXvWrdkcwQU3qkyiaB+7I/X0z006n
2r7KJJa2ccJkSHpcCBJs76lusmwXGw6A8+xyb1jcD5C85FvABZQaY6L/7vf2Kx6X
xb5zdP32jXqb/iDi2W6i1q9SZDSnyKV+OuQsM0FswgvR9VVpIUM90EFbApXas9AD
uYoEA22AWJE3LQ6/uDiGiUA+lBb2KtBYkJUoPM9NQp+Kcz9v3FCnIMQkIezXpnjq
T4KLK/puJnwY9qFDKqXWG2CBXGS8fEpvoLy0ypLoRtLKj5UmzhDVlpa/Trp9AdSM
Ulogj1ZUxU6PDie5QrfMpcaa1wIULMGVW3SbLwwzv07jG1t7TInWajP7WyqA6ZhH
2FdRFkuVFkbZPX1S2bN0h+mm/gy/t/9GNlN/V8ZDJ/vMl+ba7XqC6MzEmvNFVxEM
KuVIZ514ojOD5ToCY+spQ8Y9/3+rZ5+9r/L/qDnRslS8KOgjQsrn0P8ZV7qBaVyo
hyU/g7MnRbCovP0nfAbzZKArJgf6W2nXm+UKcgeE89bK7I2sAEdk1DRjmoppEKro
zkXisqqntnbac4QoRveIZHFymTmpZDdzVJshw4mKlOaT837v/cIq2JiDBWku7C/I
cqwG9y7v43rNVFIRmADWHEO+IojJ8WcdSLl8VluHlLj8uWVE7IrikIWcJJRyzoFU
+ofJpKLeg6QJiB9ewG7fIKNk5I7ZJRgryyLgRfdNg5jaaLmAgs9cKhBV/T4Sdb+C
fflNYKn/l8Kl+h1s7E5Id2GT62iq4ojC9Rk2DwlAdMb+fGsEw5FROz1LVxrjeamj
gJQVzon/Io0SXH63BrW6oPH2s51yQHnRQqdL9QvLNHrjwTUgLK/3ljKY9TveSdSB
yUJi05gix74iHdcViLqtezXrps3BrEz1CKY6x8x/8uj3SId1WcaZSM/Vp1ZIIuCk
Z3TRLFHZ1c+QmHv32V1DcjVilvq/+TQdEz4I3ZwA55pifd4ote/ZDyApjHbR99a1
wDw5RRY2/SQ9udm230ICTcvk4eLd3a1ijo/vyP/09YpjvF61C+Nt5fRETGvVS7yY
ihT9g6F4tetKniqrTuA1fAUYxdMeQ25dBnH/p6aOeXrwI7buimXVkr/aht8rFNsR
1FRuDruV+owhiH1y5KOo6TKg02OiWI7ATpcXq7NgZ1I5zNtOXVZn+2hpBaXC+dVo
Mah3RO81IGvvR1Hw77VbdOOTmRuBtNBAJxz7eu/K36XD6ITP6uvahebUhh7Vg+l0
MmrRD4R4NoEJdAyDd5oaJsZIBorgy4JWLHX10QwhQ47oJDn9Rm+ql9LM+CfT5kTK
rKCyfcAN7uHEe3abKrNnbsh5fzdRNHJKjfiHxOCb6CLqYY3MyBxt4C0s7vHRvZMR
MLiIjbikuc6ORALSGQMYJL82aOvZyC4fapcvQ9qchR5slydNsePjaWjNpeNe7eiO
0QyyrjAx0LcfyrY89wKlVqlx7k6zsDAwtNLPknt8K1YtMLyfOKBGapxUv4f1MwlJ
8uEfXRGiOHedWikJziyovroP3frc3vhagIOSEoE+Is+f/5L3cE+dzvmmLXJ/911l
WzUuooy0Kz9JG7FrnYOcaIRRUqT+EnpYOiUOfq3K5mz7/zpQnvbFislwq1Y0ZCvc
I0BW8ZgO/hOMePvXbCE7AH4DrOn2pnQNjd4eXnpDfb+s4GgfKjuMkLcMcgsn2ejn
28c2MtGhAWVTCxqId8FX8pGBqQDAQq01vstlWB2teMNdUKyfPwVzfP1s6LogqG2K
Od0uXNd9noBeK4KxWELjXbpkGjoGWcoYK+GeBvLTVuthgMmwK1+28nwhavq2PTEy
kvPXeD5llQZwgQn+r7rrbR91cig0z8sCOH41f0ByV1n7pki1gpB8tq9LnkJzkip/
v+fDOumYXzPURM0aX7iQWhWr9dyD5eEY2+lLIY/5K/NEMNorTpZKLDBLbFFb70Fg
al+CI3fksgoziWY6psDAvBrG8fEk4jTYf9CHi/stkR7pAoIGiy0FTNyBoa0LVeu0
tbV+e/Iu+EwrEoHXAdTB62di49+XDDriH6HRnyiBu0UnwX59WMSUzWzl61TgCXkB
bxHMDtVJguM/YIVBx+C58BxwliZCwIhhdhER90F1woAEmRRijjz25CdaquDsH5dJ
5Cxi9+TqxweBR+PyctrAdbQ8lyzKMFJHVRmy3egrjy9bDVKgd0fRF08NFUJwrhNf
UruYtcR7AA9Gvd00hru0hDu/GeVOn60k0qACb1hpOLwU1DsNvJjYmygvVzPpXXCn
DP8RT2h3mP1Oto93CB+vuwN2Za3+H0SJe7Se9UW35AbTVvL5p9h2S7w4Zq5P+SuK
HlpD+AJuOKfpcojwiYkbgb4i/e+CzKKLmzUWJeBPYUtaVE+sdkxS2uX3NuwwuOuK
T+zGiE0UQufnOjCiF1DnhlRExLGmFXWfV7ufHw0mxXOJI8HNvv+ynmjtVCfefL9X
M2ARi57qSCh5pFZim+xPiPhICiWa2QfaVk+bJC/7uDOQaLNQB8uthu3vzRP0S3DH
uDFQwvKSuSZ2g/mKGWGailrQr4E/YLyTiNHyHHDyxoMpSchHvyPStZ9ZBlIx2oCk
22UjJtAzo7AUJRQPDnMFtkfVM8KERrzsh+85VibTgySZnPjQf60j9XXyWK2dR6Ur
ZOZpJ9jOfJqzRKu8H7cNSB2XhV13wJ+v2NT3XqKQCJ5GWeXzAk+HgV9Coxj+79gE
3UtnVuBi4C5SjpHUj4FvYsROT0lum0K+9Ow1P53AxUkPG57nUOBGF3s3NobCltG0
eUManV/qMPUm35BzAMQS3q/Sh9qyqm0MP7jj79uoq53zT2GGhvUZgSCyfzcR4Gbf
v9VTTAZi5HTqeNT3I1K1FHOlO74lSKWvGf4wIcQf7M8Op40t77NY6dLN2IzyL0C9
3791BZWflR0DUkDklEh3puBWyazVWCgdaj1LwZ7w/396TO81RwaSRSKQh3BFGMWG
+Ke8vM+/1KlExWtkVVkq3M+QycpkNQbLPjGMilOdiGFNtTlW+2izfBJcUtRfezbF
RqU2Vz2TL90g7gYSkAYKETcSfx/yLFU9rfIhjSXjroVsvm0zbUksa13fiFT5hRC1
EV+XcL5Plx19QssG4lh+nCIePVrKUYPoyv2XiRVkSBok5jsev+WJXYEWTYwCtGSl
RZOSSDoFb8Qz6F6nNLaznqEXTYToBWkCh8S/jnk1rw/wQ3aGsUGF9lqjga3F+wKR
yw4ji5kMXWhI7S57VXdG+qWwOkaFcjq198kTB9XkSMJXq2KLu0SVWg2JGqmsR5cS
zuSY9cAY7Oc2PmNPRXnY7NFXpli3mtGi6lB1NIku3ckr3fmn5+VCbokO0lZgZ7QK
SrsVzrKbTbQRiNdv8E7cgMo9R3/gc1mAZ6PPY3yPXrn56GlV5BNhevek4U9frVwV
QOAx2WrGuKrwMlyUFfJw8q1LaNVbMtKtEv9zAvoVn1UYKs8wHUrv8E+vRnqJomLa
h4CNWuGuNH+FQIe5QckwOfZ420j2cFszbf1TDOiCWz+6fU/VWG5eX43id+g97yPO
8MGfNnjLmTvLhKc8bDDaEpxixc+4OugHs414rhmqSux9pTxH40Ydryx+MDo/SDzs
zASxYw5XbVAavGGBcYCXgGAWhbXwPEFRKNVKyBt4bxpPx98wuvV6Ekm8elm2ce8r
uFX1Pez3GqPdVrUALiL4a7HPB85kWixTY+OVodu9AAVRkGIq0bE1cFRwy+8xVU5W
itKHibjvc1HydXoopeURbhQPhcDAGUnNOWFXLnMuTVBbhtGwGklYGjZmLo6xIhFG
0ISOOuWEEDqfzJSftWL59JTOLEHC4fYkhFPb8kUMdkcCTeDPAL1pu7b11jtPCBRN
58nXWOoq+zc8rUcyDMeYzQZfIDvbq3knNMNvRd2qKvPIyWfPmPBRD7lsU8AMz5NC
siMl1tIVftyQ0zo4nCWjDWQyPdfrwAcD8a/+FKllpCrJ0MpjCX4bUqtmmtj3gXyO
oPZ75+ZsUgK2r+DZCJZKPxv435aH3co7qu9KGWBKg0r+VGfmQf5rak3GTIfiBTLW
tzKlWLZoGjyqur6w+jtSsN9b0MWQHrW8r8Dz3P5cnobHokXCd8RMn6MSrLjFcCmo
jdGb4iBn36tuOGPy1ZlEyUCM4s/jNdCc7BGKSBbnmBf6HLO5wLjG4PX1Ciz2XZ0k
LaOg3NW+4cyZnRWI4WSnea/IC2clxcobHZdFORLxvMnir1BkjgRA04YS9mZBgaXd
NBOLVLGD1Q5MMrzRE1FLaGSL8qLsI7djXBfPuXn3DkB4FFZSlnQXqcblyX1319i5
FOGmWOt2TDMXV1j21B3OSakPxH396k5CsO0OQ/hEeJAE9pkOJFnUseoMfkCjqfT/
6xe+4kIN1o9zKS66cYZXotVvaylQjw3pfBMRnkaDO8VR0cNI8buMRlUB/g8WcRI2
tziBlH7isrVfb/g6oRhTR7sGzqTs3sLLzMlPKABPUTW8op/PRjeAfjegXpN+76Wg
NmTKSOKizIgZJoGWU+rC6i2YaDgtwGHIlmf0HZik2nRmCYs7dkL/wyIrkpoQe9gY
Y3ByD/bobzX5EPokFDGYWeMDmz6tn2Rp0/NvA/I3nZpcSjntEvIlvpD5fYLfBf+k
gI4uYh4cqSGqvZ9N9DpHBglIkm0qAZ/GCzoLe5dL5sYV3bASgGLGtgOlZ62znxHx
vLixq7nB0Hv1fVCgJUDxpk2fwfDyKk9ySIybG850sqllHkYR736HoGPP4HHgqWi1
UBfXDDVGVOdztZ98CboQ9aroAv0IRIazzrBfFTmVlJf88OzvUocJGjI+qkl68MnG
cZtLjIlNBs6SkSqcNmbt4dDK7J6vkmKr11S+XI7gPcv5nt5SDCI/yktNTi2J64lp
iGUyZTiz0YZoRNS/ByWGUxyRHMb9f/te9NRqQ8gt02v+3HorZzwyrFKjcbcWrBED
Q+P0xvmsYj8euHueAqWhkbRm++wE5Iejx3ZoblmX3WFFLyHcVXNaKt9adgZEziQv
45NINNnQhNLqBvezZ0sZpZH1SWB2VvXVtCDnisgLzBGQy1ywGb1gFPc9v7sLofoa
KT+oSmKmvWI1F6/d+F23JKPibryKePrTnAOlQ4hpodgJiX5aIpdiKp/PKJlyMdjt
A9Yi5Opz4SpIc1X5+sShAy1OZoM46muU74nn1L+0Qbn2rxiaOhHZ4w9KCb+1c9FV
E6e/1pIg8EoCgAHa/4Ia1Pra+uBDCH2TkWlA5PvAnOgZtycgXbG49a+HJyePR79z
W03nmj5yeZBpIHh1JC9D3GPb/kczrr61SYR8dr5oQfgTgMaVEBM8FLHIy4KPpvEg
MRHrz9ySU8VInZ8K4jUCo94FMWbui5xqQnHZFWBMecPfyjDdhH4MRzfibLikVCUW
5qgcGWtV5a80/M5lsFuOO/nLN+cc8IxCyP2v5Yp2+gfuMTy9/HHfVbvRu479N+jh
3N66ep1nOXsl6vJMeiEZNWs6xsOspcxgwC9cJveohX2UR3Vp+C4wD0j8F7zSbFoc
juUkcImqO5KUdWK0q8cSjt1TB2DxvkoX/rPAysyk9SNSYvKeiA9MgloAt+ENELp+
/iI3iKGittzYrQ4ys2YZN4xGQyYRPLm+0k4gzjX6bLW+jRxYX2QEHqqHpcqcgEUf
ot7iA8T0PS4YGuSFtdWbSp84K/maVLBBXp429SGdAWupsE8DLK3gKguPoy6JFFDe
NmH2LuJ/nVoQeD/MA2gxO2wNYHbUbKCW+I7vQOChWeI9idH9ghwKBBGg/dXj3upH
GBO6YjHbYeDfM+WYIK5v76rKD1afoPQlamvAQgVd22gTue0/DDnL5cxPX8Zvm6Bq
7/JjPpJLf/LXfuB8LVYc22sj4JbOGHBvpCRdhoTdS6o5fdPVfuG0vPGQhoi0h33k
2F0FmALzBCn1MYY9Ynqi0lD8IiUDZj1fqBulXLn1J+WISOb5xIc/QfcIjeTgh8jl
ieNAQ4Pn7hlRGAmWMJ7UelD7cJZiWolf9AhtlL4tm/0y4E4solGtW7QP09OwEWNb
7ROjkxiWpWF5K5pfu1uXjHNBlv/Mfa7A1pSh8w5wlCvujiv73qSEFX8EmHarTjiz
7Ls4uIP+GS8kx8N6QvwXR2RBaowfuF0M2ymne7vKtdNvrjZHBG0ENnwIlnE+QJmC
bOiU8D5Bys5cwh8cxT4UkkNqb9oa5PSZIfaB0hKvk8r8XfKestM9MLNI+wZaqGq0
Jkp+bsd3ThluXrCsV15Lk4qWwH/DzHG8YLFYvDK4Grp8KFnVgBHPCicxjEjA9u86
ucBqK9VGnq4VhHD0yJE8tTrr1VmJkBc27N9WkH4kldHFa09R/TKEnr6e/CoTcZE0
YgShfNO6n9C93+Yy9Dsbo9gC6eV7ApXlw4Wd0TFcXFLrOaJVLpUK1vjR4EbH6PlO
e1KAqdT6v1/MfC3nFF/ZG9iKTuf8YMNvIorErohyUqQ1BIXvbmzDJn3oi4LHS+Pj
userVdfOk+27xVZwEE/A1WDSyQ/fkfgo/5rpIRypv2DIXIFDrFjmVErmCvk1DzyK
AaqDSZhTX+1T4wD2F/+Lrr/VHbudSHcLF7djYcETqdRDfFyhEH642BJoLUGkT2XR
vin/JFGGaHY2KxyHslJax0zxYD3YT8FLzzoH7jgXoZ6a/prCuRFYWFVV9V8r5cdp
uUCflC/Xj2+pCgzv+V8gqG9rTY+LjLvjpTomc5mzv3lMWoGyQQxYqercP/KioRbI
q/IagDUCA3GJfMHK2BD8XWn09oiKCTp+H4J2hEckFLMJSHpYAxiKNHkfxq7mHD16
E/6d+QQQGE41uPvDJnxGm05xf3uHa5HazxSe7ooEXsMzNCsf6boIenJVaqyN6+qk
81VV0gZqBVwQNH/qME+dKnEiNj3e/sU6UD22E3tn1M58J0S4XyS9TNq3kWg9qT+K
VBmfO1d13L5BpPR/TQCkJ0rh/9WEMXH5ki//OSDZHXUdIL+/uu5P1YI0Uur4XlyD
zI6ErYvqOXDsj9VvCpMprRo+UM9f2U0nzxRdfwulyUaOAmxHF0BJfYwei3LiXsNH
4tIlGZELk7WPsMERiOzfXfW6Lm4CZXvF0s92lY2MQA8SQsvLMG4nl4bzBVGxfuOb
OVA9j2lawYFESnFfwpHfj+2vd+9PBz7BfiBVKYQ3RIDYDzO02JSuaLj1+k+V6DP0
FO9Jl8hZZVz0+p+zCHaNAM1UVahc39KWyOd5q2hRg9oU/TqJn22B5wXranFt8scZ
pptHvf+OHVRf0bqe7pAaYZ0tbR2ORRCRfPS7cejJLAeC8j3/60xLxlUcFp6iwMLK
F+ZmxEj/wyVLEGgJEfra7ij6jWqYKBN6cLs+anDBGaYBYy8bwkOgupOHLGEmhXVI
t9r5/Noinyl6YQ+cUqr72wdd1TCdKk7IUPl63wXd7p3Dn4cJf5w4RLf6aPVsTSRM
toTyes52tkVSM+x/kJrkcokfYHLd2usBwp7gfAHD6ALeqeOX0xbFKHPEG6ePNz+j
myu8+wJyM2JXfL9qMs5s9Ma/60i67ai6UYpfHE05p6dytbYmsb30NhdkrBs8r2v/
iBSthIZagPVHG1xpFH4XimUl2p/NKVoU3KgJmIVj9oL2Q8eUMy0SUkzkoTdu5PZL
sneta2mLGj7ZKJ0FjixFnFa/llK4MnakXK3NHMUQXffCc5z2zzWSdgE8kPHl7cXk
p43Zsn65TL1N3CunwMg5G/i30cMNqOD+PTDuwsAVQDCkcYjazfH/UOtP6XyL0Tef
8wmkHKPC1OLtmGjBqzuHm1j8DDxV1DavFUPT+zsqJ1vQN6ZAgX649lCcPw1ffU8z
OejqMfVNfBNSF5hy8ixZZnFGBLDvSjlQ+lTmYi5wCTeVZvg6FShshvbwNOxik0mA
IkbHx7XXOQTvaD5IpwiT1QQ9rG7eWVCtsX2OyxbqtlmHzKVshMJcszkGh7CxE19k
eepcHHpL2flm7XvXyUsZb/8OuKktTvf9jaG7iK9BbltWGb9/OPw4fulAT3Jdof0F
w/F5oMSyBF5wPaxREF1swJ/E7aNo305eUMWFSrK76YyIB76gw/tY7mMo2hFdD1ov
rqNUc63/S1HZ7sOMDCpsfRDWREPJWUEEDxOdJcHRcty3R+sjE+2HZTuCZwWzAcZT
dVFFeV1BqjiMWq5oyccuaOQy2EWbSV76LdNMjRGwfbTbjlovGlKR6YXZ4rUA0FzP
AHQJwG3VS3PM1dTSCuMTWBmVJwJzUBW5GSC10WfX1ql8iNw9/BpD0F5o5+zSzyXc
peJJntMZMJQfkKv+UyeRLaQdm7UBCquUvuvPOb6GTj9I532S16mx5yWYYzpciabF
DcoIm77pQCCGXn7MmUJZJzUGRhJkt2A+iRp9RAxSSTPArtwx3gO2hMviHmLuJfF9
2qfTzZSiVbcxZVIR7WFvfQVhVTrTEmWgko6/jfOuTrxyD9aBIx2g2JpnrjKyF68/
N0dsUDHnrtzTur8FvSvYnIIWsCpMkIPLrtWXkaEnAP+F8Q7jXNBselihiaKujHFt
X9ViT/87kRwYhd7jK7iAhxbLrhu8/RtJJJnLqaOVKQKEyJsCVkEgO+TRjBC5ZStd
YrmVmaga3m/NDCiaAIHDt+aEwetHbc0dfEzSD14ld6wzNHQqxOcD6ZN0NDcpt/ja
Or8RiBkVSqUgb4aDlmejZNPHCJG9V5yNzUnxi0WnUFwJjYl3fEkxwzU9xY2Clndo
sSSVj677V/K6DMW0qprS6qxHgQcptyDPFvWWYSBviL8tf/0BE9S6RyDy9oPSiB8e
zjVg948Mn1SPGqqC7WPwrpfxd0WLsjNEer1jDMJOiV1vZit2ZxiSexw0MmBkgDvp
xFjxiccrg0YJnnGVp9pY9Cj/XkIjnqTo4n84VEbVMhYALoTcdBmGB/zOWWr/Vmsf
rmeGl4ez3uEtm3H8Th8NSAWe/zZVTDK/mHaBUUkMjPHNNEpsQVOPsbWPBrXQY8hF
agKUr90sySqZv+vXl8k1ZuNMaMYCefcDaR23IKEGNWixeb5hIpUxBKd8SF2s/fZM
06zwLgem6HLr7Cxj8bzGRipr/o3blbe8Axyar75oV93Ka/UmNUHIfiDZW6K9WdB7
Dblo7+JvDqDT04e3HObv7H4EJxEA75drtyP4R1TPRMO0K7Gu6FVbmT7/c03B2ekl
EzpTxq1I4jRYHVcBhdjcGxPfOYfKcBqX3CepexvTBYTQj5nvfrTCwiTLguhauPbT
7v5F0OEm4weDhttmi7NnDv3JNmpqVq8jhsDa3EVqwlcw8+33jGZWckEID9Dq4dNf
UhTUA0/mwoX32SCthOXYH4nGEpBmuLvxcPqWyrXrVt/A3Z+UWN6kYz3dLV0+kMMK
2NsWyg/Cd0q226Km++EmLRbXYhnXXKgBNGLJ+HmGN2EVUxkpxtF34PHASyf6zaaz
yqIw47p0gNo50kH/eMHnStTWvtwHK5/gaxcaVe/4ij+zQ7P9c4K3GJHhHstMyPYg
R/eGN79+uNDmw2tp9ZtTrXOTNm3PfgIKFehPj3EWeit7cFLJiYuw3uzQFW75/Zeb
LCy3UOmW4chk2LV69RwLB+G1FPluimfNMlB56h1+8OcfqzSpn2iVLFvMPMxpQku7
dfMIX6PV9jZDMdrjV3Rbudjn0Pfz18MHrKffVlYBprrWbGfdjkMUxEEjCoe5sITm
cEx1yyXVQY8foNEXfGVmcwpKU4lG+MsKKo4qiYgGFCi2E5nFdQSbeF1I8E0kL0OI
JwpeHwtpNNP6dhaVlzPRw0uQ80lWlHJUpVTy09g9PcqzUqYXOwsGkUgbcjRY9X+U
Sz4C6lQiSu6SyIyNMuhb77A+HKb3JOg7BxchxzBzmU/ShIsuY7zqG/+KKVhh2u+d
i3c3bDSzYHlDiMTEoQ0RzhJlDleGe6XDl2Qzx3PjYhVS9wGuiTrzANwpkvuHk8wx
prY8o9b0P6x7/zmpQ9haAEh0uxjKh4kDJUwiKVTNIFe4O+vgytCq9SJbZmwSxyKb
UfPRLev1wa2kxYc5VYm5RGigx4xHhpJHPsMmgOkbkD/CpVS09AqsIO4IJxD1DVZt
ww8f+P7Q+t709lH2NgpC6+PK+LkMtmXyUs0kcMMTEDtjwgIGvNvFcuPJ06h0JuUc
669Djaf2DXOeTmqgDN9HValknl1V9UdA2miktqgfrkx3NNDdJxLVehTVW1zpTtY3
RgV1HVK6FnC/D2foNvIs6dEeepBSuYeCEPP0uivnepK+uHL6Ce/SEi9kEC5nPMC7
cMcMbb3PTNJ7sxwhRCnsXACDjoSvHLbrvlMdpXDd0+LfTn14ssE+kNxcHXnhrbml
QBIkgaRrHwwni+HLwE/usZYBZ8BQRgQalh3YUCCXpJ7Pp9QLrI6o5sHP4HhsEzPc
fOZdJQ6gsN+vV6t6NxFLX2dGdAqRlWoayD4x3Dvw0VRtolFo02G+fUyhK9qmHKn9
QMFjPO4CDn8/0tknERveKQlqiimDKPPVHxAegbhKwRZFJt3PujzZ9hrg0LvWhgvy
gP41cIMJsMCg7WA18vELQqKxGf+P+kcAOQIiPbf8DO5lT1C4A19dq+FAwBT9z6ah
r/hZCLjJyk4lei8ptslRTomJSAHyLojLQ4eM+9gAO+YmPLu3PWL3hl5Z4rOUGXEE
N1eU5iPCVNhB23UBhzPRzK4H+NbL2TJZNwV4m6wVsGxTc95nIsC66x+MEo71lA94
maxTt0cPer7KX1WROUqb/E147bakzZBfW7SiGDGjXGC6kJRhtCVRisGXq72jWVsD
/s12f8RDqxOzCfgLvWeRVQeFWHUHoGZg9mLnjBk1TheyA3J9uzClnXOJlOwtFVDV
einvGtE3YgnvoTqpa/gvBPzPkTg1YPXircrG7PAd3wxxYYcwYYgXsLZKfWyLjJua
HVXHWInXPADDjqz03DFtXz42MtufjLUAG2rqMzaoEV+XG8vooG6PIhUQ+hJoQQjT
WnhhEhg9A0Y4NwWzznvXmF36l5XzoBvXu0KM/08o5z7pjuoJGZA7GB6Fkt5pm7yQ
jbFcT4o3BShuVwc8nI+3BdY6lmHDHZXyCWUw6rb4DaWFagWkRumwxkQU89uru8hr
19Z3KKrtFehHZrRKBdANNUDsAs5Zt6Aow72VaEUn8nuzDdZZjcKLSHc5xC50uLTa
ATxvuMzPjBNX/jhoTWM2V31br/JIrcv1CgYr0M6KbYNNANEPl22C6LUE38nM3o1v
W4zv8xWe2pUcuOkIpRmqHiFc1XKnF1/bPx1fcYBeKBCQzRl0IfSfEKZ/jeEWAr+r
Bwfx8ExrcWtRhIPrPrkOtBKYtUuB6nLTYi7b8BbEK3FPjeuTKqu2AhQQ+SiLJwnZ
Tw+Es944xgmFIfOkkTmlbxA6Iiq/x/Cu2SYCsBUrLmQBGabDy2C380hKxv1YIMsj
Y7EKfSP2eTIlpwmwOsQmzJF5rX4fQmAgvVgsHbbTarNgeQx2wnKxzbn3qEKCKy9L
oRoxSD2xyftsSG4zWOH+RB4ItwZJtcu5iAxxcwBaQT/Hc44+dd+KlNNdiw08VQ++
i+mOmFizM/DUuifW5IGN5K40c9V52CtPLpwTODpMg/oDVSmgXPE4//tqDoy+nJ6A
n6930ZQ6fASv1xUcsI8Cveq7rN/8BVIydk+jxqJqEIfYCz0303sMzRxMCMjw/T5b
1IrZiVCfuTUGXMURReS5ayhWJsllVvRVRJrFY5n+Wi2CdqjcieznEKgmqUEmHMiS
0CZxKpdYNxe3mKtDev/ICP3nPQz0IIrwaTdGcz9xVZFL9Ld1Sp5s+UWJpRdNWOl7
T14sDlxPxGAcCa3gN4oiBnhm+Sn5Ha9t1C9ov6i7O8EySC7e7QJdK5e5LZh9i5JV
QiQAwVf0KDRuqvnOp0Ud6i3OnOakRaHakol9q7blCD73oK2jSy7QSVFErdhPYIZo
LCwwC4UuEr2MgNa2A1JBq0kvR/WqGI1xnX4xRK+lTLSWplydjMzM00DWN7OsDv13
UmkkMA8ZADTPouA/aVlU5BTWxfgcW9rtuXoFbdf0sLHeg24IoW+03rn0EkSbanDr
2YD2rmeXaii8UJmDEZx6FeXLd+9BURC0cznOcfYn2tbe8IY76eSx8IJBdxYBWqsP
rzIg9IHgcaUxgqkvfCSDjgkkff0Uo82iyUTdEcOSeQ1v4AEHpyCSWao+wnvFBIy4
+RiAOTBp4Dm8nf7fJi90B0eOOepkE1/qqjkNaHqrUO7cPkefI5H8yZgbruTnrQDd
7u2HUrLmUi7k9Meyq0KzMksi8P7ZR4meFoyPlWLx4bOyyUtImngWOVG0WQF6Lw9N
lvUzx0MDYPufazXJXh46jqNFAlg0YAW8T8nwa9/+djTGOL/u0tQqYlzwdOfIr6kG
oG1SL74sjpA+cEI/GpPiZ02OsQqH+EoBNyMXhQEzqIbElHY2Bd+8s2sgJbXq3lrX
9cpCDib4biNgyxSVqB5M/ICosIlArYh6IBaE6LUnbp51OMN32UL9Jxhs+ayFAY/J
iwhaXH7dwXuaFrilSu7KlD7NaJifA6vCuPKwTeduc1OouurimWuAotbcfTd14ZKm
OWd9kx2eRdwhitnuiXeNkRrtcaufx3R4nXShb6+p2rr+MIIHO18b2ucjcx5VGZXs
V0DjnBTamIsrWFb7EJnCkA7DlMkrzJp2KRkLCyu/xFPMQwnjTL1VD66wkiSnaOoZ
mPkDuAwdO1TZ3tdfMi2/2pvdwHdS9wsmDjfTpB9dDoEDwyAZ9/AaDwtZfrbIeXUZ
PWStqpTuepiJK8rCPJldKAPqfMumkG3wnotNCm9jaIdyrAxBPq/b+wYaj/gRlHA0
lrDgahmVbqjPOTCuUlHAyR4Mx+WwMgTlcpLqxaJzExOJzbuVUDBlCed+qc9Rhu9I
83QVf2gqvDyk9GJKuC8N4M5VX4rE5v9vgeiwEvJevQTHTwHfeik9lpF5Q4VjdiFC
jD9RQt3wmHEFRRSoLL2rzL5dcgyNoR4144+oZZssYIlTmd1bjdNQHoLya+yl+44b
yEFxpR0THvXtP4LLNmdAnq+H9IWW1t0NLj1hUX9D+jtrQwc3mAqVgdbvSjtaINZE
bdq7wwlsXMoQZRYvrV7+0wbrZYzX8wbCmGE66efonekFU8it0LiMR9AOTMj6jQcc
PB1PSI1e+y8Xo1XIy4Oa3soP69Q3lls1Tl9FfOOECfcCSv062lQUmmoqpoC0rKh0
JmXuAMYLhfbJFNlIzF37VBJplkTtsVk2kBzjs8moS7SZzTPcKHrwqE7lVbq0+aki
KBxwt2G/eo5Wae3Bgm1c60376pLS3hPrvbmNv7mfl1MH75eAZfV8GkRUACP40jc8
aaj5MPdFMHIS19k7xSEsOiOiZr5v7ORvK/2v7xmbC7jlhALoLDuiZPuZeSDIUpN0
fWfGlNRq20kp/f/5LZMfbEMqeFRmdvG780WP+FBOnLj6qywgKemfYJFrQ5RY23d5
TZbqSqZdoDEn5OhLGlOyhrS2i2QczOYYVLjkK3giBHNoobGXj/kHHRGDrM8YWRLh
nRML975el7UT4y2OhcZcetHtjhuItrdcsOknrjcu9YkKtrDbaUyudPm0cD3051a6
0aYSYzxcAIqtlJBaWYX0NPfiex3cllsPtpXj/XuyMLbVejvZXJnYXqkhrA3CJVNP
VcbSXBB2zRyQnxhmaaa7UvBYvf7Jxs5FR/fNPLEG4JOaHsdMV4lM+ZEwuuNk9voB
oJTSdWUUgiK5qVNysxUVRDWoz2LeuKi2yowj+f0HiyQQrHST2EwcJxu3aYzIfFgg
C9CYIRgqhY2Nwq2xq264GxcEd2bqkHMcwfRpJeNlUcrkZVmYKpWnuPJorKpJBSBj
mdXUhcHxMfGIuvzsWOEiiCHRpmE6e0nx3Augj8mN5Bi+ajqnvQEfuREpBtI6GZwA
biV5iwjJ6QodmiSvWSRXLtpsR7QmjySwe2Ncdc+oZ86OW7n1MOQZvF8crw5hOjjD
pLiXsNz+3KMpPiFVoqHv48mn8/h6vV86moo2gejbb/ppm6hOArl00wt/UMyyQtA1
AmW1eVJMqycRxTnY7seG/iK7AK20SP3hKtCnJfjeaOtNA9KYuz/a1oZeCLviiZSk
n2GkHHjawnH7HeiC0TPK60rMSxY+mctItw+SsfgQvJwGsCwst0OFrbcZNvvFICKC
HGMfXTXt1k28WcSZjxY5Q8UaP53irA9FHMrjLt9RzuRqSOqObO2LKajtZY0eJvtM
YzP5D1Fu68yy6bnxOGW+bWtS6eaaXxLoInSMWHFh6vnSKbCXn3sfifVOLrCgGYXZ
Ikj/Ysy9+0HcIcFvi7KtkdgeYSeKuwge+KtmrZunpjKcoaDfzgUj+I816yUYJr1L
VSWanrPWT7VNn1ApYcm+7MRFBJc9MoU9cb0UWVV/FynrtpEB+yKRB7cqrk9FfIbk
WJOlMwcqVTWW+kZltoACo+wLjoeWzZXip1Uf6WOBm6n+ZbUVbs6CCTfGgLh/GEdP
hUOcoNVn9bfUkEPWAkZFg+HcjvIPjoQN71zTjWaMLCSHJY8n8vcMSKe2AkJncOz+
4ye/Zen5PnzNUEygW7zxOyqJN9HCZ+jxj1yLkMbogCriMqvvsAimMbiIRqDAUdGx
PyR/Dr/1Zf5sbAF9D5BdFdb3MRyAS3mvN63qjmRxIvAQLt2ikmjjJD/Oc870OUpY
PEsbrEsshICEmfakUJjDWSVxQVKnIWgiv/1ERjBoXAAVcOwemNeJYetKr9Ix6jy9
Vq7FMV4ZwEMxoQqbEA3bz/rsJ+gaihsTeKmTHc7pVERhO8/sOGk9UODEuwyEGgED
Hjl/em5HNdx9hNSotaEhk7vZriStOlA5rg+gaKdbgquI5hATQENKikEpEIiwGE3M
GqB9N9D8nrfYPlFhGUOSsBYEWt/98Q3rwHczPsSaVp4f3P4ihUBzjhau8jbiC7QC
6SYHZLXa3SKaBqZHH4IE6gBaHoxrnD50pLu8lgOQ/veCu9OGqAEPdwqL+0yRoX0f
hqYX9np03hzHQOe3cDXEMX6X4YBSBEalamW9erKCBKZJZhKvE4kUSFAqqo6UP8x6
LPoS4yLyjhvMU/4Jff3ZsFyFyaw/s8D9EI1eywozCfrO/Y0/YSgL6Tw2/3EZjQys
M6zl56M+wiTgoBYy0+ceppHiWkrUtXvNLKsGj8Bnql+L55+bH7XfqUvBzLU7SQ8H
AFxt7tEdZb3P2AypBs4g1TFcX6sBqantnIHL+2FDf8EMvmwJtHoH+/fDIrGjGidL
rPOX5TzLNclprVPi9+/SHDpD/kA1Zna91BaGWaxt1Ks4111pkB0auEBzxrkqFhzI
wE0AZE8lSLUBVhdS9O5LJ0eyxguNZjelOBb405llXQxi3RtvNhDRgKdEJ344A1rz
hJYNY/KG1LMZJCkMv0Z9fdBbIIOhxeaPsxMczm1Cpj+2MVclss1upJC+FI9J/bww
Pf/qQRDh8serpVbe+Cjz64psW01BR2g3ce6OyRlLmvcHPGEADPqLoV21gUDFrnZo
XY04zZ2W2LHRWi7vGNqTSjjR+CkFKhInKYcrD500AiuCB22mlS2H6yTXjgx9dj/s
g2IhoOvvYkE7nPZzWCyEVBAM9S4uXo896x4Ai7EUM6Hn6fLJggi9/Ja+uSSdT+Nm
CMwAUi5Oz9TstyDivG4cm4Bi9nq6jIXUjHyfP67gbCfggYnjRbQ9JUEYw09RT+Zr
0+D9sz41H9hd608q/H0zRtsAZYA9Mwm0yrp/dIZNfMzURBi6kLZTYF1peRZ42kIH
X7WEi42DP7B3XXDWF5L+CLoT2tFLQCOtDwS4GJskuQ8z9x9XXS42tDkEszWq0X9v
ZWiqF9iN5E6mML9diOTZB0zVYgmxVL+5SdhylWDy5wFxAJMVDBApoFyu/kWPqPQk
IcbR2dEv6SUOJZKmHdPcTnCl5Ia+Ar2EOewoqpdPtSsdazeadRAhSF2+8UJy+d+N
2EbCOUNBunny3kjgMZCfH25zpcwY5r9OcsAtvgpeXmB71Spio0bk2Mz04cmdRJxI
5FTiR49utTTVh7o9bJ/xrnGzkfZhQWeN6bS/U/HGZPeY92+xIuRTqDbu35cqf++X
gw+0ZoU+1sm2nKk1ZzapeqU2cdyDeVvT/f1htqX+bARk4BQPp8YZvbo8Uke4Mot4
MhnJFx+pj1zNzDpP340j3QRDKwezHPx2faOlKSTidH57xvbHljNZiFXu5ST6z9Vk
HjcyK1rIxzTEv6Mf0UaXaFX+uziHdGqbXjg6GBTk8nzQx+WEfG5Z8/pb/vm2v1zR
E7aRBKKYkQYqLroVmWPDEgcyQEmi0wVk/16TkTufjEG11XjvAm01fAUu0lUAnAwJ
mjq0ATRLE1U3wZk/d7a8tpH9GpBo37v8w3VN4H42h6Taf30BO1R9ReGIrNV8bxJs
o7/SsaP7+EHxRH7dWNU86x72bfnaa0viuWK51Y/E0PxyQOLluWLBeoH7yXyE3Yfv
yKPCFB8MBHpOfX9LKauNM56o7eFop2B0OLEo9W32deHl1kxs5AQx2+DadZQUtrWb
DOirGvUHWHK0zZB4pCuFn1MKI23WQlb7YkQJBfOw592KNRRVrzzhMacS22zQgTNF
wMOr8KMXxYa8vIYrotKEvq5+KBamWAiyS/P6JPAW6/qsQ9UXvo8Q3+Y1v7WCmunn
BbdTdFFd2KJqKH5dnBdRTfD66y//XiJDm1NZe9eerAgO6qd0DFLtwcg4T0tANtbw
XL6wvFYsQausyt8h7oSzKWJO9pTTu03m7bn/rAOxsIlojLadIvI5CttWMvV15ME7
e2d7d+zusDY1r+foTKhr3GN2K5DcMQdLiEudfH7QIxq8o7PD3MwmWK9YisdbwN8a
3LXzNlk9RJN0ySCPC6vh2aXtownwNrN9A88jPq5kahqnsoHRUV7CueWlbP12+nJu
gd4Cle9fOx6Z4pxJo+EP+iWk29GUxFGzByf9xnqHIbOVdZTqfVeIZtIXDEeFeZMm
+MSjZ154qjrNbOoVFkL/7zLqxPIDg9CZDmLUrShHalTAv0BLRmIJpsHtCiHA88za
zvw/IedBUQAnTisFDtS6ASlkKB7m1W20YCp7+74DskCm0e/7j4JE1SKOB0Ys86KA
hlmo2n4oDRnOB8vIgrCHwkuH+JMfatIc4jQKGhAtOqbgvB8TNLsA3Ez6bZzVH7DH
QUejkpGnZwYgTEXNTsI2slTBu1lj9dexc/aWXlNgvxhMjpFswk25sf/Yz6IVBNEH
avp0u2s+UUfvjTaGfMC9VKr5fmB7mwGD2nUyOU4R63wxPdC8kXWr1hCo/p969VHo
bwA+4AgQtUA2LgHBUeyQpAPQkbLxmJUdMvolZHT4aWF9RY1W3t9kvMjW2WV9oJ1X
YsBpPxj/39PQHfuiNsTFx9IiV7mZ0wqFE476zn5KLrEFASRmSArhqrysFcgg2xod
snlals2J51ndxGaINNGYhItr0VFCsfirKwK31WKRMtLGKA7FAaX6uX+n26OBloV3
Cv1vsgtaAch1FUlys8PQotkFoIPyDT0qGTuDyJbs0qKoOpewB4RfhgIJk49Lt1wO
4DjabFVQX9coOA7fLo67E+vuCziDNwR+ffkwtXIad4PrKYZ1BluuSo6RvCkWMRL5
PMtYPI8Z47vMw5+iETmQ7q13+y4x76qvWY+fFJoHnziryMNzFNkJj4z0tjWy79bJ
aoJoOK6h2NjeETbPWcSjBGKIhiRJ7EVgwP8XzAXlIv3eh/Os2O7dVgvuwVAG6qfY
RnjmzQDCYVcfAdcQsiyLDt9zqkNZ5nnvBqUp4PIhQkTCe87JdW7E8wkxJWG6IflN
72to6vOJK9HD0rR4Y/I7QYEfpbmaF6d+V6LyA1doNpjuZ2nR+cybrWBAIrzOboPc
pAIoE9rtGG/wkAUeSd9FNAuzaNMm5diZ3ThSXGvT6yiXSNeLpxWRHkhix7iCUdgE
5s+YYZxFEGaIAVWwk2fQ0Zt+tYPbt7kMkhbHLJabHcCj0mpgMYfDD6q1StKZk8+3
K+TjX5DWGq7LSPPNYOqzRein0o3qYeD5Tip8hV4f5229ckHzlHMHv2reJoWt9s43
kfOLlVRYKtSUKahMkZQ9WMfYWsdISOfyq468C08nHfmKIawV9ZD+LPCSubJ+tri8
a2g4OT00jLz7R8UE3nSanIWDxcecEVe2VFNsSYR5VKV1JFZ3aRFmFcMO7eIiEkK9
zQJsRRJTHnQ8j7hCJCbS3aWrg/Tj1ghNOwnxD/+XzFk/uq96dmsT8fmP96FXPc5f
NlhZpTU/4mbEfhH24yGNqxmcztltOCm7DrDrFpPHAMFqFS5bpx1KDf8L6Gtdjy+0
0gvbq+pGvZ+Ev/BWs98KLrAjECLUKyezMNtcSLQ2CyCm452RsYkSfGN1Eepsdr6u
GyQb80Gzp9vfjrtzBPJD4WoFeV6zroH1EJTbo0ZRh5gyG+MyqTfjUZz8RAgqqA9x
y6p4FB1BEZFstRRdCiHExAzTJtHitphgajiy7F+uG+vaaKTGnbjLV3siNy/3OnlG
eADfEIdr5Agt0pZnRpd0Sq6XlYLt3NXIjyuFgiES3BMmvzWGRgad172UGKrm8cQs
wIksiRTi5rkjmN+kNXZcUocH9Y3LfIvpGzUfPzCUYNZzOVGyK07mjyd1y0eHRhi0
Wf5cUUX3/xFdk5PhUPssoW2Qg6pHTsGmrF3SkQiRUCaCDMNx+u+kvTEIemgoaZmh
3+nO/Kf2TUk5QmC1x0xOIWy69GjfUwMhlFAW3CzVedgo00+qN8AbGW43Q2chCz4t
wy78ogln0iHP5qZkaYd0fIdnNU3I41YByI+mGkXHE06oumtuuGHa5EeRvYBJBien
ChDmLX9bWC9Q0BQxdQaccqApMqgzqdErckyyC3zAkSfpQkJ9RjXPWPWF+8tb0/oH
MGmpYyknnX9Uv+et1ZyH4Zu2iCm+4Pt7ZCeNHokMRlWdlPujY7CXClplg8JZAHoF
m9ZDIpaHG4rcfCRB8VvZ0d1y86343UbIcUHgHfLwTWvzv2g9rg0Z06jf8cmz2zi+
3ZFYzWEA3jzcrn5uRjMh7StwQpNTVwG1tI8UU3y7kRiG56Y86iCBTYlFQxQejmJZ
io+fqtPn76JiTUTdHvzNE0NVqxe11TsspOQEIosiJP+Cqnei20+EXfF2FQFHWn1Y
Ehr2D1JvNw+Luhl+UBRNk+7BMPfEsK1yytc+UxHP5nfGDT7pKZ16aH/WmTg0LVhD
htJKNWXtrw+8+eCdqI60ZHzEU11/LHt2RQ/+xDkB5wUfHSg7LRrjzWWF2msAqaTj
53l7urhYnCkkVbx4TFT7eJth89EzcFWc63YuiAiK5JnCvUPUSqzHTRJJf2LRiQXw
GuEuyRs0bs38KreqrVPRA/8vMvlk0nvP0WZSp3dGiyW1v75pTcqJufuo8nTTuhGp
/t0Jan6+iyncW6ux0NA4DARZsZh5vXcKmlzAhBG8V9LSaopVHtgPSsexT5S3t64Y
HSi4KKon76Bq/8KFG+wlP/vPaSb8taO86GV1aNXy3mvjWGf5/JBkh5iXQT6qP+xz
`protect END_PROTECTED
