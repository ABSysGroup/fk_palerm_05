`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JRQVbW4VNbj68u4i9PkqavHivR54jdQ4V2tay6jEqzWLfcnbPhUR1B4aTXn0NFa/
v1SsKxNDPIgM/iZoNQRV4avHBBaYREPPj7C0SyZQwl70hkA2IqsyoVNsD3qjDpfk
FcTYQFdU14h6UTYAiebS8GxVmrckvlgghQwZ9WsGXYhwToh4W6IXKgXgpIpAbj8F
zAGt7xMlM+DjnJdn5fwYroCIKPf/m38AsFcJjhELSpAplPqYVg1s+A3vVhGEQFZl
q1qzadpVrnoxrSYl1A+xOGr2tZLZMmPXUuuaVAE4FOKrRVThMqQTdFqnQUdut/Zn
JUiACJwK3ZmC5gCf+WLqYAUFGtK91q432sRoriprv1es2c/1RLTd0FwxI/VIT+kG
3zUb+V5TpaJ0ie5/YN9Jk6/8ubvtvYAc4BNMXpekJJ/Qzns/U8ZelBmV95rclUwZ
pILhS2Xd5SKqX2AQrXY0VBlRzz5qOhl9utLegSVmwzoaXvdc8NqHHVSa398dSRBk
FjmE/jcDRFZnBX95fsUvkwNZGfXFmO2xgQ8t5ENz2iK2HU3hNUckh0l3D/4BVq7U
LT05+cwJMb5g++pFnzg1FEv8pJApVhj41WgDQ4zVlskykE/kClp2zy592Nk0DQ75
IBVGT7iy/GbaBNzysaZjuyE8Xgi4hh+umB7BjyBWUE6Ei5JnY9vMXlS2g0b++XDk
sVeLUwLetXNuVqhUvdv6bZmD5TH9L1i7gL5dF/z/xlyUO5NhG80gD+T7Wu8N7lpV
w9Qe96VCsepoS15h3Z9uuVxJoLlRf0Eb1ZweIRcuQlGOe5HDI6ldhwPh4fDYLdhJ
T6sOVb/5IupPCROa0oXQVIqgbE3JaN02O3OW3Z84FH8oIko6bgkL1f7yxqXVSZLD
8llLdAJc7noFXo8k5bdy13EBZUbfYUY6tQjLcuAkqKCT+85gJ+y84n7pEI/O2H9T
`protect END_PROTECTED
