`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Jwb+eaieNKBRnxUgsaS5INZAr9ZPOXb7ttutDsUKHgkC8qSf1oCYSrG5rQjMeWR
MjpjsQTigYmEkj7jyd7G7B96CFs39COySBmjrQEWz94OsTApmqlbtmNOfY/OTcvC
BK9Os2BaWE0BNTSn7s0fivwGhtr0+Zz52M6Cw0FzLMnIE//dW9+J3fJO5EH6/3t2
7+ce5Hiz2X6hCXoL2ppJaRZOi4ilV08gu6ZbxQ1cop0/BdgL+cBXMN3W5nu0xooH
DGSB/v22Iq0o6NF23549rKWfosjKBYGy3oPvLAJvsxY6es4LYg68edNjf1agdPjH
rKxVKwzWCf1JtOFR3Avmy1CP4E++a6/aI0mUELqPAfKWdmJFdx/VQ1cGfP7fI3UP
4uYMfAzfvF+zFziTYMLamJJW95xBQqhDQtItRCLsaccvcK3+t06+D7spOuBz7XM4
jKeQdVmHsOY63Tu8R4++DfRUo9+DvqYdw0OVXO/wIuhdzZM54Z0l8XlapwM2LCuy
6lEwL0exT890vud+O1cOQHZTWWCf03kOR0yg5SC22KI=
`protect END_PROTECTED
