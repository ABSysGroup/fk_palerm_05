`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dZX1jmlBz1/UY/AqBqGitLYoSJgpVjk3qeo4MjeIUzSuCH1kqenEcu1hid90bp/5
k8F+3e40QL1FP0/hszmqpElcPe29HTYhlxiWYyNn2CJ0EzLo2MamqvXi2JDPh1/Q
5pqR2pj777+BlEVxandy48rUay3lxjX6u/3Du65x0RhXc5BDZZOTbdt0DZivgn4r
Gj4D9VlOMXkJFt1PZtVpkovrsrKR4XnXXIOriPqXXRKnkO6JTe5+mH/1J6c0COEA
mvrKDwi/roTnJolkaumnwmnPPgabzV5RmNQGE5lnbbizIAGNJK3Yrr+AHAF17e0D
XZLkYJUgmBADqoHeZQ0+mQ==
`protect END_PROTECTED
