`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P33aMgrOrEElLGXVRAUwQLpZm54A1lDgzPPixW8JfmkRl8VbMx2KzI/xUAwKx+cH
PKtowA26vXNk9a6Ick9bCWI5zOzi0JsihEWWns8fYYJU9gSqomdjtpz0OT7GEvCt
fYc5d3WbTUjyf+xDsiNX0zmxzuWrbfaGUpiNielO1XPp5scobfrnOQtP5TIP6Hxt
u9GSobf+/lrsmf2/HCqaajlox5l7wZKCtWASjqczr5+NqlJTqGU+IBK9HMVwNzET
7NgcdlrNxe0pPx60n/fzpoA8SxN0QIdP6x3GBRo2/70mbX2VlM78kdQ4uqZW/CeE
g5x2eE8rziWl5JUudhoKPQ==
`protect END_PROTECTED
