`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zZNgztvR9JZf/McGGM8i9725ZYfv04srPqpUP8hO9NulfO8D/c2psKmsdPOXZfC/
YzA2PD8mL9NJ/wqkUn4Mt1EhpoqJ9WTkeAJZTQ7k1rBHKGOnkQxhMfHUhxWTEuq0
bun4+gLT1F84D7rXuNaoVt+vPWs0CfEGnLB3Pbolf5dPUhm10SFhFETCWQWO8fZc
3GUKeOr9BTLgE9gAd9U2iJ0F9qDGZMKSl9wAKDHrF4G31zhdyuGWx87p7tl6biC8
wxG/N1mpSczJQhCtqg1UQC9WxbfBJINixPIrkbNlk3FnB5RpXAYeMD4LjxhzSifo
8i5d8EQVelwFr2I5cigzEcT1+me6BX+YZpqDB8C6dfqffbSbO7UflzLtoE0bHeGj
`protect END_PROTECTED
