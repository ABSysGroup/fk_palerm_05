`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ngNH96jgDfYGb2xRmoRZNz1cEJQ4smQHuuiEMvdarbUx8GbfkRv6/TeIxkjG+6cx
GT/zHySNlblqw/JVGQKKtRSXHCaK3x72sLtfQzpDBf94jef+v6BOPcNVMan45gKf
yEQiXWKUDjMGdzJRxTjUNmWeyUPKy/Cc7v9XacFFCM+6dS4HxPrEmdxLPArirIMQ
qDyBH+BMmFu1Wo/KArpVkN36G/aneI0t+KtERvQVvFQCFcxzHs+PXvBXTz+p98DK
+QRRpG6rITFrQ2/GcMRElydlH4Ygnqk38C7Qo46sRXZuUEL4wuq1JLX5lL1vhbDc
UBPxb5eZoRoXLTiAbH+QBwL6WSQLIeh7HFjId0aw19XrSYOuTYaYKEcpXJ+UnxBn
xvv0m9GKcXA0sNslddQmMCFuXY6MnXG5tN0oE0xEj1nzD4YzC14k184/w8hPtKuH
foM4uG5GQLr/QietpASPO5gK7bDVszEcd1BlU+lmwBf2+b5FogaS8KKdf9/R8lkX
`protect END_PROTECTED
