`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+GpsCpRIiRNeAQ23xOJQ19k59mABMIaj+CnkYKtmBT3dpEf8Ayj+A/RlO63vSFzi
CjdwMiE4wXPO2aNnNAUtledi9DDJJYbVwwH+/ur0FGwK6GKK6HAqe0F+0Q/LMGpR
/vIExCjEK1lnD5frIrB8b2yRzJF3ZTlosBbBo2B+KTrR9AfXOQnu46AnAPubAOWm
uY4Jn5uRgbHCdcYsqg81J8c3WDy/fNVtBFjDHBS+bMiEa/H7qteTXgPcxpm7FtvI
orHXmd7ccE8epwt4dmMV2Gm4UpUiE9X1LSLcxxs/6cSdbuJE2d42vX99gH9H7bC+
KJYLNu+Z0G9eqtMF9rycFCSXcCC2zbURgvnBLPmWUX7LkiC0p5v+CksR30x5ufQM
goJuUvOnO6+aVWsG9gSc3w==
`protect END_PROTECTED
