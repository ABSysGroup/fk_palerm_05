`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dJJchThq5f/HH2gIYBWQ5FY2Sgv3zKYuOKYHumNuU6HGb3PdaQnTolfYA9LQxThx
E423P5HDhEygSRAKL+u3AEcYEk+pl1u0VJlk+ur+t4nVYIrKWSAgMJC87jNSto71
B4c0NxSTEqPd0nEhDAC4sw6/IxWZA3deXg2ZAfmklAyGNA7tymP5vxPsvogvWL9I
N1EQrPTjm82fGbVt+bJw4W1Oa5C0RwM5+wb1EPHB6g4+OePQnqGFBhAFe5u7O02e
SluS5ONOA9LktfHU1pJJE0bxNVjNt0g2rK4VV5JFVGNonZ3jaKXs/216gKnVdliV
KpWUHVkHFOgMPjoU/uz/dXlvuD3PNXzqXfh21c3QPPvnXASWWZIgqGGVBLMJH4nf
bMbtrgNZDhH6H6flMMAWJZllwHkqC0CDRIyAVLiCCs6abHVhMbYouMjijDBGVpol
d9vqxx4ors6y8GDufuuWULgTrGVoUn2Sx1YbeyRiqmcaY47yqNMbrD6FLUoA+zDj
z/3OpcmbY/Ex3BAEjhyAeBoQHizIFqolCuKV3pMvildtgdAxBLCDyHN3DzbYDwT8
O0ZpN76QqvuLn/hy2ZDZpgrUIRGY1G96SLsKynIW8+FqVi1NCoVqF5ZrqYDvUvqn
QygZH99bNJAkyu4WiWLJoShRqtG7g3ZGtKZ5eR0tyKj9UpZ1NfwsPVdNnFmMhn8Q
jSK9rzLx9T2DjuELrcXo6gMxeruSKodyrm4znyoPyoIXjvIvEd8xf+mlc1wd9mQY
5IWyyndOjrKow3CqSmzl1sDL1wjuhE6b7W+U4jnYbFXAGHTs70wwahVzVLjA1Atv
/dUIz216UHL+QO2VEy1SoPgvMEgR0Vtr6ExMBzGYSbQzmMMzhP8jn3qxMWjon59K
btVMUaPPjNO4EVodCndCRMEEZY9fg+C5OMZTR8Ue4IM=
`protect END_PROTECTED
