`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9ImQKbhyR7N3jsqkKX96sp06UQc107/WUdeszb0+QxkFTKR2jQz2Hl7F/m7Tm29G
D+HhI/k/Mnvg0EztQrFY2Ixofd31o2DLnurTEssyWByjfvxBPAU6yrcqxaTJuHDA
KVI9l2dGNqk5f9mZohWw4h8NjQ3Ff1v9qGekpCSPndGcB3E8cajdADOJOruYAGSX
sH6Bk2QL/l2S+171EPU7JZjBRyxsPv06gw6Ux1ddMnNm3qlDTSUgRCP29FrhrOhc
F0lb/UBCMwBzD2UyuHsqLKlHbSYDIfhl4K/toI/xYLUlrhG6mUjiWBwWR3mLrWKg
20Y9IHwXgLLA0qnOMfXvB00F4hwMWGa4t1sYp1VVRjzqcmh7dPzyAuzBGvq7dc0/
R6eZQdCDykrwylwMhAhklI6nOZcpH+7Ae9iAjRsoD9wJpsAWtY0ReH52lzdEGtLq
d6KTqXE0O+D9Obppoe9oogg9NABBIdKM5gzOZ9FA6uTyPf8LHJGMrXy248+yg4u0
gDQv/79QsN7+OwnGHnnpwMEt73MQ1itiiJFHOAnSP8U=
`protect END_PROTECTED
