`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
10wNlblfDPvwe73sBDPJ7vGx4MWfo14h6AMVkrns7hmnwP+bLNNdAu+Iy6DYVylr
A31MiC+RibxNY6GTQ4Lyf9jSrI5+ZokxF5+y0B+PFSqYQ2Irm2UcXx4LS9vlYqUd
jMU8Q+s02fvmZmcn3O5/dgcr0DGUhSMEQTg/TFuIyFTlPqM8Li8A4JnyUxsvijhy
LfGki6pjK/xAr8ZIFIpCipVmoME5ZegpMPN7KuMD7Ap0oheKyMZg+Sb+MiADElgP
eY+UUgTX6Dcu5UH6N4HDxiBKn4eoireWoFPxXi+QgL9oCh0O2obUHn710bv9duZh
Z3nxxEtHgz8cHCwpvMOoN/JnFvLRmSnf2y4ZNbsj73Ys4AJ8AjP94kRsrX+5aLuS
SYzswFMXkaaNeYgTgR2XGA==
`protect END_PROTECTED
