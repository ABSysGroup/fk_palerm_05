`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F1e3LCtW6gtltP/pW+lhzEmhPCQB0gQ7jFslzBhZeKzAiJ+2MfD92/wJ3s4lWgmY
GoIpfznB2yKT+DKmoJ1tr7sj+RVUpMErf6ob733qVjw73EqTcnfdhp4T/DZr1tzM
qTBZmqcgKpLElau1iIw35IHAnmBIIoMJ9D4ego2ATKosY6PAJWb3QBxlnSEu3re6
5w+MIp+jCrpuOWjXtCM+Kr42T4kgy1sLohNAdmfx/9i0LrMKOuIjGHHB+HEsUAK0
o1OdZpi8nOMazftJwvb1M4Se/OkuYaYns5lJGaHzn/YKr4Skwdhcv7n5bUEvebL9
Lk8IJBnpMCus4ZC6uwbwZ1NSXG6rzNuKNubUMdDll0GHh9KNYifGWANW5bJVXBQ5
eLo3mWwXLD6lgu9GIfti+VR1IjfdAuV8xcW4v3Yy6phIWWi8iwxZvdXT2mgTcNyu
n4o/bLOLGJbdFg0fkBEZzi5zDzYeR41FSQDz9xiUOa6RuNcSND0Du6EvZsvDWk9H
4B/nfVf7jF42RUSWp0vDwvRH2FTO32kZjznrfKKJ5/m+hAR82NBXnjagNsOULBc4
jGf3oJ72aYOvW7wdC2oz3Ab+3ZjJWEEgUR40hVm0qhhEfs11bu5YOf8y7tmcWh5R
jcfN52HLIR/Wv1+lZjElTH9k7wOZDDmVhRNhmoCUXJehzn5ffY7bK4M9eOlXFhwA
cgESum68g3GEQ3vfqc6vVFi3Vp2JbznIV3Yk2qMe4+4b3uaoarsZrSdKcnE+umlW
8VAKnZVhFoaZUoRIVHJ8MHiI5bS7h1sTYd4grhJY3IubMdqJXIEFm1l+X5ofv3C7
E3q/qQI3i0AxSadsqTU8J19qOdsiuUfRspjjLFhkkJmRtKwxnP3oSnNoLCVp2nIm
706epX+0M5m/d3x9rNnrB49TxYFrOfHOZwoOmGCHoJwn2XC1MMXx3dj1KYQfsne+
9arEEL2O2XZAaVRYCb5MgDZkZk54IR2B6bT/abl9XzOgJp6gYIedfe4KgPq634rc
xZbhHB0dwkUeSjpVjwRfkF3yhxYqMmf1Vtk9FnyIQq+Me4Nl/xtnmAwmMhJDCcj2
ajrcO9UkYdDDtTUfQvdUsWrDiM6F1HsaOzb2S40adtzmXXWa/oiEpXcGOZORAf4q
jfVyRihpeua4jYgNAXqKqhGPVWQG2oHlHchWbW1WosAFDu1ywOLRY1R/cLE5lpza
BmkXCwe4SrU3Pn814q1ShCoadFBoB9AyO2GBT6i81QZS0R6fymr53HEiKrp0KLQx
kTwxzKZ9EVBY4toYoDFZgoPu6mRSTORatxMX1B6vs+ySIq4N8LYL1i+H1Wow68FR
JvQxG/xq15HFep7tkNtXarn9xPIbyVcZyOmnXc4yaNNDfmn265WrA1M4Z636uOB3
/zsKKCGClfJPxmNzm9o2pQwRGlN/p/Keh3G9z8nI5SCvgzz/g3D5wlaM6djz1COu
x4ZshUltR1xaG8WNEPxgeUvu+dqYL+syBjAoCUj6VbvPIYSfI9qtT5m+9PA/5Mi7
ZTYIXTT5fVmwi++hi4QWVuw9DGUBaden1BKYPcPa22KFU4En8Ekz6eZnIBJPAAuR
/qE6or9heQ9H0xjLSWN0aNkw6JKkPka2FK/gAjdEQhCmFOhDTQmiEtIsj/kuR0Jc
K8XLU9O8clYIU95HM3qY1yKDBmEtKdEjgRhhGNQ8nAljXXzyAKL0/weF/W1CikhI
jXKSz/ccBQUhdRSUfx0eagptSANKLB7jI3PTHk224JNi/te6Cj/63MEXX1tJ1tHL
RXSDfxIt9u8OSfjk9iRu28ifALXBZW2D3+JGvpvcK7Rr3vr8dBFfYzArZyWxd/5W
btupiJ8dJfGKmfGURZ9mrsFRbvV12q6OSj0dnRYdM0LXrmLdjWGu/AyFf0esXKnQ
7PizQFfgrKKU9IFduJkjLcT7lbu0ZFRx1AeRn9mRtTwm8FOd0fcnzhSUYsTHSrbh
Bj6Sut12THTB7bFvppm1OA==
`protect END_PROTECTED
