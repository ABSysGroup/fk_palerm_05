`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
snM5xvsnK21Vrs35ILtwhj+WJvLCkKQvlUFz4PfDyRnl0FjH6VXRMHkjjFNSiRTJ
oMNXNUS9bPQxRecv0tDzgbaXHKIYXO4hTOJs9OKJSqXdUlsOqqbN4Tm7fOe73TVo
oOnTTM7Dq51msC7v+sXa/k2QDfveNRAzTOtt/zyc0zWOk7SGWVsjITZso2slP5nf
GCOzrlYgLg9GttmGtTtRHSTfAa2S5MFK0PUUNDkdsV1jyY5Vcid9FU0Tz57qtROl
x5URmGzlT9z4/3lFcWJDdL6hj/54jXSEAewYDinG19y0xiKx094NFDi+9hColpiJ
0uUH517/Pn7K8wuIwrJORgrT6FkuUaU2HN347uZEv9+DeORF5udLDS+SgAQG59E7
IkVEKC9RArMLm5BVg3X+RrNLZ1y4/vrZNfPquPInIVmGKG9TGlSsETEMHJ7pF5I/
dNfV2uZm4avozBaegxE2aD0caqGWWeE3M9IODAQSZaYgIIY8CSrxPO8xHN3sgbFm
wVCQ+n9jUIkgg38wq984rlohVEvLxNScbLSPaLn8Hi2Qbo0RM4ttq/paiv07uV0f
dK5Rur0qv2lFHUgXOx/NsvnnqgoLy/IHA4lD+QNCif5d0l756ZO0HhMk77q14xtS
QQAgh4vNOqcQYk7iTLQyju5z66UEeBIVUn/W5rGNgM39ZSqrP/AMJ2vozyhHWsKj
49ubsMYcLmM3cotVJh3n21++gk5dq1fxccjNc3WPxC+bKgrf3m1KPvI8ewDt2CEm
rXwxhJGH4Gbk94xHaL3M/fere4WAYbuSMk12n4s1KyaiBofPbx2al797gmW6fXnH
+SeHcZ33wMIvRpnfqtitRg==
`protect END_PROTECTED
