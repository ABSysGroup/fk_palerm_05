`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TU/sb5mzGlkwXaE/vxClINnfKAAy3BMNOun63nNxLxyAnFmtQcJUjUvJX5XnNSTO
vG047Bb/ulDITwvJWzAK1cDTXJfgjjpVfoBzZDJrHbvD1eMQ3Hd3PURyDaIz38cj
IBAmvjli42/bA72VJJEPgptYGIYNQxhQMJK4NvGOn92x0qt/JSU/BFK33xtz9iA1
CZNc67ZUp2zx8EO7TP1Dc0xZQUYCjx+avNyZUUXdGYv/BbKLNWxuXUCfyLOHbFWR
bhK9a+E/RstihMo5yKY0/HPOgI3xUD0wGhgYcOYnhMeRvPBnFxWEGMZ2Rpzc3Sm4
udqDyAtD+8wjCn/h9U4v5fu48SUnyk7C6BHZn1rCSBt/V3LY1bMY2s2EvtLzpITY
`protect END_PROTECTED
