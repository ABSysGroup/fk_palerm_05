`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VVRUnEribNH+KEfgY/BM40Vn+ehvVothYyvG7W8Rnvu/ryZOmmqqdl4uGGfJbG0x
hoXs7cb9k+29Vq2oKeAlQgJz5K4eNvUUP1IwyXK25nF2cEZGcVSBson15Ym06JkR
Tnyiodmd+mcYI4HGjCwof6UD5PcgHxpT68QHKj9xe1myhF7AzW9igw1Yaj1fgv6G
8w5I3u2j0acanBmom7CEHiRgoRrEKGCNhw9e55zIHVAbkFGaz1ef0fsgH5axYtNh
v++07b8m/JL+AsimmHByz256yC0f1HV3cCcP1XNfIBWNww3/Zz/YmwV0FovJxoy2
fWlYxCX+owUM7SU0ogVJUR5l+u2gDrh7Pt4isUNB8m6c2YzYrNo13kFPLCXyjHOK
51V44UwQWNu65w16VbOewqtnHsxublYlU+9DiXyeeJ0mLQemfwwUSnGaQVU8rBJj
pfVCLCFrbtlcwFzFjyotdw==
`protect END_PROTECTED
