`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2h+62dMDyJghAqxC66/2UFA/NR+gDIbNFpcUqBo5qvg/+WnBDiHFAnh9pW4BUPhM
2fU7axT5kv+GgY0V5P/QUKuncPtuAe6PcpFEKo5sge9hPfZolCtk+cMJbUUbCEBu
2ix6nAa3yY0Ks+gt2Sh1rMm8hA+zBxYY6PrXwPqpRNCRYlWUI0lPAopw+OxrFOYk
F9C8WYxAMzQ2+JrM6RULkXlCFdMOZUEsR1ND5IQy47CKaagRhaAVwpYHxx03KzM2
KT+SUSP9+TSO5RbU+pc8Lkxz/FAs6dXQZTzi1P2GwboVsWDw/0MDnO8FB+Uwh4TG
WQb7JvamQJj+jUY1LHedCjKFDnrG8Mf2OrQEVMdQti0MPwCFXzZlMhUUweCloN58
JN6eG9JM4W9S69+jxdJU3+JDPhBlLJX5xSAbqAdP8P50ag8Xtdk+vGQgF0+ut/93
PHP8drIM7bC+NfIRbdrU0GnQcgvJKkYf/ss2xPsJsgDkLDgkN1fMFPYCT5SoYKE0
r6vYcm773yivxORFgHK9R78TEmZcDV2lbSYUVThxGLGzfGfuSIqnjtza6IAH8szO
ws4ot09OQ26B+hZrHsj05yRw7dEHHIvkbnETp6yQ03viAvSWPGPRE0+2zRbiehHg
4yTNDZUnnBj8uoWczV2dHcw42ny62JaiY1n7GSQNWRtYNHCx0lsnCJHrhyiLGYcS
HQ9mjxNKczi9yXaGep/ACQ==
`protect END_PROTECTED
