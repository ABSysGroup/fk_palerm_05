`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oflvG7aEFdZLxDYXPK4J/hMF7vy9MHfjRWIM8nrwZmmROVMwO47ss9eN7h3LMQHI
E2c2QRhsWmQ43dJhGXb+45D2rZw73vGWYXnCdHD2lpjZxkRUs3YZor+a3XN3/rGP
8ADimwy1Xtf7CdKCwhG+K/rJskUSu9s7cgsKyKmDcmDD+NI0j+OCBO1Kbok5b4Dk
yksS+alpNPKWo5e6CK3OSon9NgQfx1Vn7F6NcPOtc74UwsxPzgeGE5HP5TA/rcWD
/FLrhm/zI5OhCVVR23uPS35THMbb0CoSlGOjxdWGir9nDMTZXpV5+ZTcMp81HS44
LDj3ptTEwpfWJ99tdVhgXDBza7uGJX4BRrW4tPr6D3gR6zk/3g07Lvgm/t6I+KXZ
qI/iMfSZjvQanhwv0jXN4apjfKQ8LmOG38ssDNc7FaIveCsx0iy/X3CpGrbh11o4
jA0/kQNS5g5ys48vNW6/VuWaPxlF9aDmj9ou+rz3hkMebw69CZE1RtRe0PVOACPc
GWKsf9uHJCZVKihdvubn8Re3/0qCune0ohRxO7/rS+7ty+wiB0ZoUpeT2JIuuhkM
tOeOpBZFBvmeZc4jWr875Wwg5VCo085Uwxf4IqJk3SjvsSqq97cIoPi1EZEDSr1q
R3xHO2jVET2TuLksuhUUxIC1cDPXISKaB978d4awoNqNUUDPh9jyvmb33Ts6yjbR
8Tdz5YkMTbrzCSY/fzOU2t/oDGKwBGzR1J0G07/7ob6M2ZFShY/+suz8i1TkGjz5
ZPBMrvZxORca2KfPHBPKhLTJD85JdbM8qSmQW13Z6NJXytG07/QujtxL+mi1Gwde
4ig1w5Qh1+SoINJJE4i2216J1ldxbI1ldyWlxjA0o6wNeu+aMqDp4T+vYDO+IeaD
faG+sHVe4Av1aWvgMZcbWctb8jkvJL0PW1qaNT08TpwG24G4DVP0qCixXgZXlKUI
Mpmu6qeVOvPabUppcKK4MILOHCbADBd4//pBK3r9GWyXbvPiUwYEbvklAwo67ROp
2nfqZak2PTYyKCB7HjYS2lrZjmVqGEE/MLP9XgcIJUiCWbbFR45L+DGWucdW40lu
e4NrC479LDZ3FodDVWR0Lw==
`protect END_PROTECTED
