`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zk3c15vvbd3cEsykRyj3k9YtUXaEIjmHRvWXSdiNpEJyD/XnNZdaYjxMR9+EaJQV
9EQEyBjihCdmzXiengeSRV7yAtbbjQb7gHyV6+ElrnND3Dswf7jvJZ4yuKIS61rz
gGf3oGyyxfpeRWV/TUa7exqER3hW40N031yTmdmu3WwcxXRu8k3FlruIEWTl3fIY
XdmgAvDbupKh3hwWHesyrFUvUSuRs78RlU+7HJvHbgnm3m3MzyLLV9+FE++ABgrG
ffl3Kr2vr50Zdr3uY6Ye9vTFzLzMsh8E+/nd0kkb1PPNk0jh5i4EOhjNhvzGMbCW
FIhJG4Osh8+/b3nus961XfByBVJ7v2WRa4IRCrgRxOK5RzuBhNMncInt/rPDoJ3I
hGDgoWm03TS7WvOUNRwcXbphLmzFetZeeBKZYVPV2YRYHp4qbfQGMu0PHVGFmpwq
eqKd7fPnhJXZS9IngjlR2Ojb3BmZu9LZ4xglQR2E+NVCcDTAqGheA48JKHrsd+Gl
vHDtHoEfNqD6bHOYenqbdV1HmJj2r8ahlCpYNSXPOA07/+sWx9WjnU+CGvBNwkCM
FMuvbF4Y+l79b3GfVUlvn6sC40Yp4ab3Ea4tKlDHBqaSl8iSjfgHoZUKsEJvZgmu
UoSLQg4cbpW3Stdmwhyn3cj+HbEDfmlFS2hR2RdpTEztgdsGUT8tdeXTB6tMhr4f
dSCKPG6R5Id0ybZHy4SRhg==
`protect END_PROTECTED
