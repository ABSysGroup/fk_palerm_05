`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LqR5LAkR35/E9QrU2UdN5pHx2wF9rkxkgK6DEDQdztUKqnMxt6rwyEoaTsiSnlgZ
CPQrlXVFYE/r5NuqanSPwvvP2uRi/y33ivktwlhfSyXbBUDikBZR6qI4VFKaYrBB
Faz28/8++go9xHMUXr39VQ0OYwLdsur65GZrEBebx1rzZ9jXc6zY2IC1LQZPfeIE
HNwVdNLpMfAiqAtU/XWq8T78rUwOi9VGkdNidgCs7KAlUo9jtOfS5Gsv/mKSGpna
`protect END_PROTECTED
