`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rLUL82rEcyHir8edf1dN4QHlnAOhz//uWGavw6foj0XO3oseS74lP9VAN+OWDAXf
pBghU6wfcFLtFu0z/3cf8ym7Jz1HjdAyR//GpqAYxzDykbXPiNNGgDQZs/fCtzhR
C3G7SkCOgJ+cKLMVpnIECik4x+Cl+z+F342SDtV6AOqCY1O/SwR5PIJ1KgmuiV76
MBKVxpfNPGEezYfyZG24djnlMeIsvyRP6Dwu/8fEuzrgimaNCqQ/OIWYQw1FFDsB
cVQ4zyfQ1GcYUVBXvvt0Ap60B4xvuoYpjTqqM9xim4qyU/RJuA5QSor7j8dUamqQ
zqzDRBYnrYkKIUj0fI2k/IyMlRFBGXdy0njVYLcINyaba44Mb3kte4ahlXueLXbY
+7HZzDjFpUZMtThhadPj81fcep//XJ0qmC4Y5pfWc4at2Cgs43ANVFSzh5iqhPwG
XtqctaV+SxSKqLPngqQ3Gk+d8pUCe+DF5zCi1uIrkcdcEQRQTkhhHrvYl33szcJ6
Z7fz6iHcA9CV1N+/P9kSzyHxR96TBY/d79jLFC4ykLE4BZDuLoK8XinpkdTiPA3G
aYn3G69FzYY56xvxdobgzv5Kbf0FFcX/ZFGDOjA80JPmeDIs/eGtbEsnAcLGk7Uv
nBskd+cNwebyfNNqaTvz81Xixc3tdF9C6lZXd0/V4QZJn0m3MCLuOh8hT4BJq73W
BpVvL171cc8MGCaR1f4t6UuVGsu3qCrRVuUpLIOUgDXlzuZYq9pWLGtwFvScT5nj
QODhUZ1Ib1SKI2bkECP2YcYIBk28EacvDQQbHAB6IJtI4hWMlaA561A10B0NwLwM
ZW6TI9bggMX8LedbI+s7MkTu0vFgeNuCtzAhFth6g6KzeJzLmXarrrUURlDNUVIp
+mU+V5tQycGLnf5ZQDT9+xbrXCfLkxmykiv2JP7L1/GkTPkfMn3eI4LV0bwKMM4v
tr4XurHI2+67t7VT79/Fm2oikAuCKvpe1S9VsSKJ9xvFplgtneGvFO+5wUwS/Le9
RAc9LEm4Xvge/D51qwrUC1vDI5pilfPNYI0zQmKdVtaIvJlon0ld0tqLSYRzeurT
0/IC+7Bm7w506uP37v7JdMdiSCa/+a5EJRGijh6giwAPcA/OJnFnewhtta7u3ktL
`protect END_PROTECTED
