`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8zgD0X4ZN97eoW1/A4O6z7OcOfnuUARP3SCHI/Lu40D6LW7idY0L7zAwiVHwNfia
4DHaBSBecx0RR7913tr9ynrzt8w8AvcHKhNZ04iDdbcIHGSCoEZh90AkYXhy7/t5
D6yl09eEP9TdST0qXjL+ia3vCSf7FFAU50pNvQ/Zr4n2DQh7pVSRO7KrYrJRxia/
3NnPKzIn6elaRWm2yLM42RlPuEkfL7KFtmrmuZanRZDzHjp1w13NXyKpnlaVMA6f
HmkI+BtZSNjn/tXCyC0u5dXxN7Y786HrlmQFTVRzjTJ+1BzxvT57lwnjWvtZ58QI
qTMrPXTP9c4TsLVnM7j2fn0HAIxT2COxYXOdjLfOUY3l8cm4+w9qU0H5dodbMM8i
+vQisUpKxMvGXoIrdBMTdLuN7ZP6mnjoyEb8mJ6G/trTNJq677MWO4mGelzkDC0w
`protect END_PROTECTED
