`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wfjRwHKwHuTtbAxQpYJvQZw5seX336A+ZytM9DmYGpIYQLGvzqsoCEhEUYSZeot5
pv7gf3z/1nIBzYwwN+T8wrVKhEHg/dkQEHpSHYnfFdNz1NL6Ugvy0P9cHbUJJtUQ
iRHuXNj7r7ooGcnz+gbjuL+93/Zf9qH6Ur93V8AP+/TTs5itKMGYanyv1VMz5DJf
KserWFXYhyDFUjg8iq/3N8tjd8X/2ish4RBu7xE/CRwsS/mnRV7B2qkBB4/M+MGL
A+w2NNC3S4eYYCDQXPMsa3dsekCSc0A3QpJP8gZteweOTBUH980DLRq0Kj4RAXgX
VT7lFGpWYc1TV+P6i+K+uuFvjl1PWn0CFmDSWz7POqb8BQLM5OoHh+hOmxyW5rLp
fR2t4FxOmL/JKYY/ZRZeIDa3UxTrnttNQVxgsVEJI8FBCvlldPobNdZ5EVnCTuN8
kJwtJI/twUlwVuf2B1HHf87zcycBmCQKLt57fqQFQgajuO93+oLhJ/HNOIpIdZE6
cKwJoDCO99cvrVWfUe474elF8Qjpuu9NWGjdteYtvZAg5ZxSH4cOlX66lFXQPfAI
HQE9cGoAHxJkssujWnfO/aW5Sit9Nd/GAWSxwWkvhk8/lmWcEVWD3flQmnCSSTi0
5/kkjljTSN3Fq91rMRW50FZnUpQ0GbTeS1tCQ1I894CGAUyhOo7dYbxAiYtr7Q5b
58O38jon5oaFaV4mli8BDHAEYomHxTIC/CdUAy03ROxsMmFvR2V1NSeEGQPUH2PO
zlD5k7G5YZkJtKzP/NAziO3zW2yzSqhNlf9VgpGZXGhMQ+ZbAXLlg9vB0u9jcBCE
0kFWOD1cM1zqhBd9ujFKh7uknECS029iroyBRT5g1o0JlxNof7E91wQlkCM7cL9p
KOt5QKPnyHpUCX0TWwNkdw==
`protect END_PROTECTED
