`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r+9BllUPajmhfyYmQKEWvolrLzqW189q6ro+TzTDQvZr+6GleI4s4XxBzDW4F5n5
mGo+0Z8DZEo/yVkX4p42cMkDa3prVD1+AT5lQ+cxzCcBMN16KQkSkWu5aMHyk9hN
FfG+qYTlNeS8VeLND6lt6PTLOTejTS5PMvor7cR0FR8NO4YGXYzObh5FiR5I2J5v
a64ErSeSFYz0g7aezu5nm2lB5GV8OFlcVHK4h6S0cpVR2ZFB/0uJKnLxOG9xQw22
yLow+5aWNbk+gDM6OCvt0OhDnWTvMilF8EeV37/Ut5nzp7PAgGxamEQDtDxmvLn7
nJyaaKn8w6gHqEnotW5KM17Wwn1AUYLWQDVKDJ28zoT/LjnLfOOTFarmlTTfv8H4
P42QtBakWJXuw9EwP8lGQ8ao658pIUQ+KSs2ONmFbqKBOPDub5y+vG3nP0a7+98f
fmfeVUwoLX7WYmBZ6cZQa0Cc8ZQ3MkUfMcf6f8mv94iFkx+vgNMg852R1urbYooc
XQPRxSvjYLXVMZCHzpnsiV3CrvtPax/09ZrLx6Awmb9PmJnyVb9+aKV0fqdeikzU
sgh7iQ3LltrpKBUC85bqiT1nADCsGpckeU37rVAN0b0eglzScXtNR/7KUIE8loWK
YpVviVd6d4oSnyss6sOgtyShbBswDvDQ09Ztdfi0IyBZqiGFPu9c/Ga/KLDcpkeW
6OeUmv+oSwZnQT+/PmNm39WqHij+5xtZkMJL5Xr6gJ8FMjGReHpKOLkfVnVpCH88
olWJJ75N7jiHgBqTHjKhTRsQyG3u3aY6iB4EIPRTqjzBTl8vrlvG+UtVF9nZC1Hv
9W3Hoh8xMDdKvLoVPHZE3WGxuC8NNPP782ARIRkkv4ojoOpIq4H7QlY3+A3uAJhx
`protect END_PROTECTED
