`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eQslCRkGUtJ9DEiJsgPZp06lrW0Qv+91r9T+QMI5Qvop62EwHenQYW6M69yjiGgz
mpjCOnnzb1bIr8uEzd9wK7uoK2LVG/gV2KiZ/9eADAD9jvzHUZccNFdG9GXxogT3
W3iS6ExW66rEazX4h0uhmdHl0F3ft/haZIwyzN2zioXG26F4mER6dsTMJYa5R6Ab
Ewfjn7+K7+z0ZzHdVnqab5L3kWHUgH0UxOCYAAD/fcrSSAarpgJLs/L2I1vdkewL
N4qISM9R0Wwuxg8wk0s1AyPOBO03glCzeAaHMKqdxTs/8ubrCoSVHS43usyckBdR
guAmkbDobQHl2q4GIpAFjszxwcp6E7nnGutsisZJ9eT0jm9N+6aJ5dFMP8hSMNFl
vOsNCaeXkXCMZhJPYXkbHWnntLSyfd7oa6UdUvnS7Msn14bTYN2RF2bHujWNfIbR
LKUyt8algV8u0erxlrEhVqZ9Co8go2Dlsy8r+wrKQxTYH23baCoNOgYqPBJhj1Ii
JQ+XIurARj/bdjmC8V7OHwgKP/lUa2rI0MEdSXVD4dt5QUhxMIPHQmIdShiNyjOb
ylQX42ToYstZnWxMNMEJYeUCIinaKLxZNzo6klq4jeA65CU9N3eetXB469w+x7xR
EHygrGJJv4G3dWBKrbCaHAhmLTDeKhbmJ2zlosPqZcM5JqvGS0veb/MvA+DJXkCP
Kp93l+EoyehtEwaLKwDUwHoDDx7xsZaOtl9MV7t6ezN9VtBHfLHjILzpc6YHx8xY
`protect END_PROTECTED
