`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x6F65xAc9SZ+eEcq4sdzXB9zbbQ+sSj+/QUZ4eI1jozeAC+dUg57qzikvSmzHGGG
NWFizVQ5G+JddE1uIh5+bNoFe7WqWE6iZ9v/IS7dMio70GjuxY2hKMACzJ/jGE7F
nCz4OiVCYIMfDQUUqJwlB5inI9nAaLJQJGapDMNzaC7vT69SOa+ubLvYVEn7v7mK
Th/JzGq6qz/2FDHJzM7yX2CUOSCXcOORF+LPXPHVR7bjDQQEtPxRa9nQ9jE3AwBe
wKyglL3gER1GScEmhZB/7O//HyZ1oZf7UHA8ot8oShYyEMbCZpfMo3k5oQbhox6a
5ttOKaGy1WuHxYFBpBNr4g==
`protect END_PROTECTED
