`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kcsMRcPjDocQomXXSW6QPIEZeRwS6x+/wFMcJP8Crcgm5otj4ahoSF1vH2Nzr6Kx
Z3bzbNB2AT7yFjDif9llBzWnk3WpCkkGNoTx9wn1ZxLmUq3WgNpPjBt6aVx5r14B
drnWCT7Mlj/vZbgYMjPcnHsHB2iwbQ5yHktU4WtT0SWpyldRFGIyiljtHYDb88ai
+PEDoQ1vnly6SG3iyxvlDYYxv1X18dn/Iq5n+u5PfUlO4E3es+5brHyJj/6pWC+f
rvzMGbVv5v8VqW3M15GdVLSzt6iO3j3IM/OUE+GR777ZDpOmS3Gptbe5SLsu5cQL
WC01CaY4Y0Tt4jHMb7tY7DqAxtSuRF/Bpqh1cQvZJk278hXwf6A03qtK87rsdXf5
akV0bwP+L1uqcOdr22CwRvVZnaNrAt2+rkwo0C5u60lSLvN5q59TIM1C0CiCiRbu
oZPorsdGm/Mh+9ravSNbW/cBLvqBHWW4AmuGuz6+5AVMel3rKvQc2HUpS6HY/XRJ
LW3it6kMYLfibeT+BAQToXv6SEdDsxMrtXqgpeDvIqERNi3Y5x3Dj3c04NnyBxrN
+NHiQAA70/8m2Wieidz64PQA3QzHR7ihRyjS1jOWc7CaBRteU0quUHB4x2g/cw/3
PEPWt6KCmwmhOifCtZqvwRzoMo34/guSfVdGJay7Ym87V3zKQmqiwx7UyICadEyI
vTQRgDARwf3EFVpm82nBoSkpbzJKozeDIq3Bfe8tw3PPHcFDNt0L5wb7/eovve+a
QMxtEhYaT2IDdBqeCqXpGeUBo8YKXfJwuGNm/zXzuIoX/wuQEFPqV1BhUc3yqyTT
9/9cuQHue7ZcJdbGEfy8TzkSewhgRaGfZGxCZscjtZoykRevWRSGiyeR550qDPEn
Y71l7wQfjyC/HgVo/pGU6HaSlTckKBs/z4uTJ9zlPzcS5rhwDzOsFYRzkBQxhJ4V
`protect END_PROTECTED
