`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sH/yGVUI8SwQJ7hSa89+zDg9/yvddwIirXqsoTvMcj2T4FN/05EzwYRCFhhEFYFR
erC69ZagxMzGE3CXTIbVyCG2XZnGbSTL4cyGod2UnJC7wrihtl6PSRaAf66kFLCi
m2rJ8794FwKvdY3ecHjccXZLt68pQjdsl84TxQO/Em95mEtdbrnfuUk+/pgkNMPc
aFAjI7SLKgHzatUdlkH4XzjUQV5hfI/HpPSy42UhahZXTv7uJ0/2E6ZfkUXB1p6s
1/lalTYK9mitJt0cELILpR93KzuruGmPQZvO0c7hx1bOGIoBmzqbYv1RmxaoU4h3
sZQhSl25EHmwk5kuk8Q51WG2SarUVMTRtpVpGrbJGjfdJ4eAS230cVxW/HWyxQ8j
/TnF63zXDddOB3OwKFmzSiHJBjfzeXMik1bo2Cc+9iMC5LHbKeVCd5D0+YJ9ZzEV
U61Kc1S9aQo32d5q3liMoLHYBEQPgJhfNnBISzO2BjM2TzSEIswn18KCXrHRQPvS
sfXQ25CMYFXxN0sQwxKBRjtePsPzYzpcHXO8jHlVjJuhUCWdSDAr+UFnnmpftarF
Z4a1GlHDKglE/sZ9udIzWa7pFi2wbqhPwYwh9AMGRhHoRCUCtO2Ao1QnaPYhPwRc
ch7WT/g88+XH580Wfzb9jjq+8qBFrTeKrfstvl0g7kcNdnZAik07Yxz6qKFTNsrZ
y1GTKDQmh5tMsVBQQAG5PuWE0Vop8CkXZ2iupa9Uq9NXC2E/yW8mAaRx/ZgVht0Z
UyUb4B/0Nf9ANIeh6/9R9sYZ2TxzPET4PY61RiWen92zqD9jFB11hPDJQTIy2oXC
3igzZTLtdo3Lhk59U7Ab7KhjH2W/VwyLFRyMyPbuXaojUzFvZXTAIF3zM+8xDt2X
FshnDtU9FPPPq/ppdhL+EsRPOWKcjJ6JmbweGdiHzR/73IXUQDGLGYqhY/Z2iKMC
TLpVYac8clPh+/HQh2gZ74LCMXZRV+Gk8VETo+/BiDE0Oq1Cqbh/AjwfCWWcdrjD
iStzqWkoqMvk372f1OP9q50+XcujOvgZgTEpYkNOY9odDoH2MtZSboO5LGnluM3o
P7Q2vCtyCgyWnfnxv96tbYNCiUfo5SWM9U0GLv4XeFWxFK+kmGJG9zpr8W04DpLe
bJ1V1fsSyuhU4LaLwQ28RXz9vkfm7vsKFV4o4y4vlyTVSoDYhApWQMMckTK3bXVx
PCWL6ESBVDDsLyABLrsko6MeHs67e2Lm/CWGf5ueOeHnm3WlO7j7Ygia6olWDbiu
nqyE3IRFKVijL9BHcjqyofAXhAXgIaMRPCFAr1ZZ9HPR8dSwxF28fAv5YBcjogNr
JJwrsTCyp0K5T+1g2AYvCtz0e36DtJ8NDJ7bCtdo7AEJDbNg7ppL3kGWYIJB4ngi
ZPpbLxkPG09jI+ehXuPV+uG7oLNDQDlqnLvuj8D7mprc9ibNXi7WjBry2Z/PCh56
Dp+bFT1ZzO8CeYXOHa+dWskgEX0TFoleKbpE9zwasCyjWq5cPbGMcIJzCqx8NQlL
2+tKzOvOdf/NGxkRnaudqFhbv2/J8nxhKVwJeyybRQXkNGtBfWF//OimHbbLVVca
/Q5MOPIp/1QT8jbJAE1gbFJZxs9Y841KSZq3TCW7FhE84sdjJgPGHM4BZThxVpWR
KdRp9SjF5ncVnSMAqqkSzwxSOZIdRMXP0Ts3iG12ac53BNYh0xW1QOF0oDXGoNmm
P66VIIFVTATi6fP3T3tLeC5DlPFaPaGwfYMqx1nJIEhMoa6u+IoUQ4HCCgatx1J6
7eR+uOUJwp3L1biIDz8OUN0oLtYDH5g1buGt5sBUC2Aux+j4+GCPO21p9xADPt8r
/Qb6nEt6D5gtkfp9P7jYF5XFBw6oDlOeqw/wb9m+c+742SjTQZ1cbQOBH63eVflu
JnkQbz2ElW6+rXyfsriChVp+zafU1I9Pp1pFaX4ti6cNFMwq0y5p9ONtwhfAAiJM
SY77HIckuzea9+fqoZF1yVUEtXG383LnAMONNddgtw0zq+vKN2DtnEifD9KZ9cFG
6VFYZf7ZJVhe6imUgh43JT4661mYc2CPxfLP/f3kiSMZFZF01fUqe95hWDrfeL/k
H0QajXNZrIDpOU4zf4iyGe7em0McXqVqtmdA76OxOMunwcMhAmlL63MBtpwNzPiJ
/7eRHcFy8xawMydyheaMmGDec2MohHIF+AMCZPo/ezc9wviHOPtc/XltfzkuZM2i
EuF0iKeT0N44jNUbCPXZJGm/xJlJ2tSNr8KC48oJCl5mjqrQY/D1966HW7U2lHmu
HPAXgcEEj9EGW++5MzXU5sAkAz8Bqpji/EIIgOLrbclYptG5Abq4kPymu+HOUtcR
QxPanrAuOraUJisbSeHxDs8b8d+4CzeW5VLDA0aUqkRW9kFEOX+0WQ6gpHW/CBn5
At2EhH1YfsVCHc2FQeij9Yag6auUk2LyMdhCLpJnzwj9yjwcsFWy/dsCiojOejhn
tPvxa6AOXpJAyl7QBA3c5ALn3gX6Lx2H7HN5JJ3bkmmK1PiBwcu6t0cHaMz4bVnk
rMQ/6ic+OFtQ7SGvvB2ytSAmYZhL+sWZo7AiOFhoJFSAQacUjBs6L9LY55axiCKz
eTi/1wTwdVz058w0WQGSv2FZP7r5vpOWJ5LZyswjbmhc+BI6/ntjZJu5YnjupUWn
qH4tu7ok8fgA6aoluKysBE0GAqFaKGkrXlv6ckQqO1tRd59rNH9J5mZzNRQiK3TF
QG1VsAeryAOyIu97GaAysuhQ2DLbw5AMq8HFvjiYo/KhGwlOjnYeHFDorfv0KDuH
ouSVbyzGQ4DU4OMA4hRk1ObPZS87U8hBKHObdmP53t4MV1cyrdpkawokJ5KaKNML
`protect END_PROTECTED
