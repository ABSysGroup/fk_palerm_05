`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xueFvqf0TdDQ3+Xddv7Qd9HNDCb1UUO1G2GrdWkvvCHmT0/aorsRa0GvZfmLKJY4
cusDsmVlsYya47SuuJGMb7PIwfg4PL2lVWccHxWFmLvOTXO88+2tjlEgM3mIBHfy
DZnhgm/nJBP2qkTo4pdIutn0a13eebcEQIMpDGiZesGo04cUgq1pZsgFBL/+8RYm
fnP83k4rIotqkwkfmXa3Q2XzLumk024XUJqvAGOA5Iv8UjVNdo3XXCy++FmXCl9t
1LxEpgPOIL+NwDEXLfbLM4g5DFbINa2ZpVGSs+Az8F5/qGwvrJBHEziqj6qBukx/
2fgEQrgUfo/tMCz/7Ix5sa0nfoovZ20rbgnvzb22MWKHxrw0+tVz+/t9Fu/seSAe
2A3t1e7mdpgYl+zYimqTwyDp+WWC2z/QlAX3BUScydMluWqhbFquoc8YgRTbxv8o
HmBgY83KWH3UvBSLQ6tbj72Yz8SbhRxTih1YNMunfo/8lf7EikIUe4nFn6FX20iu
Ke3kaV9nFBu0s3vDs6NfSnN4Tfc7ho/WDDaRgS7JMf2dp+IoRPH4o9vL0rlOdGL3
EEDwCxF6GSzlWPfzBX/YmXvBX5rtV4O1nYO7fS+sUunDOGdZJrrt//yPeyHf6EiX
TCbJBNc8Rd+7uenpcB/P+OtTtaOaxHyA22vABuvZvYRvmFCVB+gl80avlVelCKTr
U3lPzxrAhL1dwXgQHQhGX+xlyOqPRRQt0qo8oi70S1VJwQYvqdnqGBXT+sVO9EL2
Q7yaFYXvRPXztv2G6eJ8XwOVMEs1LpCnbzt1zJHtBoNy73eYYXxa7msCX0MPZo2n
zksWtsouiYLuiWpPxOL9Lxk5SVD8xKl6++FmQRDeRcpe9ocvKubSYRiuBrhEOx0n
Lc7xUYUPKaRPDxvAe2fp3LsbX4FrvqnXq+dYDxwOdq5JQ3N5B9Dw6jpEUJs/1kHw
1lW7e/qaW7JESMqMapSNt1uK9Mn3DAfwoLbkJVlzUqhqSo2QpQ1lq92XuPc7Uew7
DLs9EfDOYknIvQ4JS+8h7wFs/JG2ywl9QoxExbSgnRDV3ABgI3C6k+FTRt8GGJgY
F/DiJFzCXlQ9eZiJ0Yk4Qes1ltiVgynnvaGaWebCXZNYmw8uQzW9rvzWLIdWs2CN
sllFk4s5PQP0mxyA4J2InQVlODCclvWcYXZ7w3whIpkcyBPt5b7bXGhNWv9NMe+x
+go4UFMBEGNLFmOURYi5XzVuwJByOAan5M7Em5P8oxqGsMfJMGKVPN3HTuBtjIn+
HIdnGdM1hWKScrw5gLZZ5sQt/DnbF5yllP0Qz0zeHtAz2E9ImVT855ZZLttg6TvQ
BhMh0c8eYP8PN+dTC14ZJWLIl3YmaGyh5MC+pJ5sxqNzAD/5BQHUZEznJTGQZmnq
8U0ONHVSdPf/asKts7q/Nt5LxEO3S07iartTRlJnkVBfenoxYRSVce/n0T+R3kEm
Zt0dmyYCu/lRa+CpMkORd3i+4hCZF2WtdHUz2R9B8ca89dAYGly3mSrbdYjQFUKG
cQfmjyNVACCry/xX07krTLjvoc+QW/58YxhyFvXcX97kddSkSMIvC+M3yT04zNrh
rQ6aF0VTdmXHyuYHF3lmwC5tsFu4PPoQgUozUTnPgf8zkt9Y+xVa5Dq/UWwxrbAl
BSHqGoIFeF5lWN2l+wKM5LzarMfzUznxwO9bqPsSxtvpHfaUv1p3Y02EoZAZtTUv
Aa66aEPulYAbKu76OuR/+fJfMF8eZwr5nxV/HPTAqanExztkyz7W/rJa7W9pNjKb
7wzSyfug1iG34m81+ivJ8Rdn9fOswyf6xGcCWX9+9lNCFjFkmOVXF338nZUdomea
tNRuuy5c7mOveeuokhZVDZ3q25FW/DG5t1cVkydtusFAUx+uosZwGT1N0zpK70Is
qf0erAPe9BgBzHmoOfD1RVywL1zynDYnbXv/Sxz/5w9xIWJQajtSyllKhxfm92Qe
RzNF1vtLQKl09FffTUKzHfW5UT/fmzPAiEZqYocOamMueAkf1h4NawfedCH25WGE
`protect END_PROTECTED
