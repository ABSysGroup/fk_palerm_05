`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
veCW79g7gWy5GM3eYGWCSVHlMz+3Ak6kEEHlrwfkMzG1hZ9R7db2NTtc0RbwV6/n
YaFqf4HAgigqWFqvC4/3OwjoE94DRyiNoKFOiOEyH1XfHCvIcG8OaF2VRhwpwiV6
Ro31xhvFd1fbFjnWajfYyruQdHoOTxwp+rkzI2QMdQqEcGY3ow6DFsdqJo8wJGIh
2Qofs7pkpagTaaa//uzekHkG9VTx/4IP8L34jOGhj5kKr02XjJJDEBgWd3hrbYPw
g2hEk0XK9uz8jWHu1lnbzrDQkOucCCBjWn7nxrSfraJ/JOadA6+1DrUaHOQB3zJ1
Py09NgWw43P4ppixX+5Hxw==
`protect END_PROTECTED
