`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Xm/myrW5QGTCw8G+/B7PUIJXfCyiTqwdStmpVqnd7UPPwW3vS9Lb9FaShTiOWVT
F95WrVHiXnmVcn6mOY4Zjqn/I68Q8bIh7RrzSIMswLa1u38sydgS3tWA454/TnW1
Bkpn1pKwwdnION1D7kwtOOBkw4AMGKnhBD0aI3trZrs4RRYiwc5nTwwZEp3CowJ6
wo/uIfuhgZUo4qPu9Pa0g2drcI5hffwUJ9eVMFqxAQJb5CJLQnaIRyIUSVsukmqE
SULY0DDAY7v63UHSActp5buVcAGKag5MDYAnNKHNzwCSS2iW+f07F3uddt5vs0oA
ttDxYpVXn7Sy91Z/wGKN/5YpI5ZY3OPnXIKdSfA6THmGzvK2LDdn5rDL/Iz0rB+D
U+U/Rj6tlVONjiiJEXLl7hAEiinrjDk3PxnGxUye3zjccdQ/SEXb1tLZ+0H6ZdVV
dXokJD2lfeu8TZkkwwOOqp44dyxuvKVlC+HPAE+tvQH3eCggp7Y1wcFlvEaieE3w
sWjYGjxO+AoEs6RbPIMHYlAXJtCX1iw45goxblXV5f0+OXQWlKmaVxITefIYwLh0
D0QJJXntcq+yqphPVdBwBSwGtxEUhgtdK6yGfLNqIaWUd7fV3B++g8sWQRWc5Goy
w3HqzZ38aL7Uq5C68DINK6IEQOUUcgUTOcR1I3QlhrBlUZPqCOg+gDyunWsIJrn8
n0otFVFsCZc49lIxZBDBQtKhA7KzmZHdRyTdpdOQFHjv7hu8IoWyzSgy+ZFTY4iL
x+cfEhvmUBoMRBB8ArxUtl81uBZXS9fAqw1A7hvUIzRyDgdIgzhGWDmCu2//DO1M
a8Qhj/ktfv1RkvoFb12+VvW5MbWnJHI61vQINPK0YIOfhaYwEIu/D2VHo0kj5hNO
j0z3PKjLvVXdq2BOUEezgyfqRaExaV9a0wkHcKVPicN+6ZQAJCqnw5I9cCfRInh2
KJurR8aiHigQHv4vUCYFX3jjppjCaF2F6A3oPuypKL6FQ701yL9IAYc6b4t6s7yp
xQnjVIpVHSerHYkiLiyCkOf5tgfp6+5Eu2gJaiR9txzoTmEEZMxtyIklUQ8PIymQ
hdd+XdBIEJTKW70hRY7bWy8/l1u5YEtfc4KrVxmagrgsAEFnoqXf2B5wInCUFPb6
9kEUNYuHrX+acHsBrAckCuvo40+ZZikJxBDQ9yY6rmrFaESFQzOce/ywKdt5Gsf6
5Qyin7N1aPl942ii4nUiu2BESmDe9ijhDIv6xR8Qqw3GVIVWfjw+qPWsHDb0ZhHB
/wnOOKbf66Qg4UNtR9L6hiFEFDszBqCcY2lLtX59YBjthsTQN6LU3cCMaQf137ij
yvlwx1OtRZqohWmuiZvy2BtXhzFngyv9DXHiNBz/u9NGVdtXqgOAmCZ2Xy1Mvm9F
KJVf7FS81nrk4FcH1fE9BqWu66QDwrIqkNzvhONqsm9dwrj272XTRWeYE77N8xQC
ncPtw9wpljr/zyXyeCEgV4rSb8HQip0kzmE16N60c9OPNqrDycwe0Bukv0LKNaSJ
+hDHGwkM2aA/qmUPCovcFF9dTVUQbGmN/cqFXSf95fgWG/PhWFCzOR5oKtXhU0qC
3jylJSF4IJkAL5Ko/7Gp8TJGvEKdjuwb9vJRkqI/bfvW3Q3zb90BiwMturkZnNyb
lTjlkWJ1zjFEIq33+JlLJLMVDfbA65ri7maVoZDlWIpdOIguU2jE+Ty5HzZeAAmb
z6wojH+VlB6z035Rqp205U19XhXn0wSiS+DGY1Lnp8z0aElyRyKvebhsl6ZeK3cZ
`protect END_PROTECTED
