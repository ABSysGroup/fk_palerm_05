`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ju5O9CoidQJmzKTdzJfeWNOQtkCFUIbN8oMWWyzI/8w/21CQZRJJmH4Es4T5+6PP
5mBePd/tlVwDGRQfh2A8McVHvI66CB/2c2At6zSr3cmOMxUUMi+XY6S+4SAV0YmI
qkMtMY8Na/rBM8jfVkRPStBrCp2C5l6RgWhXcUmfvFL7HBjJ0xd9qfAy36Ug+UJE
0W19JSivVT05MKw/TNkmpyqZ6FTvwLhZg5ce8ShIefe+MZTiE4FcbC1QTn67FVc4
KTCysfEFG27USXvNDjpQb2/duTwOHp5eIolKSdPvxT7jwGZ99s6+BcJI1Hjn6v6U
3m4hy8STd7SUNc0cXy3dpovJZA0IfTHHA4bYYitjzF5dgQrgy3Cy94VbIoPdYnO0
E+0MyMVFnFqdeEL3tuVnBzGqKzlgkQ13AW5Szm5oLDPQEc8fshtsVlPLm8rAZQwQ
T7Jh5rTQXjcKYUL23zScmHcJHg4dudbHztKFEtYNFazhXZnvfKA6oQvw2zXJlynM
95sWnBo/AL8SmjYpDsF4Ejzjnp1LSweraHoPsYl1s4CJcS2jzTwLsQlmD0SH0KgK
R1UzX5vwGhNH0PySeN9uk9QWONNLLmiVUhzdB5dH20n703n+f1FPAxbBUsPMUKXO
2n5lNLBBfBeAZNjkYiLFoChbSbkOOzocY+ioycKC9lIJpkjrxIASWEGHQ4gBN44u
BqllGZfYvRq/jNT9FxLP5kmoSIR7yaC3bl0sScmxpPnx6HPYG0jiY7a/uOAFshiM
cNCRjBOK5Yl8kINVeP4HuYvWCjLwFn9dDcozYa1AophuvtDJO3LwsAIas9/A0r09
ndaR26cIsirPUw/K32aRW7sbEz3+2HpHyN6LP5qJY2ZVVk6R4yepoTIbzIUloo+a
S/Bz7dWeWYdiH4rw/kbBITAWHMoVwNhgV8uCFWP2jTKoSVo4/Boo++vaX3feUSoZ
ub7M1S6dgOFMni5iplKiY6g9XUnpng+hX6oAbQkGxCJYrJPukY64tJ7Out1xYE8u
GqfyN8CdbByIzxWgWZ3e8zljbGZgeeHFTQFhvjTlYk2STd5tUzrJ4wHf4KUxL9Wb
4Ojdqaa0tpJOM4nTFTgoXzFY3lOcYnaob/1DrUvwNDoO83yp40xLuOIgNGLOFew7
RMsXPSAnENBpf8n4roFNR8dedTUWMi3GiW3PjnwcHghGVCnFORfah3cvyQmgfwBa
jAqsvGC1Q+9rWEUfQJRZcfurIzAYUHdyHcHvN8d5gD0Y4BNyZSajQmfwf+Rfc4j/
0ANu41y4MePTOx3VPtq2MN3+8zkzFnlBWZULmuvSGluV8Q3GZod19u9oWhqvtwDB
/6wBipat30S3MARpVVbj9rssKp+sjmU67phVIrb5rXESLyUjs1Io8aToMwNtYxkf
fPuaxcSvsNpHYRx5W9q+rFzkLTUzEblQPq+gCw8qeUUTeQx8rpkf1AktfkZ3amqJ
orfWhkwm+AAZMP34fjr5E1YElrEutJFEy5mc6l1uojOCd3356h2NcZMaQtyA86DR
IjOAJ5be9xY8lJ+fJpJdG3LEBMDL6Yy/0tsvCGwfAu4B2zT8SKf8dp2xa1hMyZhU
6bdIVa31o8W9l/eY6RPCO6VZjzv4JKGoB+2q9RticGbpXQV1nZecnf82oLtHFdtB
XZVLZFOnS4gpvFdb/Iz8OoxbOy23dkJEtDzJqVXcmT7M6NzTgEDzkJmlGDjNEB6S
sAaSQRocuEsMJ7LnI1IwrufgFa1YX/0HPB4EummtWk3VjcZWuh1ND1DAOHtsU1Q5
DKr45Ki9fL5BCBC1HYrc2QDRNJ+LRCy2Qm9riRhEi9+RsmT3Vgt8EVxE3Dsq5OxH
1GKO1DZnNe1QaqnzlafMgYm/cZuHIAsWdJKsKL/gvi6p/x3KsamNEwOJjm1t4ZJ+
F4/Mdlzp26x115k+rfz8xl8KIG1XNmHexDK3niI4oc7WYiBnbBz4bAMeLC6vDGlm
MEufVBbcbVSsRefhThSDGZJ+kyH4tCzQfXwkL3Q8MtVzWniuCgf3P6HtrlWTi0sI
nbD7RlmD5pjvfBkm5RgEi8HQ114NR5dMCPV5Q9AtL4kGE+rrebbq+jdpLOOF18j+
wp22lsXhfEJK2jQvtKIc8KtuZ8hFOh+wTvcs+pABoys1xaJNhak6ERwqa87WXlzW
FNNtZXRu+2VsrnPy74aKx3IHCtpvhxfGI5aGjGCCFUXd1FbGdSMwWAO1Dh5P3soF
aiwm7NgQzt/n8Pj+vSimoprwqE/f4C2gUplAetRCzP99NOpeedVrbTEUNot+dBXc
CE/P4O5txYo/H0XPjVdWPu7bDoTzNE88YQy7IuB4rfAtZu72mDQE4FAKxaRCS4K1
vq7CMTpL1zqZbxF0d8cBexGCWYPDcF5NHsJOvDJlCxPimzEtCYJ+54n6vQmgFbja
gj6boUL1knK4qVg1PkKCkZNcIGNx+saxLs5AdiPU4sVRA4soDW4qUgjXQvUpyVhv
LMZhMFeQ7eBeP0imW1SIS8TLW/A221+bErXQC5kvu6jmns52m8uXpt+BkZp3dUz4
8Ih0NM/tumvbUdTAxvvNBgOdYKoDnNYsxkGxG3HJe9K7QGPGMe9v65iVueJaUK6/
1ceXdodN0eMK37VD2E+hdqTPSG36K2bOXrErG+1Ah5I0RMHvKw4YoqqaRCek1ZwZ
XYSqpWtOKA/XlvvNG2tuQp/N//hUGB/eMMtYw8WQv8ZqPxYbqQyXkI1qeIh/wrIq
ENmmQXIZ4I76oDtnidN6+g/AMT8dBPbDCzoi260ScvFpuyji5t3VaArA1/Puc3Wy
q2E8lBP8PuOrzOTX7uSyocthRjulJsH6nylFuL9zfZyJ3leP/zlj6b1RVXfdHKjS
aEbZYshBWC1BlPygh7aVKyQgEPH5Aj1P69I5MQU+PVttqiBps3IqxNE2hJgguCSB
iGesWiRhaLKXvk7xlkQQ84++KCqDM+M30eE6CMu30xoJFP4klwXzidIiQbLSwRag
Ktx9mNyLKtoeBT5q1creaJqKU98NLCNas2wC0H204ediOo/Qtjt4FxrFmaEP+xnh
C7ze0eRybT4pYce6l6yns0YQ+lt9vRnEhe3WN6jWUNUtZqSR1ZvZyVn9rMmjsMs2
hsRRDFk6jmh9F5nV4QS1NXN4F5WPEfocHmlPgz7C0q4fA586Cud0guHHjoogqwz6
RG5bVbwiw6IAGHuXfLep0+pxgfE3Z0P5jv1CdvtazdzOJDewHOEKJZSnYK2DFhQ2
6DDFusUE0GdJ/xk2Boua1yyq/Uk0pNJe3FbWmn4nQDlGoNLKGPr6AeAq6mL9m9mR
8pLs6C3n27AaALleAV70PcEtRWC2YPluLHnMhxywODn6KcTkh+uRTd63ZgFKP38X
d63G2CdEQ4PyHiXfH52LswTsOu3rCq+Zd6zgFDM2oWS+izYUVd6Ov3MMxcH9l1kU
FVpcVJWRoDpqADcUwde4sSd6n4fI5YldNj4ihSI9/qq1PjGS5ODwP0nbUWrHSgKK
5GbPhqSQFTyacwceGGLyPTcEJm7dDel0aQmXRsiqPxcAt2xCE7IUgyjoV5VkbV1w
+v4OAzETUEMNtVsOfgMltS6WmeXvecaxvgaqTx+SGDtnrpBjQuNVINpUXFaI6u+G
bK0TsbIM5zwb3SiFTCurxk7ZoDaFpSPH0jFkkctE0NtZKl3HPCC+t9VUz145hrcr
duSdtXVy+7A3vv1Wr0CYRpVHfs7CIS+/0SEViGunhKuUHY3cip+KSwQONWKLvHw1
Ij4fXqg9qb4eFhqHwa+eTe1uzrxvzgJE42O1Mm86Vz0xk4SQt4nH5vo+PRU6tKx5
nMLkGeZlIAVfFTkl2qR0AGQzKbSTnKq7jWgJilWKUBuipB3rHESuS5qWR0Emrtvs
LF4y9cNx1L/sBd0XAosUAwdWsE5zL6a7/O+N6XbqiZ50gX9oXS5sQzxeYABgc1IP
4lJWLlaBvLYtYkISsTYoc29u1z3Jfi1T6lAyh1pKDwgW34JmkE79NN8xN03oYaON
4FJUcLHvgT7qm6wbSvrbz5vKvAgvYqwBWwQeZ27tma8/91WcMCBlHm/HuNcrYxEv
xtkdGg7l9zNLVYDleix0REkrbyB5O3vwo4+ytIWJWVHVbPhCmmA4wsi9OTnm0KQZ
fSLruYLEhyKN7Alt3ctC4QkQBPrJUwakqzNxIGZnFTGPrHX6yd4rm7CJwtDC6tQ4
UuyFoOz5S5CKwII5g5Hg/Rqzg5yRsRWWSgEGrHgr2Cs+6f+2GilPzDV908qEbKZF
znkKZhzUmimPlge5cQ9SLeGcCTFtSdD3sF+3EXNNRxJjofliBOsmrXkuVF3omj1t
LG2JNZq4OgJywfEO9u2nL9t2xx/7sFye/GQWWkBXPG0f4TAxB121B7NsgJQwmmfC
dQYor5yfT08pa23Bqi7OYCJaI9eLgQZq4V68pwIdyrfc+6gk5oZ0cBrF3wywoKhV
lTLrh3TzaVhypoHT9jhCJ0bRwEIs7h5NapEj1OUldMD98+dce/JNqntCauE8l4s7
ZtAjFjheFMH/17Go6lXQTTllaED6XY7o1+FRNVp+d3trr4PS3h57c8aysASXJia1
NdBWP+GJDJhpUzn/Gj+mkQpaSHuBiDjgyZgcE6HICeFljbVRGCyXKpXYddJ4a1mb
nLP37x0+4GpJ2bMAti2xtxRufuARgkU3dXNFLVlH79ENb2MIQn5Kb6x0PtogREgU
acuYNGERpckE88acICcKLfueH3XB76vZXuXtfQdTpO4+LTV+K/DfH+Sa7FG38sNk
N6mJCJSTfSmnWHZQKhwZwbReQXcoOu703u87kWs2HMHzJq4AieHsiVRfONrtyfyi
45DEpZJyA8RQVSSzPExQEKlQOUwE5Fc52rllnNCubh2Zv9lbSF8f1ZHYz1MAXmq4
y/q4IqB18EuW+pR87mFPYATS6mq7sx5uTxXXJe+ynYlJzyP+UbJLA0mU/1NxmiYy
W0Rod5X6BKdzgkroN8jAg0UZRHD6KS4UEwa7RHShpJpS7+9hjcfl5c+e+lMCLre4
18Qy9p/Rkg1TouqSDs652c487nnGUqIQkZerdNId57uLFri6EydMvd9dELROGFR1
MSTKb6rkP8dtBFa042LCEUT7o4gaJF5rZt9TY3fAfohQU+vTwmwglo4eX1mHKNj7
rym9R6OLRXBqu9ngalvCKdSbjwIDzxM0cJIB55t1/urjulFxqYvEbURUVWlnh762
xS+QRfIF7q/B7HSvmoaTCPCPnHLTtc4njXgfu+yh6sTxAg07FzSZnbsrYKz6qvib
se372d3PyNerztS/h7V6UIXTouQleb8BQxqZp6pzjKNuXc0j+TlmvBej/Q7xkMH3
kPfMrgRX0UpU0t2PVe2TIDt7baWTGytfTQeyfxopqqyqR71Lya6TNSABzn+xkprM
OFWbTseo7do2/x7yWFjZrt5Kr/23pTmGxDA7L2liblWeoHs9W0/UHsgufHnEk9wB
QbCWZ9rRSMCZLEqRNaLi3GlLKvCU5P9kNcWU0C/vgGiirdEYUQR+4EsCXrGOz7XS
llJdctSf1u7MmTnBAF9gLOBMmBe2Ukh+Mtp0JbmYGXPpPs0y5YYVRRASUadNo6GU
ZY+tubjpNx3GK2Qi/dEib+vvKd12ow2xkvLqJwrgM6Cl9fsredy7BIrV//AMF/lQ
ua1ri679cvLWsO8nGJwr+jhKQhoQetpx5BcEyNDFmQXnYXFs0iqONXim1Sg8Rzud
OUxJooo/14VjN+5tU3Ycl7V+TAlJm71xzdwjVkGch4Egl21Kl64VjVXWhuJfQQGl
/M2T/NfHxbA3zPlfTvryjw7u/mHk6/DaIXznbqLw9B9OfuURVscgF3ih04ZJoR4x
tgJXXlSy+jTophqBoGG/My6lPPjB/BqI39mzU6bjGfaB417ylX55d7eMf6Q45Z1D
dCWrZkgcLXc5L9TYkAgFFnjOkuiaAFrYxMgvahY7cbkLbfCeMd0fvO4QdVeKqZEQ
0BS2O/CN7uRjyVhAxF2FirCKyUcFMuYo96jm8c3egZggLxiXDINrDlDrQy0vBQ+T
Fa3KtlCmBeqTUckt9UaDL2FXK/90F3CjLeP3thypxPoMLjMH46G4eeS03xrKNgse
11tUGRTOQHKl8F2ks/pJPgdvrYh103t8kqN+hV22iF+yS9gloZO0YN/9aLGyG+cb
ezsNF2Dx8dmgLsG/WvsKCZaVNgbgmKAARXtcqqq0SCT3iYsdpmZuC1nDq5DuM55j
eOQIT2HPyzpZ8wd7MTnwgN5pk4bPDBEYU6ynEVGN/yhdklptUlNoUwzt3zruREyv
lCpt94dLlXKxIvWVklPsfOkx1+T7cVFwl4Q2S+hJ9rMZKo6O/FG5Ae0bZCt98f68
2Wz/uMb+th84GejtwNx52dmUMVDffxQkg+u00SPC9QDz4qOWOjCMbrPiZPlEEltD
cLfdaORYH41mx49gg0VBeNUIcaurT6v6WMOvsSE2y0Y9NuwRX/4QWvDaExXL7FDr
EiQDHuFst70aA697nXgTroWatJvreiA0YkkJHiTmr+V6oZ7M8uDiO4mADAuitCWj
g/v93JG1l1HGPW2SwCQbg3rdGHOhSA6YP9QlQCUpLUG5hkqAg8Wpbg8Q0Lzutolv
grpbTNLrLr5yAxXoiOXP43rADwKLHnfwlugLZFzYVPfXJmN61JGkGyZUdyGVWAWc
eNeL7rrj7y2v2+bBoU+U3kRugMywsPWsyAEYcQJJRbZ5fsnhlst2z/lnnroo7gjs
pdtEDZmxgWHyZravxdza8+nUTgPxjWcaX169sUZg43aBumOjHXfEZWw9zmdvWuW7
I2nYgoulNTJju/3XHZ1xGDoQ/QWssrl5MZuVcyxbj3xetTSHP1OXe8MbbqVDaJwW
GJuF9fP/cWbm+GQEwFzK5RYbp5oY/Yy6FWhsUUkbhxZLBHS4WMb7RfYs4W5zWet6
N/G0PFpeP8M1l3M9o74gMZJiSz9sNA4r+8qDT1mQr5LUOYhn4FkJs3A/QIQfDgPL
VNF6CNjScVlz8GzVTzvFS48BRV3E+sPwB41FVPOnDfJEPaoi3gjG3i2Wd5qMHS20
4mstD/VI6dXjazSP+AwKz8VJJWrRu33/XaDVwPFbGC9/8s+mhHGJRJDgClumoZFG
NB7uk3+29EP+46+vf28ApQXAEsyuEXO4PgdzOy38/RKJUNldRBegaZ01yZPS6FLk
+r3Fj3gcgjjmzzy9uPLTnFcRdOdWBwlTjrww1UwnvOond7xRl9bnTUdQBkgsBKSJ
AJxaLfijxHqz8JRwsPmWJQY+bsq1Hs5Zm3Kfx4YMbmo8CiVVVM2V5gVJmT5WLQlJ
EceCv/9hXx1EF6ymK5FMESNqEGxMfMQi9SN4wV9W/EefCyrKD++XsTZIhUVLsusu
FgCc/bC9+Fxb6wod6NAVYlDKDYtGO00S2YEfkLqclFwv2aiktvPp9G5wnLel3Y/X
8OihPLIG5fXCbJ+F3exCABKHCbErj9B0Y1XzBuXrCemO/1rkaXH0rtoQTfeIT/et
S5irSEL5A7BM9zvjnT5D5l2LUN4+rbroyidK0+WaRVsPWA+Y81OR+6Kol9AhDtc9
EKayFAk1qXm+pIp+Dz4dMt/Wok83Irey70sqJwXLAJUwzI135aoaNJL0yoqA7tRa
7Zrr4kqk65s7oKeviF5e2+iCTUBDEsLYK6A0yUyxV53VX1v1Wyms6GZaHcKwouxg
zdrr9MnJyctLvbMCBupqTm2mgkEn+OzwI7RpWKCSBVJFbtjrpWAt/NV8L7awtOqs
GomObaG9qWe19vm63C/3btykMb0pHUYsaSyyBltkfWkxkcUd/1JXa9aCdLEqlH4/
cTRh9GyuVcGFUjPzeVEhqHp5NPDc8+Nw5NPapi+Q/AibAw+JZ/lq8i0SOLzagSmz
gTp0Cd6o0nWRfaRiXeM9Dn72Uh6Hiizss8zozOIPa9VsBECxhPEdmNaX0Acf7dfE
IkIfMsiLBg3zbF7G3MQ12jRRasAika+PyIQ66WoBI6KN0Zn020b49io0iVq1mFJS
PqxMw86s3p5vs0IEhEk/90AM5iwfm2/oPJVltvpZuMJ3q/qGaAGZo0w3RfiBr4MX
S3DbsijTjBa5LFKH9JmxhNwwS1HbWpl92cvfdiNYEH+BoTlNeJQlJwqR80lJc6mt
uqkXa+04oHVH6ILmwkHD29zAFH5UTKtvOruBGbugRyYkFqdMWf36OqAXKAgCNkTS
+Ic8j+mf7KRQfNCchq9Iz+EWSE2mMnawtV1jYIO8P5DB17p45yuAPOJNZ+l40X5K
rwUHehwlLbJ75+aVI/ansfzsYSuDRYOoLAEkxRaonwtwWZk0X93ZkJqJTKrktZWl
AImiYk2zgahejXLONhda1Ovyn9cwDBbDB+qvSDtZrlwytMa/1q1G6bt5FSy7BDRG
pVDpyc+F75pOR12o8udQfVmUswrATOwNuwQv2FAoxUftwt2WCXYVe93nYZ/7H1zk
d2oQpCwUdCsEXQedjUwuGGvGIcdh2MtCAg8oXJSTWmyNicn0QwC3jbsXV6J6Nnhc
EdynNEzKR8tHBlM+lJQq8rloRJPPsa3K5X6GhNYUhue04HYnfDUsnS8jfLC06O9J
d76DFKEv1qrvkk2dtF2nJh97nkAXqnmcvUqCIZulR/DfeHekoOlCnmQ9bT5ipeLx
LW1875QM1wPuBhTZr+UOe63TVxUDFRoOsWTy01ia/MgeADrB3h2053m1e4JFflE5
jRd927o3yQ8iUj9c2kp1faM7SU099C0WMhErN1d+Qxgq/4L5GCFUd7hxlEJ3SVfn
sQc19E1Z9TIV54E1UTzTtE5PxgrqqIXN56cPL0xgtnH9IuMtnYX0orK7TiEeD0f+
CL7MR+d/XK/SSNDJRIEuVw6yNz8Pu8N/N4T4aihmlcwxuy91DAgyD+3wHTJwdgzh
WLzYhrwlE6Fdcl7WNt4GqHGbSmRyM9MZzvJ2tYocY3bPrFP7rFRFSe0tmbSdHQ0b
8VJOg1zpSfK4t0misgZvBzi4slXYQe6LPzxOvHJW8Rt3qfT0WkCJWOpGr28k+0H0
6UYJ6QLM1Lwtv2xhxB0N8dSkZBkESmHn3mKEeXd0eqOyL31M6nP+GqhLSss4WiaO
k5utFdv3sjgytBohJFeeHLQhdLkFJ1wjRRJKTKk7A1XCDjAJpxkZHV6xY3KJeU4T
D3SyoozuAbKvfoLe7tXQJmhSpElIbA3lZszK2QWij1fA9V7dO0f/JJCLBpW2xb/w
CVAHwmVp8stVN+lhN9fMEA5QIZk/lZLyuljqkgPic3hXaqxLY9mCHzIi7un2NVcC
a3kaJDrWgYYCNWIH2L331A==
`protect END_PROTECTED
