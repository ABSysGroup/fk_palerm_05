`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DJYUwujLL3M9N+NMtlaCS0Jng41VqAz6uqZXyTibdnZhUojRBx4C19AnhYAFisVC
vyjFUDfyiuo6B0J3XUdWnq1tl6EKHeQGhHs5ZN2ZkYnrGJtcJNwWf9IxsFh+/F+1
XWQe00oGs5eqkFV9dNfuiFN6+Q/Sl4d45leLcRZEL6pTnah4UGVTSbZG3UIjDmve
Ofa0OqafqE95+eBYVwuVd7xUYrqgt0idrTpeYnEnhDz0wNpyAL4qcB0cQ8V9Oj3i
2hmCZ9hrOLOnjuaVmuwqQRrdoXZX9ryFM7NaKptr2pOFuKGSCI4snAwfwoQcDy51
J2VaVOMjTcHeS5dX3iJ9u/qnc4dEiaSqZsMZ5uIpz7LqGECSaDPYy2FxlMFlIZ+p
cv1ifb3Mj8UYCvZO0bIVIz6xbsZmZVPiRxhSJuL2QNRMJx/vC1oC6Z61WkiswNYg
kdj9+SFuVUejJrgl0NNzg+9sJtrT1TvWNXVdR2Ht4hfXeC/UFwhR6ugSSlu1viZm
svPHr2A6MJPnvgt94EZ09nfCRdR/Va3XZk4Usc9hqeGflDqh1zg0CtoxRB3wt3Q1
nBHBQE46qTnDwYmdAM3coTdvbVyBTykf6F28uPT+ChJ5BW45jWf69mOm+ZoyXcG/
l3CMBS9lOcZLCbljJXlBUgc0kZu/3LCzATDee8JF8AcL7Ea395dL++JFU7vYO9Rt
+M8iJyXcbAJx/BjSw+4XOwqq0jCib/SC7xigZaraf4i+ws+FYHyCQTAHCx/wwHAi
P3IobkqXWJ14B3N+TSOU7pYe6atRyVkdnZa7pZE0ulUQ5JLPJkOl3y11099D21Tx
syaxuFG/W0QKYiRGNXLzFAFjxjrO3bEYZbYzFp1WUglT0agEJX2fBT7HwIcXjHL1
FrrL+hGilpsZUPIbz2MeKBmD6H6MGzwLTQUJx9PGEXLKB4Un2pf4jVJCNdZdcoHj
uLvO/UfBNQnujqqPoONwjAAnH+U47PWq613o+nnWOrPu0tNgjB93ftUYnsP+Q5td
T685X7zd4lYTAV4seFltL9kJYGTHXBPi7Ge9usZ5iR+G04ZjXNOtwctnyVTmfGSA
7LLwZDQbZqgfaXPPGXlHXo8R+MG6qVE4ekVzZRlIF6g+5PvA/9VFrKnJinAXFMjU
MRFb09LbwxtlnalNNQvCj3Aj9rIiSqzlkHXbAUGa8Ex7QY+Lr6Fl581z5ylGw4Gl
3BnFoYID86PWpPBuIrD1/bOzg7ruVS2ktL41BG/Nml6/88RmNnv4eiP2HcgZ2lwQ
6t9ss6WQ85U/mK1s8xz8qo50eLKx4/uPuQx3R6mnR5zUSaILIGvd5OhGypAmad13
hQnWM/49mqDveZmHmc2+wV6XCezBiIDeMU6CB37/hcd1xl8Mh9HB0ioVQ1lGfRgo
AVEB5E14ETJXyRmwr5tty06xOKz1jsnUJuDVrPdXMjF0dXJEfSL7HP9gAKcvBNj1
GF6qOND4nRyuNsz57Qpo3z8fP3ya091NJSmnw0ZsKpt0qG/XP3GEyG02IFJDL8CR
vLI8IrHLaDYU7A0oi3OoyCuxLqvUNJ3tCGnqb9nb5ro0M9V/dpeG58b+qJ+b3rs4
u77/d6mzNbZnmUB9U0HZplzUXRjrnDgshTPSDNNDY8GGvXu8/dIrn5GmGgmESQQU
76nyy2Pu+UZPEDtLyBR5Nk28bZmmUF6KUSIY7yXerImCmlBw1ITIghgxtHB3w8mL
qfwdA4lMPsQ2lixe/1JrvJUNS/IztKUxUhTQ4qcOwhbMxbrymCt0ftlSfM8hn972
jfGbP6Pobi9GSVnQKwRkFhjt/66VHN5y/V5Rwe81Im8lw7oHgcwzC3+/GhMJPH7p
PRJF6uFMV9jMX54gAF0gdeFO0adZPQvqSH5yxOqP+mmZ7fF92LFfJNXQOThHg+p2
xRcdGBV6bKxF4y9O0I6fyTeKzdnk/QG8jDlTJ+rv+vql6C3UrYKMURpiXggByqAR
o5rYJR8qkoHpcP6qUUfiK6WG+4Hkc7HeCcbgg9pqeMcjEsemof7C3To3ZH5O7x+B
GVpFnhMqf9eeqxPIeKCG9NPub9pjpAk4mqtYCAl8AmwffuZ0TDkFoWEmFE3G5IeN
qhOHG7ycKguB0TlZP6S/pz/B3VhXUswi/4O0W4K0HzAlRsbv5YfaXcIBuz8vnQgL
sZJ04A/WlLCGS0Lq7Fr720XhitLB1eNslAA+ZfAcVjjJMm1aT0z4lcWm4m9+dEhv
+PRqPKKp94qVCBjYmGiaewWduRHOvDFCbC3gGvJC98K0QgXRjzj0EWpuw4lgSGWm
kb5jxmDOhk8O93Wztb8PUc4eb9ULl4YIlkYlHAqxVLKlIgpg3/eMXgXSJGqQaVJR
vp0d0j1GSO8poZq9RZTtR7MjE/v/lATO7NFYLDZilO0koZ7R4R1MCimd0iLTqUUm
UR59g4QDGwV92OFymlgx1jZVvvIbZ95k0v34MeylnnR5In8+t7z5MHzaT3hX0BS3
vsfaJBxCAY4Kx3do4F2KdCGXFXnq/Sg3ht9Ee2EeHR9C3tOcWUyIHltCKong5aeR
p/LfNit0wTjid3xyQpwccXCx6XHkAuCzckOO5Nql0x8sOaDCAzCgA9+Ma52W/bzu
5zxzQ8hGlRq7I9/JYK5nH+Q+VmyTGxXzuHEilcXH2hhl40NPbAufKuQrgrgsdqTs
iZK0tfy8fgtD9CJaT6YF+pz9gwP4xdV3n/2oSly/QlNKgtXQfzFTar2BBWEAyFqu
Zp99XOo9fGtqFfttI7MDsday9Qv0Yaxpte8A6RRdUKx8/dazVWigs8PEIWPGyyyP
uZP4mKFVjHwwdYvg2YoxOFvx+qNZOK2JIwBa1c4yU+SjwsIUWgiKgYhC1rlQdCMD
FUP7Klh4ZsLjQmmLRI8oHsnXKhFgpWg+UNQMWtJ6EwYAPIe6MXuztAH1XRON4lrj
Z1ZMM1GbvglrxPpugZ5F1oThNvXV93fF4PVNK1jrvaPDAUBA4OpdNaJv2viOoDyG
Ez8fGkJiOMQDPjBBFtFL81BbaIEarz1XVjG+0NGafVoernBYfocdcTtETKJlQ4vX
nnNiGo4yGCSatpKRNd7fmMlWZVjplJHtxUea8drO8Rlhba2pxJd/VLBYBxbb4eHW
EbnDXGqYJUqr4rRyjdGNn/5jaBNyNNqx/bfDoQFt1spuqCH8HEa2H54I+P5dKYlq
tHT6C1SgGDFXoqBiOOlTw+ZJrmoTJ75pFx4uNATh8KZSZ4bMEGv2d2JVX3f5WWv9
n7j4ib8iYx4vy4mBuENoV+5z4zwBsA5Z1+4rBKNTHLbGnGMV4R7FFuXoGB7o18Pb
J7Eudxb4VPwmRJyQTwVbMe5L7oYYaiuLScpT52oxHZVLWH4xiH70Cqc/r4Ln324Z
5x0wl3gWOuR86126GdWZ7vwjLsj89zJbMwbLDTUlp5Q7Zyzf+SyQUZlR4NLoEQy4
XsqHfpzTn10pxzG8h4RbiQeZ/Gkx1FEAGOI8KUHusxWsOluNMxBVH2gpaMJ4uKxO
T2HbHT5B9Rue++xEh20xyaTl49g4wVZJVdthqm4z3nfbj9GsUxjMvGxGwSam1Ta4
y+DjRPvd9ArIE78E0MKeTtfNCGNZbCiRI/7YvET9NyC/VJBEt9H9DLWWMsozEOZk
Bh3XLeaxqk2BHUZN3ZgFgkYUq93CX0T6CB4ApGeGuWFJqqSyclhiwFKgpWS8AyxP
rPDfeu+UjMq+aioEr0PPcEp5GS4VXgTlRbqA0GzTja8yDq/HCLNOdVRzAsK13/yY
r5A1gVIM1e7k5SZhYTeCA325QerzTmtlvPwChqa6WKRJSz4kfOqjk6mHIim9K3Kw
Q5zqablPoXHGD0v1qFSwtQ==
`protect END_PROTECTED
