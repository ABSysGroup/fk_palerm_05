`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sl/hOkwV9WLsCydXPqVvUhO345Vsj+0FruMzQTF8bmkmRj+tWItJ9qY65bbNMmAe
TagORScpTDcmENiSwGuM+9n/PWwhPh2Suh8VYuwC0JTPLKBLRqmWnHvFGjxlo5bJ
/7OoQh29VXbRKva66wIrXvIk9yUE0pkkUTxFc1pK0JGDPojcTe9dJUW5Hs1xegbE
EHOPpqn+OKYXSRK0UFNYhW6h2cH/mMOgh0wxHeTr1AyEAAlQ44tgc6EuMDO/IhV/
Uiji1zu830RTBlhsDZwOud7647vbE+vsSwl/LSovAvVChSsKQ5r4hwRfvL8RcxG+
ZEjLtlBpcavtQGG9PzdnQ04Oyt6vjOH4orAuj2jLMM21URkf5MUJ72XRNE13UJyk
qFEayrz5KAOh3XL+pW4bXRIFQ4Z5Y3Ovjt6FknhH+wNhNs0tLhd+Q6FPDdOQThMR
w0XM2v0Br4YKsvRojuH0JfmeP2pJ8Tvbl5w71TAILWV1ne7EOE/EqOsA42TEAmRw
BoUrQSCuS+sE1p8rgO2OrlHE7PyIfYJMdS87zWXMbzsAV1Tdj62yc2dj72+4qkMx
KuHyWWpsMxwv655FiwZMVg+zVYmRDRSmUIBTv8S+9HpW8NLhdbV47zYmd63zZ5Lm
q/5EKQru58Oiwy0KI8Kh3OCiJ7sBHUs/0gWle6zDmQesjm3KXsByqr9iGSuBdToV
QdQjF0hoduJobfq2NRqXNWku3XBG51dg3GYtLiQTGzOhacaMIvMsKReIB60i+kLb
zPK+YpAG7oT+yjIOmNJX/B1AYuisCDjNZGwEe6qR1qShdR2GjtNSrQXj8wt96nPt
6i/mM6KnExKpErCKYtZVXVq+OLrtmg7bnwRN47zY32rHWP2VDWzyEihVGmhgBAWr
prU9oNeesKWmOhMkUmTEAC3BomZQbYPv5bqeV57RBmYvV4kXoErbbhhJCgk+7S0d
UOCiSlJQn5BGG42K6mHR9H/K4OcOS5T8BGW8j1Hidp0X/HMBPT4YsDkruOCuW+Mu
wji4eE4GFewZNelP1jGHFKAQGx55fGcWYN0HRRzOdbThhaTpV9wx7mq3TmLJTF5Y
r4V55DSD2F/tPdTgJvPekwDbYx2sSEu1hE4ybSPwUZHgOmuBf0AeWzpHdnZCkthg
GzWlUh9iQ4sUvwfZ6sE7haNfL/qUdud9uwGEzt0loX6F7hZQtHpj07RXGQsz9XJU
Qfi7mYhHuo8bG5Rk0HYx9RP/DiIq74BuPCyTxLQyCL7NaMnTkgB7S2/ymlicjGvw
P2Vr+Wicfmhib8vHGup2DZHynkFhzqjQ9fli2FVn7v4XLweyKkA+eqRPLZLpYmck
KaA5FJGiewyoTg16rIcjTknYdLy5SdlwImTFK6Q6rGX5h9yV/NhXH7f72sReEgdO
7IkuyOubjge3Sb+ZlfHAmPEG2rgIyG6xtemlzmWnwSK8zbZr+mAIfSkscFdbSXsJ
h3TdML5Yd82zSgd2Wxk7/yVaqr4E65ViL5e4lW1EE0HUMGGdS/Lifw2A/ObIhNJU
BiSrQgMgAgZtqjVJ/ADYWYvbEWJf0BhM/4zJJoxJVjFq1Bo8mpxmSnZtoPhvpIEN
hWL4fnVSZX+BvNXT5CteQfN/+ShpUgtpqsR1mLERHLrj9RLNRLlZcR+ohFXWxA8G
XuKm1ppKpiC78LMYTsr9AQlXwJxEymw4N5rYo+JMs5QY26ul3vFaZsTJ1YOKowZr
Yhdp2iG/EihVAdcHmoEtxQgnXQnz59T+kta/Mii1Icfejp3u4EwyxjJVcn5+ZUvR
bvx5HjhQuy+/v4D90hs5GwfNC22huOksgPciBFMRMUR0emXOj2wJeJqKe+3qeSvj
joC9AZ07HZrR4Q4tKZB6DQ==
`protect END_PROTECTED
