`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8uFfiBXi/1Wb1zjMGZC4sB1v84JB9+n7AzfdEUsNbs2gzei/EOCvosbWwBTI4tLW
oluVCjVfUXn3qGTpQ6j2/ijRn9ao13dstB/t0lurXGtZ3uYIg1qc94oXyehNC1Z4
6UgD4d7QKzW0A6YloE2OZ7UPgBi5TNfrgK9V/gpH31+S/bJuwZk+S6nZHYcAXGcj
onSopZCdvsko7re7GYomQWceHEe7ikFoztYk53qbKx7g88UHvh1emRXTgc3dcLIK
M76ZEyZ6L95g/rkrAAwhhqNFBdgornmi1GArAqXCKA9kc7JZJdIa7mBpJjrofr4v
JblBI1DB7/xy+91/d7hq5ZZRqRYH/Gs/AzRwAucNLvT8LtScngE5Ew4iPqPtk36Z
qxMfBxnnLJsZP/XKmjV8DipaA1H7FrcWu+h/IbRY0X4MdxBK5eqAY0jNAEa6ICbM
hLo8xD7xGIsVvqE4Fuk+KKlBTMHd7Hpw5Qf+6vM2G8UTzoh4VC9Bq7k9NVBK2mhQ
oJwmdjIhwSgrnHT/r86X3/NzuAX9ixO6azjQsEN4KDXPYskJ2dclXzxFQ4Fw1hQj
KlI/gFG3VKdGoD9AhTMIQzd+fxunRX4QIAD0BRsZKoIh5BxptGr0iMAbRP03XzTm
Js4stzuHvyELDqjHBghbVJynRqz48g+v1NxTAnLpVQbXaCb9VkNFdSO49UUkDxoX
hBuJs6xc4NuwQbASD2C9VBlKQ4L3pVruceQccXtYbuXIEVfcS857PKJLTbl5zWPD
WMfVLpIHsY8Ws2JIdoj7magK9xsEbroxPTtm4HkhMvv7sDR04o3JS/LV+QkDARhD
JVRBxzC9oPshS2b5SzMm0H90noEhupGcs8fBaXBrVnfi9NEL0/Ti8A9Vkx9HL8Je
6zGrDt9rzDGYMzcIumIuQZxuaJkwMmjWWPcpJRQWWJFlm4GSu3MVWnzAxdhzgKUp
`protect END_PROTECTED
