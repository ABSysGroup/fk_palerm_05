`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QKUyWJhqJOPKWN7s3DlcKteZS2ITX3SMTl93PHg88EEBxv/co9085c3StGxBOn5n
c3oxJ3h0jwuwf8wiyI48I8kWusjCEHMZmOdnUevA1XG4hZTLFY85kpLusVD6/nWR
6kO1O8lV789IWFmzorjBaevcY2U1q63WNaGoVO+YdFUMFCPdbQ+X2bORaIS+2lOn
j2O990J69loV133TLUCPqjBUrdjqRIiNoyC8D/8S0zPOdqcMNb+0BfGhK+rJYNhq
0ATS9cOS1TFPRzX7xW4ibeU5M5Se9i3nUSLCAkYscKetK1OoagEE8RAkccw75mcf
TxeHN3Mkzov7oULUWdOzrLULW7D1hnP2exMfKl4Ub+g0QjG/vVFT2emet2qmB+bL
zvaOW/Bq6n42x/z1tb8erA==
`protect END_PROTECTED
