`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KknszsF8JVGKVgvh8QdiMN9BButzAPYY4lCHAKbl2B4cHYTZO3e9R7cel5DcwwI0
SnojE07J/xcuLF3zspC0iwMgHde8/Gd4nVeyxVkVkez5LJ9tbfoFONgDveNAAxvL
EsZWflinVvkOoagsy4BmJIruxJKc/piCkJboPtYOZUk4qusbI7IUXzhnsf8bNg9h
SFDCHtBnOItQMpIGC27ATbFQY9oMIqetZk2D3zRiK4AVfTcexlaC/QHrXX/M4o3A
99P1IzfImSObULGWmz7oJITj9bxuH35wSOFJSTBdw2nEMPODFSn4HuuAxCtMqV5N
v2m1vOr+XyCO4e40gw2A38JwASZMU5g+oxf0wlL7lCY=
`protect END_PROTECTED
