`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3ofaNk8HgB4LJ08/h9pv4szLIgdyMkuaMU6y9cl1OPv5BKpsAJLc+oQiwh5UXbjX
zmVhHyicp0jnCgqE1gHdh3knUmPJQSmyZiASi+MFy/ZXXgca7gkP38YUwgxFQ/xC
nOAER22TOf1TY90luYKVG39yISEN4JN1x0BfBYbBxFMOYHygEM8nGywOnz7FSHnv
P5TX6K2sMXZdbkfq2OQ+Z6z28oa09oG1V6OL0S0MrhEFixtakYtpJsFBSSbKuBX8
zeec8mCuP+fRKZKpknibFqy01QyhL84WN7M8BhjDk66EvFNFLW+Qz/Es5K3dVwOQ
oRZtaxcjRi3YYnxnvzZ2Nd7scUl7JzuJiyiK6LcoXIx1xJ7LZZX9+EPLKTrRXDjI
bACN7t4O/Q54DY707hlGJirSijMW41lUeDeV3NxYey0K+n2BInyQUL2bjjD6jiuK
IDbDQ1sPQF86xtRrj3y/iNXNrIEocyeHj0UpG9o9vh3U1C4IvXVIZCFPz6ACOECi
stORyrU7O7VMmBs1Ex6FnbHtJhbahdit7EgGJuPYJjBXgKZVLLmtSn/FfOGJu+lS
rYWrWKaOe6ITBVLtYRp1zl9i30xHQCthiM8lVjhStKkjoJuQWOLxdGj/nzdCir6u
siTk5rKbZpaRqrA8+UJg1N5L8p8PE+NJ8sWNsNS/96PqvsVjnDRHeNLhmYJlL+UH
HzQ57suAxat01RitolWWeynK2ubLCwj2vBCLgODks+IIcRHyxcfgHaBce7NMmHup
k8PqzLsjSg25tYLhvQHBA4y0YSHnQ7WZhNVvIgKq+mqQtTvZV3laksEFi/Cma7Q+
ifWZtUDFO9djs0Ey9MnNtswqRskSRdfdLUa832W9WFqq7rR3zjCZ140zRKyBg958
kN4dgknz/FT6LwoyAsPS4QDrsezGaDqXuXJO42i9xZdN1/FShW0XWoG6k9vhcB/c
FjCsVi3wt49o5cijQOQsDriadjK70HHvPLsZ2h3PVMB39gmpNaZ23Q8bneEK1LLF
TF3/Ran8B/dKRVeAOvaEZVZeWcKbJ00PWBkWdZIN+Ejpb9bKpPl+6jTQRxaqeoVp
3nTwEG4CGvIAJecE58VqUGg0DXYnVDFdbvTZNqIDwzzngYS5XD0101mf4ALClBGI
`protect END_PROTECTED
