`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fDbKCo+ijizTgPrA6egVg2hQL18QvIA6DXSupXXJ4woeWuOOuSgKzLb9X6UL+BzL
+nPIrzqpDBf8kQkHQ/zLBu/mcfOMoi9kuwDB8t7VYdwpdZi74ojaVlE248WFxGpP
G9KXeH6tyq5wdTuPVivWLZc0HJGMVfcqTsd+VimaDPiAohhjXPngGW5U/UkTLCJ6
3UfWJmcpl51co7ybOGDj8Xx0UehPpPtJr1dTg3UaF5so8VM+TVng76UYXir0xLMO
gR2pVHfud7KnJnnEsvGFn594tC5DBtrg61Aefr+VMHswYbo0MWfmYFsywx5ErcqJ
RborEoinYusIf6G9q6fgNcPtaVgzRcLf9X/88qLoIzVrh9SN6X7681Uh3yYfiqlJ
f9QUlY3kL5xoM/423ck/1l+CcphrlpBjrflaEb+KRPu6pRgnaQPeRaO4u2drr4ai
9pCB+HtwVRqEuKVe5AVpJLtTxSazWRcxMNAN/zL+zqUnYbhMfc5KfMGlst55q0Vt
o/088yJ1IhmDMix7l2tSnE7uuFml6QD4y0nhZNVM2Cq+7LfWdJ901QovHSbC74km
4/06f/KsQDJSUpkMQxqG9aJLEBqbuMkk7bPspzZ2frrtdPH0zvAoNjRcMmep+Acy
AJHqjwVjEwjBqYhS/JhFwAkxj0dF5NaoIbnonwVTwVvmT4B3X6QcVBmm/nclWEc2
2+23G77npCyYpvOTM/XK3BQISbbzlR6dVXk2g1iyDg2pYJQhCIS5RmTBvs5greu7
Uq2WCmDIdkYpI77gC+/+ea1luFMiHVuwslx0lPCRBw+zmE6UBE0FsJpYAGEUt84S
`protect END_PROTECTED
