`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IpiFjYFjSxHUuBnxbeOE0ssVFBr+4rHt46qhI5e+oToGwbQxDYqbdB5E899TdyDr
+R9lsyxnIHMW3k1/YUYhAh9wuhfcmLoYiT0STmiOAHLqSpXepdswe91gQuPY9zg9
uOPumgrFLOLAFXo6ZSh2qc6IpyEy3uccJinwokp/LsC8Z1ErJjXWp6yXMgGP69Ne
jBmvPqylsGtmbiOHP23+r9MzXeNxeVDp3YhlMAsQpz4oGE6X/gZsBjDrsK99BVPH
uXkIBl3utrb8O4MhRMpXXA==
`protect END_PROTECTED
