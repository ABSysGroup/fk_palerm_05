`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d9MFJHUXENS+nD1uxhi/89hqMZufYS4WeiSZE8rHYBQSlbI33TCIXrDp1j6rwVFQ
DWq5T4HcuV+uVwooNiVnZsNHNZHYF/j7Mno9GaCCY8UynCMr4WExiAjSsokja4eb
feYsJp/c8+Xf3w9EV78GX7BNBPUq6T8ZUjWx/9UXpO4q1KndKp7aHEBpLGRGwDsB
boBYqniheh+0sj+puXSrk2JKRSfq5XXUO6T25SibJAmxQji2zJzMoI43OqSsGe3Q
apfbcyRR0035ZEkxpHcdNs2Cg9d5FQkSddy6meOi4+QpsJd24nhFdNwZtmwsbOkT
pCkEXYb9pxcPVtI/vuqO3653VzxdFVQ0zQxSLwKZAYX2cgeU1IP9h0kwLGNr2CH4
xS7MhUAaF7z/mb4ne8x68jsJCUhpeoygAC7na33HJgo=
`protect END_PROTECTED
