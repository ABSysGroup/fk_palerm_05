`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4k+vQ+hansdRPIN551tqLTe72znVq0qk8ZhdMCOKrqzW6jA62z8o+91SgeV6GUZM
KJ7tC50K6KBb4OktAQ8P25WZMkP5EG72PcgRSHnQ7xQHXqSepz5ao2OXxBjHaWSG
u77MvXDP6xCaKD8vLIzPw1zvNOZSp26homfyztZFMKYd25IdWcydPFVm8/B9a1sV
l93Z7TL2tYJEg/Tjn/RyX8FZ8hz+bT70/qfskrtM/xlH1J2irYJzbUE8OHN0BAdN
vVIlyLYf4qtwMWEtepUG6rflXYBjDsTbH57t5SqEkyX+J9UsmcNZi1wPLRaLyvZU
mTirHtwlFw5i8nGzQLer+t+lzLQXRu5390eie5Cgq3UZoOQtpU36uhGC92/cAW/n
4AfKTFC8PaeRmighusDUDqBectkTpOgrFxYd0/MqYNWMDv0QpOqw8GbleElOZShX
Y1MChzBzW6V738s5fS2O0ZdWXB04NMfzeupSjMYTPwM5c7ONjqRCXrl6a2DI4p2w
6lHnjd/Qn9vJtyKzGrCtsXa7ozcnHXyqoYvbJEyRSrojWCNA1fmVDrCC67a4IM5g
sal3x+c2jh2nJt2AApJF9GFfYDQ0FyeoqluKX3CLlHnr8b0NI6wxzKeP3spFkXEt
uU21UDn12S2ers/RnCyQaKtpnkPyHXMU2xg4qpb71Li6MWIm9+levT3tB3dNJEsU
0qfqus+fh9ciujFfVF7mSWi/cXtDC2j2d4vYCexDon8XkLbiJ7shShS4Ho0CTNeJ
pO9rpscBRt89zh7sJw/Qhbc2oy7ndkxpXbniPNwwcNW1MlQa1K+uk9QScvnCY26c
oRUwzjUteZNvTzAQ7bR/KLaIjDsToXNt+68deCH/t0CFIUSz6Y8QG+kAE9BN2TIs
FUdDAF//PVh3plmoP4j2mBAWvntfmmWTHZak9GocZymMxsuSWsAKhO/Rm5ZZhILg
1+8HbZoW0B13I+QeQAR4ijy8/xdbvsk7UCaJ8xTmWx+WWfJzpSYhsbwb/F+V6cnm
sj8wVy1+wrCsxajjDlS6N8boP61zFT4kFrALcXN2Jcjn8upIE9QYOVnCyE7WFuaI
BLcr7BZ5Ribrncz7+VVt89w5+0XR/Kr0WoGsSqMw/SHt6iEWAVzfqtJDSN/qolxw
/BrYWjsFQKyPm5zLLAxTGIzn96/tJxNlN+3VmR052NK55BYUTB5YX0YNW/X9hIGX
d7Y4o3+RLWLMjAnFRS/kxdG9ccWw+0/B1qwnepZ7WaQFH6/BLXxUxEYmRuslwc1T
o1j+VZhJ9alMZPEMcw7HfGulNqqNID6GbU+dqzZkm4B4fZmk3HcfDsu9KZCYmL2j
i0tRIsyGI+4yJN6WE41v8Ne4ll7rmM/VbqCam3d1Cd+nWB0g/UhOjnwxBVOKzGOM
ilt7EnxVtGjx4nBcY5MZgdVOcvE4qskD4KyzhnyZTVqt4jXFmivLS8QsSgBggQ2M
ROSESNQrIcaP50DNqCb772fpiYdXeWLHuodKAxK1Zp9rAcOyOI+jf17vfE2eMN50
mPQMOgsKXeuHEG/Uakvg4ElFHBBUBDCxPgscLRQAyl+B+licsfIs3wnZ/S91ZV8/
8iqKcFQZ970Jlnx5N9PfdUbXj8K3spcjebXGHuKvmNBPqyG8qwZgl3rNbiuXB1IX
BaYScsezm0nnsDxGIBYClXvguSFbd22Om77gzL3Wt+iNE2/NQCGMIGRnx0okFPpb
SOj7sRrFHslRo+9WdZRcVJjKj2xx2TE+kXnsTgyQ9+YGnFyv18cRTz/eGQS6xq2Z
JU+a2jat6wf/f0jT4xjoNqvol9HGYyilXzvmfzlZKwkYqHMVEOG0TwkHLiT4UaiX
Sy/lsNWfz5WFB+y3EsgCrmjJ/d3LYMj660i4Y+q7fhSpYEjaEV1flIoPYB3lhvkJ
NxnydZ/y2+eXODRe4Yi+4bvMF2jk/Ek4+rGD8kqVTX65t6smE9kAQirfg4x8sGkD
gCWBytTfxgUVZwRn4gZEa6vFa3xSKEQLyi+d3wO4gVhz4KsX6NyR6d8wwig26iFs
cO1jwbwMvlvlBnvMHUGmjPQdfiPTRn6Ypj9N5l7qqm2s5xzDllPdHnwppq/nIcjT
dD+DJ42AqdPjH8y+JEpGaRy6VjN25xT4YA5cNJC6YWT9QYzc+38eNKH939npHxPl
j6u4ev7mp6NIZRGT6ImoY/2Xmlw44y4tY9lcRiGcQNVxYQO+hAdvxsYl3SKm2dsu
qq35PQ9qgrtM9RKRQloPAFB86of/kr5Hf23Hw4POdbVMyzzOC170QWQIkUT3/L2P
rMIAeg0Kp/hn2VFToHfvNtsFNqwdKZIiv3r0CX3zV0DeENi3fKtuGJ0eRPlnY9dy
Z4JUDK67F3rfIgQVfOhSDhz0/INVtWaNFDvhn6m7KrZ6Y+s6uuSaf1SBBiIY247v
/21L39Kpzzgy1Le7Xb5FNf5481OH/V/LfX6KojjAMKlUMmlbJu4ZL6j3a+KIyM1B
EVspVk4zesvtqSwL1K+0P03ohL7fC2EwYf54XWum0qBq00ez5agnQS+m1IffpixY
WIpwDY9ML92JNCdU/a8tgnmm7+LHDePUKbWNd+g46c/rcMd6fX0LwsLlpQr40c7X
dh5COh4AnQwz+DkR62CrSIRJ4HTW6Yz0Mwz2avU/CmT6C6rFctAtx/YazERJxnkB
mRDn9e+FtywoQHhsTQ2QyIlWdCCZfZefj3/DPiQO3UH+k1Qn31xzhaepbqOysMv5
`protect END_PROTECTED
