`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y+sfs19d6g44BesCRiJH40hhXMMfxBxyskr9VSQgCmktgxxb8V0IUC0hikF/IwXU
9XeUxQH5U9vbVO9IiI0texW/8trFVZZ5mncYFzfZ19jJuVwsyZK86uz7xrkbmmLI
9qj78ay5KHjbMjMkQ53znS/as4Bv5/uBnUDQ54PlmEnKHuEh5LB3IVoHoqHNAHoW
P13jSNMk9PFaETEPncYW7XZqWuMw4FWf4dvLO8Xto9EQEZ9RPXU7DTzv2+7JKUvJ
CzwESaAycGyv4FEW+huWvsVGmpoMCWI0tlKO2KsfHvXNLqxq2rYuXFWBh2LUPHQ3
0HMDLwiHONjMJINM3ah6CPQTdNLe6pK57PnQjf9Dpcq5FfwzrVrFfhree4JuJ3+v
p4N6MKndXReXeDgqgdscrfzDXnpAGmxz2QRa/MAddwXlRKDtDZfb1mtY7Zep0LWw
tiDHA+wzI65p+sy6GbabiipxVaULkEgFM8TgR1GGq00TU5VXZbE9By40UKB1yeHE
ii3vYSGQzr337mOP7eGVlKidr7a7qaNg9VR8MiUvMLKcJx/QdSKb6cKYWd9svcap
VtdagRN87T9EoHUfF+bAWLb+L/YPPotsIdoYzezkbzA+T333r0yKG6HYK9do8HTG
IZRiQUQivE7awB8GAyMtvRkuF6QXkNJXc+t0m+2B5NHp0jEecp/d0/Ib8ZRWOyJB
NWWKtxcKvehklrOo11PZg/9mrEqSb7vkRpW72OaoX3jRAIChcQHmBYkmLMAOLrKx
BG5C023w6o/lcsg4PDSAMyzPTwWtLOz6hu3gvkRSo19Se10kukftGs8iQgfAD9W+
6l91STgkANiakFP3YY6xR1yxb8V7MdHXmtd8LYZhnFpQSVggD21rmCT2Q3SxwRX9
c/pGOFo2qk6xFeH/L0xjrcbpDmA/ghkOouRcEA1WlNWOa6TdagKcq4wVsINx9AcI
ZL83yuLcAMKjGc8b6tYBGLvLOwMmLQ+arCc7Fymos11ivB+vQCFZhV5T4j9TaOTs
J7ugYqhivC0AiU+1/xxv3ohvmBAyhnDCDxY1yZLDTSTAO18ZkMZwRc7TRegCYBPA
7SAyKB5DZeM6/n8etyJRSbJnb/3nljYv793n/DcTxqvPGgLlZJapU+uKVazhePF2
WVfqDaCB5LZ9GRKqvXce/fDwGZUDv/2ZqvDEfph74cSGi9uYWGNUaLD2d/wbHM4a
T0n16PU4CVEFZ79q2efbzufvYf1oJq60uFsLKZ9bTx+AvpF2WK24pKLfhygCIOu2
1M5cuFsEe4z0cGAYQglbuIJavryaV/csZSsp9xxU5Ti71QweWEREndvuwce5kFvX
GIjxPUyZKiOWlQ0rIgvWSie/gFO0CUlmxnTPRAAV3UX8oBYg1e0HYTbQMpMSMMSd
OLNbEWmLDnp9XJGtmW0DxUxx24750ggggI+9wq+8kEYC6YsPK6dWTkb9+TtaMJIy
8xN95QzWnCM2Jx9ouejaqwY9hL6glImkPPR/dZso4Vhxguzm1Nh2eR1MkiJPtpQH
eI1AesyBntBnjHN9lfwohOT4kp+4sdgYRuw/v/fBIHJe/q9Y5HT4h7Y62NXIdPkw
gVtB4qELPkU02UeIxQgD0sbunqsHPmo75APX/3H4gq0vbnkIwdvpb27snPr0UO2C
J5b5tDefVswElXP6TO1PYX4g5rmEeooFqbHPixSG+8UerWMYDmhZH5JeP+DrHik6
InLELWFqcKYcg07SHUZ2GfTKHANMPVOnIm0kDb+OSf+C7WrtL/D98BA1+JdQuoLm
pJXRsJ+xD9Xwb1MV8NGRW6xG9ZF0ErxiKwN9gOO7SmAu2ERxPFlPVceKTRZCbcU9
KMg7pjSte9RKvjQnAu/Ns7qyxBtbgc1mx9zrmyKoqmh9Fg5iKfgqt5QQf8lKaZmC
bd9uQoffJj+A9/p36NJHU+ih2UuXp2TZIdz+AmCP0wJdEZ8+nFIKP3E0y7vGcg4i
7SrvgTmCeeJDS7lsOBsxttLTmbgANuqqalfWkmsDXDTf0/5XAUWAu6F8zjw547d9
ux61pfRyVcs9M938bQY8mR0nWRy07iDcQhoshiiE7TiCIx/i8PgSS05sLj3qugvi
WXk/0Vggjqf1qA0+/sd6RplN1+3TJoHE7OvJ+GIu7JQbVCZ06lW4fD4EYwP8kh/F
D4+uODJnWyBALo7HNdg0DOh3IdEZmo00HpVTquylW/XesCU+I9ZjGQA5lg2F/PrG
iL0q2XLJr/Gf+4KnnHWBO0vO4JtfqoKWgPUyYnDKK4ClShwGBOR+WCE1yaB9NMDv
1jkLZbWtaVw6z659nqOOToUv+IIRmCSti+5gEcKJ9iLncups5RY+cTww/iOcNeF8
1tlEgBSd+W/mgUVuw6WtGcuDC8Xo2BsuZM09wvj1eE1mZJHVoPMU1nZFUBBfwcCA
HNK4j+g6OF3UsxXxDR8WGgdyI/swdtBQBqQ952TfbGCaFSrVki7Ga5BszsN3BjBx
Se/yUjisovlJxaA1ij5rbFx7Y+1YTsc15OjVPzK21m5L0rm/EGJ6ZC6etyiJHnyV
5Z57DREnnQdIcsIcOcpjRVF5a6a8Zy/qxbgVfLT1o2kNu9jn7OUAqBJyr2L2Be12
nKlVRvZozv92YriDXHkESLX/aaThMHVhGLqfoauqLqmgHl2tW195JGXjwBnqh00w
DsntO48P1MoWoE/sJYbjGKcmYgdUl6lPdvaBNJaGwZVWaqNQrfVf8rXPAIkMDEg9
FBFQ1+114nNkMtL1Q4WzTDQexrFcCIQYjgT10WqRTjKhpBVLEv3FWccJ/AO7ziCm
/0vCNaUcEcR55RvIvo4PcttR+ZGjDjJs4153Xe48k6k738tZVMlZ95MvM74C0oC4
lHBS+uJGIkXag58iqOO6J31HnlAm0UNhg0J/9ZPMOWY3bnNmPNWpO5GcNpTaM5L4
x+frQ0sesH4hnLfqkcTtaOW3/dUt1rWIfVhIp/K4RSVmmMybKnFs0Zy1fO4a9d6H
+rfkUcJ2n794P3sq5Tserpv1bMZbXJsk/9F4PY8URKJSPZAHXGXKyvze5UDMeAAk
KmCChbroBzZv1RZzvWOklzrSCj/wT4VH/umKsaZIdNtFwsaScpUpyDkDimRE6q4Q
dSgRC32etzayy0vMLuLw3Q4H+w3WqcpjxhbRkez0nI725y0Uo71c2SwQM/P6ZLer
zqozNaQn3M1eL9t0sXTnI/7vD5fLg571hvrnuJXsQ3jYPhRlAkJW9PAiHKW0Vqxl
48K1oEl+scbdi7kDKeA4AhBFkPUvcTfWfDcYk+ZPpOASPWEWIILm+Z9SnXN745oU
Wm+Pm5e//ACOm50zFd86ZiN3NGl1YVOtwjYARsuY5PjT2BX2pkV01WpuCbCK9WSA
pcwlK/+fZPdH2ldSjULgCA3KtlxfkBsvyqxGFcWK2Yq2RRV+Adsw/XPq+YdV9OS3
ADSZbw2pdlf9mXAS+0ddfuN6uDpK/Ap+p2VbPEekZ+yCfQzjPDNGG9WLEnzXMX3c
Xvhc6+hiQtRLvyxUbD5CG26QRvjN2JD+ILR0Ortpf43Fqt5dOzPFipZyR+pvNQNd
hXUlByhgmkRhWfEb1ozMhFo1/nBYUUoHU0+qUOcu9Ewk7Qt6LUX785IqSG+8z1Xu
VNMclDxJ47p4fh4ESdPe3YkjFuJ0KBT38iGDbKOnKNkBIJQVidIOAVg36VarZcdh
ZS5iecWacz/ckFiZmpDSeTq6CWr50Ni9hmzeSE17g+UqssE8eaeOr2JSmVFFc4af
P5rfOtGEWoiYXvNIhfITvcBEw4b1K/vbwwnKbBPsL5MeXo7K6kJ1s8PW5o781QLl
pfqSgOGz2SxRVliNJNot77+Vv8BwnTCWRRVJ85NABAcITNyqacH7S5qMFvUbMC9/
5eXkaNoCG5wwBzrbqMQx4KX5BWKC1PI8SaSIGNXcTR9R5qb/h2d7Ss43XgkGM3v4
ryRTYbNmJ7C5+qyRJgt09JB2qu/uUv6+iTnW6FDsJtB1pfx4WcDUB/n7qYj6vDG0
VYghseG8H/RSTDH4ttMRXhtiEW0tDb1D68koGqWOJOTcFQFCOUBotJLVRnNNE4IJ
q2/oTERLkRuaVcm9sM5339Cg9Ek9rKn0qUEnS291/1AtzL2Noa4jWayey3/z2eVv
FmHKYBgoDR3a4Wlb6Csah7rXqpGk7F9OG1Fd6G53lZyEAnZYK+tpkz2cxQp2WALy
oibfMlsNooTKIdpWfzxkv3qwKILZ28hQzEvNKVNaVqN14P/RhqxgAu8gc2kidiMW
9cb1QRq+KasmsVlfKSCxes+tX1Zm0cI4s4pw9DKfT7eG5qn9eMHFEGOHn5SUlu+4
DDvaCnW78Bc3xDCLo1kgqZJBh3IU4umQ2zOCuFK8B3+yBYhgYWr12AhLXq7p2Pw5
4XechX5M9kugR+r8UM+jJQaukrUQ9LhsMHUV9Cv+mBVEpUDdsD7+WdmsNlgfGZz2
g/oD4JZSPM717vBCHAAfC6Czac8FvavzDt0Sxs/z8lrT20981hrbrb40H09sRqjd
HXFb+15HKjhyrwo9YcCaZO4FyNErf6AnL/5OF1jPR8feDnuDDKnYKJcU6INAPJFn
Z/rFWjmLN4KehJY+4J4NrcI27Pf1MWqkwd6/pV6prq1EcUUneQ+LhRg3nIgssg5q
6mXqvh3sxCupaCVhtiow9/63FOgzOemiMTa+9G74jxl3TRrKENK4Hud+zPnYQBnU
6mAT16TQ9dORXuDZ0jvVOVOLJspgRu9Grazn0Ee2l9YJvHWuRViZ4ibGWLoA+gaP
4qVF0Tb/W3S4KpULAeavjpP7oNBkiU9T9IHWR53ZfDAXpsXG32z9OzOBQXBpze9Z
zKslMEWAy9E6OIZGc4B4jxPIQ+oKpaizQJwiivBPHtDJNQQy/XniULDNg3KOp2V8
c7oreOFmn4BrjMiXzt+iXgzgmuAwHDtr6ZCRhXgHwaC5OLAba7NDH0xR6fc8LlQs
OkPEyqICymrCy7XJfQ8h0Gk3nrH9uVmteF7IfWJ/rQbrEfLLZbYYEy2tNRSboABO
1FQuKjxWLsBeUPrjceOWjOwnwnUev/NiWp3yhGzRyaQM3CIWNS92mhQJ4RikFl0e
j6sssEHHDtyf5KsL6qTbrars85dqiU5kS3CkWcyFkkt8MqE0IB3wIb2MA9JvIkhj
0jn0JIvwzLj4MBGIIzQMQNP1Ewy4Ysy6uDif9lzBDQ51dKQIxVRmheutscdYAW9Y
GlFhp90ZHFe8YcohyIQ8LR2EKfLoA3AAHQId+qF8Kkil6QwA4TJzbwQ00Wt90N8r
VfQEYhibQ7rxr/tKQ4BpoSAFVYVnrxpvT/nMlQ8xDNLGZq6Zpa9VSimS/xExFJbE
2t+SfbkOVxe4o0VrSfXoidGw/Y3zHZLUthQ2y+hk6MRL0xsP0AFwcjoenoLHJJcn
vGv8jYDWEtYWNyRZO4sgUDnvZ2bu3OJqgrrrN5tP1zR9WW5l92HF/KZ4RiuCF/X1
Hx7jvilJ1XODJmtQH+WmntN0io/yfXbG5IsrYcvfv8MgkdI288nWS9MqdXK0IV+C
hjRS/xcXtBTDZEQVIQu1BaRkVON6kT5HOkm58qDE7/xiTF8ancaPRNcKQr/8/Fju
g41qFj0U2NFa72F1Gh/nHyt+ffQgZq2uBnWQdnhTGK+6aBl7fVwUlzWHHPdTBU6l
4qR8YhBW18x41rSTqURgiV+ZhpoQ322E1K887SzwV6x4KWKyxm/oKwoB0D8wm+Zg
/bjvLS6wGLJt+lYR8C5N9GGb+I7I0UnaFOEFd2h0oPD8re8FMJnFZuGjFHbmsqJY
NbMzP2tcKzdmLdTjOq5RveU2Sn6ZIxty27WItcBzc+V1Y6GYhxwbFNWYhrba1sDJ
FK7ZPXgI/b3cIvBA60/xo8WLNpBiGMoszsfnGJXyef1asxinUc4Dwskyai4T3hAX
PPlwjFS7K5SYJfOWVjNeZV03TYkzbuFpzVGSUp0FosbHgq/NGYv/WtqStXQxdWEd
aUqnTxyCFb8D5DFWd/w9684q91xztzkVVZDi/4F6t1UQhz5yjuPhQzqAzZ7kgC2h
UFNpQm4XzAavQu7U/inN4lAPSI5MzvO7n56qMUz5KXf7YFbVlfvuPEvrk9X8RpOg
pjl7R7RbIlOGPP9vaHTE76fltdWOYFBGbagydKQVtunx9TOsemtE5+mNzXZFsIEY
fyVmzxmzeTSH5T8wLnFYez/WckPhT1ITj77jEhCsHnTiFQXBpkwmjlu0hOkmisnN
xAq3FiJ9VK7xj61zdyZPYyhWotSiDumOnyRCoXwUVj797QhENGcuyq9kpM9pV4nd
569Dg1zX8jOSJJ3SS+fBoGwiXzWB5OaRPu1UtAJXPmxsQYjY4gri2Lby1c6ARbWE
ZjVv53lT/v0UcBq548YBWEICRbEoabnYZfMAifnYPBG+cw0jUkhVP6XnDKzkbmIi
4ShlbUsLJTzJ2iUJ0/R4ae5NAbAWEepcVLaq9hkC0OC1ELs90Z/tcIjU+U1Ks9co
a+YEfB4x5a6TF/N92AJZpLhmgsb0TPB49/l98SRJ6rEkI4xGi5jkoIRrvW8WcTfz
NQDd4d5xa9zMb91SQZZi2iTk52D0oyHMSpmmYKa/T21ujMQ39JD3Rw3TJlikSTYg
02hlJQRdkrR2JTnz2N3cusGEnQ5GLRQXQNfVFL0eTaXasZQ5gkXWcV7fbVhf/38I
1gGiYvXbd7hHZGqkiz+yEEm8XhDzVbVlMYLAa+aTTIqDoR7CjAVO/SPTbaYkc5+M
/M4fQV4PB0rMaU/O3fD40dmDJMDr6W41wP1V2+Dpe57GsMHf7+dGDogd38msqFC9
asNj4JuDC6gQ0BsUEDQYCfCSdhgPlsbomXTsx+Ygm04bID9RPEAiwNRwSAJ/7fr3
viOG8GuMhUX66CcwKC2SDUr3lcEHRFEi91crfQ677Yw1CDI+/vKdwWf8t1O81+sd
7YoPtRzAlRUrGpE/EP43D+u7l1p409bNSNLP7geQCdRmZxximCFd7jKfIxb5+LZe
lSQhmi9dAZEByh4TAbJATxVcMV92Zrr4i0I1TaCSpt2ff7fxVenmJcsJw+HF3ka3
NIaSzkRUhWnPlVE1CmODsrIis6stlQjRJ0o6hgPH+pFuMu9IjpCBghBTyy/eODuA
lVTsuGP7ya/+bw3j8NZArRGiqIcqPUhC4upWUV9egkTczuSgZgdKcQWm/cS0nVbZ
M7hODsoQ/Z7S0uT8bOWE24LA7PQFcecI2r/MMBkHg2+bCURJnmT5NI/rtw9+fZ5f
QUUguy8wvFhrpq0jMeRG74i2qdKjGKRnutODMC99u73zoOBBunh23lOkD/yBKVVk
DdNRmS7fGOfsje15VTuyvADtqDLEY1Ef+lydxdUwkHCPQjB4ImXhwy40Er3PX1lm
QE0jDNarF0mgywUWOKllRemFBeB6DzjnBlv0/kKXxvj7Wd5yLaNaEqPszMS2pNR1
lD5XfomfHdj78xD8GkXKcZD0TvyVWZr333vaWvgpencb7yN5VPJFXrwt+4INeP50
6+/TJx92s22LPNubs33X9MqrFU2aiT8gBKKDuiMNNtNwQEQKQFL9rsgEzc1VLhCO
K6zoDSAkTS5/D7/DpAdEv2mZaBOVO0mtWcr+PCqxT+m9zoe3D3nLNJ0/0z+uWj5N
uwSl2UwGcpzAb2/hXjLsNLpj4vzkZLfHxtG7A1ClcIVVZpHALd4XIIv1z7fprBU9
4y0dRBt/vmyWOhVdIfDfmzgELVSSuTzKRykBfB0Kk8LE0+aDIive95UtxEjStTiw
Ve5Qen6WdsIA4YZD2i9nbtNV4gN0MA4PjP3/LZC8h7Le3wh4k7IsFDCTnFjkzabQ
IzHpeZlUucjmecrHPewv1SoiuBJNN3i7+KoW8Tr2fM3jaLf/v5nAUGzrTpAuCeyh
fksVKzZJwJKVArY4f+NUvjRBf9jwTT8k5U5NKYYf3K/OPgER/FLZZ7TGjuCzYr1A
31oCOips6HBgwxzCqjhD2Uv7rTg53jbwJUwBKL15+d13dvccbeCkqddiqL86Tc9B
Ea13IURgEnlJMxxptCf0ZkMPa+SO3oyFQmTdwvHssdyW0R5aGD0xVQiDcNmgxtm2
25fIKolz2kBwHcR0SYx75urdKIJ996NRcYycQdluIGri/M2d+thNTEIoLH3oeeWN
j6XyyJ4vdx0Ms7HvR6xErVizqmBWjnDbmUAB4e/SdUXmfzJXOVntnYEOk98dqXuj
smZnUgfLSniaTd3U9KqpXu0MRVl2WImaHgowo0ahSVDiRVi9JrJFYiNY13nbhUA/
WMZNReT8565KetkcNDb0xojMCpO/XmYdEDy8sghzT4/r0Wl1ztAdHovuNPHHI5QM
fiuMIEvNcJg8XHXw2aqsKybGhu/6Byl12YVCCGMHpvbqDofSU0VfYMWsdJ4lja5i
SC3y7SQxkSBKywtcSMgZuGKjPAVjZd0Ekm/shUjRcCHzqg1FVIJjdj2B00JhZ8Wz
szyElOe/LWqnA7uQH+Tt9fAonY/S43Pd+WlXzsIPJWfQOoPkbGpT+nCB9TGDJ78g
rQHy0AvfxgElsJaexQ+475bP/jYzTEU4RqJWaoBO7xD5pk7qyRxHwGV4eKlO9dv+
+ptKs9SZmM3hsLx8Q+6ejKAv8/4/ZC/YZL2KQ7FurIqkT28RE69ITet1qA+Q++Nl
Hn90jrryAkLK4cC4WPY4SQDiaxvw1L0wztrsMCj0xaTQ/JFF5n2wJ84OTv3hcUyu
qOgvOp2kQk8wQCd8NTwmMZtsuJYme/VMkcMiqoXbC1HsBlegcTsF4CiG2K2SSBxd
ZKR0UY9uyavq+VAmwCQphUCJvgXRWNBjMKULYOGDzBiZIozZTx0uVmsQezaTJe03
x/C7AyCtBZYMaArs+jXL8eIM+RqH+JavIWaBN9S8DstawZbJOjdnCjz33SJ+1z/R
AbxWvQ2jPtPca/vpuOwl2uzpSzeOepGyfby+olpXw3bo4Ao8DON0uOIFAnmij9Wj
lNK2m7FOaeCHIxrFWs3deJRV32kpJ5LWRV2M7WSiHw9fIQDkKaJhYh9WhY3exIRn
COu8/8PcrZUXrfKXfVzsgMs2996SXZGeqozkmnvcalLaynU+KI3bGspnQ463kChC
orp74NPanNmE+2gk7ckWynq65OK8pIc2UxXkDO9T7vX4eSp8e1UpXy43t4ghQjt2
fnh6+TKGUi74/ORKf3Go44ZEq9OhIHXIE042ACi5Wb5rfIyd2Tj8JKAU24+l8wN4
qdCOwFtkLVa35RdBbUsbOu3jQ6oRgf02+cTmYf/KxKBTEIpeR2YoME1fero873qr
UwcisOTLPHdIFglXO0OVf8I/sOuZu9cKYPX0owBB+3Uif8myEShCvlmpjQmGpoLi
1B55v9ARcuRx92/W0Jfqe5a5UftkPIAxP2Kuj0SJnv2pGaU4IpedMY3Gqu5StGWT
Q1HOMMvGb+tGnhfoPc3dENo763UEPAUkF5mvaJA667UV8qnZehYPYe8bnIxM0mnn
FFFS06+y3uQ5CX0fvAeWIs076DIplCQDPJqvy5lVykSTS3Ut4Ey2Zv6uFNDcwj2g
J6zsYu/WvObWuTusBGnxO5BUylz4zjzOMRwaBWwNhW9E51j8ss8I/Q9WDgQ0U5yh
tvVOjUsd4nl5+jmL4X2Uxy3sYA3qADXRfeoyoZGaTRIdw/NBzLSODDBdVfs9m1SK
by3kNxp72T0OieXLDEcA7jNgljlZW2oWsPZ+AmY0rgT7wjqrIgp39qQPh51jl/25
PpUC6uwpwnhyJgSbry9/uUmsIbnLwsVHiVPSw5VKTCQv3DBZMmGOMbJhak4pY96z
GaRpSEtbgKAWbCTlhRweHGOiolZyr7HW3oxbiV9HwiQU9mnTIVC/zG245WBodtz/
Ua0KoOnNllZdKvOqJTj60wyd0ah1fw1b9qgJRVAM0kCReOhyvyLFaqrGjxAg16NK
vLl6Hi76aNYbvVWmXJpCjudeF0Ejll6TuYixOEFr5iWYP5v/lsW851s4b2t/01rM
2g/MtHX7dE13Q70HifgV9FUdJjgzeuaQ4rUdA43Ov7Em3ZwkwAqi1UmuJFdfPs/F
g3Xpyo1a2UZtJPA4SnPE2G0//GIhnc7vMcm8NYxe/vmHm5aJ0+mi3LW0/qhn7p7w
Tj4hsEuDTb1hQ32SyjCX2dAKi+1UtiloykhBzH+aJhlD4vO48TXzWmMvV9IQpk8M
H9id5ZpOKB6bciFdz4pEF8EZZ9LSJw9DMDmfFIodw6xxBbik6SaH61cilSGcT8FP
ZbEpGJIFtplXH7wr7g5rqOTKsnLHjW+ZKjGiXxVgkIRi9HVCAkRyiN8qznf6AVCj
6hFGDXXOmE5PfWp4xL8CREOgo3t27maY2sehkpnBJVc7A5wKpyV0W8Q4y0OIHMzY
sG+88rRHwPCfQ3ZV1XzYAXHOyDOa9s7igGmLnipub5ykHdyOgVG1u7IJROHLUtgI
adJSrTARdUJU3lIMyJI4AoKGlec3JhSm33mnIRZTBC64T7ROCYi1rzygh8LDIRJy
K9O++oSLFlpm27AseBZip4RocC4XgkZokE/Fe9VOFZCMCZqQYVEzW7roBauP9VKH
negH72ddbRX1MDz3VAuQMUKeuQ7N/rTcOLINg1e1Xa2URxAgqtqXLaCj4QjurpOO
NnwZ/m/CSHCmsGs/7SC/fekVz8ZhfX/DLhNw8suj9yO/WcxiJmHjVe1va6g1CiAV
S77p8FxYEexp7bbA3odQaIykpE7mHwoivxv5l/5qdIjJ35yzGHgQjZ5+wcR+kujI
zMqZQ2hSRVmbxj4lQu4Eq5f9qGrZOJzn4FnRleGdUHe5MSDQ48G/7dG+3Fis8+o3
baO1xa78YNfgLDmpflhLR/BC1vUMxArvULyUSo1a00fWhP202JkMyXLJ0IutQk5j
6LvfrCHUaCKF1VMh5KDcz1cnFcnn+ZnCgaYPEQOqE0nHPv0dJlxmyCZ5BGl+nWo+
WaeSJpdc4WB7NlDYEldryZb5hsA0/A5QObsZjW0Pk3wM09VWhQHIsyG3L+SDsUEY
Xp6RMmGYukIjWeZ9by1d33s7jGHXioT+WMVXPWC+sKUG004TipTvghFd8TMg38XH
Qw5WYSEbHCFCUkvGkfUJVfC8GQVIOvxgYC72ehpSaanwJ/M83bP27r0Hdhxa/l8w
NQObHjxphncm7s82oli1o2Z/TzQxM2LsJTtMS0A7PKj5oZgb6E08GwQLQnCNHxu+
cI7tdlGsoOnCtO2WcGmOxpF4qhPKF0OQDfZtNr2oqHZ3LSdzRi2lyT3a/wUSItmx
i+HRYUBwJtJCwdVYLo1W5BZPywfjo5viXgTN3sSh2nXUoW8LEGaN4Y5W6YOACdoB
WDwdcJtNwX7gxLPgEwuY9Ol0iipokNkRo8ig/bn1OSIlrLgyDg8c7gaG3NKVbtz3
Irh5+o7NaAvGZP+q5YS7Qdg4wcPPfwZTbWj644UN8d7i9lKEddD6Ec1qyvi8q7JL
`protect END_PROTECTED
