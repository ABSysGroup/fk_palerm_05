`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4h82lXW9sfMzB3DkHN2OT/C3RXcA74Gtl9YDEjvBn664rZ4uV+RE5aVwS9WTxjze
ERCHGD1kVDEuS4C7NoN49WtwjzjN2fVt2zuugdqjuSDsJ1Xqbo+3fCrY0ZGP2i/u
yITKoO5u0Ct5sfuqC/3rULM0RtqZAibwnDgI/bVfVKlUuynyEcSAThf6clIoGhq1
Y/V5nNqkKbLFax9NhEwMp0beusz/X3ReKmRIj/emQZGqtlDTm2ISC1bxM0WkIQA9
SF6CKhNkWDgVDFXGk7RhlzCGelSxXUXJFk/hCOvCz/A0AmrHEB75+L7lFdX42wa2
HVxrH340kk4RxZeHFGGgOmYcNPvT1Pjm6QCsPFBvEH70vpq+t5t+QfpIjtJiGeFR
dq8pdaUdt+l28OG9GyGqpfe7NFF7bGYoIRjeZ8UjfsNsS8htvIVJS0ire007Z/AZ
Gbhr3FGnL+Ebwud+pOM5GmA0tkHHTfPmEZSMraNm4QJ5imr1Zc0gQes5w5JJwpJD
/lckgzabPtej+blrfTTk9Sq8E9brch++lB1/nuJEUHhJERCEGE/hwYtGHBPS0uiU
l1LmHJ/0X65x6kGw+5CO4z+OtTvPi6TM58IBiAd/zYiNyTnSEuJoJe/esNCBIiGh
TD5d373kOMsgsz+RqXVz7LWyg8wjIcD5OsFgW/0PqnLvk7+4P4HbjjljnzB0KKpa
mWAI7usLeqOZu3P8c66+ini/AJGp8JyWOAjwwmBV2NSsGkpXDfrIqeX9xCayYHGj
eT68sZkNkhRvyN7mlh9tM31qDUr66is4NbvU1FYXoLBBbhO3yryFdEfu9jgEBFQO
l3uCxo6odmoJdIqQSAc6T9HuHo82ZB31AatBkyrDonR/doTm6yVi/63uF43s+oRr
VwKCRSJtOAOHbILwyywzVanKHtnJFLCy6oina/8XGtmBVnOZS7DNW5tp4WjugB5d
oCbyFOmU2Cy5npmzioONaaLA0Yxx4vYdXrVJGlDXeiLGd2HZbZlRMvGHJFJ8BAv2
PW0q4H77bQDiD4iqRtLquvsSC2oTtCiWTc+AtFVa0LayQJjf1A7NIgdfzf8mNhdZ
ZsWbT6I1+i8+AhTIMbAvJaEbUGW6Ulmdnn6TWBVqiSgUEYC1D1als6u3bY4YJ6Vo
MnfD8gFjJ+N3TbhLmrRwBQ==
`protect END_PROTECTED
