`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WpGDV36mWaTqrz24SCcH0reJKZUCcsTKU/HwOISBRNwaGgjvxPWcAG3hmAfvko7f
o18A/uugiqkKn0jdAog1MMhZX5abmXl95xx+GpcUZLdYfuuo+7h3pB8dNcx+NdkW
qpDv4EuOZbz7w6Ef5a8OsTSN6p0eTRXE5vo5W/hyHr8cqdvnziZvLsV9Ws4gmo3l
b8M7G+1IEd1FrRYO6YPP2fF80WqABax1GD8klNTzYTXIHrKajgRSNFtPUIuTaJKo
kt3nfiWjnlwmCycUMO/NZ866plGqkUubGMHHv2bPv5o6tjuuvU6JG6iFQDnoyiUb
M4x1vViGSRgGT2UIAV++75dtrZqt2VLChVDePEQ0hbe/eAo50Bh8ck/HZqnGIvjR
MZ5Z8QBP9aES15AUQb6QPgy+WlE71B+WSN1dDYw8QRRG/siV8O2PbB8Ptss3IjFG
wjnDEdNMLrUfceu5mWrWSCj/OFArnXDJNdUlMZGTfci8rXRB78nUQrz+HopO7iNX
2Elm2I8T7dzs1mpNyNYDwxYt3SOa4mqc/wqjxwdh47vxptyzzB6AR8CNTPU8ap04
YXG/isEVLX1AInEhVu50uIAdv+1t4yGYMakeMKBKOA2TReYQI4T/nIQHcsi7fia4
QHh3vsLWjIhVsmSweJrN/m5WjCPXS6ibpn/36kluLlEwb+W3IrOu8Wjq4oK0z4+Z
FXri62JxqQWGwTyHkIVF52VqX9kUlUbc1zKGt/5bgVWU6nT+VBlA2qmP6WtGFBUU
+ks04yYorzQ7VjmUSwFJdA==
`protect END_PROTECTED
