`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2n+Wm9+gY4/4bQ161K13uJ5uuPify5uGs5BEKeape59F3J1v8Bt1nco+tH1+oPD6
Z315JCag49gQ/BIq8vuCYG5hxXgBwvEQj9CWt076uP9lyLf4feRRCz618STcUvpR
2RDajychBRG1PJDFsxzk+AnxouU7+69fjAhLX7oqw/EcIZtGrXv89BzlVYV6y4Ww
qerbB6bg7TWs2s2Y0STHDYGaLp1tC/uwJseIAdZHJVZhgjbzCY11vkAlhLruMibL
Hu6Iw2KiZL5k+opS9to24f8IC9ojdqQk2wIccFif1/9mhnShFQEWc6YoPzJcFfrN
13g9YALuyJplac720/1lGmtA4wXF1+QcMmcRyszOssMIV1/UG4OtSaB7fTZ3RPVp
yI1ufjgMl+/qwybQiWYtlglTvJrsKqHLdEnyjVpDv2eDmxvuGwRkH0cmQgGGFhG4
f91J5/gPd6nWNXeD/2NhAUBl96K/wAZmkfLyU90SmyW9S8sr/HxD7Ojm+9u6fNkd
uzSKuYkKUEgbUMOJQBnycV/03AVvETnnpU/uuAhTMJ+oaawxMTNAJHFMFydjMqKJ
qgT4qSkqwkt1XsMmtp2d+ZQLnrHK6JgOkGRv516E+zZKpiQ4EEywTaIQsqVN2TEZ
8Bt1RSq/l77VE4T6r594xw==
`protect END_PROTECTED
