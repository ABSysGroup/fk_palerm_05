`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EbBPsbpmi718eDe7Zaj6z9MRNaP70rX9h9ES93omrrrMl4wVOaXn/kiyErUaJsfE
1WXDpynI+jOplmFOrMr9DQhvh+raYBrzJkFBd2XYOQttpRAmiK8Cd2vTvDjwmKfk
pImrx+peNfyuuT+KqlHkBSYO42cWVuiihZtmQyddaDe96wabrDfAs4qfwhIgASTL
+HGJOpaPeCS3WVghVOmn+Q68dV1AMwy6p+beFw5WzEqz1zTqi9pvuzYtQd4YQpqG
m2Xn6qNbCuyEWSL4t8DIg+Ar9XEw7xZFa/fzllk6X24pfbCuikXRwlQDcCUqEOCj
gazjhBkmM/bol47b+2g7xA==
`protect END_PROTECTED
