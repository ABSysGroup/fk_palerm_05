`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gT5Llpq/8D+e0YB7QqbOUJE09yNvVwmCHuiNO5dMUBeAzf09dNr2dxrqBdqINZ0b
YT2gw2uN7LIdXQnSB57A5xKTAbRAfr6ECSwNZvT1vWvHjaaiwzgL/+5/BCFaC2OG
uRtESUc6h3P1mOGMLVLPuuX6mUbP4Z2mb9SxLpXI1uKqpM5pUrsErsCSalJcAgiB
4qWTIf7Cm94O4Gccac1CNY1i76w1SLlr6jjawdaMOaC0jYMK34NqTjpBeqf/HBDW
gjw/kNaju7Oh/rCI73vABEAsDZ0m7vgdI3J4vYzBCL3veMOpaM4R2mMpHjGFR7x4
t24Ypf0gSsgHCXb7tUQilQ==
`protect END_PROTECTED
