`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MDCIZLAGSAxIvDWsY/BoGHJFfMuijDQW8VqeRLD+3i6Nce446ipzgNSnqq6DPXxG
QXkzf7GJgJmgu9SysnOB4kVGIsyMvOTre2OUQALz3nV97yyPqP2W/vRS/N8h06A0
g6NK+hoUUvIsQJIhcGRxl98H6OQ1Sxyo6cogHuclt2yTTDTsFgScEy+5CWZkr/ae
nw2nNYnv4dMbYzf9985NbPZ+5ImxVt+1+tZO4ykfsJ69B25YC3ZSjhkV4JnJBoFG
CBgkOHkVtK9jFJFcLRxUZzdfuJyUJ3gGo0TSlyjwmRrbfNmFs/setQnHLt8w3opC
ZJYej7770Jwg5+udC3aSbwNcq/a6Guam2MDcEki6dok1JGUt5iSpg5XFmoblCToL
TqZXsiJUgF6HCpuboyfGeVnsVXbFGrjVdH7Ul5RZHE/ocFQSj3lVYdh2gR9qdOng
eTudkfqXokYb+lQmAsuSr5LXxOcJMTSca72TqdNp0BRHO1WjKe2nbQLOJksxEsMi
pM2n1qJsqUnh6vBW7k0NBFcFRycqvDEFqMrJLlfjUzzwymNo8wOI/yVrUx6gOmWO
N9sGul1ll6x23Piz6tHl4MbC3+3AqiJXcr4vOHJfdmXjVmB1W4ZRFeqE3gV50HT5
pwkqDPUg3tfb9Jrq/sNE+0ZaYxlMecznwRl8yCDOX8QXSNDAcPZSpIdSvRlTR+SL
I25okoz+b/eMrIclEkyuSmBjh2SjT3WUFe7a0TrVSsdVoR2h4AITPxq8PePYZTN3
8n91xyWlh1UPCLMZlju3RhwGNbtDyWZYgyYFId0rzetyYmwWCY1s80EaeOSQsCLb
oY5tCKmkxDgIyFEqWrVGFTpH3TkNtnqDG2tc5dPs80RcdpshiMh5S9qC8S3UU8VH
B6Bb8L+yIJzMAKMgr7qRQtYXepPy3ruyOpE1t8GvJ7vNL8d2yKyOHago8Vy4PiNc
`protect END_PROTECTED
