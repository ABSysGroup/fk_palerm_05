`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k92IIRveAH3HKiDiQnstLy8ixGQJj7h7hUgCOaw3p9dAMUXQkIuuSdmUZB3mlHsn
DRxnODFMfSX93Peem8i2z4c/GPUvoh3bcPf0MXODqdeKlj/6QKMyIh2Ax7CUezHH
UkWV/HmFFuf/ALTv7la8sAF0WmqJ7vKnre0GN+BnHDeFGf38ckc332qK7UUgEo6j
dqrX5m/OMb1GVe5H7KBfDx2bobqCjVXT6s/zbsVGRH8XZUVeABzI315B1WgrVwqh
iil6SEw7xaFLHVFsXfsCGw==
`protect END_PROTECTED
