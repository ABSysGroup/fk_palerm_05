`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
evRSLJHjW8ojEIkRwyMBhZGTkqgQBTzSRDmYKB5T9XkAbS4Y761G/iMhPi/M847+
G5ZNE4+aJeX4dMbosBPPjjGzecfRxs9ZdO38017s8LsVjJkoqDuay91iN4rCtQbr
FeY9A856ABOdiPFRpWL9uROh95JUMxsdXtIOglBe08a528AeSbMslzv/7JMkvzbA
ZXDNBn4bcBU8eqOLyDFORS8oxe8mCMbfq11iTnw8Pfy4CMClRzGakBpmWNGgo6VH
nKq6mzYTX4PrZYvgRLqQsxrU1UjwXugz9PqwsMi5ESXywMa190HOEZPlVCEHc1SU
quwQutl0HPlvD8zQmbyUs5A5uQEh+eWtGOv/gnYfjajPDNPoBYtIM57Qd80ynedl
ujvrsDKQgYvRbAWkrFa9H9p1ygbsDSEN4jpUvtCSdwZgIPNeUi7WMcMsGGZ0va8M
nAlGfQdVEfrX54+sLGpY1WpLIHj8bMrJ4IaG2chjTzcy/R4xBe4C/xG4BOhmCUBd
zzHk8Mcq67nXtRKjcLLefvOTl+QTcZi7JQc7uT1F3YZGspeXbjIibWgeKgUsDAC9
lo1PKIBjPRJ8He72sCeo4JynbmB6Hz2XfDoO20vEmEsAnBu7KcVlLSODco7SzwCn
cIzHB4wTivV/gdmaWv/hmkLDTNTxV7Y07hAyWjZUNmhlWySnHovdwfStVJk/SHfL
igFIpqaOfSgB9KZRpWJXBs6wbmXOA3trEbpnk6FTVSOyZU7YYs56Z6gFIU1vbRnY
egS6sDxr3MWXWW9KFQrfaIwZ4mTknbz5mnT6Pw7MbmAClloIQgsbtQLyJbEX8bm3
gr1TcTOmc2MLj99qNFS7VlJkOKJ5aWPpI9GAUoaI5zG5hiPyLNST84zWSXYFbQBT
aRmm3seiTIyousb6is5yeQGgjoWVvi2kOo4szaGTLnvcVR2vfLSi3+iFhdP9Tz73
FmARNgnscIUU0Q5EdBdouRSNLvEl+Wx49cDnnWnK7ZhGxDE6kmg7XZs1JvOVNOWo
dyOwVW729NW1q5Ic8vZzmktb+OYzDiTv0DJ35tcQcnjgRhNQ4gx81hbsyaqcVP76
aXkB6ZIcMiPT2HevwfEqh65oJywcAhMW1Vi8KO0bHpdjNnVcak7rOlCXikdr4ynf
sYCJFKS+2hz5lvqeZ8C6F2+UQVj5rTP63MrjqeSu9Kqyk/kpPsHULOrGQYdBxIkD
Ibk10kWhN9gPOJJMaWFUdNlZT8pcuoBUJOzamGoNMIX4W5rI3QfTVQwXgFehQ1i7
6o2yzrjgZuioWk7kdFt9k996M1ftSi2fhN7CaxdNoDGUZ1Wq5o9dJeZ2+zNrI8jE
jOYq9iuO9qxAOntYbUftRCkHe1lvYjcatoQmmK+pJRdFON4jixKhjCCvcBpiFzNF
xN+Vnb72TGpGpq9V87z/tMmpxDrG1DSlGCaGh1ZWtsj7Y8GeFcKEvEXTqhYBgB2R
JN3glIspqtm9UGmBBzHZ2aRrD1u2dJ+bT5+txrnnoZoQg3dzoz6sdIomWg2rx391
4jPjnZs0OWWET9ICDeiOKVBP3bT3h53qrHiP7uBfm9ZWqlHDZ2kOzzBNIxHyk2z4
ivODXjZAgsrD/Lf+GSyf4sclPsN017lW6CjoDlN7eIDKrVuFKN1NVB2gSFrcZWAl
lFL/oDSgGOLzgESC8UA30W1q4liq1TEWvCzBMi3Xj+E27+TxuJBqp8/zIkWzPt6v
Q+x8dOeKZcuoY2wGqlVn5rEsqn6aez8PHPJ9DoYgIPu829vQYZixTUp1GFPRyaps
atcO4otlnedzrlLdCI0a4iszqUv4tkabHMmLddb2Gr1ypcVocFT9/hcoSARLA61J
H1z0miSQ2QRnWbKl0Ol/jT2zRPLcFCx4k/5GHmRgDy88UXER1w4/8gZj997y/SSf
26owK9kaRTdr2K3comufA4xFIflXlG0X6DAolPbRvj9U+xBXtLUC7RLzbc+ybF9B
n0avACPUPCGeWnL7WonUesOvYYHyUDSNd+yWiVvcGVQXDQxczPQOOjkGfzVSB40t
WRLPfD2HY18rWH/nCmJVPfAV81mf3G3muKY6NXmg4JIWyfoabyGU9WlWVg4Cqvyj
CWsQ4vFOdQG62/IqKdOHLDR3jVmAvKZF9oUpTQcQ49+xe3IizsQCZQwAbUMPRTi8
yJbkwT9G0ZdeZyXEYLF1giARb7wjaeGVfrvbw23BHyFL3A+QmNHy0+eVrk/IXlj1
UPMYs0s81+48SAMQgGlgysKgugbVD3tTw8BoCVCXm+2+FosFct2GsrWfpC5qK/ra
MoNC78cwDh0UfP/SYEg+/8/6aZDtCHMeRpzMg5AHqguxgPl3XlVMxAsJJyVne5EQ
yl1PR7dQ4tKbMmQUeg81K+kqbKT6t3vwWAHQD2UvPFhanAJicWGN1ybuADnrVYRF
wbczXhKWyUaOXzMGedqqqDcPRXK4YWqYt7wjipPFiV6seCNZxJSsvkaPcpAhb3uS
Wm7CTd52gWmD5OBwkywsaCwNtSMCW/XlPFCCUjsCJJTmub5Kx4H7Vt1Minf1wHkU
GmNRtcmAUcATtHvt/RNq96u2HOKD2LgMfNA+HFM13m7fa9hRub+NTx+pe03Foyj0
3jG9J52pMiBRxe2yJWOVgtAXk/UwWMGbIM2job9YFD88ECL2Y6jiC8V5ULCz4Mjt
Gc8iwEwKr0OEy/sbaLTzuHvbRoT6Rb0mTAHHC+DbL+CvZLIhT5tYYbdBwMrvSUDZ
LwPjLWDu7ePx25Z3xmHRyBREp0WI1Vd8H3GywogZgPqpmHA/xBuiRpwAzIey6MNi
Ig+ARSFSzQ11O2PixNbdUapGYpZOar9YgFzpgqNOdh+QS0OXmxfc5yp4bwhzIsIf
JdUc9oYwrS8hGC9Ba7/wBNifcOCYvxQSfDIcLJRZbe9EF4pKXJtK6my/OiEj6kBJ
rLRiBmlg+imbDjCDN/qPsXs6IsBP325F57KpDzpgEqq4zGbVeOH0LIF+gpa3nLfe
GMKV3vo/XcmNxnvaKycpuLgKglSeCmFq9O8v4neP1rwdu0YO+7iKwaXvZKoVRtaj
LGX4bDR8OegE1Ymgywgha8vslx9HY87Nn3rrssTh5GCLBbjhFSHhd9G5oumYBqK9
uwz5AEejIvVuozuht/Qez079NM2LTduK7NvUKUq+nRQcHTAE0jGzVaCWPEsZzdbQ
kGxiLNnl+BIv666Z6mxqEvXe+jhx634b4vq2BwdBkA0sVr8dPhAZh1fKSP0eOYj5
ctsz+ElvBmazKGceY4xyJr8KN13kqzj1KyQTCP+oyNeJlHyipKabRf3aDlICkvfo
94wjpmLWfuG58ZTn9yWZt0AfPylGHtAGQcNsGE7G6KsHSdWk0wFA5TdvX2UDcvkU
mfmMCfmPBOEeAzmH5BfAf096gvuSTLcp25pHGcznQ+KjEHUezZ+fFjzgLk0jMXAQ
2aEmRAKDcA0eQWvGJAenKfl327nUd1ZBW5ADAVKvUSR8NQV26uMLXBVfpcHqJs18
B8OcYIJ/WSw0EJd7pgfwFpE80bzIMC6n/464jyj93Fx0HqXp4m23dPohRlZMcQS8
cTbBP8PPkh4+rKzadHQXNWENnDoLRs8xE6dpBxbiSsk4pzcL/RBFQDYpiaxQrHIH
whBVNycWIWl3ttYR+ByTUOsSZwQGbu0RCApqtIHPnTCfN5ctvBd5GF6ZmgIrM+VV
FaRvDd3r7YiiB10PaJXBYJQo1QZaVEISP2V7w5MzLAgDBj72Q1xv+oS4yxN8BEGJ
RET26T0yOlRYBJKjEdovFOJxLRVSDnN5UJZKTCH8So+Bwcn2mjFLWWhQwevGg5+p
tJcik8p1EgdnX95+isMyS1JxskWEa/O2ZmLKNp3yuu6Kh4s0WS4fh6Ftw4Z8j16+
TdAXSJswv0Xn9tFypAiPFb2ca1y8Y2MomvevEwDiR0tfn+ANSrjmnG1Aa+yAa2ff
hLR+023O53jgZwbpjCK7oCVFzdkid5Z0UbN9qN58VmaebrrO23p33M79dkomEjMu
jgyOtqw5UHJ4YOx9F1mLSAcefS9wqlKRhly0Pgwlc8+39dokIL7AQIerdFv7MC/P
+XV8UlJuv9A4zrNu8RBjAkOvOKl1x2SN7F3vylvpk9pGukJd8WNF44h+5mmW6O5r
547taDrOQvZvKw3/Qp/U7RVSxvPashrPUuPJPTJvYjihggAtxtd0jRKQW8XswA2a
Bh7r8fwm8KdBnTcqu3EJDWKNRJ9U1bHycw8ux5KWEuXl1/SglfjJOBLrk3bU5fHT
a9OiJnKK0hamEnmVwt5zAbWkbZglWDzb95AmQC+xzSA6xP6FCib8NPNawc5ylS45
8rKW86qlDngKSAJtu0EG3jBuHkHdAgeOnH9xJeOcgNGfEmrQtGOzeaOPN5+mAKUF
z6ZsTwwuvDSenBjDyVyh/h+4SWedZePip074Bbm1Z20JYvDIAfmEE56nDGs9szIq
UUyItfDBogwIMLJKTgmZUcjeNk3n9Ar5hN/TzYnRKv2cPp5cMBn561m3OrMNa828
S/Rk23r+4vyz70PUQg5O18W9ZVA0HyVSCw46Ubn//tZrmPnaI3rrMnPFOBA9kbmt
sF53ABh6mMK8M7MpC322v03L5JtAQwyAMahx0o9N5mx43NrJHakyHO2dE0TA93EY
pZR3dYSwjny4sv+NePsBXyNAfQFljTfd4xIWYHF4jbT53Vdq2Ff/7yla/2oWx5+J
AYYBbj0PYetLlbhCpYYpzDENc6NsdV9Ie7cxO4m6mUsLKSkGEucioCMW2YDOCN1/
vHqc6KVJq+MwWfPhFmx0wO2knsqy9LJR0y689kTaQFGyVP3wiY7dZP8+DRbrz2Ka
w9LwC+F9p9C4YXha3WKxFSDZt8WGh5CwWuAUIGmnSwf2gZd4NFRKckkXCggDQAi2
NznOgq4UaCTRhFiFgZNsyhTOOEfeLw3ZhoZDo4Dd588otuxgVFKnp38GnlCiv/xN
EXhMtqiYRt9Ud1s4Bs7fm25Wc8h1qUo+gplKizLLDfuMp6Gotf9Z+zFFlpJOvMo+
0yrmdmYbAUfHOOSCA56vZKuXKhaXDcTU9l5QjWcsfk++iZZL7hGEEI9NVR//P6u0
LBuizUo+eLECioP/oIuk/FN/Qk6HLCMEakit4JshsgpTImDNSTqePX1+h1xg29xx
lgf00HYsOKOsm2qbNQWvP4P5lKqTcN5Qq2lxQu31f6g2/oHynOncVV2yjhdVblUf
ZdKFFfbdu29ZHsqU7iLT43ZAlkS0cb43poiPv+TmyCT9UZbsdmCwRtlZPVW2H1ao
qHMh3i5pzNsApk9zEksCMTdiH/KTK9i3iCDqQyg6ubvfipYmYvOpLN/FhJcksKsJ
JkeTS4cdyKokhBP6icH08FqSUuSBcjz601dtkistT1qcebDRdb6+cXOZbItpchN/
J5/a1L8fRLGxaRQavnLiTro3+Vvn1espSUPuutCX8KY0CrQT0/hwGDlkXlID8M35
VR2xnyre9LpLE1eZ0uN8fWMbKibUB6C+4v36JeDoOwCzXs+kZHVg6MmxpOaRi8ay
/dlx8j8MNYNoHtFBlZoeBHUUKTI6ZncwzrESBci0euJDei0l7Gkqiopwo8AAs3hh
4JB2Y9bdg2hFnUX3aj5aqi+v2OUctI42sa/NZmLQCHmcXIMUbY/TeZu/GuHTpJA4
15htWMR33us8LBu5ID21kgC/yrlxhA8HIJdOUvJ68TGN1NLqtSKrXbF30Z3DzE+1
VEzqw/yYNrMsEvqPmOTBP7chMEN6GxYtyj1RUlzhoSFPg1YC88L/oa8vlvkcduXp
H78KNlxmXPA2+CtZ57NPJJ69/3hTiTrMoVLuO7FgYsUBZq44q17BEjRDBGbd0j0W
Nqki1hQypTIZemuAtcZ/e1y18fC44C5SKDxUQ+jhBcimxv1yO7gol+XlWF2TgN2m
1O0z6fxcuLCfR3sf7g6p1qhyjV99LqeELxpX20Zb/FsyArZ6Gk6tGLNvEnCW6o0u
VnGDQwI49FH0zFBrDU0tMtSQw5+kBGdMz3DJABmHwB0FqgJEE5L1Crn2oBM/CmiK
LRjIXpHOCMMZQC+Vn23jPzxtuWwRPHkiwSWP5HcJfCxlLaECMEpyZui2hN4b3vCI
SiMOc5ZrWE22oH/cyldlrGJspf/UBpKZ8S5NXr9jDHaKK2IP2q8tYuso826WdFsF
tCKnBJPpoa6F5+wsYZeD8obSG1IIT+ZJ80D/Xi3IyBxq2TVi94i7pfAxwNhEeUb3
93aUk4aTZsYbQsgkfVN5Zc7v24weYB1ZkUlo5aT4o/QelykDPVcYpfsXoy0KwTi/
6OTyhdsfO6NWP4B8YNqH7hUSLmO00/j/sJcr494eWxKqEc+8IHi6Ny5ts9CKidpD
ilnBBfMmOo2p4Fp4X3+KjCV1/nwHdXrSihlkB7BXuwfZfvrimZSmDpSoiLjtCN33
9/zT1H2VoR1J/ZBtjltk0BaS9WhTp0rF/ODHQyOGUzTl6IxSM7e6pZW/KDAg86Qu
bUt+8tJ0lIe+JhCXUGLJsj4o28j/aUD5ZrgJijAhez+AxRfYTJmXe7Aifh+A0EKA
TfLNyYHpLnieI3igD5Eab184T15wp5MkU3eDi7YxcwAPKNQTLKd3mrCp5dBjt9Ls
BxxDJmby6TlLmO07FC8Q8bF0TpCIPF9iPPm6Q5eGKqZM7ov28pvdTpRW1M/6TN7I
1O63j5runz0F61ttMeoZiE9Sm6VsEdpBF7lNpriVpJZbW+SF3Gze4N6pNPAu7y93
OH2RCR6gLB5ndkK0CH9m1++CCnFF/nCOtt+FGwLYu+MjsdDXA0p0SOZfTUr7+mmv
vAabySudPs49HvEFFqasuasBHTL/K0tNMrsFPO6Tk8ippy+tdHBYeyI+pgJ/ZJPM
r5RdgUzvSUTzKqc1CfeqwebxiFP1IRz54tOaYPR2ccWb0iPyQDpY0XiCzrSM+tD6
UUkpYGkFG2b26vffLISPFtjDfDcMTKIq6OevxrD6IOV8YJfI1z/zxqLBowtZ4Y6d
aaPMi0ZsOVb3/RM72BQHuNutSbLoHkgn7ABmhSHiTkXJEtrAlJWiXXSpxFy1Axg1
ajgeIRWuTt8MIuNViRAIhtiqLyiiDoAAk0i6TZtF5Kf91rWHNnbCTi1wZdfPxQLF
iqYgg5WluOZD/dVojVezUPTw/dZbwv6WBeC408+1BzfpjyM93ymMhUCKYTQN6k4g
w1FcSI3gNVlK7Kjxo7IKOKR+n5LsDOlN1oXVh+S/HN2OujXQRwf34SzE5Fpv3tRh
Yqh8qj8l3YwmGuk72+xvXWAvj+n/azc5naTRWOAAXPi9x6v1WzR5ZqwVEYNXWFYJ
BWmauSzO5sAAecjaLFslKmGaPoO5UPmrLc5KsOr18Z4U+vkEcZqnevwCdfKbC/K/
E6BwSlEHBIs2J8PKiFM8Usw4FbKLV4fxza2wiMoCKvyj/LhxK+stZH7BJSD0N7Er
zsr/zVoJ4qjFoLU1PeSqXOB/nnzzQrywJsOFqQvu7ZxeWmf9iPrhmH2f+dRmtiaL
cjqW75RhunPyYRgzVQEywS9KTZ3W/4OMNh1T+rRoME3ahiDNuWVCJnTalHBCqzb5
u1knmwEUJVPgQzS1Ykr0hXGhXnEEiWT7mycBwRY5pc6o/xLuH5j9cRaGkOdPtV7m
5xhurH0fC+YcOHp0ob5Rzgx1brlnfSaeNCYGUSImPPCdzrX/fGizxoRaDaYMDGZk
mMaJwNH6Dk3ySvAjBZsmhw0AGykFCWqX23DqxyFHTafOx4FbS4mu6CONTGGuRQK1
sx/zmtNXDMnDuzL7EzwmLTuqwFdWlsNM1ON3wlben60vXI+VV+C+zP5b8OildOMY
NA5RwDBAtAtOvEdoeBHWHZ55DjxPpcS2jQCElpkp+re4uik3n/C21urmr0lsYZ8F
6lzB6DpRKDzg1pdf4EyBZevC+K/9ePDFLvJSyLvB/CnnH10CXEx+VZeqMxCCj8fM
YHg1DUqRr22Ht1OD/vcerHxZ+8KiU3ZsnxEovxTtn47UA+Q4kY3oM2mETY2W70Lm
Ltp+yV5cmHE97rYF5kbE96foo/3Ab06pkt17rca9xxAZsS+nxDK2NIOW5fxcbVWt
TwUFUxEFsVtKiFQn66KOsn2WlpbbSgGmVAeEsddP8aaRTvHxwLNyItoGQdTx3Fpk
m/zxvbKOj6yGr7Ny88zrnOqSyxIaAprZg9oOA4XRiJ9kE9opj0+qB8/VKAR4J9fw
2hvNT/Ge5855AKbDs9uuHGbmSHLMTXZ/7fVs9STrwLr2097P+5qEdVAwAjdyLUte
N8bFIsNYBIfII/gQ4cLr6LmRwu8fweID9MvC+v8di+0=
`protect END_PROTECTED
