`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
docuNOksWjQJJthHGwcTMu0Pmwtc//mYtNlrYeQsu9Tz5S9jU4qE5CRnbTSTXCt+
t59K79Xq5S9ggs3uSdhkqC7AcXIALYmc4rKrohHOWgjohdq/N2lyGKmyyIg2ecFc
mvS6H49C/PjDpp1l2kIrGDIgEeveSMkx1kcfuTn+GwzsKnNTMAcZNdptMNWuSyat
0sbOlfeuR57vy1xNCR0I8pSCx5hEjkdLY5Qlk7bQ5AC+VQoLkvRoSehCgcj9BI7x
zZAIoegFV0sb4MLfNIg26DGA5SXCS5zs2FrmfbWCM+mWcYU9hCJ+LoLd1zLm6xhy
AvYLiG5uUM0yo4hSJRZBldlQ2+/jVqorWs6HU/ysok+zfmJ93yieT76Oo+R7IdmH
E3mxGgjVNKrhwsMWWI2DJqDmrNE2e68sAAwNiA3MsZoSBycEu266wIlNiXaD6LUX
y6UC8r+GQFKc6B1oOPq8UMSTel00j0P2r660EoPVqo9bJseB4orudSDKQ2nNkEkt
UgSvralvrlVAmN3ylMqhw9bGdBtZzJ1MZ4KCxtDTBRycHTAGI0DL7+JkDG5LHjSI
xXCasHCy9xksJ17Ll8XIQbCLSQErBqtuJ4kcKF0Ti3riKuuYNk13nFa6y1hRI33j
dRBCuBQfco5pWZn27H3ncbbYviWAYR+NTYxTu+i+nTnB6kA+GXcLb0AuUjynY1V+
Za2Q8AEsUKLUprk2Op7C2sbgdqcSgSY5GntxZfUb/9XgRadhValCeLlo9PV+AuEl
0FTSgXWFsrRoSpZRN7xE5q88E4UVbpOzOCib27lGcaJWOYUiKEDjnSgvD3NFq5cP
TrkYtYvSxZudQjB5QfHNMc17feDmC5yq9/QbcJggsrtJLA+l3nT97+oCd5ThMQm8
H2XKzBuNfFtcy+oR5w75QSJ+3Z5U9pCTnc9sSMVg5+pt4oBiVbBYDOUUwu3QtgqL
ovAQp1FtKL7IfmvCNeI+NKs3551pfRBWFM15TF/wBhVHZSpVWf5oI10a0SwgUTff
6sJdQBdr2QGBe7we7RQ3p7qqZhSaqjC8KvObPrdsMrYEBwzJiWi+1ebUkyWGsHLx
d29dyByX4TS7AEW5e9UPrKEpaKwvc6QTGFDRkvZHrcFbz1X/jX2I4yDMVP1pn/84
8pJ/uRNzBj9KIalIY36+Pke8t8fCnZHuQPzK7x5fCea1dyuLURrRr5i0lVl+1f5Z
dS9H+EmUgDUtKss2IvDuwT3T6gztBhWnBABFWziAn3c5pu6eBNBhWsEcdO0rsVdF
eJRyiYUAcHAEoJOAvOLZIiPxV52LIhO+uHvRRcyjmJPqUbj5yDJFHvUxAgqDVtvM
CVCVJCMvYNErrXn/eMcmwMUTR8l4jLHMdc0TpBxyLywCayPY38D3+7W1L0vE3361
+G+SZAhcNSqwuwus5zanO1PO+DKy9+5kfLQASJ02WBW9k0v9LNLUOdNVoQWsgyEx
+8ue5Z+EdDa4wqFJA8j5SAA77FhZMshlkzVWxuUmwkIPHzC/EHSxm/0Yy/9oyyTO
nfv4KaeViJ3+jSxB8PoOi5HEWzvzr1Wt8qWMuPjeKELLRmjJ8tvgrdc+ed66WwKj
uXWV3BZPop1siNDWBoeMfFnChKpooVKlfEzYTXt7MhwbVH96uK4YILU3gk367hFW
bJ2WWUOxgr8RIeW5Gu2dbpxLEWI01r8bSjQGzNUSDAOcPvKbInpkQnAze6jiafxU
Emn+REWbDJ3QBthmfV4V+gUr1hBl3lITiNEcEzcdm/+H/CoI+kVIX7McaHI/lDU+
i1KcisTarjLSXSFVSBeLHHtUm2GqSc7M9Ikyf+O4Jy/pdR7mv42QDhclIbl/JgLA
RxQpmBXGjDJpwqa7OsZ2Ra3QQ7ZmBjWCuxJaiV0sYVb7J4ueY6IVgYhT0/nLAOc4
pkH7w0bNVpfPQVpe0oPvNu+fnkRezLwnq7tcxXhgnHXyLX7PhUksQP+fbyU4PLFM
VWlr4nLw2nSST6mCv9UN3lqIGbCGn8omufdRw5DK/hrfmrzP9O3R3u8dLRtqTqbN
101S8NKe4KtKqgaNwwNNNsCd2Si+us7RJqHQ0vI4dmphf1XlooppaqvMP6RA/1zM
tCDiNi6GrQrOqWuHNsSKiS/Kv2gDXTFxxvVmFyHtlBVeJOW3vy83pimauNiuufKo
zfJO+lIPWcCD/ZLrU25GIWuQ7FX7rJbNM/oraM3ewWwdqt5QiJq8oEdiKFUi1C/m
mJ9QWLkSp+U+0vn2V/XbwXK4l23AxSd4hBBlrqZsiCK3gtcz4+B9IWlzYjuvcHPP
6o4qHD5FCaefSjXWw1DqlZnWBR28Rn8wGrj7AwNu17bJZ2sQ5qeYKnQmeOMFDffG
GYqIz1ZBICAkLWPfdICQwqBYiaiGIXf1pNgEpRLqxE8BdKUmLur8hKnBitEf2XAt
yUlYm85mRUNsPPJBSfojLbd6nu7YTRSqK1hs1BWldgr5OMMtJf6pfYhoVHIlF2ZR
zDZw7+YGm1P7DZu1TZhk2XCVMGRHpFFkDwPH3NXZ1M8BNYrkroBHTV/IDr0l3fw1
lWJ2nGafWhEEW3ubRf2Jx8265AKPKFNrSsKpWJJVSww+kOGpGeaEGZhAHM/dH89r
wVCCy+Ttg0yfkDRhXOOhXx9TQCn2s8TcjFO/9hu57sSMJ1ngG15G8iUYrwjHtf6O
we0gWm8tEbz9+KDXC1sS6fbTleaa1ppHBCTHBfEgPikn3yELiNovbs+WsrmiIERf
faQOJhHgn1t74oNxaPvjW6D7InUx+dLTfiMEvEkWPOt+2rGWUCuwuz0l3QNzq2ez
zCR0YejwfuZt5PMf4KTzYFOU5CUAQalhQHSzNaBdhGx7THUmT7I4pyS74os9TMut
e/qTEiQSm/mXguNX9pOvrLnAynD5VOHmuUXYeaEtrf5FOxp04Q//fDO0VXVqkZTb
UaCMqdNiuzbg6QFTwYeaA/soJIJLZEljoeVM0HOECvrkaMgkv0k3x3xDNDKIet6U
B6cWOTy4PZrf5CPsg7ILd2AtbX+OtarkePuW64/UHZ/YQsR/loY/Mffpg52gVhj0
iXb1lsPotaq7Muo1J42uNM/+n0RGXVhZQPzerGQgL7pOWAS0u6xY3vzH+Mt9KpJm
F3argQdfL+KjYHF7gPjHOT+0SJpTcec94rAP4wjeaWARKtrv2guG/9ZR/O2cu7b2
SPYuWEQpf4pSWbnMwkgbnq8ak05JUEBUvzt+caHnB82+zsBw+saB+UNCHN2mwWqE
5gsoLy4CL7NeFy8EBm78RZdRPxTFsDLslpPiltZKZVPlR746KSadPNYBopLfL1v4
gwGvw92UfRmmkDDb4f0sXrnoErivg+qI8tfEICG83bnZkyA13AL7nIBLVKyXytRQ
M8iKBiC/sgxXkikkZGF2g3ueUbTkBE/YZMF6YeUYX+CfAOyFVOQIpzddGLieko/s
TzUfqZnof17BOq/CbI0ERuRGcRPjuSLrRCchgl4sB+9Wj5MD+maa1khLuZ3yKCQz
+Z0uhVz7YWBwTOcCtOT16r2qHy+grNDDJ0eXw+sUNVzuTcYYKNL/ZgUeJw61fpZT
jqwyXNYzyFDHWPKrNZIYOHUr4fFOo3e42ttBwAuow2tZmkMX9KypcF9r/r4n7kN+
+YFeGq8hsjezD8vqOiZBz/IJApZngu5sTigLM7/P1xfMKNHreJSF2WPPRDH/NRfo
qtgIeztY7GR9VbH2Pjli9N9yNcsUUqncnU1c6afgPegDg1WyELvgv5O+Ub66k2Ls
gGOYukBlRXJ6ZoJdNwBatooamQsZdQmiZ+Eld5KBxcCultzHliswaLshMzipJJkE
M8r4hSEahEdz/4ZYFSgBFWXlOayHJ+dWZLzNYASXPUHCbP8jd1LGiLXlCwHWJACl
yIbfR6SEDORRCpyBZqscxnvuzLv/aJsOMEiKAywPRm7YkSP+/Mw8VbazaOH+X9O+
5q9Nu8ICqXllOl5AQV3nUdiQrDK4Ph0UtaTlCGz63kdHieBEuIhoETPNZh4jAj7L
7IOwDL7Ws4o9EMvS3wSHW7ghpK96UCE9g4cgbiwS6tnMW+NWEEDf3DUGAfaaYZn5
/NuQp5wYekcgShSHQMf8Dwg4oeSv+iTnpS8rF2hJOiN/Pq7GGljQe6l/74muVlhJ
7GbYmLqddKjZvgOR5kb0z9S+lDSoSbhOEIptSBIE6BLVALF1by/di2Ge1pH4PFd/
4bo6nYgCnDrILLBZXhEFLuiX+++6+iOYNOL3Mtin50myQLzFc7rNtnBs39O1lJuY
oZI0B7WabI8zglWNJCnuXhW3qNSwiV+XBWwzfIwzdCtecQpg1YsWFF3l9MmTxSuB
Z737Z1LBHGZGYV5EcIxUSUeK4nQzouq5FRtvd6KcvJvgJsoQGcpP1S4cFV3gw5fT
EgwXdze6Fw8xg1dPvbxpTbU8Rwx/R/FpRh/emiiPso2VwIM8mkiEw9s+JUvWzUfI
KNJQjZ3RQgy4VqM45gNmwB2gAn4R6KhfmIZ2dnE1vG32lcMYa8GkKAHRNiMxF+F8
bS3A6V6xLUBqQaqSWOnNAYLX2rO/HHb9kyecJz1j8Q0PMdjx0WzOMKXJyT4OIY/6
YDzYPOFD3bB/itUwlL06zrQEcSUt1E79smUt+a9JH3JQ6jvWQ1m2Dv2Q2NZWSm7e
tgiCI6gkKwDr+F9zDKWZ3YgVk0FkYSbwIatx7UkjbZ4=
`protect END_PROTECTED
