`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lUZxdR85IZxQoMdYMAaaBTfU+v8brYsuaTWDqLDeRldl6aWEqfc6bczbPi5T7m4D
GGX0/cUQt6A+hIlNK2mBH/wdB0Nd3kUXfVkgKaWnYL/fOrPB9TdhgpjmdeugKXI4
/u5SUtaY8KgbZJRP2iXJOetB0aTkv+dFSxu8aCir7PilaY6tzcQIXKNxr2RPPQfR
H+LXzhaIlRw7k3anHcqoiXZin+GzOYwi8Wg8R6MbjUQC1MgqIwwXntcAebpCissJ
qiuszPqB2j0SjsKNs20lvNXO9T+h64H6UlPAizofQUuux+rlHzlBPvVFubcXpyQ6
INr4MsZkP1CTy70C0EeYMrmr2zV+tIMA9GDBPqFtcraP4gJ1xhymIqUkFtUOomPq
yvRWaqnWUqf7sRTp4mu40fEODdXyjIZHpXg1SpQMddW2p/2Y2gU4V/V8wr6Z4en+
xaBklTMu0Q2udYO1VJPWGDUrC+cnwfQ26e4TuvtEXxJQR9xqCYiAU66C7kL3n7o1
1zAfCSZ/t0aYo8fKf7UmGsGIHWMb6XoT0HXPmQV7FUXq7D/RPsxPVeqET3G6sT/L
TdG2cI6O12NV6KYmzj4uOjCXDp/XEXTK+FZPDcjVJG99sWAbW7PUZuU1mEoDiZMj
yia2xzZzcJRKkOYdkgcNIJTEYX7nP8s56DV4/LLMH0sjUctBEfsPoU6hO+t96UFo
cSTOy4mvpKUzgC5HY3JPHpiFeU8PVFu3hEk53VSShfsoNdy9mDT1CiZ7IOC5BMze
IaeCTEyutrf8X24xzFhYqO2pS5qs6dVvQeG3cSX3O40yMn2jYLjgQYPcx+hF8aSZ
/+vpM0XY1jiZPalhIAauwRbI/aYuTxmdOTRQ4d0RIrkeUp2/egKEFdXDJz/BwLkG
iDCbZz45LP1vAK6lCGJmuPR0adwaY3Oyfu0qD3E2spWdvuF7u4pQ3f7DKLdRfMUr
VqwafEUr5J8/3u3HFXn5f5nIsnxHVMVRILlfR+9FMahIur2O9wRdYBSltg+Wd8aH
ZZng+jm2PLyhy2X1bK5rJ8QUOJs0T0QPco/+Q3hnZYxs19qMP5CYAeCb8qXmHVcy
ebhwKSehmpEP8J5NAn21R9wC/m85MXb10biHL3WuZ6oivD19kqsg2TcPidco5wB2
2LduhcCaFG3W2iuv+eobj6B0p6QRTLXXiKXZmJWiLdvDce7FUxOkMgcNQc/MbVXx
Sisg02VuztGmEwX6V4mwBNaBiiDpb9RlH+qXWbPRMPYJGt40Yl+ZNq4gHGf1HXz8
v0xaTjnb/rPspGzD6GCMocBe+iQW+uT+UnASSIU15IDKLvYFtz2POgE4pZ3ofclr
jIsedwFzYSyftnHfefW68T2WLuQmH4Mj0iG6LbSpqrMtDPW5RfMJIXJxYOWppzTC
5pwABmHFPPf29EWez9x5um6xFqDXjKyc8hFyV+PwAqRcAm5h12RQCCL7Sm9pIswI
qdANQ2UZslhNkKb3vFEHxnJMaGfVDrgd6+qY0081vzZfmJ8TxKiaDWxaIfraJVgU
JZMVv8TVOq+skThZSRdwp32UDVNeHlLdqA2kGksqeHAmzBHuin62i/f8wyYEThyn
OhOvZHBOep18W/ScIxTtp3PAsXexK3rm0e28ywoIL1ydfMGymY2Qy09L6QBtGBbt
TwrfeOiPIyQeXaKrSih3hDLmLi0DDnls6Cfag1kz+EkOyoPxFrFks4510xATWlvU
4CLS8Qx/lzVJphUIVd0y5v5L7wq//Nk2Pf1rLq1t2rTfPGflBSFw79mL2TBGpzy+
wJtMbMaa0TuKzvNXyqdVgNGjG0UpXQvPIzY811MqMKuCCukhTpKQ0oVIto+ZFFwm
p6e0CV+vL58jHCleFJ4EJjVBxKbYd7PW9MyXWW5GEZvjPEJZvo7T3yHW7Yxcyobt
Gm/p6d6Ka3PtGm++6ovLrNnvqOvDKQQBT7+CeRC+6vi/YIW+aPig9ONmbDrnnMGR
U4g2kbzVg2SCBb+k1kgjTYtyio7duhhgy0hIE1ek4viR2wItqgDukQZGnpU3L+fX
w8cVUnYrBy9x8DVgm02d3OqzNV8QxHUsAT4CTa/ofzB3x9rhpdzNGC72kCqxWP4z
hxXmnQvSKK04YqE1di+/Dmx0YIEp6QNqqHDRC+fhSrXMqeyetd1xyc4qf0GOzqhm
1+TvvBCkeitzv/DGvevwOoW4pS3rw1v0ZmwkLG4nHLVWWi1ImOxSWpE91hpJ1yLa
h/VdYXddujFKfrwfVsyQdogIgHImn5kkGHkhvyysUQrdsgBdxVvXaK7C4ASUDx1H
rVQskIY7lcy86U88R0WxOvU0+qmQ4QOcTWxKwdz0K25wjIaYZJQlxc59WwKBSHKD
cE1B9XaBf7Qxzrz0I9VVReOZL/5zeumsnm19O+Bep1J9dwP908zxWfxOinoBoleI
eczwZnBNSRIUbjcbgdMGZYhwA5xDIJTFcfuw760wneKueUJUSH9li7vc2dbnrUIO
QfaRk7XWVb1vuDTSwEV7UM3BvWWLPgx2kJeKmXeCaDRcXb6KiQ9AyzmNuSr0l/BT
sOiZSvmGn6v8ZdWs+fiX2rn0YUkDMLdzp4fQxwqkgC38e6ndEB8sz7b1vea8kVd+
2h8i24s5+kH8FNWgJM/xlPj/P7AgUI55uUFCv+FFuEV5YQqBnTrMczjm2vZNI040
qWZCJpXQ2iycBnES9QadnhGmgdGxf8O86DMC6QpYav7b/zBKujm6h0qHT7MStkmN
sb7fcBF+ZAzaEhk/SivBK+05QPEg4pt3zQcP846b5PGFOd0+FOSOpqU8T7L6WHev
K7UaZi5qzd6kg8GqlrJAUFn/pMaFiiP1uDPi4CCRrm+/qyuzN5a0YQlAKJqxQEoO
aS+cDFNlQ7nT4/SL9v/u5vgDXgFD020HPSoYovMnE7elIm+Hi2716uw02UHVa1xd
2DKGlS6ClqJZhEwR6M0uXFj23sBn12c+Xx54lKe73RdUblhbf2qky7zKGyjcvzlg
3xV1zBqFmubs5GgW46Cycwdon2kE6+bxdCrY72+dW6XqBG69rcD0+6gk0UdK5rWl
xFs0Ne4xv+TFrAbOCVBHvGpKCLjUneUR3C7V5cIA2lLNKUTGZ68axpOvyLmFfxGq
dCPojWx78jPYr13q8y205KiLHZWxIrctfwUywIxtkGzbO6R2etWxMICiVxnpycqE
/xcdQzjPa8xx3ykNDNjaYauchPBxNF5qVVnOx4YFmwivd/MpN+jtCt0fUdf45a/p
n2DwGUk7GEbRLg5MQ3wIddHr67k5/wt5HdQInS9eOAyG0N2KQvQLP1mnNWQzFtaE
KP7Kopvq7FJA9t46f+JO0LqgTOzuw5YEOzfnLUSpWVHRd/RWEdKQ+CpW+1IlRoED
sgQSY/NNAjF04nIZfLSgQu/8320ABkCktMceAT0jm/OBbBozII6xQS1zGVaKlC+U
7wQmpaSlCqPvfuES2oxSqB6CyXMmQfaaFiYgIkIjJrJRi9lDNwr6af0RKWND2RBN
CuM+Y+OSxyawPHbv/Y05XaR1e5i1jui24/8EqvM0sntGO0yOAfuWMiUnQ1LWu81t
ypEOr+EUWsKf32qYdKGPR1+TEsI5uX0z7jM6CDiD/QiFuLs2CAkxG73I3YThA1E1
HRYuNdmz/5bMAaZGW3ZPpQjko+DliJm/rYzQcr710UbIe3auoNgALK4qC1MQ/8VK
9XuSPedCa6cJ7aaJDV/KVCKE5J00D2fyQNXF7aNUB/MZxcYJthcU5s01VABn0+pv
Bh+F1j63tAI/VV/yCvN/MSp03Se5y7tp69kT1y30nHyYj5NHKeLuUOSYXx/wm5Ur
wTGp+gJ5smcV7rcJOVs1OsuAOU9r+XyLCLGx0WTiXhiZyPGdWOJ1g4bSdBhwAi0/
sVI016iRfcNUeiTQFtkEXclu+PN1l0YMzfvEayOKBrCUqpeLhEwAQcJacQeqleP7
eUlb5KnpLar/Caes7327Ptl9XoQPeseV9d1/SBeRDtvH5OvCEP13lNFBlfiKcEZk
gWTE6286tERSbNw/njGVi0qTSr9SPIXpa3ARgx7vwjE7Ry2UEe9V5y5wt8rI3ODh
xzb8Pl3HlilE9U303qScPosCDqhnS5nxOo68pun/dZ72Bq0gilnglgRrdylsZGXx
+lKuUZBeQmo27oKpKRzI+T/EUwAxdl2Fk608smCHoqKbtJgIVjfQ4Ame1T6QSlDs
eGW+jiPIxOJ0n3rcf1bRhXd5TZftQOsZPUYteAIftEAotDJG8hknIH8eWLaxLm+i
0u1HjOFRvWl8e6Djfwbc5kKdVU91fQXeMp+PSENZ0QTx8QmS5bT7CvTOcGOnLXJu
FbKt3DMApMMCIrf91O/cKTMqFcdywb3G/E4yZC7rnHNMdnS84bXH3KXq5JJgXo8S
ZKkNCAUvjKqxYC/WzLnVe1mSaKIoCcve7fqh9dLQagFUgSYXwrMnL62dJaaU1ubf
LdAg1J8AoAxHlfZCL43mRiE2tM4FLZmTWcI/F+jzcTuFfZVfO6rK+1s4qdphkebO
IYlO7csyViS42cJBKFSs73PoRjbrqsTG2lxgGZ6W1ct7j8H8qYjzE4OjvpHZADzG
FvIjtbKq2S7Pt8nV/fyc4QjVM6a5/vBxzagFY4IBGEBM/ADZUpxwRPcx940EIt2H
0rj3b0QyQwKvhOePp2B87LN4gFbgTXT5OqdHPTDrCTfdH1Btj2mDdJtcvbKkNNQn
wdAcP69Ju8SvVfsQAWBHxrURuRywsCvOpDCQW0MiBmLOei0+VbBQL6Jrw3oWnNwY
P6L+Xp/cN+98VnqOqcQDPjk2l9vLIsVhwT0Gk9BkQ0EYfPs21WM837cR4V6VooHl
RvLt98/agF7Q9nzGNP1opC7V4YYOOZIV2sz//t20SvlEBXAbAZVh6cXr6QXgNK6n
+QVfyVsqiOtlKCkp3WnejPJZ5CqwmWr7/lkFfrrRoVFnnf+ZshBm0hpbxYgyCpbr
Pbf5kZW3TbGLbGRqSNuB7WITjsI6yVhD/cVi/mUOhsDCngzx6zthAscPAZy3MwFu
AK48fmVfSP7z33yXajoiLMJnRqwpdyneFnP5Tc3WMByExVjxkNBg1elCqH2dHObd
ZCgNXvJR2harrGWHqMYsZxqnkfdy5z1twYRSEz32ExcNcCS0wAxCPswW601sxRxU
9QYgCesoYI1/foyXlb7MmSm9rqzXX5MMFl5mGnIbwiDrpbJZq7h3YgucBw8bei7K
Sd1/Jj5kfj6en408t/kgk9QGJS/5zNxWt0Jos+y/RUvi2f9aR8Zws+dFruNRuECo
HSafZtsd/0j5iCewvHTTM9hnz9fOGFNvWpDoBdFO3wQfTByqcCOxE3Ne0HfLON77
J/CfIQ/cAV6dSL2LI+lk0YQBnCMGeVTW5CskKzu8DW9/xzDZaDLpgziluxX9tZpP
8QG4XO/6D2s8FiCDV5dsi1BayPOTcyo8/eC4XE4Ta3cAAVRKhCMGCBgNR1sKhbWp
CA6MrMQ2DeMXxiYiW87dunMziW6IDc8BKw4jx45acnsYp3BgkFLGDEJuyS8957SO
MO7Wn0ADvUhEwCbs2LtYyu00tk99iRQkNnTnnXsRSH/cH7QuMuHCXplY2sgvlFyc
5doRmiclc1iGGEbI3uS0GqdHnvwo0TKLU6Jz9ov33Sg17DFSdCvS8psS3xG86sWs
/y5hldDrIDetpapNe3/boZUmxZyEbkeTbZcHmMIJllyf2xRlB9ZyTy1gxD1PgdNk
Efv9n6FAHEi2uwwQ7wqRYMLOq2e400iZMYQMsQrnrrLDo427yadruilpLRBlNPIf
E4zkPOH+NRzqX4+UZriTFEFFKTNMFCtNDZ7GAAuILgEB/tDVaHxWLNJ2IA94m/ne
E8whT0Ulok/aUR8VL1nuOmWkP5/jDBTiAryI5T+SidyQVPHVM7FZjZhue9LTzjnP
vaD0/c4nKl3JrE4ZiUeE2udk++qL/TUPFhZ4cDdrmMCNTGcKBgC8uD1SuU+/quMK
ztXncgo9NoWAp6xarQJh5C8ZohAFs4QOdpC2ll9kLpk6ysY2Dc9mXRWeUBLFZPzL
oU2fEtP/LFwOIWH9IRbyXV/IqafAaSJYjDGu04IaFcvlZVuqAZi2xuFi0zoXKk5h
GLbPGjE3JAu/jRwx/UQeoK5/XDzK3fsoLFRXqNox2KItjYpJucIf8TPdOKVWKvAC
5k8Ph56w3eoGWRDfezitECF0pveF9THEiaa/9b9g3mlczhCRiRQ6rNWxopUcIEAb
B1pKlol2kKPKnv1Wub7ec20KBZsaIuCUdjOFoe52/Mr48Aq+oMROYTbnJmbeDFyp
73RZnXU/txzREysb1YE87ZqIggjfXOgg9Tp8OHk0WmsGofSDuss3z/AjvANaLT/X
/nF6u2qUmaEhxDh5AJM3wc2Td2qWE/FPj9gKysK50/Qg/8b2jsEw6plt7ibkAk5P
wisB989dfepkP+F/XnjLQeLlakf/zVJUhtSz3TrxWrcm/grv2XlZsWFk0wdU9dUC
cKbKKtU2mMAcX/mn0yDvGEHdGk4+g3PILm1bY9pbBJm8iKt//6bGIBEgUk46mB9A
vyswhlmhofLsYTAKxT/TbQ9S4t9kpS3ccwIQ+T/rOVb7Tjdx5D2BcCmGlIr+dQL/
0/0uMHFmPkaE1Mryz6UlnvxcyeZxrlOrdjOocXW4zloacRWRIZrB7UDQwq2NKtG7
lDE5NYUeRbVxslCX4szbcw9bmO7+xLrWzS8WxRDB0THtkDHJbdDx479hanylqYvZ
C3wrtHv5ln9k4WL6eshUC14qoWv/P7fluX2sMVpcu/mJxBPysGrt4ZObfQ/3pvyO
9Bz+4qwRAPY/FiTB6foxA2WW7hfpn33GzqwVr7AoSC49cpeiNClCAbtR2jtt5v8/
W2ocppPpeqeaeSqfHUqBQP0y+kqHMmMq5TKCo6sNR9WsUAfcWambpE+8p/8m7SN3
7LOutzvnFqtAgj+pZRJA/7ZTgx1FVyTJKrVf9LZfGpk0GolnwYsJOhi1dgJAjoGx
zjL6WHb4li9Aas7txZpQp399VHlSy6NQlOVh7cTcP+7BRDb7rLWF3dxgTgSzeVLI
7msmmdApPljB/9oRJgB6Lyjl22la07248RElP54P1axmcvNDTjZc9psQlnxlIPZI
mn9lQfcFc7rdS7ODcPeceklDgYa6hlMKQj8T27WDNIwijxfyNaCFTj0KoQ/tttZ0
BW1CUARRlBsUvmoP6ZISKgFefCFB2UYwe34Ki3a+JZwS7wZaj7qlYmszuLMXF7Zr
fAy8h8hz8oQxbUG9xedE3g==
`protect END_PROTECTED
