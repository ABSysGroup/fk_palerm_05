`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RBlqDTKDi7gedU5n8FygR1talCmovJUDU8omZU10Kg0fHtdKDb1Inh5PjcGsPKT0
Y8Dl9Ph1ormZ2jJcdRmWJrnKuuS4+Kq2tuC2YYpBnbDeKaNpiDflRnDYXewrH214
l5xnmGsv9J/yBHTOJz34zXC5+WZ19T6MlH4nbPgI3P00+7NYEWhBQG7z2wJr2JJO
AOaHrOXwAQ+d5Db5NUBxv31LgqlLvPLCKdtUX5um23dEsycZa63P4QCtq3s2h1qL
XE3J4PpD4ygLxMP73Qrd0tfxPgRiFgvRqWhVqujC42DDVsDU8Xh/eWeEOMk+xBos
7rkCV8l64MLEEMoHssLrcijj85XOvmJAa3o/ok82a4PQBidkk7FkCegJgPsIGM5e
7Fuc09AroZ136nHyAKonA1aqw9YxYteiDbc4K380jfcBUit38ZZPOqvBKSceKQp4
GNRu4dbf3dL5bd8y8L9/dhtfaV2HyPjEoEg1a5aYR3bfiYkp7Nw+wSN2aFiX2+b8
c1fERDGweWyla6jQepzdnRhNCVwMa2wQrIQbQLRvQzkdxeJ+FnaUTSHEN/fRhzQ+
AQX9DLVyndtfvOqsk7CYf2TrDK4ZuMjxu9Hk6LdxkEs3T6E9rBOzS8lpxB9eb/1P
6QyIg7YPq5kgC/bBS8V6gJ4PDw2fNtHoGFB+apcmf/4N0Y2c2o06uF+htikHOi6p
tEPd6Wty6QNEqjkCSJ3LJi59GdeOnDfTTRRmiUFRxjDakgYzHP2YdZU0KQAK75BE
pr1NYRrMuggZMq4kZVlqwLsJpPaDzMmvKgcmIbAffvC5tl0QyqxOBKQCCtNw0TF+
7bkmNczj8S49vgQHXc2iItwm3/GglPzImXVh9VU+KIL7jFVGthCLTuLArKSkuedB
9uDexe1jBQ+xJvrXHQU0Dly4Q5L/DHhI47Ei4+45rWD0tPci185uftEoMcQ+Woe9
4Hk3bgcO7y+aoI4hmDZnRz8smXny9+1sJXHv5iEZ/G+2SePQsziILUefzREyhczH
cHs65J+RRq3dKnLQRazjYsBJnGRwEWLKrfTI+KjrE6OBORS+5rkeIDhHCJbvazYH
T1D5jkNYzSqftlXk2iil2btkU332lcKVwEpr6AQRuHvjVZaeFUEIJZApjzTX8r3p
ek8yzeG0JdKe8jCslMEov1YwQCOs9EmW0u8xAhnuLqJBbInpBgCHZ08LXbs2QZU6
AbKzOYKLvT+r68+89B/EFr1VcrYr9Vc961DtEKZPTcDct2wLOc5yigX/NWZ2RDaS
fCm9Zejbw29b+s+6JOOou0JOEGLdToZvoAb3kBxSLvJGEXem0gggX9ZT0txGwLRu
QUzec4AiL+RhRRFEy2tkUsX86dVA8xg/5Z3nvFvn6h2OhMBlYfnKX7cpEYSP/RcC
9yuUE2fciHeETTSL72KStaFGbsa81nrQNK3elteuZ4JZJGNO/tN4Lm9x4he2nKKh
F6Y++vMHSvjqUBph/c+wPoZhDFqJo/gsIToHgEVKlYNmtuZzmLHRJoqgsDf7XQTo
kiVWU9d7Iesl2Y4EOovabqFeGrg1iaG6c1xWPd4dUq8Kr9uzm6AaZtXOtDRQI3Vs
hopdQi7kD8kHheF66v3OZlqWUW9PIDbJ9SAzFRJXHwnuB3Zvb5jaamRM35+9LhiC
OgTUE2mDu5qRiV0qfY9EkTFjUp8d24bRWpiBIW6vjeu4AD2QelhbfTSGh5WSLI85
EuhcRZITyHLFLwrrhx5hFu3uSJS6JHq26Bszt16Xx5TP1zNUkjIYSWvKOw5iTSRb
Y3d62sLCXCPh0MMLFXPE0vw4mnVWWbJ1jEoBqm9L1C/FFhN3rgmASDGeYKTGsZ7B
t3q9LlzQ4EMSXJHGr8pmjpy4cHuEj5NT7AndMF6IfZztLs2RZBnWkGZPV/GLzaYp
uSmDGhpMpFANVJ8OYT3pH0OrHYs/8Aj48jEKMTUTqpoIBsQ/4MNcWOQTuHlxEZdn
6KxDfloWCkpVTYJVSCFAXOkOjIQwJ71llxOERrobWJTLdx4fkcHCi1MfUkJav0pB
gk62ceF7Lvbcmun/w/IivgDAmCD0Ogtg9jUCiMO1l0hqF1TjCC0czZiJlpYWQPVn
vyL72MQytxdetD5jpS+Tzw==
`protect END_PROTECTED
