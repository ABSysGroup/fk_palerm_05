`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7eyQIi0L7KVahtrA/3bNeCIdn1YH8d66drbNO3uEfAa8gf/taxmb0kFgum6DmJHT
RMMk4HsD7/ZOQxp5HI9iskO4KJg6ApoEskY5a+em1TyIvM8E4h2R/WM0spKx2/jp
naoGErvgC2VLaC1/TqSAcQlEjPDi7Cbk90yL8hqKPzRN7uId4Afw7m2ZA1vUrDFV
bOd3W+Gf033EZvCOGxWXX+b9WCHjXG7Y2LYG89XUhWo+rvdiZKJTDnHkjluH6jms
utBCODHTG9xRgpyuBoaYq+bOqANZ4IqdM1CrdQz322vnw4b78vpVejukNpxd4cuR
0IfBHpqR4Svu1bTRIu1/DAcighhswg3nz8mAvCG7j4vtIEXaV3r8PU3XQqoqnuLz
iZn0WWs1XPdGfvOV4K/SCL808lQUxxWwZl4QPW2yBBTSK3tD9zg8RihdQ5VYQAK8
`protect END_PROTECTED
