`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yBKpT0XDhgsgssyb3yT2sjK6cZpIc/TA0R9UgE6FExgJ0fXtqwDtoLDbaniQeQ0E
urFvzwCvbLiyM1tYa+ROfmufekNkilz7k8kw/KTsa4/ZNq03MEuuq/oN9NWIjmp3
jlFhEh6K2+WKvg3LFOM1ViYOMS7V46RfiaE1J4yEg4vO36akNlJ6rX99mdkBmTAA
DM3EVm195CgfwrGIUx7UUDzsYPjUmQjOFh3FUyHz6akKl0AOCnLxmR41zBOvNoDT
taXOfLWhLFdJVdXjJFfYcycgdb+kBg7tcNNZTa6chXesf6B945DsDhMhc71/Sa8O
kPmrTH2YUGCsnNGk9yltpxEk0OpM8Y+xGA49kXq4CODbuZJMZ/mfYdrC7EB9Zi0e
LYYzkz59FcqICLaN3leyr67+90dNbIKDwx6/T+pFWb4Et96zLm9vNqNGbyxBYJca
hOBLiT41ZEOKTU0DGj95GPov2MsOJ09gJICxLWBg+jfRPtCduh/nX5salcG/on81
F9Jx8uMwn7Nipy7/k/oY2BWNHzBgESSOo5LkNmw2VjS4KIXUyh8TfUV81YQLlzld
+nH7zD8Fd0lmLa8+ZKvumhrNp8nzdpQ0uhrXSfjrHzFR7kUcYw3jiqWRY4n9mZ9T
I6mG5P0HtIJzDzDmWtLOOM57KPXjvlQmceGCorQvCp74FQTRojv3HfBieXJiD1QE
WxobjWPECKjrCOH9jW/umT4xnlWCoIXbsfi9cS4imZnBK8j3AJTYsITFZ+ZjTjWr
LEzO3Vn76iZhW4pMRonF6g1XGlYXnJa49a/c8kiQzROEXXSMHhhQ8eL7eG794nQD
hS8ogTHel3gC3t0faPy7ixg+nC6RksbHkJxWAKEAoQpFW2zh/yUJ01caEgYJpcOW
QINGGBcLTah8kB4H2BWRYzj0kt+RRXg3bWQZItrB4WI6/BDqKA3dRUsenrh+PaXU
`protect END_PROTECTED
