`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IjQR8RwKGUwIOUzADkTMK7u04ZA6Gf30DwutRNz04lpWcVHXnEZwaK4lwagtDFGq
ElhhrCTqZSaesPoaPFZhngzkpW3rZR38DIyXhtm17DeyNnZrxVLrUA8G9DdDY6Lb
sMVZcrxCxtKzQ0N/6t9u4kS6+t28GgKXJ9Qrv1qhchxI5u8mOlDTxQcRU/sYAp1F
4wZl28q63nAd3MHv8Wpt2bxTyzKEXRkYZUo3QVYddJbG+UTlmhP9px3ywvlxv1HO
CmlLcwbrelVQ9HTrTGOJ2y5cOEl3kS0IDTfB4a0NVCkgsjoczVy8sMNzdR/r3WM+
VDT9hFaWyzlUwm6kpqJfZGVs/n+31BnrtqxeLfbCVrECzpFMm67+K1P1fHbIAzIe
TBcbdkTxq5Q2HgQfUjP9DhhbmRvwZP7OBISMWQ36sQNMx9L/EZisklzW+TnnrohQ
tjTDNwonLexFcfvqtpOJrrR3N9Z3tGFuV261L8egoHbDX2ng139bmHo1UEl8vGRz
LYWwiWMaHz52t/6PYgSqvLWi/PFLavGjQP46Wh7HjUeIGQO3X66Retunx916ZEYW
wtDU11DOpMBi+a9YCY/3PD4PPN2NnX3FifAdrcdMamtpw59LgbxbiCIPkFWmqc/V
TA6AKR0lGkvWeHT/+qoVj+IlpQegDWsNDQZxXyNWo8z9uObvs5I+Im9dvr+PaAQz
Fi4qPMwHZ9AD3doRb4p9vg==
`protect END_PROTECTED
