`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sC/8IKJxMoNz3jpEaHr5XOgjN7D1a2V5yD/+b4HetwNjr+C9MIf39K3I5y8i0eAc
2HMDeOSN7jsAORu5vHIrfp8Fqe1jL+GC8ZXWkBC44+Bu436DsU6Z6OMVPNFFP2YM
OScdjUFO5sJ1jhrbgnqQ6L7C9nPzaFsJfOxiNQ5XeBqj8ksGNihFMbXTgJhBi9Sz
YIVagUgjQzY128hgyYVOEQg7r+lV3QU4itHdt7oF3Mt84yUhKvsYdJGXVLcZK1Xp
lJiI1V2S/iMJHUpJZqOSJSCd/wBfGYE5le7LQKFkpM4V7Smz8n7pQ4SW/gl8Otfk
X86SdRZWDLJte+Ajm8u8inAXz3MG16cwj7u2cgm2HDh+pv6VIqUQLi2KwpRJo6nG
L5tRw+bSPca8fn8WNfqyhzcyOrEjwh9bdNB+GOF7SV2zCvP/dzHwd44zD8+STj0H
Os9kB7i6/xIiGCcsGYNF77HYgxfteqildbZ+HnvzycRzSlxPcpPm6OqtnJnr3qiT
Pf1t3h0f5gUu3jftg5M41EX8hDDfg6qSFp8FmIzEhRKCUd7PmMN2M4ADrKPWBE7T
rQGJ/syGqr3hrjb25Alpgtsi3sHxt4KJFlEw7dBU+y7wEccpdsAk0gh/wRiFRnaj
YY1+tYmxN6CE70j/ECM8NiffEu5FNmyAtqSzax/8TMCjwdPi60WU36bUo+64Q3wh
qDCyvtqTMgLhQln/TLCNvtebL02tkNVR2xQZZ96jDmqsa7ZZ5YNT4R9gUJFSk48l
VpkQgEjXe5r/kXZuxj332g==
`protect END_PROTECTED
