`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hteq0u6wmkXs100z+BeOa5y9NHQgVBCKX8fNZnnOAt+ilsAcz2+GdcAPMC7LuiQi
tceTnh3D1/tKVz6AJY9iL1IwdetCms9mmyLsrkabWty+TFUVNnCcz/AFtjKAyjsz
9ga0jWpfp0a6KtJFGF/7JIns6trvM9kBOT40Qcyvido215ghMiQdxPuEeSSRcLY7
NagyY7vp0lAY419JNoH4KwQm/UUsuYlo/sQGMta0NQg3hU7FHOWTNyy5L0xFkuoY
DprxbEOaplsWP73eq1UmwxGEq0FgyZfAMHMrYEHBp7Pi/THYh+Nv6mcucJ+khLFK
RVgPUBOCN0+dTmWT3LXSRx+nLlVnW+T+GsgL+MmEeLeF4SIGirUoW8Js+vRthP0Z
d9qIHO0atnfsG5SziPraNmcAL5RPbiN8CxYsgccQn3+qQXLK0BLEsBpkNLSZCmwF
7FOpxOFPS0h5eHP/IjzLKPhWIyrWoE4NP34skDiywKIi882Q+NCw5zG6+WdlRu7L
jO5rdvh0Zyx0Vz+M5RXWTNvWFRdxC9GB4qRg8mtk2N/0OdgVun9MwEtFvU4gdSET
LoRridYxZFcJ+bcg7Of61444ao0wtoQkd3m9/HQHTX7n7+6pCojPsEgIF/cNQcE0
BZI8m5Q5i1AAvGiBgqCNkZMYwWxkWOOevQ6j0fNv0OGA1SnvwrZkbGOwTaAH7LxY
a0Al+eza/OxYxrR3yX2VBVySFXJ1nRIitD4Q74l4F6oZeciCjr1HWww9QhFK4Dp5
csdBCR9KH0pjVE/fSXJtQ2pz4MNDST41IzDPvBYNQYo+WOpwj2msbMgHhxq2SdR6
WjXRhEcLku7v2ZlbaA3F1OVey8nhMAz2YWjiqIMnL45GKkUOkQsBw5/1MrNEHQDT
lh2wbllDuDIwxceAmZS2zy1qlK3mhB/ys8qcmTn1/ayc+kuoEhv4DjT2gCqxWYkE
1/ByjXohhkQiPgt5LDMBkHYW5FFRgjD+sbg51cwlhXE8OuXoyZ5kCc2zasEb3ZbV
CnyoiqPLlHotQ6m2ArQD9KioyTMIE8XS+2L8oSI05OFEztYySTb1oHb3w6/vjZiS
R4JSkemu+0LabuXlG1K8eHa4PykHzPRvRfS7cbWvSVX4ees2+kudxoXf119ZmgHs
duOwAHTxoDGOHyOulpDbpyiJa0g5ashZd9DKa0jX9y+JxQ3JOBbFV2dfZEseDuP/
HomhKeoQvme4m6ksxNnP7pmCjcxBB84svldZ4ZB1CyCPPN8YwHK9iZ29tbXg5RhW
y29VGmB4L3vU339m+ULyxES9MwnVeJx9r7tUSMWtB68Fv3r/yNIzu3aK5JqA/+W0
Rz9y92gTJ0UPcwuFZ2TPtQSz1WQPCVhGZHpyzhDs6viK4ToCsvBoz781wMcNEApL
Zd8XcT2oRNnKp182ZlOYkcB4ob3HvnkBaoUunC8kfWTyhhYj6HDdOR7L8Rj6Cqxq
p21MsRcPIN4mAd37YPlIFM6RJSG3jKGYbyxzD6RAKUSWWe9JHcXp4umD1QIOheaP
2r0WE5sKS5D/HLge1eGSsRvlBrc+vV3kAOcJAgSl7lCMbs9ECJvgiWH2EPa9i5eH
QfcB1eDLX4EuLwEgCXFOaU+AFjvBdl225tQii3l1+FI38qeeRKHF6plYj7aQ84jp
pxX5oLWdi2hFtJ18vdhwcWSpqAVfL8i9CiKUDd3v3xbEOtjFykLYrkXMjvqmBpXy
9C2yjageJ3OkE08O0NfzCXe8w3zo3d+r7KiYz6BCjWTYBxguTKl80Fs7DbLk36Kf
1aaY4YLEjf5AyhzjbooXtLYGv9WmMEyOgRXCQeUhX1VFd0RomgkS0Hz/mms9AzuM
u4KD2qppjIkCaDzQ8uI5cXBzWGGJORCuSZNbrw9YvlVStcjkoNw07qSkrFJQVX/D
ZuXsxtPAAqEFrb/Z5fFPXzz+yPe/ZoeE4WFTa3wl+HZ9lBEo9hk2VdUUEDF14hIh
pQI5w03wPxyJ3QprCXOuaRQsiEh5z7o0X7D5g0I1D1RUQn1rxBi9jrcONPU1u+Sg
0DPgnnGiA+5xtafz6WKrcBx2UV5CLnhaGKf49uMW4IeUk12pCn4UsL9tVQUZ7l0T
ZNEt2fcvWnoSzxoi0LRgaRYIf6jvT0mDd6b1wpMx0hxtMOruX0ZVjMcL62K7xFTY
RpaaWW2NX2ZKGfNMDZPMkmpYIZ0iWL4tQwQ1+n/bZLP6wysVZ6AbYwFCbIuRnolH
+MrTYroC0dBuXOED2HXUocW+y+i8LooTbGj499BGYR8i8GPMAWc2osvLEvUSK5bd
KzCrIaM9/BT7tEe8tHuZAZayWQDQjR7dphBWmcxMKfWpYGG1KxAZxjhBh5iRdQzW
HT/d8cvqFrcAAkHHGUu1t8RHEgponq0d7x+2wuioHCpTY0TTQOzt1vsjq1+wkqIw
kDT8bJqfRIxn5IjfxRq9lAqEu/Y2o/7J+OuelXeKisJanxgCflHdovB036B3z0vL
N9oDPTmmI0gsD8LX6VMw49aF6/T6pNcXSC9bEEn+rD9ZUNIF6jnn1McgTCJ7eRvn
00DB48JSiIfBJQzjYKQzKAc6zv4t8LG0h9WC6P+usbXCVOHUHWAtpjSII2p1VEFu
y4otwd27PSK0AZvsqv21ik+VI8e6l1fr0HwdJ9QqGS27L9ziEyfqZuGmPOIyg66E
j9R396pzcZvMe/Pd+URhzEiGxtl4ghbQ5a1UuIOKx2YnHTt3zC+resBYavtN1ZUF
8bD6Te4lqTGG1XKZKwMK8EPugHAfDKQK/XAd2ap08ftNzrTVJOua6445cIfeCjbo
jhvgdqm4kYlUKj0ypH7XGKNKV1hemjPG90AWQK+oGhl/QRNL85e4MQQCglf9lWmO
66yPCYJnYaXsufhtbEpwxgVNoGJYwtmtAP8O6k2EVAAj0CV3Nj//sEXfSrruUwdr
PINpa4Sb3w+npimCwn0aCOWOw8x2jr8OEX5qyrR/QQEjS70qi26nZ4SOjUJmRxV6
63H4cc5eTIUJ2yGpfeb8tSzKXSY2Aze9hG+ogIg6wY2mysbOMpJJs6SyzyG1GZi4
30Pqac5WYZiL13MxbIHZX8q5siAYcAUQOpPmvOC1UY2LneU0ADMtjeSxLokGl5Vz
GtgR/GWtRAq9my0qysnCA1QaU4hQOrh3Xm+jU2L1IzzuTDyuXuvO99lKMBEzjk+B
yZ2bz2GDsr/2jHPYF/8N8+V3dZT5YV3KN9kRULs2ojz4Y2RBr3kH6zVGqTkrFbkJ
LlMCzxwgoJ/Qt95NRnjyPsKZb+YSczACiDypifzZUaTqGL8d0QHjQ/1U8mt0Kyns
5FN2vUmsrFRy8pPQGxmlpVBjX9kpQxJAXcTMNC4NCSE1ySHqLN3ts/oMihDAZxJx
R7q+FzJn/dimjCOBIgjqQGz1kWPz1ObPd8AvlYT0UjSzF2y4XaE9+SCyExhJtZ9d
KDT3Sx6SZp9F2hmFwospBN8+tm50LnXAT52YLKsKfdBhOGtfJO7/F0aAJuJMhHdM
zVhkCluHnjbdjsFfwGedjnJEQzgRno6Pdhm6mmmNR3lz2fnxhCEhN1Ve6Msqslqx
sVB/fyK7kC4QwluTP3kn2DtR9XjFGkIaHXXxBywpMcPQGuSnkjKHA7OXXXfIZh/p
q30amA04Q/8p3IEMb0jV8iL2AgyNkrR9aQgH1sW5IrIRf3BEqJ8D4wZApWHcBBst
iqA4fOA+G2jRAxs3YbCumkjhJ3hU+mjhkSbu0ekxzsFC0kJu4Cy3dRH6QEd21wuO
fSeoCwD4tamaa9kRQzq3WQGBcvgUF/YkoCTUyDW/iMC7UNzYLMtysRn+h7ezAV8V
TtmicmoczVpkHjj20FNB0km3S68eKzZP6hnYUk/2FJb9Jemd/vyQRGVAPgBruj/t
o6NZSX6UIBm6CEKeF3o9ovv1xKIEmt7/zpeUlRU4O6ks/pNdlzTB0aoWuGDMHzmq
dJoRvAWTmq3Zg/CXacVeQfhvh10odPr1bCeQ+UL95gEb2RsNkA9KRIkz80mylrmJ
k5hWYOjf2Xj5OLJ4IkwdXdsKXvvSDrLCExwzYgaQ2BWjtrhugZx0zqehRZDV21qQ
ntZPrIGTgIQ1cRFu6pNYrwXtFK2XUxx45EjyHlLsXB5hrOEFQgNq78l6mKxfyq/6
FP64X4jvkLoJwHb+eSp7sC39KU3I0SklNzjf2pRBE+Upq3wRhMtG0mXhuYyhDN+V
JVIN6g5VG7CXluroOmA15z1Z0oa59TKFwbzqKgKOkIUPVVoP9klBTowTcxfKhqWR
oQ5awzDY0Nxnc1ZiqiE+fld1ATnMJ7rhyrQsqpwqyxbShu6l3Ya7SUAXs+naUJRz
PiGCziwURjXbbeh1pmnWl3/5Cn6LkLiPCfnIxYsw+MBz6yMu23EGCSsWRDs24JLA
vKLa3AKnqH+oJBZNBXEi0ZfksQUYpUm4Njw7dA5PNBs71lfj4ZB1mNdiTz5yuWKX
zwwDNh9+cq8ZysHFRtgFZ14q3+UWS3eP5cP29T8idYpVoqrkeTHGKp13lkG3TPI4
mGfPF0aaEWnrp3JnefVQ9zBDhSB4gYw/4quzCiMqvJBrwku64mn5lywB5ujT424j
1VFzqZhNz6fTobv90ekbhTkfP+rIpEtkFMmWdtlLw7666L/d/v3RaHlFPFzPAWIk
YB3DSiI5kze7cIf/geuyevS7fg9ffH93EcpMsj94MSN6sXJa6gZmPJJeVwwleZp6
lzTsadOcR99VWB1InaAURj4Tmx1/T3uc3EsMDDcIeftM6655CRMM9y/yUz3tip5M
GdcAypmYz8f/aefzjsJukVzvnJ+FlWWhCn2cIV/Ykuh8n5oY4jgABxOlRKC3pPNU
3mMGDK5a/e34XK05bMzxqndl0JyYDrpAJL2QmdwnCcwE2BEEwqo1BL8gsscYs1B4
VnCCSVT0thr5iWEtIZ/Y25ITEixJSM/eDvovC6fRWZbS8yU9rVz+Za2PifxghR01
2fRiMbvl8cUIgpJFAUVhOLEDJQCJBEKZxmAfg/+E+pvtVkk1riJBs1kRrS4Wv6Ev
oBQqPj35iQbIgevPxc9YlB6mJU42w+4cs2JBOoQcsrLrK0rOnjbjTSX3snUoTBls
rYDiT8RsEQU44XYmY89jJ6H5XF9GHCXFoR3TzzvdXM5JOhhgfzF2eZ4ja9Ti+w4j
UnUYlDn3cc9nnTmWtO9fzuLpIrK9NDV6DLWGlHIcUDI59CXuoMX3tLzns3ByOSaH
TtP8nGnMOsu63FGR3hCY1UWipIQEHwTktdS/CZKCyZfT+y1sY/i33puyBNYPCnzc
kGSk/LhxOVN1t9kxLfqetZ/cgNd81ZKnj3beb7vuq7mkTqfGXOXsS6M62RxVpcSQ
Ho+O2Y76xXfh13Zn40BG1aULmgBD2wag5kA2UiAjHVWMWXbR8FB48Mj8OIObdf7E
5XSj4eHgNr0xIyeJbm7S1qIwpJrFxzhZTf0edgqd/iWTLZnmmAeKEDS4ZEWIwrFO
pltL8QqwzEgoJoBf+m8FMESlRrVFefevVVEqSdbVmo9inwTEch4VELmr9dnDEFuN
ih+5j3ywHVutGDxO8UQhQlJAJf6oaHiYomHLHbhgAby56F45TidgyelmgpfU0obn
W06G5+w470hDr7yOAi7Lu41p+jj/Blz/osow5DPyW4Pae9Tj7VQJ9NjVhn3lDsIs
lW2II6OVNpwpKaW1buivOgsxjgw+NdcriXegpndJKbSU6fBlUv4JV87A5d7QlhnB
TlG6VwEnbtUzOE6QZVHPVJimuiVBQS2IrdTIP1nQnc6jsnd6X+jIaSWD2YgMwFq/
ebq+edofEXMkfwmgZGQNLjx0WfT6XxEMYdaxk45yhC1RFa03YzZ0B24rKSwAALBF
Ctue0fsfC9Xh+/miFv868f75Ms3iJWxsYkMWa6eUqeH5RXu3QpBAfbCzVVS8tK6+
6eNQ9UjtavErGWTwvssJvZ4htAs8mbbr4Wfe7DRgb5r7SIvIs7UoL0O0yDazEjOL
LKpXSvDIjtX76WsoY1a5WDuVcA3UoLfh2EG1GwPfwjfNQhk1TPvhN/5glnA2eRNv
lyfxJB/6yIA0Tf0r2UtVI6+42Ky32VTEaCm7gexUGweuPunmn+1iw7B8cpd8MUme
TeT6raIZs//EVaZxEnSYCxT0Rpdjh26KoSUQ4HMeEtyLRlsTt3yTqrGBd527MQ7z
SZMInILtAn7HlJ0ZAdBmjwgtahA70iLOFsChGpZRK9GdxZjaISMgOV5F/ygaf7k2
sbbqIxAAHhtfqmvmJ+7PEvzYJrp3703bJEhN/zUnp4dSYEm/KFB6DY1L4ei1dApD
1adf0oDVgwoqci9UMPvwIv9gNMumgKst5aslfCS5XeCvI7F1ko57sr3Wtn9sWmEC
bn+KPrkGeWEQobxZN43zbl00WblsZ4+BHuRhcuUBsZHrspPb3M6GGY+2EUGskmpr
gQKITlbT3GQG8P4NyMuCbks9E71hCUeamURH4bqCCF4/OgJ06L7MHZgJc1td94U8
b19bK3Qke8djXJmub8dCyXlbnN36+Ab5KVS968IAjS6OCWNyMeXIWa+J0uLf2Sum
Zy93w4WqiNLVKweyp0I6USVg3/pU5D7kEJkwmrmWBjjRF9uerbNOf2HxwdJk7CVV
BcSyKbJO0rWWeYCeiRNy656w+9BU7yngO/dh3f5vSjpuEifcKTbAUevZlXLLV/JS
5F3etpuwqEiAxbDWu+ZURnj7/WDS7AJxGZ7ZOQuW4ZeAq0OMvnn0w0KPnx6Z00MM
wyB2eTwwC4v7j8wXFRYBF1I4EF294iAIZe7SH1B4xFFm2H1kcbMRTQjHNdY/1RNJ
l72i6tQem7AAA/B2H6P6dVPH/iyy0reOfn/7X8K29w2NMDFSv3uCY0cJFnvWhEO1
2nkMAZDvBuZXESSMgbeSl4pNaoHwOUk1fj/gXQ8yh+qsJr06W51IAaz1ZqM7bifG
HGGnlr6GD0VlaL7z3UisPNkYsUKBHtbn3dqDUX/B0+fomGxgMxAdandDHaZ/m6hq
j/jaQ6u8Q9y9Ckdka7Ks/J42d9fTyGeZXgVgkpqV8mOXwCP2Qkbr2YHksPl1NeAT
MNIR6ti6yVQvW7V2QieNx5z+ZpResyBOBhVS0ZLLYb9GAVuVNYb5QKQ9lSiTc0OD
SRgCxqZhFRmOqG5nqWFdFWxaRNfj596js0m9UXT7KnNP8PP5A51AClg48AQdcJcU
g7CnnwkEMAExqWMqXgqmkKRum5hbZPTUxVfgc9G5+2Mk6jQzkvuVkdzQVj6K7Q6l
XRaigV6DwnDF/YihNbEFrJUm0qMKynX8j/eO+CrNcbA+RTas4YxF0e88AbO0LLUN
krg0hA9+/Qljkq4PYjmgps7POGHH0nw8RoqTeeejBsz/aTnmio1SYL8pODXqDdwt
oWwtT2vKRuM3Njnr9o+2ltwTRIgGoUkf8E+hns3DGhrd/rHrftH4aPFiAhvcJ2Qb
vCJt3IYFXzsOVeKP09AqdpoSZ0P9I2cHGP2a4UQuGZ+uws+fUd22kQn4m3bYrnZ1
ulih4RESHfmV6GdXdyB+mFgsG1WR8qIBpcqmDwjgr3MU2I4AoavLxDZUURSb6Af4
YcJnZVqGB7e8tuKSzlgQbgPz8g+FbwqvaVxDjD1CBP+w2FHlf+1HrCo3fdnhePKP
6ERaLusNpbK0B16F1pixnSWR6Qt5fvA3qcBYgYhfNaoCoDnDeRwxcLUUCSmvPk/m
0o0d7k0AsR12m8l80sYC9tAEMhfDmx2f0pyZwK1NOxpAPiWjTUkpBsAoevg2sJ25
9eGWEK2rZ+6869k/+y/AzxDni2bWi7MxSiH2kEdExBkInFUR1mwFrubKQI5obk4w
eBsjVO9iv8szh8/HjwuNWQtj4liwNcSarV4EAZaiw/unkI9FC/k3+FPuDWe/377J
krthkAnU0sPQ3k4oKi1VCB5u6Ix5YzQj72PGAU1SVfwT8yfHaaM9VZ60UqRdLuS1
9VCVxqTiIM4Jw5WyJ5vHzc6AY5KCUnc7YMI0br0N1IC8jprWc5/1GsJT1WE0NXrV
2yR6cDQyNpaG8uHenygcHZ7vcDQOTfZhDS1l57sDZsojJgSkeFvefXI4M0py5n7A
+NUvzfgdeTLIr52pzmtoavPs68S00Uotf6pMUyzW8SEcVbB0etrXVEkfzDikDmbo
TT/Uq0r/5Xkt7E3c8U6nZiNSyJ9s8TnBgZa3tmSpcWSPJ3uIiF5onHXfbU33DEAc
kV2ogONbhPwQfZQ2DpunJ27A33Md4XI7LXB6FJkRQdXo3NCEO+gEUgBxYutyjggC
MTRJN/eftA/MpNMI0QmW05bne78j0MMPUMlA5G2B98xpn3UWo+QP0Im0tf7jL4l6
Prfh6adJ1DQ4eK07ahofpSKFG+x7pv7NslwsfXDeTRfgDPTF+0/lSXwCZXgQhAB9
Yv+SU9RROh6P42fNBKobJlZbkd9U2d4/1Ih8/lVyh6UHPCFPX51cPPWjZJ526VZG
9Zfm0u6zRqmpV6qQgM3qOq0lvYCJRZE5BoVWv460HpioP2ohO8AvanK0WUZUj/Kv
1t8LdTjNSiQlIqo04GVa+m8vGdhDKPN9+TRHYi4X7r6bYtpeDFJjomYL1T3kdNiP
XHxs/hzm4S+fSVxbK5tGZhfVXtx/QIxVwDgv2sFmNLklTeB4HSatilwAPqLT/9b4
MTeCLhcodDO/OsUKR96e4ZCEkANcvDaDNATQ0o9MRc103M1oguwSAopQM5EA1Ao0
jLy2P7j9gXmBUuXnOnR2PK03M1KivRqeE1yLQwX3Ly+KilbvwXhQMk2ytisUE85j
wzwhXtlYnq+mCU0U0UlSmuw8OqvK0Of0xG1LMoc37HcNfGsUObiRrJpOP71mGIW4
S8WMmmAmo9cHoK3FcIzVlCPM0qVCFErsW+e++aUNAEO67R3p0HJuZoPo8mDgSWdz
EG+hADKnF45HeoCgF75HVMcihCQyfHL14+OZMB8bLmGuloOG2cnypcB0hsSW0VH0
loNQnsNPEZ145hJf37SJd43gdRzX4Ys6/Fbx0vgOFuYapzOuUqXbiV+5mcbXIhaI
f2KshzKMeVZhIJyjlOdgAjJYUcguPGwN0VXnohPOWXyhf6Wrol747000zLtbbknR
+FMveY/qKlIo8LULdpWEEr18pqjfZv/G63XI/CM+12rm2h481x9HFt1xRarXdqzW
ssyMvUAUucxGDw3xxbJAk6PLMYxE/8zfyOCRiXvrHczK5jE3V//7ql6StmUOeAzy
saevvZbGTTYeYGpqOV4L/UK2h/cJOciWSKtFJAKKwk1HUc0gZkGgsObFUDvlzp2X
R5VAsOp31KcRLml3xuL9Z2JCsaeHUrZ9Dpyeenq66XzhZRa2zztRGQo1dY1E1Vuc
LMBoE1Jz3ExKSrZK0LuK49gmtwMkxBOlgpVDO8idUH/H+sfMPF1qwUby04fG1KrZ
1I/8DCk1jIJ3U4b/+zFCrK2dHqUKWlmD1P7apn22PP41vjzVd9Q7aDln8iV2COXn
j0PcgR+2cNlEAlpaUhd7Akd69rkQt+BgdBO6AHIhsj82mjIWvL9uYfCxADOWyxFb
C73lD6A+2hIx+MGA5S7s2h8yDx3bVqenOeqsM/hDwyWupmdc3RawqZpC6brT4RS8
7KME9GgBdXFm2jRkq8WaHlxlQaUUxNYj1PsKk9Ml4UzIipnbhf1RSlqKhUfoTRuI
GSFZNOlLi+41j5adSuoYxLqGrFzUqEY1TFnxp0mYZu+JUPH2Bkc7F2sIjEjYIyEJ
E39cxtRqEhuKyQW794Mpf4jHsOhFV1fEmjToKeUlPkPiOZ16ZG6IaZaEEZ06IVRE
9Gr2Kqd+g+7I9l0cCARmHtDu88WAuwJ1FruFeE+Pw4yVqZ7Fsl8Ops2o5Ep5a5p/
WawFI4igZr0qA1YXgBnrN16Jq+iICZ5uNh99nJ27mMPG3plio13TPlJYXS6AlsU2
eveeXUUH0Sl9P63mUIjbUPESceUE+JbuSPGtaewvqZxPEmYhj0WS8x9YerEZDs58
7cT0L+59igvJBAD/Q5dyN0ocH4ENxFf4RY5Ly0ufd+PTTYopXFe13D7oH3dRVaY3
vT/dQNo/BG/d51UhaXLUGm8WT55EjZMpzXtodSgAfimD1u6TRWlntEXa40OgEajs
qWYt3R8bC3rJRwd3fJbRvFLMwjNriDBV6t5YYr/X5XStRvjN+JxocLzTqEND/D76
p9xTAaQxnWNX6UstTb+eUeMRYVhGHgFtr20Jk/puWV9tXMA/ZNo9OnBzQgryO4j9
NOkAzdazDXmMMLrT8EYd8kQTOaC/SFMhy4AMiaSEZL3CrHtXNdb+xr7cFyqnuGBQ
xCnOrZJ/aoe67Nkfsv0esTdD0C5tAskMMIQ80DN1bh3VLQz9V4qT2SIzTSW+vqzL
Ej9zUMTp1ulJZp1SKdnaQcLxNNlOweFyKnOJ/Ql7UAHBAplOO1H5CvLYgxDqKraP
P0plU6q8QxDjzX+WnIURrUWAEUtZmyuRJu4sQoNMoOuNK948Vb7GaMzyK/exASDH
9y6Zb+u6y0nR6YnCQwWFQVPJDvOk7x1IilE5jvRrYIZH1OA3dbZOlzFykcF63cIa
pxC4/7AQnLwvlYnXosOFrXB+8AZSmiX1NAIEVulinMW1vmNXNBeVuJHpUzn4XzVN
+NjzBqaxJ09D3xebSW7DfIws8owYJdjMSymY5RuMmaGIMKg/tNnYyuEZX0SgYEcM
dDC5JxT7GEHNbb+wob9bTjFeG/s3HGOFooRGfHpA7LY+JmbkzOzTL0p8raeLVg4G
0HW0I8JkPE1qbjGaYNSO7KR4txeEiTbXur585mNaDVQE0OwhK4BobL77yN+BvAht
/wey0bj8/rbTk4TJO8b3aS/0fi3L8ZAQdkayRCo6DQSIDeSuSnWzQIdhQZQybJwz
3Bz/M1c/RYiaZ918QI9f/FaUSRKDdmpFFeX18HLswDLvhywH5mVTDAlzFbpfC49C
nFrxMm5Iqd4RH4ciWupFUMIjqpIsqLF61jVHKtj0I2XwgN3sycyeIDBmc6Fmn/e3
qF2PtZ7cGp+9CA4nBB4zv0yeycylAaMDsVThJQK0hy2KqQHbm/W3nm6MmA2JPKG5
eBMohoY0lEaL0prR1+aV/WqGi/rbjLHCab8mmeoEf0lcHDduJBAjX0Nge8uqsY6C
B8ifVq+Vktz4Ci4ZAVo15Uu/hN1FNjYlGOEWn2nVcO9X1/ivQFW/vKuhd2yqH+tG
bSuLFTqTD+oRBmwJBE7hlej7L0thNOYP8Nq9qbQFGKLFUpb91igbq0eHahtqh8lN
WkB2MSzQsUySOykpejiIyUroUbMBz6DdzBc+/gRs9xDhnPhVRBGLVRgjUd/uNou+
G1q4AWqT47CpxCxM2xHKvMKEHSvoZbs50VWSaQ9RcG7X5TbRnMf3pR6gazOreVLa
xYLt21oo+t+tu80zjooyO49Fk4392NNd8ZeGW0mqIJgiA9CYHsJKpxhJg2siZzEm
fJmVCjL02MObTJh1Pt7fU6kxLxXzcBsySAYXAYs4xX0ISH/KvqHIe/kk3bXSsEtu
hlbOGLtut3b2zLMe3uN6pOeo+v7u21xHzk9WOZTUwCb1NIy9jgt5DbjS7LrRhoNc
oqxx+vgdO1vsT1ld/BIdDtetqOZsStLzSMaRbW5JjZN9aGWJK1pwEumBoVrNJXK7
kOFTUaATvwbdpQh8uTavz46w8X2hrz5k92oIL2deaNbJeAmPb9LCPI01MN0JPXO3
uNArH2ZC9/XQVEVjdYW30Dqa3iFvjSM+/ctKPYIzdefuNp7m014On09h77XPahDP
9tNoW2r+cxOURYD02OaYvZcKh5wVK0WXn/a1idlVpu3/vfrg5Fqd2vmX55e3OfSz
BxwmIA/C9qHOzGvYKxHNhp6AlXhGFBn+aAbyRiVGZLb/Pv6DC2Vjh+HbCGmTojOh
N3I2ZjFrBEADkmzEYe3QPgNSMyqgUJ0VwiK81yJQHf3OO9QVZeDiu+uLBovdb5Dx
PCi5nAXeWFmzCIFHAsQnGtOKxDwphmF1G7sUq7jx9RXtEYFaOqlpssMs5ofhGtTw
rvqA8VG5X3/AxtSiGpZBQ73l9o2PlvRTvwNxF6Xs228hFPaL6NS3HOkaomSJ1Ics
I+PJUZMasTj+fbq4k1OmFjTzisZl83bnuPqMJM9B8p10zKVDNWNJe7iW+jhFEDhf
txH8goWY7PWoCEoFEesV+onfQA4MkUTvri24zDkZAHjznHGf/ms/sOUujnTiOdTX
E4jgLAStayUnp0oJC7w66fNN8SBlSbZl8Gmub5vbkDQeIFozK5anxsU6ZqWFCdQh
JIGY1y9ecgsYBPhrYtMwiXG1yDVnsCxqXRX7TF+JfW0SKpztDTkn6DvzS3pAqDmJ
GiV/ZB0Wh7LFcXYv6YOZzDFEzelikKFUmneY8YzihMGVg7XczamOmXShOQGZkf5H
axAfA2jSNghInjj4oplhZUuZnptcfxxucMLPCNGmGYAjIo5GVVlWonR4E6coaT74
SRWUhS2Kgzn21koMcscKlF1nq11FC1GHFEN/R9h/5wrI0EVFQWC5v5Lqjmga64wl
wVS17aQ9oZs8dHGu6IiGl1I4o4Ar4BlxhUd9wcw5yLJGnGaqptPtScRJi5hU11mW
JkvxWgKzwO5jSiiX+J91EqncVvZ6TJmYmcmU9vMU+yDhDgd3NoEO5owKImJshJqd
cJeIqU68jXg0F+Ata2QSDDb4LwAJN10A3S25qf+X1gky3nm0lQAglPzgOgaGUCl0
BpB1lfYZaGaOq4i6I3zseqZkiEQbRfpky0EYqAKDa1QOKK4aNINq096nmfgB9PI5
yR0EnIAMxVn6KJM7Srtz6yxdlmpzx85JHqd0V22mVYp/7bwEFw0Bq0vQ5OjlnXTq
8b4s6wx3xJIIWgpA7dmZ8YR1S6cscEavrvNJM/cmkZg4tP3eyjZcqgiC0AaP+J+q
rGl/zjv75Y3DLkODeRUv+XmMsiSEhp5T6uH74xOfBX7NP7fkE+monT4PHTSwObK/
laqPzuL6Ly2UIWJ2hZwAhyh7JsLhYi4HVUJNE7MEmfCF/bFTxYJAfzJh51wUComd
W2B5dxI234bqmPiR7Pv4lWvfULxHjGA8nuqXCYnhovjrgP3sUwOjqd0LjrRzQr4s
VBiD6dOmBNiBLxYb/y3AbsTUbYRXg5kUUPmdp2l2K0Q2wJhnYkhsoMjSdthZTboA
HeIOYPlQfOECUeKsKxEtVOi/orvEoQlflunY8cuEpRh88rAIrvbDAuwi8bHJGL2q
6dwJdGj1wRirGav0OdPgPM5BSeoxLh7lYAJ9gJiveX+SerBsaeaN6U0e7QnxpjEb
tatxf3gxxudVCBktIPdicw0hgG6qOtCYB7D0UPRj6oYfwVjBsrm+obi3pa3HCRiF
22E0QyHHFDjHky2ztVnzf9SDfVw1yzoiwSXwnyv2VPPDhJRtlemIvX9EMeQR96WU
DzVCBcPPEWBuGFnRRZJJGIRNUmcXONNM+E/uJdhQFHmPV0Z09794X2w5gAJJPXMc
CATdoa1nDi10V/E2NNnydEH/dfeM7GOeZR9lW3E6Gc5z1RObYS3mEfRNNxXu6tKT
vbpU/6LDLsf40zYvpeb0lt3XZSsoV6zjxEajFCXStWXQvIhUHNX/NxFjSL9SDmOc
8bkmJ7cMVANzfbwY8WLIyC/boP79MyQ+FDPktpI2E9RumRTvk1t7NuRh6FUh5veV
rSNKZQxMRCZpXhs2LnjoELMSm05ILTRnGDQYkcp7lSa17rN7j6zrms5Al09TowF0
nfcacL7kua7IoSg6cEieaMqi8DJ0J8tyIn2+SwZcMukLd4hrJerbhL1MJxmB/PfY
vwqI+MeOS7lc31NBa8LUh0UYPnNvZXKMfNKCGETfxo45uzun25VdUDXBcmUXWo5O
tgWeXkeuIm1730UKhvHVAI1+IweagrVlTaiTN3QCIpmZv9C1Co2390ymNr/hENs5
3LwvmuBBhhqMBin+IWF1P+ySunLQL/lvcpQCt16p4BTvhpZt6q+n9Eg9H9RsAnpn
lETkdG31nhjNHo+13ybErMUEnNQA9rLajDQaPJzgo5Gr09rtMTbAlyVchbRxJ1Lu
ajK4K5EWfUChCb8CO8dpXg+44bSaA9w6RSWWzoixPaQLNk3UGsE5QKFH6NF6lHqj
3xqa3I1Wjnn7lLzpQHfruh1hHKK+S9sYe+wsKUg0nx8JUYXaN4Av2FrlBSDOJTG4
hn6xQN+Rl4IGWkQP/KO76tqhlans/PJznMbxSN8GD5lK24OyT1gtpI0kVEukjzPL
FWN0JU+KBkHMG1Fd/sOfyqjmEZx0aGmTv8C/Sgyvva3uZwvrtaFqDm2fDbRPbq1F
iQYTqAIk+5frdimj1T+2g/dddwUPJQUzxBU4jnzmZ45wrgIph4axqULhgoKQhkWk
nr8yKNCHII29mcoh3TBcyhxNOIvJNK8+9uu9VP/wThzBTStZXD3PkEbeHfe01dIW
djFGyYKQxXrGNU9cuAxur1DmdJXEpRR8PmKSqdlV9LhB49latURXIkoCS+L45Q8U
XUQqzZqFCvoWaK6iKmFjoHxDHtHf0i49scUmcY/9yoHdq8Q4rYN+CCKCoDOB6lca
8TAQSHVHBX6WBJMHZy9Or+/Rwi3s5Dgniwj5/3ZNAUBHcx7pZDeLGQehkGXbHfmN
GvgT1P2J8pOhgxddRkZ0Tz4W+ggPv2ivUWfuBYy0yrCsbm+rTjV1eLTrbiZHS5N4
EcohFmW7T/qy7DYnAP01MokyeZbcUB29Dc5kTYjvMSlqpQQtQ20yawW6teZNIVIV
9/TITJxGuKJHusI02V9LoxbLq5YW7BZZJFRLiyCF+wiZEI0LLu0B63ems84yViYy
3/F0RRQM7VSveIECvumepzhlYk9+5UT44Gtrp3w2g3tFTgTp3d975nDZHWQhyeBk
bkbJCBZ7l8MEajM5pEhJqMZwwH5u7tIzZLHHzsLzVwoRRPwWLodWbRB9HyRE9ceW
jnz+H29zuGuVAncFq/+yviUBY0NJhG+EufFxa05UdQWlhFXS523PxeunARtF+ZGQ
XCFkOvKg7k/rQotJkMQffogC3nGKa7dGNXSnlaI3A5uzPraTCXIldS2bXOeDSGpL
obEzKiZbNeMK8Rab2apBMi0i8iOFZPDNbEAofkec/FUzuWz3wM9rCECqEwY9OOWf
rdVCj6AzvK4CAlUyUSAg9glp44Fe55/cMJC9tV7bDXmk0ltV6QUmT9AOm3hDjUuT
5kZvkn6HH1nRhxSseM04/fAPPY+GFUZar7xknqxIw7nDUuE5b5KVGjq4KQrMVCEr
vBbwNbCC4rR2WQFaY7PqfO411IUzqDtN4RslvM17BRdcE/2RjH+DVA5OK1h9DXav
ERt8Qt2jI0IoAQjF2EkmmIHVbfPjBQ6v8Fvc1ClWiNDgc2dkhBsfIjx7gV8AVLq3
6ET1PO4XguedH2qVn7xQ2Ty4A7EU/HsNMIvUmxjlM6ZyS8H+JkZQfjlIusK+Twci
GW2nBDzqhcgpkUK9mK7Ynkg9XCnFPRsp4R6fDMuYuPuosxgfzYDwu5tU1/WHgn8U
KMJzdyrukOTiTzscvIITL1jsL2bSICDioS157PnTXV9vpmlM308w6v0cgoX7B0l9
N9J3czQhYJwx70Ky7SOBhzcHx3/t+AdvM582vnMTIml/NZmeRPUkrPIS2Lu74zga
xPiMi4I9KQl5w2Zb7C6PvcZkCi9QOovEar+G9sj2fIwYyj/QIgCUK5x7KXMl7ZlZ
JC3wDkqV/BuOlSc31BTqGifqpY4cxC/5z6Edczgk4wOGU4boocEiXe8pZvbV9trH
SaJU+UfqCpJnEx6jPOBDdLY09NEqQPiBzq1z3pMCjdp4njMUAgxNqM6Wcc7hGByv
qdU4U6RHjl8d4dMSP8RIypO4z+1ANATqtEAfOIwyQSGJ+hGm20W5f7krGurTDcVX
SNZRm2pUSIL2drGlNhWgau1qdKUQF7gjel7iu1UGZXC2pbqmaEx6WGBG+qeCs0oV
9C/sEDBxPjPLqrMZ21YzlwCk23M4wl505CLfpTrg1LyNYaZARw9jQadAl777A44Q
qcOrMKCgoRv2dtNLpogmuCvmFPIGq7BZ8A0nfBOed6hMUq9IAFlIwCO+eE9UXqOS
R81RaXJkLPyD6rACdMIAIFIxFZJBRggDx3BTi25F90bkeHyWmtWST8NZJhjJWbYl
7fpNFHzlteOHhCwOZFvOmH2p5QUWM9380NuxeUASEoPGLxbtfRIyQew42+ncOT+Y
qx4lJ8V5486vq9CQf2el47SZLM8sl3qBoSztPmE6asuopWYyrm/Qzs6ToJiURadD
iTJB+h4y+IbMOtWA3G9pR63T1q/Gsz24udsvZ1EC1Fv9mon6mEv34A+DAyQQz6/T
5RCP5I7c1UeBU0VFJ3QzcXnnokm32rSHEZnGic3G7qQtIK38gdldYBPEZaiOlkHy
JSZRsB4v6UKDHht6syjaMYXGvZqZfNb3xYxI5no6TbQEaltdhmF6QKCwqUuFjLzk
8KFQDBoADqWqZhQDBiWUnZqvGhDUfvSFWeS37lNqUXCYJB68SwNL50a84pzw9vJK
SbDz8OCUp9YlizQx5t4zoYQTl6dEtQkT6K2yHUMCgfShiUH6NkwWDqH4MTc8gsOa
HyoZOFPH8uMuRtz0L33kG/og8pf8wb2KR0H/L/RxbD9Z7w9d8XTOKltA9Tb6vH2J
UQGmAMxjPtZvl/qvp8RaE9XNZRy0/YYuf0UXn/Dz8hIlvrzXasd8kY1OcuHYvFG1
hlA9J1AQ3dlSsOqf8xAQGUHscXLazPf+OVCozoO1E49m8x7i/ZaB193X8xtyHBRR
xe0yeTcKyWufBRx1BqdAmaqYTVzbm7Hb6FoNIKzYZUJTs6oM+dI6p9b+U9KDb4/T
5pWDBYiKYHIPrzlgnvzG9YV1ZgdiCt2jz8R+yDju0tpPCvgM8W4V6rOrgXLqol+s
a3FVf+3pnB2wMp1cZvs5/DLRTmN+Akdb8ExjWbV90FgHjpkr32GPFL1IbfdTmcGS
dVvbr5h/T4J2+tZ4s0t0CgXjzuFjb3cheZdEmajBYmLEjOB1dB/c67ujbNoj1E2m
QVyVoq2HXTG8KYFbVEzIpX7qaq3+W+eEYxJpIkOMVoIcrzO4JkhKLrmW2mMAM14s
55YdIRodYHKgDBKt6JW1Y4IS++ayDlVKX11DvPJV4fEl1IeUJlwtFF0+fHN9dirU
12ByY2Xn2yHff7OtNpE8+mQz52+DajoqIphVQ26dhHrStacSQvgkaLKTgETDbKrI
zFh2CaykJkfCQ1byr/CDNyowTnUUoVFFLbUPURE/bXQ=
`protect END_PROTECTED
