`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u8VnbSgBmesUbHBAYLYHYfu9gjzXDhEN2V9FB9oq11T/+z9laEraZ0TCwk76iF06
C/AXCY8CjBkV32Wf4w0gkKCx6BSwS7+NhasSl28V4vKTNy+4/dsqUe0wNW6347Cy
wyIkBq2JkMyiK8yt2lhuTX4lbDzZEr9v7vVpCPwMu+Q7jyQTbiofERzvoXAQSHTC
Rb4Pv6OgcQBfWgLTxE7IIMv9XG801AGjZvOeEDl8uZ/p+DSF1WY3ivXejbkPtxuE
SMyoum5YfnV0iAFxAS15wJ+JNatG2aD7lC4MVpIOr12UdRLaz2rqYocsOk11qH+S
n0jS5zirc71SmiO8d4OWF06Br2WPEZZa27E/wKpmcl/xIiou05KnW3Qb7PRV/bhS
DlWmzHbyx1CT3U3F1OV9pxM/qpd1fOwpcKUZsAF0U8z55z/0oWcuyHhpDCECfbrp
OnKxSHAdU6sWgRV+Sx1pxmbJmZphnZzDXZ7jDmuRuOImFmWOVhLx2ygwnGIZf7DN
ChhD/IucR7+q2U0A18otOdoVbIeDV4Ntz01G70QEKZ+ICDeLojfNOu0nGoYoJZXZ
QwyawLVMISdRphNCrfBScv8qCL0x3T90YF1MZ2Yti585B/lsTSfaf533rAs6bOm6
nq8md8cMp//pfiR8M4aDTMrmylnvqVHFIVp4u1H3qD4pRdWpf3eoeTm7vemN+/2P
nTHFg0BNryGQ1bAv1/hbt/V4Hyo7aUlmwVYdvzqbBJCS6rL0U9qdAHhRywuD54Hk
xdQ8WWvajfVxUkSrVHilSjD4S5JFjpjA96FVi+pFkk7YV/fMsr2xrtw3+97DaPxL
JAavcbyguc5tqxc4kHjAgytavJfykZH0KAm1OF6Nx9ckjRk/XlSL0dGYTeMGc5f+
jpCA2iL+hIqsFQ8mhOIXfFe9fEZE3lOj/wHcHfjymDM=
`protect END_PROTECTED
