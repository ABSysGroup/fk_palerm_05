`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rw3TGQ1aFQOKYdeaSrRLwhgWT7b4vUzZs3HaZxELOPkrG+wgzQ7R+uKPlNEOyCCk
w1oa7MzjceKh8+584JmedpSz012CKfQejrsm4+DY0Qeb9srWal/9Ze4H8Fwqj64R
4XeVfaZW4fbeH497Dp7K5wn/b/d32oFaPuOBpyDYxFBgM4Zzp0lTCbue9uFe7bxW
JJGHzieFyuPm3ewIUop5GuwaGR/E+LIVytqYsJ6Rv+8l3VYNscoMK/hygqjYDk4Z
Cyz65FuVAinqu5ihpQmuCW1QcIkTjU9GLaKBitHpTiFNLqINjFKCzMHKksurFR6T
VzLgJrub+BND8eTuIskV9EK6chvmXR2GjagsCp5uUPtrLyuMNJGT4MwMUIn7yH0j
T4aaCgWCtgGRNgbWx4L2LAaQ3BsU61ZaI7sOFGuTnH94jr3qB6bs+hQJzv61fEcV
jyxZST+4JhPtGrCeU3g6BekZKavdUEuZI1sbOvHde6SAQdtyZI4B9BWUiWXwe/S3
pSIb6wp1GGp5yrrgVDQIPera2eUjPJRsPxu6+wlQu4KQjhkn6zdFJkO+K9o7xBk4
phbN0+G+G8n+jS4G/lvngHQ2UEEgul6fFrUF7PBrWrN4My6VqyWrFu1iUYUkMS6O
3ZyTpgL1DFvnNDYEPXwoMyRi+sd/KzFO6XsfQ5C4+hZQgRagPzAaPPMWlWYmDjIY
dIpLY6AJ/b0hqbJ5mimsivLYgg9Fp3yRIko/RPinUdxgnffXKgZwnXY+qQmaBjWw
/4SMSKkaK/9tEAJYth/o5gzaHNCoj5udjqO1IEsFXODvkzn18DRoiN6juXn23Des
WykVpgX2rzIwpfr1aUQ6s49fSkjMRsiSdyWOyOU+MiS4+0BM7CIUmUPIgd3uoV3k
O4xVLgMlCMZ7gPbVTM+DFBkpN678UeIdB61PHoAqOaIA5RoGj1gFgTz17KJzfkNU
jg0oWtLwdAh4/Q6y0xWaNpDCYXpTGeaVr84nsZnGUXnltt4kQ6He1LAHp5w9Hgjp
oI565CJKleynDcHmCRbGgCZtywYEQCY/MaA1UGoYOfcjB1393xOaOw58KyeRtiEd
TshCt+METTJlgyfXF9xr4yZIzmB9Jibxq5eQEzJwO0USJulATuYAO1JSmwGWlWPW
nnRAFZ3z7aznDdxHrp2w7Zy5XqXhRd8AMY1WKWfdZ4G1Z8E0IECdJXHWS5HeJUN0
CEwcqt4IQckJkuEK1ZavpVSNBkqfQ6c1LWllRpbnN3d5V1FjfulT/UYp/q1+PT7b
cre2FJaFsz0TB8R6FC/FBKekP2l0RToAxQe+4HOyEmiB7p0WzkdO7/1wZLYjIxi5
8tT6y+gUmdg/b8S/LZSggbP0gGvQI0MqeXFDZzhRJjVdy20GXtx7/sjpcx63Ti8Z
uebp2KFyWcPgD6FqG/01T4Ek8J9a7ZunxmSlhJ3kfLE2+i5DXjSU22h0+uHZ8Csh
PfczlhYK5IgRJ2G5ae9wyiK2akKBgUt1acOhOBsOgMb56YF3XG/zoNFp4mCqskYW
wjM/hRQFcnQMXSF7K2Y5d1vpsqwG+dIpUsfGTQ5KNGx3ZITcRFFaHpYFGyVuIMk1
oO/WWTDGctdFAutlLSDRi3rPhxP2MozWDvu8YK75gqBimB+9injZMdkYhEJPYDAF
sgAhNE3BwDL3aIuPO5C2ryBhyYGIcTKtOigrMz0kB6q4R4yxyPsbtxah3L7mrIiQ
Le6OeV4ggbytEbhIpA+c7XniFXVJc6eb1ma9vfPSJO0bhylIQRsj4gC2LR5OWQ/+
zv9Gw3VWNT2b4ahp66GsXasHtJd0LsBdmIHM5Sp6lskSKbJzNCGc/K1IU78aHoQe
lkLtzqWGi4rnmKAr9JFgXBT+ntqTO4RQr7j9/I6HlJjhnSy34F3KBMQNGwZ+VVPo
zNEZeLw3fP5DLb7xSRH2I6CglW3/1pF4Ya/IW4+5tqF0AFr59MxhrOZNce3eEnFg
bGgya8ocFnj5aXPU3kPGjRhkEGgfZKV0oHslW3fRJ6bUybh5LxxzKTNPktRjAWB9
2UbaCgn3kCcGpNRAdHjZ1s9S/AhIpirtEzyH8aA586opktX4aOtV9nBA67cT2U4y
+4NR6S0WmchP37O6dlttnNwLF6oZk7xHQU/TXGfnnF1VXbe0yQvLR+tglH5Mz4KS
0NNDwjDFfgBjF7Fi/HqtDrsP6qLjRrkeSWSo8i67alUC6Pb7kMDTHxvdafrp0+NI
VAMaU/9qyKQKAlJfFjX2Lnc2p0KLV/uDnK3a5mmx1gtzGBTZtcbS4/k4pDU/X3cn
zY1Ml+qPxTZFd1+LZokSR9Zw2Y3r5VBm+nEM77NHxUxOAeXFlMlDUJEvlncuAGHH
DAC8B65Ysog9EcPxWvxMdNwPTTIStrN+ZouaUJfZarFRs0GHJCTF23AnWqJeJ7lK
BY5msHR1G+l6EEraMbMXp6AAdt3FzQ2YNArn5+EZPb58VOHVmiTgMBBW25SrfHoz
9WMhaISLEi3vTMhBM4/CZq3GJ2B0mX8s/g5o2IxhyAP1lhA7McPusmhLDcDYqRty
VcTuIY3/zhMkxJPrNmNENqQDx6A4OrAMl297DMSunSWAV21UCoJSWwJR0H0fsLIs
AzBVqXGEso3YIneuMUbaex8NyAHVxkt0bLq2DYSr9eJlgdThbceeEWzrmcPZc5YL
ruhDjfT8tLf6x9qFfnY19bypypu2RkPWI7UcLrbh/EXohZ0TsPHfmeX8s7mzGAAR
MJsRLroT2b4ybGOXoeuHnmB+ngP0s27tmlMADQ8eNSR9Ur0VVV/eWyJCSGaB5Hgt
PqQdBOIj8DOGGCXbLBg6JHhmSyKNYIibeYBpteJvnM68/V+/eIVgPva6PnynGdxl
TDcglpqjH0VFJ52S/KheIGYGEedjjHTImcPCSdrdeLg=
`protect END_PROTECTED
