`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l7bedPZuaaOGl3ddII0xcP9J+PRsMAm1DRad0hIXcPyL66mv9BEK5W8v9TkExyP8
W6nMXM4jst0zYv6cDddxELVp2Sjt9sgROgJjf1j2pZ9oEhAN+axX3mkecK2tyU2x
zd0mY+26kEFkcij04Bb1VwC+L1+9APgdPP31Z593bDCKdXXrYNJ+x9B9ErZL1X4y
FvrtVAeJej94VqxSzu9bpt3xtPceV3CweBgsOnHylM/9AktJeRt4cG9VGjd1VPWz
6U44XZCaek+TpMEKKWVjE6UzxWJ0YZ5sTFSemRL7NGTTnEHDEHPHKds0n7R2iHNw
cIQ7x15bdVnYopgYAxG/7Q==
`protect END_PROTECTED
