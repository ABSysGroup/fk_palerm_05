`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f4CRCzswdcLimBb2yAsRt8fWLeeHi6aOWBBhX015W4vBoSDmiyoTeXgbkz/+pktG
CKmL7B/4Bqdzf6HbO6HJZuOu61DTB/OQSOr2JcpVZ+8Ks3NRMlmK5NJWALeegSMR
Fs+gWUQrGRrkJx8V5sX54jTrt6qRaT/gWa8ubSiQNIl7GX6Z9VsZv43nyMTGGbqM
btTj1xl05VCKplM/BnOnGwzlZkIi86eKR3GRHFnFpyaUiU9f2Sim/T8oUAaTTpEw
1XsjnI+JX2druae5sNrL2FsbJE5Wh+BSMMlcuZCzRYpSPdRuwWMJhxUYGsPbk6QI
NRXMgclWznCOAVPYZB2M2eGTwRr06MJ139PsgULJoD3kh2hTJxEvD+AZ6CSLFULM
Mdn7W98O8Y6DNK1Ra79ckaBCaq6GRJc0JG2/0gypaFnMDEKNEILxe3yH3S7YVZ/v
pYOjLk8lXHrgJTGcKbExUbGp1IooPkGy1QUp3oYLZPnZcO1xeQR7YV+QJ+lbIBL/
qyT87gAhTrVNJW3/+yp7lmvuhfUe4bPdugKCcUiYQaO/+cO/2nmNHVlkzcpUuZ0C
OyLhAFwKVzbE6j3iyfEisAFn8/SNvj9xlR9I7JfhAw42umjElrVAg0eivgoXqZso
SyvQ55sL8+wGKVUa/jl/jY6ImS0Itz0+2uyFTseDgteAyzpW1h4TDLi4MXdCYoSO
mSln5suOopztgP+BdykK0rzZls/8GhYrtT3m2nadTl51k+ZPnRaOEboe/LPsAG6w
mdvIutdNTYCAlXHuwndNMkyRYGhZ/ED7pjobfJRVKP7MRqIJXDHZEoBc7AYfln1g
RR79SaD2buyZjIFAGnJIg6hv8RBtUkBRWFIi2XzXSAv+Q7sVrhtsdu2FfgDxyhfV
BxrUV5JhbLHJuvOjwNqhJL8Ou5/65hmo4E6RTeW/0nGlRlQEprQPwsVCTYJQ62eR
e3tpzIZOkoD48G6ZEM9mO8UFMMTmL8qOZG+eealE/MRTBCqF3OtsHVwl9F89OPqk
+LMAaLb1PJE9S3hjQy6/HaHCXoJ4J86Z1Xe1WKQLD8fjXuPXNfk/fiN4vnvXqtPk
sYwcaWG8YrIaB8o223L2TDZNE1173T6OhVZDl8H0GTQGwFahdtX+yvo8cZM88u68
hKGjQC1LFeOgdY7T1da4XfvRtYODZ3Ej2vbPlNME8UUCHTckKuCeNR1kz2QAGDrl
hiNQarZPgGyBISL0xaJcjodqp7QoSf2VFaJhpurDUmSBRqpk+eQ0OOkWRd86NGJD
`protect END_PROTECTED
