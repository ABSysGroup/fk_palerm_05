`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MoD9wk04jAUMqc4ts/yzOXspZ2meHOLFCJDlcF5tLcXtpJCMlc3uGmwCdjX0WWcV
LdeU2JnInO7bD9HK3NHsqB00b9QClD0tT+9fxqoFs8NVVMbFZddYAvMnd2co4iVV
FjoZJ6ouaD43ZCPUGciqoU79uo9oFzVmxqN3XGaROAi3GmvWtk9bTgc0/Y9IvwZa
tVgnfHFSZrhR00BoTLOfQMb3vg8tXgefsVnL/gpjbKi6AUD5tY7cG4vglmEVScnh
H2026iAa9M/IZz0KR+lXoe4Z7ezOLdVdVAE7cyLtrbW0U8pH0iWbqtN6K0OUeiiD
HbuP4znitr59PMon9nYVdhCvxKkruewhaioBChUv+7z/Wmzi818TeA0M7+P2zkcs
zavLu0Ba0Q++71SBNwn71F8hOCsdtC5BqMbH0n4tfAzPattgKlYQDZr763l/sO7L
tnUr8BTD2WiaxN7ewkSxM5wwNXlChsDcjHrSaPHoQ3V88aTGVJNdI2LiKUL008Q0
DG/4XIqLUF8ZR77HaSu7dtEN4RuPvMk4FPADbcy31UDYmYzsvmSVqLI9WMgfFHEY
mKcZOSYaMNtcPD3kCa7D2t5YxhZE3eW89ajZ0xWZk/rwNLP/wUdK7+TAKvREGLMs
`protect END_PROTECTED
