`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ctcqkx1vnCcmp/t89YQmF5gU50KkRtiaMVXFrrVo3ePMV7GtrAZurwZiKAfj6Q/3
CzuBg1EYeUzKFMI3wjKOTHfk64Kcbn/CilGIR4U6cPzmWwJ/+2YgC4C1k9yFlaO4
b6ojlMWCkV83vxXDyaGMK9dKgOT40u03pZDoYOop8f29ggtHG7JzqsnpfOnYMEXX
7GzuwDkL5NZSNDCGr+STmam/A2b+S5XXUdCAE95Fi55vKPkX+5qPR80HaxTE3lxG
sFmw3255zPvNF3dd/KKZsJ4vjZbyycRQ9jW8fbc7Yturxk0Hl8l/9embddfWWcrW
T0PDntIzqtJ8gLvyI4h7dBUmDv7oBwqQE90a0FGKrRAzv+d0NaDGOnVxmmBWQPyG
+c+8/9O4p7bFMZUyFCUhwHcDIBllA74SONEkF5Ay5CaUXmc7MBUbOh3OM7UF32NH
Z891/koxPWPjXVLl2bB1PdG7KpECx5se/WJsM+irhGwaStlL4q3eCoUTD8qS/+4R
EfB19BtVZtVZRRgfvdEI/HEwH/e4T9N6pkkuPy9K8/2iYhDdXR3SaYLZRQQYpCh/
9UWO8io7Ok/EiwpZzpT6rFbpZHOt+8fy2Ks+6avaaKoXZQlZ6LS6AE8sfAxizgFt
IEGIlYEMzqu43gOilh57NLcV2Sm2TU01QJSeLuFdwRv0Arb85K3m5C7nKTd/vbrO
XameLUix32l53OzwVjKs+cyMJPBtoboLMiUVlae6w3TxBWI9xr8da2d+M6TWIMrF
7BmPXZ+l7CYk0r2KjvV1wsH3FD6iQY26emQqaXy+OOxNkgbQnyVnHZIcXQzpjckc
81fhUM2FxLRGjdgT6VYiLhg6m66jWf/xiBqpTZcaOMesWdsEDQRh9BdxJWe8TdWP
D812D86+lZZ73tUkIWvYTmHcCFXnVtJZuc1qfRlM4SCYN+c18iJ9o30phAg3dL64
u8CEo6VtvaXeN15+8Yl3cAPGLsRqXpfeNra7sWbybof6Us3a22dyd3SDxouCcDQx
1pyh/gnQxbubp31Iux14BIvcFzfaY//W9HVPoz2QYdS2AHkAqjyHJPq9ESlipGty
zcuUUHzwkm0hJiVK+k+il0bDUBCmb2JvhDr66HiY/73zEVjic11Xmc5R9LOMaq4R
8TAcOU1oAgSir5oqhdr8iSu7G73chHGKoIG0zRJZi7UiwauMTnQ1R6BA44pmMzf0
bwR7D5OW+hVXowG0TUvF5cnhiabG50tSYwpoCgcrJV0IfUsfW7Thm57E5pPYfFSQ
gAzbydsfpTw7jdaujuybakzKfp00L//D9KXJbCjSn9d4UeLhsq+IpOHE7eiCEr3n
Vz3haaNZMizab31IR17HVkFz/sEC/qsDzkoVyZ1HPbXPTn8mJi4h46lbhI1Sim9j
63trLY31ZgNlysZhAcwv/m0nZ7rKLQg3aMKlH8d7/0rUjuyK35w73c5efLGLKWim
LjQ4fEofBdTT8EwVP0cfkMowaL5t8FMZZLeUAR3n35jJe4ky1MHAG2e71EAeY04k
y+tTK2KkeqQrT7u6KbqotkCs79+EXXM4FaOdZfqC4mcTnXnmGJGJ54lOfr0lEJOo
qtPklSsKj/6N4Df0Ozz8k32+NZl6JQi+cTmyAGIQNpgg1pf/KTx66EemPUprn5QY
x+0qxfjTZtK3dnkh4sQlA+JeEcgS7txjJEf+sHsJyUWKc1sg48lk4bE+CghgpzU/
6wvd17KQqVcjGPXCfT16fRpuUOVLsPw6T1IpwY4XYV9TTa6Ec+C955qXvhe8UqVd
TaYSDf5bV1UO3vWJHW/piCViy11jU29tUlmvSI05Gvw8gXcZqd6eACMJHpLTL4JL
7uVsiPHSdvq10lhbBulSO5HOPPMBnjDcGzpsHeYjK8tJi7TPjlb8PYNlvHhVN9st
519e6W8AqMhd4xQ3h/NDYjH+AJ1RbqPZ1RmwD2jUXftwDEqp2LsXUbbC70cehMDY
/ry/9tU9qL3o185YNNi446VFJGEOamlS8mlWxg4ymn3Ehr7557/PNJUexcQxQ+rk
+YfT2jDyJwPh4cusjjqoEM2UBAsKfHqn6JzuCPNU4dTnj3Ky/5psDaTk0a/X3ibZ
2oyjro5mZd7zn+LNAN3V9WzwiKhXQfbVJ87vejqDwJqkbRa2AEkygqrcBWA4CATO
8YX4r9xcCr4I6GzNMLpSTjmdernDNeaRk1NJDv1rsQy9/C/i+HWJfLTFHgJPDNJw
s7Xy7X8eJbJecriwPAsJ/C5fUR9N1LkWCJQdwVESZXEyZLvBSaR9rG0/VsqFs5pH
MjepJyuWsRsk7qA2qIuzTbFrmZqnKYjIiTyeBqhC2qTDCn++omTU9I+ubDfvAI55
uFMNkFhRBk5cvSPhymjjufqecxhl0A1+3F1XPowy7zOcisSZtXhDZw59WvPErqJh
EVlDm1Fpp9Vwig1Z4VkbkzpNT9JpeeUUaoeEv3Ais9daqvAnHUxfbppBMlzPpsdQ
9VyoDkaeGrdCTiRflVlwUo/jW1XkknBtpY64eQKUtEKAXZYoBbwXSpcJdwjc9xaI
lybLK28qq3M31YD1tGVyD8yeaieew+P2dYWe0YXfo4hTOi36T8K7mhoM2TBsR9rz
JQx9DU8MB/L7L9XIHaoVr9Hb3uAXQ0IYV5a/71xZegeyVSvzLeKw/Q2sIe+Kgjhn
V4jYq8wED99dxEnokJY94ZTm4S7q2aTBJabJ8To2sxbjEDC6ZKaRFK2oHXr2XihM
lObpG9YFKWH3A4fSjW5hFQSbWXfjT5f6MZahTGvv9iCPTXmRpF5+ePfO1qgj4J4R
5GoZM7DcERqso2JaKAV9fcWazdjZLtGex7aYhynIAeZUlu4L+0tvlG7pEOVblzL+
pKmWp1PdvnmwKP+19csHSOMVHBKqZf1ElZs1UuAZklGrFzw/SYLwKrY7mGvK0NsW
TxLQ/HMNcukFvwOR637Z7HmNwNbiUmYfOqwMyX0Wm/Mbf5+STiOUNcEk9aiNcQG4
P1cmM7kiCDfk5oqeNBzLUKTeOZtsy+R4Uza5zix5daT4rPhdTcsegMIPXCCAjL48
0X7tJVpWTDRrCIf47xv8i+88P4mZGhoQCkIi+2cnjTFWZpDN+vHCLndKJsag1i0B
8Ko8PZp9fEh1a8z+uUhKcHK4L9tibUtcWfwWjnw4g9w1Sxo4dfsjWKo5Be7CXsvS
`protect END_PROTECTED
