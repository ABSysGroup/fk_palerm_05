`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fQ7tSUuTMW/fL8KZG1PvC7KJjVYcV2GX1tBpGEBBpYDvOBknYm3Wbphfgu5L3Lsq
zk3VApGGbsdtihYFsJgPTKSjidiguDDTitukWpXd9Fyu72U6EVY2mAi8DtNElxLg
J0Hg4bza4fXzau1pKn2Fzzz2wkFhyJtjwBupTGsPbJ0YUSSK9CWetxmK6i8laCNm
yxPw/3zm0Q5LfOomp5z8hiHZq5Yn+FZPmKxrlGuOj+FxuucxJavI6cCA6KJT43Db
mXG72gmInYS3wcY/gq5TFlX4Fkj18FF9Hg8FlKWvjQ7fjz5cFBDDZD/iua+ErW1y
djrwV/ytQbT44x8aOB7VK/BjkjLfGTnQYgBtZ3lK8l4=
`protect END_PROTECTED
