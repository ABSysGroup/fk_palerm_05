`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/7rTa4sYHT/gRxxrjKxr7CIRWDcrrwdCeQ4qm8AzCZ6CAeNq54eTruxEtg6F5+Rt
FNIunQzfAgbsxCX590Yxv4OeViy8R9jVOC3VWYH+8meWApL5haJfmc7hXOyYla0/
8vhuIr3wzPR7CZfy3Gh4G4Gx83PmeZFTk4gra8HGtCryULveZLQh0kpOPp6FMEgd
u8H7H814nJkIBXbzNrwKq1qvQ8TWNMM87yl4LdCWJc3VVbwYlmEywpfQHvb1VLGD
8E6sC0+pUU5L8r8pBU648vLmpjHMIpqM8HQoeiDq20YeTQhsTAnCfsjoMnFdnwz7
V6z6hv8TC65vtLw26hxl2pcRmwhw9WQAl4Af2la+VWI6bL9xE8CUe2iso8TQR3/b
kHes0b90v4NwG/a4EaXFSF9+q+USrjhfFEFNCXsPKYh+Nqm0c0wmTBFAkTJGHf0X
5ISVFYu/FfwFFAH/Ci1IGGD6qzWPYLmUUScS5jWZk+E5GGjFhKy/9ZjJ6azA1LMF
gM+dgAhACuYhe+GW1ilgom+l92xzaDDF/tXs0C2M3PEVesrUecinq1EG/ekHp9g9
5+tLlnv0yHha1WqtN5vgO2OnyK9mp1zXNRvidYfApsNxRl5oMkFei6MInvUhe2QU
5HITnie+MQEAwjlUAh2IShQtpguRDt9sbrO7IcISIWNhF5Bk8G3uWbjlivfwClhZ
l6Zk07xtGg1ykky0RR4gROrjA/rFmNi1EeKcTWh2kWo=
`protect END_PROTECTED
