`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nXMx/PzEBClDNvr+fgq9Qb+Sn9Qe9lX1W+9XaBcIU7ojnLGTUNgdd+sgtH9ksGD7
WoeBWRLVhtFThEJN3eqTB/6aYK4FajvPA3U1nstWIm/9b5Dcody5Jd94owl4bs7s
6NhzwI4JeLlvIRg620XLW/CwPZ+hON/2MAm6jp6E1kFTJ1/6nwsb02wY6Dl0ziQt
WA6YBIbWXytWBwTRtWpgfFZaTdpWBSDJqvJq5aReCSfcPyT1dp2IhbXfZrkUtLOo
4TytWUODTuP3KXI3g/TB9Q==
`protect END_PROTECTED
