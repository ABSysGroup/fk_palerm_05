`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lR8M+kvSRC3CVKX/ab1OKDnbWsDGOOpv4t7Azey+A0qoEfZ5O3Fw9T7LyfjHO4zg
xt0sKzY66u4eUDrlc7KiFx9WQP80Rd119qhkzvbIQDyTp7116I3llBkfCtb6PHDA
W3MNOHJ7zD3DQQsL/C7Bx9mEdf3MkNWQYKW9bClRZurKYZrMCixqWKlLXzGCcKrE
VzslBu8eeCegl4VvcdiUdpyfbIi8tLg1MI13JLC6yDV75gnjxONj8MXVUTPpa1tD
217TjQwPg4goYkBO46hHWKXkN0sS2x2hrMd2E0dcU3iYsCJw2eaKvTG16GBNCftc
idU0epJ97R6msfP0WKv0so64GM7LQAru8ahuAvLaY+g=
`protect END_PROTECTED
