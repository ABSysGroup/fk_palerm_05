`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qs2Pv/i3cI7qNo/YgZuxXoo5KR3uX0JLZ/T9EgY4wWKwqjqv8aO5jd3/ivGcSrVD
2tm61SbmoibNZtSd6DbaAvzNuD2MuoZASbPF7xOo5XBda+650fq7yuTR33yZepn1
llx3JKafUVJXDTMUUi7wUXqfv66Yxg+JBuRFYo3IHzojUWXSk7P/zlP4JIzly17K
HTBhkLh1KyLx+Q/zgu+NKUHwnA8PRf0ANXgTpjl2w147Ef+CyYMh8HZhEBeb2qg2
J44nM9tn+kgEt0otUkN/WB7/OEsaqZL/Jmw835uZQX64yQ/SmlhedM/1sCBYMWNs
yVMSFbrVJmpcnQYP6UQkst1P6oBenzAhDd0XG6HMk4xmP1Yo5uSQISBxqgdhOPgR
9SrOyVC291uD3fvh/madCcDtuzZa6xbTzl3Kfcl8V4HlW/QwAAayp/j/dYw5tfmn
LWIVgLXwI19odSD1EYwAjX0hOWMSaGjn2Uoq78nujnJj7HPFzveTE9JAWJir5ABY
bTcjyPE6WkJLa7FdbYYa+iaMMzwV9hIf4889kCXIGMdQB6xI4UspNIyR7wu3lFrG
F3lgA25qfTHstbFoK1IBV6Q79BWil5G0YroLiA+dBkumBgnS4O4TEt56GF5cL5yy
28w0rn0HNYotJOeoCgFIOuYWoXlRjgjLdaWK+2FpQgj8LdbEAUoqHTLJ48uQ0hjv
ail+z7xmTk4T3nbBomIZ7kSop7Kc8jBR5vSt89wVnqRdXo5ozHE2X98v5iyVPRHf
FPbhTUSB8eT3LTNdTGdFH7bQ6o22QH/IjpiXySOOSC7xpUhCakuHY6XkDHF0uQwN
wKe9qOCJkQKvYEuiKseNvdVfBzEztXu9XInR+0IHU+TAyDlf4/KJy3q8qnKkfFwW
a2Vm+zIS9JLWqhi706ghpDEMRdGsQZ4AXvEsik2wIpVqiutHSUbo/eoMjGC2LRGD
1bPnHU3pGd3vUuhrjJX49YiAl0zwge/UuDU73NNldmFygDTdBtv8pB5Tp5j+V1v0
`protect END_PROTECTED
