`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XUB8E4iVgPrVVp1K9OVtdzf+KT2ekzwx1iso3KyKMUQ8F+WIcYZSWQ00/FMM8NNI
mpUg160SiZB/dH7GkLZY7fc0mvOZc6CWkiQw2kQkEBUtgZpZLDwh6gl7DhGAD+RL
cUx3jWymP1uZhCeIKLY2cmig/th+RWn7/3crUiVtGL0Dh+Xh29uf07Pc5VCQEnaa
ND8FalnlKXNUaTBFRnERvHTV1ma69s4loT4zQBXpUOxJOybqNRF54pYJMgVGb760
91L3KLRFyB7kQUZPpVB/Y9dlVzJ+uV0BtAYS68iQi70KaHJlA1CXMX3xEJ0XibyG
kYa5kOi1I6b6NTdnXoGIAAcPfKBKZJ+NYhkbonWaXoqK709IUe1bw3MPgyejXBUd
PECFKmq/V//79mQC5McLJxmy7IJ/YBNx3IAvNPs+7L+mqU6ZP8Fx3Ii3VmJR0QN+
O2KTDy3iWPC1lOvq3y1knSBgm7+dTgSJC7BL0RzZASKYahi0IUk5q11nLe4KH+b2
iBs6xn207bSg1QW45LqWB69wuLOxOg4KKQVktS4RL1txgNXvUeYrXAW2Hb6lXV+x
w9Hevvb93p7kelPS0J8WzwjGacXAJJvCby+oOCXgmwslF+iLZUUyzmg7Q0Gn7kgI
VqeZW9EaHZ54chy0G1tOui4DhWjbcAKBbWyTq8R/KuA=
`protect END_PROTECTED
