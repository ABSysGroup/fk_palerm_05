`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nk2l6ZeWG2USYDHIIf+ktdY0g/lLDwj9CownfLwb40DDeeDzpJc2UZ5apzpoHCxJ
0sLHxRUqG52czz/XBlgmlAKbuZf3jGweAu4O26B5yk2EMH5Sh8j9/VXdjpP6lwng
le4ZJe9BCbgCdWr+eYytANPueq1AE7vN3WypY4SPxR63AAoapsBVS06GU7hQY2Rf
Pa84aqmP4/bTNlyrKBW8hFIX73SyzPbqIFG52G34pujzqMwvfoy+V2T6twcH2E7d
yMN1Xvs5V0BpaFR8LSOMXHtpkyVmD6ExvgOANIWz2gte+cSZzo/dwdQ2YuhCYS8v
H2JeVP/hN2Cifp6vBg8etUpqfY2vMAKMcKGVwQTf46aR1NOn8zX77Wl4I0P7nO1o
c5DvYFgLTC9YXsjvcf64YsewK5eNxcfwOwBSSWu/ft4XT//6NfpjucCbCp5+2ZHT
VzINTuGQuN8w81Vscq76d444jtdwPj5XL7PVmnd4qt18bUjUv8MLZmeyALGb399P
s0dkJ3TrQehfttI2Qv7w6qZpDnpFBmFCXRd/6PRp9Bh64jNI0x/N+6Sdj8NiBG9n
Q6rr++bEktfgjFgWk2TcNX3RhaR/nZdgW+mXn+v8FHOxU60ZUOLcH+W0eWey1V+2
vDn4NJ0CdNCxqCMri5LS7Xhpr6ngw3GNq8NaVHTb827xtVLbWCyxx2UPppXwVskb
kxJBJJtyqUMJai/iHznNaQ==
`protect END_PROTECTED
