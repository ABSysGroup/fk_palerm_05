`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fNQkbsPxU6gMJo/AZTrCY0e8voHA8W5rnLuQgQQRZ9fGEXEv0l7v5yssTGuvKWS1
EaNgxNpwSOY9PTna7YcjEQh3ezKb3+JVT/rWUnYLHFuIdZbOBC8n8ClfI/hccJWB
TNgBxnAE+Jv2i9pMLYo7qWHqm/yV4TagEhGmRzQAoiGzmeS3/TM5N89mn/8LcPx4
V3QFEYhXxIf+DvfVJb6UfX/olRcciiO+rQK9qBDUHakMoY5h276ojSl7yrk270+d
tmM7KWr/qwlBVBiBwktdVV257KfxbG/wuWkRoew4JYrKv7IwEZsntiP28FuyvwC0
QPxh4htsrK0jo0Q2jkjIRi8xHsll8xMLWDsMxLpi9oBBrludG1PN7PFaLnFrnYHp
v1iua+EU8Gf9mO9d0X36ykOGbkJt5a46uj16qfVnxpk=
`protect END_PROTECTED
