`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oizVT0UlkXurSYqu+MX59ILUpj7H0isFe7sUdvlcoOc6lD82DxZLLtoPxpMIGLDp
gZjldZtPzkIDus4OKZ1eBzr2e0jS2It52RWy552dxBbAMBGQ7vXZoy+P1izN2WBe
pZgUMovTln12zdP6VUaLTry7NxjPrn92i6T0oRFTMs1q1qqGqKQ2cMoSgc1ulFAS
TNVWyIK3K8+0dcnuDswmFBwqjJnkedM21Rgqcsmfk1+1dDTvcCMZxysvl3SZHet8
ZBAhfjZzYIPyD5eRv4If2Rpoj/3dK6B6xx3sl8wno4OplulamnkAmSk9rltt+/t/
VvvrWGLVFWu+V/rbKPS1ROmtFsvySuLGKwurWnXAzBUwsbkqMgn7yzHltioXLI3S
pmExtZP8v8lyUA85Vjv95qe2c9iRMJQxIomgDB/smPVGGLPUSfbvuQaqluxTQBdT
Qj1zrOrLURVd1sTDYofpB15+mSpW0fHdUgcA9ft+uuswqNhAaWJLsD1tyNhcJ2cb
ov876Z9Sx1ML3fhOqsOhArAWR7FHN4cfhaYaa3GAr6dKnooEk/lWvmqEBy8r1eKA
tKJRkHpE1mKLLiLyOn0+u12STR5HwvmZAJOCGI8ZX8KW5RhZI0S2ntlCvC/3OOTS
pZcjod7rSP6VzATp8dW4frkNG+npRmupUcxnSflad0VXJ5CbKevVnSyEiNYpYGje
yq9/yPN2sNdcvNgbi/zgxCRdCbwu4yBxUXAhgp0KFBiUsYfsaHlEEHzyq9qsSkej
MMSI8oEqAzyD8hUg7GRwvPLB49QrLKcZySI3WsyLYRM9mYNdme0Qop18qxtFHMso
RQ7+jI0Ig92LrNtuG7RRAw==
`protect END_PROTECTED
