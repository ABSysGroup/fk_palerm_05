`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZErsDPwG4njjg1Ztr1WaKWQai5BEiSZtk5n1Y6DwTj7s3caVUF/Kyug75HVKPYGk
EoGN0K7sskJEkut0lZgOdcCVUNrzTwedpn7biGBNfFAKHIK7bI3ZfKnK5NWlLe2M
nXsCFz6Ku7Z8nSuXBjZEgFFpGveWlQ3lrSAG6J6PLHADsycF+SCEqh2M2aTBss/q
H5XDl9IlFD8ZgZ/FBDWKjirVKouTKlyIoAAobBDuBpGOKJO72dkJeSc+Finyd3xJ
l1NRHLU3vw0Cqt4MANVkdG0tA6L7hcKCFRxG3HYGFaWE0zT526L1DQGrlXXRjECN
RL+V/QOzxZVf3n1Sa+1A2pBUHIjc9c5xWQ41dLhb/M0/ESw0SntIrElFjhmMg2U6
TbzyXmmruw0n1pQWnpqXiiIGk6IRvlrGVrRptLYOXNHRhMSEVYGoSf7oYjAGAm8f
75Kf7NHloQQZD2/+10ueA+Ni6voOsgWVcAITtCzJLi+/xZSeTuZL1v7YT3v0Nqqw
E8ewEYtXY1nk67lCkYg++8dxOFslAiyi1ch3HhVifNEDTX9kEmskPyulTSTZ8K9p
`protect END_PROTECTED
