`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3CPpRJc2xwyvvbO92eIQNv8+Drmk1MIOjL5vmANZAP11dja5wprR1TDv9azAcw/p
nJqKLeFKHNXUZxzKJjLJqf++sIxzjB0aJhS0LH9ZJmbOYzcs72L2qfwVKYzyEdfg
fRt+rjtIch9sqY5+1vytSqMj4BvKvd3vA+yBu9byj73jPnskXRJSuzQSrlbNlBKM
qMvW3JM5gRvm+ZstTcDdLnjbbZsQAaI5HB3h2mKx4/UbSQnd+Tem34I2AoHTRzi/
I3FBFHgx3N2iQjG3iFAT1eKsatYmeHHF0C8oWkZh8ptifUbkdORTe+VzqL+r4nfF
dHYuGceyS5p/vBeOecZe6KZxM5E6d128U7H+6sTYDfq76gTVxIUK0btNdl9iw8tk
BOOPAZ4GqKQvVQIHl0gEg0iNllWsmC1SDxhUbe0ZiO0vAoED4wDHCmEPfhGupIOZ
`protect END_PROTECTED
