`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KangfSPUAVAk+T27oIrWmhQAX6goiVrnA8xsNp2z0aM169UtBwvd89qAtldX7Z46
1Gow7ElWUHIhMHBujs4aRkO5WuL00EiU+DGN4oBW01fi12rZjMnnuiCE0y9tzSRY
Cpk6mB170xp9Y6RZXdYUXuk710goNGh/1jEkuC6/HMdEKU1OzdSL46j92Q834SzU
/QmYiA+5h7bt7ZVLq0RyivprlQZmI7FRPToyuurPaoq6F/mV/81bj0uK3xvhuqUy
9h4wofa6tCU+9fpaVp4lRj7RJRAcX0FA7lbZET+MDHARPJrKrHly7DCIunSKoQ8M
PQsLkncgY5MvOPTeZlVoj6npBi9EGrMupuomYzafnbMsQRcdh3pcDBQoefue9BZR
H55ka7B4Hid/zmGb9FF0XjaWkADEEZzTfJrz0wdx7EtStS4uX0zHxILvYWXW+KQ0
XH9NY0YmI9VC4xUsPN1SzPPA/KTGmdcYU65sSR5pADrqr62RJC+jm8GvqToWDega
GaaPuR8nXukcCI0AUeHUQociOMjQ8ETJXRMUjbmut+yCPHDvvk5IgSEbgdPG/m87
vRnj+Qq1Z5CYpmQFAmWkL+HzBVOq7xs33kf0zh7Hq4PinAA6eMsFCZLnsMqXKfIL
3ixf0gOK2Fgzkj0nmac0JOxFJOmw2dbPTwTdxu1BQljKMZ0nVtvByUA3ZQ6YyWrZ
accoWoloSx8PaFO/4o934XibFdYOH6wlWu79awSp9iz+WfU3xuMJDzfOWpweiXRm
l46ClQHBm2dBnUX/X2yWgWJuv3QfblxxKCPACMmhYb1nkSewp3hi1oA2TOdo//OY
`protect END_PROTECTED
