`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jhCVqpOkQoibMAJWs7urWukKD7hqrBeoGVeBEVQGSK0rxcl3EewjAEt/cXM4zFWS
8OO/sjknvjpkfAbWJmilc4BYieHvEenHzCIH3LM1j8kqP3fhxYTN7Or0YrVfq1wu
cJgqcnyaPJ8uVFzjjCUpO4ngDK/iYmcRWQreMzC1dY6Dqexbo6CIZ6mOZEHtPncp
4ez7YCd1iFXQlqOF76VDNRPOuqcqn8tjHt7TkSMLsgMATFr/usq2UhSJbYZ2veO/
288DfmG9HNnW11xIbMTJYJXB2VkeSACBREs/4GiO9n7Nk+UitlRzoPZK+HiMD8EK
p/3XuTjNcIiPOwGlAq36ifaO4ErN8Mf8PZJXC2h+vA5FRXRo2SGMTBZz3M6hC0Vs
zbOmeJWmDuJBkC80XRR2dk0bU/Ze5lF23CHALTmn/TBFcDpgVtrK1nTefxuTQ3BN
SOK5i4M6RCZTLRsv15kEddiUZRfYVSPw1fWwUYUkw91BV+/fcIDfHmH1I2kqZ/z9
jWst/QTwmAkEjnNkLMtaegCKF9Jxn0GQ3F7bGNAX8fBuR4FhuXziNBeB4Y5L1R51
pQ24T51pvqNGX5aG69pSOQ+rqHSDE8r4jnbNoizhVxvGR+cfT9hn/ZmB77Hhp4Rw
UONjL9O7AWc9NGIxt9vjPQmIxQFFGpKLOoQCW3R51lhAZHY53J7+8nlIXpf78Q7l
GS4jXKPpPAwr6Foc68FH6fFZ8PGe29amk6T+fgGYSpclL2oKCIKIAIf7/Nft7/K3
HEmIVWw+q6ese1jyYyP1SbwEfmbp06HtGqiLu1jFaCLsfB/VU9rnvIj6eb1qPzqs
osRuF+kvInkrXOV1KkJsuFtooiGkhm85eoaKNqkzIjkYsfMRywPllVGhvuph+hjK
tr0sHDHZE2jGAgkpZtJZhKQGbWCJrmOyjVB9XU/P5QNWzDeoEfxfCtrq7ua8Ootu
0UCkUacjyO4XB/W/E6o2Pp77/KPjgAJXtPMNF3g+EZN7XnyNEM+Fl80RFWokAz8p
VuaiLUNTKb7MyKyTDG6NyN/aSoSVICY0N39Lu8tEnfa/D5WnclyvKO6qX/+/siQR
5fDP7OWxYbEFI+1v8rx31+U7A8EPsb1O73YM+H0XrJc2sLo8kqQOUkyyP5YubCvv
LUz3G3ijBbKPm3aGd8FtelH3iLPbEd6KD5OwmCIhr8EXdBvs34UZef1nhpMWQWcC
mVxWMoWqjC03nDK4IOYgJBMBF0oYbYq/nAHcplYqDbdw2JDLj+WSflkxsgw2wk9X
BySjqnMANo3vdYccE/5kFwL6vWb5emmFR1QWiY2kkYqrv++J2UZt1Efw7omnYTxk
e1CPb4D/Dy0+pCLat0nHVHJGHKVXfeX73u5xXTW3Un0x0qmBlKcSWMTacJ6K8t+0
qWwdDLtPX5huK0WCB6mHb+VjJg5t/sZbM4vlLEW3hz0xcHG+4lUzkDruz52X2oy2
kK3Mvkg84IcaKJnVu9l8vC3hACYtN9J+zC15H+5bcgH9Ew/9cbuAMcUIQCW9jxZq
F3SnleKMJqKZlWCqowPk49mEIzWSvXtENJB4tO6VfbITgufsd2EPGSnZdEEqQJeg
qWA9pamGvagDUbMwSzVB4TgQ0GyvMZvCgw+oHpcou3BFqL/dVges4RIl73d81nlj
F8TU9aHPNan2GPZ+5WVXUtYV9OIy/Ee7oJiatfyZGHVRdvfT3sqg9X3RjXO9/QUU
ytsO+3WYalrGBSE70R9vbo+lS7dLjpo/3o7eeWX0ErUc8Pht2EQdaOy6d+VGQmbQ
qkFgUpcJ9IsU02HOIDmxcTlXJD5x2y2VeviUgwEhtIh9apkqY0miWbODQfJ04bX+
zpxPsqmKBDMz/LAoHBQ6rdiYWRrOQ2MwLt0wOGwDUfELXxOdn05MNEPEcpy6hLPe
tp8qYz/QEaJWa6gkzpMrG/PAiZ3u4dOsbz7obku10SZwcc0S8GZ4Eit+9IOdfrIb
08UqrbWzysNzG8r2u49AaYjjCqgKHlh+OKsT+H5tBC2nl46SuuC7Uy2WeWF+i4Qc
bP60277si/eBm5if0t6zwdXmRfC+WmXLuj/NI3e8uQIERG/tMfPmMzAlKRf3XOq+
Gvry9SY+FQesJqgG8WJIwT0STt9dEGMunFbWortuUJQGpX3mAcZDS1+FBN8UXiSi
6wjBiEMJyDhsELlSq+k8CyP13tp0mWVuK5f9DzbATSFe4I5p3Cl0iUSl6YpXzKMt
P07lyy/6t1t3pPVVdq2leoVWHhWvMwbXQ/luBkcepcENRtx4U72fSmdlnQk56ytg
dTerOVV0koRYcDCEj98BGBKqsraPsMD6AiKAlrlH089XExrlJpACCvrw27NoTzto
hc2W5xsrL+AODiKzvoZpDeOyAPZydu8NYRO45i79cNU9WOsk969fYJ+BvykJbFw0
OA+GNxsoj0jcML4vFGXPXYHzG85VojPBixHc/ak73DBsEx2X/39to+wYCNhKpF5B
jPMYsYVW7gkjJSYSsmBfPLYUJf2v2GSaTZbYoAlZdHhOl0aVSm0l7FHqE45t9I/r
jybFicp9LHSYKWFf+QlhtGRZZc61JRGPW3NwYjMpQxANDta+86p9oFsdIXcJLDuI
/EgtuxAX4reZjCN//UbqC3BEUA07O4K861Z6Kv6rhuI=
`protect END_PROTECTED
