`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D42GUMeDofRRsX+gmG+jEgYGA/qtb6z3EkczOKURHjnVuIkIy8S4rJIcz7qotxLU
9zee3pdZgvvR2JLT0ioc2ykOyJ0VVJciZ2CAY2E5t8rZUJDmvxuVFW7v8Womi17k
yRX05klj1vWfGOd/KOcOx65iX5wWISpYivVXFraNfq32FtVGq2gGClvr19oxVbwd
7VltfRZO3YtHwZcbgMEtyF3+YdbSEIf42yAMqJVq1U6SPMmJ4SgLYRMoagtuYqZ4
IEt91GBAx62XKnlXbxvSgKh59dP7mcSNFEuNe6qnWdGzzkyctIG7w4CYwcNPy/uM
/h2rG+npMV01ZDSEEe/bOHo8XZYKzTYiEkYx6JujHfP7kBjjFw/eWKdR5Jkxbsqs
e3xf1bgz+7f3CrXp/Xn7hNdzziC2yvn9+t6aKR4RUm2R3bsM6CzPpvn+mG6BpOKI
kwYm7WgNvsHAFUXsG8kW7JyOJoIDDAeVIHx+yFEkDXB4WI6igN6C+VSFrGqWapx5
c7g6tnmvIwWdzxgQCzWqATabuJFbjHeWgSEG9fIewtHcgKqBbqXPG7md3K6k9aDR
YED1onSFbV8EHqaBeccGIw==
`protect END_PROTECTED
