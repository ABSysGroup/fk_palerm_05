`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xoYICPFIjL/yclGutEHgw5bgRFqDgBwrU8bd4XXDuzlSUhv2B6nfpS6wN0MSzQVP
GiYDGzHEwgsdHxhy3JxCN7HYhwo1MWkHuFFJ+ho+oAxpvxdoKCwW1L9Winh4o/wB
NpCaaDLUylDRGtInzxtPg2aPzICPFC98vblaP5bMB6nV0Sjxr7apGJcMP/pVh0nx
kEMKn7WNmYgCRo3P7dO1qiYV/QQjDP+hvFsdOr0JEdLXofV3pHZGjzygfD+6n2uK
3tDfJkVCK3U8rIq2gMwqSCLAoHf6CU7NQ5kFdPJlgkxBPN5QwSXiHdWV/AjFW2cl
djGZRf3uOerEwheX8akpXstryeUsDg5kg0vBVsZj6YiLYWrzigu/PokIgVARF+tc
BqMlKl1toDuywB+6K4TRBmezKbSdZxkogDJy3kawMIZJL8wnkn0IlYULe1/8qqde
iavNMn72QiJLY5c9zO/w82vQpjeCkokK2UiUnS0iBOEm7HAwqvjLpuUCWVCo695n
lV8PCHmGeaY2WuPm+kQvJLlilewbGvFehNqS9tHyT36a9/z5rzHXNpgc3UG1PQDu
pIGXz/pRuNIIws1gmszAgahsdzeGOlY3RvOBizDC+7k86yULzzFLbnUAI0G1ZJAB
qN40hMsK3noHE+hBjHElupL7XkTnZP2bRnPPvTAQhrdASB+1fVxFKnY7Jn4ugBK8
P0ENTyiu3sjqlf2nw1Wtt95zj0dMfsV546jMPRLoQQjLR+53F9EuLpxtVhXDzWHW
n2pxCntcC6COjH2KUoROnRVeQZ3CNluxY0qdftO1sGTpEooqFIeVrYlXKWuqgbQS
IuA61tJ4PVNcR9ukdYM8K/97gHUqjaqtVzN5sHx2pM4GYZPkWEc+aKTz66V9I4n/
gRytkvb1HQLxpSmitsEKVnKe27mKb+kquXt4qZkTtmcjciL0I8ARCuAxAYS1qNKy
5k/QlkXleNnHV3gse/eW5qS8POyatVOenHUdmZpIgla8luzdYYll0nEr25YuW5Qk
hvRjSvE9L2Ut1uErQkmNVUNSZZym+O3zwGm0WK/o7vHMo84/5AGkuYXp3s5/4/V9
INmU6mEchknEQFtP20m2L+lZo+DxXUGkOMeSSJYAijhx3ji5pnrbevzAjoYfEkeg
tbqEuMdkYWM7kllszAA8mcrP611ua8MH+pVNt7DkkJmWqzM157z+k9FJNWaUS3Ax
lc1wxEtU0k68+saxRQS0maz/v9jQtTVQPcooJYBGg/MGVH0aE7HvMMAlYLbitev6
g/WO9/9992q90ys8Q8gGyo0zCMwi4zmlDR0ioNZ+ThCHhfHkEkzyF2wA097yypGX
hU/tiq3wOUlYhATLvrxFuDylv9hX2Kykz6BgTE9WdRKhXY2WC/hG6naRI4KqxwWc
GKfnkk2DP4yo6uHnM2fHPlULrEhvZsz32cxNpz6ii/yz2qBZLOYNu3enPHNX/Ife
6u0EbWzX126AZZvJSxSlrsKxeoymOFx9dLKfFlziUFG3UUIgUGPDVm3sAhxEnHPI
7eyj1XlvCT9ZBfDz3GPR9Cooiisc5RPGKCczx8VnRUigM7O+VhH7yFakh96+KiuZ
6RcFOge2q/Y4/lkiJINa+tSGhaGyBF7wNqXX3hxVV16E9N2papJL0qvfUfCTyRZg
Tl6EPDfTpdkENLUWqXO5JHDzwOjdjHgLG74syDkwt5wOoLQJTQnGlvKkXHCbb+wp
B+iLLqlowzyPRqaMNJ5t7MYgiVYo5EfTdVod1Ncdnd+Ob0mIxGwdfw5KWD4C1b8q
mVhX8K0SXtJOGR9cgGS5IYMfAoRvndpe8zXB+91YQX6Di7aF+laWF+7WHaurWi+c
lGzz8cdi+1V8RFKwjDX4U55+wc18ud+FPG5P0m4u9MoWoEJd8ApAcSIsQEruZE4P
fip12mHGb0iZvSRr7oZKkK2rKEG5oOVsMlMULWR83gy5XwhQ0vn24kk4f5ymqMKv
Wh6GsWiipFvo7oGBDv4UB6HcZr4O6q1KVWnNVJHgsoWRZzm4slE280hpjukQt71Q
vnGesHOqmiW5BxhNNz9CX/T2x6d1AfNRTwNqm/HFy01NzD64kh17YE6D52hrMCJV
IWu32H8EH5BZPMt2hIRLVjFcMj3xYXe/AGsIIXbXcDCh0+8afZG6Z/G93zJ+Jn9v
HmzF9uasfm+f+yJbmmXHnnu9e1nt67KB2O98ODICOaM67pulG+iNOPczQonqICEE
Pw8tbMpr3QeR5stemOT9DVePVtS5Dt3rNq8P02ZJREY9GXuYRwdC9lX4QBvljzbm
BfdHWhH3DH6Ejw85dGTXt5sJ59yilAcxhKAa7dhilQGisI7q9vplbL6TEikHPh0c
BPwuktsdJApWy4KcZg4D6qgBXCKAN0t67YzF1R/qUjT6MQSLcUzTOkkt0HQ2YaNU
LGwVa2VcOBZOnncZJd+nwOpZtGPaxVrZdXQH8R2R0svPS3llZO2eNfDlc6zxrd2L
hKeR4rSLzlZiFzF8CEiEddsRZjLpLaQiOA65MykpczNtgu9P+I1NndRqiFSqqoNu
QGTmGfrnCJe1qHgbq//UIZ5JlBOLG05svkuqBAE686WTC5LanobpOiI3Y4qVLm4U
lsdJ6C82BcuSe6pPg2pfkr6WPj7bwyg4sBsTK0dFl/uqr58H7o2n/JQO+VXvq75L
j/lrVu9eMs10lFzNCX+LNeUEnYGCmsbHqBu1LmWsRTwTew7yJ3Dg4OWR/oG71qD7
jgY/Df4uz7NIY8b1PwvwTaJ/2Y+BpMkgRDndufhIpRz2E5QFczZYZ+yZXaGRfsTW
fE5ouhwMtmrCXXpW5h49gIxIkbzewsuzg0MmT+y+zIcvOMZWdCqB3X9K48gSxwqk
AMN4HprZqfGqdIMEb6Ye07LDCGAx8uqT3afywrfY6Hj3SG3XwrE9Yr4vpNWxNRB8
JGhemfT5SJuKJE98vnf7y8cTITPAHjxfr+CKdgqop5lcBXs9EIXRrcTZDsYpbiym
vjJpMLr+Jrfvh5wD2FBoz3kjMWCJLu0AfyZ5+EnNVLykZEIzimbAf6mXsRIzpQPG
MWqtNVcH/DhPVa43uHzw2Pp3KWwk7qTkoina9NtaGbG6PszrmRjCrCLUjQMFY6zE
FnW9YvNckLHcPOPxkrJ9UKczLs1IH3kSQiUQmB/dsV9OKMZButMqtqqnZ5OOADvc
lucGDt0nVRwUMG0J+hkNyc+OPQX8s6HCJoBGhLXGNbFMdlPqr5qi7BjSCAc2IXde
SEqPZPcZGVJ5GUL5oFAVpdEzskaGbC8YULu3qLIU/EXhRs4X8C0OTFrmOc7hrxFt
hLGxCeoYjbZog7ouCA0jk+vIGDE2ZhjRkhxIiclU7c572kAhsLlgq1cd9PMGzJmg
yL+Z3NCNALzRYSt1VSnAoPUiX5SXAOZf1mxk7gNwvaoQ/VxEV3fxwY46nqkrmAKr
kHik6on5hN3sOCXmOZCUxSmjk/Cob7OdEPq3VSvah9pbx1r/4PiN+f5aZuba0PmU
yOC9Xrh3BXVtytlMOtV09wik3Mhqi2UH36JCqKpLolRKA0Ln2m7MQUkvdygWvlTE
zJzEBFt+URN0E/OkA8jcBzg7AFJQZEdEhEIJkXCHyhrLhtWXNSXsV7vLDqYxIn0x
9s4E8OOSpqF4IIH4VUw9b3PTsINTn3WhKG3GHuFnnWc/KOMNIza9QFbF3yrwZ1VM
LF0BYz5+OFn8UK4qA4fXan9Q3DeDPnmdhaAM6CN7XtuwCuNHA94RzPScBipBI+Ff
xcx8GQJMenAHxpQ6Vv0A1qy+1rS6VxSPMi38b3/jM0tvwCNNDdgwaHuwXy/JaokR
SjeSkR5wTEbGPfaVbPIR1Gz6SJoHIf3hse08hY44Cg1lsnEpZbIEisNfBN//SC6g
yuXcKwJeAuuHMnsR70CafY5SHzQcfhLKrf1t0hrxGNci+5xj5slaGeMUxASlWjoo
RlT9GMext2Pv2yb24npZ2dIHhYUpUxTBMkn8Pp7/58ZbIwLKoC5gZo0Mg4S2i+Nz
dcfRMesgMLPKpv8vAqQwnFDNA6KWmI6PzH9j8lMOlvvC8OKY5QLChA3bCN4aNVRO
FxAHAz4gTV1x+6vm5Zt5cy0rYR3fanYcm6Od8yHgIQ25HNvdWAPAw8gcs/81Jfkv
DOtzJhjkHVjF/5Nk0TbMH4TO0YEgGT6tInaArBSjJhNGRIIv9MfyYaus2krmpYH8
pPyPUqJjDYxxsMd2ExmLk3cBP6WnXRoRicowNQtw7ldFGT/fMi2UEFYZ7tyIVN9b
g5lPjrFQlXA8GEZ07yKZ9i3AKRBS6K1uWJVYiIcsoZkbenM4OYxO5hYan8ptEwIT
gi09aiePfOVaAgiE0sbTBmEoIpaHyeCKqHUE2GiU+zZDpxZYpTCd73Us2Ihv0wY7
GSn91h+zabLD5ZFLiCGJ//MejQ2WjJnAM0f4QzjbyWCJ1ASeckYD186+veoIr4y7
S0KKWwm+S0WbJ5sjXmgbTuw2GhIlIW5SYu0X8npH+CO4gykeLYJDT95A3INSrpwt
C6IBEEyXIh9ZpJNfkfJTxsU2X84uY3kvLrCgBs2bEJeLgmHAD5ShMdhXjOrYnxbX
04V7fEMueKwC5/iXrqHMj+CF5xsIoj5xzKmOelVytrqKuOexLSnphj/IeJn4KOGj
6H638v2Ov3D592Xd8JACX2Fhw3EY76DSMwbP8YaIg+zJL0iB/buPtR73u9ckQOrE
ToP2RlvXLcyAREcEcALC9X0ndI7pUauKVj/ajBUj96voyXATP/ROmu4YW+zZteU+
/8i7FRRmPDTXEJqHKO9MHflmlrzd9TZVqRwlysfSN9zA0oWiIisL3JGHVhcBUyxP
GCaorq697fByg7YFjQkVm1QuOWD7xzcZeWSZksUSy0svUWHDMA7dxIauia8skJEc
AkRnpfG7c/n3VmWk4RBB5q6BFvEihCP5XcG39a9BQEECDqr4Dith9VSNHgXFtDD8
pNNAJBZrdmykHhD3f55REV5dBeS1o6GJaK34A7KHJ6/j6f3/0zfGatSqrM8dIxhU
GBZ+kXvKKBa6JzduW53fsAv9dufj8k8T2JRuncGnqEIen/EyQLZLWtT2qWLU2Asc
4MaWSRioQzaJTPf3A7N/CSPT5Lw9DDZRdhONGg70s+sgtZcLXen8aVF4W53mAGDn
o1XF7rc9VTWuJF8RbF7/KXcrbgOvN5U6D3o6KoFaFh6LDeXN7XlSyywjjljf8l6K
E/Ag32oSUDMbu0cLf0y5cFhEaSTgUaBU0xdszG4mS30NJfiv0k8jstQGT05gHxJ5
UznyxL1goV0wEX9GAV4KNiySXm4QIfKuCrf0TNuWvAoHWJ8cCjjluZjWe9ISCalC
1oD0LZ5S6kIF1D9fLNyxjMTjo5G2ATMlNBCRQdgKp7tO7EAxDhK0mJJ1K3FE0nK8
Th8JHi77DEZ5DWrL8dJcqnOKrvDHHr8530JG1GGmT5+jdxr1/y86/maP5IYKZ8GU
8QxJ85ShUuJFqViAZDotG5FURS4rstiJDjZyPIOGbY+UkrIXFD9MLQ01wcUj0jgc
+5KH43pau3QF2lK1KLvZ5lSWLss+H/6In/p5n2nweBV6zSvYVBuM/Wva2JaBpFM9
uRyuYUThPUQMi+EWz9hd4ti66QElDtBW4QUSOEwruaFP+BOCa7DUbOMnDIxWpE9z
hasviF+69+LZV4Gg6TXJfq71yRyJ2TDD3/JQphadXreK8X/nGk7baRo1f/JDAaK8
hg8vN/GjdxSQ9JWGfQp/sfaf1OIXFAmDIW0AtTgWOVteGO8maovss9yYKfmin7ca
QtiyYiakwjcLnkhoWAfWatiWHrMKADJfgzdjV71hyf1dGIQK6iL2ldyh1YjjtFoR
wJau7AsCky+uUdXDqd/dUvDS+Tg1Wv8SMSsgK6wwh+a//62HbztVPCBz9C+tfBgI
9JrHJ9B3XBc5u8n1TUelf+N2Fq9V3o7cnwKtI8REK1kHtyAHO1xXuv78L1brKRN3
bOSSpByLAaa7NZ6v564bD7Wk4mDzZJv76+jebgbu7NbRVGG6N0S/TBsRSdkpKVTf
0aXItzN921AODPKtSQ6SHb48KlFOyILrT8RpBjXncsafrzwzbZc6ogF2EARPcIdX
hHzHBqycBBpsGoLnE5U5XATmqjXNjtFtC6/QE3IPgf/B+MYOKZ3ci8MJ300yt+J0
g8Y8fziU0EHTk8a2WZS/NzlFNz2yQwHxXwTBi7mNtUWVLJv9EJbKKPgIgUkcMlLt
R6gcAmhzWNFJJbDkHIzHOtoDSVtdEKStK0zBIn5ENjzkqFvxtzChilKIOUUmtDwM
OavBwDxWFIweB6eecFymTB5u83aFPKdFISMfdMqV1bbPsb5xptWdEn6nOCuI5jGR
KsxDCmRszgQ+/lS8IkBEaBQuHdInalz2M+YQFod7odplm1GYJTnVDhkdOG67TDQI
kEcxcVBNJoyKEzzq9Utq5K6P/vMcc3Wlzoc7Pvjwn0fuCDPfVp/5bzHfFk0an++W
6HvCN3caO+l8p6Sbb4jEkXIDPhEhRlmMwHxMMzmzFMIBpnMAx6GVjrOXlhv7Mwfi
SDfndEdW6fy+wsBMBHFZO4fQju8H4eHjpRKlZiPCEmGyth6K8ZcKvbp4qC/r03Iy
Jy3Ucx/ggErNjAg5Ke1t8+xz3xriTVZsoCfWJKQNmpEbSbcOsGVDDAbU7Yiy5EFt
Z3SYaidw3czmCstq9lzEXzAH9V6DO7G5Yx2NNeZvvReMz2L/uq1mK64df5FNYn8n
02HprAw82ATpGtiURupntI2mm36xVPllmtC9SiydHlzX1xn+cTGuW7eLTEU3K494
H8YncywuhEnG607AaUhgP1vPU+gLYbWhIhOGrP1ayBRE/2+qtG2FraZsDjiEXOBu
wyj8B6miXNbLmYvgS2W88bdFwDvze1x2b4KubMGNuvE3bd99b7lvjT1F3WREbP5G
LkxjWn0us/BqdtT/E7iR8gLzgktZFkjvue4o8mlFHt3MzGVxyqQI9AhFAvogSkxb
vqxqbAfhDpdZFc+ESlTXPCHHRbACmDncTbjf0rv6arf3ovqgmBHBFzBmtFNJkxfY
cNZtcew/c9vhfKN+t5Tpd3XLI/uZJtL4HUtI94C1/ycqtCIZBfO/X1+7PWdROWtg
BU5H8Xe/8dDGPXqOM+XcG28CeKV1zvUM0mwT6tqbW3d4PGpM1aq57m4EHzVlVOvL
UJ5kBgzBgVUjlo0ETkcbc/uCdrUtyzgUATlU7xSPIE3cfm17aOssi9ABdqJAAm/8
bNa+ZBclPNnMhTVHmmS7EH2CgS2YPSOrv+OcnZ7SA9tE7FGUsarYWTEVISSGHpJD
Wt2skWE1b4Pffb01eyjmSjY2nVMqa0dk1sO6bL9kWd2hsrpJYeuFF19x5f561Fr4
SU1f2Sg3RQYILH8mtj7uh/NdU4Zw9KMTbzWoEmzspkBEP4TkxyavvwkL4fa5CLYh
lUuFg+2f3El7mHx3MbnTQvZ8IWNLnbFIhpp2mUlF0XxVJ16Zxka6e6OA3cgzMmhs
0wRspctf4Q8m9HiQAjm1zgK5/laOLapI/4amvH7jzibHnUBwXaZ6k1AebZBkxfVN
ywQqxlzwZg6qdoT54O6UX7H/MPF70SH2nSyByi4fn1ACF7IVxBT87upfq9rqIOmN
lqyd6wZo8RBxqxLQ8KTdUoBralyi1qMfGFrmKugZl9fa9+SEzxOJATy+gfjZqhpI
Mw4w3eLmsG5ayH0IEC2eqBliw6rJ12I8QWnzg77s1dYTl5TYCZ4rBG1ElMn6Vcem
8RbGrnWFZUfsg4Iq+/IxaCEXrGG50BP9TDGbcWpeu+h7G9TERU76dR8e5VYyQI+A
KuW/CV8Gqku9czl7vllqfoeeFGXp2EVtXuE7SkoM2V+nOaySwi75K9nJoLPEOKZz
SRUM2BPCPXArRYARKOswHfGqbEVAGjXeV+fb2o6kGQ+yTmaRUA8FymcWH3a5yK3Q
tb84p7huxWN9YoWulgDuOP732fK+BJdIAYocM7Aqs26r1GqmI4eOf1+Fr8Flx0mS
P/Fa7laciar8p3cysY8+SjcozUXPEQaKdyqLMQG799OZAGHpEZgDybnVePlBIw+D
zfanBND8uY9y16h+PBUbyGwV6Grvp48+zCx59DnAYqxC81jkZ9V05diXGgxxQpDs
MSAHNOwaCaTRdByoZH6hEKXhQ0/CNnZm+CGCOXuUPGMulqWpdZXdsQpOyOgAW3dq
kNwRHx89IuwcWz4TmulxHYYmtes4uMZ5ST+E9X4uAzmR3i8M7sWk8ZeXNFcFUPO/
aV86Bba4x/v7cQsFc4G0aeDt4ez07GozWwVhREy5Ast7jkhoS6t2a/BAbEGRurXE
DsJ2xc41YgIhrMFzjcuvnxMwDGKdt6B9qt0n4/037mhMkmIVUlPb1sXczbqk0FSh
7SVY1BIpQt/vM5vPXL+p3XAUL9XJsTYmPs8RpWy6BrtmlSIrNafKLnxWLzyv3bzg
lrZw683XuItwFUqK94BIqnGmy/zvaxANp+M+XklAO5THrPOxQWETv9wPaO+APx50
vaMSZgXlNR9Xncv2GwNv7IP1kscHPFrH/JbyGkAjNCUFHJqK/uSCp1sXQW8zowno
6MgsoFhgZTGCvMHE3xj10NHHEfJYUCttLacNfZmhRhoVKPivnAmwUEHUN7trooJz
v/Kh0XHFOxnafuh97YpWgz+Ay1k93T4UWvXB9+LwKwkYUtxfBQrfRnm85xPfcuUB
dBMUOblMjNHQeAbWRESunsc7kMTBwCF30/03DaVC28T97PZW/TRQyfmHQf42S5ia
DSd0yPpvN3lOksXnWVN+P9Id/EQMyLMGDor/y9BQwKNl3tycImv1+vxaYmYLz4N5
CMRL3hWJ1Z7yMTjW75ouaEds6rPlBufcVgEy9OZ5EhnIPRNh/9/lFBqQ4qV0sDdU
U0VeSz70/s2hrvJEKqGP7pzFVT6xvXyPodsn1cexlCO0MejXQ+e2RVVEpNWtvFy7
acyPZ+FWe1InxDgeaaw+GGEJIzNBSoUYGIJmKVJuHRocAY56cO//wOzPt51C2EQx
kPzuHhEHW/qSg0iowSR2G3imH2YNg5rZZMVLw2Z+oE8tM7/AFmTGxXtA0fi6bPjR
2HUJ32780Cyq6ZktZUlOOancppBCegL5xoDqwkh6YOwkgbPF+xWlpaABuLm1AUbR
thBFOOVD7vlCE+M8wOsiCbBRKRPhglTA6rZ/DzE4BGv5r2NjkxqrpVF/N49h/qPU
Oj2OtiKnZX7LXgnB094m1k2T8LGu3KhxI4SByPY/Wm+Z/cerm9gPBDVfwfqcN3au
wSP4WAIkUbLSvqoXOlvAvjXTCqvKxfhYbdzOokXMlFoKWejto29L4qbxpPvR8vGz
g4W/UurA6UwVHnF/xFM9FoMJrMrEYipK3819jwPgCHr9/t2wGe/LAhrOL864lBW+
q+EodL234yMhGjBD+zvbojjMEhoEKtf+hKuOLyYaH7uHgT4oaaovtqIEShbFdl44
Jb2FYn4+jkF5N/IUr2aAS0jdl8iXJJ0qrtpuZ5gTVwbQgsc9iYiAuAj26ORh7ZNs
zCCAx3ILuRQtHfj8spSnv/BV24auKFEPASSNByb4H8CLmrsd6eIQoqqVBD151xCg
d7gqzBiTYrj2R1WJyDzAns/hneHu8wNAQDon2SNeDaykHPutmR1ukQXYWWt1NqNA
PEvnNRjhr2UxAyoRlkGQ1/Ea97PhZTmUTeAIj5EqI6pQbbckUlflmRKJJ6k/g5jI
VXJakgv8Bhsj4UIaZH/u932BT6KNwz2w19SM3gW8EVXpi28F/ywOnDcGtj3rpU/Q
H74dN1azF2fnis2akKIKHto7d2h5VS/zes+BRsjU2C86ez102t3+QAC8k/dLu3LQ
MkvTsNPrz6/5O3SNYT2eTArDwhUuOXuktoQxT7whdEnQ1CLpira+WorCH6dCZRAe
qpYxiCiZ3YySgN+cuI5aHOKwFdENSv62J3odEUQ4w2zXnljNe4s9pnl95zN37LT+
3aVkGObUPgOMWiOB5eEIXVS0D19RLovsD7b9NSeg4FKaYeSKJuwyiMcxyfHkxCht
ZwfsgRHZ0AgiLzID2HtQj4XXwWJObB7JpwdjZOZIaPqVpE/youEKowt4rA4fnz3S
Vwm3+fY7r2SZQQQcuN0H4kZt7hhUyChvl+CHcz3voeWXd6fmz1N6MCij5k3lRnf0
aAM/+tOslXHpVfpU62BIUfP1a500ijh2qn0coVKU87DYeLHs7vVVPjXzcEf3aRra
m/BPAHiRlM//KidbXZUfm0LwoLZI5FJ6yxOj39l0tn/X+yQMsZhOGayiRP1hbr8+
vrNSE7a3hOZ2fNxkyxK+z4X9OAesrxi15E84uShf50/3AUmK6ACcHqfuRfa9UYLt
mK65xbv5HQ8UXMJMSsxYF3bc5L07lmW8DN+2WKR+MSRHrWSkcHHu2TuwwS7COlY4
nhZIqsbk7EuxD1nozV1PhUkVrMqvBnaAlTai6mBCHxdeoxcuyR2FQEj++E5YIBLA
k2SIMct8P7Bz6C7l5jOf168NWMvGlQjLVIu7wT8a1NF+B4nXd+eYYfh6AqVGmC28
9uxBkzjD9541wAcq3UIVOmcROETFwnlr2k3dYhJymtn8RytCzKs4u67zYT5JLHyp
0GvZPbG+1UM7ZrixPl/q1LHXjbd36KLpR/iWOiBZd4/s9Hdbnr4BYtfzZeLk5kHY
t8PaqoeQT0ANko7e8ZM8ItjGOgjyaQ9i4+nVV4MicLKS+1ynHDTLISVw0f7ch7D/
aBe3dKhKytTGl25j1N5RPKm6w3jogIU4qAGLQG7IxvIGL0rteajdaGk5R/2nEKwS
MlgwYTMh3t+5JddeDfjS2JStZ0GaXt+CoCCn16zJjQIx9++pY29yejG+wauzNRYK
wl0HJJdFhNwaa+YkIGZuUV5JNss7RTvbHjXNGlsKZjKY727tTUoFqEJWN/+ZS0xK
UZ2IhsrKDhk2q0ZBrPOrLHNiOVPiWs+3O4vaLQDEqpXqsD24xoCpNni3gKgzo10i
iNkDJCPBrSgelebWcorgoHq8bDqN/58nW4LfXL1ouuvGiLfUcTBNZv88+5YSIBmn
soAVDNGUAAgFjZS/FJ/fVkdDvic8IFW+wcy1REx0UOplwzJE2oWgY5W/MTIKHrzN
bZPt/LshFxc0ZrdyYOM+jhWZucqj0sDHmWuyAg3ix5d74RfvRtiGLGZ7A2WV7HdZ
zZhx3LD2VTD5LU2S7EtT2Uss1x3lDFmL7ahiajDaZ26Guo7txgY4XOGisA5BPBT8
GVLbJ77goVi/OGkbH2xdj5JW7ZZ3OHVIy1GxI2ArMpTgFEp2FXMOo0jnHtRZApUO
pbjCRM9Rt1vR5/uVNJ6sLnk9mFCPvbqORV67ASEVYrlsxnwNHekzwBN+j7SI/tpm
euu52wHCC/XsUwnbec6ck6mH8Hg8wIKOIuedM9nw66EB9hITvmQo8kI1fsQRaOEu
7c3fGSWLPz+5UtXLIDIy0ixWnE/YCmnclhgBq7U9oVCVb6+LDzxLq19SaqI7J6AS
e4DwcFhPsCTNUTh1sfK3WPZvajxxS0utu3Me0sZak5srmUIPg8LsiCeZ9ZBXOYRx
YsdYLboYPO5S1bAGOAsF6LfCPTbWjfiQhVcgYbhMwNBNK6xZ3m2oiIXwHduXVhNC
G1vevsac9sWtc5fWrKJM6E97MFYCdSmpwXvc4zZiYL8M6nw+Or3Sf+ltAlMxxn2b
TkXLwDeBxtOor4I6mOhTeU8uo3R3Jds6zPTqwDX7TE6trA2ooNDOFu8JWnmKDoAY
M2k/R1ZeuZBcJSC/rNRHgneTpqmpuzY9oOTw4fC0HWsS8Fd9248hq/JqG7qbpzBd
bfkr5h+uE3VD0BWaP6OqNNm348rCPAgVpFXFGeAY35jEItwVCZ0YYo/d0qjuUmTb
vmPd+HVQDq4pH/cTkdm9tsjo4unMeA4mUgqMKgDqH9oZFsV9ceeIsh2HvnsfezKb
CEmkcHicfMtw0t9lZxyL++TJg8Z0hwfRpuFk92pxkC6iLWNjwZ0u0Am3MMIx73tj
GBfG9r2aGe2t0eRwE/o82KMyZ1B2S/Tw007vEu/Iko/mzNif03L/AFreb++nBjFW
Q7z8X6uI3C9x4us8sCc/7MiSKDo2zq8VwEU/NotcGHHtTKq87CHSmp/e0rc6ZqO5
nlAktDcf6FHmXtK4rnk8YRC3aLFTaPPl1GPauAEqMDAl3JI7RfSFODTuPoacdJ4T
a2RlkyKfxyR1aEhGj6295UQFz8o2B1/3RBJ3VJH/qGO1TT5fXyXJM1smbcapuyl1
Yl1KyNn6PDvdEC6++is12ojYwhcISyi8Wgf6v0MKNaqHHL5cemThIekRwbVVi0Ri
qG/Na84CEImZJRvIBMg6UdM4oWC/zuUVRNIU1dsx+nx+scuYBgkUasE5d+9M/pZW
U5peZbCyFLD7lgRxT+RUPg/2TI8CUCSiQEh/C78NzFVnRRgHDcQeR3/MaZ+WC+u1
+8PevTw4f25FPVNgBfYrKwl+fHLa8cziI8V2lvR7rBSOtI54BvPtrHolqZ2GeZDo
AfKtwNDv67zMs0drvhwGKHGkKQUvxDCdkVRlbMR1y4rCttjDj2udzV3qhMpCmjxf
SHOxwNLfTAClasxc+kxR5hujw84DBntFdbKqucwl+4/tElvrmrvqzttYXKyFBIXq
am5Sou2W3WUyHeuJ4+w8BL+3t5cVhJK2dgDAMbJLHCKWD6+UZfIAiiH4FomTBK7d
O+PFyh0/ulA4NZfqa25bg3glsODnsLvAH0APylMd/hnFKQ4sPA9F/RL86PSMlHC5
pufo8z8eMOUAwkfHiDbS5RnRpOgjzzfpI6SwcL53fobN4u+yOBohlmAXKQBsICyA
nhqCoPwNl7vXEhq06TePtkr4Iun1du6fieRRZvdXNRq/miwsmGlrLBgQo+SyBNLj
3wBYTRPE0NMPyhkISERrT0MOr8HGFI/jxUh8xQIqH4Dggas0Qo6H1kBhoc0UF1kp
Y8PglAtYHCzETEEbohc2nMyoZ9UGc0AvN94hEWciqtEQmIw5aG6GYja7IkBwotLs
uKBmjcjS/Y6xnjouDqt4r+12ssaamrTdSA+IBQFs5Hsi4oKNg1wpz5uEcF1NckHI
Zo7NqpX7agZ5iPZld43MjaqWvzyxRwGIf0UB8oUijlme5wmFZf7QLSeqChnR9RnV
/9pY92XRVujq6DySFF4cQUhLoMBs92USYVwLJ6oU4wUz0EKgunF+cH9IY6PbOxAE
wj/IPa2lt8aDQZiU0gsInjsdn35S4f3sFgeHioVVohjZ0tQQ2fwNuznO/hdb/5hd
2wfuV2t5/A1PNooTQ0IA9jq+PQtN3R160INkUrTrdcjfPlBL5PteYFoqCWPmj0QZ
PZR+gE6M7PsGXEmzK7CcVveh/Pl0PgjNJeF3hJniGOEZKo5MEKVi+jc60ehFZE05
4YMxboAZwHxUra1TyvkagMXv37lNRi1qy73SlHSrQkkMOR20W8EeATITvMv2ZJ7H
2J/vvveYv49PAhu2T0BROuFRCidl/TpadMBIxGYG3qbx9H0/l9YdUFdI6tAWmF52
WXWTT2cS95QmQ7XjQ9vbsmNowS0K3MfB74j5r5gPcnMB6FyRZAx9HrFdgjzBtyDD
rQPCqW+6PQg4mGSKbPwvpUVxuBKacvIrDBvPtTDBiF3qjTiNeQfhnvBJkhYBl5Dx
lHJkfzj1zv1aqzn0H+Eog0r2DnKcJWZzQFsJq8r169Krzcf9zXkqbpnR5qcJJ3OG
PYMSyaCf+WMePc7f2JhSDGvwDlpvXlWVSYSeH5j00ECFqP1+2ygGiqBoG+4nnzSZ
RJ9AWSA/KdAcKlrGlonlS2oN15+zCk+OSNxHNr56lEgvOucl73xHPd6a83pWvn3i
bwesVO7paj9fcSWLnVAHlK8iJ24OJps0Im2KX+nWWeObrf8KIugzw1WmMCH/AXVu
eAUb7PGvAh7WBR/zoNQ7XJJx4KYGU4PayJoIk1vbVt4=
`protect END_PROTECTED
