`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qe5DTYT9IL9U187rZD829JGBd8WgzAXVbtdM5APwTE0yOw+1hH3lY6/KwWyHGQ3r
k3P8138Rf3WBe59sdG2P3yEKJWNjs0kv5a6Hxz5jBYZwhSonuDyU//A5f18HIcQI
89BC6hXhEbkCUrAhJpxMRDcgHLnqWv/gviWnR3iYya8HWiqsyCj4VV8fyCz0XkfG
5UaRyenuWWJVOvy5Ph6CZtzCmAkSf7czvBOhi92AJYv7J7q0jld8CCeVxm5eEuRD
7tqXkQs3eirlUPv74WmxY822rF83xb4NkTuAu8Dcj8vTPmcRlP7vlfR4gYBvhZgV
GZACR8O5U1MfJIamHmgIhx80GyhSPaz1M+79DXIiMFvJrSjA7xEA2GufPq1Uv40H
qhwcVd1tw58gd1g/BjcFnK0gx8PR/ZuFaA3U2F+zuL28IzFSxN1/KPWUD/IgPFhO
rAZuYzox7SvC3Od2fXVdQStWCBRAUfFdhEgYiPfVpB0K0AjpBmcUDXsaNbKg176R
2qr4ewV1KbiPyOaUo3YvuDpx6C+erBMEPysRTql7/TtDkNV9Kdv1NvhrsPVqYmy5
bEYZH0Cmv70WE1ahkA+hQ25c6L9cqP7gM2hJR54cPYkHPdKOn64kgpuoVBBrx3Ii
ENyd1OKWkrRBax6kLUto18LvLAxd7EPPvnmrk8iiLJz+rNfm9PmOaDndC0g0+zp2
0wOgS/bjV+0NXPat2Dg+TwWmz/x0uuWutszLM0XKDnfgnZX/mktkblqFFiUBboWJ
LsbvuSeJBrgvICHmC29oQoR2A6x8XVzWXFi48VBHy4W70dzNKSx5lWsC2ITgnSOe
tdytcN1qybUEqDJdqTsTNQa/yKsxU8ENcc2aWPfeCtRXIA6AAJPcWV0yT4N/pwOD
173c5+u9jW2i+fbGrKpqZS5WPF2mM6eIO5BJm41ojlqj5YosQEMVVsw997mBoEKd
k2ftC24M9Wlxw7pkc8uzCOcSnTYO1b84Ppobp/U1w3HMZI8sXCozrXfH9H1moaMT
hh7HOoiZCl+dUG8RqlILDmoPJWEObAfeNLp0nrIlawGXQrnDKEW8PrGJQiSv1v2R
4BA5h+W0G3CWUJh87Al7JSz5P5cyKimHD4JzAZjjg8629qjBduws9pZ4VMwjO2pG
mWXa0uRGwFnZWuC+1fjaT3rVVL697rfvnzf03nIKBhY3sPJQQKQJIXgDzUiXJwK9
D7HrOJiPMNNETkSh2L0xGFG83SSyg6Se6TyxjEXu9ojd9nrz9ufQb9+Shlk2lqYy
CoLd587dFxv85VRHEv4TMMsF9OehG4iWr15D96FROJOTnnrcp9AMHVFDIuQ5Xykz
hcArNQcOTnFDoJiEdjGf8/fQDDFsvSvTDqZMaR2XPxOiM2mvEsOjKRjDjM8Oty8x
36wkVAfHzRuy4Gbn4KCzeYQvnu+qZhOZOCX5L5cUh4nBXhig/4aBKC0saXViIh/t
El8QaEDB1I9H0EcAOtSusbuvZrHPNNqtBk+bqOatIfk2EVVDP8bNZKgjWABAAhqH
FiW/HlXN10rMh7EEMTZBfcMp59s8fA7A3IYtWGjReLvR0+Eb0SHmOXQEQxx4b1d3
NkFK/ga1fNW1kGROxpH5kJ43Rq9/zlU/tN8tJ53FjKV3767Nl5DP8563rivo8zVp
Wnuvqqe/wUY70aoPFCn36BMoLVCNs73QuI7AetYPSPdoOvwQ9o4vfQ6fTNv3Q+d9
vivRxulmvb4bmZYGXcPkZ4CH8qGwg0KnhYJWFbHNpH1DWL7jGM5CSsfALu1HnU2K
MB1A573hreJLShPUffFLaIbEMTnMgNqx7wb+EbmKZ7WX6BNPOoAoXPEwbjKKgPcT
vzEuuGf26gH7BXEDkC2AOhTo0lqSjYKBX5m9F+1bIfjmQXzZGX8ubBI1CcYbQKKR
O7O5tNRzCMMk6rkobuZ63xOESAE4wTVg7P9RCj6UQ8GRbiQztdS2ujzkvov1eLYa
W59CVuMREUyZE6mHQxh9M30fKq06uKIMBbwRtzQAu1Ncj62QeTk+DcAZNBkJWzNc
TVt4ptVA369aqDKycbWz9v3PGlqQ8etl0bfwMjCAv7BeYDYx63HlfhNZvN49hfZA
8Mq6zHidYg8PmXTit7OQME6aCN2RzNowdn2fOj/qaFff6s0SrCtpnjzelcMaZeXr
Cch1qPy5WJ827OezgpVP/Teaz6UHidOuLEcWvVW/pTchHP3RVnF3mUF/2dZH8AnZ
DyJ7z1EM+zO7/ZeHrQz639ZjI77EbEKKHDo/FULqPUCdretO58NqDqRr9W83zmh2
IdmoNk3bUxSn0FaLszY7vHJivmK+kzRZ2IdU3mXhVLkXycmtlNx+/LPuDUyJTuCN
oEhjiPivjYUWZcsYzCFtj+fWUtd9zvlAm/40aVueTxEV17hMrC2iJvg+EVr+7X00
m75/21CX2bB+F6glu6SHB+9R93bVuKrrGHgptqUUaj53DDGMG2mE6cYkzyKQtdhr
iNiemZfLiHBu/lrcwz7/Si0IKJZdzJuRbhvlo9cbBuvprfuB2t5Nt5Nk7qVqjoTz
HokgEz8+6y2D4vAqepWHDKFIXNxKGcGDm3U5N/T/4ilg3AU8BIlQmrnsqSkBuxkJ
jInyTfu3XREwtO1QQ49lCIlU2i38aXUrXLfHgFpRqB7rUe5ktN3t8bsXJGHFNNRO
MbR7iM8chG12NGSj+JxEZ2H5OhhlKvaTS8x1uisGwnk9mEJbH5V9yiofZgdkRT8K
joaUuROIBNflTcsa7m/3mRNvCuGQ86wB9UNEsUP2pgqymZFIfeHas4wABwd9D060
++wYGJwQhSEI8t5V4fQscqwH/BxLuEleZbEdBtiOtUKWAtX/TrrdtQrFZVqhMzJ0
+9Lw/gFvUaehAGBZdXpYcGGGAXHUKMWEVFlQMzaFycYCbDki+8Sq6bWfe2/YNjMh
HTkKFltSDArQ5zGs5FCpr75AAIlH/+3DZvDJEMzMojuW9AXbFsNb2mAjwLOVLe/M
Izapx7RF/4d8G3zkV84U+WfsYvireeeazr1RCdc00/VF/kDSBxfpfrwbP51Ys335
wWcqNMTMDhJdiZRqnoKM8EE0WqU7l9giv9q4675HbV4jGk/XeaUJNu+IpnCI+KFY
+5UbENhotJPHLPAVOvuvH0pW6KRz9qz5rtaBco+tsmi3SsomUMguLnoYv0mZaMsH
nARYSN18oG2hKtwBLmvY+dAfmnLLnpJRuEwVmxq9G+QidS2X0fOz9ww05AFJowIt
U6jlTByxAs3dOHfw64J/mYGnw3mNEV51h7/m0xMiGLXp8pr6N+IWpvxLRwzEk1j3
E6TcHNJAFVF0Zva9bqT35F4XQSamevJ58RdEHEpeOGNtK84xfhNn6Yb3VJx6hKvr
egM73UHIBGrQEbRNLVDu97UwYbPC11pn9NT8+UBS6RvANdhbuKFmdBwz7YSW8FTR
pP+WEMtz6esqwr5Q0icVjZV5BXYevPwj2j3y00WazGZ0VckCsy619aCaj1xLZnPX
ZnGh0YhhDCKbCHJycBlwbtcjcHYqyrwD/WjXyj1vs7RsdEh8gWeW7EkU2R/Q+wG3
JN51PNgINK9SsELD29q0AH7a0TOM8PP7/1DU7JIvr24/xO+j/KJT0Pj6BT4cklYV
StRn+AN6sMrjyAN2Xu44b1sbtPhPA0vBjfGZCx+1x72lF9qEwEoZxht2ddf4KLz/
bkIQGGCTL/9QL7oIILhKhdTVrOagKcJUuzS7cQxhf9eZG26XdoenM3ZhJ8sDS1g4
uAL467m/lvuFMF7c1c3UNJqK59WwI2gP3TSQduBFLdCq10IymF/DNWLQcpa/MaU+
TBT/StktC5sQXgZiGJnMxsNPxOYz/6fJHhhBJJhUotjoiowhY+509m+79Qy/COdO
GJN1sPcvfQoyFlA7bIzSSNtJCKA8kLgNyFzT/gFBafEt/Sx197brdNe/pc699Ile
OM2RO0I/Vps/9x0AoXLviQixbk3nQvRbpPXX6k0TmlJoCsAchEBKAAQ6/2uEFzZO
jRxzwl2kJYPODCNr5LgmrFZmDD23gxgLqL5fJnvijaqgct6SAWdB6XUwd9bUazOz
rmeD9CVd4WNu3WxvsJYWJQ7H7dNrHQledtZPAgg41/bVNtRx16J/aTCaV91sGEUa
Vx7mZmUimLxQVCdIwjflpnzABWMKwxyTuQJ9yU3imQGnKZVf7Y68m+si1ahvrrn/
bVL1mGrZVyufMQ49XldHcyfodCM4eS11oAAc700RFLEToRdPnmjHVHelNIyDLLnd
6oJfM0/Due0YI0Iu9iW79TRofPnv/tRTWYnLAydDDxpdhTcoqJk/LSLcAjV3dOL0
w7tsE+6/M/C/E2ZsxXJrHZQ7dFCmVIeSCmeRlPHi29E81hCN/onzabh50LS03jsm
xbDygTcXZUW9dc+yw8roSxdjaBj1bCO72cxdTBGL4UuuhM7JJlQLb27iW6+Wc7Gv
BuiwPWAB7iwRh7iHk3B/cltnDUHM9Ksd1pTdWstY2OWSu9hQVdErfJrkRtKBvodS
C9uG7rXVNZEG1OzAZjVrbErVl4Lp0wOdEbd7Gz+icr0X0X1DxYH5chA8iGfi3g3r
VfYzVXN6OQsa404TDBvAxfgONBUZ2nBmc0Y4QTX+5WD1Ina5dqV63nSsxayM4oxh
6AzrVlm1nfUYmMaIfVutDsVGUvlrHM8hBYTZxm2kjI4o06AfKeu1AsKq2PFlyZiW
kocglJffBcxIWL0B0DqCJyu3OLVmIxvaIiA6Kv44ZpU=
`protect END_PROTECTED
