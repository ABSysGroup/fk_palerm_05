`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MoN1iO2aDVzvrgta6tDQVLYv/xiB0LOXPwD8v/TIQEKHl2EOFNd5DADCof/L4bYx
EMbl+LtNIYKORECfHVDnYCZsnkJfnCMvzQd2HXLl6u2F/mf2ceC1gQpJcU2A4Kl9
2fBJhVb+IWYHdt8Mv98GQGepoP/J294mA2nCv95sD6ToC+Cd7bDnTnTBnCsFmAGN
T/gXr6IE3VRWR9HKZSvl5JgajZmSfUcf7TCfVWuoJ1to9hgQ/mbLzRsc7ifQUTex
n9R9E0rTvHUGaDdRfiKHJ6lhNppWZmexjqeSG2c4fUGUma+kxgRiKz9OPQWdEra9
MJT5JzSK3h+SjVLK0PEWdlfQDuvGhnv0Ga3QecJFsy3g/lWtzqahQ3ZM1F9p6RAk
09QBmOfi5LkccNIEP6L3Y99J58yy4HEao6fYxG3hSdoMq4OF4c9cMoOtBgCTQZbO
BggzaFqxwzQVsVZl9B0levv5ad1CvaZzmtksPA1SbG6eY36oNjOkuKESJ+Q4GhNp
Hn+WdRfmvUZmQ9yK7in5jJOOBshEJZzlqgRabmXdCW7CCTNrIUyOJmrv1a9i+Wb4
Jc3g8rxPZ49OimMY3ONyU4IvFpX5e9F8QiedkHhKv5vZMyvP9evhgecVfoTKl2p7
8jimtTXyvlYO5KuTb7nbbkh8H++pvlN9hgq505QG2ikimjd8J+VCi5a1wVTC3/Ls
8T7Z5trS/IyV/gMT+vXn5gcK9LEyEbPc8wxCaQatxShgZYU8VCu41MMJe8IyPytd
oUeGU6r157WELK4q541qm4riAgsx64cZpQzsyRAti1CpCnrehw1WExsXDfaVwOtI
tgkKq4IS/F9gHfqZ67OeGgaGLZFfKDEcur09A/ntI/gOFBfnhGbl2J/GhR/e4LWu
v6i2cqaNbSD+Zo1D0hUrsF/diFbSc7LQhBbeKCnOgwSJNMyXhm14pcpVjc8GmgPy
9EFrpxnq/50e/RHwdHKh1WKQgpiQa8v+mbpWNL0Kia1hkRXKJqlRNNriQldmVUki
semUODxy2gEmz68fIqyIdBqL2gIEEy9Md/3QRDflN9puvdpWsU7bunJwk6KgVLMa
2FQf+ju5Yinsss4D7q8azln++QU7j0ckkCMK2vVIJVj/L3+ZlYp1CrhP+e+t1osP
FKtctGigbJjAc88pMIeq5g/7YaGTPPp84R2TCj5V2lhMGw8bR4wcLV2G6HLxMJni
lZiP2gzK5dntDPtyaZpoGCc9KrQnSnHRoHrr2JnCJ1sBHETTlmR1FCma8WmYWvfi
dTa2NocPaOnkRobbdee6k/VIkHH1ikBhBanMQ3E+5bS4YPnUsSYBwqtJ94iNlTHQ
dFxKMyV3Bn0PRpwb+wDKa8SsoqhXvar/VggewbICJPBFHmlRMfc3kVs5oQE5LeQO
fYic5m29HPARZVhp7jNfMtrU9Zja7lCNLTT205XK7R1ng9qKCxTqfQxvfqtowloh
UFAY+qEIxhZW550nJJHxmGYybBcdcZyRYQgQKsIThuqL6Fir5jwm5GluMRs+xhch
6TvPUNfFUmLTcLOOFITLby9t92fXbBUiO2nE87fX6YrgdAX5/PZCQmgxYdZd4rIX
IE29mvQvkfnhwKn95g4/N8119G9N+C5k5LekoKSGh2XewB8DFKJkWiKehy2r1VcP
DkR0qv2QtQ9egyFxWkx28XTlAv/+rkv4DBeyG7DXX/UaweHng/JstZqaUY1qTpaW
zIj/5ETZVB6f76ZuI1SuwvoEc0G4/fFMgSj2dxAFTSU3sdJ2zJm72dNhUhKcl29h
rWMkxg/uv3XkEkfszSaSiyonN1CM7GBVGjjSY2NsaroaNzOUJKrsPlCsbpGusEuK
EFCcRW0Fb85/wqrHt/mvkdJ9lYRWsfYGBXEYGtyGq6E8mXaZFRqmN4xAsvbjJSOZ
AQ+WFkwqnvAVYeFcWZmHXoY/VO8jW0+bgkqWNe87oO2QzKkE2WYiRSUu+5qbW3C1
59oUNbnM1PH7XrXJ/5UOOg18B2Ojfvo4XM5LSaZ4zwmtqQ6CuGaRLRRl9mBtAsZZ
7/8LdwUYgHITOLQjbQ8AFRJg4oicamck60e/9s9IP5Y6f5+a/4XfiUcUmDtwocp3
UEn5YGXf2Wkuw83p8dDy7YNOag9fFhNMoUyVZa43BerNDUg3tLYZDa6Ww/IU0bFA
1rruDOtj+ZLLTbSBbE+cxM1lVPfqGxP2vQgv+ZIs4nTKr3zH4nHaq9aCuMdF99fl
loA5Ge39P/RfHdMx7mkkgPHNE4K3XTqLXU0XAYbX5Gg3KDvF2/Ct7SeMulfAMSA2
`protect END_PROTECTED
