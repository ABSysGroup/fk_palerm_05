`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AxaZsbA2bgewGtKi8cm1JMRuYs54bgbNmVN8uLruNGkH88EA6IjFT7cVdUQP1l0P
E3wnuvop7xXNCPHF4vC62dc23IeOTTGbdghJotK/DifWZtqdhoN8igNF2Ic6DQ/V
3mhzBTCBvMgCKfTbnzPNpmFvsp+m7gLs+sQKWaxJoVVrfeSUt5uVpdiuAxqXEvJT
Za4Nn8fFjiIbt8BpizSqFvg6Gam1XNrWefwRNJ3aoenfQg1gDtBO+v0Xv8APoxMr
LJ0PHVQraRPJ38Yvm3GZ1muCeGx0sVsnKCJCaDSgvXewvNpENnAj7LLNkjlN5c3n
t1tAx6xpwqTwI2dC7kJmLhpPfDZJQ6OF1Ltpj19LUIAGhvBCw4jGdg5a5nEqKsEN
kYt9k3noaHXMO6Zj7qgc6IEGZo5y+waf7JliqTWLHvdcJMihYiH/qThZlJq8CDXj
aENzUbo1BMQ9Sf9WqUgU2mXRgUNxNx4nbJiPLCZogAUSHC7ZgS7IyPnsr4SjflMt
1QP3v74VvDaJpltxtgngcWfwt5tGTAmgrk2AxGd0VQJ+PhB5Lx1annm4uetDbjiS
DNivZ5SdAa23K26QLOHruS/L+x4D6AOSK4htRa0LfnkWRqWrK4Ex1anEYahEhFYX
ZbTAAWlmz6CCsMJyoytExoljlJY678XnFQhFBQeSdB5sYz1aeiNEsvNoffvcaD4R
/CG+sylz4nSZm2a0qZqNx+kHXfXU7sZnVtkRBcnm7WIh2rg1vElNPWhpAAHrjpY0
wlZh0+LS6Ti1ymHvnCrXnm22dkTdL0StuUUpSTNmq8XN2smg9+8sa6VkipsVjb1p
B5QnB+Ca++aW4WkHOKXG92ymss+ghUE8G3f9rN0CFJfGRGy05xyNT9wHbhETTDaq
ZAnnNcve4zZVqvIV2n2P6RVFW4myd8fqpvl1HWvlLWJYZ6iH/MagruOnFWW4DSY3
vWvo21J6ZYEAHk6yTLz4RGURjuLj4lYryChsVi54rhFs6mH3eWnyXAdNsuzE2vF5
lHqptCt5Y4qtO1lg3qAyVnpcqeMBLgN4iul79ipwZmmXbnuJBreSxSxP+9MnhMNE
9tElC8LxnILEb73uC2zKp6hGSMHWkhOd6YQjgzW1HN/8erwnU4eauj4QbYPhmqHG
bmfW2LCCexkg0YUM17wJO0v5aRL7uo3xGVTlnDpupAyN6NpXu1kBzltm1kQykMgA
0aE+w67nyhouDnpUi6sKTTMfBfRybqreJJ8slib/ibQejvV4lEidGj1+8RLQjuDS
ObQ4sGsMUZ4pnODiFDSwSrek+BJnxtaG7fLviLKNMo3De+BwiC0D2NPFJ9VBjyGk
B0uaph91KkPaztyZ/SuQNmvZi6SSnoKE5JZbA5Gdawih8k8jMmi3SIFNGCTEVx08
ZVlS3UOYK1FWvdYB5mdxVFNpuHu3wEnWaQ/xCo3BO4yfJzCHkNYUY45a1xK+Z5rI
lx84+Ds0qhqPHsScATqm0DKH0JaxXdLwVwooMwzHWXQPLgYWY8z0snRvo2qHdaQP
VULxSg5B55SZtOMFS4Fu/E72FXOwB05Wx4FzfnDk1gj09kF5GAbaqRwMnihnYZ02
HzJynGvdV9eJDgpbc8vbjUjjQt3pAtaVFLgQ74iqsTUkwGLsjr7a7Po5PzpOg5L0
OFs1mXtalyaaBLX/LpXfEOu8NFOC3vLZW7XCmjUZaeFnloaxNRbX7eG8CyCmuyCn
TtlcFdhruCccDaXILZwA9cBK02/8iatgtESgVar7Y0JOe9rP5p+6Ar5n+Dq6ABBc
DPh9XDpAlWD9aqy2yh8XA4WdekGyB2NEk+MyvCJySKXnGw590lKT91rzW3xsxgqq
CB5le0NvjxX/gAfQpuJCFXy+TNCu9IQe48olSRmxga0X3+MTpFdSQJ/ERRbnc0WI
n++/scV1k2Qx5kfF8xj15rbVt4sKUFc5OUHrw1Qd1il0OgiFEd4piqqDXIlG8wKQ
SrWihZakZvwEzH1DoEX/bXGteOApg0wc0kdbtf3HKO8HBKAsb+I22wv5KSlTTgbN
KTEGzRTSLmBNz+nq2VPlhUgzsDcg1s6IztJpGnh4UAC3+wyGqgMhBDaNNAZa5iel
KWSCNhqXEgUnE219dMh9w3+2YJLXoNj8s0byntJYDT9UPbuu/zDELiKp7xQX8Yy7
sQHUvCQEDGhyIvJamQpMGMIs4l5DFOOsRZon5hJzlBl5KeF5h9OWGnKRIPLDiUGL
4UKYH51yL7F5EB31mUUcE9ZTgUn4HomgpGqlrjPD2hjF8DEBOPIOmLvV2AdHFrVz
kHFoOO25iUeMeIiQX7DUC7yZ+h5LkuHucEX+r1cfRJxIfX5BO3sgP+i/adXycYZ2
cEpFwzQdITEfc5AbiJzNd5W94tI05pq59TzWGSm8bC5cnyJtX0Adwp8uE1Vjauyy
UnXpfpYk+ewYU1kPbbADm/JrgdEzV+OOLjfDTkbeYBb4zOcMPODnW8ucSc5c2NIs
qRkJYupbxOwB9goApRgVxxszmJqAhE2IshiQpJOWYjQa/udChavvLYi3KtyXANjv
GomWpEkNn6JStu6GiG8WliwlEVlfmaPfIBAom8zfBk0Pk7GzWoc9mPwJ0gCWBSLV
K0i10nNFuhatLCRqhogjmFUlM3S+ZC2+SUnX/Efl6+/ibuG6fxs5f/EaDKtbVmZJ
zOVQEqKVKc4y5bKbfxrBlmPt+3M7H4Vemg0/FnfxBV5jYJC3G/yRpdFmRuZ3wXUF
JW0XdVVCI3JSVdLYI1O/Q1lryiK4GXzvv/nakUT00yTeH50L07nCU6Yw2Kh+TapB
G7ITz2H46PHhs+urkAMgVeZET/JpQP6BPe31c5aYACCAi3X2vp4T02Fc/drg5kuB
ieZuC0ogwhFkuEbDr9xoOu6BEaAMnsUG/gnf8b0rH3Tpl1UampQtXCEjbm9bNRtO
2EeV98x7r7bJat+9Z6nmJvakfwY3aaZehrxqg8XgbfchSenY0q9R4jKv+9fsYEv/
sANRCcXJZ5Sda1m0S3m/Uemz/I+g7jwQbSO2ePHvJIA4n3labccFCtOaQOY5Vuey
AKGIGWy9HK4bGzLRW85v/ECkcitzbgBXS+pHhmDyrK7EMO+thjN/OOTcn9IFkPGo
/ZhqP/FabxHQzFHs3nmKyK8V6Hjsqku74q/U0D5CNJTCGS0PpOn3hdSnm8R88YoD
v9Jv7XkO0cit11WxTB9KdVg1sZcH9tJbEmjo+6P7CY3lmDvU4/V1FkGY8TLZu9+o
xGDdv8p2gqo6M44OVLVXxxTLioiqnlkrIIeEhjCRcrbwukX8bcRSZskPXoP0lRb8
6QEk+mcO5xuVg2+1mYYjuu7CvhJwv64fLTVJLHjnjwU=
`protect END_PROTECTED
