`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lesh6Kl9LKFBjvbqreYsoA5pogjH7zJaNCATwDryvj4f34YNCbP8j7MPojpyBTdt
/c0uyfZkMI73eom++rXdXys9F5Koz/8Cde/T+fGKDD9YBHfM49jZQJpsol51Fw9Q
td5YcV0kp/k5cwpqPkAqn7rYrQV7WrFbWvzfmKt+fol0adPmSWexFFnijycYf3l7
CYKtT3I7BjcSEMV8ItH7q/eF1vKq1Gzu805N9qNxgQzzrjPAUse5+cU6a+qOG455
BFVAnCjcZqPedkR2hIz7OWsG5ReHn+2eUyn3JJlhgspvXe4o3/VGOacrl6vCB6G0
QTMUrwPu0Wnm9U8/tE3zNH2JqEWFgkcTDR+JyV+dLE4btqiO0Wd/Rj8TZjasrZPr
VZ3gbHGdVIazHVMLpDs70erh8DziDDogELE3oer80nlj6ztVb9FHmZfu37plEJlm
+4aOoxw4zdcHzLW1f5/DzqYyNoW5n/3+hYKibjF7kDneKWreFatOWvtl4fO58YYW
FZHf/K/jZRY3L772BQEuzB3L0WUGx8dCkrzGCQ0+7wpHWBXRvlRFUU/XpfIcQo9q
1LXNqbZZFebVMn/p5hUk2vFU6nbA5DxA/xX3NKGFNfZDbGu7VeuhWWaZxGLS+jYK
HT4nerOWuysRCYlNp7XxgAoCRAvxIPc8SpvXGZQOwC830EwaEELia38dexNNdXu6
mnLG/Zz37PAjdbhgdu1Uy/34gI7Q6zgmYmAp9BCHMhWv2x0KhaKBKtqHZ2sT/31P
MPTnIMD4H+tJOg3Z5ni00kSip+fy9hM9jfJ2oOe0S+T+oi474PoGCMQ70jrjRO4E
NanRWkGSIa0wGjuYAlZED8IaF+mmQXVTOgU1FH72pRD598rPP+uDKP0tVx7NX4p5
R+aM4qcPXJzRDV4EMXDKMEWQyy91Bk1zeqsAZ34BiG7xRqnyqrpkaP3Xh/gVuiqq
GV7GpJyDPDagdeH3TOZ0hkkcgAbJHS1ZWRK/v5bi3Qb79MeiiLGtW8uijVUkrvpd
Lxb5KqHMtLNaVbpF1DDCKGfjvYJuTlWpk+14gpPp92I/McJY7kgqb5LLeAystBv3
xUFJbXR72PbMmYWl896A1ANiyD73YzMgOHZaxxVJLJlhoWW7gmuR2BiISMH8tv0n
JcWKaGt/2CZ4zhNvlERjcX0eE71bEqpTFKAWl6zinTO1+E0gRLwPh2/Zr+oP1Nqw
qaKAuydVB9/vyYW6hXbX19ADBgXFXeDBafjDlltguSqYQkIWntDAz5p03PIIi2sp
pSTblF6eJrtsXKX2J0uD7PoQbGAl7CDrWgVvjT23cFC9AwhjGd91xaEor9EN6142
UMzuL7Io+DaLMlZo/VVaE3Kv9wzehERztnsJfJUpt1gM3aay3Mv9q4wPn7FfN5af
ASCz4/0Qw4hW1D2KX00oHiNmwmvVHinlwfpen/bYZNDBmMX7g5T0UnuUUVHn5U/i
lE5ooa/N+n89H5emtTy72Lzplw2xt9h9gDTAI7CORsRqRUVDASBVSr+xX6Y1baBB
eRNy295HFu1IIbD68HbZb3JQpIda7E6GgFlrbJnyvPbT7pFbIFypCSv2m/QkhNSY
qstT8hXFxM0j7TBMnD3MjNYjSRTK4JIKcuV/z2+ehvEWL8E1ss0m265V2ZczdjjN
V9nXGx2xVymnYKBYAhw81RP06T/2Vs0InP7OS2pItH4/DlE233ud75xLgRmuDnz5
5KYS+7mzzLtYWToVR54SUtum70NhyM8nYMPA8df6eE+/Dra8vfmmGbKAqSgNrU0Q
pQVDdJHka4fmB58CarROqyB8zIovzLOgHlLsQNDfjR/Hn+YrM9LPMnzCpA7cHv/d
OFEIn8ap/pAYx8nwAPLlXNd01HX1OlAOOCMXSH1g6fejMatbwzUdbwwbRmH9aiNZ
7LCjTxAt3ZU1T9+9VrdANIdMWHlei8D4lqMb/toGuON5frEBLmAWIuEea+3gXjhF
mD3FbJ8wZa2feWV3oLA4Q3h87G/Xhiy5S4uEpEtFNYGm/KePbFKfv0rQEwH+O6XB
SYR7i//PWIJIz9HggFE4PIOov7i3055qsHhHkDwb5P4/FYbqw0kFbQekqqHVxRHR
kipuRc1s274+dNhDGrxjEHt4dbGqvZc+eaAtreduzDjqxX/j0DqO5e4/aKPHqJkD
c66z8C02ozsr31ilL91JhrtSr3fyavGih7PuRFUfzbpIufv4fMOP2TZVSP5s+zcU
BN+7BMZ9W+hbfAXuySHwX8+pl+CqEbSZMm5sWd1TWOs/cHo+Z4/CdVJGcL6G7PYt
5s5E16wAr3VoFA1uJJnnwJ3g0Og+j0j6Ml56qr+KCaQmbIL3Ky/TFSTN5R4ay10I
2eH5bFDZTbp5KAelJv2NEiSS+MMVyTEWwryEkbEKINzOVwPnC1ACKaIUTCsUZ6ji
KdjBXAOvyPO8zpoxcpeKgyjtOaQBekCy7e9BFtSVGZe94TyUUXNEoceQ/CMi+9Cy
reH/o7U1e2w7D+tLBPd5nLRElETn9UNAfJscrHb9kLxakmpOIlk5ZjqwAEELJMIS
K6EbopDa0wbbREdNgYgMr1miDlmqsmUIz4s1966UPY5b+POw+bE4eQ9Y514WVQxX
JQ4HO0HEb6PauvGr9n0rPmWpfdWK+6g1gK5ciE0jO6m30wonRuHB3/aCrS5Mmoz0
QETNrn2DlUXPGxig5YtdbGzzGceS7Hd8Tyi8v2y83rdLohwkPhBGDQJoD7Be2se5
cyLEjvNhvTDqRuDGbguwF4wEacIuwR8Lry/aYCVHtXoThjxKLOx4mQfieWnjDzpp
cPGTv4Sw891jMGz3/m/PqD5q/zLfEndZ7Ctdn16hv8Va23TN/1c7SsXXEZ/CLQ1x
g6Z27Q4sk80mDsfij9SHBFUofNTivTS91OtpmfL2yf+hwa/VzJWSUj1eiQzkSV4x
WYdXtETSoeSGJpRxuJuDQJKeZD00lqomgPqXPaLZSvE=
`protect END_PROTECTED
