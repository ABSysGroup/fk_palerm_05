`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VBDb7ScsTAkvBj6BTXcs3PhYAX6BF90gB+S4MkEOHx0mZszckHzJeSovpM3mj3jU
cA7tVJxIujmKyfbB+23x1XZLXUYJ7XMIhVEDY41fmBeme6UykB8ehNZbEAfGdCNu
ZJUu0VXam1BSyh2Sz7SxRglJ+WF7QZR9DkLI7HEFqLVzPgPaC9sNkCwlMI2UgdZb
yyMn9to65s2fisgPyd3+lOYaFsSSrf15GnzHnyYdyHBmcYy4OHYlXAmWtwJpxCqr
iefppCawLW6k2fBKKAm2fvvI9pM/fPoXxkxghaGrVS3NqWElwXKNig865rrK7nhj
ulj/aO5xxjpvQKtp53mUqyvdLFbSN/3QjQ0VAF+OagXP56z90EpAhpjrAxjh0H8z
G/aGMVzUmMxPih0IdhQvh783A1sz5u8McF7Yosjvq0v8RSW7OwNjVN2LJN2H5GOl
`protect END_PROTECTED
