`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p1BIDyNGsbKkGUdJ8VgiJDQjjVRuZnc2uiHyp5HC9cmgylqaCP/Quz4p7LAEBOgk
c8B8krnLVh8RUOLzvO6WK6tGg6EHSzVWhYjkK2QicBhMhgF8aWYkc99VA827LqwY
wzSScJ3b7PM/uXAFqdfLg3DwffjaTdBYcTUZZm/sl0Ai5rr53dteEwCwVWybITY8
FKm6ezn3iYmAQTDu3ndfCpoy1EBpo8l1LkASKArYGZghYNaKypZG9Y2fOdcrJbg8
18teVLm8Hwh82sW2WljHJqAe/YouzWsN+z5ZuMCglAiJ93Nv2ztVgfASD5XmKU6Z
JAYSYyAHPtXGeDxcqU4hcauKK5JZIaAMtgDFKKuOgUmkSyDCd1AYEsNf+MZTRat2
Aevq1oOPGDlA7jR5/1ztChsNJpkaI79oOYAMlCNt3BRt2EQ1nVByOqLVLprr20sV
m5Ks5ekklszwMc0bIiqD9w20b1+Bqkluibqy5tun71q/p08/ZGW1G+KOVJdRjSxz
crjuMmkYKcGgYjt0vqd9BxDvgGcwMn0RgVzNrp1Bh3GPWChzS21tjil1MYf09DwU
E1tZqzWHvjJvMGnMvEEtkTvdahlkKGXhdMhmDGkEwElN0EjAx9sC5jk70uuW2lgJ
fEyhJGTwNZGbfYSnzQj8RH4z/y/KkLdMVdnckxIfSNtx9VdsQs5bVnvpmUlpxIZ7
A3urf7P7ra+x7/qOxZ2anS5JdgA/nJxjZhpp5R+hKIlr/z5m6BpApR2yoi0eczWW
laYnHsUTBCr8j23i3oR0pdkcWcw1tOByqJHahBzhoIzuRBvy9fXEBDpl6uj8QfKA
SJeM9vqV69/qnOy7+4j/9u/iNldXS1BVuxH3yfyfww9VmmCN22ZP4C6sHVUTdz8c
yqS7iEIr60XLK2q8qqi6450+Ftaz+0J4j4FQ8KJEVq4jG2C/eM03DX0b7UIsjPVq
ZnUVzmJyywzv3f2fLQ8VPL6IbixxR7OOAAzSA6PRvZdvhwnc2Ym/4b+BRkw63TgO
SMDxE4zP+6JbKEuULSiNiG04F4udKgASZPpb5tC+wlLBn3acknU2wtP5ouWq/4kV
IPwtc8ZlrJY4MbFHsXed0C1NygqJg/NvUF9g/RXVvUGkxbKqbjM56oJGdnn82Dfk
yaqbOFR9s1v7gcZBEdfppkAouK1Fh4v+2STXSF2cIaz/OViwcDnc2lwH25LPIpWL
2MKOTWjS8zbprPD5bK1K90H489fz/ionP6yYGFzLFZqKcB9wYDQmDcG+I8jpbBzQ
ph3BZ69hl8I5p2FM1Bbj4mTH3/G/tzGJm/9ok0HT9BnEtGABNcG5q4XBusY5zeIK
C1DmHTzgq+eCqd882lunby9YiWEMQu9tNulo3h1k/Lxk8w0RFEdwkwDcwb1eXChz
5hqQb7ycF1zuD+BehBoAjkXkM9vus47pCELhIFzzvnuul05YvkIS0UW2Zdhmx0ek
Fao2YQDYnmcjkUP/t+x4ZB08hVM2NKiRRhbKOc+jHpQeiblPWMJltduTFx5ULGqm
U7OZlK3oYsTryqtxoRzPWlWXEiFiIftqCMHLSddJMPYNtLnhLYMni+73gu6HihSB
8/413T+lZHCDZv2G7XTehRYkKVdN4wzyivvYpTNAXmHWKCn2sXsVnvBZ8jm54dUv
Ca1rdRmSA0DSjcBwSFz+mg==
`protect END_PROTECTED
