`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KH+N9Aw88XxsQnvXpek1DQBAhKXRGi43uCPPnL4L/HqeSdBrti1rM/KHKpMmn7YK
+SJUM+CZpvUPsQRdsrPHVMr6joWiXh7lfMVQLRJCr4l4u7gaD9nUthU4O/7xYiQp
k1cJHuDLDs2t5QeoLHaNZfebYhY413elVwkg6SBxuRoqUFRdJ0P6igi2T+m0qMma
xUbpCKhZ/IM9sUI98FeYWxdBfxz9ioW9w2gzC7Yovck2qUPZuK3ENKVraNeot/fK
uqfxijBz6N1KWXTSUKCwMGKlcnm3qcHZ3VOgh3Xc5TqX0lYTUVHGzvCfh3U3rWhI
t601TG1ERpyDuZGPSOFIH03XZYBPrflQzJIZjZRSKJjUJcwddshBmUIreEZPJXOB
kWlIpFBrnoNskKG44kBUg748Bnud+OF3jV2Be7aDZjdi0G67IpcScL627SLyYj3K
svQDBXzQweyBKwk/aeXcQnufL/WuPP+OyzdeoEu9BlSNrQMZEWkPhnbQNEA7A4Hh
DIkdnkUxtdTG5R8yycrg5utTMSzmR4SFztchSMJABhSTq5yyfAD5YG+PWBKPrU16
`protect END_PROTECTED
