`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7aI+WtfjuyhceuAhX5ROutstw0StewqNZJwExoObxO/7nkHwOMUq01B1gPOS8bxT
vbHVzEBjLOvec9lOILRA8UAO0V2NaWGm1HJEORvCkF3LZiTuLGhHIsln/cICi0/I
CLXC8gnxGNXvZ8blynk7rBKCI7X9AECKoeXyUhZFBdisGFDd9e9CfVK5MZXxJZxU
RZMPjbJwtiM7tFQNxQ8YHKcLJrRj6mYwhnkl4CfPN2xrsIozHHxLSZnOduHSHAnq
ibNzyoyBLSnqFjE0Eszy8chnQ5Ot0CQ0nnNA9idppbvXSslwcvcechJwYmCS0jGg
YlCPZRE8cEP4qkS+FdkBm2eg1u/jjEgCrZsPWr07+GdZzsIUw/9nrdc8QBAK9rr0
vamfRQPWF6iIAV2aUmaG4BmWkVAAGWZxYmm/nBj0bL9IVr10qMP7icKi2PL746xT
9LpIojc2PE6iyOgkW8+OiHMnBu/Tymcj3bCG7Jzr3FmO+hgxlMVAo9FL2TWqrw9e
6zwlWMDK7WkQySfvXlZrH/35tTABSzc6DQr7BlEbguMNTyBDL4rI7+Nn4s5u0FQL
n2Fl7W9Gi7WBMnzpRkLPhS8gfZlJikXyw6A4du+37/5kvSweJicOXrQ/tlYHRraW
6IyZVHVQOh7cEnzH8VtGom25KBYoI5Ut4MYOD+cvt+YUUGuJlW36SB1g0jctizDZ
W8gBbQx/xHHv9BEXJ7VE/hOvBgRjxL+7CdLQLjVRP5WZGDG169DuwnINVD1TG2FH
K7a/leuINKLWtPvpkthTLjNuA+cb1R8bn9bHAJAWCl5VnR7Z7wSSfwQBkCburTR+
nD8SLS0a7iZGOpUR1GHtFY0MMem3l/+uiCvd5ECM0I2IuPkPrkbF7ZouVCoWlbJp
Ug8M4/j/CogKLjpX11d71BzDZVAw+X2LGizI6wRJovctk6rpz0DsCK6BMPcphvns
cqkgvvdTzYmz8V6P7b/QT1nfwSBUWSPjcg7pI02fnLXeFbDb0Ixy292nksp21/I0
qXPdMxxVaFsW/0LUDuMcsCZDyr3n5v63ddkJ0WsEIX9UzAvgVJLa1JkzFRQ/o+ak
wsR65LEqB7b022yxEhmZQcrVWpmsoGLi44B/+1wn6B9WsN8QBp60Ze/7SP2ns1Tz
cWzKs6bqZUGZ5dU4tKFu3PRib/3Bxo3uLxkL4UtWZoN9HpqIBI0H3R7xohmCjo9n
gnj1i4hOjvwjFRRV8ZMblYGgAGSGIJXIVi814MNPLgTTn9APd/Ce5m89pO3VRwlV
gXvP8C4Uqd4MdMmccX55Z4fp/M+LE/hUM7PfxgFfkQRQJLb15/FPXbY7vQPGXspP
p+ghwTF3Ch/yy5dCDGIn0qzk0hjYFI2F9bfT+H6covl8tvsFRc1fk3GZTBE/6qyY
eEv1JNp9Ba4T6Jt3Wlsxvh+sD6NItuJBtEOrkZ4QQlyjz2v5oSyQyh1vN5rwFa2+
XOmP46zhIxrYguoS+XHUa+MRPUvL93Ni7zt/+CGTe1VMqfqPI32J4KHfW9rvq1IX
b0CjV6O8fNdnfaHb35/lsiC9cGGGMH4/zhET5nPZERda2EUbMs9+HcxRfl9UKN92
OTTrbWfSk3igyPNUBM7loUZ8Nw1lMZNDAaF1JglsmK/nFtBo9CH86EpGB3bYrOkg
OV1/ClTm/XL9O1u/YvbLUN0BUYGsS94ocuFxtf/6EaRdbA5TR2LIq1xP3o1TKElK
jK4kBoo3YIZujX/KM/kr8XiDClonN7sdq9eVBC6mr6F+lp3oWsRDVGLHvT9DrEES
YNGRQJgknxhdtOIIEqVhCFee2dQ2P4e5yQQryOedJ9x9MOOjNOiUGN7UUC9ROK7U
8oFAXKzaGACyPBlm8ncodQPQyaT5KxNWhU+XWKLYthGpOeiNhWwL8U8+PXKZffWR
0IeWuNi1V+v4aEkpXET5zWrU9cs/A3WIxR4vX083YkjDdBQpt+qSvXT3f/XiMzMk
ojcYGXxF+1pZhNpCx6L3nr2gAY+XVPTuuzx1DH8xpEyUHDxq0lWh3IApygo0+2iG
WmLWtuuD7GoezQ2qlPUgpc8KeoHyynQ0oglUEID/FDKdF+Gb1NntcvqrcuxQUh6X
kQb7L+Y8DakwDo87nPgckaanaDPp01lTBQLJr2u5BzIVoZqoBERJ/sgaFgqf1uuq
gFQ14iRtnHD36ZZ0EqI66DJrh3uPI8TBv+ggoGse32/pgJwZiYo6JbtSbdvvMpjk
raiGU0jD3AdO1Y3x/pKXJZ/LBr7zsYnUFumghku2LEBgvNDmINMhMvEDaF0cPfhZ
2Q77V9ZwmKh+fhg8l7EZGlf+oGSRJrzywIwKbuPV4SEJYVJDi8u2v6JHEa3sI6Tk
oL16KVsTDSX9H7CCODLqhQ3HfHi/7TksZgbjQin/AuoSJz+90FtuwuHugEdY4XNh
wstOV3528LKsUhszZPbEZNuo/vFt5+QnEdgtBz2MiZtixS/YITT3AUpdmbba68Ne
L1LmWWhfr+P54q9bBk3CHnah/lGbdig/KCrq8mhWeuAO6gD3zgn2iq0dO26a44h5
PwO4W4eDW7a6oi07vOumB4SzGFb4Sxwvx4zZre65Dk2O7rFbEVuYVCPC7951Vskg
L0cMM87y09eM+Tcu4R9muWQsSW6nNCaTQuhxjNuOQ7S1htgmY4fmPXguKrnRqhhW
GgxSMoyWNvsPZaI9nLIfoMOiU6641w6LQkxkkX4OQ+Sh2w8KndR2jC7g1u1WwaQt
QVuTgMxU9Lr6AWziCnKrygCtqEkVfv2rzoczFJjqFGMfuL4y0Lr5Ip051wloAo7P
Xv8lgIiFViIK7ZFqqECC69WLq1+0Eg3iQRV8beiom3uLm7Im+OoelFXZ6Faj6FNr
tUIReDadI2I8SKFS3F7WmHzeAexXqwa6qIeBqpB7GCJqpqKVkz1CHW0kvS4WAdbE
PAe7FkHuK1W/WrjsHpTqHU8u2IfPYnBISTi12pA1M799dibnd68lxxPJHTpHRp89
uBcflZ1T89AEGQXh6kllaZftYC99P2alpa+QEKOqrkIWgzpLJlmUngC2xI8uPG8L
lmNTwdlCVkHaRyakuIXSHxiIrD8/uAdhmJc+PcIbAU9j6Xlo8fQLaxONwegnD6tR
NW38mLmjiXLvJPDU+xJ6VvZAjU9RDrFF5hcO0H7bbQJvfF898w+MSmRJn6T5JCd1
QwtwkxGwm8ftplPxg9zpV1hwqt3NZUnk80qPjgyBSZPMio0ei4BA7AH8+Q9JXyGo
yAXwxJ+E0rRbeuXZB9Lk5vKbzNd/lnfqZTmsBx52U3RKL5e85N3ouV2GfAw8cDO4
03l/pS3pfz+2thPN0GUM+EY+ROnnAjsl3Um/+z0ZajOcQvnlNjPl4tnSDLNuvBHZ
1mnZcOHd/RmghCxrmBZnAXUws2oF/Lf33soPdgmP24SwqWI7Sl4d6dhDn/xTegE7
ejiCIgtEu02VqZVwMuGhcVR3mQWXsX7xaN2eZA6ZFM7qpMdZCPG2OafEEYmlQ1l0
Nl6lBObeYgwlA+xrmRQRGjdBdMeBdLLnEPIuTZUDTkCfG4qhVwFtAnzm7BfnI6fd
Tz6nqHfdFCu1kD9wVD737u+3K16Wb/uAplf2/wSw/tkwNaCVLGQZqILb2dTWAAWb
hXXZfCv55NHGnC3IajhvjCD1S55It15yBvHt2Sc0SxHsXYKfdgOXIvZmOc9/Qv01
JNNIn63kBuKH8w19707p8cmUDIJ6zLvkh0vSXWGZkafwD318tiWSqPV7z17B8FVQ
eEXiRw3DH3lx7x8Gu2Mv6Q/TbL7gNTeeqN5UrztMqgeSwn8FqGCmvY1tAyoPHvno
sYcQ6qftX2i1G9j0RtE6XGs+e6oINYaGx7ZaFX37NQv6hNquMlUDSy9FOUpmBwrp
r6NjO3vyr3jEhRibhgHHk4AZFQDjhuPTlxdt/jpoFhFd+B8c29yIzF338YaYMF81
LU6ufS/dBM0quoZUuR4G8MW98QlY0Oe4cwKEAw9LVP164NzteMp5SOhrjSGAmXha
NYKxP0Ilp+xhu0PxvZECaRdohdy2AI8ZXaSV9ytulqCa8PpOAmxkaia7Q5PtM8jM
udz3CPJpFU4MQDUUikENa+wtGGlojReXEMDFICJhwQ2o7hZ+9igXSCuj+uM+W9b+
9VdwzvvaOF4njd7XQlUkfL81OpBTSGeDpYGFcr/mYRW+7zHEVXjaiEeLqow8YhWu
2iHhopac4YA8M4ozMQr4aJGYrGaEj1ubG65sjTqMVydBP/kg80ikmMsWh0hbqrIq
x32219hDpY0NNtTBo/JOGFwnhs9+8H3S66NPWCsm8U6osvtSPlCmASDua+XNDKlC
MiRwHGkb46pBZZA4OV9qQ9DKZPlOjJMzJABgtrkz0tRvKQXTait/H2vyVd6gP363
GsVBEskFPyYxnGO4MSdu9WYQDlPOIdMe2ivcjhi4xCxk9NQYYvoBWRTRCMPKdXnb
mZcKPCnd6ypkYMg3Ge5Y3uRtlQGmq4hYE6nsvNGAbYoyJ9/R3cCWh33w/+U7a8N4
4bF6WJJUmk1Qm0BH/sY9pEXKOXxbja9FmqyajK4nhC+vElqZjyGHdLS51AS3Mriu
5+rw27UxRxW8K6M6i8GFSXvtlJIKXIlEbOa5H3TM7GIHSxcuIE2KiQNaJUfMvSiD
HaWiFxzOiZf8nEzEYY4iG11/l5KjLJYI8Cwaa4zcvX8ElzRm6GPvPnVbcNZ5JgYN
600W4aeb364hKtUv7v01HBPfVSbsYs6yfzbhX7Ct6xciQLwmtLWZq5zLBCYVAdH7
T0oilVrbn+tp+yci0moH3PWYnxGy2Fdw3hRm0/G2zJgymnWEqnxzjvH1DdTJ39jw
/QnA8NF6xe3IFmTnD0hiZiAcBX3thjIX3Bqf6x+R9jsYM/iDqx5MH1hmu7sn6FVK
Cg+U20YDhDSavibr8aPppmUiFBwa/JP4xVxYdMGGKKqNzp/iR7KpNw4YuV1bEG5i
SWLfBiUCWkMLzNMIWOw9asbrcRdePxvirc9pFC1eN3VKuMbv3PeBAT5l98tcqnte
vVpqcNj0ihVzn2iGtvgH5GpPxToKfM/2YvjTf0A0FhuONWzeY8exQoxmaefhJhSy
qqhExqBL7FhXvDrPV7d/F3EL/KoyqEYOcQqENetq6bI7FObtLTrjxwLOfuuPZ/O+
M9qKHlGFYdAENMQRAOjhep5TW6ylNOJN/lF74lgCb6WcJUs2ICaGqo1IQ/yyjP6I
yqNxhdd7Pt7TPaOksV0ibeq2O3Nfn6aUkeJW2flrXH3FESRVQjWmg+EzCoLwLI1H
CzV2w42grABiUmC0NdFu6zyiN/GMSLKkdieLjuv6B0+7zLQzWvNsyd276A/jjP/P
tRUbZTU0vc/HBOp4dMORbn/Y2iS2CQtv0w61LE6W3Rp9993VWXVOKQGxJ3+46UyQ
dChzJHw/U5wkQf3PSa3jeTkzexOa+rYGhuCbStnN4cWrUPI/e/4UGdZdK9BsmtJ/
tEiw3CdvzeBv8vDdeplrDQ==
`protect END_PROTECTED
