`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rqe2UBWY3bHvWDFK2vOE9qWvuJZBfLjW1yDH7z6DRza4hRi1evVVIeo8nSXY+Cca
RXnpKb66b2c95ADv219Y+g/GSv3YRL3ToaFXJMUlMx6M+6eroml9ZaNErT6awDf7
gRLGl/W0syBBDAdxGPIRt8iAF5XbiTmAYN+if/yrgaJiNCPqC18yczvXiyntrTNR
LmSm0m8mckt4Ormt4vFVRhH+W0uxCs7HHfsa9XzAP8qz54dKT4sv3wa4Jlp8JnIX
kPF09+mmFli/pNh//QcyoJYBCWTyLQ3Ccwsxa2dRVx5B3X0uNR/X78P9wpozGTuB
thRxXc8wcYiEYikRCmK6qwbHoqO2RwChq5Wa7Y/gL9qjAkwXnCWwdwz6hrPpSrRP
95SQ+j48gL08tGM7I0K5mz4EBcajtN3Aqwz2vyPqEnW1/b2eYFdeLy3s0SDXVmIU
ZVI7t+i9zX1YauJ5Yv1Xj/TV6CaC5ByayCOiDf4gQ492iJc7+xJHmwSgjfVJmIPp
XKKXPKqaiZaaibnCX7cA1A45pj3vIJze+KBSE810q368Rxgcr9YoVQV1VJgVdsR1
/MQLtqe9hghuhrbsZoiWKd+bbbha4QUYwolWKa7TAOevKMuEEJwaaVjY73Vnh0Ns
sEV2CPg/+JaCL33tGCRUycxEDzhiHiaHKH0bhKOfrtaI3ZGX7B+ocFPLYHEx+YC7
F4QDU/cf3VV5Fu19gs/9sjkq2R7XzBiVSrs8AakMTSRWS82cKATPfkq33Uf1bp7a
YPFZBcM6NO0XqjYGTML4v+r1rBDxz9Va5mWjcctxMQdtazyXbI2VE9sgHCnpqBfs
1/PV9rLrPJBjr+tEcRCAkvRFmVR/rto6/TWrhVoERopm7AZc2CU68Vrd+tcOobkq
w4ERVRcdgLO1dB95N9RSvd1kV/d1R1PX0VbskRK3jGoAMPO2vo4MEovgw865ccli
+lPHTXAiToAaTESKKkwL2itE9KhCNP/T9jPBNHMgTPr/g15stZLVM+hHV+1lkxCm
/Q7RsKLRuDTSp650gm/fNOWyUvHalGKUFv3FZ25hcw1TjXrMpQf+zXga4/SYG+A4
q/jJ4TvqJR/pTiAqdvA9gLy5Qs/Qx/nqs80CAHwtlADw3qCKFdkc/7pCN9gG2f4h
d/+qk+nKVlE7nzkWYXK2cTq5ooQf4oD2Lsn+oKycLUKZValds+CWhkUz/zmUWmft
Xx17I+AQMyWNxXAZ4DwgMv+G8pkJRKDjfEHVufFvApmgaAg6WT/czQRxtwrY5ccu
oSp0ZupAWYlWEf9B6GpfgPFHaTS6h098mMZ1ZSEpwxCRkzGHRu+q+l5WDgk6TxMn
LctiDVzh6oXsXNX43Uh/ASiu+ukXMIeDrsl6Hp2ZVwsGwEYdyjz50HsFAsdt/b7W
Apw7zudMPQ79LxwhExqjmo6enOzuMPQmqVidBeOzUVbfrD5RygyA/x9X/XBl/67W
YkwZwRnXS9rG5k5apx+o7WZlHGVJSdEPTzlh6DuiB2E2LfhVhFwLTWcCLtQlrDrn
zCF6zNngfXEZRnepykH1uLURXKmQO2DVYJ3EhGhv4IsaKyxZpNjuD0ba9mGWrmTW
2uSH7N5vgNvLsdZmzerYYou+JaKGPxoTK+zjupVK8OPwSnniS8pmNa8guCcCCJA8
cNaOMnYSnhtdSKwte3kV48SOCUeVajer/Z21h9KOQSxe/ulNNTrvjpZAnu4AMEpZ
YevUpBCriUx9i4DCSAvox268KnNOCw84P1bBjJKwdK+m0bYsWJ/gMAoekUswlxe3
S6EJjweeIs2TKZvv8GJRbAKSgw5mFd69R+OiJ4Sw7zLcgVt9Nwn03WYVW3LgXGns
puzGXJeQQcA2CJKmF7Ew1YvI4d28cNCeAOSVJz/s8MOZfa6t6YnaP6ASYAQo72B2
2rRrl5c8uvTiDsy7bakJwRRGSQc+kzsYnUposTpm8yJ0MFPQ4BU8ruHI9LewmOl/
I39bzYS/RtC95aZ1AsutFT6GSk07icexzcwIcKLuo10ZZr/t3hcePbg6iPYwi6rI
ARNBxLxBkxb7uIw3KER0jwUv/7f6MEZxUTA7UcQvvS8oApbmN0TTR3JzBlKAK5HI
uF13Kr/ieoA2sN4KolXRtleG0tvJTr4ZEoWkeNpTDMbQxVdbHCe4cGsoilP75uXh
mHLP7NFvDf5t62PGonN6lc6y6kvhWhlN71kOF6QjYaDHJcU4uwiMTFyICobcYnTw
Yzze35szQTERkUnblinuYIooKrtIUEp/TQGr5tQMJYGkfOM0La5mUQpDfHidUJpR
oFhq5HeiPJ9Rn9EQw2EV0tRp7jogZL9Z92fEWb96QRK9Xl476GOl2OAU0fc+KMKT
8z7h5WD82EU18G/obP2GgkEiDZmCSyjvXWvyCZZF8El5afnlmcG1H1zuxI6BHfXT
A5rMvslsIeAGiQ6yhQLZZk65txoerJqSs/EvbyVC0NPks/PKGTYRTywrtG0GVp0X
BIMVcKS+8qeRR+4VAEYFlMEWi20bCXLFBqVrPmHhZFZJhsVWvvMuPSI3Y4UmG2lE
PRvZX8BFrnVfPXN3/w4Gbv951RsAkfNVY+KPL9zoLOMQd2HXTqV4/TgARlowJ2o0
1guOW4dRmp4vQDe/mjFunBruS+EtM8N/L0JAtn/q1B87EuUczrffy60F96AtkC6E
/vgo/RNuEJFuMMkP2rsNJfX/DPNg/Bed+sUvS3QkeSPVugKEm/7ftND6WQQXhcRf
AnLhDZWjZkDzeTI9YWYvIABvmYeRNFm3TApBpuxr5ask+/mP/o5AiWLqBxQ73M+j
ol/4txpQkJ4ZsRECqukyZX0dnNJsMG/rTea+xjDj0rc46grxgpXodypspB/Uorio
ZyoKW7e0I3mw7FkxspozIdPBi2kWhHbfzWyimdF6ZHGXX8iOpycawvgVHY+zhbYi
WKGHBsUfYlWOKxzRrEVPpYTcqkocuPG1ONEuHKo2WEo1Rq/a3sG6x9b4gQvJ2Hs4
DidVcBiun2oV0Gxt9QDwByUcRfOptWOJgwVN8RiiohFTBa3Yd+rFLeaaogUoAdj/
Nwh+aTmWNeQ/jmVqbpkfNsE+a+X11L36gO6Mz8by5aNnYDJVQKWp4Casvf+XkduK
ob1CtomVABu8ptPoFJ5+WgswYSLydEV0338ioRo3bp9YQTtIsWEroJzlJJralkaD
23bYyKSdUr2i2yWiVZThcJti6RglgMNuglbgVre4IRX9g43bs1knlShAo70AHKGr
tAMvyoFkCj8VJ0VHyuS+91imocm2+MvjUj2dBMnHlUpqvtNhdLtuSe/dR7U6hWnx
bDqEwWcriVqseKbJm20ezJ88u5j0uo9xXkaVyP7T/ykkBjTH2D6EXAUqxqIuBdDB
Kj3LLGz9TaGG2OaKiiTy3GQU7T3LqvYadWgtyHRhoZjqH+0csaBQtCpMpGuihJ9g
5BZp5FS43eHjKuecCYQHQFx+QG5QOC4kXtMv+qKBib8qKETQZopXs3RPTgEvq6wX
JgYVBEg0yAbrabQtrT+HUyJS78IqJtHE5ijXsyE7E4bwYH2gppAGcjfyjSiGKYPs
VsxzbrfXLpDfmMPb70dihwWBxk8sNdUln8EQwWt0VeA=
`protect END_PROTECTED
