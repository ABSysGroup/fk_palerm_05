`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fCEIaC9hVVBNmBZo/AUYJCgUuvpgDUeXfcFCh9Icnyy5jdFv8hWR8gwVSMCMXt0y
f42/EqlAnLLeQJuTlU9EdV5gv6x6IRXF4WG2N3Aj5/xT0KfbEp3XH6GPJ1bfz1nE
wPtVkTkC3nfOwnlp9dx321SvHgdEpinYkdF5MJQWUmY1zVpGzdoVt5pzuMCsHsr2
MAHDDPocUxJZYUcrMJdZFQkxRFL8peTSwAJU3P26kI42pvLekmEY+7e+pwdpIVJ1
d97JULBqMrr30yFhN7XMOtrevzGnt+LlKcmyrg1BhGLPzhvAZX/AvEIqyzQ7VtO4
kbgGqckhzyp9ZXO22j/eTM6rg/Mi151huSoyNP6Se9RgwjbbZ5r22WPphb73/D3A
Tfxa/A2oswbrLLI57O8X+gCr+3MIZf8j3Jv39b/CJZqH1TcZ+hNndsjjAMpPUvSi
bH+BkZNNFdN1iZV+mUkcCxChbmbDlfJ0l8YSlwA9Py9FM4WwfwmEE8u46fFwr7rM
t4a6Ut3RMq4h751jPe43kGut1c4FMLLkg8ONJlPxJQtoMrOzY9L80qM1YBGnBflk
E/N+GdJ4t7+v2VbdgrzomBjAeAd2TWgq+UucSCKM9giaHnXhsfBsSyLOv6HGzhh0
dGDDKhaL56DSGaJvU3PzBLCftBYQ11eHG6adbBcx+pQTPWMxbq2+JJbcasywjU+W
xFvJf9Yk/zpUYEstZc6rbyKiS6NvG3uWCbXr3sKLom/DC2JZ8uh2d5Zw8IC/6hKx
85p0708CCIYdbaioGTR4hVCQm8ah2gXKIW60o3RZoFezJP2LhknaiFFxBH3b5Urg
j14KGCUXCQufI8y2dQoeGS86KWOohRWSclwlUGZLtTyRhRvZN60ONgPR+WXCjUkw
DxhRQ5KIa3G+xk3TnbOZiOIbhfzCEb2DNC1WYvZhhEaxVl1rigVjeU1i+8GG0Ruh
6REKJ2RVcOYhSopHUCLAoKZZ4R+DvqHdtxLFo/InkRUCpB1bAmLkkuZQ6oA5d7Gp
TSB7v4n+s/9NP0dneRLiMdkXOgITGRVEnFc8dBV2Q+Y3zA42DHxiKc4wQuyrMUY8
hGQXyFcNDCMBLTcZWhAVV86N7rZCnQY4wn9vX2Vvc7OuGNs8t7sXTL/636pn7jGY
UpE689PtHgn4ACeOgNPlMJHqPZwWaVy2vAnzOFX4R/JuYbTRUAo6gH7BAJNhxXJl
cKYCf3TvD02p3jZjWwOdVzxZenKsMABZ8FyD1aXflucV3c/S+3GpQvw1Reu+y0bH
tFdACoDXVmt4nOeAZYO071LXuveEd7bCzvwP4XlQMWziZpO1eQuk4wTksflOruYS
gB1CWBGZGj22002EfcNtIl+0a/RjL0S6MRxQXI0eJRdi5NItgESL8Y/okGcSmT/j
CGUO7XUNudYKlcfcJmLkOhflJg/Mq5/s23EbKaPvY8D4oN/Oht7f+uld0N2GTh8F
39/4afmw/XgDLJ19IH68L7y7VTF+310ZYQyBRVVal9703EZgaCAstg3NOYaT1Tsq
Blrl0O1xBQle5OQJJ1ZqkN9zHBUJXw+TmfH4qvTvVCg+nb7JvPafUOL67kW74jZS
8hbZUZWSafbVQd82tVXCtq0YdsQMKuYiwCgrfS9lM2qx6qvuvbGH8dgpGtR+2Py2
5/4Psxswat+zUFk3+L8rMmorwcLz/TBjbi4j5HgbsqhoNjHk/cZ4/8oG+PVHLgwB
GmSsNOGobrpeDcVdhejoGSiK52z9kNlI1TAcebfH5ZWzgvdZksLGan1kjkVrIy/F
BLAuF8e8Ug4aVaLuOviNW2D0/typ9ekXv35ABmFvaVQVzcNtL8fuU3JPXMmTpXzL
D2BbcJdgVizYYFqXqqSAIJdrqvuDmN836DkQnkrViTBIChoCEaCwB83nOrHB3w+A
YDoy/3sgcu7MrpqGtvYd8RMwid+IEgvkc35fYABmmpxkUtOyZNI7vmg80bWF6xek
9aRDF1Qnr7dsfNNq8S74TRYU5AU0kEQX2a1rww3Q9Opnpo2xruZAHbvsLneoqJwm
w3vT+03HJi71hwHNhZtxgH9VUmgcip3bzQV4teYTigSwDECB4MC8izdTfUUDwY91
JTO3jPnYrPEKplYgxZhfj7g0whgYIhuv3aEjyN9acyXvmaCv2OrAn2FuhXgHL9hn
BEb19ettsau5tXSNrl3xe+MkxvRbngQZ5v6qMx7sz0jGg0RioyCkT5H+OJ8KW15E
Y87I/3B9QAycF7ubKA6qoKkG+j7yKxU32UKhDj0serk0v0Qe2H4pQrAMGsUzrVSd
9suTrlvZi+2EiyjxVSPsR2iDcOqn6xFYeRkCTq6BWGtRmudnOiNuttgRo1pEIWHj
nIdeX+5Vh0Y5a9ZfDf3q6gNnfKUNTkxW1K5IBZf3SZsEIjYUXm9CNyMLJwTUx1sZ
YyoyXqkeo7CB7raydu0IhodzxWE7HovpKlDSewBMQb0YmTQQcArReOVXuEmv1j0O
Pb6bX7AV/2dE/KQ/s6Gf9aac7zpOSQUluJ+kUEoXIfYysPEN7E4pWO4SPGDdBHsh
Fo8WvYJBTUTESYR8ZWWPRI2aRb1fgcaOGj8JhgZccrKo/WyxcuvT5a+ahCrTDTa5
Jz9eYZpNx2u4Erp4aYmPXDq0zKoY7D8d7BXamKKBhPTlcC9WO4DMgUOfsHBUlWR7
rCinQ2iAXyF65FdIngie7jOysPVeV5ZI/pu5wSMRl4SfcVKuEeFrWmZ3op4l+h38
ZEmHorUW2vAZkt8Bt/FAWPtVPMTyzjchDkc3iozR9hQ7NznaG7A8Xv8DW045jRrp
VmUZFZ8qEmWce2vPK++67L9MFSbXXtx2VjODNvo++N0uIKwpUpU4nW6XNr8DFgts
TMhujU6DG7a5TJ2d/gI6zzXsl/gtKzqlPyn0TIRvnIPik3ezE2i3WV5rcoxwKpWn
D2SOV6ihLnShzCN4W9MYyVGhvJTp47oXyQ2rYJxKvWFtYZkYrBMjgsiGMu82m4fl
Yy3RvV6LNqFBawehOjC4wh5vz7X6XzpFS8bA8DGK50tGY1CaX5C/SZB+CSgqkkp/
9tnBQti5rYjf9Mm8xC1Rc8VscGu2gaxB1ay4gOIy1Em9RVpDI9Z1/+N9lefTEAbh
gCPybCMQGvO/NMYPio/JsflAwNEqhUkX84OHUioVl8qjyJAY923g/ANoxcVq2f8L
tto+/GE1VdQQfbUTdoV9nprWE3AT9oRJjjB8LuCO5i34vncUuJaWlCcBjkyVanox
E3gqR77Uv6H3uC75ZD4Sn9cBs7aawkt2nwcd4uwjxnaWO4KzDtjfCzyfRptleEQE
fDUB0ZEYteyZu6UULZexo3NvH4GcmKEEbB3TB3yaJiKNOgBAe4ACpCwv04N2n0f0
y9oU3t2hx4K43taRse4wv6urm7O7cM1nRvBikOahP54a256iIlHvOnNdHTYkG7XY
2LBj/SW6Sdhe0jFl1YdIA8yp7g4rRxODpm++yOlEYwX7v36oURzyskHna39efzmb
dlq2FFmH9c++bqi7NirEOdMRG/MAOZTB3n/ppkBMrwxRlXDTAl1jjlk/g1JTlzC0
NnuSDZfHs0H/FpBuN4HBQdtZ/E7Iu1z1BwSCABM5qrOLAtcXh6u6TR5c34wnQwBG
Iclfx3s7mgcihRo9gXv02NJ/k/1Dvv7ZdzsBcItp0xqwmDKfo4IJZQwux6AS0Zrj
e5mFbEy2m8c/RFQMJ06gdWe0qI1hlrXzEPCxotlGuyfGVzOurEaVRpEGIEiqc68G
akj781hYr+8sK+pzgzUcwJiTb4pHxP42hNtUpRJ0FSi3BlONUPzIoRT+tT2cTJiu
yZtuepGlglRG6u1KM1ZQNfQHLIy88Kmsm+kxVH/qVzdeYPIuo7CCEX8H6U+9HSab
KO18ZxhTARfEbwXqfFP9DSxyUIQ8OjeuLY+jdPoZapfJfzv89KTpsme/y0ej//3B
aH5Cu2Ry375Q6D2sW9ZehBPaL/7a+5UHakgxrAMzYQ1gn6SFUn5QpOjIRG+JUks7
8h2FBlP39vTb/d6uP9S4FTtrzbamLX5ypJryPInE+wHkWlvXA+Ix8cghWDqh1YO1
HB6WZP8597OnI623pA9dZ5bEAR7zGKp4MHE9/HLzHtXboWl2rtX1wUDJoQxIoPoB
7+FSFRJVwbIp5forMDMAwQ==
`protect END_PROTECTED
