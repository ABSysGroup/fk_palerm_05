`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
36ad4dMuWHuIgdheV+shvWCVb0iqW4ZhTp44voOPsaqk6SgAbaEzva+HrqVCo32k
xct2zpS80qaCDIxNqgQ3hDjNxHbcSJcOL2nCWfFzZnuobQPeNhhiesO1ZKxBewWj
bkMpcx423CHJtgNdjrfe+d2vXSsMvK/uq31gP+VvrZ/0AMEMbZjwUlbKJGTao2pX
rMEMUSZpHXB3TJPsD2IXQPtJO6or+gtjxHU08EFLsNDVU0ccws7FNTpH9OVK8NJV
tuqIB/IryajQxLhcnp3+rVwWLtJS/9ZMPkSuL6TSD1+Bi3/bjvcSWxfSyq8k4Z1W
B9mRLikVCMLvxd8oDKSr2UxcKa7JboJr5boy6hAUVHcWzcjy4I/eMID17lqR0dLG
bLe8tsz7L5kC7eMXmGKw718andBU3TN9lMncZtAUR76U/268Vch0JByXqOGcTfVV
OfmMJ7JOMi5IRqqqRzaPlhyZtONQyY/RfeKYSpoPUnQPrZqpP3jKnBFjBjlAVYAU
q0bpS9t25Ve0g/dUVnZ/mg==
`protect END_PROTECTED
