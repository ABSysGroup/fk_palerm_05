`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6N/CGRQOMZ5Px9LPF+knHn/XzshoZ0G2MtZQhji+7vGeH3PINArE+Y+qTeGJS69X
MPRvsmWqxP+WiymOsN1DvQkTc6byEN8aTK7IM/CKi81yyZjMmS6TcHCLgc2YgcKY
S9DUkaGo07GB6iTzn1ROuNvm98jge12uiZ4OTCwQtyhg9EMmMcWGqlAL25Gl1xWs
2JdAQfT1I9+ZAiWzeERFG9YlC2s+txJ6rBF56dQzP9C91QVup8zL1IgMb0jH1ylA
vXUd4PjbJSkprAiQbTh1qf8xAzIx9qq2AU3KUPoh9ecFjYsmn4iFyGtnFF9us4UK
ZrdOC9d2mquPgPyaqK92xi4+TI6Reitm71kMmO3p/awZEVC0/bfbjSd3NpkdlJ+S
naKN+fEuwaQZBvwPevD/GMg/vWLqktWTUsfsqw5o/+fcn6pvW4ohChokc14JvfFN
`protect END_PROTECTED
