`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bwzrAK8MtYr3tsvKQ4JyK1uJCErnW2grMi23mC6B2l02jxR0hmnNbgVd6xcilUsy
1hhN0xEUpNtrqqbudKW2d4LfN/9JoVE4y7byjs20eRHKdzCw06WqOb4vdSe+XuyJ
lIZXWWGISWvCig4PZmQaBJQPaQRNOzZcK/cPZ8muYMFuoARLpo55zBOnFIlZmVQN
iUlvWvgmm3WVMmZG79DxLQ0Znw547yu/qdRM9sCR+WrM/jgtuuuiK0nZV8AF3QHC
n2EKNngJmsz7Zd/mGF5E8v2B86HUPZhWcogeRvc5IhEJ95oes5lGKUl2jt5YrbQM
E3gAuGaoVpjP5EBD4s2anlqSzBQl5L3W+NCLN5pF4nIUUCXiiRLx0zPk2Fujg6V2
KTzmywM2Hc5r84RTk1/GLHUuyFzMlPYL+3xQz81K2U12TOQeoZFA4573cc1apQ8C
du9paLNufQFPLUIFkBBXWejzHTWn+p22taLX7SVNhCYM9Zp2Jmw8/l4nFe5rViDM
1cGv/JtHUAQ+rJqB0JwraDtoS2xzTClJMolDSpShNCk6+6nfSY7J0LGgQGt/ZtnU
Y9ZLEIVLAqWD/jqXe62u4jYexoy7eZUtOiZOwtUhwqi9nYhy1rUUQZ5utjt8YstT
/aofxMoCXRdouyyEsDeNEtYBR2IRelBJ5Gr3aYkIsW2IIz1Km9SyZrzbL7I03pbF
SUljOA8GZBl730f3KBEpHJz7UFf7PBu5Ic5cHa8PH4mkQYOCRKf6Z1xr/+IJc9ik
Lty39LkkYdvkeSfb/KOirlVQw5VUMCY2PaVJnvWOM4SJ9qrqlj0s4vjka/4XAflw
/95cfynQwbTtzL/6N8nUeSqsYkMAaeOasAVhCS8cCTDc8arpwyT3LWrU4a01LcxE
nVzXGxXoOwGW0sjEXHUEL9NKyIjy/5prreTn4TqjVAE35u+UE62+IVeK3kqp+8E9
`protect END_PROTECTED
