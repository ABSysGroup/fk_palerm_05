`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ED1yQlvz38xDOK3VsZc0b5ZIO/zRA7d1Yc1QAMHOWN/6ILAF1HoRrqcM4b0JRI9j
Dat5r7EmX1RIhn6iWLqKTiFMuofGc+n+uYl7A8y3Mi6G6t1he4/gInnOSQhYr54j
RQpgoisRLkCVW9AGKqZRg2mdgV3z5L6zndusGjwstpJKLoRAZctSc9ytDQpMtdLH
h/dNPZKxLEfT4fB3kkVE5IRwD+wvVuGQi2ht6kIccfBLQ+74+Mg3SvgYdPalczjl
RW7aoGn1Gia0Rbgcdw9fc3zUE0xAC6uvEFaNVcimaNUIfH1gVWPPh6ppGmJXKllz
F89VxGa1s2pdLpDilo7zeQtnfRlYltRGUp85FkefttToMiv1qYqlEonIUPvxGGSw
72j16bKhRK0gjS9+UNnLV41k91F7Ds/zQNqQAo/dlx9ZFADfVFZsgQA7KmKiqpZj
dkc5IeLaGzTg3BpZv08MrIFSqgs635GYz8GHgocv3aevBZHDWEt3YWjqBDvMpD/x
JfFlJxE9YZIudqWktwztkW+IbMRN7bZX1Zd/qqCqfnniyXTyKvXw1ahD+qr70IXK
vlQsuIjeYhKtfbKDfOc7PHnjNdWwFd2/hwfUFJ66nGEp2cGRB1w3Hb5Cbljg0q5D
xmKzdhRMkQuRLMnGkAVu4pI/bY0yYhW2Mji9VAZ9xqPzBbc5EkDUFzo+wSV6fszR
4O8ppFBIAVv4uRlhOUevEWevfbaJ2iHle432b/sPQJUZvh7S9iUaq5F6dUB9fq9T
HczUgXIREwIvFznSMQCRvIB3MA4OQOmEDRjyESh52th8Nlki+l8A/GeNZwE/6UkH
eh6EcJXc93yW6KIJrPkg+hyW+d1hSqjSV77UpUEMCRG0T9LdogRnonrPbi+Upxdf
X3V0rRZBbxoHg9ZGtqNYseSzsCq9fKKnj+678qd9BLXNr9TXJ+xbtcV53VRvPoZg
aObHR3SU4oeCdccyAb2LCQh9+0luw3CDZMBA4GC7jbe21FXrP5cps2W1rY6a0zMZ
TIoMh+aUPJiQ/JRrjTNAugacxx725MAm7agq/4aMBQqZhTIxlrP3bL4QJxZSNqyp
fYaEw3tShNVCJyd/FcSqJHa/r2ytp7zTqH4bu+h3ZKOoEyV21CQqBKFcMxpscu5C
CTtsl5mr9SGNCTzTXJJzwAM7d6tg4sg8g+d7lqdU7j929a4uiaq1RyEUxXoDRyeq
yg1PME4S+/UGWVAp2KsnxSmXFawfmm3JR81grSD0zGjLueTwRO38+7ccWlal55QS
zKL2ENcL7xZymGMcpRKqw9I6hOjks++t94Wyzpt3lK3BqrCLtVHjwmlDYbbSu8cF
ETeTyBhK17zx/3DnuE8NJ/meuhBn2ln/ToPHrmBzyrKvHuOMd7g4JLt8jAC6YY5R
0rodkG7/mnKNA7Fqj0nrwCRijzB3J8YSbDtGdWboAdIL7RZT8fiLLAkUC9M5PX7F
TuugYGuoMdZCTggtv6aH4Bo8WM+0BP80xM3yYS1fwlsfoScfD37UXcJrV+6COtvN
QLI3Z8gRClbe6TzQOSwsFZEdTxgT69rOtmTZ2WYaDgH/JcXMrdMvwUS/jQGOzN6u
Puf3ynZa80BEd77d5zGJCWLFqUflXVyJdn1KWNQgq4g6Od+Fqn9U37rqACvydYNN
9tbjGDETlFT86aXfnB4p9dK9kC5GkjNDt/P8S2IQB+8gXCdaTe5OoW/E3ZCBUHbf
abiSvbBVcdzXZgUuD3Xx2xCOTtEDlwYlGIcttV1pUYD8O6pTRI0I+Sf0l1UWZQ7t
6Qw2jVz7t/cjGEmM4xGxQ+W+jD+z8fIMxgmL1YIH1y02HBtS8HgCyTqnOkZPCg+q
bJmk1gz2y8OS6NrKTdsDMNHSaBOyN4InraKc//ofwR5At12wAgGGWuqPbohEkcyd
+wHCRspSUyrcmtZIFgynf0Ll39NVAy3q1bNFbjishi+OFxfB1/cONAVM4kX6iVhI
9dhP7Vg8vnLJBHaGdIh3TVVT1EDRvvt24g3faL492FpS9wluLpRdYckczBK61rDK
DXOvjq09fSt4M625UN0Ic4LXSo2hesh8f8rjgKY9XfZcxdwqHMfTFXryZQcJqmR9
t39dq2Rx1AcWQO+/zIREbSrUYzPgSrpWncaxOKwJoM7T4n+FoPL1WicwMVMfQGVS
im2eaPfdWe9kJg3UTYh30lYZFe7ZuK4kB8bM33PJ7TJnpmOYkwB3eDa6PKXe0WUq
ewYM9LXce3vCco8I1KkKUFFXFe4m4Q3nt0rh/wdl3L/Z3YBu2zL2oGPO0YU5hXgx
CEYg313R38NJRTyJWVQYM2KHuwRbWp+1lKwGNKsPkQdn4kk2tfqJXrfwzGO6dpx9
WpUcOa3O2iysLzGn1GW/oV3v9lPAlmUjd24xJfj9XstNN1c9+FRYVYuNnOkkQZ92
YuWa9D/3ztgGMn6afBPZIOxMOLKk1ZXIeyneTGy36LhKW4l0vpUoEjygSA/U0kaL
+OxV6Ay6wXaPhAcIX7vcFR19ZnMJW8BUJ70IHnwyQY3E5uWE0X6nn48hwAaOgbjP
`protect END_PROTECTED
