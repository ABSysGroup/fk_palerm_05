`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wch3b3lNPswDnQbqWFpDAcDS11LP/sCV/sOY3GqRgcmcS3TH7UVLZH5uLHgUxBvj
caUktdWzXSHNoEusj8pvbPzwkIINOyyJSDJ8h1hZ8dn6yHexbkzQ5sgF8wkCwE1L
uTSyC6nKsSD+eA7eeHGIPey/V219HPWntShvAXEl2bFDDlKBcH6ncDk6eXYJuzTs
YKRpr//wVjvEV9nfItdCkMRi9lElWt+Q0NvVs4SUtiQL+RBB21qrqW9BRH0Ct09E
2WKaiQnSXcLzCMh94v+AkUa2AdXvX6Qf2RLZKukvhHtCIX1JUZM/uRzWlfwcJc7c
wLmfusiBZibmgJq2jgROpQ==
`protect END_PROTECTED
