`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eprkRG17aoglhNCCnjzl50Uah/t6j2CXkqaT6P4VQKe8GIS4Psd15WdZt4fcBx2l
o/TtBSKppRJxFeUHJ2wTDMsNJx+f8sJNWwibUs106gGlfy7417ZZKaQxpVr0pCfD
yHu4TABSYdFHDzTeeeZ3OXFvmt4UCPGvGLJSXRGq9JAMdyRjFp6IzAdGjNIP7HVv
52bMS6Ej4Sv+PE7K7dDOMesfq2jRyNcMWepT0lZEItwvfNerRv79InMR2WFdR34d
B46tRzAHPVb1DkADP/OQcapN8WY5qnBe5/K4JNJFeMBwZXYQzQCxs2OxCKyls2B6
1KzkOy+cKfsvCRO8YBpKv12x69W5KP4V8uRNivZjumEfO3ftz2JKHPF8R6EyjA3V
qjo1Ja6V0eiFZKQe5GwPlMag+GB5Ejf9EPY4wRuDKp7VyEx3rnMzzI53XOtgjeMU
gdc8eZE+gLl4va9Is+sqtNV1WGcqAJO8/GO4LGCT1rYM9PsRLcN7pQpI7xuhevgT
oBzjJCYMixbierMqv4UXmm4ngfB04zXETYe0shEYBi9AYagnCsVfwBHco7Wpk+d8
2o3ZLzH4kToDvFo/crhDiNj7Ft0roR8g4I+i11s2rrDfA5Wmv8gtgAnVv4vceazB
A8gNxl7tExrq6wB/6XBRI644tjwAxzBS0l7bHNtUlq+QHmzba9G3+UBOCjmoNmyf
Q3oBbw3dPgjRVQiMyGfHots3R4SRKKG8OdGc5auXkjpuIGXfhi19CxXtr9hSqRxc
7ce2vh4EbOXJ4nkhdxUbrC83joZxAMRUSkvrhBAAqE5D50klI0tUjraJDqQpoPky
l+q+U800RU4rPrOivOV2Er0lXkwj/5TvzgRBKA9ot43oBpSSlSiAiSqMIwv0IURl
b/vP+wMrzW0D7nl6Pb7+uHEuAH71w+W7KG8cw+le2uq+G3BeJBSrSbPWpNn35vDK
gH5NHRB4GOFeqBKNBlUk3vT6bT7ziGqI5GxZefVRyzl4WAwJz+kmMv/WaHw58kGW
qGUuQ1Y1FGynYvdxxrmFx/trS4FI7zMsy1u+921iS6LlBqVTJhYlU+foxhHD3R0U
bCtR9D61QPD6HwVZeBy/pwtOWe0m5SIjOLoAo12YPBgaWsz8n/7WhzswHO4zRqMh
nMs1eipgJDsAt+zLCc+uD8HhISXa0PkjT5ncjWqJjB+rGIpdlgkyt8PsymopJWXQ
hahsgoY/HwCaGBXycBKXhBvbb/zUC8cqt+LZu7VDaowydq2TlHcDGzH3uNk7zDkG
2Xh9HMwql5WeB+FA8VB0AodhchOJBT+6YejfnH1cc3/JU4RBKmsiFvNDcDp19Ism
TyjQNin0SNzMgbT/cwidDNuK1+m7ikUiZImxYYYs7FSg5y1WwuZdqNt1yv/qaii4
b7j8jNjg3fe8vI2h0w1KLjfAm+HXCjkILEg81tcNsRbpSh7xpiBlPFwPkuwoSwit
KPOcpgF775YMN19Ay7mz7McC0/wChp/cpi3kYlPx1zOMTapqdy+zN+8ppw4+WAJA
bZTeHIXnVJjVTNsPpVc6GEnMoWDBXuYmpfMWQR9RmJz3bLG7oE7HMl8HeNqxTXnA
PE0dlzJe8JJSisUVUSs1ySCYjvai5KHfQI5Mj9nklOvGcBj2sMoltjGy5w81BBOp
l9nNxqM6oh80i02f5SnkTcMv830Tjzrru/X/RHLaBkvao0JXhSodsKRz58d7vG5c
sF2b+ui0on4sqB8bTpOT4ox6dtR9S+Pmims/ZCwJctKtIbaVpWvKU08jFKDSyFdC
i1VAFLcTKB1JE0KpbQ9+SNxBLtaO8AbXJorSO4LFG8vULmoHAyHFuIVODEQu7iAx
uk6b7xWOqi71FYOikaxo742XT9jGfaQ0Pk6rea1PCQ9bWXlxPyrxhRAQjtd1FmDR
WxTilwkFObBtGWU5vto3wE74jG/aXmj0qrU21+5JIQexwUwg5JL7LSPa3c3m8ihM
ngS+nDd+Ue5ooKLiaNYypdbjYZHuZuYRjquHAozqVaFtP2RNrZNMjmtQreeWY5nB
HayUvHIFyIoP6XDhqdp0d4ExHFkmP8ZaQ+YRlt9L5SaNy7zeIsYCU+XPi5ntm+kR
XJ+rWUKvR/lJKdLXGG5L8uPqe5ofz8ukYgzFXS3bqce4s9sdvggFcwXRaTkXpDgX
3dTNREU5kcLzcQEpSU5xCzZy7RTOrK9va1NF7uzCoISbK9OH4etkHHwjGjrGnN4G
fkxYDw0wEETfEcfEVWqCmpkDCaapDOiwJK7mWCs87l0HEpnVpP3P0SWM3gS8GfPd
S2/SPMT90X4jinZxBm1g/qvRXZM0sJ4mk0M6oRSRj8vjcxiUbUm46uezjzWLEE+l
WjduFNiFHYfZSYR17KNIdvZHbrFLFFZMbkNQ16Ub0+/hL7yP6PO5u98GESUSKjrU
5oy35ucW+dMwhQdYxq7vtas7hsvT+qD77fD7DIXmHBptUOTxCSl3yHMD27lV0ifg
4rkAJOs7EYdF18gPnHez/ls7NtxlcUcc0k1jg4nj3tmQp26bZ/4hfvGIpD9nNy5x
PgVkpCiSaikykzN1vW97zLZe+IQOm60i+3QGWuT6mYZSP0/F4AiUiPRYVCQHlQ+H
d/eNgdUnvAznzqjljT4YzgNZeTdK5r7QjO1o8eZm5Op/weTgtnMTaK6a9yIzibTl
lU5WlhHmpJDJO2UbPIsCJACNOZUR0yXuKEl02OhdVwFYIoYYWzzDTI1f/zlaX8MK
pdw6BDPry4I/3RzDiG3nLKQkm/UimkYElfLoiPVQUxh7z+YfGJ3TVTBkAGCILGoO
vFtc3RVYVCN5QfdF0rTA3t/+ZX/Ro1Xw4QsFgQw6YCZGViRcYw3i71ANq2L3nMAH
vyN+4DadFK4MP4go+Xfl0+9qB/k+Qo9Sc/lbw8LIz8iWKVeg+gTYpfUEOOACw1IP
ZZXPZNrvP20AvwFyyRi47iVIJXv6bPjgS024aEQrE6QCoUG/7+iEUMny8Jdv5c08
X7Ndq0rWbLo1ZjdByvngaPxHxAPmE7yu2rHcIVzQchxTfCap9EZ/QDJqF3B+dpag
NN3y3PlnpmvwGaQHTNpZivUJXzWgIvfW4AGMZETRh7Hng6FzHcmEJodCNL2j8NX3
sl2QJSkysNu3/FX5ObMntDZ89VQxnw4Ua30h9l0R/XkU6yblGIiV0z063GFdzqKl
e9gxcDIVlirjCotxHGfLhldY7TUgUarcEM08/h3IVdO4y/MSzs2PWLwl2ZnUTlPs
KSelo3kx+IdATuWa18xdOhfGnuY5iDpPS9ZQBsWLTfXHIPQM8+0NBuK3/+x/Y+xa
e+It6qiR0mRZ2P2UhUKQYjCwesozobm1Fg78iqzxWRJV/zHZL7aOOU3mp11HdOGf
MEJrpPm17TXBSM+Jb7T7LSl+uYV26LjpKaF9P9dVJkjCcJEzBqAkUIMU6ZdTBgit
6MXmi1Nx5hK/eFs58r9YBaRk/SPpVBWsKgnFgunVgFDex+SExoLsK8RpmLKA+tGk
5ASxUckqnaw0l1M4GzdIUVpUW9wE9Dw+/+3sV0/psiMgLakupnWSOejxz9gVf+Vd
1bawRf/br9Xa/Dfrf0OHHdzUg/h7UZowwjKJmdpghPIfFsuSEZrcRYlW7/f6qiDD
y9HPQkMRC4gvmdIXq9mumiro0s5V394OppCtZoKTknjygmm3oB9uloZr4gy0ONbK
3z3pTzeTN+kL8MZKG9c1UJ9zQJM+aT5jHTp8fOBn4mx5KW16iQqS2ZooJJ5/Pjsx
k1fvzVhVVtsFTY2sb661881Nev3WAgAMQudOQfffXJk2BQ8UEpeMbWpTHtuN1A5k
5bYZP98EWRoUG2E3MRJoAz+v3/iCL6hpZhqogxYt/R9+hgfpmNAci07B/nhk9EjO
uDyTsErP1nYHhrmupF0dmDysJhwh4O5CFRJxdfonG7MC3J5OKfpmwMMkn0Aqu5bF
QB1XKpdVd0wiqukUflH/Zb0Q4TBtZblD/7v3Z6m7FIsWbNQBQpkIILF3v9S6zua8
kKekkkkwjpaaskd8jwKeXr89jeKJuDsXcoUamYjsc8jNU1RqX59MkMAtBoyGdwNH
dfpEbasf8rNZ5u+CdcJZPvwRrl89PXSOkD5pzaqAgLQ+vCA5yfsfF6FJmbQutl93
v/DfuLXRReFWK2txl6S0KaSalt19OSgq+BR5u+/60YYYUb1iS5iB8P0gxaZBUs1z
rQC7gncrYFgKF8A+/eXqP3DUljjYHqYM3hG8SOxWxni3phiwr0/EbsTDkKgptX1V
RaKZkAwY7ZruNJVHWglklWD4QX8Hv5lNHkdQlPMaajJ+/8FBIOfRjrbtIGisKvXr
y8ZBkSs7fFKmHEZhMOM1U+h89saXsiJbbN1beq1uRff1jK0uR+vFYAJSc9KGg/32
qlYm5yxezKOBImKt8XuvYXfihpmM7anOSgUhn3C8XqG+kkLrkSZwolnikT4x7fwy
1a8i/ZSgz4kzqCb/cIuFelvKH9JaYCB8I1571vyx/MuUsvJSJkqhlK5PBmJbJz12
NozhZZuGhxZMvG8zP1LmFX8DZZBD9rfgpKfmRwD881xvhNj3LGJD2MQRxFaKhQ/Z
yYnEIEqLobM/a5bQ5MQ0/X7ib+EqVHwNLxqiqztumEx6YCq8HRrV6TGpHgYCdxqc
O/y+69VppAQ7YyzLzlkBRqH3i+A4jiLbHXqt/hzIgkBcLQbN1Of2FNm6rtUJBXho
TYl+7kcsR5MifVk4r96G4yVX6mY0vfVh8yp+CoBQZQwc5hwFYatmMurHgd5emE8H
Ib4wLh6hpshMGWYzvdPCOevZqIh/JOwekRtD4b9BOJdTmiJjLWdg4rNKEC6TUimL
cbZ5pNnxsREQkdv9s+G6ZdsDvf0aQjkRi8Ogh6tb/P7x7XVJfTDaB67LOLCVr6S8
dxyt1bwx3qVj8GPr5BSWJqKLUMbt+pa5l41T+XRaoPO52Fww2C/8xltdTmqjuU0a
Cm6vI3Sp0a/OZCjkYVs2cpt8mFOz/NK/WU4CQii8i7hBynXTc9vlnNDx7A5CRhJk
OK0vhEC82LNpspKLR+yLZX3xmhEbksTg++65/knZc2Zg8Eb0wwmdHBzQE+Yma6lt
p2RQrzFSSFrZC6mBHe/bsGv5pVRvyPaHd5uqSDD2oIigKhPGLifTEi8qzjEe7YGX
ggNCr+jpO1fTkdeP4UoKfRsjAVlBfq2YV7dvtRsxcRjMOtsr1mtP2oajKrZ6qNff
ypfGcVqN/WoBPWk8IcsGWLFPCkljgQLHjNrtmCA+tGnNstiuonH27AK7YyNLUUAJ
ghmD25KAtImuIcpoQctlCluqOZCdziwzsilUaaV+PqlMaQ16gjeg84Xr9ce5STKJ
/2/WXMSpeDtAwgtVXOCbtz3ztqy27+Sx0nDAWWBqg5wlJZXippkYWwqnpbkfhE1U
o1S9pRe3+MzGLKRTH9sZ9bOUuh0SCmIMMF5YN+6mfRG1A6XYa2wF0HNP8P85PESv
wgeuVfE2mGV6j6ILakKORqX210Ie3i96pDb5dmLQsCW5vdfFfToSoUdURehDZw8r
LeQJGjTq9P/UNISz1kKl9gTPFnNo1dJ6VPa3KWFEslahwJnXp3VtMe8WO8Q8qNgO
Mk04l676NKKor0yIFtKRAFc2kMwYKYd9DJ5zWm7YwGQTIGTWjN0nuTQBfKJl1ivI
6PsuSaFqxqnXqK/bJ0+0YGoBBLH9K2WEB/Yc5s9EHLePdHb3W9EFNzypqeWKPcaV
/gSsa+V+oi725pBYu4e5thQNkJDhBniErKek9OHYOi5VmJSBKHB71WERVKIbn6ar
/WkoN2K3foLlAddMWJTq73DjhfkEWi4pgSR7hpepj9Xa/eeJvzj2zbxGl/utRb7i
TGblZnJf61RQB0NfE2XRg97LmqENhUQ+qGjrgvN5dUh0Zmk9cwamECGXjFAr/rqq
ZoIEZ1AnSPk4VO37+2fJP62SPPCAKgtvr5jvCbbsjtcit2HSVkeu0CXuM2MMX7Iq
uKhMMQfis3iEaab8jNssdwCBOHa+E1kTd2KeKwJqwwsEXl1crvMv4DvciwQFAUdf
RE9XhVXPtb/JCYYZ79pN2tFQaC8asX7TbL3MGS9KJoJG1KpMlcA08aswLBPl7ksR
qWxpaUdSdPWLGFpJ2KBuJzZ9VI6EdIp3xATdpoE0ChDtNaYv9GLK0Lu67zl4HRF9
vEDB66Zn+UMOQPUTVCicT/lMIXNZlBSyQnx7VjXGNfRjja5VWkb+pQg/FFKNPgYx
eAG8fTjTlFdMMExPGr0cEB90655+zJQ8eb8ICnDbvqF0klnht4EZ/pdyvmAIZ+m5
DVgZbLKCYNkKA5nH6aJb8SA6I3RlEjv+vf6VoF7lJ38pavxAjP5jmKtiBr88dFCs
L74UABmYXd0UE5DIsfyx7r8RsnZ8dA8UP6M5oyV8BhSdmlpff+j96ZnQr//5Fotk
/i6xdd2SmxpjJPazumNo5DKip0U77g10cMy7UnuAV99ZmDcDjp7Ar5tZJLSZZAY/
u9lGOa9NHl5lpyEZcENTMqnQjLsUjyLbg8qqpXABhdyDGOaaZhfJKU9Tg7VGrrL6
y9SKsaDKnoALlNicpKvb5MRHReuhVmv4gMh1MH5zojgnoUBpBVY14lo8NBoTrLMn
qPG+uOICtrUZ0QdtmAOVVFDNQ1YTFFsx1YPqW84zTPqjWyvxIvQHoZ5Yr8Iso5qN
tA1Cv4Ld85uYtmpdTJYKs6GxBVMKwwSDBS0b7FJK33LYM2ARdiOKMinpKdJPJfVK
y994Hp16EtZJi5uS+9hpXQCHMoqmBjZDhSec6Vz8WEqlYLhUga21iPexJdG//5xz
KswyhDyzTos46dSJsMXN1pIF4VlwpRPFQrQrakRngxzwjpE6CmZljAJZquj4Wqqh
BCOvjabFy8hxqFjr1NoR0YpGHp4ZuhWdu8PDEuDtQACaUAPa/kvtrnXvxzBJUhmK
vfkyOPe8A3vJY/Y4lxOX6yXy1hMOnhQh4vsYwCprH2Q4iW2sRKKwJfEOnvyNQPBM
R91bKzbRS4JScsN7CwX752YYf/05TjyUI/KfIClSuQf5zhCBjAgVoJ3jqPJq4CBd
00xcFG6A/gaLnkG4UOCmhUtg+RwjNT2EPmzJAIJrnqjOE2NIH9s8Ky/zH0MU77mg
sEjNfa7/o55PPxu88V3mEcnUD24YPriXL1MxYk7ddvX4rZHJbONTbKsZWBgFTx2P
/RnwIoJex/pQRpAqUu4pPR9/q6QvTnLs93XSjhCdIpOooOfx+fAY0UWw9PKNSyjr
5CvqbDx4PmWm8iitv+T5gQQ+IzdsYxmiLvFlwlfsyNJzM4oi3fazhxflMvFzwwhg
a24yOvAtvwaqss7c/zdvxrlO6APxTJrZ54XBZTQWny+2+eWhCYhu5JxixQqhT+hW
2Kw11exm28N6C0iXWM7GZoMNHwNvfkLTETCqNf8BN0rgb8J9Tmr3nYZARmXxVdaS
5OiKCaiSc9ksv6mUuaYdGTC6LQuLaYwJkVoPiRUtBef+roQDWItdNHq5hJuiwSdp
qjQdLjHhBiCgvjC7/VwxyI9q3doUbvPv84Jy92ZKiwGFDcSrEDPGO4bLp4LPXwIy
AysxS/fJSo4Xilh89g3RUajPD+qniP0yaGUpm2Ae6SzX5seRRrXQ7erxkRRxp+H0
1wm9yidckWyom8b4s9MkuMiGfBdHpRRD+UsdGEDTiMUFzV7FjTgDQ/Mj7sYmvrMQ
01LGZ3PSPEDQIRdeIICIofD2Agsc/QtGSLFGU6bZBQJbkt0UYJogoPKFsFl4z5CR
s3uESgv7PFetO/vPQAwPHsDS+L0L5ZM9y0jGQy2MRN7oBeMhfVDgyOGUMQUiwxtg
uw7/auoP5K67ttu3Mrjv6E+yJYU5f5oVVckV/5LEqyYAB33JIAt71bSmMKaZrhhW
KZR0vTHD3hxI+dxt218mlRGEWw39g/NPRdMNgLc+J6a5xIMvDh/CQRU5M0huJ4I9
0L2BDeS9L3rw9CDgNaNGgvReYteKsFYRv03vUwE1Ddx7+WBVgPHwy9OdlUSWPYRU
WXeJubblnA9FMHpei8Tj6MxizHiNaklOWPdTH0ZEnn0HncJFJUAIk91kQ0PK/xSI
TN0C8F+gCBgqLhaOrsPGFGbde8XFt9tT5Bylh1s/oxo3EK6nZpkEHh246gWyqmi7
aQyjbts9oFs/43nBdvtLAWPtUsHrQjmrkqIrjqgyE+5IDJpz/38HZLu7w5sbb4tO
WpeZl7gH1I3kMvTlkgkI+5MXJN0uIkH6g42y3FHDUUEBpShrb6AMCC2XebT0Wdvy
2eHziPqI+T4W1RaNApakZ8mWs5jQ2pjpLTDOYttPblDbBwmHLbMc6S65naEjkVrp
5/xJZOhQBw97+WCVz+OSu4wf4zdoSgEvCZf9YssrRBmUrGj5hcooKhXiP7C9jT6J
uJQ4YrArxXMjcParnNsK+pdIF8busRkTo4pIQJbmJz05dM7ZGBJiGj6TB1KeatWP
2O1zfv/xeQqaZd2AiJ4P0mA6zCahxZv2ITvDPhN9g/iQnUowe91WMJQtg+WyUISF
XovUDf9xxJajkGN2bCYXJ5XkQHCcvBbbteWKf5/YkPVJsa7Wy1eSfITmcbenqKNK
WFgK/CKPT8i3hl4Tsvv3XYY/ZcTtX7VD725x0HuFsHte2YEU4Nly1n9txDP+Obdw
IBx9VhLMdZnvfeWZGq0g0f5/d778YEUtu+e3+RrCueHRb+l9+Vp8Ye+m//e1drGL
Br0EvC5GO6d890IGP7IFUBSxELsmfS0c+PgoGeN9he/3XrOOLm4hM/HkCUmVHZM0
u+bt7DYAX57xn4V8DC9YPc7SKlvCil1EySakmleYqxt0Obe4Io9uLD/1zPbKR2IZ
wGG4GHOef1Lx6ydpNGs8SI0xMTViIe4CqS+iXiTu871FhgO5Y+9Dzr4A1j18pXgN
/4+l1xZ902/h0uD+V3kwOmmeuouqk9A3sKocD4CUBxn0rq2Uq3/JES8u2eSlQXia
OQXoyweJ6Lu+nmHTg7Uf82UF1tOi1P3EYssjb2r0xELPsW/FMkW/ek7o6AWsKH2R
Z404CVIP2fr+rECHXhZwcVKCwFzC/7fEefysurTbmyQV6hzsrKjKEUs3Aglvak1D
XBHDRyRc7UHNkgKZH4vk6FqS9kYTy6B12F0Ia0tQ/LbAQ+wWg49+jUmJLulFR0wx
/Y+7YyCZ2Ql1llwjKIInKmie+4d8eSJpt0siBnMey7DysVpCBUdVwqFFw5x82g97
WRrngqiffTekwU9nqRm+1M5JUtJH8SOjbWQYw3PICJt3GBrhiK1fCo53foUgwwkd
ct17wsgz5X09noygWKt7EUYNbkB6tlN1FLBzF1UCs7yHWcd5JohmsT8hI8D3cVDV
YsmEloVB0Bsy/kOC0tjhttqVYAd51J92E5lCpwX2Ffh/OVkx/R4PvaPa0lVwC7r3
7N3nRBsVMNmBjJFZXnSN9SS+BNqbNyC2jXg9KxZ7PzHqwb/xoU+83q+NAP1Otj7v
N2lHXGWXAsUZh3SBBDNOZx7tgJGcnoB7o2z3a98ecgdBwmgvwvzI6B4w6yUaK9n5
ED4FPEfwbeOszlsv/kvOgy53eDetfeKdhdEAqbxlQi2yXqFmJwk5/QZZmr3NfUH8
XdfdfaF6GzoIIR4TW/T+s91S+rYGemrKbhBbL9OeXmy4bMB/yTTXrzTx085ojFoZ
sisoj8XxEy2BuqZsXctgCf5TuyqbUe9S9o8g5ZYg1YOMR82ZvLLsxxZ6YqrVIGRg
1URWmPetAVKTqHRK6q98PHkuBE4u5Yj64pvlb2cyVQa63bOZCf6N30G+Fcj7HfXx
Dy/edOi8TAXISP65MZR/xE9M9V8ysKyXfWGs1RSpyt9gF7EsZKgTgc864yxumyAF
IfaviFIxHdS8FRxH9osRNgXJO1s16+CJjPOB0Hx7jBfVi6U82hI5i0/WkLZwtzqd
0qFiMLLGHLbA3mwZ+gh79GpjaXa7AIujKGNVNTNopR3gQSUIOPy6KAW24WenBbVz
vRtXz1DWCINZjDMQuygDmE3H1Bsp7FShSN/OZW0knI+QuH8RXakKfPKdV6n+1cCc
KOp3FJVWTGohjGvjyvoNYlLvNdcmpycFcIHFBLUhrH43FbXt+1cD9OCS46YGRsG3
naWZEax1jlsZi+FKNriFCdOKcPCBO0TwSPh1GJUNvQ2zVfwN7T/kKQ6Rbz6Gbc8a
AR2ggklbqYDOLRjhItwW6me6HscZpQEo44McXCY8OVUKFfnNU9RV30KUc1ifv0QU
Q+BFiAcJY9E9FTnmMLSLv7E7NG95GkqTjKfimSOnWt13b7xS+809CmSpXNVxbdC9
ucGitRrbZAECHTLc72NFNSvkmm1+EBEAfgo95/UznzU/aa8a3EPPNcLTlks9BfH6
NtCVaDDOdx3mYd/Uiqv8QSTV6qrdpSXZX3YOIq+sDI+p1t9yzCSBFYPkJCXIECna
B6oHCk4YdpB6S/IOyjTxuVig//0kiy+V5zFXMC3mAiBfioJIjdkfJKyir/YifrSU
bUxY0w/ZasNECtFrLXnmqrOiJtQ3j/63T0DK49eQKEuW1JTMC6z4Dv9mL47fed52
ES/hzhHiAT5tX5Ql2WxJlGbyOSLW2X9Ewn4TR0am/m1G7E93QvOidwKJ9TzrPfPw
TyY937L94vmWsX4xpF/uj9BCpXMiCwJ8qONy/A8tShvX+fbwwYO0ywV2K663dsN/
ZSaJZI0bN3HGRc83H2lm7p1hqTB1I+ld0CPwJODxVbpkw4w5ZiweuStLKDT/oVYv
iZckbh5dNmV1fYk6W8wjT0Fm0IW/j7Yu7wVTm/jkrqm+C1FVwQLke25Q427/AItA
fC3YWF4YxgIAvr+wY9bLtckNn4I1hhYMoVzkbv3h2FgWlidYa2gsyB6s3sQ9ae2E
RO6JRpzJT79xSNRjQLc+U/SMYgGrBgrTzp68hHR6faNL0YWdD9ThJmIOMfwix0S+
x5nHDqcjHhuePN+9nxkMnevIDkX6hZHClGbu0kdssVgksMpV3ckM6VyO7ZQLkZBc
QlW40cwrAMS8Sn9VWDveRIp+656J4gzvg5YF/skY0TYJmzhYsEXMDnqBUyeC9kwV
vxb21Di2/FlCH/W7J4y3/1uUx2eZKTIz6p9N9wN/gdInxdoOk4bDbhMjvAiXUI8R
4SvwgFBxGjYmCnps/zOsNJFF5szFIJstC7r0gxKapN22UwqtLq+IP4k4xSmW0Oay
YTrerx6bJgUXH/Tu6W3SUX+xTbP9j70Aw0679qN0FaBVmTRMfudTtYFO8hdXIZSs
DY5AVUwnmQQ2YmSFsAq+MAMW+kDJVYYgETsQqwu/fCg0W9TbXHMLvGpRtMRAvPS5
1whsCssGxKZURE5Q8SmvboGzAXXPGHpEuiAvOXMgWRBrpJ0wj+WkICYfjrpKeQIO
IeDxTAnV4atBFKBncnv+cYi1I+I+nLAvWaRe/fjsZl68TAbf2BFNRfoMIwDGbgNQ
Q8iwBU1OA1KF63lWZBTh/bzwY3hHzMTD85NvJx6fdJcoKyTQB3etogW7P/7tWwMG
EZ291tTtQvkinYEdREOUaZEaStRXwqVy+zIGt5qwus46KHmJ7i68zQX67el3nTgJ
iRveJDbbXG8yQOYFO6I4dNrAq1zx/JODdPVnuF9zmTuNPjbqhBiOJ1YWYGTenx9T
XPTDPzurI/IAS8TMnw9nD2zKc7NqEFib10NuM8AMuZza9DFBSJB5SSgEdJlEPwDv
pShdkUW2W7kqNkNwVuWHaXDNaKRdQn5V2O6vna1BT3DMyZWo2XViNoro2IW86aaO
NZ40k3dO4qOZt5/LxzromtYSehtG2b/bzdoZxdWNHKT8pr9+Jt6oDGzHYzEiFPYN
k63GPv+WG41kvVkiZNN7R8e3+6JIzwXRG93plyCMHY4sUeyaqkPG1d0p57/oabpT
tBN+ZL383APCUvVjy2fklSe6U+AQZwv0Lp1EbVSkNGr6Nox8XqouMN1p9kMtC2Mj
13hQ8ctynsLIPm2hU0c2IpVe8f9sd3pHJWMwl/ABp85SH0RKGIWjk3BbBdZdd0Ly
ybOZbtDu1e8av2vBl537g3pJPYLahF9T5kO128bR3VYUEyWJAIe/rVXn+tkJICX/
9NitSW1UJoSxckR9d0MzxrJjq/OnNQz03vFPWd/k+znzfe12ZNfDO4JzMbWf6CGR
V7Ke86VgPdb2/SG/w+F02X+3gqFnK6FdMx0VF7qJXvQ71VcCcRUWr/i9G+2lUeGz
h6dotp94DkZxlQQhKbshhamaUBBhV/WtEXZ6/d4Q/E5Oor26pWW/Ev9Rqrjxq1HC
LxKRbeSlgGr8wE7xYt9te3tJM/SQO03QS3IO2IPahu6X9neymj2kcsCQmy0cII6K
PrOGVxwhikJ9UcZeVdRRu3pwV5e3Tm57cS48K/rIwFZvUnDLou9Vl+zXlT0HS80I
pg4qU5v26OKYJHhy6MupK1sBEhJ4IFriK5y5VqN5Xakk0qQ4aIMZgC43GjM4O6uz
ZbFMcECoGlugXOHOdJbYWgC5omdwH0NyRqUsvO9/W69H6iutCUBBTulVVUmsa0kx
`protect END_PROTECTED
