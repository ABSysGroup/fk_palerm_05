`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KBHtcnDmO4DcgzOUAJaUVWHHfpsKGiiIuM1ioFzCj1Ofdz6NWJMl50pqFVdxhWjG
hzxxv1HJIILMBeZYQfp3BSg8yVQ6OhhpKVHrDJfP8tsP4BC4XZ4j6Yoi8FXDx3gB
kKtt9t3vBlrMbgJ77rl5ib6FRIvsgfij5Fd9Exqi9Fg7+I1UsB+4PnyfYtteJL1C
9DcfApI1vyqDSzUX5aIkouB3ihYbUwJVVbsR6D90cpkd1XMKrqRrPwVYaaVKmHvy
yLKVs5rzDo0TYBxDvKjX1JE8vHlYJxyyUg23b5ctcklwm2zcVwMGuHKtO664KX2q
vlUltBCAH4diR4zK2IR3HikTWJCPBCfvnOTmHSKsfA+pigpmJa0JWpr5t007tdrC
GZT2eZlfNeDy0jhmDYnUs4OKNcN/LdUGs9gL9NyHTZoE6HFdjCoeUHTbC+f/MfLU
Db/VU6HjlFtZe//5hEIQk+IKBIDs7/zF0qIH+/RnInOrQ1PiXTw1stK6ksAV96yf
kKwJL3tDnGXYRF31WyGdPBq7sdzWn3LXOOX9VnLR+w8TzcSnxnzTtmcXIOFXWRjG
5yrXfrUB2MIRV82NOuV5zAbF4+KVvYKjel0dq+LlSC1zK+zNH1v2XpfQNaYOgKzo
AVjSBnc6sXrVosVOh5yeIUMW95zvw1hwk+NfPA/S45x6PG8u9oRVU+L2dxvsTTw4
yW04Q5A1TgsuryhysFgziKqYuOgCEh0UC9C9Bo5zLqj8osOHRpszyDS69IP8nZGP
MgQyv/4HwzU4LmrG5HIrMfaPAO0rqej+nCl0D+Hog8IfYQMGq1kbPLsweXKf5+AR
`protect END_PROTECTED
