`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rU3HEr17f8qLTy8jKiEImn9gwcr2fYp0nf7KPVKMmXoq7/GuihVQyeC0EPlsd+kH
kFSxKk/Esq3JpVy/fXYlKdZihVHmJgt2y277SY7tK31G9sHg5c3GkBDFVKvDNccb
DC6t41GA3M/zgan4q2zMgBW97pO7bcCSpxLmtb8EtX0dMtZxk8shABNEnEsJSNLA
LG0iwR2CCAoytiDQnsxVFSpFqzGeYd12ZTmXJzkGb4AUrv8KNeOEh+UlIxmCD8oe
bfn+fRLIWIIiSHjUIwHzebdad2Axo54hkVRFBSOAAxknHqcTASKjgqcjIcrp+S1b
Q4KyxFSZ4FOJqfDkjfLIVzCCDznnmNM/1BbKLH5DIBjxLqOXPr6GnTm4XqTUBBkb
+hsSIkg2pLlmuRx4qleQOaX/Tg6NF+UMAZorEI39p/5N2mV//AEIn2cWpOgjiiyI
2b4pqGsclm7TjAuyigLFHQMdYQE6Y6vSJ1hIQBJPRmxExYzXnLNpN3XlSl4+jbo+
K6gCCbTRRf4HvFTM8uO12Wzaxh8npZTTM/QVQubpl37RMuumugtsqMe+97gng6Vo
NGDHc4s7JjvEuzuqC+C8fgWL4fgvrxDc/EmG0fGQ4HQumOlTII9Hk8L+Wnnqr35C
ucGwkjqiKB71ZFFo+A+haG3j7RkLlLREu74Wz8Z3Su7IC3O89OKWuzu9aQfUahn9
FgzH3uXAZR2L8zrV0JjbKqKAr6HxDMjeLVIWMOxVtpeGo86doHjVG6gJ9+tGaZjg
FlKfQXPHGDHdfwspX3iHbq8nMUZrn1eUN0r4SxIXdSOb2/DgHFWixCO4ktXJBbC0
z+E89UXLqqQPvM9QrSZ9JMk5yMwKefL8tSL6hHlwVpG/hYwiO+byc9oqJCvmDXst
EWZJH+SbsmOATVrnsBPL2XJ2uvzqS/wAavjFlGhE9Gj7EWOpR0VhXNPV2N59Etwy
`protect END_PROTECTED
