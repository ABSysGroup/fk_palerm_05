`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BpnEw7q3BW8bDL4e3SM1QET0qr8xvPSqvRwDdWRDXM0QmWwyhMyzcfwCKYCgYRk4
05G8AYV7zTcmO50McQXGHBmVWuCG4BxV/HGBkAlISwiF8L9z3YMW5nJVkEgee6Wm
cTDBJBu2oipN0r0mZFzg6RWwtHXK9CfTuTGwRPdhvC5tlBCH5ids2C95Y1LjUc9x
Tl/hLzDpViAc40KYgedBF9jyeFuActtL9BqqXa8Y9ohSXYpE7WCGH3CrWEecCToX
KtnjZzAfsBA0sgTW2pYfz4/IKbMvkmF+zfD0mCiinqm++Xp9Nc6Bp/XFOzusqR2J
2d6uOBu6bidRRESIgDfs/IezCNtPBsh3QuEeogvndwK5qjlCgbUGL+mAZ285n9oU
yPEu26EPC+n7wmCXRBVmRYDtW8WqaxO5d25hoCxOTOCi3qk+ncIUo9z5Mp59MxKw
08BvSJR9stMqPMgeWqTIY7NetYNvvk2wrEfXn0MWm+gOedF/tZAlF+kpsoy7x0vR
kQVahooFb2jXGh9turgRoIUwZucyV9RTmb70dCeDM4yaZwXwpTZ4H6PPjwLfYT6s
wTdOagYViIj9SeHNf2hDiSFOhT+/sl+HibgACxYWhoj+KVdCxgXJCSFCs9TcBzmy
qUh7uqjk2FetIZxK+Sh+ydhybcaBXF4o3cvXYscdohQgb8w8FSeHPGok7pWCJTs3
ap/1h7zaM6aDsBw3cfoIfc+YHFyqKFjv/N6RHHNtOBXM4QepkyIHqsbxzjqjLlnh
/hBbnuy1oRB2YaVpECPxuQGmlKQKl5frfScHpGWhspLgnRbMdj7law1sCwslUiti
KB3ValRHWi8mYATW+7/QonBuI/UGCIDUIc6rHSpqLbEYDx2B093U78B1j+09cHXT
CQWBxI0FaMAfLBwGqOtCVa6u0x5ZcuC+w0fKLPqdoYdFF28kxZyAVozRn7M9tIRh
ZMNGvSTtnFFhGhD0pFVijvnHD8H5NUd9n50UeMmdf0fP5wv9y4f+YpMP4D4aoVzs
7q/zFzRqNC6WHXeFqn+OpRdP7BYDRKLaN05aB4xSyNujbZTcPvR6gyDW1PH0e5Ch
nv2PhDrjLSxaj+mODmwrw3oPUpSoh2wVLXWllM8s0R3t6P0oKCc4QDxb4dRqoj8L
Nn4+qMdHTKrBJ0PnZd1dPJvZUuByboy+lFXbFZUvxJLpyOmgbN0By09wv41TaYPH
W6qjrKyz3Z4aDzv3Zpoh52tP1gqzrLgEhCtsqONfda94YqtyduAjOXvyCjjiY7XA
AAUGwGfSC/AW4kFwrQ8kL74NG0mSWljCP78fCN6NWERFp/F90y8hi7JT+F/JEzpR
cTSJPfldKiSHdw6pp/EPrRG0EY515Zy2A9NleTHe2qdDJGbwHs2Ia5QGKvgXxgEW
gRFL3DbWecAHoDJOUL+dIvn7/xPgYGGSpp3nrDIN/9pXHSKvEt8oEJKSn4zWeoaP
HHXlRRLSQmzsO/Q33ZTyI0cbz3AuP5XbUHQjGR4vsp8HchNnX/JiHlzyMZeSmtI5
qepLYmMTgai2RfNPoEtUdBFuZ/RydVg/FlROJ3oF5IcC1KOHUZl/etUbbgbdHqdM
r3ROycOIzqUAu46kpXCWBXUKVV8ZHb/8CGz4/FdeNxRLdlPylSCRKLRMDM9/JA0q
x3q8rbPYE68wjQO2Uh6JT7pgZ2LUOSR3+4e5V3K/8C6obJNh/tQ7Ii50KZx5wb90
fHeQip1RuL850clSwgj83mXQkXfuRW4aGjz7PrLKfjJX8Eb6IabY9OaOzXEjdfsH
0cOEZkIDSIlNXvkZH4qRHYESwW9rtCYgxvGDvZPhaYCFaf+Dqsjyhs6BG0YvPTck
2PC7BU+lkzd7B58VcWPyugjpjQq4h5Q5jaATu7swAZ4q0QWAWeA9SsTeiswMJrmv
Ssf5T5DlOSKWjfWfkWJ2yJAvblosh/r/Iu47e16iDR5L8CnTuHo/3YqaOR2fbbPr
SNONldGy1uE2FrU7EFrDLiGM//wodFrv5dFNTpkKDWauiqiI7t5eJlD+7ANJJEVR
7Q4YWjmmwRfeFyJE3PxaH7clBsrrMaINhX+zEXFGYJA/elYAo5E7f2XXZVZJVJz6
5l8PiVmEPiW6NDwHLM4kDBYqCYwlgQ28HZE+lJSg5IW7guoQHck09ZEtDxaMz22s
7fXe0bEzsgh8Dr+IJKeIaHV38Sv1lPsATlPjXvIuqZRJ0ql3RVbTux1ntDeWvk2E
E0xlYxQvOxQqBkfRPHEajgE3wdu12DN4/Bb2Z2+Wh5hbzjqtxRqofnuFxX6OY5d3
94aj6ALleUUpjBicC2O7kJR/2Lq6j2bnhHCQu1D0cUKQ77WvkGkaerV+TI1IwXgd
hmx/3ZtRUMyr1JW73bcyDiCgHrUqMPpu/dWIffpbvkejI1mEOWHzvON7pzh8/Cru
RBZ7Kb2/FKbEPWxwCHFIS4EylgrLFNscOAROVDerLhLWvDnLsIAhnkBD8OTf8IUS
qRq1HHLeA6F64AUse7zPvg==
`protect END_PROTECTED
