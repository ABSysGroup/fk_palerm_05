`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MXmjvnRQq4L7/m5MUrPRCnl7GQ5gsjRH6XOjP6/SKpXkhdj37gVnNdBQg7qBH8E5
rc57aU6CkSWkYodJyog/t4ehkmM0bIDTP2aL1VpuF/ipEuUuK0kMrwY4iWub/96F
53oAvt1ParKkQDsIhCC2699PTeo4oURdNJzucehcr2EE/KG2kmBlQgd8SPYNJkhq
qEpJq6tjedQ6dlgvXNf/1RZLIeaWoKM+IDr92kJWMPErP5XAqP6k549zQ4QxnoEz
uZIyTSX1G8IvW9rg3fUGNFUWVdrE233vImVHbsHp+3k3yWysbNdJPvX1FKcB2DJZ
lswKfdgBHibFTFHHMVRfrZWPMFd+32xvB3ucyid3maCiBuOCbheqOE3HWV4Epo43
jnY4BPju+sgMialPn7837yr6kj0NBOy2CFdcD9BIyFBnhrHhcw26kadXZsypCbXy
O6czwVlcBBsRtkZ+YpNoqaJJry8zQB8fJZSwtNdJLHIsPMo6YFH8/ge1WPNlxtUb
huR6sKgzTv/pAv8WLgp+nkWY80uV1D8kAady5S3s6zX47zuEO3ip/hLQaUXayKWy
mMx6rcLTJ8KpujVKxcjF1HdIzdkdg1gyuBYMdP87/bBR0xUjplgL33cF/NdnFSuj
PmwFIM6+OzZczSGb918ribq6AWjb661UkQlzcZM4aBVRY0JiUaHq7H06eSCFjp0O
GAuvJ/mVNbW7IuZZCRQq5Xw2k7c3NzV+hJREH9sAX9HKYcCjrwwfIZYR+5wE7gj8
RvsRnecgf66mRLqGdfs+RqHaiFsyKDSNqiYBtuSWsWCTgQLmB0m+TW/SBiTF2DEH
3zTOcilc9hfrFNx2vF6Yuhi4lOq4UB/RDZyJU2pd+tJxQkP70PUaI/D/gTIkQDhV
77prCUDzx9SJhe4hh7G0GlZPifN/0FK3OOGyRpwblKL5EKwp0A/uIzZCY0Nm2k0E
`protect END_PROTECTED
