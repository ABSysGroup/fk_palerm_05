`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1X9EyxlHtXzo5I99TYvA7TV0PyYZUY3YmZydHW3gNJKHPgjwJelJX9IPhxkz+12b
TgDs9yQ7k4YfsUboCXiGw51sDsRhuUxqj9dWz9CUq0jgX7yC9zemiyD3qfGIyznL
ZNe7iSdt/Yf8mooAoHWSR0maaxh5f4zINPTMrjRzsuD4Z9FhShc+yS74thJsfLKe
Udu3tU/x1i+17lTTgfl+vxj56d3npWCa40akcl2cRgC2Xx5iYeKpMEWUGNI8VnHu
FFDh9yRE1NcGv6s4Bue1enRSgOkMRl+dhBeLoavYEIeuK8bWchPU2HQqlmkYD0mK
IcaDyM1mKNCSZ0Ke46MW/zW0JhZQJkTWAZH6b9lP5fc9MBr+hu87Y3os4OVAl9x9
3fpcaINZkZ1tt91aTGijeFhzPCZaDuMV+cqjkB6gJlk=
`protect END_PROTECTED
