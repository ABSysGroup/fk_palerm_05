`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L0Laq2Zz5j8H0vFaYVH9JZ13gepHehTGZ53De10dmcJkkd8xOBVpym+Sr2XWHcwr
lFGYao9FOcgMfxRvs8mcLILTnrE316SRydBah7l4N/UHfxRMP99oKXIAI3opCo9M
gDIgAA0z2HicDg3aiAatPp8fMW+kpZCZ4wADr8Ws+yAU2piTSPr/MjuN+VUpT0GD
Ux9MFmHdI2GTSTHvBNsRunAZePQoss3xLN2+ekHPzMcUW0q6ENrW+X2EJ5n+lvew
J+LGcZ5jnORNd+5p/fhmWuKG+Bd+sWUN+BeGkAkak2hkSeQvxUik6YbndgRYmOw7
MJRUyZv1nLGJmr/mkq6rcmqRfMlA2mrMk4nHRrz/4kkn9d8r/xxU/RgOknfCm0Ck
KsFqY6JLctZCDa08mMz6TdbV9HJ/7K9/4Xc7E8xX1QrLPN27NZQvo4RtguMZZ8uF
`protect END_PROTECTED
