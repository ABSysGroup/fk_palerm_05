`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L2xgF6XDxZfC2aN94h+f5Qrumo6VNxqqW/no1nEXWAuI6iV8SHWyjqEVf7nU9J8S
YyVkzlu4qp9sChnCqnhWqTysWr1bHfFEWFPqQx+FuXuxPiz1hVaafNZncwIhD7//
IVte/6HkcSaO8C2U4jsj1R0Sas3uZma2NhfgJnowPVs5Twx4A3oFmMpE7uWbeN1o
FujS++BZd8j0avc6JSM2Qx/N6YGpjM7K2UOrycCBBPFR74V1eqCRBMrp8314rqzz
s0QjXUBODGEtsBOHCiRaGaGaka5fpyvNgmqH0A5hWVBbuDGMqVpgvD3BfgKW073v
Xa0A8pbPAtqj5M8A3Uid54No/SJJt/sdgLoJNNO+8ACw2WTT3xU0vSJhQxqim5FI
FwRalMblTCK4EH4ZcMgxewVqtArdnZUYLo69IEtipc88o4Yr6iH5yMPXLe4g57BY
7Dm6EwOJw4Qhl6IG5ygfjcwJXNXxGap0+Did4KxF58WwOjsq2rp8Skeb7RaO0xLl
CkGFQzyQWTbHCJnWD8QuX72RHeE4zkF8/aYzgl3Wh0pA9i/6tTUVG30nj/RS8Dqh
GkmuBeWo3A1994Ef4aFmqrDrSOPwl+E8HmQwExRtL5gwDaJSngJ+pX4rJ46uUtxF
4rbT/k/f91iB/Q37OoE9XI81imqoxBMPqfWoJuxEFEWb4G6iKeb51ZFYHKBJvlKw
oH8fstMisZddm0cEhuJe9ooc2oNeILu7W/8pLOIfrmXy5tHBy1Hu1GT9zrZR1eAC
7adfzY9wpicOjR//CI85Wo2WGbXC9ZoZbw8FPHLUfljpEf1iGHMPYr0oo9by0/Zs
Ys12runCUwlNMy3CPmjrWZT4Yu+Sw0PXv4jp6gWjDoar5v7KgGl9p5/cyjO+5LKV
wLbYiwTPoyPm1LAbbHlYkRe8ccVId34p+8nU8FfrA8zqFKG2kO0T+cpXXs7EdWqU
v7ADYyaDy7YXCGtUIEciRJz/AIOiGL+8TYuiCj0zPJhmgEiUMsgVbRjKLZ/zmU32
BO4U0v/M/QBwQAaK2Y+RaTC/aLFnRHGZA3zLnpNy3KXA0oDBmE9GVtAF/WHclOFH
osbaHyugPjLZjUzxDCAOsuPEWjpOX8CmNE7Q2mc2T9WvB75SEqjdb04ICOr17Xxy
Pi8JxhKCX2LCeRPLXGP+MwPils9Xlst9J2FgQLis+7P7P1KY3UqLkgjsrXvSDwHR
HfMC1hED1gFtKopFGQEe/PJkSi/vReVYR9HpmKndm9b2v4tOk+L1Hkwk+SWK3nWI
lwbXAYqbrTXyli6+xsw7XMZYNVu6RFeEQrtmkBGM8A/ujNK4c0894tlOijQrJnwL
PqHFZLG18qGcPqpnbRwYric1GFXRvxeBzxcIdwz7H2gsgHVVp4r+s/j+RZrZ03Re
hFZ9KRy1T9OZWEiWk9IlaqwAS5wK2tarGOFoh9skp4p8eFCosK9cQftWEck8bUqK
CD6c/yuxUk/EzSfjDQ7bpoRkXq6ENMLSH3ZLaghe4U2UZKIaXrkHCsZohBZPsAAs
i2Lm+Xwt+Z3Il6v62Pe1izhAyfqWMV+8hPZo1W27qk2LuoJl16tCROHWDim2/5xt
zo/KxlSo+9L8n1yKr9ny7lSCw+UEv8HO7EXMmI6CpVwCrTtVxgMQFFN72aD6rJ/B
VO9S7u+cHdR74pVaqZ7RQ/vXUT0PZDsCjE6+Fl9LV1xR6q3OBrK9lwhLaoYj+75F
O8BYgCzOYScTuql6QcpZszmfUrWcfncBLKuvWjL2PABIzuu5QNfgzE85ipODMccv
bxlb7L5xk2uWmUzjcx81Ok4dxD2+mk09fbBVMz2fpmWeXh4UQFqqtDnDIx+GOxW7
2JgkJ0DkEUiUYxNqABLm/bAGnZJ1QDoiBFWJDwdxhfYI5hB98XC1nky6VE5ZP1nA
qNkfBT36wkm4dWcMVHvgnphgAWVo1k5X60R+C5OPNMJkEhXhBovnYKG6WicM+1KA
TwYluPECNmywsz+93aTywDD1bUNhJihvbw4hhHj+Bav1R8fHRIUreD/Upj2cX/L/
rWtKyHQNMEhmG6gPhFKJQfe+KF2FdVwUhzXw1esSZ0rzFs3dBxgADsjLPf8xBsx8
icR0a7LSjFvj6+FOHpiXIQvtKeLZTlJK8v+rUE7YXyWTK8R5K/mdam31R11goMEG
B17uEaWKfj0bZ4xx5j1Kg0qZ5t3YzBR3kH0Luu9UbXOvOzDWisJT093TOAmM2Ths
hH9Usuap9ovxCBT0Bujr+DhSrOQGcqyyxpoF7esKxZyKDfAXW9N18ajc+SJMZAgb
0xmn67AxBnW6x63X6BNhRCDdZB62C+Cw9LSqAjvk94m7S0yXSTGnbjBVOLwhxnLy
RRsNTFZ74z/HLFFM9T4e2bJ4fKyaSSM1Mb/TIiwlyeCDAom+DH/6jK4XQCnkZtIs
gDxoQ4wB6YuMyZ21UwpaR/3M4uyf+bv+QdIxPD+LtwEiFXwGUJZ05KlOyyJ2arTj
do9Q2SVxyQfVy+Uri8eqfzpdkfaCyd7113z4cKGm68H9rmdP5wyTfJ7sMz+HAfVf
b2UGyQTDJ6QmQwoBkjHqkyc+/atuhLgx6ewNyn5FSuUUDGvi7aP2wvxuycTjWmTV
uCneqU6p8uIj6YOusLONtlh9mDRfTVSzUzs9+4yT0Mmd+I/RzOXH3QIk8WLrvwcc
kb5v1+enZ33KWCSZ5EyEyC+hSIjBYOaCfaGDzCJ21NcTqu2iWamkRtZ8U0HfOTOQ
Tan+yXv9ZAHipHl10hdMknVJmqUkvLePDjJqfk1CI2otaYEluFm0wXVGoU9XLHZ9
tB6hCkfDK4mRsIlIoBXxJF+2k0bKghEJwVY+8l8KTfDT0Eh4N58HfPudmbYquiWq
yTebQ+vlfU5K3FrdLYAyqUiGeZm4mHL0zbI66lOpxu6IryM/llrzlvCBLNsI94Wo
d8vSGhdQ0h1lcoPyqLtm5EcyxiIgCd5ijzHHqr+9R/wOz7vMKltZHNB3Q7QYFr1i
yBzdehbBoc3nJbQcK5yRPoFSDT9/KNvZOl5UwyE6Kac99Yq9OHN3c6d4A7aKL98r
NAkyceYeiixZ5KrWTn6uUfc27NXvniH3yjxwySc7FzPyew2/Yb8O06QmP/G4uqCB
DOXRmallxO9VD7EmSkmO1ubZfnkLp06Ve0lZDTSwYr6kRxIiJgA8oRcz8fmR9JvA
MDsOUwRu9mmZwCVPsrogXkKledgj7mJtGSLLcl9MusD88fEFvyHvQF+XU+vDx4l6
ltmXshaSnFhciWb4mUh/FiX3YRMZKrxrqYPgTG5si1RfdhKDb+MkrYEH5rMAyIy9
p544DlykzK5ca1dPZJFpEaB+zkSX4mA1yWv20GwiqEyRAQTQAeNZF8jZckqVYmzV
o5azZN5Q0U+lrwxxULu23r9Eay+0tqgZp2AKFHpW3wBWTUawM5ag7kzsTcihIJsv
aAAyvIgSwMfY5AH2taRrKRihGLwj+sHi+idKcfyfMf6ZWBPmgb5mqDw6S2DIqwMW
b31nDfzZxAY5ln4mSoij7blWXdxHu2fruCmXExbGkMkqu7/jY1f3/LoFFKDIq0UM
1ncYAPdDSDE9r+kRt8gXgREMcUkLVz7B6tDoWHTq3X9oYEGJZjjQ8BFwhGTY64js
gGLborPCbsMNxN5/oewe2oSPaesCPi5zs3mHXWz0s4UdARM7yYv8Qgj1GFRC/zTE
tj6PGTYPu4+6Sp8+fUbWYV9TRDrowBhLBnmskZdmMZ/7wSP1d3Jxh0sGe10C1NfZ
THiURlAHn0672qS82l14YwLY6d3gj25R+RHvyBdKpzGLn9Wliy66qsafx/mo7JJD
QLlU8er6KMo0iYwxuJhfJjTBU1dFofYoJakIldBYhi+il26us+KcY2DWdc7dJOhG
0URzGwhFmSw/JPKIhDpnYKT47jZ1KPuM0rNaSv8tp65OB+pG2Btji8dwvGsNoduV
xjSszT/v+xrANgavVVaEVC2u7RvH+2QZdMWxhuLMYi7ni788KmYRBwAQK9fqWGYK
lFQR23t4S+YuTBSiBn3IoLzBQcUBljYuadkxv8lVI8TA4xXY88m+EReabaXIDvPZ
jYtWUG3BUGaMrivqN427JUHaHyrLmWYslr/NFiT1+KUWMeem9PSS2JuahgwlpM6r
wvrqAxySD4YZ0UCv1U0qB3FNN9TgSMDoSDPL8LdCVzmhk315rlpBNYXSLusXyuux
bjriX9qOCcIolcVzXs7w4z8loZWVUKj+EsK70g4lLy6Nkn22dW71oHB+uZDCpAYh
DVrUqRu9Qj5o6B0OmdfApI3CdgKguG3+wvTnE/EBn/fi1guIoBPglbl5SkTd+YOS
FcSUDYY4+y1eoYGjU7DmK7OmiJ9z5Qhmie/w4cv2WmAVxsy3/UNplNAhxwrxmxZd
2t2p7qw6cp5lVKvSSrte2g95PkZjJZJ/x0xhHMFwjenUf3v/wBC60cSTWttxMoVl
HDvQJLFb2DORHOkpnIq+DViDdCiruSabZok5JFqOyZ+3oCTW6EpTZJFUelk9XLBB
8o5EJU3bDfo/3Q38FcSlReJCaafvAWcdxBdSmpDlBj8AVM6uVXga4vfJjY3tmJKz
7iG9KFe/usS4CLRC2QuTN/77UX8hhrlAZtIvPHKR6IX7G/3uEhTf/SE6zMLH8QFv
lFgWQp54O9YuVP0GJJQ0Mo/9+JPLhXq+YsILY/BPXpXALxcaU8xpkrcFU7BSeG6c
K3tIMOpYPgWyH8zcWi1jc1iR6szSakQfP+M+U/J9upTrmqk62ZV0YBw/PZNdBGPl
YZKFVZHFy0pE3jJUmCp9Yn8dzCGcHOjMfzO5V0O+PbaMhkGZKmKQUidHZ0NJfA8d
NyrkKCCoAOECLx5SxfMS9zRfWrBSowXiZHi6MW+Gahbeh+YZxOhMgsammjaKPpoy
ghgVnZOEYguQnHYy/lvqO7+YYnmyObbJaQZkVbvKoY2sxd/2dRsqQ/g2CBujvNOd
7zWhifE262LXroW2FnLCRT+mcPOqK3zPMABCnRQkmN49i3de4gH7xfHGbgn4Xals
OaKGAjM0gDCny+uBnVkwZoKpmfEKMfqWXxPBTbQAbjDiFal8qfstOgpAe5PVL20a
6mdu0QwnsK6kX0J+2qTnFdfEebnqNkMYyzT2lMUowQDHh4Lm5U8YjrCzVj8U76rU
oPqTNZbcTZ4prsouruL50RjiRf7iowRkrpo/QbMRenEsJ10BDF8LsFQpXZyW0ZC5
RyQ1IDD/+enYdbOf+8JXDiwE80RRlcJPOJ13KmZwvZAHS8B8eJh1LCjhegfbHtg3
JUqUMxZJxkAQTEXpBY7hntg6xxzkuSYegU9VSueidx22kJ7s8roImnytU141xuWT
ioeVjSpoJXwlZDjixzYdJmwQl/BKnbztna5A7jTS6/cd0mKNXc8Ny1ai6Pp5kf+8
XzBFULhxrB11JzVqpzhogpC+fBFVQp6a6kwO2/o3l9F8ijaAbfGj/lwEaeMny63X
c6Gfo3mZVAfOSB36q8cejKKlZbBc7kMnYb07AOyBq5a2oKfHlDjUfaVZ+wRWFFD0
Pj4sBJOmESBighf+cShSEWg5gbrHP7CM9rRhI0Tbp9DFS92fbv7JTI7IkF5IQ6u2
TKZa4CS+ImB/RCKW2kOA69l9fqYztovTvFPDwvQUI/7WrYyQ9OY9z3QEyjI0S7ab
PE8Q0s9ssAavMaieNYdlIs7aRsC0fsEo3gariO7MKkbvCVDan+9KFzLV2DPi6JNB
d9nvOx2VS9i/yi5KLIyYZCM/PqgCcnxXFi/7OzCU/swWt3XGs/Osl+hqArcb+LfJ
1d2NnUa2EcoABdHiEiH+Yzl2nlDK4yQvbNxkb94/lkL44+mAZZbrLRTRzhzh/44H
LIQJpU4qNlEoPOaJo9/1iKqPK+FU91zcqg6wgzg2uSx3i5QFRBwN6KMC9oxTys2i
zxu5abHjnCO2luNEMKAEYYSuoxeiqMxWhClXjWGzeeFnJU5cHWcVfQDPHbJ9D/6+
JmzrBFALPmccMjILPoZuMjUuDo1BgeP5omliVqxSO/Y71XiZYW3PyjJSW/oDDSKB
AdbfwdqmfxJB9v0fPOd3I+cLRHNqou4g2ZE9jOQVWARYiI7VO/L6dwOzSTacHO2O
FlS2nHFCxa0jeF4xX6basy8SIqAV6t+G3D0UGwlQC33JX00r0YbI7gl8yjQ8HK4i
mVBX8GkeE9Rix0PZYu6pP8m7jjc4rGQMn4xL5hgBgKM9/JhamANUTjIaup+rmqBQ
2+s+TIqe9f59+XrKqBvjD0eaK/7C/+Ognn2DoHoxSNOEMGl+rnn9lqwaEYjojYs2
BlZxWSNO9uAcoiqv4qYKH95ABARkk4J1CXO9lBgMSBpE7yXUIDYTxGvUl65X9dfx
hGTok3AFurlrrqB68lDfq5bX9d9wSM3xAWulLxeGPmOlmJHrUZIsuXD13C87qtij
4CkcMGtOLFK/zOmubpaML8ByDYzqknL67j4iQQSt4te0nFe2D3iy8ZVdyuRMiU+f
wehmBniND+tzGLJP2k/p/Ju+kDZCkqUlh7EmZVf1s8pQX5/w8OJEKD5m9452DrvU
jgytdX/hGy8rWiaBIJ0g2RQy5ZQ6lN3Hy4UX7tHlDYR1GD8mtLRihd6+/L2twrZg
Vm/jk2Pa1z25vh3JPkjehoW0/QJu9k96ZgoeaMZW09L3yEVGqFIamaHlTsdYupSM
j3vjZCPwUAClaOVY+mmiJF55y/b2PvfVk4RtTbxstO7qiDjpHsoHACgPxyKRIp45
NFgSSrA2TSyUUTVKQFzAcU8yoqFBcjHw6ely7EB772xW/oXaRNydYvHhgAQdnFDW
ww+w8tkjjJHHF3Xx4624hDVBHaMTHPEeM2G6zOX6/HTDsGuf0rG9HuSOcl9ZeDx+
nQqtlDnW/mTk3zhb++CVrM4dk5trjcF+Zmt+jyF/XEEqdkRt4ENfnaiD8XuQl4hU
RIogiIUX6aHPWoqtS0B3ORZFc/J9drtAQHBUoLSAsJII8SzuLqlRTFvcBLw8df2g
cU4trXF5y2FwGwl3r5M11mhcjw5dcLFmOKY0Vtgv2YODs7Pu5T7B+D6FQJ8ZzVCZ
5UiLfDBRaQqFsuDX2eeNWKV7+HtQsKk0Ha5zYVWuHgcTL4QaqbxfRfXX18VmhYmQ
Qj4kOHAbYm3MrCfTKqGg9xQFZjw8pjdftbaeTYFlcLHvlJaXLbIAJ0Y23umyw9yK
v/IKQfjBECgviWeFB5pErh9fySPC3gZLCM+cawbShvgK5/G8wV0dbrl3hQ+zfwi3
W/LN+OTmo2PIaV1FfObxlFvK33z4rCq7qQc+iMn3IfGd8BlQkcoblYqvfozn8e5+
YSjEBiKuEpLPd/MmsGMCw+NF3kS5/QHOIEZ5duv5W7Zmql4/DAoylWDmHP2IAQ5d
fb19FKxUjpKnvkSPEt+04l25n9J/xsipdyYyt4Yigl6M3MdUlhQRoMpgJfwyghG0
obuFfP0REDEUINm1g4dV5jFvrXrbkOYEKcDNZNdwROBHbTY7CxX41GgiXu3N9db+
RFP8x2UL5/Nu9MP2X6KrxrZCMLy1GfIgPFM5F8soijCFCm0b8tQqWWvgVYghkIm8
9vujF05VOnE3IRZSy3+k/B6hDkDCVAZwHsHRG7ovcWS1bGJvTohzkXFDMuECL7yS
EsLaOyUF5MLRAt4/qnNz9+ZCycA8CleXvyE/wbxL6A7RFVHO/enD3xL+A6awK6Rj
7ifF7IElab8Il+Sv/YAqk5l07oHtbl00zi17fElDsynqHcWenh6qlPJXDj7iteHI
9SB2G1jqXtXTZJ85r9Jgt9gleRYDXVFexorjkRzhm4nfSw4Kr7B3ZCbiEgnek6KT
/Z1m5OSYrcPSfDAUxqhI8zQb2ZnAgc1Zq0JoTcjukAC4gb5oEzb4CeWLqd9v3LWl
t0j/894c3KoFOjkkXh0wFafaWucA06rExp6oVb/WJI5YVX8oFj/yXa7wk3VKGuxD
Q/q4QKaX8kx0JID/2bGHjdfDGQshizwByMttmaE9GT0f0lawU/FHTeTRfamWrv6z
jFMzyPQIc21aQpyfGKcVFK5erJWQNP3h0t91tRhxc+si6TVUDupeybkx8yw9wuvQ
22qi75QmhmCnVqpjbC75b3OF5ewhescMgrYCIJgDo70oLd7pSr6CFECW9xyBtBXV
EzmDrIF/w7zO9jgivhZaysz9XEp6wjon7/+vXgpKSqSkDNkDP9OgQ9chGxZcX1YN
`protect END_PROTECTED
