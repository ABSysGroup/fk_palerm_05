`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ko5b1hLPPxyhS8OOqtXt9G35s2ciS+/XzZjjNW5HUNO8Sy86WvIIh/JiFwDSVWel
ADyvWCNt+t24ScwVusAjLb83knc8CM0G2N5G3jJfE3I51uMDCfTPNFaVs9RjT9hD
uHqKxmE9OBCIs1NTUGO+MFztJ+1MVIAbIgaHfQ38hptcxF1xYOIrf472NVa7MGIX
ZJ9787hxVKkKHHFsJmxkToVzPgLUSVqkmAg22/edyv/Az1N0vlgOKNtQsPGFGGJW
7HBoOwmUAoyggfDfWrqbOPHkgBQqoOud3RtHLBbgV1SXMEC9AD1picnHNYhZBHfC
gqWPFW4+fH8iW0kPU91d2mAEm8Xf5qsGBB7DuvT1Vu3LogoboGtWpooPAJNVGirh
RTA8BPCUDnsJEDmMwMxiWdeCNJrmmH68DeAOw/v33kCDZqwrterP9M2ltgAsBdlL
vCXTZpfjrPhm5K7pcwzk4wiC5tYc9UUXHovmYhEjb6ZGZPldq971JiCtZyTCVYsn
5+X4JevXA9FHXrg9TB7w0OkBJ3e5OagNsMOl1Td5wnS84PTy5lRaYEapC16L8ynH
Gn18zy15JRzOYhTZFdc9seXkaKwmprmCbYkDY5mBKcSLByoqIelR4g+Wl3CCKKGU
wtl8Fl0RPfI4dkXEm+VjpT6xpNs4hNm/1e6447JAJcY5N1Y5FhB7Ye7KFI4B7vLl
q/LMPfzhWFupzlQiiNzaJsQMXW35B6BZvLPhn32BypkuvMJWmY6h8xPjex41k6BL
0Dcxz06FPN5dNA1BgKfwxcmgg/o7VVxDT1z2rROSM8tXRSI8K7Lb3l8rAdvgwX57
mxytUD8bsqOIyFexJC2dP1D2isX1yAoUvDP2Mt+Ff5F12rymp1kENjSwzOjFhqdZ
1PwnWtB4l+g4GpVSHFY5Vf8GymNa1pACHl7t/tLoRtLpyMg8ZdHL1xh/6zpUgCa2
`protect END_PROTECTED
