`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rPIKYvVSPCheLpq2ye/KSy8DLBFl8rMVVsUdrbuIiCiS61XW8YlMO3+Vbnx22/si
QS7LDBXCR+GcKdqSdf50opgmNt29oyXt8YpLAyVSmjuzR/xoTzdENTSPOmaN1zXW
c1F18jCLODH7ZsRUu5VwnvLjPBGmmXWrqvIESw8P4CvHCJlm9juctYJBXLGGPy8R
IDzV5AvyZbO2iqCxWGuA5MdHwdneXKRPnWoVUoMx7vawASLkdhsIY29om7N/sc1h
t86EAHaFRiwo0zM+iDnLEm6YaAuJAirDg/5iGV3y1TTMRwfb53q8XHts5mpbGqn5
DC6rRC1cJTPi9d22IYTVJxfG5YlU8KJMb+GIwzFf6+Cpf1Oi6VaPxS4FPHjQZBjj
FZp6602iJWqv5ahP3o4Rqh6BIz6PqRDkBBdDd9BNWBRg71moVoMCSvSvd5aHf4hq
pOymw7oagK3LFHe07ojkTD1zm1e69uA7216w9Iu+Wb7Xa6g9mrf65iP91myeAjyM
fmwXCdXwUusPHpwGyEDdebMMuOVswWETy/u9oPDh3fQdLvMckPCVHNeCk8mo1Fab
UHImLrI9fQ8q/+yfEQtqgDyurih4GJftuVR+x8amaWjX+zg2S83WUdUBFK4CZoh/
BBLUaLsoaepKFG+KXgCgbKxrC5IXFR05gs56S7DAzw0FmPRr/ERx444zp09YTPSo
ZjLzFXvsbfQxuSDOu0yPosrqtUKUS43WxlOlUe8O9xNcxP2pds/c9wQ2Kp1xHQ0J
q+Or+qOQrVMclOm8mYpS6C1JIzzA4CN4bRcDTIg2uEc=
`protect END_PROTECTED
