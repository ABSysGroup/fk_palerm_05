`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MbXFqgjUzx/jxEIuOhVtpoxr6owJF1OwjvRR6BjeVze2H+ObLrHCmTv//S0t6WUm
w+tXXPE4E8GrUYi0aREMJ+RgXHsfpATzsVzmqWH/kda8JptihaORCVyb1QhhoC1m
0Y6JfbIt5nbCPq1N1+ywCvtIEwWBntzitGnH3ZM7/uetDAm91OCn2Jfv9U29Rj24
m4zzm6tZNZd0BsDtfRFUUTJALrthRi2xS0JCv5gmju/QEDN3YM2pe/BBEo0bmMSS
lKW3/vrNF1Iaoi5Nifkd9YswwsverRCXCZIvqq/cLLyDjmyaR2keCjF7RngHxaRT
T7eTBh3QZchL2uW9SiAtU8LUs+F+ZkFmu5ZXHzfHKTTyo0rJZXEt8kDBuGPqaAdw
XhvjstkW24LsGgPV2Roez1/MlPLHjf4lAA0I5twyvv5YloL2dzOk/lQUgeNP6y57
rzMb4PJs85lzmyQhYhPuF81qvV12AoyqLujeZrAmCoo9mu9Hj9oqPFkXZCrkvkVo
yDW2S9PMz5PRpPHIpDBcPaKG+LVMYnmMu1nJm4Moagz7DxtDnK3LVM1X99YweR6L
ScY9eFBbVGYAOHMcnBcQkLh7DMtaZZNLOjVhV/2fm9Pi+wgKNT/q5ArJgaztCi28
y4LcM3DptscFIcgYUaTnZAdLOGgALqPdzlXzj2cmLg+0I2QhrWVpJWUy6/ZamEGH
LjwNX/RJFg7qYx45aC5NSqxCuwc7Pqx+G5wHc/qb6Tz2SPm6XNDNsHcmMXwnxgDn
zQkODqUgvBx9UPnGjDCyGwiBqVkFf0BBpv75ElhGMxpmjI2sn5DKngXiJyLQ7A1E
Wkyn8YW/ugR8bqneS+nL6G52xcSvz0lIKkgD8DzuTKB/wUVxuXi2Vj0v2fn61PFE
Ili6QJm2uyLyRCKEoWh+hKWabV/UshXnJRNIxKeZYsFuQYod/7ylxDk9HnJwWPH9
nUXFBLliUizctkECwSOT5DJxAFXA3LBvcwncGSzQAR6t+ELq2zQqzXQiMQjpDrHJ
`protect END_PROTECTED
