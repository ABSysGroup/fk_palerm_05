`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KwRoDYJ0SP/523J3jd6ko2WRuxLntTdoax9l/288BTarYFWDq09Y4ZB3tX95+EQB
6beW7B93vWP80SjHvZHp199zmGc4ZFkBXJvgiOJyTdqHAoChwEc2jdIN80NIs78c
nVtmSkBw3hMNC1i4PCxompJ8IN2kL9LM4Cd/UpyzObti0NZ1O569pDr27x3gcFoW
6R/AMC63q4L/H0DH0ko++0yM9McyIWJNlM0veVkvvqt//EitHb5ruXbBVx5V86Jz
G3q/RZDKyhOCR/GyDq+gKbLOOKQo9NWMfi6tulDyEG78Ot79vXZJ+AIisjWKjEsk
fD7m1Lkk/iSGE8NLTymQ5hStjYQ0Hn4Mz+VaCmRQ4i7ycglydNM1FMcHAYWiVhDe
pwUfDKX8RrTossFsyxTVew==
`protect END_PROTECTED
