`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rZEZo1wrx6THfF3w5N7GAQm2yaksWLBgATbJVZsYi+Us9JK/qVVaoB02ykKLlPjw
zMKQMpZMLbDa0nMBguOy/2wbudMWErtdftEnwidEGyBV0ElcsrSTo3ZTM9sUedKL
6dK4L3meOtN/qHxN0Q6zpkLhIWyvSe/Krkrz9kdbKiiFsLsRZ+InjSUZd5Ww1nhl
CW53piwzFLYD+P7TJXokpDWmLCD/kL8aWiWSFezZBIgxHepzuj4LJ4SJYLWAnBO4
m1dr+R18fazq2adcTpeAXtELfQ5/tyPT8tQDBuMTQclM063y6gnx0/Y/U+bON4Em
LsWvPCc1z3WbWqFtXU2eBckdQkpTMiLKyvXVOHqcthBtaZeb7YzG1Yw5TSNISZwY
NGVuwf7L6OrU3E0wlhRllcpclcRrHcu90B3THl93sxsNXuNpDMYcsAJOUfmtZSX8
7gMgUwdEHFiVAHU/kE2Xkn6xeHNyi4/P/+jcBSK82e6BUMwGOj418CMwbTWmgQV9
j2M0DQiT0l4xLEyyudzLd/yy8qO8DWrBiBawUXkOSAQvYPuJpJQyRWCAlRmo25UD
rTwutGnozAfQe/UX9kXWZ+PARDzaD4GSna7QsnOQTxzx1zXRQHBXU5iKAV7ppuFo
JSR2G6VHuKijqvzs0atQnA==
`protect END_PROTECTED
