`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S7g9BM42KtfVV/1VWsiaaDnx2aVC6FpSd4x+vgd1bRtuXlLUXqWhrbwGb7Ylyt5E
NuDGW8sXHObYSIttD4jfpAW1vlOS5yam3hbL/9y9rxC6sgLZeuWn3l5AqO5c0ZlA
rOrq2gPCVMY7sxkLb5JfIaMU5SMRe8ijyRJy7gbortXhvTiZOicIW1wwZJTAP47L
kf6Eb+bP7wjWJCj7iFmfTkUKqB5cgQkWXjNKdmF9BBdqkxtAFmp+MRjQXGq2j7sT
PLqSkMWmTx9VaqC5bR/zFcCcZ65vwqbYKHxW8ud05OP4ZGlW6pPfQ6RM9v6V91vU
hBToMb4/p/RVTaEYNLFaCNy7ky0Tqcb6XCQYhEgOaP78OHxr4R4waRFJrtMptsaI
NVSgZG9U1NlMxCIYJlkW/wd+rcTd/FkrIWm4IC+paIgFJLkTF826Ur0CAdAT4HVz
Yb6iwdAtQv36u/ndQRgpjYxdaKBA0s9YwJosSZVvo1UFEazoyHJuwzv0T1HLuCxH
ZMuQhArDbiwSFTISEkLUW4XKY3Oh+KvPa7ErY7SDWlJTpCg+w17KezRMjltx8Sbb
b16aK+B0ka1FpFKquMciigoqxPEeCf65UkqDGKKGuX905SDH4NlupP02WEnNK0Je
UQ2L3mMNJSGYcaT/qwPuXfrxkUWDhwZYac5aMlZXJm6NOcTlfUoxsyXI8HQj66zt
1icuptut0drQQ2udFYJPphB5RHe6DEL8Nqsqgi0HCf4VGT8hwccFYRGlM4CJahk2
Z0eVpA96AE7kGvGxq7g4oDg0z8FUllZiPaxwTLe9/cypAUoW3jrrX4nhOxbG7ORD
shc8CxQicAxtEJxMkVi/Djc3he5/yx8kWUou2n72/dzEEXeiamJ0gt9r2COfvy6f
3R0GTE+ak5SpWScu/p62haNaeqVGGDwVp0YiZ00EjOkZoftng6VMaJWfa8Uepz2w
GrPqX8URKvaP5wjYX99wPveW9PVBTabn3j30+mcOl36tMt5rY6nO6ZvWD229dJ3Z
YwbXW3G2YcVirhwRb26EpW4WbGw5bB8T9gPbFjLSOrHxkn6A8Mf5FGMQ736moZyA
CxNq6bwcIJ5b6wZmGiNslFDixtDY4xhNh0D8XhRcY263XVznO29zcR/I6kiNzcz9
xKsjIJiUnS9g2+EPAq6tVvaDE8f2FPaXEiHHUHb3wjElTyOfi1tGboSsbIeUJk27
ZIo+pkQ/6bWMglJnhv1lnCJkgr9UfEI3Kd2arZFCXEOR2chIl3CpFBK6Y/ojKTZV
`protect END_PROTECTED
