`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c9H/Td9Yw4pfH2kS8pAarrEHga7Hv6w6g+JSMvtF1BxNR5JL/m2o/3i8AYWco1/Y
fFJqzi41vPRPfJfNbfODZhiUmEh3xTzVDzG3N273rHeaGE2WpQmNUxhxUs7Rn2h4
NbxqsdiOMYrj55CmleV78R4i0VqUbxvjlZm+skxOG6Z74J6CGMxkVMUN20hKktbp
6JHXEc8Q0slgDM8BIwvJ5i7muaqsHDlXZp0vl2l5jyNaqYFOXQpY4Xi58gicpsyG
jjzkH+igs06mzzhYfnqaqVNqUU0zgX4lpYGwmS9zmS5kW8G2ipuIDCmYuFXsPPPi
q9fWfrxzBxECB5+w7oW4EK35fZc7zBABRoZtC0mcd2X/qXf/vCEBiu88095IdHLQ
wG+NUyo/F+2NS8HVbytym3i6VGQXhpsAL/5yQANIeGw=
`protect END_PROTECTED
