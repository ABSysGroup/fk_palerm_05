`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qlhX1zFSed5dUwU6TimviM1uQCVwcQYahfHzAzXLAYwIAresfQsgkG6po7bdqh5D
4dDoIfwrEqLQgt3o5g89mYcnzH6Ke/qL5rXa+hYlVPe+B8K1MQQ6LxudpYSRSals
ToJN5tgYU8aBka06Qa5xKcd0PfP8IUlX/el+FxgwebjloiQ8CQDu1r5MZhrEgt++
HpvJq+2o+7xrVTzoMOYt+Cfo3VFaq2KVDC9vcXEgIrSWz6TkQqTdMCCjniPKtF2Y
AfbP6vRpwzNvmJPNi90CeQ1xuQc2U/0AW/iUsbzeWvXsDEnPTM4yO4Cy4vedXi3F
yCqqudsmOPDtC35OzUmaiDKz+K/jD/MiztH4ubNn33qegQB3LmLRO0cZS+VSI1ER
BkBSCxvguca/GJN5VmQ10NHvCtlm6FX8H7cRLPLpXY8nl3x9Ule6DwSV5O88mZhL
sFoVpgqtUetihBTB07iQQTc9lAPnILL7C++qaAYj888T+FVZgBFY/Xf/z/+bWMdw
UXY+I9Y6M3cgx/AIVt1pzHCKrzhVz6cGPjoaANcOn00oafKu1bc2zj8/RviQyT0f
6ZRvsv73Hdlr8wXbleISu3aWmjx6OosXtxdLWYFFtDmWiBHQ4MVJrXMykH293UmD
p4fZGsfUxaug14KE6rH+r57vxFdq7M5gBC1H+LtVfLIfHGqimO0VEnawrZluWhF9
omYuoIyJn3DtSy2hZDSefMgHog36f38WPUO4vyay+8kkvUIq0gceJnDSBJOFjcOL
iUva/kW9AGfzbwW1sNHWMGU7RCrNDojOHGpvGG50gCaSCVmVgaKDIEowxtqkcwhR
GNuWlyQG6SRE7HBbreHG10hbwrbGVhfLuDZwKuCUE91x0kNASaYArBpzY7TLBql3
74+asiOQmQBCCam9yVbCrjJT83FFOJGXFMHuJZjUNNWjmequAE6a/B9WGg+tB9jZ
w0oBWd1Yj1gZ6GIQfUwPOjJopL3BIsTO4Czbk0ph61czo266udvpy3jmKq4nS6xG
5EugHMmjoZfxK1BkOAV3z/0XKZ5bTrxntTUzSUdqhqw=
`protect END_PROTECTED
