`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7p8CHNv9EkApt+HXoviEAQue8NzSa5fMYRQ7dC4OluE0r28K2iDQaz30LcTaVzha
SpfpIhYDFoYUs8buyvSOH2wFrzhqgjadBmzBpukDkdYItphzSX6dX8SZUalo6123
yU4R0pPmu7ZcUoDqIvpxZeuGUWPk6+QldD6h1zL/pumK6ZRDRSHZG23f0n9AbjOg
hzGBVNhQTkXu7KT69iUnZno0yGD30Jg/sZxRrwaF/+PnQNIgWvLpbZu1FX9TTsjx
dyLds/6zclvXn1Wu34GAfOQTDrfL/hHRVIoIaBcnDZSjI+HcQVWnde0piXhseWUd
9AdcQXxDCLAn2zIwDh4MlSpjdWoqCjqTU3YAl6EW7hSU6+kIu4WNjEJW5tgctdBE
5FPUnAOBpYgNc1DbhQh8cQRNsuncyuRYWiA7TOP77HAfkQNKespaRVPOe33rWaCE
uVOhL5Rnk9qoqf1jo+XMqcwcR1pfyjpbJtZRYkNqbNP6uXAUjPKKVa4hcVkP3miX
JpjqhgEoiM/j+fHoEEpREl3iYn8wnZx6oDS3ZHBPJ87JoG22SoxNI46gnZW1fNec
R1Zk1y3GxIpQ9gxPW/h9eCNY+UcbKyDlL8fJmCZLrG3NvCYYYkZd7oQYY0zRzYoX
/7uJMkABxm0z255Fv4Ldu2UkDz3sC+MzrwG3NcqNNAK5NYkoVf5X31685BcxrOuI
C8b+o9Flhps9YWNm8jbUs4NmS58OC7BYD9mOsiDIj+7pNBIZ6x5qIvK8Ijhz508p
MsqtPN+QIEkTPCGfh8cMKF7kcdDfRlYTCGcKmC0x32/kiEw/9CyBglekWxiGMxEJ
Z8cPJ+Y7x3ftOQg5miTFWccrDBPS7h3Mr0szUAAm9vNK+OEr1DVqkGHffgEQiahy
l3pOSF749h1orjOJL9KIaLtjtORF4DYkG0yxhHv+FXJVX205upgpVCwX5X/7Vdai
wNAy7kBfH/RHH3scaoT3GM1Mvrt7MIpwysK7eIsSYIANDV8JOb6HAslai2Jbi51w
xRec7QOrQAthhNLT7YOeV/T1DsRRoLN8z1gkEWMCVvmm5iZIud7aNWLGsn1VdM/Z
svqoLNajQhd2C8sEhp4J3KGydBQzhJT/uwqrAKsoNP3Z4RKpObGSZvoxTVbrv/V3
0tXisHDOAkBGnlSvHybdU60Z5e9iJP1yNqU/fRWaK4utnmGntPYXiDjx/s5AIR/C
5a+j/pzxqhanFEa9HRS1GOWXoAa50qaKsJ3pHG208FUJgJ50fLeD62NEAFN6oGmf
rHLDR1MgdxuY2W4JOuZQ/90TpHg01q/hMk3l6pWrm0f9WZeB0jLINDdJRlWiPpZe
8sr51xZMm+5PKlUPyx/PYOb+cfAU4+IRQZNpL9ZSv3pg2sJCYwFqUO7E/H+wnnB+
E1ZbCWm7WBCqGStykeWdMnPvBMNcqD4uWFTr4FnaK5YEpLjBPj0q4w363SCQbJA1
Qr2/DfH4CSf3L2wxTTepSKXTSaFuMxjIgxAQRZYfrCqzNjuEzvWXU21GriNnaI/b
1ERIiSZd5zm8DHJhTES1QPh2G0iRwezOJ7VQrTHHe5oJMsL6qs4QmAHYgg/DKAu9
IeznZ5dmCmzh88W0TpuVa+ZH+IFyNF2m305yPoX+WzqPouHKZHn4sXzxiDq2lR/t
cP1V/3005gNa1O8fIu0mpaIXbx4fiEwfVB0mOOhioaxe+VPpeqdfEjabMAqxHgLO
b9SUzzKOmJWIJmdKRYqe7Lyec7pwe6h9D83VP4KowVqXE6x4jq3YBQJEqIcSrfwN
37UtPFj4ceoyQFBIkya03t77uFmchIfkktOv7nfOhvvVJobpJBYh2tlTsMxw3CBT
KriWFSZ1Bfd3uuzaapfFc6SLsRQUUSzqsgYtd8CvUy7XS/R3BsmGrynvMoofR7v9
bgSZ6CDAP6adYArOWI4lqtjk26RAlbLMTc8pbwewfu0gMlBRxkF4oOH6eQIjTcIi
k3k6hOqy80/b+ZcHUepjBwOl+24lcVskHRwB/ERkukQ2SgMbZkdBsF9a83HyBBVr
lRNAEo9sFSo1LjLmu9CnNd9BxDL5M1EWm5ZN3ZWhipcwoD64IzsGbtvFxKnA0GmD
KTY34v0qVf2TgZ2hEkezx2Cd6gPLP0ut/NpUd54qZp66brnLhbislvpKr+aFmPNU
ep3J2X1vXM6aSnNx+shNxudLHax9LJUDLyReURNW9fuFDmgnKsetwvOdjjS/rsXs
2NGbbixjOKgsAe/3rJCKlzcWyEUrAeM4bw1yJzE3neUEl4rltuySUeDlZxZD0Uua
KAcUaT9yFUUWJffUD2CpEsIzGvstISua/Wz4afb1LB4txV1KfOuaSC2lbkfOC6to
NuurcVsyNdedXRplQoX3sCHj5Rev9YMVB8643eXRCPBfy+55DmQ18jxYtU1eVKh5
pudR3mjaTXbzzNPA+C7Ug/wa4Ke3QGkep1AY3egnzVZjxASe908HW9qoTN1tYTol
RdlxXst9dvpNLH1p6SoGDohzrYrYne/2SG4W7dhSaaBde1atM9njJrt0n5ZP43Au
kUSHgG5tB6OW7bI6sjK2HwIBdoCwAGgiWCJMuqBgTOAF+l9KymcMR7iPhTlHU8Fd
BN6OGcpaSGZB9QFT+2M3ykYuml/rOSqCsO4xsJ1qu2TgObFG4aKQyI2/a68VwPYE
InFWuQzgN/WVtyiqIHgNuoxCeTqqaB2ZRkSOgxEdw/SwKq04cLWHAwFEFSzMY9fT
C8nMMHn08Ba/mu/tTeIyYKJnV1RcDKRwR7mh4WR4Enyuqs02I6/FveCZJJObrv0G
dlV/JYrqQ1+VqFGtDHgZ5hPP/mFAL17BKHwhyWqXHmve+vo7EADepoez1z0TdGDr
X8gbLEg2IYet5iVOKC/EJI3TBjeQJ8gSRUzbaIbzaU/KupvuoxPzPUVxEdyW5lYz
mphS3bKcgcERo4mJI/L10y7Z6QF1JcL5wMs9fk+SSiSSWpKPtrRc93S1qdMxbH2B
Vt6yB9mmE5hE+aaiYFabBSV2l3D5aPIRBV9lj1x2MqZ5FTFVxazcaNuXRQ1d1Uzm
g8cX/F6TxkMjmbPQwAthw8NR7UHwNzEs4fKghkKa5dzjesUOWv5+RWojKLt4FMsx
FhJWDP4WMH2r0SK9ClPUT9K44ZIQyY8a81rHlk0tzkM5ajIFSW3LaQpQJzc6/sgh
HdY6D03D0Wb8a8AiNLtPk7EyMDuKjmH2UYO2HyJfCSdSbB5gwBV4ZdbXj9Zxs9pv
iBwQ38cWS4p2XQ/Zf2O2OY06GapnPf6Q6FtivFqA5jGQgHNvn6s6Mdds6frq81JF
SCa8ZFOzTXCWppI9ukpOJKiCh+3LsqRgomcAgArIrD9oJJOYxSkf6WMwAGb5m5yN
03hHbdbCp1wx69y/ms1jjxeioPBWhnjkVpt+zCorW9jQGM4mAAjBnN9ihi6cx80D
Ce7zw0WvwdZpJdpoLSYZnkh9kfjNdusLNJ6JK/l+pU/oAMtZ/JLwoopRx4dWYY4t
VpX98NlPAZcGkqcZ/ptos0eNuAjB3UuCdFxfjqkNNH91WVXAHay9+w8S67zKtK/q
qeS4+oBR703szu0lqCMJBCmJY7HX75xvEIAostu8jd3l2TrEBSVNoz6hy/DdEPfM
ulP1DyXLwhZhp90WP6WBWG/cSuV5io6QZE2B16ji3zwQL/tWo+lsJ2LHklk5SNkw
QyiXLVY5EWTBQzT8L9wKU/kb8PQaMS9hKdewOyadTPK0pcURb5q1L4hjCeEWux/I
Vp/D/5avnO6DPkm/QdxpCQ5yMfW7tlMfLSvwYpl8hP1J29MCAynGDPNXbqqgplvt
lJ5waMaHRDlFrN9Rh8LUpFOWxRcsSMAKj6Q72xgV0n5LG4GcAsQKjFPPfXm6r1mR
8Ja/UcKaC7IX4M/X5n62yXxj6BAXgJ/AFV6cgkiuRJMKxzs/sa/b50TnCXdUwR4c
bLMNRN4D4hl6yZcBAOP48Rkmx0AZALrXNaJPto/ky4vR5nzr5vyTDGflshZquztO
LvZvn71XwrK0+5qlkpvFaAF7/Gjtr39xSdo7X1LuvQu6gkt5JdG19oDiKuMYy575
WtYK+PChZqWAwsbKA5JvkB8xa0fa4L9f1EepeGEwaLERW6EAXu0omdSrPMrLdcLZ
+4YuVdJn8JEovdZlY6RSumTmnC4UdMQfy8QP6egrsQJJQH22sL1v9H200jVVj4qh
lFNuRw/3+4+g6uRLF6nKOH05qETcDGb0lmKCImaurEIVapnszd3TVLISH+GEFTS9
`protect END_PROTECTED
