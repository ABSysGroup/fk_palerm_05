`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v5hLAZbu3hszCwnxax48IgF0gy89NYPs72wYuhIVQg4J8GIKZsCdwAdF/xzYj/Nd
f7Lq/NKIZJ9lWCdM5bTlZkkV9UQng5g62uAIWV95CMwsXyAcwU/nz6LorPwFBZCx
rux+a//r4XuE8cTMGnKrpILovDeehpOome1blXUUJxVDUuj/p9Bm4qhAgp4WwnAg
ZZ395verNGiLrCTWITlO7cwMDTMePWelzE5tuyGFnv1vQI2kJfkpLj32H1f9ti9a
5cyP47e0qJ/rSJkkTNDTm3+FFAkpe0vCCoxFLbNA4xDaU6JqdpsPginLRPuZf8kV
4ajhu9p4+PGvlD8aM8XyoQ==
`protect END_PROTECTED
