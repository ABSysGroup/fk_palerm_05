`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V5TC0vIFJRqWAjHg77phnB6EAcwfC1OFg1etnMyq7/UEuGCDIzfJ4gMHRtvXSQLT
1/wKgofuHM9Jz4ngBkudd+iDcwpS45WUtsbnxVHhs4Z1vEwbvTa2zeVaw659adKo
ikzjsJ8+yiAjXP7tICPWhdiwbhgymazR6LsDEMdxc5X2iKNtWZ3qgyOKLhnmOzAM
DbamM6mdpaecX/Sm7tKCQp8YuFnJACWdO2AeOha6rC0cX+m2lUi5Ks2JtTMKb0+C
2hnRaruiQCfS+s8LyD7A3D8NMnl2IGYBw97EUTG21ei5U7ffrunCbGGwLoI/mA5V
VWKRd1a/UI5GV1L7yAi53V5VIQxNALSLlci8un7m+vcNfa4BnH7cxP+EMCry+XDT
sfMkGKVXLdRmvnOMG6oS5dsMGevKRhJU1YqjoM9gvMtEapRom1dxiyrQ/V5PsxDd
coFsCK4D6/wSM2QCQTVzfV+/1lbR4aNAyRaBMT3rZf9VhyCFq84NRiRPput2KV69
qInpzvwtGuEfxCjvNyMwEVyo7wn2z1P5PlgHBgOaTwSNyOauttAkBfIkYXFY0F15
e+3oMG/KYoqDBkkRQdoM/IxiKpgp+XV7BZaBjjwDsNnA7c/P/VQzvQHc/ltviXGf
GEz9Wcy19yXvyg2iPl0vxBhSud1l/QR0mGy5urhDGzjROE3bIGWeNLZO+yVuIXXi
5WTRcnHf5+9lN47rib5N9jd8utomgUnIMnEH53h3mmjepNrKRHDU6q1Q9NlR7Po2
ETbGZQsVqKQS0UbfQA/2pT5m0RP6GsATk7vofiSefm8BQadeyeztUa0kTT914OsJ
sRFuwVNqo/yaQV6gTfrvHzC2ZK7ZGOCu6LEqnKrfEns0iqsuFCzV+hec6vA17BHi
GvQER557WkbjUl5XOLiT8mIq+mHSIkNLEZ2vLPgAzR/bpqvIpYD/5jX5sS8d5Gjg
rCWQ+BbFrbN2w9q+dP1FI04K5309om0GSSjDFYgLs8piCy3QHffV8ud0Ic94bILf
FuKN3fg2Aqf43RyekAGEU6tERL8AY76xXyYBoNaIF+BSjmEzEtP1JrrtrQqWOgiK
12a/kOWY1WeMB/GL9TnHiWLXk5wzjh2x7+zMy9H/YHbQngasroPp2+ymxkClbXRY
54W7DWY0UFCIoQc/k1Bl88qjIIeTMOGd5vTbGo3YWWLNMjuJPu5xSkJbMxZxoLx4
8O/ovO/maPgDXzlRkJ30EGYBhrUSCIzLWioMEFQGCK406b0wFq3gfMF4y4ct24dQ
CmCtVFRBlLAiXbr7y7mkbMgNM5GbVmM+b0E6b7izGYw09VdWVeuaX5rSq8QaTMtT
IGMgAJQy0hV3h8WDbkfdImIHfYtqZdaHvNsglft7/8zRx8FNJqarS6aiV5BmqQLM
Wv64dBtG7jTMOI+6hx1gOl8VtC596/V8DzA/r2SSAGOxrjwZUmiIhJ09htN7Le/6
`protect END_PROTECTED
