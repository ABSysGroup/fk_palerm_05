`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TLpewn3dYjkupvQCijNj1O5BpqvC/04nnwiHYICTI+VTIz7ts7iCaigEF7sP6rYc
7VYy/5KdwLCXlDDqr+YW/uh+4+XH9JEgiVLJl4nFHt7+imYZb5vev6qiTZTXyrJq
WXtl8VV9m1jUgLnFss+TKvi8p0aS09e//gXvIzUkFr2i6GtQq6jMkgchHvDoDjDh
8lKX5v4ZjNztyPMHex2T9UhiCn28gRh57DmWb6OefaC0nT8Ny22F4h7KxNyzTtqp
0rp9AHEpIJO2n/PfPi/2sgmd/v9wauDVvaXB7V/BsVJus5iwAqx5fCV7hsAwppNU
lbS61LPL4PF7B1gMOy05WA==
`protect END_PROTECTED
