`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zzs8lNmkNV36CABeSxEaxTwULTd2UMDLYxH6VWPy39zoMbGFgy3RtjK8lsw/LhXD
Olkx/RrmryCTlZxgcg/7EcXb15ui/goEBlQK/2sb8bK3rCHiZL2YyMS0YDC7prDc
hCJqDHeqcnbB+4lwwYbZ9/obcCc5Hl69c588bVhjW5ItrmyK29Mjv1yt6OgUm5s+
/Yn8e1jfgBdOZngzFdSURSHWZN7/+hcZMgVmZkXU1agBXNUL7NsLgzNOgbOtLlIy
EUcq+cPrXsDdC079Xby1xNEoHwiM+gMw5CxfVyMkrM6s8rEKQUSApkd+rsSyAhgJ
8tMKO+szUMmklKu3fWRCIJ9wsCg0f0320gqP4ON56DJbERopv6vyhZpGETaJWb5B
3JihS0ikOOyDijRaog/2TIT1MvF/AnEA2neJgrSG2DUqyPhRvH052YfHGy4klMXY
S6Kqcpl4kAtpvtGc47V7owfWeA1TL9XfxiYE08p1zExl+yikRe8iDDp6lqLdUgZs
2McR2Ph2JFK/wlfCRfwh+2XzwRsI/EcNZqBs0dNiERijvxGamWWU4qDxP0r+CmSm
UaEkTBrln6VqWt0TYtehH64KItdD5pFpskWS4m7Z4copstWF9tzESvyp32iu/yat
vYuPE7aJM7DWSSRK05VSohPFOMtA4lsN70M3RSZ89IoYFow9faD6ssnJ5G7FeAmo
I7hoeC/z6/MRLV+UxsZ8JjcGVtnu3ZOLB1hq7QMfvdKPU1WoiJNNXU7HDAcUBAWg
ePQvkgjY6nvhab41AtpUM+k3tOkbxM5Wix/FGYs46YWkw9e0CJ7+qSLe6plm2zv3
q+mBvBeQ48zkG8CAkECeVbAGnekuPmKWkXOhkPCE9qFGfJnuVIZDAcgBchTaNjHc
ZRJD66KDEAypk1lPDyoDma1bbh1qD76+udZ/2NCoV8PQTzzZsgrcQMYwyoWvGg+y
vBEZIgKiwmtZudvvJS7gHkMkvH3wSn1GAZlmAB4x1HrMqEuvyQfyauqBHtRZDu+n
v9kjC2P2UWB92AdryETv96hmNwKvVNyvkOgUjgeGj2hUgh8wSMkI/vS5+31ZA6W0
2okHoySoCgmaxZ/6cMY6s6YWd4FOx+fNU8engH9dD0pXBZpoFuvQc7MN/jGJ4qc0
szPHYSri9X9IMtP5IVauPcJkCPz9+qfhfWQ2y++pqp9ticqeIerZEpwngjaOkbG0
S0/+U1LF8VA458KdCp/SmQ==
`protect END_PROTECTED
