`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RN3rK+30ktClDPl14GRvhVOYCzid3cMCCwqU8cL32ohT/CudIegYc//PBuM7eNX+
E1G6KriBLWTKO4tLXgo4h4ofijMWHQOMY24waFfbjVUloHekMBtrSfBHpAxppkEA
UBCPjKUzqnXLztZcaq8WI5Q5piCPzvW/mvDmnqVjHg5NU3uSuOywdLshUJvpQTuU
0X2xHicUah9jfrNaLD9j5VVjFGt7AaR/u/8T76IpC92QiUP5tOHo29N3g3RjRdQT
PbAwkY7tGUY89F8yq/5JbBn2fU+CfHL8QjEc0ij28js7mC5ZfeIakL8cwkrFqU5U
vtzaOsK1wPeD6Do9E7hOnXKNmp/1CJHiEKmLHvC+0cpQFJMqyt8vYD0D7wPeu8ot
DhuV9TyuPwtjdQ4nI4u6XTzvQgz4IOqptAiwsBUA2i6XUwVGsjExPtCX1Cw/kTKW
`protect END_PROTECTED
