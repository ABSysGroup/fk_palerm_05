`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VABmW08vXfJ381savH3qMIeJ+sFLELp2veOz7arlLCS7/J5l4sHF878op6BNcZT3
+iuZEFYl7oy6m697AZg07Wh3+l7QUGpJp3uchTcytlVHNPunIGJhKY537ZDe70cD
UrlmdsVhIdyFfa6I2EDiYB1zoJI2OsPCYL8SQCLHaJI7QEKtbOwP+ry6xZ+Wymp+
IVr03aQI5kZOEyFhobwGPutrgz7a9nBfRmfjc0YL5RgBTSFpZ4kYzZQ1qB2sTfHM
ORgEhbr8j8Na4QspNKG4MI1FL+k9MXtYk7zQdFVml/pItLJW9FaqrqOEG6A8vDXq
uPN4Y28dIwHbDqfI8tUpunVlgfXTZX7jhUH9cjt/EwAuNMUSMQKw0rc3/QV5HFfb
23OmO9Yxvj++uAjZ0258Crb2GmXPj0eYeXAoVye288XCLOA+kHkcTO1mamt8K9xr
En7LyxndUDbnKZG2Mmu1W5f8minn7/7sHNQltZl27IYv4dmgOlJd4FwuMbtqPgjV
oa4rrgBVQ8QEnBiWatpVcjw5rqZcoEEir0y/ic1hyZ4=
`protect END_PROTECTED
