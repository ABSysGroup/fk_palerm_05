`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nOVCUCRGQAN6mmzR1NpckJl3gX5n7ekoGfkeBSSLajwTZeDRp/ueOkPNAwc/JlVS
hORK2DA3YgJN8SgqkOErSpcffBVSR0eX57iHgBzmbDCVTrmih/LQvEyddizoTwIo
DBwSkYIquVF79LnoV2jW4265etu24QZtvp5fMf/EYciZyS4bQUnb2Q88gjF/p1YM
rf83t7DBbegtMFxdmX5PE+F3S3t1P2J2zrubm8WbOYJBR3FZ/LUkRe9M0OxuHkmB
gFQXyOi9Uc2wjYzy41KKZoe5V+70Sl2W84imiTKm9qDnhhwphStbdmrYHlkGty3o
TNTsefJ/tiXU1VShoUkBjA==
`protect END_PROTECTED
