`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yX6mxOCmkymaGvE+K+7srAsLCHhc9ZLpwFHwBZsM3gRpVK6BObINazNlJoQpq9BQ
6LPsq6OGmK56cHHZVTv31gtniyzrpMGV2Ay5Ee3wvSNvtCkSlfjZ9z06SwsonOtd
Pg+/oD1xmiMXinwuY6FG2vMa88yTAAjYX/ok3MmhzH0pC+5oLFRc7xdl2WXUloJM
IDW6KcU26XpLWDjwHMv+ftRcRMTGWW8FNGwEEj4juwTTS8j/f7jNYhHnsoMyn7rd
Mf0urClqWaqhKPYjCC9VT0C+SidTyrJnt4VlbRWyglFTAJE2NVQfq7Dn/Knz+oVD
b/2B/MWkcisUCtq64KPY2M15LFMspx5eIHspB8NS60A=
`protect END_PROTECTED
