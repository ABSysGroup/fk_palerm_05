`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OWjaSDjRYNE0IwcnRsH5KU1efNM7RDmqDQgpYgH+i01204MK1zuwTPBZ0kNgGVu/
8ky5puKty765wG0UvomIfkLE3/w4qXDaeQCbeyZ6SMvq59CD2gAVbAx9bMTlBmB5
MlPzxiG4/LRaf1CnHWcJi0dnp0nhDOwbX+GmnsyTlJk3NWXs4VDGcGQJPBaz+HPN
EbhsKzmVQDstgLb/TeRcyaqV27zdFCTqkCNmDfLvcnbJvHGGObx0tR2Jjx06RS3E
aLzzRsyAcNx7/+yDgqal9gmagwkRHQTaHJzUFzZ3n2g08ioysyZZG35aRK6B3T21
fwT/vam/oq5a7xko6hihrqQcLKKvl9bNREzAfgT6GxVHKLTB11evdQ6sClupeung
oMK8WpZD0SFj+m2c8fGalw==
`protect END_PROTECTED
