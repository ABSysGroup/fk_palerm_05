`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ju56BRVDNhd8t8ph829PzM6uPbB5J6zuU96tYjmPo2q5ORXrn+lQCvf3q8VQKdcW
JkXk9m6dw81NWEhsTC9Z3V915MHjhk/HED/305aoyRjIaQnPNHqZ33bAQPiBgK7e
ltRwdkO6LwepKBuEXRwL8GR/pKzAujueOK2bOhNirvWlGPEgoducTS5Sf1Dw0YpV
pYfmkrqbhdFsNqMT30WFlcnDPjBZUjb0IEKv4oVvr5BLaC8Q+6h0nCxPMwFB01tj
VpLff0iJPfTX/N2tOIkAmuODxsyHTvyaNIsZHBky8RgHFHEHvXbXG4rGT8y3ZQe+
1RMTbrOO7ho7SWD69KzVxxdQ0yI22bd6I3WlJwdUD0vJj6bjIRJ75d31fGyuOU79
XvrM+g5K+Ydeiht5kRPiQVtQE9k2JND0W103Mvo16NM=
`protect END_PROTECTED
