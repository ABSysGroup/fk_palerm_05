`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kofTSBXQ5oCcZ1avpICyraQb9iA1NbfC/RfjFMmoWaOwkuuFbtbyqPD/fQGotxRJ
o5j1WH23KNCeTU0F/OyrNoZ8mekIMIyNhSoYNA8ZQewylhaxD4miPXJSizU+8nOX
DY8R5J722RthTWPvG8S1ATrr3xmXrnaf0CzUba+EBSCyOfCO0zSuvufgEmmhigIQ
Zcqs9tmv90kgz4h6hbjoHEjJE9CbQWQjPSWFQN3gU4gxgXSRJEo0tUFmWYmUUasE
kn3N+eRUubm+wWBZnnUPJXEB5a1wuHDPTDFdneFXZDwZa96pFZmZg++nmHyNZBSr
sOc6nSs/9XZ8qo2WcPlNCZOKjtP8dtf6DVBUm+Ew9ifXHuCnG+df4pNfZqKEsBpC
2iq/KSP4um3AWRFR7bkmWS1TeyuYJGzEU7n16enEb5AH1zgYtcTs7L/jt5jE/6Wl
VZ8FPwEqK624PlTogKnJ05z7k4pm+2I2X7lRs6gun3m/n8+aQ/qjCmnYBXNl6+yj
meZ6wsYA47MnriPg4Xz/Wsd6zN9I+9AEzmjIP0tyT7iTcFGwy3p67UGzxjB5QSr6
nXfacFSScUHMjC5DvG7ss2jtwOk1t8tKyDB0NAJjKl8xp6AsSuBd6Hc4ro3DN3jy
M4BiDs021eIXJKPR038jOQ==
`protect END_PROTECTED
