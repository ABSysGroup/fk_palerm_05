`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b6j/EufB81QeiQySnxMQycnVcO1vklXMYRDrGpB2j67XMPL3rLY+Fe0nJ6tVr7l3
kLTFMPY7hhSjD0AtZ0TLiC+dyQoVL42fh3QLnkiebay/UPoSOz7m98tYIspJPoLn
5xDi7bm+47cO0JFkSuWqsVYGRtnLK6jmP7a66X57gwTNjh9XW0hv9zq/ogcUcsoR
Xxmgy+sk94J17xMLe2WERl7jJFCZB32hcHvOndNfqtMg/cpFwSEuClsYgyKrHdqE
RDEuXeIyzLa2EcnO8W0jvLxGEDxz+MojeGBBBq2C0VDYCdlWhta7D8g8WBqCxhyR
DDXkKeY0YbkqJLNS4BcvIhRdwfK79UTlUUQdt0G4CsS6I0IejvyCQLTRSliO7p4d
SzK3zbGCUAnNNTEGqyGD++Cpu82MJCJbfeV9kTGi+LiMZO4tnIvBjd20bEFuSK1N
`protect END_PROTECTED
