`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uj3PdjOcvwa9EWxQpYz0k2aQHF6cXTwA9PmVVoMBuxoXM14a2baTBobKo5FWLCoy
7ikwxas9noMYZXtoNUe8z4fs0c9MpCNOj6BGJ8cbsttGDVsCSUqxgLjwSiirSylI
p76IBBQvTtjXNht6TRlXt7zasdysJJuIEtma/d02CYqAj6vr3vHD4IbUJTR42tlg
tcdlz5j0+V4ouoQa3vvKFqMQAw/d5eZWhrFQ7U6POYyfdn2ljRH5oJ9xPXtTRM2s
Z5VcGNDoulNofyehOl28HUsvtmTd/d2eP1npOubI2Q4HOoW6G+bgxJhjE7h+ycDW
9+AdOxCPAQk+sfH6O0UvJA==
`protect END_PROTECTED
