`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Fp109u4T+Umn2704hrklGYTiTSNvn/Hr/nyz2iTXNuwS2aIsqqkSSBBVCwWpRQe
RLau38Y0hnq/Wd5mydelmoUWk70kZ9GWsxnNTOOyj3RKJPfb6Zhdfrl71nLCprLF
c3ady+N8niBj5qZokWUgp9M/imG/sMnfBLumi8QYLtsLX7jq8cmOrXGzzYXohRZz
fzPsBF6sTqJQZnL/38puM2bjeiHVpQ7mAjHKsOtWgZJlJ/rSa30C+Gueyt8RJyDT
STej/q/jiOPX3BLi7ThfiAMpm5HXpSqDoMrdy1lUq4VEfQt0M7gQrZoKVY1Vc/tJ
MZbcrk2UaUi5ffB8xI6fLFbuTd7RVdqysI9BqyM/CAXkl6sV+XbO3WILSFXxoaq2
Ta3O4R5uSS9nvG7nI0wEL3wegGN3E0P8uKd01mrvoEA=
`protect END_PROTECTED
