`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zemxkMmoznPF6s125JDEXv49FMRlXCIMwyEa4KKRswz8c63VxvDp9SsA8fYUPBYk
UXM0SyE61j0UIMAZ/XyOSdyw+jxfcSDSHAB9k1F1ANLGWs6Bsr41nXJi+aEL+2Oo
54mviA922AuiueioMqvp5daM3k4Qf6vfXjwS9Ph+4ji6RUJ8Ge4Exely2xBj4Nw7
uAmW3MnJwdj3F9XVTd1qPDQy2tblhoCt+qyWNVgyFBxFysCOzDLbAedy5Xqpwc7O
dU5x+/IUKnNeBZWKj5FqcjGX8+RCeTSSgngBfvp0G0zdv+9SxUAd4W0cmjrDaYqB
5LOvT3tQuemF8WPvsZ+1/ILE+ov0bCh+IH/QiU1HSB+8FVNBi1dB5w3KCUd4mL7C
I7aRYtXqxWYGu8h+EVbLih07zkA3mFr8GRxPFyNIbTzNnNo/bqprxwA6jxuaubYX
ADTMftGEizkWnPAiMjb7ZXw5N/FxI3W/vF3OcRWZ13wnYzMF6bko0ekhQ9qNzAa+
8aO7xEz6hNw8kwdH5KguGBL9Cie1TVBecr9bE9gI5obemjTeJty6d66hB21HN67W
GMGWoJV4H+ks2FPLHnzKRGOGVRCJcf0/t10l3AssbrGcVznZaztQb9wRzEeu0rRx
vs6FzD2EIOC6cLhOWb6lgJbpBHUeuBBTdIRuGFGC4xsOyfDkpYH/a1Q9pUpiyMHB
F9W47AFqfms+O74+JkK2IE6/OL5iSzsuEYLR3W50YhW7z36V17Pxwjb1u7gqAC3G
4jlfUQYCoZA3orVnYGgh6TA/yagyBCQNgw3pXniLrO2mYzuR1gIeAAQw2SD+DQW7
LgdbI2dREburV1EeTQ4oaWZSAHGbwuM3cnPlWbdT3WfW20LnMGDHAMRdn7GISwIB
HxnHEGaiIUOHkc+bKxzddyELab95Qf5TjacZHVcLjQgmpF+naWQOLsvLk2QqcV5C
VvS9yPWooZnOleNdGUZT/2fInujLZqpRJlOGzfablp8q5hV/DS7E5jKlPeXBEcrC
`protect END_PROTECTED
