`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q+tx1Rx8sA4wTBtyzIEcfD0S8IXr1SuSUrBnGwkUQxedOH+oNP1ZwlpNgw82e03e
uDbhyzkhqkIQk4ANuu59C6ogijMWRf3Zcs9Z5nz0LgkpazJoLs9qyn2LhAg7NeZk
ryBUpcUxVgEVyRk07aleTp8JhkGI+G/XJImu4E3zyW+p5TTeNY0owB1qjYwlkah5
fqDfvyYudbHaRiAAhjpFOgLfl/mOe/iYstsOyILAM0RCC8iKQQMht0N42r+ffJRv
yIevAsTmKJupRzqyIl1ugIiklSp8b0zIRZxyEA8UPbkVXYoSBxrFzzG4VSEXsCGO
AXl48IbCKFIsvnXAl/mbyw==
`protect END_PROTECTED
