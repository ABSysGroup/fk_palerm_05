`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ry6wovXavOCni5iGIZSSIyxxdH6fsBPWHLfkg2JW0Mg2uIasBbaniWnZoRp6aRd6
kBeoXwj0Pud4jq0CQ9TIIPzWH/7qBHX2+fMMjp+TIcJErmI2pder+NADuha7GhAz
VuX6xNKqcBReg6qrdiHYJfPe28dyWFNJjZwXI729OrphFny6NaTBb6E2Rj/zcwBU
MD6ZLE2ifn9eP6+HpvBaJ+PUDqa7vf76jvfplsoxs7NeRp1soJT3h9U4cgnatfAK
HWNEYjj6X7dJvvhEqsWQKFnHlQ4TRpxYSz/fVAzqE/hHvdBAce7iWs3Uyuqhy8GV
ld3vHCwjBzSx13219pMDPYhb7I2qxHELs78m9H5gWIHEuTFhTYxbKQsZhlpVFc+L
evYW7YTmjXzL10vaTcZI/KM6wJCUB0KBcPTd59MbQ7/WHgZhF+AzhnnMXy633YoO
0gXO9EaPB9ySW4M9Vm30iwh1ZjEjFXLTUUZCXk/ER9LEPHK80dGbc+3K8FYt0T99
jYczFOWPbyeeVukfUhX+jgCJoP5KXPYuKUMqj8pVhPmn2ckDWVpcGUlnyH3Z3HEx
eNKtpMR9tnMBB4OKXgYS6uoUO6xsikZU82uVu5idOvWPeFDbxSlHa59aUUPLj2JV
SIK5SEZY5350+15b2e8oxCN3Q0YPFpGinGxrSomcDeSdbmJ4SlMdiWmkM0uW5wSR
KJnsE1UYtaGYiCDSGmPRc6dU4rB3fkWD2gko3VzuXnG40DhaMlbCBMzzBApOZoY8
SqC0/SXrsuDYuhTsEB4Hb45xdpS6xP+/55t85Kjq6Cr7RmdNnMo+yFWX1OYNL8AV
xKquP7+EtfJmnCp62Wn5yo/iY7mlAEU7wTpVS+noB/5hl3kSbCKOuO6j4+S3co3i
JK9UaOvV1TvwZgtzfA0p5csobsp/twel7s/KTGUtvvVrvC30xCFWwlN9JHviSXwn
i3W4m2YrMzYS0Kn7ZaWu3pyNxKwfZnSywBcPzZ7qrWHNTfB8SyyWrdFCUCMZXuAd
gnj4Ix3xJoWqMj4oMpgGas30b6BDgPm17NgfDj9QT0v6+//PBM1iOAutlLATsmur
+K0destIAXHtch3U4wExzo4mST+zKY5cenq+62ZHVvu030j0xTVPeIHLHoQ7+2eI
d5ZOoItuz/71V7L19Ov/ZSUxzGPzK5j1CX3SEO06FfQRiJJ5qOrrf9yys8KrRGzg
ruduYOiDdCephijGtJ44BM23hRiCBI2QzC0U3a+2QktWkITSrLk1JJYBMnavPSix
2Bd8vkWFWUkOQIX+d40dJ4NjJxvM3+WitnWQFcrYCvOALssgtfgckiiFoD5xMaTW
zRDeExvweMbCCXK12veVE1wDKZDcIGpBe4aeNVkdewmiZZjmlTNAtaqCLg8GmMbk
jsM+3mbrZWS0mNuf+WXdEqNcxanJ6HQszBXkGtuItWsSBDrUBqD1rb0YpQQp2JLs
+7flVzOK4J0ld3nykH8CaKYJKU6oQSjkaFtwcvNphdfI5Ny7uBuAsHZ98Im9PweV
QekTHOjp98Ctyvp6MSjQp1XamKvBa73NmAMCe5IDBiZBYk040PGOGaBWmwW/dlA1
KFrG0ivmDmkOlVkSPABEG5AK31nGnnG90Jt6++NXnyI9u/xa0eC61cioHIrHi1x3
wGCybG907CWedZ4cAER9w1IljhLvQIDUF4TESwUA7k1G+2S6y9jf13Tysjc16ML+
um6qgMVa5Vb7OilQrPj4uxCoaHkaDrzi83p5nhR9hjnIBQvccDeRYcvVFy/cHWdg
/T/hH6G0uSHh3pDw4Uz369cjNYeH+sT8yavRx14TO0awZOPNAIqVID1OfXBnEZFK
wSY7dnHHnkpPPejiyzY95aKc0YE1xDg+gU4MLoTdXsHO2CeyZ3LyjpYbxoFFtUrc
zqgtrousGp2ApKSoR6l79Va3tQ07ceaSVpshMYI005PqjH06p37BST1UwIDM8tr8
2gRQcjiejg+O5PZ8T/SFHy9BPW0xT0HOpZ3bcPizNGIU1yQy+c2VleUjLGcGsGhM
mexVbnds+V3IXdbGIqwMP5alDjacfbBmHj9EdKwCnGVhOKL5XyvLWevq6zkRJlsM
RTtJn4QB9nuIVmkzHPvk4YdAI2PvIJfYi9m8qccDYooy34Z3pNflU1rqBUJuEi0i
hBTeoPwaqyAYpS+gGOYnPVbbOT1/X4DekXq3bdgyPcmuyEuTqi9LcS8Ns04f3IBB
iWsOLZMoRJA1WsRfGRpDw70cGIeqKZLYPRFYrmnkkfSTJko3HV+IkwOGbdkQ6fDE
zxpJ0PfJCPBGeuooRc1H861qdJB+WaXm7D9gxhl4t50pnf6SeSEWZVV3U+srieOj
1CZH+q0vnymTLk0/ItR3D6Bar31cgC7goA1XqFIS7fjOyyzH7Wes4Rfe/P74Y4Hm
C/l7I4jWS9CJlNBKPzTfd+ymuc4FdhloOTk4tdODztynh5+k/HsDdHzwBgqSvoz/
yJBYwwzm8VLEZF6TCBwxWs+27wHqyvE9s8OEAPInH0ZBVt30Nb9Dz7UTSn1di8lH
b0sOOBk3VcWNBLP5gWm/Z9M0FdUinnEb0VoJaVkoB2aJ2syVHU2JTxAw1hxMe1C9
3w/0SwygsuEMmgFQ39kp1/+8l+ekVBZDvrFU0xgwEQwTOuTAMqYx9hKMajN7tAtz
1esiJXGuCnEilSotcar8ijBxDxVWhidPmPVr5vega6YFsliItSyIbcWNi5+uQmBQ
HkfEsit+FBUAP9ohhd8ejWSmzn4Ln7mid3Vt2BqxBxG4iiQd10nZsVislqnqAtj4
uTMVLtdZWWPzIIJC3uO8+fKE8R1x4m5P7cdpnl5Gf5a2FNGWl1F7rJP//Bgjbjr0
cy8FjV26T/BHPVMiUCCsZVmatj92YFgGvtb3Zb4gwpm1NEaQaSAczj081qmIPvfU
HwMD87WmjvBkgBzg2aE6ZaoSkGxNqeOhd+7KD0CbN/VGrbWf1b81RVsZESq2JAz0
YVfIj23EOACoz42WEtVlpMxerlAuSLXOu8yvO5a3ZyIG25YzTe26acoMXSmvXsLy
rqkkDY8E1LP4/CBpVbjDTJ72NXzWGxtq9PhCwOY49cXCLpAgtaus5iE8wmoqd+Fi
c//htgs4pn6R+Qi8ACgwI2hGTiCkwmLeniHBy3PgA3wJT0uuGh8Zrw48ngpzuaBL
2dglTwj1Fa1gei3xotOznH50ND2x332Z5rcGEO9dTp4=
`protect END_PROTECTED
