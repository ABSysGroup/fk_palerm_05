`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vck8PvuLpA4wnY+ZFwIyiGiA8QSg9jwovscqWaOGjrtDzpW8NsQDQwYLFnLqFthj
vIlgTt5AoQTVIG75z4QK2egjsx1UBpnKkIe28PHQVEDVLn4uZvjrfVQTQInxCEP5
O3QyNxK5pai69hmW2qdctOO3Cg4lEw4KC25+pd4OkJMt0is/J1eFqdcM8PQjCTSq
MKes1RmTHyj8zbQQoquXVpLUHAvFfjPwaBa6CvjLxrV+eXdv1kwWEA4k9s7655Go
znYSQJ/66O24WgOD8BCdfCD0QUSmdUJxrO5RjoKyeH3xnxsmQ1hCAHpUdbzoOj87
QLefaU+RTlGusq5nqrAP8w==
`protect END_PROTECTED
