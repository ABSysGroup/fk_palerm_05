`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qQZPqrs65Nnz0OMFErRUq6FbRA4uhpoabPG5bs67fxZySvNKTfiHqGY+wNbi3LTu
/niamyPazN/L0zPeTlg/AGDleZ49cf5as/KMEt4xOhRWiG804PWREq2Yez5m0bTJ
Au41BM7ZssSXlblq82J+yZNhv7evpvGl73F2mTWnSRKUXwNWPn85dm6FmJrh60Vj
lDD1aSH+86jSkgn64Fht1qkEXvZSEl1n6L3Qc4+unZvzDMl2AIuGdxEAIrnItY1W
/VEhbHnS98b8+h3Qo4JP6xxrt+ycBkTmmaBK54x0uvbrv/BVFMO51a9Wcc7x9W4V
9/VqgV1lKniG2DO7ulL80jRo2742TYbHikHcKBuXGKgWMZdZxvBRVA5SVtaKQXKe
HaTU4hYihYfZjsL3FvA+WIimmada7QakFVj6H4GRB3aRbZ0yYqdYNkKhJ/nBUxkv
jvxlmqvLMNa/BYpUJzix0nfllQgoNC5tSb/A5Vj+pZvPyDEOzGVdR7Q39C/CJ1DH
q4cXzgrx72b49qksmH6eEsKNOAIqiYFq8VG8eEvFnvMiiD4zZbkTTAkSJl6r/CbQ
FyrAKLyXwZV2CvnwoWH3tuWX/7TqVMdPGXc/SG5u7/xxyyTcuUwnSsVmSdQPSbGi
VOP0Ga5jOHsIcuSL5f/d8UKwDsHkZe3lXVmC9Epce5upvAgFjQBaKhUzzvR5kOio
nhiFlY7Bj+7exfhfzc/WzyzHimEHIB1StzuAGDuLIXs9x+0YWhjUf8fEVT7r5RBZ
kOTzV3sQTag8GPrttCH4vHo0QA3CXzjmadhclfuX5IO+dPv5GakGENGm4wSJQHOv
EwDvABMRzaIlnqqYYZHwtYpCI3d4F/wjnQ8C6hkIf9AKx1F7LnWJlJE/VnqP5Qi/
ZTU6Bgc1AGGKw8nfHix8pe+NcNAwhsjMsn5vgEKJ4kbOD48fn2f2wTuKNAEL3zoK
BXaWtwpU3q7Ew+8mi/ZBVeic5YbGP0Kd7qAUp4UMArURy8Xqc7QWUwZIy6L6USfF
wPIBoc+JWb2IwkUoifOIqlkWA1GSvXRQkHOWXVDqzAey4GUSwdVFmjWeEN43yuMz
DAb/BKD8neNSp43IrkwjCZ0vnECAShZQdbFAfLYrNL4o4OnSfSCzmG3KHDnWMDp/
5FmBhMUYcsKSkJeBualjpMBlqbFU89993fcC2SOAN2FLbPT6o4za2DqUmjALnKwW
cUzPZB659aGNXiwrp9e3KgJx04ycMlXnRD83XOdibylGMAHkr8iGpsRGk5Ktc9Yg
0TmzRMaVfzd4sC4smaQWdhRGet7zNqQhfYsO1eqBgdEW173i55PbPsPGqJT/gYbh
i5rUd3+f0Yj9vOodSmIZCIBKqwfq4SEtvh9JHS66H5Jr7qtgjZ3HDfYHWYMBUl0q
q6pn2lIBNbfEGmdHiFqFXRybPiXFUS6tFx3DmG4s8TOP2A9AvoRkIFWiPokff1pa
4cZ2vd8qw4Yqbfp87vQY2tT2wkrgxaw1zr+WFNTADQPrKbrv8QX8s8UYAyMhudEk
BklgZSgcY+Sb1DQI8Rcd4JVwqNKrz8NZnqx/k169cf4TFKTQaFMb9nLJmOxCHLGk
UQh1wUJjsFN7cxYbe9ntyj7M7cXs2KTVlYSNqnPbHemSwDl8wudeg91wm4PwsNv9
Cuk1Zu1CXfG8pv0yU+gJF1O0gix7tGo05P6FpyJe+BSdf2utflGZTxOygm0IhKRz
dVNYQZ1ERhzwP6800C/DKRlK+Z8s0EGKfP+EDzP1kNIUpB3Vr+Sqdc/scBhre0SP
56vsd26LP0gOzDggxZlIS+Jlhn3yT+7HkD+i8AkO2TflSwSZAafnQHZoDh3IMq2G
xLtWhF6L1TaIYiFeKFiqhwvq+KlUZcoyUNugeREjVEqJ3Bow3+ga2j28rA2za2Ch
6t6KNd4zQ17IhrkoYOgvb6zqgfzE62Pu1xGTEEU2TvHTEBkL0ljEKRJmbPyyqazW
QD+L0VnrTCPxwgKXj/81WOHuycJka9k66cx3hrIlo1PqwzBa+0dcdsB51O4l1+ym
k9JNwCyxehqX76pjOC7Y6QTS7oBAismOzzWIjBEFDgUjrg2mMb1IT2TeokzxNq3A
SkdaaeftsrD/oBQYNj0i3h8k2E+U7N/HnGvcrTxAF0/GAd/2IesRXgv0PfCZhfi2
u8pFNU1ZycPGwDU1nThLPiKPwk/GLoGWbZsgzQIrwyF0re8J3p04me1hIjoeg8FL
KNBeww6Z7pn/97zMyNZ3gPYkVUITL/a2FC6dMyqOvVmZd/cND4BdblDNLmJPOsJq
dni1r1bhAK4zvjk8c4dHYQLwXxCnEyro0t8DrurBW8bOH/YSVCeUGZGXH05Oxjnx
Z9ndpaiPouQPm+jmziEPneu3wzyfA66IdhtAYDqMwnh5M8JnKlQ5vxGTITFojqOF
azXpuT4fP29bQUEnRXR8ZxMMxBRu6EinE4BJFcZ0+FkGVnOr4PY0IJZ3JAKd0I5M
M7O54Zi6v9+oICU1R/VRilRfehXHsmkow/6XwuYV4LgRQvy13r0y3MDNo1efY+zk
l0u7h8xFIdjQTsC5ZIfU2sZFlhDuJPwIEz4rVPIgl7rmffT7yN9wjMr8jQGca4qv
l4a9ggkz8iAJdZKzy01NeGZ2MfDCpd+G+8X61aLZBYldyvOv0tICH5N3UzgAdQAi
OwpVJi9q/IYqndIlgAoS8CiXpD2GGRIP+kXUSs1whOwFtW3/ZnFe/bE8rw61YFA5
bA2Ckoo7n3zJU7Gjg2+h+21ZhKf+zk8rozjy5ELeD75kHzJOZJGyL/g6inEninEb
wfYyMDaqTpGRZPeyThutS7E+fsIBfKzbZY6+pJTpoJR85hxoFq+/n3Z4CWeTN0Mp
`protect END_PROTECTED
