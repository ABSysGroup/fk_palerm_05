`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v6tDfXVaWoQkFAmkQw02x4Ax1AuaDsh669NKRZmFw9IOQHDgc/DfgNvJY4MS6Y2q
2olg6fN21/a9Nc2TTqdgjJqv9yDhcP35D1y9zmYkceMkaTHd1azvUi7GRlJ6Mu8Z
rwsbn428kbjlRQOB/0y9XjjpsphWo+H4x5bDgGZLkyioQGOg91k6n6Nkw0kR34R5
EmyCbpHjcGUW2AYlIkdB6+GdzSfm28ggC7lEKI2OFGj4YBhUvMxiP91NCQMUsuAn
L93+6ldTGdr3IrdhGvJJ0ei0gS6wHjIBl0MnQeJ3fjVYUqy/C2RB3GHHGYdBvfw7
Euyj6Fdq6npLgwhs4NHqRRoUGzUerhHf0NwomFlKc1wJEL3/im5SGJ2BidkbOqKO
i4YhBYqRkFMJHGQzZx41jOoeubQDRBzdo0CRig3TxFbKVnmruZ9A5nAT60SYIXEa
ElKQNovOnM9qqf7qGeF623FCsZ1r1aNIBgYSUFCEHhIbZ9OrSXsvvo+cgj+NL2h/
O/oK52nPEbUei7EsOOC/9z/By6+kA/uFM2Kbvwwlm6kEJ8D76JF7ocfKZQvmFGtv
jhhNiCSTEGV/agIWeImYuLUf0yV21uf7tiZcgA8EhwMd0ti/stb/0n3yuzPOVpJ1
flqCoymdlYaY3yZslurN5uzFEuCzlMLtJzUqU+ois/E6gVNEPdK3ZWOzme3LMEWU
U3tmLmSDF2AY8walGbnMlpSYGhwlGE2jKUNoU9C+l5+lh4e+6FwCQEQEmAnVOosn
ew69H2tQT2InJFhCBfHcwc6AmyGixtVIjjyN4Eow3qE5OAafbra1Tb7GVLCZr0op
hcoMmUyt+bZcps5OoH34yG3Czr1bv5XDv9pFgbyfLrc6f6OjZGFWq90ucMiCCazN
H6+zgDgKrtsJRae1bVb0bXoLV/dg2IMVk608qiyYjlFU8QzWhpzXjlU02PyQTWn2
k+YEjyfP7A4bSvLo1Pe9XDH5ItYYKrGy5OJy8hDAP/3CExwe9PX3PGziSYrrhOgB
e52+gyoLcC5dyzvaa98ACxVDfOoWgQUz5aP7xh5N60myJhBJ7bB6rYT0fQSohqGG
q3si9hCJhbY7FJO1b4nlsLYqy0soJiGJBeqjYzV+/nUmoCVnqhNbkDao2UNEbUQ/
SkHfi50WvGdwlFSzk1DRmE2nxw62HmcLMTrPpdWk+6Hnf1r/y9OlN+oZdGvzqb4n
sVyi/J7bzao9JGZVQk/0FVL8746OT61myrOmQWddyiLukxwHqnSBxCmE5oxL+QmN
uzHckuRCQ5c0uN8kwO0lOtSYh9+c2GzTvm5vL5ocKTcVn/eosbQ8/c/hb25y9t1l
ENprVEhEda5Exk3WRpoWP6DotoVSbeUQAXy9rwJa7Jnu1DCYlgmaDYzIcSq5q6j5
e1rmmWXSDhyZ7UNCMFSKsK/tpblnyymHHHPvrlFO8F/Gj6cdLFZVf2O2HskwB71F
NGKW9QPYzpk9o3CE9utKSpP4pxzH7JpJfeWvV/GfgejUuC7P/IhRzfZwaQ0equ58
7eOc7WHJK7yStNqEbbYptu30c/IBbe2jnKiqI8Bq2d0xcmXBf3iMBpJqBmBtPf+7
kI0+zRNVLF5Dy6/q0KVv6RirFfxUb5mubGebEOeBROLIV2HQX150OmilVUx0xTZZ
xhz3/eM8DtCagdCs3xlpM6R4v3b1NY+Vvlq8La/YOmDuTSraRut386mPt0XLGwVz
BjWWtgEotFPAO93Qy/dfYbMXvtE7vBm/RsfyggE2GUsWpmIYt9Kmu/E+ajLTk16H
6VS7xGVc+B/WFaQPmPzKjQJy/Yd1s0yaWzJRYh91kr6fYKqrBDSjDs2rFB+4/wCy
w+tIGnf6DZuEZRC9IxvBViCeTPWiitMJum1DuwY1nlaD5nBr513vesNwnyM1J/Pg
YfT0zM01fk5QFBejjqzci1HLzGcEDUsqVaJTu3gKqMVhEGPJaJda0bIWT+YjAwGM
xRuD3U7u+oBMSNfRmlhkBdrwTDLJtb5b1BTLgBPdF7aK2T1l0QNqF7osloGOsmaC
8Lo/sWZyoTCbSLm3nXGYyLbHmOqTRrlafwQ7kKJqipBYxgIk2Xn+VCuOPbMiv/Ex
F+ByoUFAoYOyBXbyJF0ERWumU+Nn0onURIHyqSSABU0HsC8yyCQV5HJv/NGNBUJJ
9CSEgv98mqKy6H/YYNqAuz7YjEf9WCkjDtbtxjP33eM9QvqxqGBiemsVNLGQ0iSz
x6yw7/8S9PEZgEpoqSoCcJtNZRvIvDjwXDHKG7xdhEgCDQziCgkWK2VXCDCr159k
679q5YxiFZyKbigUNhuS6cvWionzZpY3JF/3yyiOkFWQV3YPqi54nNMt2FxFfRVA
bq3dGAUyZ/EvWyk3twP3j9rgM9uox7GktMsXIxn3J68OPtn96hy+Xg8NkF/Rh5iC
8nDPp4vN4qrjB/jXFRlQnpLjOrFpRngSkB04xDJR0oGJgqg8gvWZGbCJI5/ryBhl
PjbM9MCnviQH2AJSZ4jKHUim9FitVuZOktH5upK8EoQ1cZenR1Greofa75joH8GI
eWaPEpHhtYufkGmrSl/p+J8P0fDuVfp07SZLO3t6R+4VdNrIY/8LwQoQVrGcD1eK
3ahsqo5Y3EMcCEO9+vojVO0EsC8iXXCzaOkxDikOXSvgBDBGburgdG38H5qBTkaI
EqelTcYwxnpx/gUHkMbqatawEt3tFlzjNQFfCGsUZ6BEcsjHFz8RyVaygp3OefQH
hBB9e39LQnoDKjCGDi/n/g39f0aBXM1GSk7FQuLezTxr0nU06f1V7YHQg+mqiuuu
c2F88cVj7w4WxDvxIyAsIqbW1G/pm8qAyMe/wLvXil62tiAO/+MHjY5OszhtKmkT
eMkqLIzaqX6pTvsbcgCFvh49QEx9VUKu+xHYWrQmEO86yo0uJKY7J2NDSuw9U6ml
X/VNUSYG2tYbtH7e33CqJPNSXmXhL1mfP5Qcy+imLOkyj38IF2nAkngRIoaUQXnI
VyEulbPvIshgYBtIufg2BRDKzH+JxFwNC82MS5pRR62VWSQKMitYb3hx5bnAEpWI
WiamLqUS4mpNuQF4OCKNkW+pW0TQbOGCol13CaknFlZSO8IoXIVSDeHoeqVBHIMC
BqXfKghSo0crXxRhbyZ124AdkipgqpHp2K1MWrZpznRjoS76m3kzxC66dxf1NGwA
9ZsECbRRQwzoBvr+6f5LOOAmuUXz+hwl6sp2W+NMs6OmuBnsbZsfTWbHN400FyYa
6jvIyQ3ZPFNz0RtznFBapN3VEdBYpR0Z6fUSez3DTW0XUT+rbQAXco/LvC3UtZ2K
uovtCOx4ahJnYqX/yM5eNELy24iLTaVkoY6Gu/SbyKREzvis3Ga5ipaNLa2LG1My
/bw9jUfdR8U1upGQbBiH+xKR5BsGtZD58dy+y0T/GNDKj+oeN/tbN/ccme5wMG2x
P5GCAH/SihQkm3rfleIFLdJfVF9R92MKepyQPuIz60PJJN1Sk857WGM4LKmt9Dsh
rytoc/7jTdE2s6UQcQNp46+ffZmYIWYchPOuplOZ8oah+B8iBoAwvD9B8nF5b6AY
/rJ0AkletjlTWwwHCpHCmr/Gtz0j/n+NvnPXwcIQVJewt8CEbluW/8mEyT2eO0Fn
5zmhQCAoB/Pj99XS7/w9zXwwAtgFc33P+N6OxJ9a4qPgb5DdBh4i9ERI+EDYLBz5
LYNhe4/gQ1Sh6+va8uJctJqr/iBS6gBr7+02p91eoNMKkvO0OS9ODMWtbiPlT2mp
GKch9h6oMtLEIn5hK6ZU+tcHpWEecr9g0Pgj0wK3WPEvzecSuBA9nPL7jNdv645z
Mp2VSBbgdgaCg03gLYkYEcuhXgw47fP87Ed2+iHDFkhmh0E8bHeUtOGEw4lui052
eJJsvncDSluKyyWudgsqyDi+no+dQfguGg+89X3jVUkND5GP4TUnFtzpxRWzF8ok
pdZpS7ZgVnH7Zp4YimCM932gLu3ZAT+Q2rH9hR1GhGN1+sTVk0azetblPRDSzeiZ
kl3fxQoCxXa0wSYCLFHCFKS9ZYc5k5BfdSasaAeoMA7pkRYD56V7VFFEmAqLnMsZ
KiyWJ9ak4OZlDY3BoAH4LYLUo1dBtPt5N+ZovNqqYig5brQsyRI0fj8QPwa05KRi
+QVHZRIjoL5858D9ppI6WDWHv1UWex/EHolmJOvcvSxVFASKyDtnaNt9GyFy9nr6
i0PW2ZTrivJ5rSiKQyCb+202jVla26K4TPQfmhlDKpo+8EdIdmXw4WqX7CTngMnX
txMZt5hf/rWz3cXd63prLrAOysMAWjnIC/M8xKH1JFfy6pSPlMBD0vyIbZbLE1V+
2bNKGwZWKPmj3aMawMf/PicmysCYiig6WQQxIj6r0yXGkAivCExDlkTwujgiZjTm
`protect END_PROTECTED
