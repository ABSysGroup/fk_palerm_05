`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OORga7/7PlK+1832FSqY2LpNaYPeyX39HGjIQQ77ifkyTjZCGbs6tHRJJX1EE5nq
vjuQJakhPMiagq/ayYAD4PdVIlC3O+m7Nyb8uODEydKkNgjA++DtVlopVWTUebUR
0eyd3hzvvx5Ie83Lk5UzLYYv03DTjlxcChUAkg6nizbxYQ6S8btDAG09gNefVWHo
6ut1xWoNrEz+y6a2k3Ahd2lu1VwVi3XSBK3+iyMWVPdpwbO88akqaNpCkYe4pyuQ
/C96FDTq8j6G+pgTwOZl4g==
`protect END_PROTECTED
