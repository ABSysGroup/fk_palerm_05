`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R0RbupCQl54XZhChvjz75n0JFJb5oof2N9mp9WwUGBjOe2I4hZ2i7TMuHbQwIZBS
+X/I4FkeStMx3zsC+cZ7q5EGwu3HfGPJfSdh2M81drFnKTgGpFXW0JXoFojDJkf+
ZpSHzJhVZt5ZU6BuKO/90NOeZ3ObVT54eLdWOxUOqiAn4/XflgLGt1rF11F2Tgw2
IgOTbKVjsBquATFBUq/JGLClZPo1/iceBN+pXqRTCmgxaDlRUY4bA+q6gCU3HdPL
UspfNRMer5KEfQz5GyT2JbRb5LjMBp28qiuyh2Vm9tEC/LOeSaxMgyan/RsD0aaC
LMRELpBQeRHLsMDyo0HK6bg+570mOen+VaqSoKY+M981Wa53p7bVlnZlg6LndA4m
WijSl1wuAy1Hz4QE/V07gJgRJpzrm2TUNDjWoxL79TqM+YhrSa89VZ8ZpQASJU+u
tShXU1+ggP+OchUQbqb8/D82+VAtnuR//XRuLhriLpXoORs5Hm1OlIOpWhRxOC9T
ZW+UOI9Urh6ifIWUSdJ5v5iVfTSAHmGC0ji19QgBMGnbwOpVDorM4/PW5Zq+2VWe
MQ5uA0cNzMuZsFRRMdnzGMcfGQ1LmQRS9RjqalJIDut+poQ2HCyJKuHLApG6rqvr
hK8Q7RM8d8Q2pPJPZPd9iglk30mF8sh+ej8va6ZTx//RPxhyWoLooGd0TijhYjbb
8wLUBrdq1zkoQ2OBZM7XaprEC/Hq6g42e1lPRBPmjWFA1Cl5vQ2QC53grBn0RtFg
L6C3q2Py2dTv3PFEW9JAVA==
`protect END_PROTECTED
