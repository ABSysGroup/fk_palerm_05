`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VfrYHq0h44ERmgQk1KQOLq8KNd16VEyrTN0ymQuQ8jYNwJhzGfaguM0931EtlpkF
RUE+azQCLLzcLkU1RilXERWmluZIIs10wEJOj3mwBK+ygdj7Qyb0acOMDqAEmeIz
gEAYtObYFB8I4zR6+mp2gNPCjBHsXvloeRp+pleoThkk94goOb3g8pJ3AKLBp/yk
3zDxqactB86vnW7pVuu9NWy6h+uIP2rE3tx3efK9/upIDiUq8M7Iexvgvv1bM4cE
bTJi1Ms+SbVieYHvPSAH8aH/TTei3EinfIUA31SrJZtZth43GhDNhmOPDDEzDKOi
zG5PdAj0TsuPkj6ItM3ksvcm/s9edkPT2gWSU5XEP5HdV74lm0PyD9btY+ZC6BPa
gcKb2h1mjjnhY1l/kDwXhLJf7WfSpi5PEPafSJsUhtyY089Tr1i1eGPUetwGw5jX
k5ZJhmvGUl1xLLFqgYTw/RRVNHVFgViX+3chn+8wEZv6LN4EQFiLcHnHGy+k+bdM
vRdNV4UfAUKh14W8Htfu2tzHiAyO7psTBHoxiEDPEAp1UO8BEuiboHVsgwMebyuO
AuEazx2xglxaATWJ60+XoxFcyHcR5rGbTEaVdJGV4kpWho1H7plK9DibMb3V03L1
Nxlum7KtmTmtbByohYcWQWRDsUDwPVxbe8STYAY4YxgrkQ9j+DpuOfxO79DAITHG
7qIC7uRrT+zZh5tZBHgVkNnsTkLzSHp087AANopGhTb/LaJ755wUJvOm6ha0568F
aGhmH3L2d571Y5A8pVuTPPAolCe0OQHLG6f6EU3vxIxE/vPdIjueZFmldPEesEif
AO1bPdpIUAC+2zKL9knWYzV2HjZ+8B/4qyi/zjXk1x43hwbgkRkMwjwC0OPspOQ1
Vw1TGpD+IxI3lkAcOAL/dJxrC3mTYnddnEB55uHH6z8+2zdmTgd+ZN0sBOY8MEN5
cpHfP7+SXs4+1AA51GkQtCs8HB3YgI2EGRzMxD+tTNCh1CPSF0wvHghgINxz8NgX
tOChuQ4q/kLzvEhNtL1Gs1GycQZq2U2xLzpI+Bx5cmHJiEj+6QmJlPqSxF5+y+Yd
xi9G22I70RdHqIvBabYNcgBO7yAfudx5nZNhxaVUPZXe9Zxhpx3f6RzZEOHzOAf/
RSS48ioj2U04wJNwp3WwpFbyMdEhbeJczeoPplQbDDX3v1ng6+tX9WeG3Bzgm17Q
rmRDHEYqum8xmTjBmDS/jo442YwR1A/H6D8CDxJyFqw0HYLjvh/97xCx+1ok1WyH
4Q6T1rDnbJV3Xxm4KcwIx14FkdW6sCrpht97m8EO0tRHjxs1RPSDKvfE1lj1ghsl
/Ban7T/9VMP6plN1rDnVuEH7D/iMZber2YQEFVZ1IVUVSRnHheMgg3A2zTKtyNQW
HceUuz4PXGiEUDiQZhBMRz8jPxBSnVZgWRPskzNeeUTvts7yorhNKoeBebxQjT1Z
HmoLh/l0i7XBvjHsdA/NWtx8uPXN9U5TF6dsXnBPb4awKYIH08/Vh6mRCTr5SXjY
2/ZDTxQYtGzZJL+C4j7oFhzx0T9rLI50IpprfjuP72gk+Eug3tx6zA0Cap1Zp+v2
nM88tPs8xefwayvtZd1fC/+qHTIgO7M4vLURXKbWICbIe+pM6g1oRGAd1Qy8YrcV
0sFsoVZv1CRPKH9lciA1Ci4R+uO8M1kitIMWGaItqxffylMBgLiZZUNMvyJOapXi
QuTpVqI3IsPuYODVeIeXZjb6euOTHUidcFlwmgeg0di/Sqk7zCMC2hfDglwy0T8N
jiXqOJ6kzvGohuWxFqqtTNdo6QrSyzVZxRRWGXsHg0iVTocwD7kF9fhVTcckbz8z
c8Zv6SfEtQYcMHtJ5/vwiB1kmz32GJyLQNdLQiDk9yFPa/G0uJ+KXkhnaYks/8ll
lMCQ5xcRbo7FZdPZpMc40/tadtwbS4ThoNd9qc3hSg7MtCVsutJXhazM8o5hdrHO
l3bKxCEgLdHG26FOKEgLT1qFB8Rbu62o1uWbGmOFz93FV37yNr5i3RZN34Y4EYmw
e0z2ljcL4evbAljaSSOh6/6sgz1d90051aAlmoCNNTphfQgnTGKUZqEqZaCNEblx
XgAAR5ip/hJ+2Yz5APxWJY+KrdJtsZya39JJ9EnmG8t/QtKr3c7ATgPf0h5ICYFM
7C5K4YOwFsFUz8j7SkCD3YeKM0aCi1KrWVMxtq1H5AyMTQ3V4Arjuu3WlA5wvnhe
HC6xm9g0FwjLWk74+FjBnaJ9lqrMFafMk0uiHBamjRGcXNsiAcJ1bmotSOOJxf0J
gs6kds5lhsBnVCetmnyWGXMCslahtmteKlXXR/6yA4T36AqumSLPpiltYvFkHhRQ
UyXeZKsPPFDZzH3d0WOu2RpYFKeInieV429yCzFYH7WPoPFUFjrjmcFENCA1Ai4T
83ZVEONS0wkollL0nbvMuGgX64WoYPUcTD+6CfiZXiBDB0zYR9tST6HDpM2RxnQ6
WDAiCmBJi67VmCwkmG0jfdki/wPWCsKbOgvg8B+kiEts4jo9DfWQ0SeeJCfV0uTo
XTAwBvinkuATsf04icThmBB6LMcky+YkW9zhPYp76q96WnyrTLO8huRCW8aruavH
+W0mtXFak0kVVVrhhDsrP65YPp35IKF0MO3uCJVYlEbPFJwH1+dWSaxjw2NVdmbh
4gGVcNh/3fafvzPWFDRoejZMS7NHZcBtJtEHgH/ZhnnZOubpzJVJVrX2Hnevs2Q0
Dwuz/lNme9zRcgYDdedvchEzCTqi6BmMIIZVwpSt/1aCpTpifbXcuCbAa5pePzc6
A2mVosdJXHQwsW0Lv4TO2EZibDk1YA+gDnUgZNo5CTGqaeoNw9tSP0MZjnfV9Pms
uo+gEgQ7KrJG8B93615mJjtxe/f3H/hQD9CMn38C/w2PEGIIU8lg8vmR3Zh45mdU
ZZzfQoHT9CJETPaMsbXl8p97aKbnSlCLbCOshtbufpi2zKcfU5YexTVNzXQqPtRS
5JqV6naiOcuPwHaCIL38L3PdlMGZDuKL9wq1totfa/JeoZwWmE2hZkiDUm+QRffb
JQHnP5pSEfxoRd46tszJRwNEgkr6IPEArS6c6K1CCF5mQhtXQZ3PJsY7M7lNmgCl
WDxNU6T79yHMvo0Yl7SYJoQAmSWpTk2cRBFw1MHcKBDlDLboXD55rzVxWy7KBTKN
PS3W09VGQDgn5A2BgnjEurWUJZtOQKuZTxfT/fQKT+DIQwKOO/rvdQz3FgAbdvOA
mXfRdHMcjK8abIF/wiZw5c1CD6vc1UtQbroPlGJZwtwZCGjo5yPeZqYCPLXJ5eB0
vcg04S+WcVOJlMPigK+MDCpOt0QkUVDCrC80/ESY9dww6Ceo/GCfPrtg3BGoITb7
2XPIT6PkTQ10DsMFtj7shPUuSvrsYNStV1TCF2QlPBG1vr1qY4c2dDnJMYxLXM2N
5vM/MyR4UampdAya6IbFSgc7oAGJhH5PQoE9ysP5uYIQ5pbLXkFtql3BATQC3S2h
tQkSyvfc2CVRWUSVQJi4yXKu/coVCUuro5upIaFmmOHiuQDzU9uokqE9AGwYg/Bk
pK7IzLItbpH7QcfPFnEBX1+ihwCmFuMGh6/klZYgq3+00rD6TCEP0BlX34LFt0Zp
DxdU67KUvcu/pU4ZIpWDG0dGccR1ndbUNUPQbak8KyduB67v9WH+flwb5XRVmBzF
MAfwDVGxMKrSXuvBEtxdVX5/L8Pwxum82/nMMybnTPav1wis/FXrMPti3VgeaLny
hyhU1u+lGdfhn5As8v5E8CmMMMJVCnlQv6WdGhcoQNY2Tu18BJHPjxPieyQITCHS
3bH4m6iVYdh3kg4mVW6CzDpTyIA+pHvJ5WDolYEaB52gLAjK9dfLfc2h4bD12X3v
cYy162qjNgIa+MR3KW4VE8B5RE2zymB8DlSwwXYW0Z5TpSonQSTct/JYSmRGPqpe
EfQI3RIqlhN4X2cW9GgVKzz/cs7Shrt+VxH97qMlNDYrox7pglgh7EMNMyTDFUpT
e0CdOcbibkXXIaFrULZEkDYhAiYHy1nsIQ4YLm9TrwGWi+Ix+xRS80/vORNUx5bH
n+z81OwleZ+aUe9z93AbTW7dLtcWPHPNSm/lxmsKpU8J4NJwR0UBLzCJcYuz7Wsj
McY1njoWMLzXZ7UUVLfte//GQAKV3cP3yiZ7LufVY0ZNowEb3tjNmd6urzogRrjS
xzMjU0dSk3rTgNdFDYMdap2rjN+IKC1GjlQM8DTdBZsEDURnh6kYKl9Q8b75m2OQ
BVfog8zvyRGCRbZ+d8VN6Bk9V13WHmxlZcT2GOWrrJVk8gwTms0bLehe37P7faEY
//MdJDWawBlPpsRbHb8x5SeuRA4CF/tpkwGW/l7oUugo2VFBYZCm001v4UMuDI8P
wWmYCtbWYHdkR1GB6jcvutXU5RJOsS2l7btppPNFoQDZ7iudFKGxwRmTITosQyc6
berph1hwilCA3flwYonSIYF6Xa+8Hx4o24n9GHSne/bUPy83g0VvH1aGme1ppvfc
bu27r9lYScG3zLlP3g5Vqs+jkHoASmu01UCfSzywHMnc42UQsdGUJqXiXsNO9edH
EH5sn6UvDu60MJvsjLwwMY7GbTSTzKYSdMcMry1uT4flcuZMGYa5LIFdjNCY51op
MC62B8B6DxOAkPBC+SkqqplKTtfOOO3azLmDGjkGrRuarkEFJZawDpvPGPx51TGY
V6MGFHKqf8daYOpPfzCaIE2sb7It2NShcCt5/ae248gu3hZVBoJvMQXcZ2652jt4
eVEFlwgZTgZXNW3URgpn6EvTb2rd+ceUjIGmo+1ZtYzTm4Sj7c9hQ7Gbih69z5qs
0xDYy0T+gRqFaJaEbsxbp2mSluxcMJbBOwVZ9kF/hHr+DR5WEN5NHJ/Dl1XLNRWc
mla8kEHEfPDd08czvL8N2x/zOSQvNj/l6xnsWEiN+9p3+xghhnSx66YKC6oG8klx
rlU8Kx12gi1dOGM4h1JC9gSZJQ3eo19aPlWq7PIYmaIxvwHoUsnIQCi3GLXnYIgq
p6q+ZB3HLV4+/GVaXkr8ZfpDZ6LXvvGA3xPsuUEz8TFkGCp7EVJ/sKAHgTdxEpLE
afYu2kYksYaYryZiidVYAPisR79S/pWPcmQaa/lPZDYh/JgJeHy9RE5H1ncYEhdW
e7UqNCtVWIgnbeVEDcj1dNWgxO1fTUTOz/JpHTCI4Zz7fw3OQodL2V9xEgcZy0/u
fAcC/Qb6ULR2i51LJCxPm4FsMgBG/uqo0wUmXifHIJKZ/GufICL3eCWQjipjfKWT
7PNThDAb8LWzpmerLt7XBQ==
`protect END_PROTECTED
