`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N9lfMGgb0TVjsG513TT/aySrDzafiFhMQJ2VTiSSilBEZVh0XTRXGUcqxVXw/3cJ
Vw4jZKUSQh3HVBk2rcYEQRScG7eXhnEsDQAWfG89VhSAK38nwpxR9sTx4UdkGEYC
+fHulrjMPrvtihQnfcxpES7+dPVKdGpihNCZENskPDHkcBSDl+Zsw277bta+1Rms
G5th5bIfLzjQTgarx3Ou3IbP6+wIhDZKVg2GjqIUSRwxUEMl9uMm1UVDu8U6dxde
5zitdTwn3KEg3x575bc53Xr5R/7LAmA9LRoDvuoGAGoLo2Tm06sfUyfm96AiKnN2
Jhr9HaAqirUkE+U0yB6WLc7OvyeTqW0bSGpTAEHfcZW9JCBH8uaOWs+td5czmi40
W8EfVeM8FDxSJ8sJsCqwCfEjVqgpqHeKnNKVaKvWlFtiTaDxn51bgR48hYZh+ls1
KNq8Jj0KkSriBGX9iWI9UXlGWgOtaC+R97DOAZFgFmyB9SE6yTt0e9HQSi1OsYyQ
4FwtBvDDMqnsLE16e3QsYlbTedCjn7SzPSkxUR9c/Nr+z/UNl68vtsAMfqLhLZoi
cnn0Il1J8UILoNTFjdfX2ONGW4PR79j1EF4oaxW3lsEeAy0c2/N4auyx4pMk6RVu
`protect END_PROTECTED
