`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IenrOCIRDtVbLJm6w8S8JGXtxZ+2Zj/gMM5hSsLb6WSexfchh7obMB8zJAE14J2h
Jld0XZgdKmRwaH7WUUY+2OFjKboWU6/QvNyOPkw8kUQF038rTPJ9iMj67Y4KWdYf
f22cNXd090+HcPWMckJ1nYsEg0gLgigANWER1aJqpRhd8wSewuc2dry6t0GjW3mI
9Sb/tMwovJz9cvyvlQn5x2NrLZP8MQaf1xk7RViUQh5JdgHm7kULCSTNgUI16yBB
MtspICRMtwQvhjVJHe58cIWTxwsf7YoulskOWRV8Y7nXAaLeutJDzJ+0RZXxWAIh
erJSXRB0qYjLyVyoT4+/YoWMjrUioN/Opl7zM3CgGi9G5vSRJwWpR1K93O0sIRiG
qvyGquP+lRRTcn3PD1oXh9d1hubyn+1InZxLjmSqKo4Hjt4qgxMA5/L5b1gQ5QaZ
TdfK3gARYtrXhaw/tX8iGH30E98bkBD1I9OlhN/JO1Jg6+gsoW2mCwyThYuqVAb/
Sqx1oOtQlyTwL5OVDKK+RuefRyQkFChBAeubs2u503qQyhEl1NMHsjlvMSDPFCny
9QkThLsG3TFcfxu8UVEueHM01xjo/zcBvjtQOeQ478k=
`protect END_PROTECTED
