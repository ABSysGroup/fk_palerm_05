`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+gIQ7m8Gp8PxNxAiFcqBZ5srfLUbo6uh+CYXQXBO6tciYsWOgdPymWH4Qxe4tuU7
1ayqwJiBOfpe5UfDJXjb2A21kXsPs+yIsaeU77S6YlCPlArdfXS8Gu0Jc6fixbtY
97AGiHCovJQ/9QE+CpQlYJ/h9K/EzuU57RD0RnatUhlFVC8fLym+zpT02tkv3n8G
+ImqcZSaXp9uWDdtDYuZYqxv99kJyLyar76R1IiFCMzuzEahwhhP1uN+IKIMsf8R
Dc2Z7qu9B+lRm8uxor/ieDsfKxPz1quMiHBfMpqnU4M=
`protect END_PROTECTED
