`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+BBHycwmawLgxZqBjKDQnQSEtuxNhq7tibiflBRKvZ8urKdGpY1ecWP5pvSTlVae
9D57231Cic8qIMQ/uk/EGYNwZfQhM/+d0DGP7k4GYwhaB0aAwCkt3EtMaMVJrpck
ZADix+PfdwwDftRXmEyPygJpUNkqORoW2piedgYwKYQTkbepZXX6Zc4nzpocOMQA
3WAmPYpdkTOBZiACJTpjm5K4uaYzWhebFr+b0SpcMFxDNJpKBnYu+/gAmHYUCjRp
RF8/ro3A+Zp+O+L8UdJfRLHuzIMB3+zYrysYvPADlIKOwsL/CPeGkSLggrDDpMul
K2wasaEAlDhgVdwQBH0CX8UxcDbskVHKbY/pNIHn8FELLBmBcPBSS6QSdqy/VF5B
S7qAQ4zQ7+pszUyVBGKdq19b0SddIfQj1CxaFOhor2TMcjmRIfj7a4EFSRusqlfm
n9juPP+hU1oX93zH64chUdiSeR84CsvhcZrlP2++HCaJlSaYPaPwkEEmArcuzRp6
XQmrQHX5IIWdoNe/2rklmLfBeqT/E/JjDKk0fMKvUpPPnHVF1k+gsjhER4bztNdg
rpZMwvmwtI3o6ju6qymkwAX1DnwwElytddfHFk11KxH/98xTT4EatsfNgYxcfGRZ
QlJMZ0LP3J0gb8wBMRld/Qw3S6boVop9ARTCHcsHmwrIVGpwjRmVOrOKum426Rbl
fZ2jNNj2aeDArDalDH0hU3qu2HnWD1cxuLGFMft64YroEfe79OR/qrEvFGRkPDBT
e78smuyqfb0VryapCfn0w7BrubhWxF87LHBsvu6be+j3WXITYTKqwa4nK3Hh9uo5
i3KqPxToa+c676BzkE/4JuimEojmFhZ/UKRn1B8Hi8+/ON8Y9jvfY3v3YUBQgylN
gFLBFBLE9N/pENxBKZr6T9zE+BbvdjxkxRYWsD3FdwyI0zyWAR9XmNJx0Rs9O3Hc
`protect END_PROTECTED
