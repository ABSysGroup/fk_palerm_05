`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M5eQZKKJkEPXM6gjuYr+0A7my/MkHJmaAzu9Zhi9wxI58oJzZ9Q4qforYx/IAuPu
0FtIz+O8mpxPzbjk15kaEvdR92U51/bOUVRsFgoORyO2b8jwgOgt+a2ZgIkpG4u6
BJolDmwhqcPaVNQ55RLTxYSEI+oO9f+JbNhr7Md3lVWpgBQKE0BGDvIKkiTlWp6R
mh+vBwdKBYZLZDDDtc9Tb4JPX+pbWHuG73SAkOZpn5zpG63bGrO+wBpfI+sgmdDk
FSCoGIZSW8LUglillB3mIwaaMtS4E4fpRwfa6vUL8iLtBYtA2iDBjEy84yXIC9iU
NDGCqZGETCNmx9byFYROyhDE+7TR/YGvtSy7BYGUuVVA//EKiYO0RUiE4b+o4BSw
vMmQ9jcFgAKFYfLP3P34C/73eh2RtcILVyRF8daSyzWIaIbimuqmvllBiUiQhNkC
VlDbnx3MjloodNj0BdMMa1FMbTr6LnuxMv36V42L8d4xhZ37uxjlCfh9Hzd+4PtR
eyWH/Dekq0TktCI7PQrwcJ31Y7jaqFDtz01SvLc2jFB6YV5Y4g+b4MCsn8fdu3u4
wbeZe+0o62K8bmCkoRRH9wuSr+8nG+8Mzk0YDnjP59GObphLRLJC+9ptiVRqk2Or
/ROlEwzJVirD7vkl87yhlEswwr8iPiuHPHThUXnkPsSG9V0DVXC7WdVxhfRYIaNx
nH/tlCqSQra0WGp8G7RBvfsgvca5wSQ+JX9Z1gG+l4MnnZt3UHnEGEqfF1jNmoAA
ol1Ww9y7gW/9Xpj+t68qmHey5TzsqGYr8HXx8XMZuqtqUt7VeIgzJS6bxV3VXWFu
x4trD+Rnn9aBuhj9qh8TTOZim/hKnyOcXWxy9S8JbKWsDl6ZTVeXcWwmn023cQQQ
jcqGUsEotIGsOgwnHFeYTjAYfnOHrnbGbnZ+4iyDpEB9BVwGjZQZmoqglnAx4URF
OjpRTzN3lifx+y78mowDwfVkE8XkZmttScyDDcOAu9JxaC5wLRL+fMh0V5OHRfNo
8it+DARz9xvoeW4UV99+DM/dIFwvN7XsTIPvIYRycuEVoTEIWx1l9Z41CHHv1a1E
6lfhPZt0QppZLwbYbDjF7En2RbzVJRN6rLF1N/vawolyxyhxBIUpLkvUYbHDXtLr
nYqK1TA9b7SUbz8EXWF6H6lirhqPUDpNwUqDTTYFGZmtjfRKIXtZTdwIHKoRnG9O
5OOVeDTVV2F5xsWtwqTaZMGNwqnLb3MWS32+YMn3V/V4UDjJF8iVveihIjaQhWrZ
N27GjAvzhQ9RX9I+h0mqHL2DTgMIpTgm5dxX8K2KAQUOZoZHVjFdO5snACiG8M2n
Cz6KUEjSpMx6p2el6HDWlcun1lhpCDSHBWDf6rHCZPB8e3JQsk3/zfszP/m8RZML
aQWRz3RXxoNqLLQ5zzVs8f6OnHfUh7/qWXa/4goEf/5Nwb3N5IOI3TEhivIQyEdm
S7kbc6TJQuR1K28ssVvSwJRLHxXId7M/crtkWkXi9NBzOUvmo89eAM9P+QmAGhX5
zFj+88MOgxvlNuLUjXG/8SOAbVibidDzlrlUARYXINO5ODkG1twtTo+ojA8rF/ec
/oEgpg7VaByr7spg4/TrcN3mS7gVVRW4Y0NjuhEANDQ6ySeeYz7ErhfFyeMIJ9PS
yvyFnNqwmay4g29CpDVTexfB65MluEJlS6+2ydS2yYWSqGnDF+Il1JQs5Iw3clGR
Ky89iRVWLADYvWDso4Su+VbjeggZJrDtpMbL1LWDHoK/pHAAsCInIrfayorNnW7d
D22ys6Y+DdIn/0OssLgi0Bqz8muaT6rSXP/GJmMpGHhahHPUpkYcoUhe4IRquTVm
JG+9F92eVOWMCVIIE65yWZeVwSjMDENpug+yry5mz35pnswDCytYlP3rRph9soXn
Vm3ZhDO9WGtsYy23c9DOxMvhQQHAFZciE9HLLdvnM7v+Q1ULx83t3DmnhE29hf0N
zVuRjl1L1zbov5SpHDvdc6OiEW4tXZ+CHp+j4zO0avMarjmw57VSjDQNOmLJJ6q6
ZozRqXbF0E7sKyYBN32IOsp+oznoeO02WzFX76jFL6n3Vqm51xtL7NBFx6dzwElX
Hp6saLHhCe/LUxaxi8hxO0sZ1UDuTchYhBO0ttxh1Dh65Kg20vPgWzeN3fir/slU
OM+9bM1RV5lSIujG2udbigCVbv/ybgNShtTpiCLCipcpi/9BVDz+6BdkBV+XiBVo
XXIMIpWSHIzx+SgQj93+t9gVVvwatxG6JsveFKjtHpPLyWOKND1eHjsyZKd8VpBd
HBnWkfetW8reT0LcSMcR91BWc1aDpg2v1nP3NmB/HCTHd6l5kfHRjX0BN8xC1SAU
wq7ARVuIMb4dSdAutKiJbtE9ixX7r1kJgh/9aeeW/p6PvmYfUy10aVFBB75IN6sr
8WYWxekwA1nptE8veyZO/tvf3XoLTDB7BoYAdrd9LUOSC0o9HDuokntqhNu4U00m
LoPf1dgPbIl3fX7Hzmqr6sIOshMID53Drvednr5PV4EPDQ4gwn/KK16LkiE5NnAF
r2a9oam4BEdEAwQ2u2Njtrzp41uvrYKkyLnaxvCqm7hzfJLTGQQlZx+dkEA+Gtc2
NZIPY58MuW7CmGv+EoNAm9p0jpAyMuqALhHy9ledupmaUIxq+lCjqllBCni36fx8
g3TzKb5nH+X2n10YAcFgneXDqt0LLbBo7s934dIBso/Aw49rXpqtp7SLJvPQg828
RMSmBS+OlDGqu6yr7ui23+Nyo8fp74JYJjQ5RTtbosPQ+OFr2PoIvg0/cQ/eHuV0
kfWiBJeZki0f+ZOyzKiZh1+xeasrPmVTdorHrRh0Ub2fLg5Ywry0VZjOPQAV/qY9
Lq26uH2a7eLkh+COJVANg1E1b7GqJhvpNBqZxYN6uOEs5sQSW9Qj3dBXwzMzUb4Z
2kqtTDkE9z2ALPG2rHL2AfAPj+y/SEifqKCe+A6Gg/9Wr/5gafSz+wLA/rjM6QOJ
TRlK5EwoSfSJmIgIvRKdLqAZtII89W4sAZFdGk7uLlRxdUNQlWb0IfAZUNS1ehxk
i1fQJn8KW7tPH69BKwWV9bJmoQnczkclzj2jE/xPi7WX3Pv4k4pUmL/vKD9C/jSL
ec2DLTAMPumxz9HX1YJER5jrgM2Ky13ugnYeGrhb9RsZWvstHewOihT4CTOmDJDT
+4gfC4TxPMXZsnqgqoKZWa1cbU1osjI0GaUtrwUHGXd4pwQCPk2uIKpxOGZ/wtP0
FD0zBLovxoUTgRhGJlRir0ezz5CBiJ+Jel7YPAU16C5EDr+ZgoYbQ6CJ8yIR9jEO
oVv+xazyfkWpRRo3ihNd2hE8LV4IIdp25xL9ULJEFNuJc2l4y2zeyDckoRJd3PuJ
xXUTw9PGpbgLQr99hxXy47l6C7Sp1d0S/WiCAd+l27z6WmHmUscaaZEgAZiyTW83
1q2C5M0RYkAR/dfI3jWUbJBDFbps9QAMBLqNavgtoG5PUvR1+66HG2nUKVMi+sD2
xpxDq0dp0fBZWHO5uPrKWSxDNDgWMxoQFNqgMVankhpkC4iN3EAw6lth/2IIreXr
3WURRCvU1gdF9cvLpGtnv60MygIqwxW8GZtBUEIVn5MmY0Q3jV00vYgDST0BrHIn
r7nv2vQqAGRlf4J6x4y9AcGUn2mfeVR32mmqu+gBGyQB0a64iggca3ERTaq0ho3x
bq5xKwrWMO+cDJbgKARsjb9B/GYcPwgIklOihk+9fESjuRqGyFQTF4w2EQWOdH8P
2KrkD+TfthAK8SM91/dp8JTNc8jJvFpejXSN49qb1z73Nfu9/0ucgupU6YzqSUNo
VNeZzlNtmF86T4RMrpuiz9j1HJNOAzCf7BN6m/ekebq9U2PZPJcV+hiuXkbIH4TR
8zPdcKKdHhS7wABZjTbmCLS/yNlnrxgcJwm+8DyAj8ro1j2+auoqEuQqsAEwQ8j7
mhhYtuYdHiGVPwTDaR9VTRCnWqY2Q/Ux7eSaoxIrxVCI98YJnLjNBO03pl+PrZ+j
tuM5igaDypkCIeDrBdTuAKuIZAN5LyPpUUBfAJrvDir7TzIkyuUlC12skrXdoiMN
KflJqBpTY3Z0DgMDxNIY3NVUGbAslXTOPvquDcUKc7IAvXeyjdwSxLeoBUdpWdsJ
qdxjEKQ7Ui9XtFbTKJIm9fmbqizLNaND873utYwkoo0JBFEeDj+TIUIeoSARW2p1
5esE8FzFnDk8sErzNbp+1mqpRT4BG9TrEDhBHMg41/BbwEKNrXrlpuQR8WUWVmIA
0S9r1zmzmAdhYbhpm0LwkTE7yYhXtOARlrUwCNKvfbIEz7e3es4SAY/kpGClbgsp
wqqVcCxEb2D5GJGs6iYNMRX0sukCHFcddLyL3EpFeZn+odmUR3CYyISR7isZ47Ny
axgTo72/eXwyMMERIGkBE1ZEUupSbudpav0wuF53ql7R/JIES65A3I2nzMgM1xdE
IYK9DL3D8qnbM8ldiKeNjGvnXmUMvnm+WGt18+1le8rJ4UHVmaU5q6X3cT4CbQGJ
/eHTsB0vYCUQb63kLe1tT1sbdZSzmdyfOuO1cn0Qb3ByrhgenBWNVZfg2hDDf59i
sk3/wX0C4wfxl8DEfdmVKQ6Tws8ftWoAK5OxVUm4cysUSIhOjO0pgI66BUsAyRgU
OoxGBns+HmfGtszrSBMKgo6IQuUR3iXo1yTRLizv8KSUtPy/e1bnkC3YEqu0LCsf
MN/I+pMga57LLm3szgDSzaxgOPXH1DbLG71aTkU2ekKXwbxSkiLQRbAOt3l3bG1Z
RjC8AmPKUSr+/zsT2FbZGyUn8vCYdKIEyQ9l3A9xNhA0tnoEmZFHB3Oiwgx7Zsvg
emLhSAlhyecwlr9hRwiqBpI9S6OI8jbexWJaatMuSR9JBOz22Yi1Rdc5CtpROHgV
4f4gY6tL0lmyhtJUCMjEIYy1LviqBKlDnadHd/6vHM6n6RiVYgCCeAv6me6q2YUI
E6JVxDBUhDNdGVbGPBqpt3Rgjx2VS0HvxkxLe4RMG8EJX9DIthcbp5+/PJvd7wUI
K6aJWjhElPg5SaqI3vWaWyZtdlizHWJdozKX69MVL7TAe91mH8KaqMAXUdiUp8Cv
oTD1Y80uV7ECNwoGYonCTLPAXEQoU8sIKDiwS5xSDjpFWnLGjMDiUrKpVO20Ed+a
5jsOZSlaRo/Yyj0zKKaU0XlbCbttXTVt+DEQiGMY0OrChENqfAqZb76JV+IF64HR
JpWpJzXhgURttekN6b8etdnQ+NpEOvALXiuyTePryjKaOchyM59kUEzFagfRxlSq
OeBoC/++W4KoIPHD2qJvBQnnWSZg6XcBMRdBdlCaB2K6dgZ2gOdhcCo5m572LzJw
BlmDRRweQvHspBP2deanL1XNw161oCu/ns0tyvOjmHYCwolZLitxgHYV5/rFhr43
VVx6wMa2nCdT5gyRGd5HNPQEgf3R6WrDglaHl4Kfw6RDhR6uYC2JLCqPtbr/yQU8
6y1DDc7xfXUEQgsKJbbycdHFzroyAgeWEgtvSkGbg4m4f1yudVNwOGtgbMkcYXuK
jtIziwY2437EY/fBzSg/gdB91mZ4N+viJ4olgoVAXGPfs4On20OFuI1NeirygCoJ
Ri2xwEzsG/f/U5bdi6JeOI7RGH6HLiIwdWHmkUOxi7lm3zr+VbUQSBCILhet+LqK
z0sCOT1TpBsDhzX6JJf6J3T2UffaAE2O001B6nYsI/ubbNr+FXroWBMTY2BNS93r
ikpxaU4ce08enoJj6Rq1AjzwU1sZcNZ9ZnX7Z1GN2dzAH8r5emdPcrnb+2IbNCsc
5obk/Q/IQ89ydaqacWFLRAjUvk9mtZUt4vjr1A6V3Uw2kBOQ6HeK+AXpeoQZbBjc
YmIA2iEZMODDTjE+huJl7W5pQnKUKbKy7/7TKvU9GHiRmAo8bD5qXX45t8O/L+kE
Ju+BA2ZpHPGILRPSxmh0Mrb6ktjPssicDPyeOwGj8nMEwCh/YGTT/XOSS+SMj/Wd
JV09/NnLfb/uSnNRgjFS529eEpZW82x7uu2W6/YJ4hmwhClylGsi3nxk9wlV54vi
attfq9CP7Gn7q5HKZTA8MOWYbwsawPfQtAi0F8GSQMWIulCe3npA6dyO7KVqarwo
2xEpu4b/ola9Yki9b/UIORCr0a3fmCR74BtXm7Hnb+aX9E3WIjGAPYnCLpJZdjR+
YzI4L+W5R3A2nUHncIgcx+kd3B24lgU+f20mfKiuw2bSU1YHx4vehZhaSDDYSENg
oPqMj/8BF8xWFl9fjr5q45Rgo3Zm4GWl/Fdcad4799wNvaTeOA1PZg8SZQoU3UMQ
QOQuLtHbFXzDFHHG2BN5ffAIGhkKPVleALogmOpdVToIoR29UIr/wymzhVs4aPoJ
Id8jtI06bcSnmdNlwAAy5ZZd8pnZMZiV0XXY/cc7RMiWX7gBxOgvFqZVijtwJNl6
20aa5YjiCcrTWRC6r0AB7yzkk7C9GkAxm8oJI46UL6PGyZikLlupX2ZW9boUk4u2
dgaB0wIsjdn31pFXJSQ2b/jq6qBi7UYnJqDk2ESa4I/cHCCqiXgOaVCJHt8qjHJ/
czaxlmK85PESH14EeLwzpIS5rFj/9Ytu8IhRNtOgyjstWnA4/6TFCnCQYTZo/dx4
tBokq7SG3a3QGLafJpFpLlcwrLy40SWWNNcS1F5xgS4x7qukMPZteZAEspEpwCHx
QnG4OJNt092yf0r88VhiYQJSWoGBbwbF6tcC2vqYdGm+y++EyXylbrnB7YA1z4qy
khfT81zEvRVsA7XcKgxT+mwdQBZCiYSoaSdlpaC5iZ1KtML/UPdduinWU725J+i2
Yr6hOvcAjnO980Zvo70BUktD18OHVwYN1CAbm5CC4fP6/8CTJN4IwPrD9Mhe/7Gx
joUeWR+0HrUVJAZKTfbUDGdkgU9sKJQbMtKKMNWCfzvOXhKTvMM0gMzw01pp2SgD
nf1CmppD9/mJdR/C8eFYJIttbqH5/NQZcsbYCtI69it4CQapRS5m+/PhqMv09+OW
m5zIhBEIl/G9m6ToWJN25qMpr7N+kP4vQxht3v9TYxs0GLOsK/6KXJKbm6Lzlpnp
rlB3TkgWMON0fwsyABXHzNU0v3XhgVhpCqrWsiJJ7TJYtkBcJmvtTSpeKrohouIL
vkLHe4eycxEoVAzleqrwv9pM4ma38+AVtq86MdeyL2yCxIcQlPXyGbhiIH7AKeX2
e81DbZBDtkeaYF7UN0lxs17nwwdCxmpAxJiKZ5pIXsDxTgyK8bT1iZDQrVIbhkuB
jUWPP6Gt9SQ5VTz2tVBpER10FTFQLfFHPhdXnidxz3MKRhxB/1lr6RCLPBd2v2lb
cZaR4EtCECYuc/vZKBQyBS9tQZqAO+pYDmVh5l2LsqcPlaqTwbQ6SKymPc1TwRtP
izcbsoGmMDXbgitFTUyO+cS4fHb1IYnP4gU9qr9VrkBl/rEO8p3vTZ6vKDQajfKn
vkNOswIzU37q8+s5jSdCGkDnLKPTz8QAn98G2cCR0GLdsCWFzv4GxjdC3A6ixCdb
iDWaYpmIn8Pl5kq2aX44JYPlb2aXwoQA5agWyCdqkiZSQhKh42brkwarORGUBDKO
XzF0//QpQWXilZIIO4n+UoYiiOYDIsD8x1wksRp6G1l+nGpDe7jS3IhP0jQYIidh
DHxRoRbaboy60L/5RqI0NXBinwMXhYMfKF0hqbt8enpiqsHl6OX4eODoTZiT5fGY
svJBI3qpAFgMztiHtc0dmXyj0+CAlsbizy2TtP52f2ElE7gshateEcSBtazgAwgY
izEw8IUnQ3iHmF+awHsRpydyN9F0Szhu66ttxQlzHtXVcnYjDPkyn8s+tRasSQ+g
hpsWTCuAvukIagrgmJOZFqib7eXH51TwH8pIGDMs5F08s9xlynfG5UrZuQQi0Idh
wWKbq6JgO5+gHsra08YlNxp+CeE1T30cP2H4YwlkgHqFz1CvwbWfX9d+g3A2sO9g
NjJkUmnRjQvwMno39vuTl55kIi91RLFiFPrDokuLvHnVVOMmaMVT7mKKZ9dRYrj2
Ve/JnVFN0zxVgWcVx9dkeS5W8GoBzSLY7ZwUdsgh53/lK1ul+eVbNvpdCFEiUjPf
ZRn0XbGpLtfWlEriyIlA0Y+0V7gV46kIs9jUjSJ0bicdS7IGVTYdJETt0TyEUZMW
nXkjfKyRVvDdxlMX0veuOVKMzFSSDk3FdwAcb7fb5j2KoeQJD8hQaAupiwP778i7
oxRq0O5NTGg8BsHmzQ92vJaxqndkyXOsc3O1EpCVHMXQ3XviUjrcUjuBHiS6NKSM
VCsRHP3+E4tkPpN4U8bimkaMXuAgItrKApZySn64/p5TXteSkCqHsvu6v4SJfWWG
6dxRC5Yo4gK/4RQd0zEdkPZPlpHRe3HwG+FZLDZUMq5YESbsviVN4VCT8GLe0uPU
VIfLEnHTLjSotV+cwuiQ8H1RJ+yPF3s9pnAwXqdZh/y6U5qRAx5Gk28JZsulHzsJ
MYCYwpKSj8yep1qMAOobRihbH2psYCXgXsMqUUCGUoitubfIbM65iqrQmjaOI8ZR
3XwyEKX5SkC5uphQEm+2lFOdWtKJY5vUrfAojR5697D1lLuZvERO7F3g2u4exoPY
1MpHhPU6m8LEWhU4etm6L93tYCZE4nVI1aBuYFBlDfTrvj8kldaxuJHRiJJq3Md+
MMdfdq+uIIav9i/uc9m63Pcqa6kVABjTzM1MDzEBEFW4x9W0g2mpD/Nj4f6IYEWR
vmuXcJfzt2+YrJdA91SCyCKyeEdTOFEVCwuBqTc8dY0kkP9cYLfBUI0gltNbLHt1
3DNdW7lPDhr20YesW03vKr74AgpSWke1HazcESEYkH9+eStsdRLCCyLngD0LibHu
eR8Wkan82jk4oF3UyccUNiUo1+sWhcuXlollfhnXvsidKKjSWzh6Obl/CnhLBV3q
u2EW97XgTH8FOj0ERkqlYs+zHzvs3m4ZO+9zSl7FzyYPNMQa1FYV3n1VBVAfN8fV
bkQ7B58rwW8aqO13TF9gBUTIa2SEFBLL1UIo7t4H5qvU55hMh/ne2LZLi+f8FQPE
pInBjdTqyplZnj9E8JinWBV76qm2Hw4PPVvup1hjbKinbcG8YO2timHWp7IylSB8
5T2qR5EmBS6b6cCoe8P2WnujgfC22RNdzfa1Hy3yxJb5jkCCcyatYhEyWSyt423H
6F1MVxDgGaO+N8AXNfZd/9p9tOd4/pKodUBBKtgdwkpCFRRACTevgNPLLFpxQE6i
hQKJNh+vW7jXlbH1PAyqG01qTJLM7uBW1ah4Mpz1Lmcg+RU8LefA2z24MhNOah0V
tHOnewtvKwqg/q+gVPAl2GBpTIjgHkNlnWW9q3DrbhRuHg3XyVa1zXDbTfoBizr5
nMvfK+Gb2qXXzESodD+285YOZ6wLQC4zP7npS+sH2ZB4bMz5lPXSgxXrlWDwW2Xx
Uw1LtEiMgsgGNLSsit4gey6XZLSstqTPL2IDYKuyl/HhO9qv5YmBAwF1h/dfbeZv
O1hyd7EubNIz8WqG8DDcOL1ErD091gf78ApIK15vjWNASkTHURCQFWjFz8jSIgb4
y5igaQTYTrWAPJFblvVGwkImpAMo1z0wY48/zZADheEFGey1E0DVucuvn3LniOqb
rjyvgj59wOFtOZfYdkuiRCDMNq77+xsKLfHUQiFudFF7yuL+5zWnQTDA6Pv4k+oT
dAWypdDdGnIIVFy8h5DiMgUIetWSMLDoFZa7adQVQfl5ZQQ0QkFfmQlEpns6gBVt
Binw1Rj6oFKGGLvLAua1I6C7OwUX39OyeQReC9HacQHsO+zviwTK/9HiDVlkr9Ac
VXEBTq1NuQ413tyW2HpqoXrtYIyIzFB9JlLsUnrzUg2RE5NQwd3cYek+Vert2Pvl
KjpIacs0A1CV2P8nsFemH67diujJH5i0r35f/CUjKQ6BmtkqmJvF1HpYOklcTqzb
JgXEpmC/iYFRusKZcesY/a8d4rge9QifzX7mxhTktFOCCLGyZzG3do0QqzG8LMNX
PNf4078Jm2B7BByjSKV7xzGskaLeb7wusJ3XcZrFDqkww3tz7kpBmwKEOWEbC8FR
e4jQaJ3K2oSzJWy4fP3PZA0OTeC6tCTh4ZyNYuSgOBkx/16DS0c7TB/dNpOD1aVc
2yA7NW9cHGIn+nzD5LpldZfKAjz/2i2n/BvXjiG2N4uUPqKLwIVb28cTYPJTilkC
5elUqJQOYzFhmmFbxwx0pKpkIiwjAID4QYc1eSBdVA4UkHbW3J/Fj+LUysFL2pJu
XAFQqGXPzwfuxrr6sKnhmQDbxVNrrd+luniJqNgVHytRyxreEBQugFHg+ws777OH
OeUO7u3Q7qDe/4jJmhPf9ENXlvVkG9RcP9CjgGWqrkXTyOssnqcTVtIlH6VkTCEZ
XRplCeZ4fIugaYbqnPoHDJ52cfPODanV8BOthi2HIfajn0fpIu34BDB43UYFtTGV
viIrBf+vDKtXHnnrIzjWtPcqz6R5oSYabAq+jeFoiobMuaZHalYPHwOSJmAteYWD
JOSSA6tzoxrfOZKUUNJZOZB1+ND4vT6sMDBvDqWDyl8=
`protect END_PROTECTED
