`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wg6TB6NMAdYStyWLsGG5K0ls9QBzKRHMrgidsrWnLi1eaOZumrk7UcAZU0JNFHXk
P+7zSHAePaOPumUQOHokHtSGyv6E7ZGCVGjx8pCpwAmcuCNKRA7B+fIThCaHbQFL
L78he0yivtN9pLomRiwHH7AVq5hYxX537sLBMubUaPnAN3YXXN5WAP7Hkk7dG+g7
n04X4Z2gS8o0RtVG/NOH25k7z4N2TSMJnoPRz9ed1xEH9Q0kqzktnp9wRFYJnRQV
5KS6957E8U2OcqnKR+pwrr72purtQauVhhIdv36w9lET/6OlQx8lbkBpIy6Za71d
1utYu2kPuol3W6siLNWb3rgCgMrJ2IVZ1MUVMCh3kdoC2Ji7yCYO9g8uBhSye7fv
6awWkhffsT1/2/D1hR9aYbLHClUfjZBJIA3XFrpH5a532w76s3Jmgpp9Dzy9Xkic
javWRHa7HcBDLVR6NivFrUYtYvvGCKPn3mcnmgDaKP0lYP29wl/D5pCt+bAFzNgW
n2AA8VwCx+XA5OagYHtaj0TbPljDQtYlpjaDLnOWzEax7JXuFoDUc4XgrXzIc0Yn
Vjgw2Tdpv8eWssXGG9slx7vN3b7IKno4zlUvRGJR9RTTe5PdFikNvW1S30Ig/YdD
60nGiq4GX64hPnGSEMHzjpGR0nsGqgyCgaPu79ZhGI03ow7WGt69e+k9EXZ+dt01
dKR+vA1cMrf71HdzNvpwioUaif7HBKsI99MqiD95lwzicqzpfh+ouQ1KT6gtafBr
DxAV2SKSMuGUueV6y13VOynML/r9dr8FUy5KqHssqplqjq3AZupRRCIS4upa3klv
9HyUQK+qaQ7dTmNjSWXWjG0gq4q8WwHtdCSYBL+Nj7FTl6JwC5LoLWQ5jXYc04GS
JaWdv/uVHsBAZC7oiatXcTBH3kkgmkrBiINaG1Zlbs3mJ+xmIjp7d+gFpif53sB2
BlFmlghMd5F+yygieU3h0y0D9rRhvEzdxJ5XhZHO8D8rZ7wuVy6Cj+6eTFwupZyi
Ewx0mpQngoCJfSvnbeO0ukWkV+89CVr9Wosxa9q9YZLYLvIBYx+wKdvUA/UHjCco
IswC4UPHFWqaMVuEJh7v6pM0mmHvKp1728ah1XMsyJenJkoW7LH8zA0kFhdNjHKx
i2BqUsWwTzzqe52ogP5RCE2L0jFIVImTuv/bCdhqd3eJnzJgD+D1EXlM08YOWbHJ
rPS89E0mWEOjaID2Rxf8L+1m9rTcMkeESnEp92ENp91XvhF4mmTgrr1/eC856oNU
ha1SbMfJfBoWpCYs/CWY9bKcMOMJM2rdADxTj/EPDN58e/JgvQw/T/ezuXpyNZqj
9dyhrqvtlUDXztmuo5TQKAJqfGvm6rrG/IOmDZwMf+CmTmo4qXGBhWRdKJ6Svzo1
ttFPN3Z79kBtRR15xDTbKnP4xeYktXOVm9ktKQxgsjUVeTd+fooBy28X2+SFZHAb
vghK4fcWhiqYER45OSZm+yXnGzCaUwgDco5+v8nEYmJrajyeMLgyvps7y4JfwSZA
C66VdtBM9V2p7tUBL8zkCqMz8T+Kj02+ImxfQ8g2drtg7fM/xQm5LJmOzTwbd+3H
wvlJALAr4Yncf0ersRLvzJeBg/T6NnaoqRe/dtFuRetz1YEJpNIW23da46jCBwen
np5Q0z5UPwAtvqqNPLetEsy+J3YE5cfFC69SJy/+9+n2jPECkeltINzRSSvXAeM7
1rotHjRi27JhbRjdYjhstx/nvx1WT/er8F7VFMBvBbfgDKZCLJ1Unze3WAaR3O2+
qSrUQ4czar8fqxoIlMcYvTiVUYI0eTL9Ia665NWrMxLp6BxXFtjMBP92T5I1sWTm
5UR6mCTAs8boh0qIRZZLHp/8lJ4woqLEz36wSLZcjaEJPPtC94yHN72WJnZxzfDd
LL5lrG30LuuWcMzxKxFftgTJT00qU4ddUXewvXWRBSMqnLhwhEvlA66U3pib/sKX
2O3kTLNrVK093IfdoQ4LjqIMoYREzfFK++VGMdsqvyjdvPHn9z8oSVh/q7BPNqxf
XAmVhnbGsinTkkS3zgNJkRMwrcbEUJ5hMJOkeFIyhdbWygG+s7F5HmL1KiHsD42a
OB2espbv4VzfBv3V8x0oYHhrwzITSbLieiwnSF3IoybLmauM4vcxXF+eBI1mFGU0
X2aiGbbYFcxRQhlyVu/1eKmfh7pMFI3reoBqG5euoXsJ0JRbhrhVBUwZMiDi6C6e
jG2r7+/pyrSv3fhHTpJTE/O5LCKHZHCgAaKhaqMVU+R8W47XxGH5eUi8zVtGxU3I
ufbyRTzu3SUd3+LVhPXSew7x6Qz5PCQCsTS+ZccpWGAc01mwe2tbIYG0xrjhHsPI
XQSxoySbH607N1P0n5XboR/QdxaMCNdP9qfEl7nxkYp0tq/szs1/bLid+zlU4JrI
BbyrjRD8+jEz7urCL1r+JYzjLIZ2+TVavNZNsFKX9y9628sqtoHlSrypJ3rJ8qtv
wRhJDzYvQ1JUOuWqGCl8s+VMUGeTZCWNdnGtojgutLKSGZxJovHTWPKZ7hoMf7D4
KFHaaqB0cQT9PfDIZ/7h98FwW/2szXucMb1Dn3O8qNjUOVIhyMD8+u/ZDe7LTaN/
hCtfopGlS356H4unCjq0kEsYFGQoBkq9Fyu1zAJ96DJcXmDa1kV+GKUcwosGau+d
p2s9SJfOzkoz0aTPDeejBlKs4/12naxq0yxc/whyIaF0dZP7TfWUl1ivhyXH1Rpb
2FK55+lBZWEDXumkeUlFLVwRnVdm4bwJGgtqE1Y31lspavmDJtwps0kfTe651qhI
8M5z66twAt7+373LqXFMbu4juTaY1v8z+M2dse41E9pDcp2DQqD/20IooUR+1gVY
vaUYjIpR2vJBK+g3aybv9FstMHmiuZMO4RIrg9wtzClJ+MkqXb5jpQtCQlt3/we3
PopfM3ZTz1vuwZrr2ExL0Tgcb7EtMN1LDQqEDzDR7YEymqceqyUaa/+HAbOulP8N
T87Rb2ZrY8KwBGh3WT69rqdX2pjGYyRU2RqqL+p1cGI0SKnVoUfvlbUG5qnHVQZU
5O8HDdoriHU4QfjOLOKwjUQty0FxbE/S92ctv3wldEcHo0+BvCDoIJ7UypjkbsOD
rYQvrFdbHt3XwryRm3tuTU0wqkHSSH4QI1364Uwm9ilMEY865+xaUopUXLAib+2f
fQXcO8G2+MSaz11Dme25/FvFlA9QgV3fzUrM/nSGEHxJuRGRvHvIGs0+dyiMC6GY
LJGk6w4sCsy563trU+XjEs7pG7e/deq+7FcfnngF1OhFhsyUjfginwdd7L9XxWD7
DkU6kdRVUftYz7Ezae/NrMWBABa8NgIoB8hClJkQWSPE/gqmw7pT20yN8CebZzsX
s5CZ6RxwfKT3oh3PuKiU05tb16DdLao6x5WNouKqZ+U0VgItsdsRcys6+I5od+G1
cwPcaADJSF2+suhpRSBeK395ipNCJzZhAvLfdOl8p6Rxn54cWlxcg67sjJr1rYXZ
vuZrcKiogp3HTIg8m0iISJ4Qg/VqJP7EW5fXEJI1xK3I1qCgxGF72hza6CZ9HoFU
lbKXrI5vmsRVLiX2TRF4tAf7klSMAGWzqTHxAi8mbYS6r8rRhyfpGneylnjNFvZ/
vac3a0VDoEZpWy/pX7AhRCsLe9I9oVXwpC42o7wQkLo5K8vfB+PAEft3u4XjtWoU
/BQx7as20NrWmW0KL2SO9+8Urq2ySHNQ4Sc2gzZalV+OPZpUMmF0lwvhb7bYRXz5
BRRHhfE7jOBLrkxc4sXLwRlRyHgOpWj8i9NnmZkXyOmAQZjjMwdjSEq7jzci+3Db
3v4k0wZh4tA4RP2CCnnxM/j5G1qnyRTL3vRcCtsRtO6utEkGC8meT/mULoQR0PGc
ZEnZySeRBoDAv9O9OtbJ3dG3j2HX9Ay6qw0udMMiEa8aVi4ftW9FsTE3FaM63eST
C3X4WOAxQp/XKEL+aZlc9I9z0a127TLZEieZj7spN0vRNXgik0ivHNxGdKmfD36N
BPHwGllZ/eBk5pS2Zd1BMeBCYGwdx09u8rbTCMO+dh9/GlLbPJupH/K29Wpbrp9O
qcWmagGn7xh58BojIVDjbCsxOzKk94HCL2JpprVpj8tz4OuJtkzcp/iw6/WRgVyg
qhCcRb9vDZXf4C+58YbiqhcX90twLaM/I15115xfHeMwvFr9D7jjQ5TLKQF6jQJr
kX02T6/TJEeQM4jUopUzoX+OsbYCX7XoXyoOX/erZ3xJz+NU9GjS/9Ju4I48z9IJ
/CYpyYlr7y7nB8QUw+sjDCpZQKKpc7pfYzUyvweTd1kgzSCcz+hIxaVIkLvSaG9a
t22jKvqQPdVMsGKWHRJH7A1ks0LrBBuh0fVnwHWeBIZlkoVcdhFPBM11vIkv3zAc
/JFuz5SFmBC72EKnFsGFsiXE2+EDlWpJxLXPUTqeC0otY/Oae4cx4bDjQvOnR1nz
MYrxZIaFGtW1bs0UFnyNXTt26B8vKlE5F070nUwwAdCYHCcnIWku4WubFuVi4T/H
MKNPJ0q1Ij7mWMZynJtxiP1cfuCeKDK74sSFozuKsjh5Hsz4puYIONf4ybzqwhAu
qzGr7M1OLg9P7TwnfGO/7dJVJwJbcDzcPK88c+1rgYxmGo3xUXwgyyxlY82XyKOC
jNp5+KrupdwFsq7VJazvu+HGGptMy2UdbYsDmNkhhmiYQgnlXL2uFC0cuw3zlYgx
nOyKKtRDnFlP53s90aiSyfyp5/uHZlW/XU01M4lbr4Xxqkye1Kib77vKMscz8yxa
jWpSMgHtw+LcARKGHUTp2Lwnazl9kEN6GFUx4BW7SoRoYuXYsc52gy72tVVtaNXx
WBmxQGm7uMpcDvTXdACOyQn2k59gcciYeS429Cu/czE82BR9PF+kr542WocHo1MJ
Wcxk5Y1MMEVrbLPYYWnlReUnlz0XacTW9bvkpvffwrmUebxj+yr5hVBDZO967Vib
oUvUaUGDU7foUaXQk97c187fEVj5Pim7Rhl7+Q7BbnrvuqILa1XTfd0vhzggLR8S
LgdI8/urCWPpcy+61eODRV7TklrdEHOFlm1Jh4IdY7ecb+DNzJi06FKEbEv7yxb6
EhwWDhQvwBSx8gjJmp5Ke1UL6cXe1lGycuDdxn+xol+ywUr2/OAe5fOoj6wAApAf
XI+rHUIeSVITBAhDjrru/ftMfzdXhPxP+loc9aiGZeqyPGaR0SF3nQAhq3/BqkAm
sVDmyeklNmn6IY3fyjgYcfUl3NadUSWNhkZzHQ9A9RxgsNFF2rwinK5Cal5ccUK7
qKdsUwFxW1M1aBBftyMjahNvrjgqFJB4UMSz30ojQqd5qamCidJc8Ds8pXSMSsFB
RQlQop6cWU7jPbnX7WQFHdeHvYnkswND7ezBEI8jvpD4iXexI9IDM7WdJcp49Kq6
m8I6MTsa8/3XKBmWVvuvweeGdCEfyJt6TK7rUTI2sYBgKIVyqA5T43alyIpLkODX
O5sMfSla6vGYbez8l7Pw7KLKRvzOSCgHlSs7SApB6KuBpIEEt3HmQbU4+O+PVqZe
61lrcIDCRQvinCW5XxsqGp5m3A0hKmPUcSM20g4/NxfL9aYxD943Vm9EhajBdAO1
8+mJotTrFb0FyKxPEul4WHisSpIE4nO8/NM3zNvM21ACREeckBqHlXS5Xq3U1ZrA
ciIRo7S2034yC7GMsPC+OeEGu6243jtkc4U/Cqc0foADb/Ii1Cb8NpnfMJcP9uvE
20D/AwPkL2Qrdr55Mn1Noo2xCk3d7X4DpL5z2TmnjL8jSPNvhiG1aHIqmnXJHDoj
noPNV/Y3Ro9coD2dFqXpm3LITi/MeuNjv1aKYI5ut/yQFYHBS/0rS9eA8fKvwArr
6RMzS3FZfCc5ymi5bXvdFceglBT5/oG2Tdns1jLO2NZRMxaLjr8pv4AxSWzYYFq2
h94IOB5VmY1zIfmMXoNZppoyB6GptKMu2rZDdYyr6OY74bLzbVGyA98joRzChZih
qt1+3iud3cPP2+Zo4o9nPmcTUpQvsL19r97eqbcob1MaNYonkVYRAWXJ/afkX6+O
T8X/rgJLkQ5H0WZh0/rCFB4UJDb5/nNV8fDBLBJ0ywkjQKFyYAfa34L9VF+CtIHR
YKgwk58mgKg609h9ldiniOYJCCz9aB54OjziprEAi/oBIuSH8Le/hqdLQTLfVZyj
b3D+BDbtiYOmp52kZMy73jY9eCx7DcEtWR0G7lFXv1jX4IGf3SSjqzAWjElvv+4G
ideUwS+fq/hhokgGTvP3Brb4TencZMYBe1qLsPQIWJOGkycEP1QypP4UKB3Ldbei
bSKxmOkL/Zx+nLjOfCLKX/ibJO7sqBKqit5j9dFaryRLVyb7j+nIjHi8qFVxnSsP
d+DRC1QQd9Evpo+RnLcvXijYtD67t73ckEqmGz35+1UAes0i7RDv/d4HIiUh3wKE
fKwI3iCBRM7GzaR0kcRQ/HR0GLCYepcGd5K2CuEe+v4YgZO0S45cihXtzIfEVmX6
1N0TD5pfQE1whNf9MQlOmlq2Z2aFUiIR8LC/m6oaA+IHbZZA1ClygbQq0YeXNwEl
Q08saQ3ckaO3QBPSPAJt/ERWyOcZz14Fj2QEuEmxopaBpCWTMXWVapw2o1YgrTx2
KzMg/RJWxUiZr0iUqnne6JwnwHykT3+rwai0SRQ7ft/c1Q+YbHQnujEg5wdmPRM9
JYFr6TSK1sfIphzF5a7F9nUuw1NP6h+/0BRCvtAPEt0ks7BsyNxkw7iGrO2g4ejj
02eOLcZEzoS+bmDduQdcUPyMRfGfRnXIvSU5sfdE1GrgnWpzpgwustgv/vVyDd49
mvHEJkZKL1/xPg2tdk0TpTlKNwDk6XvIpx8h9in68u7Ni9i15LBJKHzRLxff+ni+
0GTMPDvlALnl/WHTdh9kHGh46L6L1DleBbWy2EEs9NvoAusezcoUAn1G+7al4wK/
hZ7dApAZmpQQCNiP/vMNiGQ9gW/GN8JkG1kU2rV57VH+5Iojpo+9WmU+eQt1Q9+d
PCSeGQe4P2cMU/Ha2BKUzs8AbvE5e6VO7yL73SZel3Tq2+vMG/0utJjqaeQMnQzl
gBmPwddtEwp5jl3KxpigkUKHLynLmaJXc8+jO4Ye7NoRQZ0a3qzCcUcCTe/HbAq0
5+8JB4rVIJWu+hKEQjBZZ0blxCdr4lpVGolxRvSz3aYy9PiOLAeOLwt5s0l87X7H
j/47SBoMTzpRC87HaqSvRFGcTDcw/G7ZOFSNAd7b48HuI5i0FqMYS3QCl7G83uK1
ph7eI5vtCW2EDStE02DENP3CRatoBjmQwuPby838WJ0D1qQDgt9hV21OWKHI4Vjq
CCUubnQl88T65MV1mjTIdpWkUeDzJdgovQaCwnh33fbEg0qOoZ7NE1C3/AxK3Lkn
RFSa/WrMPNBli35XRzEsNEca6vF0vYk7wAD6ktUfCJQ0sbQi8X99bCBlfU82dsSZ
d0JiU1sOAOlxeUt1YTsjRuift38VzfnzCvooW2zoqzxlDGGw/X0Y1nx0FG5DNoL7
xR0YXeDU2O+xdubG9jCYhrS/j2lM++qpmER0dOAaRNMTi9NkXBRKN54KBH3EtHW9
PlefWiqytFGf8hxparpY543HqJpxI/ak2fCm4QH1NAlPi/07/3QT3UHp6DIV6+2d
+yVUz+ctvcOLLQiythIWThMyDV4NVmTMTk2ZWyd3TDbLvt2btdSsa6R8aNkUNWZc
8SmphmqC3SEWQustRusC/SRFhEwduJCWRcXb8AwoCHAPXkVHi1+y6qH65hQYVFto
7cscGclZNlp8l86zpk47twZ5PZKBjin8AJ65W/6nE/WD/jWQyISO+YKYvFVxlZK/
7hjlY3GqVXA5igj2+b0xsJtW0xlo54wVSm+XsxkK4uy4gdgCuzxzXeW4iK3s+4Vh
OLS3Pt9xW5kjmk3wr0tWCiemV0Bad4QgFZLTTbU7sy9OiphLHepiCdZGe0psv74P
Z5KgrBDwaGvHN2NUxSFnvePx9oPy5VKDVmcQEQtZ9j6HEjRbA6zHl7GQPw9uY1S8
q79srcYsC4YDMBIs5EBOe+IRNjd+jfeAn22TWeSoa96muLX9bD3wFwN8F3yei+U+
wWu1PNb4QiCSGc07+HqoaMiMFDTXH6J/dAktMK3Rjcisbtpx09vfiEznZeaF+CqV
22Fe1fq3zhTgjK2x6ljtsVNAmGNC6lU5JdrXz6Rw4lj16Ep1VUhBTs7T/k+EjaPx
kmIS5mNO8e+TA3W4tkOzzRCydXToIT0hjQRkBtdEsBtek7O/nW6SOJnaxoAKmM+2
IkQHpaSWw71Xdx5B0inzPgDzeX7npUnx6LFEyozj3pjoaqKfqGlhkigByquU7Ah/
D774+Uq7U1oLLtYn5nAILLyK0zlcPg5kHo2LL8jh0Ajip9L+PfaNht328QyOhm03
zF25IBVtpAW2TF+DiJ34nQU5gTL39Y9xLsVCe3JqOYtM/dJQ51QmW0Y1moeuH4aA
IBkclQwrnCi2HPBN+kYue4YvDY/x4hwgnMaf9QPt2S9os5ZVW0dTqIzwKj4FPFsA
LuYVlVtCXxCkG0sG3N4fux5FWAhzu+zd5vqgof9k3nTlqj0CyheHwQe6o8VEGNSS
wDm6LirxZrB8z6RWAemt8pR3ao/KFm00ucLlryrpU+aZuiTpV23Wnb6ulohKL+Hc
3Qcsv8KukfhanN8hNwolZtKYxz+P7OmVgiJ1qFcMX7TuM3J5/WqUn93IuUsVGEiz
uSr1uJ55c/qprnEkpb5YMb1irizUisWYsT4BpvCJAjurk2ykQwFYBOtTN4JwzAnA
hr5YXA2WGS2NUS+BM+kdx9cNbeKNefCnJoZUoPNA9utM29lhH/hPCF7FXYteD7Eg
Gzxo8qR6LWMzcWpdAMhXXGwqSsKuk4zyxi8wD9btg02aB/3qDwwDhRzriN2j56Mr
zls3asikvy/pxguMISHbrKCXLi1Pgh4EUggNdG+sch9c+XipNqiWHWp6cWNDDAX+
XAsrbbqDVJ68meZEKMie9gWG8zWmo6A4/hP2xIu/ogLDt72oKc8v6qDiQIKkAeQb
ZF9T5xzjKn4XTzNRBK6tdGJqFVSCLN7JiBFu8xYq/AOqpYAPL9F8w8Ny68Us1Ud6
CKg+b0x6AHIHG9gT5tqj50XkQn1SuM/H+h1fSa8Kr5zlIeFw6zmaSXAH0vp/Nf2M
YBI6T4QtvhaE3GVX6b8l2aD2d1BPdOiTdltLAZx6k3JySKLD3N4JaRnpg4wlUJZD
k+AYc3WSt1LKDlv7lM3ia6d5wSqP7Pm50LRDh73Cvy3JdK2x4JaaEZ90ba6yfjWO
l9VVROp5NEjew5eA1oMKXHvy7Kzd1Zc1PORmt0H8H8O6ib4MR8V1at/jyWRwSsei
pc2Rs9uk9U18ZsSBMOLWDmGPZ/509IR7rlxDvrPSe0CpYS3WBkBjUZg7MPXhkSbc
RA5vOeIXoxIyG1CU3VsbwKdNDIgLRR5rfqCOF9Xi4cIvb9gTv7v9Ace+cHlvxCYl
AbnSrKI3O+UHETjLdEDuXiNXSw23yCdJAX8cmQJ4T6kw3pxFtn3GmhVgMquhiFSe
GL87jWghQb/K4flQxHBvh6Or+d5aLrJKc7f/CrEMgAk4TA20ptKOji0uiDoj9ncs
GAGvZoIfEwkpAj6V/L5DowLu5rIQic47F+hfDkNlMZsiZLZvN9zcj5RnjgtlPVzg
Dv/eTJX78Rsn6cG72A5QEijlA4E/aysDjSxAogey1Hqiu1Imr4gIxFKzs3jgaqh7
qjTDdyJthycbkIw1kOqGpZuZwwNOD+z3nuuae/pCHqigoptr+TB1Vg1u0AoZD1Ee
nZ2T1NNLUHfYBZY0taEYBJbM3S1drAGZycMeq/Q2a+gFnKic71rUZ6k2L7+Z732y
MDWEffIqrH6WKCaFb+jjmRoa2/QNQNhNkMuylt+yKZqX/U661n90Ij4k74/qBndg
oJs++TfWQsMlqIJwxaVYevOzCAeaeFETkFt5XwuuyDxxKghInn4TPpc2yNPfEgAR
bNo19dZQ30rjOUo38tVRzJZXiGQ1sSx0XwbCPXBoQt8BRyRYM4n4ei48lp7eGIIU
uQgchxPAoQojdd5IdSE+Yh17VEf/h2YVEnQxUeszY6WF/XykktEMVQPn7hqt94vu
EWtXCfgHws2uFp/klH5rHXMgLD4/IDcqQlGWifuMmiIjNKQpFXe7m4QlCp+WEqzD
BEHKl0zYtMTUp1n9uX6r7dYgby6O2NOIHaoQiPNLD4mEZVTVGbTalMYT5DWjfF6R
PgtEwJlDi1VRNk1qa6Ebuwm3X3BJA/addPZfqTwnUerYm2PmyM/Ik6nc4tUl+q2b
3Ay8Bjb9GbGejj6eyEMTQ3lPxKr5ss2GSeGvvz38WtcABIH9THgRFhxL1MYH3Ugl
pvxoFzhv3mz9YGyCodysX/uygMBj9U8Q4upcz1q8p2t7+Pr0d3IJ/yXrksW/yCH5
wT1bvbY1EgSbn7ic5TGyH92B/K4DT857c2AJ6zfHbkGJBN9aTxqvUDtSbI7LvLy0
035l5YIBeHfnm5znCyPvdEde8B+YMZOaGgy1wDpXuK963pQdnhCH9ZrmEhNXX4NX
oYiRnMUzjh/E3un6WD0oa7XPm4l6lF0muulJki5O/DCBcfQtmmYvTWXoDELjbPOb
ghV+TAXsudJVWk7I6oTpnYcZyr4qxoZoU18c7ra1ygE+dFlNbmBzMQZMCLLDQzhg
mMr7jAuAjzX7Emc29FobYiUtnPDkGkHx9rtwTzGWvqRzCQckkqzcAw6C5bRAzJxU
g6ZpuccjAohmAvUmiDAD5mdU4g4a2oQ/i4tNPsvFhzGFsXfQFHkkDQUXca2OhZF5
Oj+Ar7PbFwgko+vjrx0yc62b4O314LEaqthlHwlFG3n4QNiCVBLOPC0WXZKsrqhq
y7p1QhiaSvhGmJKXMoCvN4oyPxMzNkspNRQ7NCceXAhs+pwSs4YtSuIAaimFAbYW
91i4E3rwt1T4w8BqiO+N19j+aSxKkfeZ6Mv5910VVlxL2e8CmESUEtVvpQ8tUVyk
Lu3THe4iZnhcgu3ktUtjTqXUpciC5kxFUgLMEQejeMVsmwdyxFR+PlgJMhAoMwQ6
mzZb4+NIMNp4LdBQadyI9rPdYHXSwA0+eaDDTSNsHSnLE89qyIdpHp+JGUlFPGh1
ddwz9+xX1LdfAvBsE3YoVt0mmwwUl3+YsQ8jk0+byX7NPshTyOv94A/Og0I9f5mH
xAevNBXmaf4FeUm3P1cqM24JBRauijRGaabrPXmB+x4o627MCL1tuNXAC1vYxS2e
eRW4hTnDSBl54DZ3aIyXE+BZXUwYKe2i+YFUlf6baGjqvGdZaXVJ6FLfZHfuYAzk
thclCAMo5JEaFhsMV1eqTZOoAHAKA9LI3Da7c+tNQIbPWshkCXzRYHU+LNvujnVU
xtp0K6ZcEAqCjI1uJS7b9gzmuueGLFJmaWyRyY54dt5QpeSKUycVRyvF4JrOEq4v
4MpMKc0AhGAwjixEs61AcbU1Lt2cudm3xhRDZcRny/5rgkKjqB82YeaRytLSp17s
lwpfjSCRBAZADQh7UT+5O/7Yl2YYlPQdN705TQRAPCKmgP8yfLghm5Wtpeu31ddY
HIOWL57C+xcz1i2I2nLWRM7tFVBnMwXvroqfw10Rcw22QiDhLoG2XDNrrjQURbvG
lW+Q08UwAUuGErK6I8MA7Q==
`protect END_PROTECTED
