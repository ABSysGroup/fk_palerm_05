`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HNKkPosRXY2jckAzTae+BQ7AG/f6ShN2XhI/o0zzDKrOXmFQ2h951hUAJn9JdMqh
SYOJG2CpT90avOZhY2yQhHVR+HQdu9bBD0aRpesqgrdc/MQBlVA8MYkDmm1CvOtM
laUkmsZWk7i7EA4R16rRv3UQfslTrlxXRmhuh32rDK52lC2vw48TqPZObS/G0dtK
RzlZRlv+FSxfVPFYTghWsG8U8kozPiYEm68QNQO+ArS59xLBTMv1FPzObgo/yHji
XKDT50R36F8l6gwkCFxRiWlTvZbmUNkpj6lzzofxoNbBhqZbSM0tAsJJ4G55wsM7
MTQMU94toGdKJJ857dXpDaWrLTF9d0Tsw0mOF6c+o4TypFJmV3hD8uUFc/63hYw9
As7FL4Txabq3RIA2qT5plXp9A3XbpFEZtQY9VZoKdr+W5iCxuYq+gWe5qHDGMjyF
mcgndtiWSUQT6KjBozhbCpwE+F3s+3vtTg+jxRqIhdg+0GVv5x/au8FmhwqYv/vR
hGhcm+BK9t2x2Tb5tFUrHSeAVT14QETFY6jf/FLgTbp3BwGaNH/dxCtOWuaB+2Bk
pOWoo9G1mQR55xuOjUbLvV2cKFuhLytkduKqrK1pQrA=
`protect END_PROTECTED
