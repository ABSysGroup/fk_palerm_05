`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o53/d5XAtkpQtxyCmqpSjmjBV+kkjjXQX/78cYg9eabouZdSgDFTx/C8UUaQLovs
uKYZqu0kvDvMjDjvEL7ITXCPOq8MJh6ubnTtl/Tq2C8G3a9y6iamm+nGk4ZmvuHo
CsKhG8TcDtR7g4VEmEqZul+HmyBOz0mlP6pXFHTHeJqSZfQYCmkXnzhKCfgQ3yMA
nrSU6X//X7a4B66y5ebGlI7YzQhMvmGr5fi8Xtym4ZcAzoEsmFO1gp7V11+nQA5l
ThYOi9IBofpbD6sUWn2HmPLurdwbkflIWvJeh5l/Cf/u2Ac3u+vOlQui8AmgappN
Ok929gqI1qlx1gK9bXnmuVDWtRLXclTlMuzIMENgtGAT/CPf8P6wLDM26TArcaxc
vQWVrjpYcNcYxOIQBxYVpuP2XfgGmX3l92vjraR/96JvTOZUTMCT/iMZb+gTqKFt
2IEouyh9KK52MtuBKouWNfLft5gpwqiLWntYL8+6AbsO4zhN9iA02aK7b7ylYWio
LDE7CHLknBqsgqm8XzZwXYXuQjkYVrPvEUJ58R0Lz+8ZC0fCNc5dQbz4qJhDp+FQ
LC7PFs9FX7jeTdvKZ2+bYSu3Ca7ty7HqyhS9HG7cBt5tvwVfvlZWP57kzDX9IsNO
d4TJj78f5XlBHnF9dhbdQtliC/joQL0d6cMdgmZRS+HlCfTFpgEh1Ahepvlprmnf
MZvi7YelZNFe4TFzB23jXp1sh+K93vIDIs1Bi5i76jnoVYgfrrW23UPZb/ZCI7NY
c0PKz6jNEGl8cNKMhfqkTz5kr0Nvdz8zI1z26Yd+V3OdIobhJsQBiMt3mip0l9wd
WajyNzqATochRWL2sF+ipSewIzzfO+paa4elQcnySCeMQOM7/uzpkCl+Phdk3Hon
CmFo00CxyAs3+k2Yeq0pVjKLs3T6Hzlsujt6ntwG1lE=
`protect END_PROTECTED
