`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cVXDBDiS3NrHlRcQE/LZTkXTuungV90LqBjWdEbeZmor9yo3L0lqYKGiG7RpPJPc
4nIQfiK96Gb3ce4Jsled5MMmPHGf66Jh297EwT64fyioRk5UQcI4qBYiP9mPGr0i
DZtTUKawm62P1freyFTVQBfm9V5yWk3O0esyg2ndpj/JaMuxNYBN481qJaKbIO8u
vqe1LFhQ6S16ECk3cuO8kMij+IGV1AvhHY6aXb3SmT1TmGkgLU89JXaDsDOt62iP
ijvj12kSH9o1Al1HACKuP5CS+5AkLAcSUu0ULAiH6JV70bAgXZx8/2TNQxmr1cag
5JP8mMLm564S9lAwcE0gG9Eon9ZNgNmDlN48ILrenZanSSSQwyRF/jvaPnFsE4vD
9kIIJv4qRVPNCTBKWkaJ7xON0BntCYHT3DXgHOYiykL+Y/DdQ1YZ1mhJI6zNbAnH
5ADJBPcO1M12dlPq8TXRp2trfpIYjQwbyw7VFMltEr4GiAoyZOpShC59VUsivYQ7
kpUvywClEdZIKLKXytKTetkea+Pez1Mri9211XiWV9KZhA7cZ4rJvvjyBV4AGEx6
zzQQqpxXeXwHZD5rovQ94dYhIHFlNS8swKnPhBDnpXakz8fhRfS+QF4cjZovUR41
6V3wkuKvZ+EAK96R6oC3g3jS2F2cH/W8BVvqvK+KmXlxT66RSEp9x20SEssHqjbe
nZnvFmxzSVi9zp78ZECmpBp5SXCINaCM51ErYhKCHNRDZbzUXzLqLppLpmeIsVOu
brIpY79iIiTX7yIeoMV08FYt+VbKA+bfwOt7BuhKha4V7/+OdGvLhFzJm2iGA/1f
6zBk2FMOX3DtZoe7xXKzm4+LXFAnRo7kGHbjJfRFcNA6L9SjW4PICVPSKZRtzlWk
/QlKx42q2Q/zmzH3J7koxrivU6bSWnnQ165YzC46em9T58fDtP9PZUzuXBy30IFL
zt7azFmqXIqdls//IOtFU+4uD5au68BfYhFfSfdt+xB0Nt8gU3M39qpvTWPBPG80
IWF7fwpShRxyGb3fGrAVVoCO3A36M6jeKCHNsKMDm9HEKFQ9Hh8S/YiYdFXh43Ne
g5j0J6NhR6WD7F+0txwMH5g3caSteqCE3y/z9ZbqalCC+suLSo0X0LBhjAypGneM
UP8m8/0afBRQUfbSog/LHBmyxdR8ol/6P5pFfu76nYpZ6nCp2185RZwgTi+e0jzy
lTFxGnDC7XjRGvo5iYA21JK3umfuBRbQqIGSaoiUMh24sBGMcPvzZZlqlfv/HW1O
IU/927FgPdqcyvAQxD8qyUJpqybcIfXfXAIR37uU14PhDy5MXOaGa0TGBP7ncyhP
MXr+Wbs3Ct+v20y9AV69mdHJvEvd4O4rjXJ02eXS6L05AtQfK/BKVhx9v8rVZrGI
n+c5pUqnN+bmmsx4W1kudaHufX2kBcHzHK88LZQqhvQBgrpGq+VCOeIm2eMC15P6
SyPdRWBctypEXAzErbik39aU9nNpMulszMYRgw5I9CgyjExqBwXfJDado4nkr3Z0
lqc1sTrKCq3V3KNvITUF3WBrvQUzuIY8YkZrxKIghkVsmrweRYI5ONoATWsyCe9R
0P0riXxmKCtBNzNANy1aXo51Wd+5x/BDjIdLuoP5Yes9jMzEvsFWJmwBr+nYKL2Z
ylALVeLPj1KYDzkm99KCcAU5RA2aYqVmda/TLGS8LbwEE2z/atU4jiiWcZTbEgNO
0Uq6e8h4tv1A+hEkcxDzHltNB2f1nQ2Bz6FCjkwSGnKWBycFLyme48z5IPl/9fT4
fbCbgqcLF4OSvCmBsZLpIQiQ5XA3AhQHblK56aD3K/8ZPa4ser3FaSfiN8J7BOfc
EIpIJkd7EHvIZ63/UiUrlbqEuk+fItV9d1hvgCS7ie35momLEhpJBeVoV0kIYIeg
zIQdZQVO1WLuxk1yMMWqYgnlHNLggzM3SmkDc4CxPGNtNSAdnRp7qlNQIAiI++Om
ZI9mEjaKX+xaYrqivtzCy+TR8/ighpNs59zeTHl1vBlzRnph1QLyKAfA48r2zePk
NIe5UyoEHW47BNefxcTg5MXRlQLmr4JWeIj802ELS3Uh0AaWy/L8hosjfSTbilTn
XpUlsa7rD+r4Z76kM4Cga3sklrR7R741ec3GSmPAbtVy6gYRoY2K6g1ECvOLsj2F
SAC0JPTY8Ynk9mclJImeqU9TMKq6bN+gpg7b/iaSZx54z8048jMKaHYnFdEX+epf
hnHTB+ioZ32w03TUjq4UDCPDzWQUFKgEwfKdf1DGOgcVKxaj4KWbRveDG8FgSb0E
SRjIjnWvA4+Mvsd+3o5PlCJTS2G0weV/2ReummHVxWL1Gw4VYa5f+FlXqYZCHtSh
y7IiiufuqoKg4wDEAcAIaLaDT+tNXM5BHnFFbM1hPqfaPTjN6L3+IvuUqmUW9rZJ
A3+i1LVaZ8aZNIOoq73Ld9lrhFE5YxUFLCHVAz67N84sbmtxWQBYhQ80vatIztXb
6xG34JtBzUUQE9rJU/gHJmqszGWFFU07RsZnKi+HWj7FRWv/IMqDpXv8jcwTV8rK
DtloDsjopJPHw+7n3M9LVsOdwisUr2k1YDXpUpekPlEUt5YghofBzfONSA2OqLpj
fnKse8EVwY3ki3bKoaMoJF6yg0kyv1A3OPdHW4kCcl+SK4lXlWimBCkqQVNK4nWe
bn6GWIYk6OaaL/gVQICxhu4JgZWLTrNmAqGpMnBVrosJ3Tr484VgHIM21c6O/zGR
Okdkk7Fu8PhL7oOUk6A2DdsTY2Hj4l6pjqmHE/7CB61344mtcPZxBbwXS3mjF1Db
VAKKrwC5c/hpBceJeimojmov00BYf7grdQ9cLfjB0vTT/2yRz+9lD2jLuv9Ej3uV
b/UZFDiV+FwYp6oESfnzNh6aqNdXhHDatCneq6T4bqEWGPCVrq+F97TI94mfe/th
fbwsBq2j1RyIaJs/DkSQe9ZWXVka6c66C9n8EHJ/lcwf0rtNjr85BkhNEv2klOQV
ccLEx+bxaL3Cj65gFgThZiOwz42U2V4DMMcQn/en4iMpONhbLSZL7M2uiIuN2PzM
4Vo4T7CJlhxMyb0qg75A8rTDpurHcSkbQGzwo92WoY+wywm83a3h1wY3h/jDZCDT
6pMHJgAAeewu+/POSvaY1gOE8Ke4QAU6aaX6KIuIWf0lkYIlTOFlpRGC+AiYLkcA
eiSUu94YRiJhNyGhO4eQYJukv3z5Ex7dGDHahk+RzSNP1qQ3IGZhhvY2uvK0at3O
mP3GK3oAIqc322RCpSQgLTZWCAw4TJqRkwUulNKFduVRiJbqMrBUsbSA1YQMYVIO
0PzbzwK4bbp+51JqFu4bXc7WT6Nfz56DhFe4dyf+tmmrn6BQGiM0uaQFft3lupVD
v7Rg6eq5UT84aCjAjccYoU3l4zwTe0BoCOQAbUkLC3LdgBmlG23eJ7tGtwHNoiw8
AxdKFDDumEjMihfs8rw6AmmKkb2rmZwMOWrM4jEUNrGBjkTsIjJVLHvoJ/qt4KlK
yqz9DzDl7gGh32bxYh0L8xP3zt7kUsdZD/DwdUXZ2ftKSZoSF0DygZRU3o6kk65F
OSEJ/MqhJujKa0/Zbpp/xlMddT8NDShJWgOF51b1PAxqdQ0atubZq8JmlzpEqdrn
MmOXqOohDzoQoehsxlmi41lCGuVOwnDNjYUuQVnTSSTxMDV8r6VF/bxYf4IV4JQH
vr3NmhFFCXkTDk7GWSLqZCgbcmSQb/zBYzPjpjL0HvGUFu36byRHB7QkxtJuaJfW
QYQyGQMOXB6cf/kBpsgOPSSodERSZILXAaOq1UzuoB5+tFmOpYoLVRv1Hz0Bvexk
UCqW0N5jRFK5XiZ1hwxYChFXXiwOuoPjNSwWzrzJ2otabImDny2X3dnr2rnvzQg0
NLJoR3CPmpb7hfvSo6kVdAGEYX1uyITcqeeJcx5ZUkchXExi6zLliJAg0L8tGaQm
1xhIdAofyYr5QihzPMfh0bJGmqMDH9FFyQzezq/+vz22YqIpOu9tGprzELjAOWeK
781PSQqfwYtLSFJDqBIcx7CFkPo+V7e3AIKftu9D4qOG/q2F8vPXM7dvaL1jjeIu
FJt0oWh7QmaM+kMycBDloiHD2hy359VUpPzI3cB82nLEoBfsETSCTUY6YDc5ljwu
6z/K020W+nw1+GDkWI8oF3E6D/WOAlTzvxHff7Y0EmfihntL3Z8hYLBbGdokLSKj
xy6kgT2aSIDFac1RnCoXqM/9/y8YGCcZ2igN/xrt3uoYi4mua+NHfa2m5dM5/gjA
G7vaAsinoH+CDs2nvlJyfWtSakchBVgsq7zX5JmTDYJt2kWMWeic97McTd4BazXR
axAGXQnMz7pLND55fVC8+6qrNSmFca5pDH47W+pXYHW1llu5B2bhmYW3N8F1jeq4
RNRlN5grjfyM4oBGDGK+Nfq87OoVgAOL9BGsDB+Apkf6rWtGFUj5uFXz4ZZ8xx8F
tpLphyv1rFkL63NozwQ/QNqBSbQ27Bw02dEnVLSnTjQkXS4o8hmobVlvHeb5tekV
4nVTsX5JiUBQThJQvob1WjNgVw7IqigQYqaSvFvsa2UWYbbWNQbo8X3sj1e+xtC4
jkOW69nc92zv89yEf5CD2OvkhQXcu9X2GVZj32+cy71paqmLODvDbcli8VvAuJ79
m1TC2SHs5/FslKzLIyxRn9myTptaP+wVcSbqATa+LGURE6sdZkOwm8fITh8auvx/
tFCoVwn3btQySZ8U1/t1mIQUDqofVgzA7BtdUGNzxUMmJM5ga0/Q8xYZm8C4ZZzg
QACACGUZ3LOw2g7F+mlBi9H+GLwWsPif9944g8VGCDge7Rra+/SH+tqpW2O4Fblw
tmvzqyKDbdQJ+ExGprjdzILlusYiHjf0dwFRm3GDXHmRHQ5hW3Qh6WQ+8mipduBx
2zjC43gv7yWkJtICbOnBrKlTJkoQ0MatuivlSAkvyKQq7K6Z0gFN7mcchJsNTAw2
03x6BaBqQkedde0eW/ZbKkfqq9p+VDtA3vuMH7i3J4yPSjNJlUw7svziJoHyq0fh
Qv2J6XaVLI67rPAElZMcGXHT3a2aXYZ3rrztZed/cNq82Aw8ABrL1Pi51fk3KJkl
ELmaOLG0hyykZhQR3Yrp2hFN8+RQuq4G+RIuFZH5Q+3z++r6bLn02Y34lkq2PHqz
NLsWqyxNQHYmR8NbWtSnB98whnPVnhV2ecJCneziHq4x5xMRfu+zcXXFrbRVfgdH
hpmriyrG6mzLWZeVv18z/REVUBplXoA/6pLKhCGOFbGy9yIh6qqq0UX3LH/Kcnl/
/FVba+Efgke5+EfaAcl8WRsMd98vWLR0nF4e0p9DrKkwjhWPaHr8tAjk4InQ4b4R
SjlAO/Np7vBH7ZurLScVRXvMHkHX5KAGafzLa9GHGa2miHpTuof/qZO73TtT9jqf
BllCBe6E4C293ecTzZ8UFktzJu7RNubnKeDKmOV2D/oUTUwtwJkm6F4y3dX1Ybm3
cVjHsrjqcmQHTC3dCWwd/MFtgLwyEy8moDaqbT7Gpccz1Y//K45qDXjWRnmoWt1I
yu9YXQTAstH5wQbeEK+vtyGeu71tlpGcLytPhZc1G+kV6wD9o9ebPR7hX262s34b
6FMAA8h2pBmpxOmm89DOH6YNfDucbAN+UZOleG9pEWrSf6gBgAOKCHMfqp8fkVhr
wnC/4WC1COqLf2qFqZ8pqp2S2YQQzdGpt/UmL78xiKVDKa+Qa7QGl7jGGAhij4bH
ezAr774ayx4lgfOgbw7f5q0RShP51XpfYpdRLpd467pkWitBaOGRdPfhkI6WGZMF
Lw/M820XDT5vgw34BnohpNq+IONFdtAML9tei19iX68BYa4tE4JQjmEcspa54D0v
awjjvqs3KssABNvQfkKj7JsouzEeowJkoyJGi4DoGF/9HekajeG0tjxB9WIzJBiH
2KQy7oEyFK5nW2ZmxYmu2jybXi8g3iBt2BeL8xapetL2o8s3qe2R6e2Uh2m3WUlB
uOdVLYO7ICfkU/KbR8ZWl7eqq90FOSQbLGFbozP1JniKnRDKzMy6SpWyOdrmgcor
RKZOpI3vpyJLlgROtY1hY2LyNh9pOqs9RP2I3Icu6Fqgk8XsAnpzKZUtHtu0jJUi
53YuAhm6OcPpW7Ah5BjQPaoC4aw2M9+QxC8XSqvg4vnjpL5CR2oIuouDXHYPaR/C
hqBSjoG4Mx9C9rA55WgU1k1ROD38+oA4SrL4UNCFt7E9odS5TDfc+9B8I0iRuYy0
K16jNM52xBPT3+OtNtwauQHTxm97ZZI2puSc6KUTX/o1iom/+kMGX5qVJqGK/HQU
+5a2xp5rI7/DWI6PkDs9LbvJKOPUOeWjdNdYmDvga6T0VNlF8niLI3+8ZiwoV9Lb
pUtUq/QxbkeFnTADi8jFGpMCP+QzJULnCn95lFu27ypSjYrpqUZREiW+cYwAveAS
ZidrYJ0dIg+2xH6h77oDetISXPDLfWVEZgfOpCcwREBo/yECpxPdch+sMKEGWT+I
VoqxJcl6bWjMF2s5JpIrqxmYMGx5wwmSsp1Dfg5AxqcwxRC7axgDsBrFZSdAkEDP
c6CEUQdbSQIyhO8vk+R6GXc5JCBJC9RFVQ52dGOJIZa9dg2xATlwtXHC0erAPlVb
ed2cpbFVcVeO7RoJ1nIY2k2PNwdXUdNw04y9tWJB9auzNEY5CaNpiWiothTCrblf
hN6P72XS/A+7NXgo827+h2Njv3uQHdwq125I589WJkj+iZTBp1ssy0HnZIYJg4d+
3zW15KqxuHCQACPpZnN04Gv4cMePIop9OnuPb5XCYGQ+bsXFzzfuqVSTUiEr7vy0
vqwtF+cV+lNG3AM4bAnXn7YDcRZxgalEPaW9wFgPoEysnEtnIw0r1RUdBwb17e1b
Zmj1rJHpnSB/6bcRouvo+A==
`protect END_PROTECTED
