`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XiqC+8OhLaNFrkDOIBnJ273hCp51PbpOPOwSBkI4TlIAXTsdnkbrEckMwRtzKl4a
z6cQY7dOPu7nNp6b6xHIGbvaHt3y1JMwnreqoXN4AEEQPYDvvysoApWkuzZ41yMB
3V6MEiX7OgWa12fOaeqdZ796mQWrZB/gM26CrimgEIuBTZRvCJgTa1D/EO0rXkWF
yAyn9o4trkGSE6xp1HLTY0CKxxj6JBa607BwQygtR1ftjTDwkaDNuW/faSQXamvm
CFFHWsAgvF2DQUozV0K0qKvt84gWBIQhX7n7F043/ZaCJxE2eM/AAfZ4MnbhaCoZ
sjQyozIyBOvnIYdqA8UZmf/o0gE/sDhVeRTQDvytQvFzVrhpGiGzJ4j8azPTqOMN
LNt7HF3eZBocElG5FEg9SZyEpghgul/DCHdn7r1rnDwrlKy+HDckJP679lt7hz7V
gKczy/zfD+u/NPe84F13srhvdN6F3xwmB9TZ3u2HWxtZizQ/XnEp/8EcLMbLT/2l
aHeEmdbd/bBE8sMpqTIOPjrm+0ykmP/QbXvxD/boqrt5LGCJq5+wdlSN+PUx2D7E
ervpej+xp7xsKm/apfm+HH4moEOF+K9yeU7glfXqO05iElTSalVnz/9eLOnLDrT8
CqQxTIYWVPmriz9YgzEfaqLrqg6tlzQwL5WNe6rKCIQE4MlRNu1sWQfuTr42IFPO
M0rGDwTazZ10wpZp8DsxuBKhddeZ0dmZc8T43W+4HXZ6D3+avbO5EJU+SDCTUfXN
uBDPSiK/Hlf1VYJmOQkzXTiY+UvO8GdPZCcXtW8I65tKiGLcuUkZN+OKsDnmSvop
e1hjosTTobhCzmNZ3+N++F3o6hCEuRjZv6wpQTUyOurDuC5AtbS9QAJlVGnJZvP3
uXMt8d4FLWZGsfn4quglToex/WfUqiIFNjq91koC3kDyNEFeoktNqsq7Kjw+IHVX
`protect END_PROTECTED
