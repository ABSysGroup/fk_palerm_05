`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Ynig1D8X9OA4WBHn3Kqzd9PkuASmXqoszrfnEPNUz9JIHCC7YRpDFV2fKrOIRhH
nTSiy5zt13+gCveAm/iAtzCjXAQI9cgEZk4zzm+T75rekynHlk+XPvl95cPy5s2q
YE/56a6GdE9YT4YYyFu+oXqti9nNTrL5/r9bzLDJPwDrE3uYR8zcgP679skmBS2O
4aGoV2QT5pTi/1v5LVtjbY5Xjg7SEJqD+R4u5Rm9d8qguEuzSx6IOCnGkAfZmDo0
/yv33FNbkqHsFgrvk14nvKysypWMCVabPU7eaxjC2dez38Yd4LckYMnYJN2N8uVS
qtPK7NCUOhG7BW4Dv0wfONXbHesJQ6FNB24DBZhm6RhrhGBVb/mFlVyw5XoNiRMY
jZUKWYqiWQM/NIUGP5fC6KyDsGWruwGrO9xObutXxZ4=
`protect END_PROTECTED
