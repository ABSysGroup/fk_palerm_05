`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
34shxEg9JVabW2JaJMNTZ66psnYuK/u97BBn7h4LlBbOQGld1SUboZwHNmZhBVB0
XZADib/Z7gRuJLBMqWd9+nDOQEKFGjqBirfk+ks1jrw3kOqZQ8KzytGrjMlRbo3g
E/IWOFIDNGrzXLpdJXZV+EIUJ1x6hK/7t2U9762/C8xi56U00oaMZbxFCrQHl0oO
Z5edZ+8APS1mvhi3FzknO/eNH3Q4wtB3gu7TD90M+G5jp+2Ob/HEvIWTE8kFNExm
wS09T2+IWwxgKbIGXLVgev2GYv2aUHriVm/ZL/Ni3LHuoW4Gq+61sLmXPvUKirfV
nFTyvZFSIR+oQWtXvM97KdjwC1nENjv3siygzeXemrT6EznXGSU0TzSeP/MJdCtN
mWGFye6TffRZbwdQHCaGtZw2tr5oGLYSV0KTNSbLuvBMM3DUM3N8ZB2+QdpLvzPe
QqEb7EZ5LnWH6kbkEDCPrGXqJryLdjurvqekBzZyBgn9N1j/uqBFrZ0GXYPybisC
Z9+jkhIZ2T8isvYl+Whib0RVSD9V/7hkWur4RWl0lrBZc+PQexyXXpdER8nBBR/4
FhMn4+cNLyJfWNlSdkqqEVWaNl5QDLqn9uAAiJKsrm7HMKdU8ErSbPrlrRSDHuin
0ugucPyTWs006NTD2x4wHQBYKmHopXlP+8hylMXESROMZHbRUXFGO/kREH4bs4E4
2eSr4KC2SFZ0rvJKWobSdr9s4/bGM3nw3F+TMH9thuVYJQe+OYwjzoOQyi4+KMJb
f9hhzPGAM+147RCO1KRPN7aoJW3vh5k5HqPcROZNuNTn9DAlIOeNHRwgRWbDAAod
7DcXV/dplwvvlciusnZCF7Dr9/IY0DiJnwLSfoamyF9L0oTQxzXLFAlohj/MhuTJ
apVBfySFwkbvS8QmT9Pw5y7/VGM+/5pw7WZ5y67V7RAoiVScHpbGlxJVQwu1OAyN
n3a8VsGkjC+nBA4J1ZRtSUV8KCqhob7PQ19mqGk9mhkv45O7wEWhx5IjqNT9n+o1
8fmyvEatGM+M+6GsdyFtV4kVFurR0VwxPYVeBD7pnaAxuew2vFzFmqhaOdwv+AZv
VW+9JnsEjTG5OyC1Mn1XyNvgUOF0OAfw6u1fsYaxD1RGzPz/+PyFU1JTr1UBaN5Z
aueX1GQ9f0Kur7TT/rkCJHTuYNMoVkvu1aDcqhPUHZE2F2w9m3+K9gLzIudKAFCJ
CythCCEAuA7I1kZpDZG+wTghXSk189BgBMJxoAmeDv5JAO6VLEQpoIZZYLAPpjmP
IpUJuDCD0W2/6TfvaSjMv88NY5G9NJvxKgsWO1lIvEW298Rmq1zTe9E/sCajZF1e
VZg4A+gSsIWS8g33cjgd0JwKH42JO4bugBpTU0ITZPgOXMFvvu3ElhhPFtV+1BhI
gLRKdAsFZxJH+rNXjyE5UmFTZtymDvvdRaXsC4KodcgkUT2yEbYhiULdRi5qmN5V
+AsoK6CL73PlrICJnvCOsRm7EOjh58YdSFb7xa6V8Sz/NZmPBEz+mTg3N85XnRXZ
LU5z2YS61bECygCd5lbGSB3Okna8IHiT39Aj5JQBEfYvAwbrqVdKkJQ0G2361466
O7dpBZCqnAPjnZGJGK2q0LjyBmgI7dlLlUKsCs3Ory786FuVtlgQDg69hl4oa5i1
CtD52Fucl/fPQqW/zFpUGJbKAVhNf7dQWf2lSBTOuKzMQ9SZdocIbayEf2PxET9D
L8KnEW9LgkG97wQk24jM1FbYIWpgBzgVclPEB8cKpXEktNeYWtIbPb1GI/DvmMw6
kfROhpid4gJbUMuAtpZC5TyjccenajUpjQi8E83Kyn3uQFD5qpgdV+XkUknsrHRG
H08Zms2fLLOR/UM86EvU0xJNgOuvGlW9jZavFgIxMM1k6IRniiDH9nznCefsWs9f
O1IqKEedr6py8D9y3N19k3jz/Fi4tCj7FLBwTHiaKL9XfNITp99MUPAR30oKV8Bn
LsON6JLrL/v/gI3KXj1TmPqp7QSnwbOG0F/uIXNz5AAwEyiEljzM9ablX45GV+ky
qXB00qyFwNye4teNhjGg2a/qHgrVJBov3BlEv9RX+jHqa6OEzvHp6FWaAUk0fyfI
2UoCg5LfNVhYTo4BgWINvSN3Mq0PRlvSw8jca4htZ+uXm7rMp5GMY8RMFJSME8ok
SuZHZ5DcCVi8tETY3IlC5jg1X0YsLMiqH3SdiNrHdJ34odop09GWPs1JY1lio1Rh
NVYOkhB5nyZGoM3hYAcUHjvbua/sJSgo47ABzgkQB0tIu2X1awmrjsHw7bVCw6cS
MC8surUyFr9BVMq4Gvc3PH3U5TGt/Yg3x0dnaZ9B+8tpKummCVw1vBJ9CJ4SrmBc
hEWWoibNEfuYwW/NjyVhmv8ccPHBcQyLoQX9mjsejMGtEGBzjebMFcJt8xk/QcSa
iede7GkM48eZD0vmZxo63eVzeKUvWBYP9e9MM4toQbgPVTv7aCVBCPdsisulB3hV
HzyQjgRxQCva01gsGUxg8cRFrunGetTXGD2UGto/2k96PQX9YC57Q2ioTYbRIwXQ
yPounE0Pl3KeuG6QNlEf+YOTrMZkbAcVfmMZGTsfGiSPKxtHA1lmDckJEyy/uOkZ
MVnowMJgKze+flMX+EjZMv6XeLKPM1AuYwSv1njxxCVdj7du9nfC58BvaIOy98ns
kpu1ForU5BLmnWeWH1eS8on2rpOM8IFhtkvrll9d6HUlrkB/R2rfoHKSWzfFHjxg
FcmGqrTG3ZY/G8277mlB03VJvAW+Lae3JqoPM37qpVrpsoiX4AGmrUWN0nYBWumd
HrH9M5/ZUoV2rv3pDkxHe7t7X5wCrrUfIB9wNmhf7mAhEHYCvi8vuPRZ/YuzD1bP
JTH/g7EmtDEREWSelb4Y8WmAb6oEVVk4wCHLjnOpl+bPprOwEbDEyOqO88Qlfv/E
wMoTRoRS3bqsHdCwID1zh16U7RqwpkZz2kUHbYzOszaAQTQTO2lI7bVydU8d+JDf
cTwNEe3hBp4uh9yLkPh95ZHLYLq4HaYs8zuRJ+tLjoPtq7kMsDu0NX1us99h/r4t
EQK8+90eT+tmJGg6TGsvXimFHyQXPj0AVvOhN6pLwtVmwsVE/fbRSoGEV5vHu2Te
yD3TgJPD4S/BR2Ags7xypx8b2AFcCxT+kTG6mIKXau7o+YQd8KtGxV4zQftDhAaj
/vDyxEIs/5jQop/qn4iBfPPqnlOos2fwi8pigaX8PGxH7DV0nvOlAqauu5VlVfFz
TBZ9rygq1wGY/bD/owbAggsLqp/QfsEQfJLCvzzyalisVIcDz0MMjDsvfoOsxOJW
swQy5aOsjU/hHMHfXTds16+xSLKQ4Z0PfFXK2zOinWZvPLSi30cVj0c4z1KBLrvC
6GYipF4Fjno4XofNNahTumNZoy/bT69hBh2vgnWCEaMtTQ7cfWZlAQ5i42StBfRv
k8bdMnhnmk2tpvXuHBUIoOUJBVM8Vw4LcFW8f8EVgblnTal5NfX4kyfn3HCpAiL4
RZbDcBFlLSeZAgqm6fQFUgm4s9iQBoZc3n5cqiQdKL8uHCYyBd/xnxbKb/Eo/WQP
A9It02Ky8BXP7BFxcONdPc6xTccBz2obsjkZ5NxlFr/719bzROagurvI7avUAnL9
LSlbDU9qixQHEuUEcITNS92v9FY5Y56HKWwwa7BBCSRRuU1AaJsDxlxQ5MDLhoZB
LWjz6tD67ME+OYK8h7DhJPC1H0Nz2NnWI/ouyFbLiSucfDA96f6UQCW7eKsGpUAw
yc3OaxSJOeP7VsO0uJ2y6zBgze7MxVTbSghHkUHUYuPJSR6CuPfk+zA/5voKxvFU
BqId2qJEb9o4/yQPcJhRIWL9Jtx23OclE3lPZkFbK1j5nRC0gc1CreePWJqf05j5
aASFOrE2oHYsQk464cnppMSG+823iY9f4JmNL2slTP1YP8M44Xf6makzfL8nV94i
W31Z01ch8S/fu6eL1JGv7Xqq/URD/N0QwMqcA5VAbsHruEjqGcOQ56p7a9psHe98
cuHwtlJ4UGMVyq8Gz/+BeQSBdPBw2um/KwNY/T2aPx3B42Ph+l1p7k/NtlSqkBnI
SQsEhMJltdl+UyJW6mU6RWGcNE3jRHmKXfEHMmIxXCD0J4vPyMbJomWmpYfqTv6E
JEAl3FHGQQwKUNse+ikKPv+BeFCiIYdxus2O5Fi6r/MuyRGx7FbWBkJpymhKBNaO
QaRMvXesTRNI+RVmqJHifDMibhghaDfRtuSzQl3RbDVTsWZKFYJED6r3YEEoJ+wf
K1HIj8IHboQl+b8xp3x1Q9IituI+saN8nA2T8WyqqmO1ocyNGteAg4n9rit6/1C8
njWwpbGqyJpPcljq4HL8YAPXouXaHso9NbhfPWHGcVbM172RVgg5ctEO3HEnODPv
QmRRpw0hP7PnMBdyQhLOvNAwgbxbC0+gzFju5oOHYYHG0dDkR6eBfbg7zGUabIl5
AZQcnFmwIhfhVAgZBRjOjPUZTAQVN4vOHmptJmusGrg8+/gpqoxQU4aQNoHSbc1c
RyjzGoDabYukpWrcd44UiO1FiQUEIR292RlREBCZrVHTeJiJSLOnACQ5nLcQCzwO
WUW7Voo7WgNGXNm0Q8DW5hFGEGxHyoyMa9kWNKCSMoiY3zqT7hiX/ht2EXI/j2kj
JGQYwweV106wPFcAemguSedEOchaHdeXiPbrXFQYKOIpHQJQ2CWCU6gEXmCq3d25
ivkhqc/uXjyVL8zrPvyXHbTjh3PDUug7tZK3QKVIfyFwUYEU/vgtbdu7w2Si/oYl
huanrDbeWs2i1pLlWqdC4KYfY8Q3f6LdbLJlGd9tZscjtOGV48JqGu6xx+cpzBHX
pGOFY1ZoOzbD0sDI4KALClhQj+BkbS36oIk9lTiFmD6bgymD08d3eR7JuI+wPqhW
YF6nD69qbAcOhtLlz1MlHZj4CE+c0wgBzTkQ/APxSFH1vx0o7HgYmvzwt3XtcxEw
1aVGA5Bm8Zb5byy9ntzTy+OFS+nKgzV0mpX5z32qZxNRFXIvZGY71Qlm0FC8/49K
cSKhOYfiKl8StnCLOyZZSrxsGQMHfpIQszguWHeBmKJss4lZSA55yLf6+6aX/4X7
471D0gmR/LYErPVQCGpRqCr8rae8yYn79Cd5EMcAEpqkfTExUCBVCIrViGg6U3X3
lfkA/BGr+IAQT++wcm1rwfxBNaPuCd6X35ehyeGbl3xrZImEFOQp7DwjAYuQVcJp
Z5Mo0VOgkPvb7IbzuebGcS1Ug6bPqN7LiW4bdRVKMRoX2Q5LUsIN0a5jR/Z7UDID
oH10VHkUNoN1rLpIOSUQSExTgQtF6Ggg4+exmVuqZ5heDk1HHhdbLOUm8XqCwLZt
Ktb21SAHRg27JJM+PU8CP05BVRo4125yeozYNXj7dOu+m8i4Hv+yHf2i9BQT+Lyw
RFMECiMKdCGsHog2bGmz4a6edkq5aDRCfYFsHYIjVAnohT6lwO7KqNOokWJKATU+
hh+c8bUryBB1/3YSoN9m2HXokEkwNPg5FY1ekINu07ciaUHZrFmWhBaSKnSI5ymO
SrAYRSnxr7SxoI7wQe5g4Ovts6qn0OcCJP3x6lKPBpNAQs5vdPi/Ek6HNzrkAkPZ
mNvV/Ycz6JLc89yix/635nNQYAn+P4arRaM+F98DZV635iQaNPjZI3ztoynvKRln
PvgJIxxSLPNfNhxUgya8VZZlobBvxS32QMr1r+OtvuS2TOQViy5HMVLcZVWoCJaS
hMBijxZC6ESO5Jv8tvroojdYFl+NHRMvPDKgD6kfby10yBc9jNUAfn9aWiSkGXHB
flCXuU8Zwu5Yyneq1goGjBK4kCKm9wujhGj9aDG8A0D4oBX4pqGxOnY2hpZe2vS7
6sWG2zB6M1yKW/rwAXoQTVuvzbNPqEMJ1bO3atXchiT9qhrgAwjs+Rt89LaUC4WF
+H8bNzMKLc79CVmGi0WeliYLWgEK3RAyoNA/q3yiiyMr+Ekx38/uVtJ+8H0KGVCv
QS1RK3Igr0THR3xbQfjl2S7ZzsXK2R5ifiUV38a+bELDfmDmIkkowhyjBDSWszMz
dMcDCmqHHsA59MDFNVnQ89X0eQT0SqM/FF23lOJtRg1CBTvTxvQ9UfFAlKigCpNW
AWFKuNLQkQ4ULPH2aFhilxF/v9jOtexyeRAWZsMAUc6w1OW5El7JLOgFewpiycJZ
HTlmIitJ+4Gno+Ij3f/JD24Lv5htwY2C1PNz7ZUx9cM49LetnC/e0/ifNlHRZJ0+
J7yGiKNInYzdP5//BjYC5MPKFLc5t7KiIbSiLh1t4zfTpSlOdm5VT4XpGMQqb80g
HM222N2AqQzK4qnzjTCir/MMG7lzfDZjPDg1X8dtCoL4ANOUqROxaXipBIqFQTHW
R8GydNYfBh0K0GizLzAyTY/3ADsHotbeac5Z0q4XkTw6toABNSSr4Yy1r5mDmtsj
i7R61vUd59QO9pHBIqtZTqfj9q9mJ9ZCPiOFjfp3A+9X4BL43iCq2ZkfZQem7YfJ
duJMBk+GN7kUzW28mf/NzFWdbSrfhxySSbVuYc2/Lt6rnPPaWdawzgXL9KgYRr7H
JNbzuDhnco8KjdKiCFbbI0/YQTxh2grdx3wVQaKuSr40iDwGJNJTgP61ABZa5Rpb
vR5e3hzxqFGulbmqmJemIw==
`protect END_PROTECTED
