`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JsNHUu1hUlh9MiKbSvl65N9JBEgmZyAmaQMybo/mVdyxOy1tFNeu0Grbk95ySfKG
wvtMSncaOpf6fNvQONk+T3d6JsloqMzFJypJhZtvwWldmMVW27dyR7eRceU7Rd+e
/cWHYD18NeftgV/HI29478bLInP+6FgDmah0ad6CXAiOn/Ot5UlSCjGHApth6EHH
vd1hKGcdycUk655y9Nftr9lbF6vAD8VqvcNDhSbnx892UsdgYx6ZfLAsBSOq/F+L
bxR5yUzm+BC9EVVebHaqvNNk2e/8GmlM8Kri45wlno3MFqOwSysmxJcy2mHVD49d
Nt43moZVHSSclXY/Hetx+SpoTfjmI2ke91PmaZjsV78m182iOz3HH0cXZ0fTLfZ/
e/KWUEZxrHUnIBVG416u7J2DynXEdn2F66wXbUfnVzXp7PSo3vOU9+3pMC7zofl1
pTk6l9CceH70/yMoLCZu8sX0SKdvu65NVu5l5YPeJY68wg8+fMPy4BCOGIpwfLbL
4yN+uGyn8lroX5AEP65WlpZMqM4tk1X2ehOIYEM8u8jq+MrEvSsXdqQUYScbXYI4
wkizk/6TTP9TANVcAxyhVrXk5dQIl6zcfOCECevHooSQMn/DunhbbGdWNEQaM7kn
Ra/MNUg4L8/GiqHJOvrN6h5TfEEMMQ55fmmwPCArSTtntUCtAEuc2q/gydjV8pQ0
75Acl+fp7D2EEfVQcg3zY+uqLVUb/VhDx1fXLmVVlMQeHYEaOPGdmC9YsoPPdMEn
jqjPAB60l3BhndJgclXMiCIhA3livPGRqzp8PhdhD+6oGCPPLrDnzIvuUKQ4Jk55
XO+oFr8/VOg/ay6W/RhyYs2GbQaTY7xlrAh7EG/5QGuNoncO+RsaNx2PXg/K+RZP
6eaZnjiARg0pwdrCzBxe5IPGd8u8siJAso5f4fT0TGM=
`protect END_PROTECTED
