`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hGMr8J+AQIyVlTIwhDzR0Gicr7iY4sJHAoF628hPA/RYaWx8X8QgR5AyG7r+MzSs
fLrqKdfYetRZuqm7YsmeDXwyhKFi/VVNrL4UOXvGxhxDOe93EoHYwLUdiSv1MNY8
b09oVMSZB78ByThIT95c2VeAyYbuNykNpCbGmQ0gO8B/Uj6sPl0QV+5KLh1bJtkI
lenOKrJICzr+0YqSdaxWrSzPj2M/aERPic+gr9kuSxfR8dxGj4oaAwaR3y0hrIgY
JlWqrgPM0JPG306VkNMJvyQTy3VPpKn7iZA1amE9A2I7SDyVtjpbLz4Vk19DKg3C
R5EggreNG1WpFuK9pLP8dme/1hcz5t4nNpWQS6n+CrU0Q35zskf3zpnE5Gl7MdkE
iXAEJHu98Uj7+PK/kEb9lDhWwjApFCMF6tFOwhiKvCI58On2HFiUQzCRIbc0UqJ9
8JNNHxbSqaNJgtiEnbpGfr4aiE7kP1PSvzxsXJlJAcZ4kGAUV3jn4etR2Oeqk5Fm
s5WMmlJsl1TH25KlKeFGigvcREAnpCtB+62fnYxhbjJ+2yhX12hgQwKDNAXkg4gV
hZNCVz32C/QnoobxZ0bzEXy2zaL4lAzau7KXXHmgSMzLBuAR/g7TwCwpHGXu0Mub
OsiIgg9lUtHs2QvQuj01G2brop9CM8S2g21emaecM5qjjK1HsMWrex/gyQq8l70X
BGkebobfDIPUE1X6F/ikVJWCbwQNc+8qhvGzVVsJ5cpYWqr00C6R/ULFSj38GMp+
qVQXEAMPeOrHY8jN4WepvzxcbA+jmaGe3lF69owkwuqT7tGXxbkE/LDUwRJjcwSS
/iXRvoXY7dwQdAgmy4AHw2AOsxrbc0L63SQ8IZGxhNN6+YdqxzTja8zLO8aNUipN
y3ujfJCk2DdHFGiOZr5hKPaqVtzUJYfaf/zJ5nKEVrs=
`protect END_PROTECTED
