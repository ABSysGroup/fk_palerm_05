`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/hFqAjqhpixrLW3XEdUmY/nacEXTZIOaKAn9ly0WtOQ7NChvTodpauwUCl8osOCA
2vXUgxmGx/9nZ89L7mh7xX9SUkv/c7YTNC2zj/c1WjmzfS8SL29eLkbSSFFu9y1k
8OtGH596OVEnfAWmt5oPD0+klzgKX+7uQRCVcTPDv4ssSeJEcyUOsaSsyjDKiDPU
pZZfhyl2pF/cdoq3+PONYlkgUvmO6n8YW/hbmLNHcz17OydQBZcAxu0q0Y30XyPM
C6nrjnJQz6+RUVM5WlmRuU20IDebKuD1wiDehHSwE7WNeXUSLlFcLEAHM6KgLqOw
U3YmwmGMUKbFDmeIUDcjkbRyTf47TMPm0uXINpaxbnPMJox1kMrzz2nH/V7hgWhX
+6V5M63WeiHmML7FQV5sjEoA9fnyzFedSrvTLjuQ7wDyJ5q9Ytv7TLYHHJL0ZDAd
pDJZtMq46wJFMZGl1M/HFPV3Hg4dKX9o/zBq25MlI/DfU35aCeqQxfTpOqk1ZSfD
cGFGkx2p4VZ56j4qhrsk7g3jtkKciMmUJ9rsgAP2e/drq4YVMjnMAnodZiCo9qPs
9K7X0TU9xHsVqxlfAUApAIL4yqNjHGPPgx5+Xl+lgoS3RW/Zk74Kt1izC8vjmd4Y
kvR89HqvrC9bW8lB84XYioija/8CEh2jXepBpj5JvA10QQM6HGS8YBmSE1vi3on1
4Ym4GHmRfrAJMtctGb7ddeuXANmQFAft5tR+s+BFvnhmQigBmi+dOq3lSjXk3exF
Mj8kPIV0uU1DjN7hhWAwDqcLdVGI0yWKBSIRek8XX0JutcTn+f1WopApYjX1iKJ5
Le8qKdSIcbTGLQY9jfoKJrW/igIUPc06QkZsWKGTPrVerC0PVI1SA8mxkJvS9nAf
mplKb4RPzTLwy87VO4fzVoNo+GH+EHRCdKrH9ebqgo012+HV+bhv93/Ul8jzbwX8
FMB/SK09GOD0GkBw+CFjRHuiLYWDsTBZDWN7z52XKL7tqw10FOed0iYOaPDagdtV
7tCPXEGVmOcPI23MW2rIczLzlLOENTKZd1OgqGxvgb7j95bW+8OCwlQuFBgkPdLf
12zMdWs3fljwTpvr6Gi5ErzAV6BILjxj8bZ7Mm0hzGN/nLxlAjJv5luMbWWzp1c2
r7zKKmUhuHNdHxoZ6nPaxEfuc9R/MGcSKt1A7f7XgfA+ISdxqZN6ktut9k7bYRNL
xZxvegNLbwIwb4ZWJ+20LpzYU8bihBWdufgpOgGS3b9u7numocApMIT+xXmG7Erm
6j9ZyucZdgjhLKtFHl+G1DRi9TuGN3XMvb7DnI+xL++l+2yS/MFFsdjaeqOR4+nh
U4hH+aBqj2SG8Jx/JGz0pQzbnDZ0nkxkk+iVROtxw+vza7Pa+6C1KAIEbRr4SxWz
EdG4rP/GgJYQ7g/k4Ylw9Djs29uXZZ2n3iRQf+UaMedlx6qfj2S5SLrvAZhDVGPz
+n0dIhqYM5lPqjo6ZAA/PyuW9R5UYgPpgwoO8dQs3z8ZkKpHAlGoderFj32pCK8X
8yagSHa+AXoeiWBT2kI7YwnZLyjck0Le6UAW3ij7PO/WegzHAhe16WcDnvPuH/aS
gFoO69g/4r5No/aIAk1aL4ekK1PqMTBZ8rTPcsLiWSE3VQiooGKLPVqF7/1JLyMl
q2KjpFVpXh13xeIQEZj8IsUl1fWl2DPlPyxgGI2kgpI1jZ4LZFh1isH8gm+hZC5f
1NOkBdzGEKxOkIHvv/bjQcYJAnyeQTgGWpo3wNFjVZv//R2JUPCPzjGDbMxN2zVT
UEg0xMfCKdpqgtUrugJu4MSCVTHbhAXBf+d9v3k9CmTaGPrw4v5D51hiYolXSkae
YCf95/iTq6G/DiUjtYVRxEP1PKdFDGpNQHLZQ+93IJgtaYp4PyggK0QVZ9zgaKk2
G8ydsVWMkDn8/0Oz8SQvqzUP3aG/9xVfYvwlCH5OFOhbrzzoGPTma5ofD7UbtSR4
8N5IhR7bkDYmkLU4yyayZUGFf0djzAtmi3h76YEaunTeVojXXMNSUT9/DIWGehWH
OAZ+IGNGky+x4MFA8Zzu/3xs6/y6Tcbh3lnZI7KXX8ROTS7mQnC2040kG2qCxqSx
nX/0P4Rm7xOJpyvKJVPB7zDieqHGerfIXbOA+gCcJJ59hDTIr9xDVP0R2mgNup0L
C1D1IReEH5Y4GjAZxqYrLe+ThLxGmc8td6OKxo2ltTYeXymv30bTeR9q/wYT0Agr
9UrYG/AyAglFOI4bXacK7jAnnGoAYAX8HfCxuwp7MJSckuPaIb8YfHiPglbLnUSl
JpVAUu/9N4QXdtGi7FnYPkaTVCTsfERJrTBjDK/3dXf5HBKDj4wI3wTPdIba2WDu
gEPhdBCDzksgAqFhbY8r4I0okBkEgftiCkM4vHgiptDYDzS0wdN2MZroEgfpB4yw
Jd2TP9Mf3rWnFKdpNA4YpxQS6HditM1MWtBlTfyRrH16NfeTa05BaGj05a0/Ui3p
RCo+9m959P4bRuI1/hpplvuaHVXQZs0253yfzZGIgUuOI0vAxXQdt9pbL/XQsl3F
bAMHzHpIIiivl9nSKppRVDG5Lw48ILhi5vrmHlmsITRdW4MZ2UHsPbSTvIGm31kq
Zivgou4BhHWwH/Xdt8kfw+PwtcsAtBZoMlLonpnIs75axxDwtFkGMR6sxzlWenkp
4rabbceyHseK/9LO4mE0ArUO1aYdZANKDeQ7WH+yiqtHF1vfTZOJ2gJ8pRRtqG0Q
Mq2aM/BIRrfblQ44UvqSl+mdzYGHy5ysgem7LCTAHNtk+cqj7uXhqsOa4UpaSATe
DVncd+zi8Ay+x1bt6klVjCqbUtF7x1h93/2VLX/s4ObPYrRZEdZRdT/CtkMph07S
xWG9E9hY3Ivu+IXckg3z/pNkAtgttIZD613wNwz0xNJKgA+bP7c28DG4zewnDJNS
gn+x6RRYq569OZ0A4PZ0xtexu2iojqexsxMnkmNSDb7+GvDzxkCPHb9eUPhrULOf
eUNRtOK4S/EXbChGN55lXtpniYCX6xpXHNIE/xer7uKab2K4ax8hzFIHihL4bgYH
cHaGBahOA4MiEz1VYgz15ohzDhv6eBQYiLB1SqeyW2kBv2MkFj1DPHBC+HMFYdSE
NkjU4xF5eYmuUx0kfW4PfYcuR0H+o6kZPGkK5CWJYsDd8luyLHA2wU0vAdPFK86n
seN3u+hQ03cnByd0AKvXifE6cqd/EaKNGMvCwRWxH4zqj4H9djQWpHirk7XJDL13
ynreYTuwjJUap99Q0YLx+w==
`protect END_PROTECTED
