`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wbzVyrIjO4jsYo+liYrB5ku5zUeAPvbN6UHjjoSJ5X0hiT+jiIXCb1M+uc089/QE
X4v7oYhIwwVMvjDMmjRZCDemaDXALUhbtNzX0ZECZJ0WmNl6f97bOJqYRXICJae4
pygRpi3J9l7i2+yetmeALJ+jH66VQmyh5bOkABYTkgCPgbGUtQ45JPTayHZGNTfW
qkTw/RC/fccuTZUT5az7GZ+X4oRzCrqFgMj3b/u9kRbQ15ss8mdQB5Vasn73NfWY
V/88zb8Mvc8VYBlvkcfRcEpUbtQmAkOmhff/bTEX8vDbMaknidoyMNebNn4tAghx
TD93A502gqdCvN1tU4WxZQ==
`protect END_PROTECTED
