`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6vpcd8bcueRSmQJh4kyiUKbkjPy8/jAk4aF/jTg11H1n8lfV9YECSvn7RpHt+t8j
iA2d8RajvxILCLRh8MOQU9GEN4XwMel0UhZrwAJ53J/G0mPsWF/3eQ8bpe6O0JeW
EzQT3IymL61G3+qNSbBj7TOQucbaheUyuMxDLZtz4Q/svXmo6blxsWjoMKNlNFV9
eKPXAljHG00DpKxCOFzwYcS2quzIA0gTAR5C9LR3CIhVswVjvOj+Mjwa+ZI/P2lB
daZt7Ay0ONMBKp8VlAS0AYU/o6E5hU9/t2gZGjKxWx8nuksn1RINeFhoup1wtPhb
PK+jutA7DXPRhLBkgkuhZ7I+Vbkr6cIUdCjK1sUwHrOWfHMb2dADgi5veQMlPKdx
1VWC71GUeXhVaWhlNEqFhGeUmIznsUTKiZoufXTv+PFXX3Hq4/MbGqgfHvxuNbNM
zVloIg6iK6T+yq6pOIl+2F1KwAekFkqZC8bGgRl+KD+RwtUh4Sixvku7xkMWH6em
maGsavmUNZfQ5PdDhqME68SQP/lhSxyTTc8c/IV7Y+3AxxuNgYdM+ZN1Ze0vTj9I
JWxWLAVSuMbooEV+eMacC9UNyVyNMLMbjTxpyowI7IS/PLiGXlrlcYdOy8jgW5jL
`protect END_PROTECTED
