`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xsQeEL4MK2Ho6MM2Jy0U9tW7cKGVHQ7Zv+r9mnc5xaqtuxaXrBA8sKyyOoiU3am9
fnTVi5CSCBeIjetdm7nuw9TiaYGgRHdc9lMizedrrpOdn/3V0D22AM8Vpyi3bY57
HA056ENIaPrdHmbU/98ny+XMN75ntiIiRcpAUBHKdCQDNnPgXlFgbv/xFqD9IDb1
Az3TYuXlFzF5S3gkcrflXJjUdQtF8o7bAislxL+iQ7vP9FQupT/+p9EAeZEDcu5W
IfDFlIpg+uVqGYHUrcOxhZlaXYsOuH9E0qea7TG0MAlBG1Dy8BxweDmlrUOFIC4t
KWb2Y76jLDye6Xlfp4oYgWkLkPQ/+7fb34NnlventDeqdrgVCjeRJf5AuxeIa4KB
ihevGQauh+HF97fqmHMDIq7Xr54uGr+gT+Fy9DWO5DkvPPSx5NT3Gyk7GfSCm6bi
AB5ZS4pNtT17J+7/aoWzQQOBrq+6WvSldraqrDCj5M27gPBEV8GMgk0AFMeIbYCX
b1HotyhslHxkEA/UQUoUzdKG2amd1SRsgpSkdFlvVpJRFmYPRIQfvmVebCim+3Mo
X+3XVKI4YBXD2GyDIMzMB7T3Mr/Qzzv4FcS/fT5ihp9HwAthVTLQzsBekB+FVKq8
wqmJwW2FW1IncikbnPSM7+PfmBSCf0eUgy/jlgCTFLzKPGw0hJksdZKZBO60NSVL
gYMy8XTANRundyGmHWbm8yFP1cQ0/sQo8h/8Jo4WSNgOPhaAc9ckaKsiyxK2tJ70
tQD9SdVEsYcDqIRbnT8YGhLKIebOydrWbsJNvzl/6oIxB8xd62VKYnoTlzUju0NL
Ck+cCf+7HQo/DJ/IPXeO1W5W/eTJLZfFpe7Ibwt3teUhahm9mDF4xyeVrdAlUMs7
cFqpp4NQFzrgclhj8tugV7uHqOcKOyICoH/Fk/OQO3R0qVrpc2S9Ju/VvpGRONFS
a36Iju1XO/vc/ulQoAPIIhBrC7/jNAb8FbaRRaYYC5KO8R5pE85hxZR5FcommVBH
IXreYXjBXQd0paKuIpzLsz6r+HtLw8xmeFdkJCMxCbQSS9eC4TXXQRiOR+dhZAwJ
0pWP1vplGqbaRBZCaZ8pXO/cEiwriQFMBCl2wwaRCtVSFlXBYcS8z2qLwbwOJ7WG
h2yo+oSJr2muUpd0D131/TfE5SDTrpOuH9A9ZtEcHZiiWuLnDwXXm1OItMT01Fr6
ra+TWAxdZr93mGsqnqFPtFi3zTTuR47Cy6mtMog4KIemN4hSKIWpwyVpBDbYVhXh
Mvpk1tH9p48CovaMNi3Ci2b+tM/Yu76G4z4lk+9rGIxXmoohYIQbyLHrlXfaRdTY
vem66Goyo6bk9uAAUvfB4n0AdP39oqqMUMzvlCT9hjvWFtShQqYj17qtLgiGNhnT
/ROGaNLV5ba+pTrEPhA3UchCsS8UUEIpD+38SKKA2EsMwyLBIwLzuFAzbgj+8QP/
tAlkMFxhIID57dyebAP86FwVd1cLZFX8JuHPqONwSJddb6V5bfyR16VkEHe5YYGn
e0AjG67jI/hw/1FB2oQGTGT0H6tkSWF7QTdWF70X/+mDM8IHaESYaBlDt98tGGu8
mrYe3EJQOCtrHjZ5fsY5cEqwA4bvLofBwxYf2vepOAS+MaTsfKlILm5+yUhIe15f
PIoxg0yTHwtWaxSdcDvrM8eq1ulaaEL0MCAw6aI/5ZkyANfCYoD2emk23oQLg7yt
fahPnLN2CtPCY3elKvTy6LoC4lrAgf3JFrdURnpxx6QRuCO1dFYbaWiFCZAhy58I
vAcKbqgmKg2R/JMpVxHTgCoDnq4ynWf8zggd6XVfNhmeKT8vjgUg4excpx/+8sx3
aDJJA8qXgqKw0qJi/A0fhFfIrzAusjP1bVxdujUUwUobk3sUav6+7GguskbC6Yhc
xUmnWucaAf7O4X/z+765RbaWyIaS10H5pZcsX5iOu7NwVzeCP7njsd1GDpwWH+KG
t9HcS4+HYj5uova40S33L7MJyYFYVnZO0ep27OHmVtUZ5KtD7cuTYcYAhf1HqLtM
LchBRdmppWlkKSG9UWqOMPYggM/C0LS31qdSLuWCNpgBA/u0x0r/V9d2SgW9d6wA
/1ppYt6sxkVv01W07kK+IqVps2xQO9ux/P6zjqELdQUoX3Yz8n3VCYRXiw6aEVws
Z1wvRKn/4sdhdJJStCTe8Z3i/7MUEUCnH6GKzsES8seLTS0S5vU5GGHDzgBBt9vd
H//laPk6V/SUuD1SUr3UrcMA0eEskfk3+eooIunVyvRcZAe1xVBddp9qEbEgQQvO
ukK0jH/w+NW7kENNSqa0V/mQHYISFmXESAe5QjqYqofIuO1shSfRHzUuGppkOQl3
p7ub4ifoQ7NzwSg0H27d+JC0sK0slok6yg23GX04U2hSpgokPMAXYJG9eQD2rTOj
45xX2ZRQ/IAVpuT3oLvsDkGT6tOsCyRqDJZQxrSX2JVKTAZqLD+2wE/9XOw+7jBO
7EtqCsaR+Sew60Am6hcLHymaTZKb+ZETtO96j/58x1F5DEhwSp6ANgberdO5EpxH
`protect END_PROTECTED
