`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lbVZ0GAmY2kMHEcQbJyW7YblaoTSNXH0T3LPPfKdxk3Fg5Q8EKAUlXmaP9bvWhDK
wl35u6MJYMQ5KJN0F7Vlvw+Yvsxb2wH7r64TAdcv+CUeAxV5PP2kp835tP+pbCuB
nByZEQFyZCQvfyq6Qt/naqeLmA57ljhA1LXqeX2GFfHBO9BsTp2pi+PFZiikReT3
J9bcFhgfEibwKNJ9NrYcryVX4qTIFuJrLeRwbvLB7mDVpadEQ0EcrJzK3USepwDZ
Xlu9lRf6h+M4h5BlIVH9REt3OXkX3DeTGygujGIuuL6jn8lKURDtPx+QO1z8XGmu
Ub0p0PwYigLJ3DrX9E/ffXdvRWLcRzi8ZvetTEIL16aKBZuFlFB2XIc6Np2qtyEX
XR3HEQo0dl5yJ8W6cMEH8s3gcQx7m9jEMO9WHHwtVVJlXNFrfidbb70YThbleSig
cvwwogv8BDIlwzb5YvLN08bFaI+I26DMgKjlajEn42TAGMcFw8fgcY1xBQCjOcKA
Slf8oYbPSkjaupfDw1kWfA/L11XKL9NGqZn27Wtz4i77banfQjT76Q4aoH3UN0nC
JL6tFxoqPrnU0xhNhEB8FDLIEVjiRDWxr8cQAaT6YoIqNknUR3y1UHcuLc+oTjzx
O3J0wGQA4UeFaag1VtPudgTm5CGtyUWJQEjPpq5imdMA5YhSESeyErf7jwJ9I+cn
Ky4UhkFHdDwxV6LJ75eTL1v95B1KLifvYsULPUAciN2D1akhXcfu8ElY6Dxcj6Ya
Lk4ImA5qE4ENiXpeN64CS3C/eykXMn1Kc6Orlh3Ka9kaGSzXY6GTJm4acKtsOPdw
RPzYkjGjQuJRsxO9Wb9Ox6RJ8b3pA32evNYS/Bp4cazm/V8aTCfUShLHB1++DiYW
qCCb3nFK7uuwhROvRpLCnhSvisrt/LypDFk0x7fhZoAqBjPZx+nXjxDJKTiChJ8V
PVvKIK12zNet5OBhbW75gBus2KZBlL+6LvM92Cg+sMsUDVfkSQ9CZ04xgweShvJY
7pAMSNy5zR+vuAvFkUu/F+le6E3zNupHLvDOOK9Fop/d8fhm1zDt+YVEZNT4gRC0
Q0inXaBg9pRX8CkuiOv6KylHADlvn6BvdhoTnTYbtYSvosChNOCBN+FjfgGZdIuN
3E0RRdX+JZkgjIclZWMJ02zi3bFeYP+9ibcKeqCwKM4=
`protect END_PROTECTED
