`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
37nV2RMRbxP0XMoqxNX3EIqMHGGcKdF+xPdk3AOM6ZgWwRCERkwo3Ks+bXcJ3xr0
QeSwSMZlGiYAl78FisH0fr/wN4oGA4HFxSdUWHxW2Ss0qXJymKkRFXKtODVJ9vv5
eH8/V2sFRvA3HFZP7MPPn56rz1dYNF4gfBm/Ag6lC7QiDYTo3CRVuAhzDvkZK6Xq
xILJON5bvpI/rTkw1gSKwIQSX+wvQi2FZ0ztpOnYyiLDsPr88kMD9eA2t+j3FVw5
hgracwFsyzZGHB7iG90OlQNC36FpcS6eFxynnncaunqwJEsQI4dfIvdbO91Km2Ih
gl25pLFceF4hpp8vEo7w6xKZMyFhlRU+mgTgS9gewdcIAm8hM+F68J2fAc6trTMo
/uqA09VZI7aprNJUFeH/5omLZF4aGomfadHhgLROGYJ6w1umj8AXmmbo80w8pwJe
C1adJHfyN/byF3RJ0o5slQQg7noLfyCI8MkZ1uMsX9UZ5P0Br9sdtDY8V1tyU9Km
CRHDy6WlX3UE0pizfIb9FgTtvR9bZJP8lc3hnRn7vQnJyqIVCFXEwjsuQnmY2ar3
OLXfY9O0bacLvaQ9ymkO0hFtSE8svakrMprU2iL84C/6KcHHIEOgjEtyZMpvsxm5
/VzZN+sPDAqt1C2NiRgFZ71y5wet7chzr3PYncYfPNK7qxJDZ48EgV5visfeKzq4
c5A2DdVooY7N625Aja34ZaKkaK3GpVGY3adliQxhwO1oNf82hxZ5NRsmPYO2ZTXh
OVMkx1L2lI+ThlFq2vZpbLJwUKM+4vLGr5dWmwHijKJAq8fjBIDb9SMllceumfZz
ZhaU3AkE/4bKaM6wCkZIR0igY7u1HxemHqu9kghKg/f0JeA5mEAb6TOFepVGu3B8
JiieeiTupsoWm4JBxfIVbXwmznyF5kVXtQc8DXhKfmTAeSQL2zh3xoQPdNuwq+/Y
yrVha/+CjK8wEZjXLnuRzuq50aPso9Q+GCmIaNW+NGLS8AcuD9pc/GrZPMYod+3U
4D3NZ9QtKFgurdIRqq5dpfg5O1KGgXjgqCJ/J8pVlrwzYy3KNJTqK4OVMOkGdFjG
ouyG0wC//fZR1m74RowhSK4qfY/PgTvUpCW0NOY8iKsxYFaOrFDSIQCOVQjBtjVK
ozvb0KbMnM/twcjYnm313wtHjDJH4Y9NnyUzdTp5KWNFPRRt+TNwOvuqiwn4/VPW
eq4QSIRMHtvssd55VUeEeE3+g652omTh7KvkzBdqjjpZZRDQ8ZXwp9fyXqPNJwd3
Pts6WRlWaQDit6Va+Z0RQRX0xR2JpI/GUDcaT8CIXGo3swrQRF3Q3nn7fFwNm2X6
SPJ0yAF8DqPHdmSfjwFUHx+pw0YeqDSIhofy2YaqyfoIvLWQ0yuqXm4VdMxQ//b1
epMUhVhZReC2b0PnuDKlkrtlIJ5jn4M+7+qIqPtBXIU=
`protect END_PROTECTED
