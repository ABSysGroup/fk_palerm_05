`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5WtXrXdKr24aw3Cm3VGOOyOF0M9qcSljpLZ9ZcvcMZrh7zhHUYi5nC+PvEpqBema
PbmzybB9C6jN8+orJc9cLJuBmU6sYJTdXHx9XoUjepuQ2F3L4ZS20/JRoKDtQi0U
TXYIK12HS611eond8QwZlcD4byrtDq8N8U7c/h592dsWWXm+zisEzR6EOp34jz9N
KdFc/u8yHJ5SQjbq1yJh9jVKcDmnr7oP7iRWi/8Z08L82+XOSm8o6j0lt1TySDkP
OnGT2FxAo0RZEghh/u+g1EB88VmqD6oa2gpj4NcvWzoqroKGNcSDqtexxxQA4Qwy
GNSXw7umLr8O01HWK8YsqsyLscMRiszod4KqBDzeK++uVJJ1drNm9O1E77QjrET3
vunp9OF/7an4HV1HVlVUsqDOXgmMioVOkiy5ikPpPIbJf9tzweqq8+lqMBDCzujR
Sppyc+EUE7h3wx32u5KxDwgMcDsS1/NBQYzOgLnhg1oL7nJ6ksyN5nU4YIQFVRae
8P646sACoQXm/Ba3zCNfMbeUZEXs218ZIfy54K3xSe9bG+w0ehgWbSi5qujV6pZK
DcspFbkAYNIy+yJti7wpfXN6QZYISIISsCJT3/uNU8TlofC+yzx6vNhcfqZXhYwk
ZeBh0Zmb2aFp4j4mKHKV1kH7boO2VAJLGzetNyLgKQOcNGnYyJuaed/DcjPVVT+P
yedQGiv6ITzTAt7v6O0FrR+khkm3K8D6X7jPIIHOSk+EACFJq4CbmuKh3ALrznnT
m9RMAMPjw1oi5Wr8hyJhofJvpLTrKvyDi8T+oFFGDRsSGK6Z/f+toj0L17X/aGPN
sAr2s5zqWotEA3b/I9FdT0qSyn8TnCLuxUdmqrCMX/wQxVAbYXxWWnZ0MtI6Ukm2
8Uzb3/uaA1Fb1dqvT9dJVxZqx746+1LylFrYXJvrB/8+H0th7oXPDxzvyUKZAven
Xk90ddAIkHccBTbvlMCZ/o4W5FqkDaOHZR0NTrY+Ze/tvGn8AUr0SkVyvSQDZfnC
lSIJNEXdzePP7ppefwnPCU6ZVl8U4joAvHR4wENLVK2KtEBewflUGpnx7udmdSCg
eP8HNTnpfkrL2p+cOQqoACoMAlWJFMgQQW0Xd+nE6z1y+BJ9gfxc8o3baHaRS4nz
Sv/VPYN/MJbVCd9aNVD43DLzGHht22c7L52xTyNQYxyRNqDGvc0+gbCK2SIrPJQk
f6LHRoEzRERsLpIljz3iFf+K4kkkcOI0FJCWHECs43w1MRpCSnbQfnUED/lDB4oJ
PEKjvGEPCJ2BbZuQms48iCG4pxZ/g0yjPEFBJsFvsjvocHwCJm4XCxIdTj2S4vlv
w188obmLVkFnpZxQksTCeaTbOrLJMsA4Hg6bP5+osh07+wrrGG71N6yBeC1o0p5x
djRC0rGzP/jdZBI7DNhEc4ZS5dCqbbjkkmRKDlSpLttnjDt5jCMAKuLQt2AzL9pI
Z5RjTqdHGuISQVVsp/mZu8QpIbFRhIxwPc2di5asblDE2jwCcKBiklEOaaMhUTDs
1tPNJ1xQySraBRjsB8DYh0t2xzbq67tqzopsxs0pBO5MTAWGgGn046A4vpFxqCHl
2ZacbVhVnSLe3XKUkVVS56SH5bpKKe3aJna6y1024zILluN3MDuBpj+ZY4tXwnLq
tdEk7JaJ86Fubr7FmI3RgoQcvGk+co2lwhS4r8PZyKjftqQXSbAOQeGkDsqNCqjy
Ptf6UdIlfkbMUJGoW5m0gj4Yq5Zbvgz74yV8XpDFS+wB0o8hgb5G1yI7BxCg7EMk
FIUw+THkiJOsIFH21Jc56tGIgQ8F2mKg8/G7jRJz9k3mFAN3s/9fWjZVELFUQHmo
vCgN08RbqOAU+0bLe2cQVEF0eGVEDPCt7taRXCz8+fkh1/IRKSsA7LNaM0edvKU2
g0cdaVcVsLzg+aAmiTS/SmeMrWWRC6B6ERR4Z4No1gF+8SDnc41JpT6BHtDKm4I7
pUyXIpuO0SbryDuiB/z9X+I0bXIouyA0pE14QQsXqswdV7jjAK0M8AjEf/VA9EyS
FlEjXgOd41Btiv8Hwx33qf8ji7FR6t2DlfJUnTxKO7Ry2LIGvYCM+sg7dyq80v89
CnhjczlrG4nKluSf0Att7ltJ14G82dGaWqHSrElxyBNo1BMZcSZZ7cWb9FQpC++z
Ntu0prh4fcCvfvZeuv6MwroKwB3NDi80L63N8yfkUmsHrUgon3B8S1V1xj4gbh3h
71EBA715QIa02vGrWXAWi2OoUNT8u+n0q0wE+B7KYt8POhpSDtqy4MOYFTrsi3Mj
8EjbzoSJ84ltzGOh5PHmZ2IrbniWl1CrLLjZwNg3t7fnTWsc9xxxE/AUfQUYC0uu
yFife2sRFbm5ERHszYHd3gZAyI9Ebb5rn8MetzkBFRvpTTPN7kwwqjbGHuIQy6yf
TLpEFXL056ur4/o9kpmzHzgoo/lTVan2Ksao83R1/QLOfrc1mvIryFT5gLZkzA8B
9K68wawv95PjiSLbGSAQQoP/81Te/yK4gCW/SwQDu2EjUGb089xpLvizb2AY7Jif
BHW/sRIGApWMwlRPV9gF9M6l1BT9kgEFNB2ZVTFXz9KHQEAeGnO5gJNZez49r41y
6Euw3eJVE0nj0tET2FmAWmlkjueO1g6vqzMHhv04Ot5Y9i1fIJD1jDjqyFzDxf6P
dodkL3jqyhjwiL31pInhlaxEDoAVOIxH9lHUg6828bMDbIMIttyoBzDwG0XfI2kD
Q4yi/Sd/7+Nv635mkBruEsL54xvaqsidfY0PGYoPtwcqtvOaBeh9YGNBU8NbC3BR
8UP28QNMqUMFDk5UwlC1rx74Ud5QhBbYzHczxggJXcoKezKhowv9/+DB3vEg/pEo
/My3tPWWLrlNrq2F7VJdolpxwpk2URniYeFGwafLoVITYl2UtCIbkXIcf/LkWA1z
bUsiF032XNv448b3dA808j77fU+WwCx9zH1hRkB+wTJA9z+KceYm4cEPJ8WoCw5W
9vQjemqz8d+62xymOvHzyr1LgQBaRZuSLjOIzzwOyWQKJuk0+Rprie71oL6ymo+O
36yJBws6bHbro/Ry1FhqgEn4M81r+HicSQv25fBcHGQWJvpMScppeN+SRapr9hJb
ewcnT1kDHBnBsRN4qhPqMhaidHYy/F1OMwrnRvyZXnd2PgylPWsmoT6bMrBnccDw
svMbNw0qZibHF7IVBWxQuZiQuqo+qdVVqaiFhNo0+ynBjFvZlsWr58Fh2atnDnlj
Q9t7J5WQrBs2lFcxBtkqrhEJMMwa4THdkqEL5Nj891gG7+eAjVJmmzno04fLdOk3
nwScSxwHcH+r+zdPjkYrkO3I2i9aaGlhc7xru1TF8dP0nEmyGnepCTZiNZ/MzptY
ff45QcIecW1PK/PQCbYduqifDJnenmja7RMZnFZJR5z34mm4ySz+dOYaE2AO0ODC
xkxbCUFDvOJ5/YK7r4ZWzajS/ixKoiINidkPBJbUS/jpwz6UdMmnvtLLPN8TbfC6
YWyDKwO6k4Uf7SKWDgEaEEiHR//FJhfUrqV3Dkv3Aj0qVHGN2MZdAJwJyYIUPScQ
bSfNPqwO4UghIqrKT55viFg6hrhz0qNTI8PKPdTWL5u/+hivoxLm/lg16jYRMOkT
fdujAPWmDjDC1QN2sZHN95v1PD4nui2p+aX60GBPmcRS3KhmcIZr4NUrJ4IcybKZ
XIMOmZBurvTmpn1tofobD9EhDnP3lc/5RfOIvSN3EXl8I7p+OOgxSvc3J1DT92q9
SzG5ic9TK/RaeXHSmj2OunA+LunTfBXsCzM8u/bCVawCmvRAs2TWM5QrApshQqcu
GnhXHyG1WBUuRr4AN1HH+fkbKl8/25vdIQbvwz/Kw0hAuMD5H/a2PTH3Nd24tTBa
ythfGSNVQuNrVkmG77V5tSB+H8c8gpDjuEZvzLx2sno65r5UGym4h6ZPCbYNsdpp
8DsNtTEEugdb2j2+Ntpnq6AW3HzDbCIIjeepREvLbijiD6ZLGfXQeTst7LEslBZF
gJvuoMJTD9ccLOd/+hQovwQjQ2fECqjzMFwe96HHveBMZdQHhgI3eX5KtwWES6pe
ktf60T2W/v28CyWxQdazwa9cqnHvNjL5E9II2ymxNCiVFeG1KecDjtX2RL5eBn/i
Dfl4OP9uVXn+XnKpWPpLtA48KgN1y7KLTXs8WuUh7ahRdYAykhf7heQDbblgLVfy
9vR4paqYx8zTzV+7IRV9Y0CTnhDbPckSyTtsJxJ5mFeFRN0AznD3X/XgL3B4KBOS
1W4dBrVWN7fLZuQGZ5XQVZWwVLHuLOmhPxzEQ4MX9jShHPtG/KkOBTHqGxxJNvLz
clW4MR4EX7sNXEww6kXsb8Z8oIhpM7UNVrcFxjC93k3Sei18BWixvlD/pzqjfiGf
MwtnyxadNAbSmcQz9pTWON4UQOpfVweyivg5GIeAM/9G5Pm691GhdVoaqojcZZrI
uCrMZb83jg58X6ZD8FauQy1NJCuT2Lyk660SVpcaAYqGJMeDRU1Xth96ETNOZ690
iPbtUxxLxKGD9KuMXApp9l0fm227xQi+XTbo5NVnyrsYNth/lGfES7oCz+sT9uFn
dNHAYP7CtuGWC4aQdkFQ7sRXujdYqHOVmsl6Lqm2ljmRDfeNDUYrd7Fk8LTqt655
oNQrTOnzGOl9l8KMiDs7nMZgdF5I7P2YuidBImTEVx2MAvOJmtYReExk0nzBS1dI
8j7utulGHCQrA2Qy59T8V4rvyxQ+pLO3+iTXULg7MJATbfHueEIlfXPRQqhKTxIQ
46at+HBmR+hP4nREeDshAdyDqgdWfN9NDhw6N5Ag5iKc/m+QQJ8eTaIk5s/mCzBv
KyAhMHpEC3ozp7B+lFpYnoLA3qSdsQ+sO3o9OQsdxJ6ZC9RSDrypV8MPsGPpYBUO
unOFa8rAdrG06Obw0aZH1AFNJsfw/xY5C27Rg+pd1xr0ChFYG7FPjRHXLSpnucKr
ShE83DFXBj8USv1TZREGjY1JAFYIiJ4efSMAzlTrLiUtY9gv1LdObhplIkvKQpck
kkhpCEqBHSgVsQP5AKJ3Zud4BiGRrPlp6gIEMXM2Oo/uPqYyrCO/GlqOJVwC8lrQ
AicraY+sm08/PuF5xPIZy3RJKNvUbLfhF29CpEK+pbmMomhsc1HDBIzcllNf7Up9
hx4VhqE7+X2w/YxqarR/XDiFhHQfR9rajnhDut9ebjU6/hBIHwSoA5b2/lP7RGP2
ehK63LJXSeG1qt/SJqNVv4RAMMYX8gmqiBtN4gVWmCZIQzu7GU/daJAdzIJP79IB
sn9CoG64lb9p5Wnu2bn05sYASAmrlyY/eK0q/CztfK7pbzggj8VwGIID6I8kn4Ao
iI7EySnMVrx0EmgGlFC6uv4YfpkRLx/soCt4GIdE+MlRWIAspjzW8YCZwc/jZaHp
De3AKwGtTBpQx9RGMItihzZqR4IGphkq+a24K4EVE1n64eKl6c3aAuXZL7iklw0V
L8RUcn6AA3BrUXZzFWc50lQ+P3L2H/b+pgF+Tb96iJ3rO//v4LB5akZ174nO0uDx
CxQI69fM/pb4caPIt4GG68qpb/LepRfyukwjbzLr1UKBv4VkE3r1m4TeKrhzK6Xs
cJp6VFZkgq3OTtH/lsPc1CZb/CS4tLGLGKS1N58Ht31EWzPX55BXMOst9vy518Ia
N0MhSM8BKWWpD7FP3VaNzIO8KvvR762RnYZ5w5XtulPY51IWUcsbisV7fJun5mxC
e0H6ta+ay80HdBwWWyW2LlRV9NA+UoUZUarHvtsCvBHC2zQnd/m2noPsaBHEgVUm
LnZnyD13auK5srbykHp/2qZI/5qSseLScAXX+dUb6XwiKujrlKEY99M4clbIG+rq
zwzk7eTpbKIB+5oqRhHcN7gc++mkk3XMU4XYaq4FsTwO9mvJQ6O4dAXc4HfSztG4
E1FEtt+bd+uVZL4heDq4yiI0FkKd1mp7sKlPaFCPuvU+J8W2o8s+qrUuKeS01uzW
u5lucvB2xh+ULFD867+n5V3VNsuPeUmsq9hpM5iyXhvZWegeB5DHC2ZXjQgLFVfd
iyzE35q10I0K/3Js1saoCgkmJN/4adOGceRz75uOiEv92vNDdR27GShRPZNcYqlN
D9aYdUFXx8wQVVUk9nLBim2gEtMc++C9soNNSd6DFT89pF+obgsmrsvzRhXdmjgD
6GTx0kLhMS/5Mm99bY8SS4PU71VkifOLFTIZBpFBBCdq03HwZF5/G3ivES4Sui9J
UOJnjJgpPFA10wKdFwS6gIxtdQTGPt3ab9r1epxOA8YC6uvl59zykeLxXPzEvMm2
rTDk0h7w9Be52ML/LzUrFCkpanoenA4f3oLxXAVkzoF4M+6HH5SETxEQJ2hSqB0T
egvM/DXwnDaNrcsLsqwxFOYV+OnOnKNpYM1TQpF/O/P7aI2SQeQwbumwKHajixPF
m04MHDOMMowA0hUJGMbMUNKWvqVWCcw/boqE1mY3nKt1HCzB8RmMeNA0gYlkVooQ
oXDOfCOo6tThU3i3h0v2PXCdkC1sGEK4lHWs+3RSWpny8mLxxMWPYRxTfPs1dwwH
0v4ZidCrDRmhB601V+Sqx3Fdw25wGhbvO4ODoZRnOLMZd155m1+0x+H2L1DLlycT
AbS6+F6s6K3xIkjtrCbnxqg9Ll41PwOsPLuOArWjIecJ67wREMEdgqpXJGEmYFxE
uv/o9ZzFgtMs8flxV2E9lM/fMdxuGaS9yFLSTsmh1yYKk33XKcmXhUykisFCw2FL
l25CXEN34tzjxZ6cz6ci3+y2dQuPXerp1Z5f+WfsmiLzWrBWolVAaEQEmj8e6sRT
g7Zfdj54bxUW2AEMVaCAZPoXk4B9d2bTTjgYKv/R/DfCXZEuPydVsUhC6x8MCav7
azRUCCO6CAc81jTgwFPOI/IBROtJY2QYIj9HA7HcD+WU2vj6a6BaKU/WEZqvKWWT
hT8R9D0iRTnbEeSol4eSGqlE0FNbPLQxDXmr8BeUjgYSI+Qj6ZAzO559xj7EaTrz
oFApp9D1pv2UdgOPnZj8m6lnXr2ObvzOYARxnw+kkOADVT4L88fQF7vLampkaOrf
nYldwQ2YnuxFDMhUJoGy77u79mxqZlxoblC3kaJb6ZiaK2S4SxoGZbTJlc6QW+6i
2jRyQlSBu0Ijy7t8n/d79IWs9eHqYV0IKIwelnorgwFU989QmFp2Mvqq/8rjuwOU
aMg97aon8/DdeCbZxZHladhNrxaf44rjd35wbQ1arCrD+nEd/rH31dPNeYxaBl/i
+ChqVfcG8NMtI9DmM2uB1VFd3lzqkuEee9LH0UCKWGD/Xa051PKRX0+HOuZhI2RG
+2L2H7U0IGP20w1RtIfwOS86c6AJlbtvZMWc6z0poiYJeApF+o/ITShcTxcTdnEv
xlNuf8Y6XwtgYxLgYvr8pk5uzpWZTQzkE4G2fGHexkslwdXQqY9yQkG9SnRIDu2k
S1zIyyhgvuD0AKfQo1hfqL3SRVqxjKSrjx5mi4hhquBjtXf16lXdKZy7hG8Bqo1S
xK8rNW2yCNPu9weucnUOkMg72jVh4Kj53FZy2kZ+/lk2NBEnpXkxZsO39bJInzAs
5TrjVX9WYMQn0b+AJqqLWtBF83kC0SUYjaoVHLC+Evx8+AlP4sZTvILHqM7Qpb0C
ZsoW6ZlBW1MAGfC7EsrLPGX7pJd2NF9TkZkymdg8WcoMlP1Y4hxDKX11kedRLR79
jwCIhxRUsaZJrhrBY146eKo5L2WQEMfM00Owone6JTvjPm0Rn6KFAzIYCQ/B7pPP
obj/1o0wPIgtsolbBSy5DKOfVZ6bPbJwJ8WOa0C0BmcCsld+wmbNov6zrkvY6Mo0
yURT3U+OXX8AK090qwDb53wgc5mMbLZkDeeugMBVbwY0Y3szsyclIzqg/S81bJzy
/dbSD0E4sK30dHBjzZjlNuscEnNjiR6qcGmjiYzztltcMv3JVg1M8OIL4a+U8QDw
KY5ud66JxYpbPSoVNC0l1dqQb5FuRDFFPcZW4K6NRr2UHf1sKnIjcMMI2ADAg801
2IUG0kg3zqNsIyrpbWVrVUTrRi1NjqQ+qniRCDZ8/HV2wCwaU/9+1ghsK9NxWoO+
kVbFocD1IraAJ873vL/89KqcqOEKCUK91M3IyqZdv9FHxiwlw90pKWcbwtEo2/hU
OCQvWu6XJfAxIBm3wUNzjj0/1YanVBwJ0ZZ4pPd+n6IAYmNyWX1OtSPKEaMqkg1H
iM80S5z3151tVDaVskidkJNzsPfVmfLkHu/rPBseBmUoxWO4JJGWiHBmnvxP+m6Q
s7Dmvla+Da/hCjRXZORwm5VLSFuP32vzXvC48kSvQNYnGS2VGy965sxW2grSKHM+
ah1IwDudcu7DwWDtDZ25u8xzoaJVh38cG3H199hI36WH4rlSgvtXwx7t/cTXiUky
ssjwHk2gJpTJgyXKo0QvxHkVcrdgRmDZPXtE7etpSG0OJk6Ky6ep0SCCq21q6EmI
SsPP+X8CUM5htLxUvobuFdavtg+njnJBdJkVyuoGx63hp1RhJkL6rZKb1YP7/RCm
+fGUaCh0nHrEveFnvGXEdXWQCRXlPqrYcIsE/3P6ECAurJ4bkyNY1iswgyiaxshK
i1885Hyo8/9u5g3oExqRBGotSuhF3Hy4r1pi8gbdZPt4K75dMg0ava0NacLFOgac
9Bg6kMMFIPS6EIF51SD/jNeVXZBghM7BWVRYScf9iaUOQOBK52mz9DWcRq/cbiaR
Wz9o2CONj9gP4I08nKaX7pF8k2WdWgHV8ttnjJnyFHoS86ZHf/n/flZ6GdgzoYBu
islA+ooy8XU3nqqWV0s01CCS6sWm70mqfXGr5302oYFslffC5gXErBq/oRU7Fkzp
oR4GDGoKEKY2FiL33UN5prmmihbi+ktzbc44LLRzQnD6JUdhHM8gYifLh8rLvXEx
Ia4iM6GikLTujGjN68PJUP5vrDH4NZ8+6EOS2dPrbKy8EBcaqdF+PUiVvgXjP1wD
lUKPz4U+qqz7yzNdCoBz21JD0aRi2bBi5mQWEVCXW5NIGfxQ2OhXT9ZBNfTsGiqb
TpHCihZHQVQIu08tK1oLuhnHgYXLnSTMofoK6QYBER0zrLafnDyrPeHKm4ukGCG2
1el1QUyBlmhGOO2VnAWJAcZQvAuOg9kBCq7pudv131Wt1KOewAp9jgAN8Nk+vG0I
CkM/rgPitxdexi7ZObnGcm7XnkECHsW67DkOSHsGCQWaAwa2v/lX3pjtBhyxOZ4y
Pbe914JhGBwHvK7SafOcEzDRpix2v2EUALWA5J4jiByBZhDcPOLWoOGAU842QnyZ
ENh9kzwG2NzpN2cvFaWPO2FH6oWYUPQqR9u59x/ON60cnuvhm7/eIZ87D7hqAI7V
oUUuykFPsjxlF4zpsuwmz7R17ICyzFYZw0bY6pdWcocELvFImb542dw1ZPkMOzji
o9Xrt5el5jCfO4QdKaIyA4d/VpyiF+olp9lY/LbUTEXk5aK7jA6JToS5yT+VDgv0
5F9RD0Q0J0Wi89TXCAajzB3ea+fw6Cxcy8rveEMMq4evVJ7+mOeucd78QYc3gxJw
y8VwgLVIzgLX2YGvcgqKByvLHfpBQMVM5HF3Awg0BzcSPqhZVUo9sbtzDorK80Bw
L9o8ipKF6c/eqsDvnoJK+rwU5Cjlg6oXeMoEVh94OvbBa3DcT2sQzkv5rHxtLehA
qzbVV5fxx6rjTnjJl4pWHNANIUaXEZhEsaxxFegxyyNlvaG+cmO5rY0R8AB6vTdX
iYGXgp63727PwNFkvYJPZQfTUuqfxqajNo/fNCIrH5hbrSyWvUNb9pBYKxcZxrib
WRf6Ri6BBPmcJfdNhNjqvp2Q8/rYoiDhf1hauiAPydd0SvmuC7RgvRnEBi+fH2/Y
irnGEReIuVy6I8VNxLte0+OIVQds9ynUmfILuHT4BKwjLG+/v3LrGebcHF2ljd5b
t8wl1nmOMmL2NTDbcVjfiVaeezgP6jFN3i+4ay6PGU9Px2T/VYzv2vbQU6Ks/DB/
8loD9A2mSST085Uiqz6ar3gkYQTKT7qqFeuh9NNd7YM0JmXTBsVjSY6scrOI6zwf
GowuCsM2oGgjFeXfRi09nawOPL8ViSOx7DIxf921uYG1nW4PTk5Xza2xNRiCKdeD
lG3Bbib8aByMvhQZLulRX8VOREmBSBn/icqh/w6zIHwj5ScvOrmJhlwqzVoZzM20
E4BMC6god6TA3oVA0EwuWwuwZk32YgcyDByhvAIOzArgVtwnn33VIfdLYZSXjJ6j
qmVAQzN6LXC28KRK8AsyupEY/YRu3jLJEmHE1MIZzcwddYlWdc4F5uuZIr+vJvMm
ov8rp7wydlUDpzEr3Io6plm7W7A8lWT2yrmFcwF+JkZPyeqRYFAk9VNymfRmAqT8
zhC3Fa+UAM6ue6KhucJ3nf9dDO02TVTLwG7uZF5tYjh+hymXhlKDc7jNfwfF6gg+
S1+Ikn5pCoPJGYnEUqkMmXMBDvcGxeIP4yoFpIPEh/NV0Ims2ov2+EaqQWEADhcu
0mCA3OXp/lomM0ZGICBOajp1MBAdEFJRgpTptfdgU++3TOjeXYZdZ74vqb8Aqvwe
FPTvCsjki+DvYun0RGIbPLy/HD0tbNFNyv1ZWMLu4d0xEAf2yzFTbHJ9n4lGOKo1
voGoegIao3YHZb9piRL5uKeGbeMa2obOQ9Ex/71WgiAHUWqYGMaJtIqxasOx7qfp
EortaobGFCbfuHDWCxbkrVmQCxE8RTwN363gHJsUPC+rcPbkoyydcaPh/gpGH++V
EiH4HLtDWkxPsJVmGjfWp8BxE/QXOFqhVPDzdt8S8BlwdudzpfuZMaCMWU6HBJay
dBOeUCo8uE9ndRiwP/+fPUGng9XsLsu8bsoWUg28W1pTbLO6ronpfiRgLpfTg3U/
jRCibSSxB+gc6BUNQpFwsMKuStb7CeXWVvAaW6VjkBgQzQamVhVWcoZ1BXiBQJcu
R3O4+Drzm+rnp93rFdTgCVIrJa0st1ibX0zMotZm/Yv9Wt0G/tC+Qu7or3uQ0pa1
HcRRTLFAc1MDRDd36wESOCGhsIHANtgAEFJDv6Qp0ZxZ2ffGatS9Fh3TcLmEEeK8
xU4BwuTYENkU8Mm6ZYGwZJjtAwVKxD6WEBUYaB/dV0LDcBFRFRJzjaKtaBqU7NL7
Mrrtw1dE1qq/hILE1u0kwoyLmZugltYr6ZzhbCeHNudvxA1kcw6ElHWVKcxbguA1
iafB+b5Ba6YjKr3y8WbfH/yc+pivz9t4qIUVLuhB3lg8OMNmcu8/xM1uKVAo9cf1
sar+S/wBOsZ7aY7PGSldZowadsnyHoLZxxjPb0gtCSdIFAVtpkhros1s/mpF98o0
QWoe8XHWNz+dg0KYSTsvhCY8tYu+0rXU7B259nBCLyfe/W+zj8oHp2sq5+6srC3V
SLs9aA1aaDcCxlbyG9655o2N8MAaZ6ny3/zNdU8bz/V/C19CUXnQE6llnrK2f3Zv
fS16H6dAD2B0kJooPP4lgdxQ7+gLbjIb2lZvoOfyLy3PcgRI74wdeAhOcySNw2CU
lDL8IbT8ZGH4CjEoGPZ11g2ZVI+367WDG4bqgGCZbnATqV2VKWpP7HLeasqqPTzv
mrFskicvhI6Jb8N9lrs2Vc5phfAbDb1N0W5ZWWHpYnH6P5GnG/mRnmjqSqlsCvaH
c0SZc0iCMyIRpYJ09OiTc1cSWhw1AP5cJSQDGi9oP4JvCLaVSdjtvGqfraAcWTKR
qJOirg7mjyeoTPuUJkK96lW40Yr/a3Be0fI8uIPsmpzKi1gS9wWS1TnYnmHRuH4F
4O0Bwxp0WZ0k0OziHnW6GSwqi0fHsw0mR6SYacXYNiJBzqBwB5TbESVTM/wfphgD
R8U5ruaSZpzmUb2PY8zanKv1pZURMjtw+3jaT2YBYP5WaD4Q6ICsdJw5TVo66eEx
VkTdvEVkZL3ePu24CvXJvDesdl8q77GLdHf649x50XeYxh0bdEvP14q04I+eI9dr
zKMmo3citIihW23FtXgeUi1vNKfmsg8XUo/suUXplJSMXHeLSDQ3H1vLtXVR224S
QFPZfI04kxjHSNIcEL9dXWPsKQZyV3VRVbhy5IHghRsMTvIcoX+BqVHdx1izNrDk
z0V/2LgXbjxZUyGDaa8kO2bI2HuONbdzDr1ZnAdr6ktR5Mwkz/7QyioXAPT9VcQi
3iJ+Ad/f0OTOUjVPt1DkA+Ic9XPeEV1jKDNyUPpdoNpbepjNGGV8CB28szmggon3
YkEerTFL/La/E75d/T1WcIWUKMXkmWu+kdi6oYhKeIvxOji4fc1En7dI/ng/Blw7
S3cW3FwcSXXJ3O8HXGy1/sc39Hb4phv51O68cFMj0P48p6eqWmNMxa7wG43BOP6E
xeaItA/kZNQ092Jc1cAf21GVLbosTjaXsD7jpBCD7xgpYr6JB6DpdkWG5ZsmF8qY
+9De3KtZiDSqa0uVHo4ME5bXKIX/Tu8ilfAR/3aXwvPLlw6b1bshn4ZOtMU71ZdB
YZ2/zf7e6FPYvoO47FlpQb44NJZJ7qLTuTJeX0PZIMyKQfuZ4CKinjQ99SUQLQLJ
Jgqsany1LayqF3UdamTS1gV19DZzs/76dVqMb6rR60vy19suEQtxjKgogrp7VvPw
PKu9/oX2WatJknLvuPD8bJN3RzAEW8NNaOqSS3oPnzuM2VLPyVb3/8yqEq5zFpNJ
FFPuv74jNa7tIEhmO9XccgRynuMLenRQQVJMhV1WGfnqFicHW9uq1C7h1WTWgbZq
8uYzoeJ8hikGYEgdAXpYBFBywrUH6cvy9Av6fveLdzlWGaO5WN/vk5TTT0qGzsvx
Da37pWMLGJyz9LmPM/dc3gkiL5ExIruoTU/2sKaboJFygejZqtLcWorV/QtOiaup
9P9yTMN++wjqx+BjIrZtPGjwgdJZmGOisGBGxQl5eLtvGJg7ZTCAOh7LsVZkDApu
9XO8i9yktt1NbWmH2lCj+MQJI7GshphqLSLNy9IfatbPA7H7mOzkuVh+Rs77mD9H
nW/HMUANSDcZhQKak65IJpqgpc+qu+F3xXHBp2zsr/QKTnluTnGfK4mqRlHBIJ94
nZyN2/u4soNwjx2Q8iG+YZW0ytEU21DEcAXMR7sVxLDMM6CR/5xG03cidynaJtRc
EaTZ9kfFFw/kws1iY9GBSwvQF+ZXNRcZgBcJZCwu318c0tNArbw8S7MbrTovRngu
nfj5QdPzXD9zEJropYlU77DbPt3SMJmQEk7H1FitNGMokQdL95E0SoS/7PzvukPd
2ZuTpairl/uU6oUNNgb3Zt73TDsuIfNnRQevHbVdEbY4F/W6T+n1pXXPJHC/rpRn
ZkQoSlgxboTVGW4dlVGwQ/rpPkizPpouTnz/LkK0GmNO3fylqAefak/79Zvtb6Ky
L3SmrkUKVZxDKDRtnxKwKDnKgQtpVT0qfUvtgPreDlkpn7J78oXbES/XN4JERIe8
pJo6RJPxFVC56/IMHCUg9B7NFHUqaNC2LxZEJbJpi5JwzPz7D+GGe6IeCQIVPTQ/
r/1cRSLB1goWxAAsPFL1RgRwATEqQC9zNEchgOIDgq+eKYqfzT9xAIg1MwV0tpNM
FmI4/5J6MQj3n7PJpl5AtYOrYnkp6yCunIxGDF+x3XACvEJIuHYaojIGcsUHfRMD
L8tl3svJgPDzxP3Y/wDNOMxdI8+0JPJKrFYbiLuj6qM3D4xPzbb/gNYttdrwnPlw
PYWgXyxA2pIwiVDtJSrksOp1fihhdNXczYU83rGLjPrWKI38HTe+AttTP2OufwMh
CPqU/OVoSo/KIeCs9/1yFOdiyEmRWemTZ9y9CWaxmkU=
`protect END_PROTECTED
