`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tFLLyl7IwnTQ+NgAJPj3EfrPdsO2+YV/4WV7RhijBifJJ9+T0Nl911VfcqIxw91m
coAfSa3X6d3ieQydLE9laKekBMNR9JNLNo2pUhIMmwEMsw7+ZujLeEsQp/ghldLX
HpEn7iK3VE+Ovrd4E0GpUXr+y+NsUem80V99L0eNwv6rHqRqd72JQo0fRAw8olZS
ra5XsViJpBR8cvUPCWIxIhM5dgo2wH7xEtpwkWuu4ioalm/mrEGG/Rl5tCGckkw9
bTDGW3TT2K6uuhCdUVk0JPjWgwRGmFQYL4UbBf3xHKuFF3iQ10TFIYVI0UNpBZhs
z9jzqzj2/sJwLCEge47fAtDDvUnl91grvoAwAvzSswGVxcowHQUOxyrMHraf0qjP
Brs1MOBZHe1o8jXksRLwMgfIzXM9exGpEIbYihg6Tgc3goh4/4vk3D0RSzdOWfb8
017vJoeRjvTsYKRoHknVLhoHQ4zQcTJx/lqdI7LvTKH/fZd248x8c8gAVV28Hixd
nITiTdbIZwEEaFa4IwRLld5pAjzVsuOwQxQsAxPWi8EOjm0Zwk0supq4lpmH0RMN
GNQdIoNfWjcstT9hML6znf2Z6lqS3laR9mdb1bWlRKJywb5tVOUF6O434DFMjjLl
x4tjEdLnpvS7Eu2t/Kw5Tk3ozOsIU7EYqtTyUuBzPXBrGjTka3cRT8yNo53I6rn9
DD7FWmycsvh/xNMYH6ibTeh/UDToSnjudP5Km7yr+NO0Tp59xcf+h0sAunmFgsnH
z30fSbia+kAMPULshmBqkM/KPd4NSJLLBO7kVKb3SDGT3d8wvase0AWZsIcgB0+t
iU3CwKUUqRShl+8hCunMtrRpNA/SG8LmayPqpWEhCaL8qZDl8ttDOhl69ABjywxL
p9oRaOQO3mhkjj62AhuQslGJptacNT6Wz8Dsx5C0IR6XRMYX+dKYwQqERjlsUG/J
IMSlnLZvPMBhOTnsagSxExp4brTOBGjerHfQS4YcLrPDnG2tauIt5c4eHgccYGLl
V9Tpcs61r1QdWqiscIpePfHX+bBakcCJY+75t2z56Pp4VMrSDBGWaYkgtyPSCkeA
H42hAUck8P/0tF42ZtQG7+ypXDoOi5YBxiCKhh9+8vLHfZu6TyAIfge317BAsVRq
5BsGzwanHEviqfswl/G2qw5b967kIBW5KzMcz4xZ9Q2KwhJXB8mLAQaiJNrEFFsu
5E8U82ca6MxSagj4Aqx1WbpdC1e2Jkblq0dEugTd0ivLEDfUkp9nZ2Wb28iNtUH4
BKo84iK2SSNZLSiVGXeaO0gsQSuRhJ02JIieAO10o85dYWetAR5yYomgx50rcYWO
1OT28GvLkoXYjDlMKlvmf9aVNwjDYUp5ZUPu9uYh1/E292JH4/opDAlwGXcILf/m
9AhT+OIxbba+P/kVO6PmoCjaUYT2Z2qn6kcR92EX5c0ttALpvkDy8Pj0Zq+sAIsn
KhQ5f6/4WddEg4wiYLd65g5OXdrogtQcqYiCKd8/P32Shqt1JR7jdTp/+ZA8Dlt1
W/WFskrNJAT5eT3EFVH3AOvSi3cQuC9IT7Xvq6wwoGRx2uXAp9ufk37HZrt6Gtc1
xpY0ADaL9i2AkDIG3IvLM/BKNIMVBW4z3lSl86VjyPJRqeCQ+/qj30jh94cpUA4n
yzmcnE+cS8oopx5mX8AXMtDlAvl1T1NvWr4TPVLPiGeVvWWDfePyqtL0MiBWi2mG
FHdlvHQl7Fv0hXMgqNpWf8glhIwlOvnUVSL9gsH9K4TuEc7hM1FKjEjjqtHR8huj
tcHOJu05whQi1/yfeMZe0zlIp4S12qZauDmImt6Vby2P5WuDOUvdhqBsk1YIZxHA
jcVTl9DXtdgRhFpN7v4RyYZqL8hisrjkJaaSCSXW+iNgXj+zeEfdFTekT2GKjyBG
wlym6xhjObkLYtfjtitrqo96LkG2IJTXLB6mTqDKMYB0H7bK+H0eDeA13R2PBjS/
`protect END_PROTECTED
