`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0jpF6GNLD8U/O0Xb6HDtqLNqH/ENnR/aGiNu4Bp7WRY2hhcQewLeosogucsflK6A
7TUjgXiYNvvaK9/Eku/WEI26mheGQeAESYFWPJO4Iof/KhuXbdASFWGjxizx8eJB
8suHNnElD2TIf81HIUzOVRJoxLlDM/kVtc2NELt+6WsxNpQcc+4PA0499ommXoeq
/S5Bz2rizsnQx6/mE8uxz6UG6TaYf2aQEpNU39Sm9lVxbBFpXFoXJDHTQrpMrBDI
t4imSsia8ilKpdGAfLJoDADtXUfOMSdHavdXSvvtM0UwMm/Ua+A5Bha3LoBcpbEo
JSrCRufaMfrVKJQWukBEqwqX5KHxIb2VeNKM6bFQMWVyLWJ+JVn0NDnn4Gv/5Hks
ZwWvDk9M5LxuDidWH/vkJQ==
`protect END_PROTECTED
