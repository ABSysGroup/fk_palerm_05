`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zlR5FY4HskJxCIsropgeTu6TR17xC1ZyrEvkYJe5F3TYXDI8zYd4Xsx9+Lii0znw
0v2eJZWhAAu+s4lPd7rAksGGrIzj8aq/pHKS7DUcbdg7tbDJq5xz9BsFLwpUboq2
XO1uGtoEqVMBfhHR+OwDYHdFwNOF6vLy9actZ/JwLeNWni4r1QVClESKRYa9hpyB
UJXgrQHEz36ByWOECGOFoOEMXXIPxjDsmbK5/sGoilDsxSlTk6LbxoMebrunuImd
2/LU5zvO8X92hypBMUF+8S/FS1Kp91iBUcMuzvf0/YiAzBhVYn7RkT0a+QQO9qQp
S1DRi4GIjpBJ73pGWWwl1fxCYMD5ZH/5HdonvXg02c7ENCP6TndpajJpEPI43oVc
jbkn4IrryXg1x/4lj/VO4ZEweYN09VyvAj0uhAY072ZeMe5staPry4Qgt2h0AVAl
a6pYIUrYF8PCmoDK30A+ZdrCmEUDrh5OaX+ZTY1nsgA0a+73lCFDZ5N7xZbv4DQP
OeKhwyyPpiMQpUudQzeBw4qeKSZ52bPfv/sqSRneB3dFn7OxFCgk9dU5RYuZT8YN
lGFgFy4luyp5y/TLZzdtQat9EJ/9bzR4qSAYDZUxHe1fD4WEZfW7OCcKbZIL6ROt
t1YQjsfTJJXWZ/MjPYqFiNhV4czcdDTBE2dXe66kne1EcgQRZpMMoF2lQHMU77ev
FrgX09TWRUwITJWQeidmD/TzVygAPgy6dJiXTmrohIApucCYjmBYJKr5oWv94gu6
0sTWrrWad/7sJ6gpjv7ggv0C3cikosR+N7DxpaRl67N/BrLpl0Mldq5R64WqaL3m
QI/tfe+MFPTHeb1M+QPnkavlIpqSqYTjnPxlojZRwTWZZSnj33iJa7YYTL96jHjE
OpnQ6/gjvF/a25dRB2hNverBTH/srFBU5rv7X1q6SJhSQEAUmgBeG22oWRl646su
uHlywSlt3U9iMwIc354j7DXJpAnfo+6D4y13xZFAdBXqOpA8kCk5pqe4cIdDQfPW
0O5gPsWpTuOgIE9KAwh0Agj35yXXTReCyYUvGd7Db4sKUukbXUfjginJiLd9vrKM
/9QcIUFqgWTm9GcKVdivIvPeXKOaOf4m/m036rzW6RO4AKu3AHbb0VUqWh9eZchj
TTUnQe7XOPcME7vBAoiomKYYF3OBJbHu6bpkqs6gaie04wy0mY7oW0r7dbTQcAF9
FLLTrD+qcc0O0lm8zRpX6p1IkClnwYKYruJCgeTBKHHG+l+5Nrmc6DzkDBeK31pe
zskljGaZe71SJkgz+RSaY1ceDTTP4RNyNoiyG49S12jOaEZ8f2MX7TZ6Ykyyek+9
BDXVOmfy6MfTStRhVYNUPhfD1ChRTjXejvLZEweheMIQeFgYFyOK68EAjcsLKvVy
kNEpX6JNTvjUTQIwLQubzIGMqMaqIu+p+u8C5apdkCzU2WQzE217jnWgshYYkkoH
mFBlkHVqoVo6H2IXwF2UISNGyVZKdEmW0Ck+ifbnl1/w4NCbJhUpOPA7P/dJOxaz
QiZkf96emvGwMkaJnMZwZIEAX/b7UZsBp2HmjdhbjoqDsdirvWMoulzGFUtkn/il
0KbGpdTx743k4GvOxJ1bApKrbKllMnL77SSl65wCja3HXkrgGqVkIybDu6F1T4UB
ERVyFJ8/k5nEes8D2069Mqt7mWo3hAVPl9w+7c4ZenAizAW+YgW+d9FiQjv4QKn4
lpr5W2BqQeuDC+nNApZXcpNfJEkWs30VU37Lyde4DonTYnYPF+LMhyVpslP+W9Ch
dhXiMvb42hIyRvPRKg1bBSeV+xa/VjhcC9ELBy4HXKT3/WQh9hkHnGpRokh9/04X
WswiQcXNzo2DDq0s3zB9ZKKfZAal7yvsp/dKQRs5RhhsKQ1EqBb40jCBt7P82wGa
WEakF0JdvtzNB+dxr1flmQJUmfBbqSgV0EvH1ZvTpNK7sPqzIV5ADKBDhGrwflIR
By3eY2VngD5vRv9DtIjjlAr9tpbaUx163JUTMnzACoq0wzKySCsmxrKokLW5loQw
kEmBv8/8UI5deXx0gEHh0cA+kTIqtLsVBAxOKEzAQSvPMdv1mrHlHpOvhJHnlHMh
TeAlag46/JqwK+7XJO35sGPy14o49m61Ay6PsASg6MqNQFDg4yWa3rrynuhIG9nh
nK5pEyszUpkjpG+/u5M5J4HFGI+0BBIWKgi7SuGeMycRTXgc4nhXDN5ABmHnhUeq
cOz9xZWn13KRiU4umpNQrYjHknOBEN1/ZwvhNoOKaywZt662c9bcu6IVllzQZMNL
94IBQkziZvMX1lGl+5qtCszH5sXfGgz0q4qQ4Wkm1XvBGEy9z1PswHWqVGVJEzn0
rPYoRt/r9OV4o+ozZD6RiswZUlZm3OZ2bsSvdfJJfndROaO+rQhFKmrwReBqL0PJ
H9izsfRv5UEDbif9zPDc3GDIgiUpVhbmSPWPh/oqlhGH2Oyf/PHRev7eVPAdHqfb
zA4HLGpb6pri2sHRVE88fF79vO0mBdZsIEHyBvGmpmqJ79kXSOGfcXpundeL3H/0
lKJDjeXave8rismK7DmnsDA1ZeNeafzvhVKyOXwCI0V0JRrAopr4SPzBYo/QbPRp
prSwy89vnk7TnSGEWipJzeKGvrYHn3fdHdL+o+JdHgOsvRpsb/YRn6eYpeuWXvMr
wd7T07WbWMoO+iA9kMjxa9QIATasqFbXUR00Ho7d89E/wH0Xm/I6h4zKXSwMyQQr
ck70dlfvSDVD8jrQwUZ/oIMSuql2PyOM81L8hAkh99iJ+p8gK152xnaQL2kSnrxO
KoclasfV+6EcMyW/QQVk8fHue9UsZn0MQUM454cYPkFtkp0q7AA6reHFi2zAezEp
KH25YosfbZvRiklAbpqveTQlnF2AD1BhXqekmv6iW+DRNA0amYzd/RC05U0OoZAi
/xSa6qgIWnS0HHbaUyKIPEZt+dUhQHWYf/S58/odpaqKZu9acgC5Zj9jnCDIvR7l
UYK7hpzNRc2N4m2sLUIt1fho1/kexsSbKjTSeU8aOARMWF8FOsx3Un7LiFBlARj6
cO6DIzXjbmzFxHBbzKC22AKimRdhBcycdy9yy0Sazah9DM2Kju897SdQByNL6pNk
36HONi2shXeMWpmq9ub1jiJZBbS09a+WHEb6/c1OizQ1eIR6JDm3lQm4Fh+RzY0M
1sj0S74FVd4o/m2wbYHLSM8/Oi55zOSjeDVQq/p8TDWj6jb5JFX66N7NKLgq4xsw
fi2m3N/0J/gj6Hxih2f0HP5A+LLzdyY8AOkRcTYxGKpGigCBwnneDmTtL0kbEBjs
ebG0jvdSgZG2orFw1hfJqEVAHLzETvU2UY49ZnGnnfy0CfePP/UEITBXZAIcCVsL
vXaYwP1qnmAb34Tm5u+6krZvaMo2/qUgkZEvZGmSTVsfjIusAZ7L4KGy+dPjMLGX
FamKF/u2Q7qSNBbh1+v42mE54QNjR6Hx3lr82QSQHI41vf1K69vvtmqdWNmZT8D5
tAF+lSZkGwoAilwOaP6Ofg==
`protect END_PROTECTED
