`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G5UHES0eEJf1RwmI2ohnh+8ZXmZHCRIxMV2aTXX+tkTi7yz1fH714bzdZXdtB17k
Szs7cKecsGbjYa9YO5unhb4M3jLL8/WE1BpQYniiV5VW2Aym1MzGtkiV/cXGAtw4
bsg5A7yAL9hdEfHISCtLQjkiLOu7AJ4vDTVstOVEU6bpFy4mmNY8VZF+JKWyk2D1
3eJDYaf2ajCsZ79cYGnXkubvGAFOhq/ZEt+GMQtF7p2FmCTZSEYSYTKFrRD9ETOs
GOFZRAzHTXLNED+CCkxrMdh8CmL+ZZqOQR1RdsBFJxSyEVH0ZlIusd92ZRQ+uDFe
qu1AgITtBvW2o+aslBJwL5aHI2DHPQ1tHp0KArewn/GssT/B1oa0QvDTJENDrYR0
5CzcXsjnbwTLTXoQE5EBL0FgKiVGa02rlvWVYMSIHeUbCdwO6gwGiLT9V3FgxF0C
`protect END_PROTECTED
