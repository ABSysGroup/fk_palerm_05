`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
03h1J/9WrBgp2kA5WH3YKdrYkl8L3PaUGQSbViWltYeQx7qjWIZ+La6oq3HwD5t0
+rW5Fh53xZdZbn4zsxemdSytex9gieZy9WxKLs6YLf7npWrodU9sqk/sP/zJ58rs
e+R/8TM8EOb1j4v46X9g7KesDqZoGMaTAyx1xohqcYlk0bohJquf8Y+nlvUQpDJh
2tyukrQbijQMPv7EX4Ggft5mSLkjFPEQPDhGh4vN5Wi8SCpUTcKmd/9taCCiO+vj
HQo9uURg6Kx/eOy6TkumUJzdkZJT1TJkuYWmStOR/uPhs1/24H8yaYji9jcmMocj
z7QrGTNrdK20FiK8iWSeGgt8K0uGIYqUjXQNKEQJrqE/AhxefP5oxwjDCrqdgapS
hHMoTpPJaHj0qSECpc55U3AxBE1Pd0hPMTnLL8CNgVcFNmupxDuWZ6kmWY0KgaEh
tphpb18g88O7y0BCgNa8Mjgu5rZlYYSDIgQVSiBfs2Y=
`protect END_PROTECTED
