`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IvAcv0JE6tWpMIoEfo3hcszbu3L5P5hod7PwSOaYFJ9d4cWyo1RBmbtnWhZFZpXI
RfKSe+JwfERqT2Cwt6kA5XF265qLnek+VPO6vprAIDaM/4nHTTGzl4lYrWz4zOVi
a1X2doTeIvSMLKZ00UFxADx0lbekoGSJ+KePU/KDC+Ogqvdr5BccOe4DdBNrfp0g
NScdVAZeS6AlbH/yYfNGjkSt+h+5huzR0ipEn11RrbiszMsCErbkTftQcyk9RCXt
IKryubkXzfPrSwzMNoJ1IhvL9BveCYKexx84CFGMGSs8BsxQsekcjJpip8Z1E667
/idPycS4M/HcY0Hq22BJZwIf8xX2aE2uS0jTS8T4tTWiH0+gX+yhl/vSMz9H5OWT
md3q894B1u0Jo2Wm4zU4xVyj4nGluqw7Cr0hH/7TozmW4hW2OM+eZS54Ii+lLYwb
ICVN5aTHmk59pAbpSorf06sLoOMsb1wya05hAHiMZoZ9wtokdqmZ89/I6GyqlF3M
ek50T51CDOoxTha0H0mp1c/cHv5v4MjH+miJjMjtpfGSqQN2owYaJsTf5YpzsYoY
cVh1kHRGK0Q7LuBbDNudIxQtGtHxpq/nvY83al8T/58LiNL5FjFalnmDoGE85eWZ
w0CQCUdv7S/LVDnDN8L3d1z3FdCoyS/CMz5fZ3/nptznfl2UMjGxnYP7pjSu1VOU
ZzxO04azrJ+KdW4f55fFT0WG88PX46hKPqwIVEahnzwWGxete1jleigWTiu4wfFj
zf5U3H1oMO3j7gq6ue3OU8csiaSSMnk1fstRszoECqx0fiZ5H1r/lXLZsis2N1p7
QUPA4R/BOgnnJnp1uA8rIQ==
`protect END_PROTECTED
