`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IfET5hDWjRY/Z+Olzfa4YIcTEGzbKYSGBYjQuF8CWxcVjLbUr3s20TcjiLxL4dvQ
buDcWJtxhLEVb71KTXmO6e5qdKVQXT1TrX67YZzAbdb/6vHwE8kQFdg6i1uUjwP9
bhmeDApo3zz3AOZDkuKEK+K/Pbd6uxKShfh+z4G1DbTM3YpIkNgJNxiJDk03yto2
+W3XxQ72GC6cL7qZGUm6q7V95iC6c4KMDQH8lylFwV87ESlmmNOjJM4lJR/aLn+e
hvpxvAx0SRtiKhl/FemOJ9aoPaCQuh8VLQb+sCEU1D2fZGjzi5gKlxOuTNfDy9ZV
ZNzZcK83//q4u7CyQQewg6FD6I/vYNAPBs/q4RjuXhy54UP/j9lQ0+YbyRGiZ++2
O4eSQ3ocCc9gaCedwOOaI1Ev6msQeA0YPdIRsBEf7lm/V1TsinFqrcaXaLDpDvtQ
RhI7JLD33qVA7enNsDo0RV2uFbV3UcY9xkCPKUQMsMwL5cVyfU1aA12Bna8/VCvL
aeb/chbsvoQWWX/kW/Oxlqxwcs8kgEL8NzkSlro13zqmMqjmMI5yD74VyRw+m0oo
QZzovgP+FLSbxubDA1RQ3w==
`protect END_PROTECTED
