`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7mW6bU2jt4GxehZOPjIFksG0MGvIwPhAP1RozQTX1t6uS96NaM1coZpZMX82UNq+
uw7JbqIHOtMRCMktVhbmjdfI3Cun5sW2bd6mO35O6s00MNjYeREY+4zqZDGbcA9I
ZFxFFEi1CvppvaZeSdobX9s2k06xImPHZxZPiGB0QWSCanjzv6M3WHTz9zMCRur0
CvQFNcI0FnZC03alYwvEvPIanlUKkqZtnYJKaRlQEKc6MrWTrP951MqAUU7ZZUBl
Lj/ophASZEa8ICRLHF0b+xlZBtqfRMLmrQPgkr72ORjI8vbDd0e+Pmhs3lBjQvmT
Bj6qsjUZ9FBDgbHUnJjSazXlRNBHztAC2VR+MphNwX5QJj09JJziD/UNfRcoIiRu
4elnF7Y3Xc9asJ+g7DToXqfDB43/B8A+iIdGG4LPLUXZ2ddqfme9ItkkibhlcHXL
nF6OwcH+Zs7TyAwAoh+SszMk8AWYGlI/yX7or9fBgxqUYRy0B1kpLGTqHxWq1J0S
xgYKuUFFn9pJwFbjJxtTj/aqVILl0oX4nvFlrDMjJv2WyD3PSZ8f8tzy9y4j2JBm
NSWDHt1+OQ4sBLn5GRfhe425XhIw+XuylpMf4GInHo6X6PChOPhusSbGx4g60JR0
9TXuJjtVcgaa7snNG5ZpF4KWa2STccRrFi0738mopcOPrkNrVG6HQ84HW4nwVYS2
rswovKFz2LmVdujCUD8wfs1t08QzhgmGYWtd2c8yrrmRl+oUoOm0nWie9WDGLK16
o7kXP6QWzwkjBnyABgIOfLVNJQAg1XVJvrN9dh4sBd6eCDNZr3z9iP1D9JYLqB0H
hGLRELRxpT8yRcdDimnawrTz5gV+/vyzdfDSMsNA1nTntFDLjbgdgoEtB3+jHog6
Nebzh10UjVJPwSrKFF5/cc1Ztb8ChOm1IE7TmrNhMl8QNTk53WQ341e+L07hbaEe
OawcaOplUrE+rIU8WxGhMIvbocflJHuLeW79HGH0B2SnNCsFI+Iu02zfXJsdhk8k
KvxJsAqR74mfDnGJr72jWVjF42Lbb+RFstA4MFPP63uDXu+EUO27R6igx/m74bz5
ONdeobJE1GMmp5KCxGLS13T3pS0OiRn7XhYn2wTRqHz6OsQW+ySmsjjLxZ+NPiVT
PxecZPY3YiIS+ePu39srp4VqdypVn3JRgumPVT0nCB6UoKIq0yeiHFOeLB5Q2c/m
PtqfbuNYXQnNwvzBPoYLn5uzoMOvCG0Wy8lVjGL8erJdKxF3xA9qTlw60fTceaCd
Jj16fexVZG44kGWFtEPCadm2f14X3gl9RIhc18+iKcRvRMtj33B+W/h/WJwY+xvX
gKMr5gWOIMj2T7ZEmv/N9IxLAnI+s9nxcRDlXJuVp4002JfavDqTSw1MoPxwztv/
8WuR9EwKWCgCZtqVNMxgUB9/WlBa0ZiBtGCxiSrqd7ejS/qae4PuM32aDo+14qsv
2hIEw8mHbQz2fbJSafYwCttdnyPsacUlghmSXHRZJ9i/BR6dWtmWNh8adTIudLIM
wUZgDZNbVjTcd81JF6Ftw6X9S8d+Dd2SBFbj/EGjq9LuvdeFwGc/Akl0fnWjiHaZ
sn862eOPVscqq36+ADu+Wsir+xlljZh7tNX4FsJVLMwTSor9KeHmOUFn1ydB0ta+
6j6jwMSqifmjD6iWpFAF/iC47G5bV0BQ6/hW3YTiz5C3u8PUH90jYIp2cRXT8bxf
I5qt5OIWArBCz88JCHlupGxjdnV7IL3bG81lvAArbr6liykSDqdF/OUv/OLsGVx7
kbM6SeutSMMsyNEODLluPlOPkVWfYbNgnPswtmg6xUBzZNZxZrA0AaKjDdjeT7hH
OXRRmIHFwJauem8JzEMBQBxH0Rbwl1b1dzcYq/0BeKTsRDcUwGhIMWYPLX/ZFgd4
ndX3W17JuWOkLW05przuxIJW7rlgyzcgP2ohAZ82ssITjSR/n7UV3a5tj1ALPV7k
98s1XN9OxaYBxlICyTJ90IoqUnPrkKrQi35tO7kNtWhUTsv6NlYzqYsfq9Srujt0
NVTI4wj+8X33hrkJ1FhB2IsG8WoAiKnFI0oWBMnjY8oPgVD+fD0mb5SZIALaacnJ
Rd/yhqZnasOuKVn1d6KihDv9rkuLUbbpmgGvMwoW6Y0yJ+wNKlfUjjTUgCfDWFaR
FaKxJbdHTdsVRNKU/5LFSHY4YzowCVaBCTGPgyI32Daf/tcUFkqYCSrW/2ZF/dwu
zdCeE+EIa4uFXcpg0dVzX0a/4p8ibpjsHEJ2AaPKOCtPGaSnEYL8TfkWL14rtaUr
7qm6lwwILvMFNCJ+xivkr7ZK+7e5DHnNmyYE5KMasSs//98iP8t8X+qaNocjGhJD
KLf6SzTfwdoKSiB+sr4bpaUNAzVeKlkfkAroMiBJg8yYC2AKeNAqPMFea33LNCo9
3H0F6TnEe9ix4O9VneLXBHfDmmIOF2VjPNrmgIp+g7A0Q73tlETT5IrPzBlk7mdK
Y4nEqWpx1PY06waf9BMpzcnB0/Zq2NNEBMNF1J3iiotMj7ZXA5qcusCVz+YlEKQv
Qp5y2wBZPmrul+AdSl15qEfavHv72yQ+xVB64i6tJm9qzWkIORuIixVz3nyAVuX+
AB3y1tP68hKuPZXspE0+2Ii0cbYJ+4DhXI9fxVyGi16A5+awoZWPJH5VY9/PiU5m
UUJHD7cUMVzGxFFI/S/uS2Eb0H490o3E1ki1A4uttJzAy1py+TVExXjYAm4/5vkX
aFTR8lQ1E6UY9Xw6UoFuH29ewV9pUyrxcFh57rPVcUfALFGQvpa3tfXAY8hFbmcu
c27ci13KL6+99O3fS01wnrP8QXM9hUHGXg+1MUQ9mJYTy2igIkpKiOU2l/2ExE/U
xPjo5zPYYJPYsRlHruLxrVQojmZMQBQKHi+nn37cmPXGuD+xY8mG15FbTWqdTYoW
4YWSdCRxqrX+91MarlsfGg9crAeR9zry+hdY15L1XJb9RKwyH1KTU6L+yV1eGrVv
GpSd5cEPKqizcB3sngkmytrOqw2xb67PwlVSa7RLDRIcN5ASPW2hS/a3AGpyglj4
fgXZbK53klCM7tfqJaakvUKdY9BvY3x9/bmm79v0S/eThPDl1tAbTWSfUN1pHpn/
S74TPiOvzj4xdrS2UresM0zjXsN0o3FwbCsD3d0b4Hp5wXiDNKUN+s0CfuPndXFX
/mgnyIC4YML30VMCf+AGpd2cr2dv0+rJMON6HoFkipUBr3UKCdUlbO6j66LBXqvG
pFjP6xIIxmfnK8kqTQBgpQGCkacMcKRDbgQr8dfJc1muDvxUE9p7pZ6yaZ421G2b
SPh/R7IeEjqIXEIMr6T+VpyUR0M6udYjr3tnfVRgBeAPUC/19NFMEhyoshbOAviA
vmXqEY3uXd/dqWIJzdlon0Al7db6Kh6Myw60KD1E9OVWbddy31KpvnMrrjH3Dmhb
ZpnJElai4dQtVYeypYfP/SaivuERlolalVtoF+e+rGw1STTrPzIcyW2xP4X+9ZPM
p1AY8He+y3Sau4eVmoVs0UVB4QqlPt6auRCMrdMAiL7AFS7xtjo0oI/ZjMZAH2qo
3sF1ZYNihM+LTg6gFPKRl+f5fT8VWOngltOxfvvHjvQlJR1o5Z2PJAcWI22hvJEE
M9o9ju2X1QvT7tWT+kBG0LK1lrcCh/tTegJ2O4ET1RRq+EhU9HHIBkv1qlpC5959
gxocBIYGkbueB+tC1XS2Hx5TWUGsAwjyxN52eD7NKlHRhraMe9X9zApkE5c0gGa3
7jpvv3LcwbiQw5ZG1oPqclIyz3BSjfjH1FnfpkPnec2ssOp4wXGEKhSwA2ZUuzxn
Y+B5cz5LYCxpGycdK1JxCWooZGmZYdNFXUv4cViFzIwuftz996fcQsFIqsFev/n/
dnhRfk+j/I0j1nSA2I75cI00bWKegZga5m3pbD5apjpLcWcHWAtvVnWF7h97CAJ6
xOHxvrRe2iEzDblY2/1s9C/dLEa/Lj6RKR5GZTM6sCOQZlLsurJq/yIel3YTy2Gr
CqBykTtDcstWn9ojJQ17gxn/KNWXjeY/28eZzNcBmLxPEOW4nw99k0+sy8hphsaa
JFKl5irL0RxvRlY513NIO2dn3wfY/mYVhWOHCk3kLcqyywQFlnx4ij2OptQYy0Tb
dpbL6j3Qsrms6W98XscLX1+HrAQpvDbVzuO9rLRXY9CBxzLpNZQS1ER63APKdYKy
1ti366TSBmhrC63J9wBORcVbhQVgSsw5rZV0tbO/wG3sg91QLHPO7slD1x0bvfWH
LJaoAauGaSH9pl1C+OXRDWp9iJimN7L22bBhndziF/zbteweWrLnqaZoWuKgKCum
vQJL+ta/eIQXLOhQ5Z80Zg4Vo7BS9yS8Is3fd+3IRr6R5cTf07ya4AQ6fpgOmez1
Mut305IiS8KCgJRtdwAfe4Mt8H77wDIBzJa4P/tkEqIea4073uo3L5euiCo8uIxw
4gQPTHMKFm/MITUpc8f6JazKKcDDf0JS/2hnz43uY+PGiaE2cjKd46Rv/y80A+bE
nsPo6UNkeL6fQe9+DJQQwyBsZs7OsP8g7IPOAZw/LfhFfkoPU/qsUFMhfynz0ZYO
5+PiPu6gHrtG3RZvYlQkmOnzK07nS7se5PMmp/g/VwJaNUb+y70nQ7ODnPUqT0gf
9RgJFFkOhiL1/TG5SA10KsKTmlJEM5pgy+Ume8cnPDwZwZoyBo4HNPz2jyrd/SST
iQwLE9S9JRDnaBqePXChb/xlPaTRgxnzrbw9hxlS5P6K9Elb5gQZBEbaJOsE9SQb
HtdDUigidFaigeCd4+lFkspAORwa/yd3WwW2nIr4dKhmSjNB3G/hUbzfj4S/eh04
MJbUb5+e6+b/BewCpjtmTwu9FoF+cIxGldqqo63S3pxxPXdLEnQzIKOCVx9oXjEH
RArHZCEosvRb7wlaXZk4R5jgb9epXwA5i+6u7AMg8gMHRn5zys7NnbxVn3xJz0eD
nnCayswmcYgv14FkfldvGL7Fo2gMayBb7QoB0R1BQsauZuu86i45p/68Ebshjus5
7r7ptas4rA71aFA5bvDw3hGjlJuLxyN0CyEq19J3QLyI5zcOoJxtAh0DjUUkpy91
chOQJsmrhAdRQqv7We9E+z9VYtDKFU6Zf3QIngQ3PHpFCudJzgGlrLtqRwo97YxS
TPhTE4cmYSn6oqIYnjcpRyh2dy/aZj20dOHfL+jJ7wCzMJpLJ86JDuEsLDVPfKAE
M0/qt3vqbs59qfQg1cJHTbw9HF4i41uJVyWE1lrZnGDgveHmxIFfDzpWVgrAupUI
Vey08yE3AoawZ71n1xotpVNEaR6plYUwpaw0pWHevGOzs3rP38Rjxo8eRe5vpWMu
Ok/wPIWyuFpr44IEOJj0iUp4jpgJ8Kr+5ZHk430o8UgLzFXbVQ5XJsVQj/yYXnqb
26eVCPKWwSGhxc86Bdrx6M3A6lZoF7vBXXmtdGtOzSph9KXPUE2xjmEfyd620S4H
96wqUbCH/OF6hwm8U8fURw8MlcJfgfJEqxq484GY2mequAVxghIlBiDI4Q53HbwP
g4IMzlD4dXBqPDwRk1Mb6iszOBxTxGJm7X00+YacKOx39RHrzNWzeNEroQcQYvQZ
mrnhOmCcJf6c7XddCy2u8oLZudtGitOb6teYtnLYB4oeHnu3fe3hbGGgsV+NhOLp
/BEnW3t19n2pMpOc4yxnfw+V/tD2awZL9qvzJJu/Dy6/PrakTEIDC33AljwABY1/
CeHWlnNlu7acfEOMRNqzQYGi5pgGvx/jtD8EZBK0fV2ocCAvYRQpATH5is7GsJBn
7hHPHpFC61UZuhuQ64gO1/SGcQOtXiLdjWoRwV5WdjAqowZep+QKBK/sxmcQOWye
9PzuImYGdGAKXACH35ViU5HjXJzqIctMWJ4cI9RlJVkKalk0inSaI7Fp3PwLBaCh
ww1l8tXLeuPA4PwJWUgScXO/uQ4o86wrB/dPWaJSQ/S8iesLrV6qOSt3JSsVsnhV
O0c07IGFxEANJ3CZlIieR1lRAzmTP3BrLqaPnLRLn9odZGvAHM0XB/pzQnD0EMmM
Fv5xJloBLoyJMOLS6V8sCq6EsV/sD7NIOE3Dx54JHXne9CFdBg8yLz4DFJWpRf8y
k1mB2MHCXWi5m99N3ckUIiPKT1f5CZK4+RgZpHE4JqF299DphKz4vB0iuXDPl9zg
PVh6PHEKkPz2K524UEGnkB6vNwkvO6U6Z9TlfMS2k6lL2kxza9IT2MrcrbYRmcVq
WlkeIBQI4fxHG0B+nJ3qEicTL2sFy5R8PcCJNv/wTV/ifr0TgtyU3DImDoKZZB8r
29cjGMpV+9PL18IwqSiPWyCcZS91HVd2HBA4AUyOV1Un1XCSA6/c/YGmCBn/NtXV
1K5PrJi7+rslOWHkTL23AYcTn4M9/Lzl43uUvd4nuyGo2+DnZB15b46rS7hSXNZP
TVJwA428MrssewIMfAUTxaPmjzh23GzwBMlOnv/G3tAVJJseR+VbnPFBdTZE0cB1
tzkTmAo3v2VO69sOdZXzT7bqkbVmLrsCkXukOrdWL2wa+6Cy1gdEveomDns4iz59
guvJpBs0FztCvC6Sjx99P4uwC/bQVKqiqwMsCzenXdSW+b7IH2jx/yKTawmaiyIX
xi/Pauf2SQXmxk7GZNyvXGB+ZPLGq8d/Uma8oAqKduDqlugOwDteYOMU+2Kg40Kt
DDpBLvmWZfEIHQia8b3ynrlSk/OIVeTdOOMMYsh9lhlwVTMXPBHAmDnnEubfW4sr
YyAPGVIcxss4fohic4vRVYbTuJ/odkhj0QEyF9W/KmzJHB4hfiwmAEuVU+uwEa38
lZPTrbR6G26sfnI1O91DSjUpOmlKdJQn0JB8SFKcG4HUpfS/PJJW710f4IMmyTIH
dlMNOCggrxj0h3mZpSUbwA4i7fflhnEe3wueDFwCekvpkHlOwPyKSnYY2z9YRC/v
nBxpt4MWPjLXMEY2d2SAEeERrQWaAdPCg9chL45xmCaev6E5NGnO+5cLGjBGV/fW
FzMcxZDpSik1BAsEx24GmEExwqo0j4cY9vxlnVBn0OXc2qZWgN4Hvj2g0uxxxVxa
GRoe86N8oN4Gxtr5B3HKq6s0CGo6wyUrlp/HhiM2dkBt+QuF9nPeDzHo6IDw0GaR
DUepQr3SOz4/ALPzg9u7zlRmFJfebNG6q+sFNsKFjuOsq2KvHweL2GbQZY7w5fKJ
IOf/nyCsm+BqbcDd7d/gySpsbI4l4Rr5ZoBM/sast4LQEuwByZ1nvwVasjhX+qYV
T0+cqK7xEGqO8cWWlcv/e0sEr7YnYtaSQ8g6XGpQtyv/PdP5PiR6HXjb+IEoZjhg
j/qOfdxx01Dt0Ul9kixQ/ca6uig1YrXcnj/GbAvoSmTWGcUseMDrJczUwAqgExd3
OnhtbPyleZaC8GvL0av844iG/CMnmlPfELwByMbGQIKCNlgYc3PFBU4A/ks6yr3x
iZ6gqbRp14dyTlIzjAorXzrWbbexoB6rL2dfVVJToLMvUyXros3XzRF1MIwTshhW
Qn0CWl2C5nd4+6bLU0txl4SxjNTQm9+U7kI5vvhIgZF4R39WDX3P1S13TzpK+hHH
5gca2lOlG1dGKasgf+9MvpxtKbT/auCSEQvyMelYR8xFNmZDQ0wIwhnu294IJmwc
1hhwQ1lZFf3jIVTcdOHE0guRL0ZEZZXE/q3npkfSLrH0s8ty7iK2dLhLrcflC7GO
B2KIS2LGfeHV7gyJyGRDUsqTXtQxBa2pQFcosxst4iwrmRMoVcnWUpW+3qoPCEI7
NHuNAOLl1b3SWLGykzjV63wgWnoBTYpDALNt/J2RfwAucaokq0JcSd3BwjV/fsf5
P0aRevo36J/wkkZxO3RID6TYjsapH7SAuVSskH2PBprGRuhrk/K7QpL1VZXnbni2
jNtT5mhc6odh+TVIEc6bZzIrGNBCJTEJgjYoFwhIJMFBsKU8DiAuDonRd4EpUR/q
PKI4abfxVnn8PYreyXjeEGuiqcxLMFBXdHdspwfik6zVmrD6Xxz1xqGuWHm0mRB+
4yNaMbxLfWyDehrDNdftWXC6i2QweOugKH/Z4fkCQa0i3YA1xvRg7SQr+Gkrs46V
Z7ilGET83YnXvTHXAyKcL5Fd7rcd93rHnpTAhh2X4IpWvxmF3lJc05LpLwuX9win
yhfT6Px6NHE+cniY052L3pJ1JmdTcPxMXBAkwgBfPZYVP87eIj49e5QRazXEY8sA
KhDE9iPxdXO6X15aA1a7TL+3TevPzTLEahWwObk5JbxG6ISjGZDEPE7XNEIBzwhu
V1fx0u4UaNxhTankY/GcoVtmqJ8ccrKGDZhFE76HJZo+ugyq/q4cDRwfPqi+JCbL
tTA0ZreCG0Qi82ZTCdayEAooXjktw+oNv7BN4pJ7oOFz1umvfbQ2EebfihMHYA0H
ZGYuCGD/V1l2hbHR/ZtAcRM6MVbE5jV4/xZj4ZZvRlzeb6Y3qL0lKl7iJ0ZpYPK4
7/WUxigzBxXXEnyS66WEMUaKzEFLww2tmNtptUKKLeXu4oKdH7jtKulyfMMphH0k
m/3ZqpkEXRioYWpGcUqilZEAItlUQ6VapReEM19KRilBYJRBIjbnfClhPBNq3BjM
6pNP5oba4/Zg4QXR6llsO38oPA6e8mNRaeYDRowxuM4XsENkCEprE7POWFmu1ooG
34L2P/3rYjbPburWVV499cTe91uFbum+7IjDYPp51vWYrcjtFuKdZeU/kRnrqgpn
q/IsDMEG35QCcKV49TT04PsJrDCChrUukb2hzHRxcoyDn74YFpkNBc08DTga+t1Z
F2Kpt8Q+EhF9aWV+6i173k95RtMjA+Py3p4BDANszkN7Ou+AvQm6wS/Bfx0hgJup
T0q9FKUD9X7Kc/YHbd9kuBU2Ntc8/JkCTRpRbrGMoCgmZ1qdm7J3qj1Sz0Wi+90R
pXYJnxMy3X1nse1wXIj/mT6eRi3w3I41XbRxnW9/vwmC29Bem1mSN7NCaUOkWE+w
rptfB/Wb/+tGubhK7ljwcs59NsJWdowoJVM39SWfavcOcgQUwnM/ez/iruV1bOU5
9SsEwcuaoCjn9yYsrB//XDyPjowpBlVnVMSLrFy2ddQ0gN2WRcXddDoHdOj7YT76
PQDJnX7PI6flRT0ygDlbeC1QbsuuJnx4tHnM1RSetLLUdAJ4XbdMUg/lFWEZ0G6I
XMYPnXZAoZ2p1xHBa92HLg==
`protect END_PROTECTED
