`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LIrU+gGUyqy+LbMsX/R5IOmKdIkWMf/Vsm+BOATY+JhgnXMvGqPRV1313UKXPV8Y
KPhkTRuic5nytaEqbxhsRbzkUGC97GomMba4Rm2dXSQ5ZdABaol+AWVpIJTUf5YC
2/LXF1A7VtFh+Nl9Dwg972oThb7RFOdK6u/Y+I+btUR69iHuwXgDVW9meobeamvt
Gaw0r2VJB/KzmyWDkaBa3itDub2nf/Fkjhd8dFaKeFg6jWrAeNaCQpDWQtI8b6UY
Y56BV016RF5hDUoKaRdXjGAawoDU6xRMDho5uZsg8OtUD3EBwcJPDLmqDGwCWtjJ
YBVU9LfurfhBxKQLRPI3jVWTFHz3sc8c5Hwc4vrdSgUruI8WoGe3qyw15VKZhJZ3
0sgdAgvb1b8UF/m8GdW0ac+dLjvRPrEq+8f1ja4cWoARWNAEMbGhQUEkQ8XZp8bt
1fgs9v2NXVV2kp7OqfN77jUdb60Jflp0asf0J9lKKGTDScIsanz2B/czuCnfLfQg
KHEWt5Y+X6Pdpt1z1A3uRBEujvT9s9P8LZlcZWw2FJxQMM2fYT7p/q/alSc8LyZS
InPdqCJRTn6gdU0wHLTP8U1KDJEJoEEHDi/nMcxC7RR15cR705w4xh4iaOGw3NTz
Ip+6k8LCjqFo7LqV/mrqWg==
`protect END_PROTECTED
