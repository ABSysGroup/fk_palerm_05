`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rsa+mkXDCpBCgJbd76mIMKlmi1FjEfvTzEK+/EdE8AydKP+KYI6WDtqgURbr0vPu
olZIFiHWpMINl9aHaGeLN5N+PkMd2UviI4DaL+P0ZABgF6sUDfImghHE5U7hDOgW
jww4VE5yeRV6CcRuT1tLRlXtchsQC1r0vMPc7DQldQQ/I3mm8Ck9E8vY/iOrLIxf
BP1kNkgA7FEeTO86B5yJ+PrTXBye1B7carhxr7/Mzu7IToQJK4mlq8ZKzOMSCSHO
E8R8OOxBwnkJr+ppLm7AgKNIjnNq69h9r9DFT5UXiH6z7OJ7cAHMMh+ij0ff5L+7
NfE5QRKJCucqA/S12UzQfg==
`protect END_PROTECTED
