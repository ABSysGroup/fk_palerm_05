`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tF7rxW8byx7CXCilw9sZDmOd9oKQg4NJ/t8r2gAFTF3F7dhoDEqZkFBtdvfMNZBJ
95gzFkZtXGZkU7utLcFyKxKUJwsCCq/2XhQE/8aqQXEZ2erccXT1sLbV18tcuUe+
fV+YxHjZvRsEb1Ls0WCHdzdZlolcLkAt+cgmMYTl6PBTB22+l9TGi96UAQqeo5LY
iOKu4BjJJn2Em+y4J1xyF+1OutSE7WpfT1S3KNL4Dxsj/GByMD6qVJdIoCV3jzgP
g8SpsVt8kxGP45DRX0FGqkUwxJLsboEsvTN6TyXpO/yZIqzedfceRh8ZuvPeLtE8
tgEyKoS/LWK7TG5zKs+CKBdnaN2f6tQ4SLdoB2NdGPkLXpslUaRkQ4TXev70KOdc
6kv6ARCpmBYjfb51SdIABqSoLHUZTt78AoYrQUjghtjqfk1+HLsRY5yAKoLhN42B
fxEBS0quGFinUlRqgAjeBMUU1/TenRHXdsCuUp0MT8XmUqefWzTyBkaEX/JonmBX
7ScrOQaza2ei57+k4NTC3Wv38KRxt9yH/kZfU0AMw7r6yt6ggA0vKKewlItEEZTU
RWxA8sJoLoXRM/F3V+JzopCQhfRzvpEz/97+5+Reg5+BrL8x5B6hhBTbS7QESr33
hulgmK/+VnrZ/ImYx+nEKmYTJ9sBhZuuV5/7VUd++EOoi2yx/yCEAFG4M0w2fC8P
xsr6b7T/lnBFj4EtscrZkBX++Ub9Vn4GZZm9XY504SjB8cB6E9dsx+b8Acklv/Xl
1ISMJkMwfCnr8+WDlQAoElAjtRlofeW66+curtBXK/mxqWEk1c5IaRbyoe5M3x1e
pnRxHOGBdpWrWmJPPgjDJbQU5iv5hAwvnb27SmqCG8yH8OTDl99mHkPE/1/zMZBI
UwJkLgErdQSVtxUOOPX13IeK4hPWm+307m5ONKw/H1c=
`protect END_PROTECTED
