`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9b8BMuEc5yTRcjO/fNMiAnTxVYPnQk26mi9+B8P2SUf163sDPlBglNzwvPhjZJF5
hFEH4d6mEJdlYfW4tmHKhLfyk2zzKYYADiveLe9GU0M607W8DeK2P762SDX9xBJU
jmPf7rqYDEevotbkufllGprUFmXEjMv9HVHGRNZmU2Y+ExKtmG0WNNNleeShOMxI
yHYnGkOKvNjflRY/LPbqyhLz388w1+14TLmSAtzoe8ia68zfh17FyvC5EdT97hPB
dIwfXtppluw5j1mAUXkr2ari7klw+e1opIN5zKDjYpC79yxkh7k/1o641i44/USk
fWB2784O9yPjGtLqSIdqERFtt/9JnLBhBgwsM00z8IunnigwZyVFZvWuqxiwVnGq
oOQeVOTqXXKN8pxXUdoXGJYjZPbkl8cwzLH8xVQeoRZodsKGumYpPTAJq/mmcUXz
BHnCFLM/aD0/3+4zB4ZlxLeUhrYd7qlHRwExYGe7fyYjXvto0J7bKtEm9cHWmWtY
CbD8r4sgWMUwtKsrIZnhU6vgOO2uVtRFs8CjClletALDADVvBLyjDQpI0MkvuFI/
6430kMehZRwVhmI9zFmQ6tB06O5LCzd9f0XxrNcsizPO2Yv9OaS/yo7Za8ZDkDDl
+2ynrK4KDvvvvhvJSCgaR4vbhDBICbc/8wS7fPHz8F889tujtoxuoFphxT+vpraI
h06fj8yXrFumHroCmSddLIbLuKppL8L9IIQGkqu/qCd1zyXHq39oMXOcRsRw2JKT
/5jYZ6e3J2FF89uokIfA6MPGB8NbgfvfFrKcv0k5Lp+5TLrRnxs0nCpoMjH4rUmd
YxSQ17iza3x3U17iXjvmAPP4zbsDAyXL1UQthZyilN1z5FtR+dlsC8oW7CqNTs2a
jM28xkDfcOZQ8LMBCfF8bSwS+ELoLhXsUVr/QLKpO5Mm8d0y/zevkBhRaSYovxuM
Q2oYtMo7iNDZaz07X0zm0RiH2fn9gfj2BLlBAKCEAcuTesfNdWyBQUnZp14h64Ho
b4r9yjrkX34JqEv2dr46oM8XnT4KNtharLd/cQmn6A5X1RLTQqfTiTfQxgFnNw62
3J2FZCkvn2xEPMIQaJmhr9ncmryr5zV+NEIM8VbASYpF+6DnvYMyOXO8t1OTEqEV
/UjPgPP9zvDdTDsyPqyYhPTD0KFdSaSQESZTpmit1msL5C1rRhd4tRBnCCBxIdsD
oFYsoDey5EBkDuDFsYDGcapf6Gi3aVuYt6BIUQ8Vh0WXC8MBNFQ9YxNBhbOg29PC
z53n40Es4Rz0FwpIEuejkOvXWqRROG+QqbD/I3JwRGO66r1Ry5R/kyIeGb3OdWo2
ZB59jY0vIm10l490NwXvjjjG4Xi8Uh61EmnFluWhFeDOFDNXxOmO7AalO39qXRLM
kOo8dgbNVV+I3wB3JIi4a7r0VvqYF5Z9cliq5DBFu5b7UP2WiZ6MeOJJUOQujD7s
AwsI/20HIMmUhE1CAzIn4yybx894j5z8CfZyhqVAQs9ua3o9RPbrCIp2Ro8oqLtd
IBNUR/UTE9/RKJX/iS5kPIsxBcmVXJ6I48JmhZwWmihIjbvQ8yzXGQSFMrMklSjH
/n+MU2GJabxeBeCa+npvWxH7qD1vcdZlyCJTzG5crEKfWvqMBbE966LDwxkQBSAT
T7y/34arnz1dFEb96WBFy3hL+ZX8BjakLNPSh+vRRwG/PlzNk7GxKpyO40VPv5oe
mTNctaHFz2E7wxg922v+OZNijI0xtmt0U4mdFagKkichzWYXj/3qLGbuB6zoj678
2i9avhTaT919cokiFWu8AysvRFVGXFb3GZVdtN4EB/yqTCkZ5WDrEL++EQQyb0xw
WCBMzUPKUOe0JbLg/vrE9Y0NPJwS/QQnKJq133exmldbVsFY+g5/z2TThAirertS
SGCB7v7cFiFT3kjop51lsh5UPGx3DadpW8aT4zms93QMJS+jMIBlDbo1LjEgpyHL
0AnsWYmY64xBwl7OtO8m2DRsDdktaxvnvVTacTSRVBFBCI/pNZ1xzLwEOnX2dyZI
OTRVBCDfQM7bFBimUeVYU28HnCAhkiOhEbSsDWzfbbwX8F3V+dFo16RSbowu18+I
ajeEpn61iyKdiFmrunopC+Rk2JNuF3AQTfkTWB4mRD+0fEfWmYHWuggnIrDFgKUc
IB/owBw2BLsTJUA5PX/YX8DKn8UCxTmiC7wZq2wAS/Mt5EYLp0A8mr0cEpijBl72
ORcAtrBjOu2EgB6jQRjgQQMRdskOC7aapIGwDoNntMh3WY2IX4ayZ3RrBQUQfEzz
NOvTonuG/E7z+shIAryPaW6BtTp7UWmOlx963I8dxXJtU/g7lPsr5ABa1gxJwBiH
Q8oV/F3uFwOWvf1VeQxi1pePrThI5d/V0t20qvzxOEn3Wx62U5Bca1THtq7wEesv
VqYW0zT//j1BfX0ruwInNV9042itmqn4EzP+TwBcv82k6cF86yuZzYMDy1IXWWPL
mC/bZ8rxSbXNguOUlzTNLJ1CtyrUtxLnX0Q1mw/wcPzFx8b/Gkvoz1IPW6V9OrIV
FmE721gciLXs0q/g3aRqJNvvB3gqdJyLEWx+2PgXmuE//fPWipxiYs4EhMgI09x3
fMOGSemAQXgCq6XO5558PVIOTEUcs3gFYjs8otKno3dcEs4F9MHlxVPq9GOcj4+8
u5T9e8ZQpLFR2cXXGsc8zLAfvKAb8iUDsAjpM2L8pBvgv3XEUjA0bjFhjgs6CY/Q
BgZFHxSW0WoyE+GetrxPQmX1JVQ1U7xBAyNKc4Y+eEa/zDMdU90oPa2UyWb0Mqgm
iKTgKxEtQ/qhauriyGG8Hr1jfirObXrebXzZbRKotag=
`protect END_PROTECTED
