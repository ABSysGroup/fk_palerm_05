`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MC7p3sl8QeH3svVDPeOLRxiMssf+HzUQP8TZsyGHNbDHEubEwG7hupMb3M44lPQX
QhSLX2a0jpQCtgMRmitdrfZyZjt7b72fbuSwe/9pzWdfVAcCnUh0JDLPp5VI3b6d
9erbJyl/i9DsSdo7go3/orE/8Lbnm7drKcMo3WTV62GyQNwFGObPRKCffRnwVZN/
pyknmGw3C+rRCN/MC8/2iFKCTGUQdIam2fDeEXznlKpCufA3ESfOw5DFPWN21baU
g0ePpabhgEQTyru+iJR7XdkETiddIBP8YFZP35X6rkTsxr5BMRdVYeDVdGWUt8xY
SzEcdwTHRkGQrrVueUnJPg==
`protect END_PROTECTED
