`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WNkVBvgpmoXIqqEqPIbqmY/CLIyABkmpGSb4ApfZJuTyCc55sJ3l1jnL9F/4DOZb
5LHUQl2CWMR/uxOty6c9+1i08gZgJBYf/9qnZn4ONTePcabsHewmC5F1VrZ9yFSE
O/N4TfMnvRQCdOK1p7tNlEduzRLmvdqtPdsfgErlKDdAJf6D27vMrVVzc7vCr1sQ
Z78rC9YL6wvuHaxmCGzMtb/sZmq8endpKJKuajcZlZKYyX83XF1evhuFX3JV8mUq
7UdsFXs0EosQhQYsoJHdPOiAyIbMtWmEwNUlfbl55M36WdFmIN23lGRnsYHGjgvo
RGBmo7b1KAruEdnOAtAszCe8KpTFJ3U97cKCaYCIiEK50J5Zll4WBNTa2NmTRBOI
aU0eMrh6bG0NjmqOwEFQTid5LZnK5CtkfpghfCB21RjB/hFXlbaOUB4074s8EQt2
WrBEXOnYSg+9rk68uUaWfty940lQOi1BE/Hjfh0x4HEdNEzv1KurR2YNuUUtBPsj
LVcU6VOughznE/WvuJ64gD2/thzSZZ31O5/j3JemNhAswgdKqidafa5ufWudJVs+
dgYmv7/DOmCDA63e5Mgl5hvJjlpaL7CMv/xA3GT9Skjpa/DAZUM3wYUV0QdhOwiR
QfKR7WQThgZ+QWqvzKYN2Q==
`protect END_PROTECTED
