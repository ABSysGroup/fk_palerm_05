`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pWfDX49uxN24B1KRiN2giZXK1YNEoiFg5faptOmGugW0dcNiWfkYord6snEAeHWn
DFRX7qS3f59F2J6HGfiTQ/YSYxfEuDsa+hYf0HzSaL8qimeLAgeZ1IecO5M2aHYQ
bMW6rjRdxa468kIyINV33SLnF/nihlq58PNUviBODG4cvffWx9E/hvxFPbdIeuQT
2uG9GHZQOYkzXXr7jVM4jCBV0tKuCuT6r1CV586HpuAG1bkEVBXj/3uMe7ruo6fe
/7tOl73leMCesM9rqXRFcCWhMgzKsMiLYaSqDT4tog8aSITq53nuE9cOQKVpWUOa
EU8Tz9j5BY14E/1gs4c5MJKUDzoGWtxbjn14cq0s46ElQq61t5KspsWGM3seQsLr
32knGLR8U/L/kVizS7uFPvEKwkGsgH3tG5BPkWyswmB1ls4oGvbQj5iemrJyZ/qN
lETrC/qZsvwCxj0FSZB7q3OuPy9MGjf7fVoTf79KP6+OUZNI5hnNpR+ObiqxAp7a
RIFN2lz/ZVvBGIYPtWxEn692fSayU0PPQ3uLLRZv3CGq+YNPVO9eA0lhpeVSygHu
Dp9pCjproFxiINJ1fLDiKc9xfkqWWSIIo6uLsUC6S0ghCiFyw6l+WPpH9lb0Dje3
b+fbh/lbWcuZYiBDVVXxL9RZiIxX8UwDU55iTgAKQ3PxSqBgXY2RpTwqHWMWQTUK
`protect END_PROTECTED
