`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5R2uOT7alyHUQqHiYi0Ch9HdOkfebvIMW1492FEKsD4qt/3f/fAYNiizSNGKDYfs
6JiY6rQW6WhoMlEh8WaQu3CuJAzqAUOVWbHC5Ig4aIH7kNDiFzEUfKTXLpuFyQC6
uu7UaHtlqv2hdhu1H33NaGWa++jbX135v8Bm4Eyn6KGLBO35wcGEJoFYxEHPHD9n
qguHIcaoBv6QDgp5+ZW/OdyH+H0QOPfPhYKoD3pjGCi7GvDqK1hKKHMC9On1BuY8
4FyzjLYWfujkjPdqVbvpe7vQ604ErPTBD4AaU4vkSB7jTmu0d4F4U93A1tj8YpIw
dsJwD1+Wawiyzs3Ko6Y0Cgvw4BAtiqpItdwC7fFoJwuQ7M7QmdYwA8m2sj5HXwnm
`protect END_PROTECTED
