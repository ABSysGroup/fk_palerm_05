`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vNQIZWatBSA+3oVFyKRrBxHBhPRr3sXcyn/6Fpd9liZuSgvCo19SoeH5mQoIpWfk
l8OBmJQgMQ03ogIYsL9Gmv7fbiXSmqUXiv+y9Xk9zK714ZSKr/ZgNb6S2p7x/OQa
HGt+9sa6WCQT254rDl9860rtc+O/MNt/SAs4/6NLkIxK0KtUWBn4/DReHpv6rnHA
DBKh9SqF8+mGotypfhEyrF28LsRcIklMHU4D81dIjRb6Hd+2B9Ys9bELuXK1sLy/
tT8IWeQwk41b/YGjr6BdEUXt4fT+14T9vd3mUpRd6/OLUYdxfM4xkz2NG3U3Xi8q
OPiNAaluHvmaDm32NrtCZiCdJ4tFpC/zW3ny4EigFjN+o53RKBT3oG2giJNRWYbY
gRAYWHNIK8ybeUaP/uoS/mL/BP4wiqCfTxvxiLTZiNZ+g+36VsH6+OueYAy3Qyje
tnX52wnkTKA8c6hgRKRBMMO7aZbJOBIecq3k+YmYFsYlRBitIWY0/+aU7zCodqae
IuBsSZwrNDmhN5Y7QdJPWrdrz3ABZkILmVhcZT2/+Wg9Z/cv6lCTZXZqE2yIMQlG
GNDzcgy3x6X7SXqBWJ2HnAypd84QLRlip1BqGeC72h5lvr0MfDGnRHkabns6pSXs
ILAaCyFE4lnp8kln6U1PGHbxasBYkKK5mDOQqZv7KZ40lZSrwKUB5xtfZJO7J4lO
cJz7IEUOiCs9myOjRmmu5g/iUANXZpfw3XNWBUJScn4Q4CDfXpK76cuYjbk4vQOC
JMBc8uX5f/WzUx6vC0UBXOP7tGN7izyrhzBk/Vwb4DgQrjjSM3cJ1K0QFRvREGxD
oorgZNA1TxL2bITrXaIBe9/+m08NLXijX4Z1DpeGSvC+qQxpGr27mRNLnzFKXI8W
xHKNDP4Ekmpndjq9PvizgqCUNxCvfq7eLgjn1XxWX3cllzs4S6czGBAKd6w/Op4I
TjdnXvEaMTcWASAFNPg/7s1THk2zmToyugfREGrcQS3B2Ii6FwaBhRmP+ShMhVT6
UMHyZiOcWgp165h/WdoCBckJpCoOJOZ85x6FfS9aurPrzxxocUWzpDlJQ9NKjJTN
0Uv/waynR4AwaiMtSpfBp1hpmTszkwz6PjKHDs5LHiK1Zc5ww0ISKOBZMMl5HzAR
dDs9UyBKsOaLMBKgXhWGjiXa1D7mejC6OSSU3sOW8S/AVQHzYfz+9+iQVlAxBWTJ
9E+ThlUnnUx3cgg4WpqG0SyTYSPe59S3F/w+Rq12sSfnDPc3Yn0IJtfAVBIdphHs
jP2c1zj3+s8JZu0/k/oS1jyaHjqsbHWEZjxJCCqoc8/kl4mib1dQdPE/J3VvfvA0
VSnKgbRXBCpG+iTYHwSSsV/SJhyskJX5I/43K2qi+5BAz4WOR0UPsdnElx0FYiZj
mVW9O+7jHfeon1dj1Yccng==
`protect END_PROTECTED
