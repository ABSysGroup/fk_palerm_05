`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SQI4JcYlvDVku3FB2kyZAm7t2vHJcOvwHem2v333RTccP8StOHj4unkWrTUMUsxz
bcHeBzeR6eU2zqFln2aKmnOQec2CIMtLIZJVoRtgYrShzC7vQuvOlDI3b4TyiVVj
C3483pMml5JPTE0VNOQR6WQaAijALbbCYS1SyeBKe15hkyhRXkhPrJwc+gmTYeYG
BVEh2iLrRNEEbfwmI9o8TtD7J8AWsdfFAn6VB/wEBw29K172/xNLgJln7elemBjX
kh6sj36WAQ2e2uv31AgfFzaB1jIr5eKinG/1LDBdHIS2qbBebvFb20h0AQkXSGiP
HHDEhSAFTr8SiNzHitczcsGzWUwFiSnZwDk/Ukd9FFBrgFmozHabR8ZSDJp3zyC/
PUU1pW4hLCLiJ6HkHpSDp6DH5+zyhRYWmdl3/DDcJLYJ2oB6IHlMV4nMyoui2SJf
eZRONUJcY4pI7EGvFj3pZ9iUq7Trc50uIFgI91yARJ92QeDpRpX+i5QjTaql5jxf
LwO1ygKUvapvo4eh+FtqrP2iIV5JLP5BIhj42tFM0wUpKY2vVFj8t0t9RisoZ8qb
`protect END_PROTECTED
