`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S2YH0ByAJeLpzocZvFaSHFsoJPeIlG7vTXJT+sNf2m/pDgDqlhQfaD7Au++XJNde
J6mhUxR/E2bPAfhrV51JJUZtGqn2F9eCAyQGLHHa+PwWsU4kYzyYYs6D8Epd7CEL
0SRpNAhrurOry18xB3M/0YSqs+sFE9bH7ujp9dnI3DT8n7PqFfXhRzO7QUgBHfI1
whc7lWUfOK4QO8TsiotodccE4u2Wmu6Pf+LAk11x8f7K23qHAvIu1R0RqLpfvr6t
+r508YgjS0J7jxMJTUaE7asny7icKkbD62HaV4DKYAR+8BcLLjG1Cu2PRsSHuNow
VYU/4nDwZcAEBHvhGmrUoelViGxJ6Xr1rnqxo8cmUucQNf4pDpRwG/yutcyTIk+1
pLXUuFDgpcxEuKrzQc+gaizGF4PtqDhHnXfGjvyBTltjDAFT0vs7Hs3upNivu/5P
zYNo8lqJquEKiL0kKmw60yjmRBRgOj1sWRpC4oBxU1I18ZXU/6ID1ge7kR00hrXP
sJ2ocAgrHe8LRARHKo4c9qvoh+CvhhI2ExioNR9lpmjgIoL7mSM1gg2F7MJeH13Q
sRYuUmEdv/ZtJzN8pwX+YA==
`protect END_PROTECTED
