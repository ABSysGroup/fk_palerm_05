`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wj85IIXEWPtjGMVKwlLSUdfIBaIfuwPs0nnEui45eWiZreNVGJUcq2JmC1D4k/fJ
wN1gDOK0SbLNqaZeFms+nWFlvOv+pFBqc1qgDzSq+Ddd+2laOa/Ucc0A/zjIJVKX
GtGvoOh/qhXlIJxFxCTUqn6Ak5FlB+JV3VxkMGuSAFIUcbE8yQaqzEb+TqbA+ccL
0qKnxZGdR+SwzR81B52ZFsW4kWQ780m7kFzOL7VGAnl44VWj7abkbD5tCJzwk0uN
EVHxlYr7+zOUqWZkl2WV6LTl6Y2oNUl44Q7Yo8mwSElKX83uJ/ll8k71HL71RYqG
93pWoJ9Gp5FwH2FOqGbHvpSgf5II3y670kyzg2Hc75LPPdy+9fMz5Z+nuS0z4HIZ
CY3cmcpABK0f3OytoZ421D2MlCStum13MWqf9CX8sKKKxKkCXJNokQIFD2uH7WB8
xybHzw1pTQhTynm5XOPtHlx3DUlh3x/jXidYVvSVBfihY46UsQ5+HKHD3ynt2g/O
PTCouUIQipwDKPVC2iFrzSOXSetqMUp2gMN5WxQWcFV2gFY10BNCCUzq921OC0af
6/YoaxSTBQRLFSMNWtk27zuoYDque/b3QczEUcMLwQLAbg1OcDo35UcRbSFVzgIK
u0VuvqOBWtTeHHXgxM+8murVMlJFK47YGiy7EM1VgNDxMWllJ7EZtGnZ0EzgfD30
GpbAGGMkbwQ0eKGtxJGhabHPAQo/iJu94TSijPu8mabwboTE5SP4pRuxcXN05qGT
fDUZ1gCGQMPfcV1tn+nh0rhgFD+7IebcSkGOvA3whjC1zx/nGxXxvPWGNcRQQ8qm
C5Y4Au7qzr8Yzx7ryoI2uFs+G6IzH7rzW5a9E2IXnQGJd+z/sSZf5+s4fA2ombR5
fqfMLFE5cXEa+g/QVVqXdNGHSA7Ai95EupivqRhwMOyJLrdy7lpQM+KaC/nKi6QY
Bt/slYbqY1t4DowRgjbiZzdP3KorPTYcgrMN9WaV8zZVJiMtmeESaO6IjT9QWBWt
SaCAdo8YajKCe5g6ide1NyXk1y1CRpLR6b2yFD3xk2ykjZBpIgcdTLXMGQMI+b1M
GZNXWiQ//OPD/bfEP1paBl4kYeuoZyoh3UnEqTNx+Ay8JuwzMfTcTnJ9RPnI4nSy
vxxpIjqKOXRbiIKdVZHZSfaoeIQwBvScQpKS0WWTdu3R+6GR0X8De1MXGGQZRqfp
sxKTFAnkkrxWZxhInMFDX2Jx7dd7cYT0fR6EJCfvAANgvu03CsuCK5Ik+QXRt4tY
iswRPVljY6M/yRaGogxz46qpvCYL2FBGg0FtfDa/KM5MQdVmSW64i6bGx5GpBuGr
TENRMquCOYbFMMSY/y1bEuFVuMlYqc8Y8Ws1fv3E4w7nfyGN/D3p5NRyDLHBh04w
yawhx31j+7J+BCuAK821AFZoJ4XIaH68r8Z9WPEjioAQglOmHMgCuyLrM5NvxJi7
j5MW5NG4FLM27wvbryezCAViKjeZdTJlKFrHttIV89kzZU69Ehwj+rMjmeFp+VcV
RfKrxjzseUXtrud4pM7DwTmTg6srLMqn7AlTw9Lb2btVMaLR20+2lBRhV+9rkp+C
pFEHZyydNZHk+//UtPTOmcczb/9yLtT2mc+R8zkjIBLutbCrU4QQ2h7OI5eTSMI5
Rv0Q6JDnH+hzJIjJY/xgwrn3EW8ElzhptF+RhfhlFe5FsQSnp13V6tdpfdelZPkH
sRTrf+ItWlh2+b07C8+RWvEhgHIvTvgUJj3ZbgLrSOSRerJUeUC671eKgI0jCqxm
HF1qz8+zLDDShmHAOOgHS4p+/sjYrJqtKxE6EgNjv8scwjhI+ghpOAlWiHtvdcHR
m6BtlN9BoSdS+nJ0xy1+WMD+5TgZYmtvsYMjAFnYN3a+MHiISQdHV7GuOJ3U6GQ3
PKJl2WLEjB/8LtCVdcYYnf/Az1h93n9EWausArgQQu39fuk5fzSK5bzEv9tGed//
hpjfJtT8kDw6XEDF/ni7R7zfqn2GPO9MAA9goXMdjAA6r15xrdiAv5DvV848cKRV
d5/8lTPHuYOF1CQXjharSlDpxpXpTUN/+9OEyuAqL/Q88I7ywWc8yFilM66KY0e4
EWBqEXjuYhkqKR2nKHgX+2xHtqmx7doGv8A/6SG1WN2blESCq0LKJ3Ea4VMiZIzZ
F4nS/9+KABJ+GErhmc86QFBfDHRmw9/IjBCjsa4awbBrqvPjWyMSzm1nvQ3DlZ92
JB5gh+mT9padv81geWAMa+PUFUB5RINygB74k1thY5FGYGEQ1+w9kj8jsHCjj/vO
gixrcPtJ50eUxzUUvgpOo096Y+/QZOXBbDaVdm3bqRh/CoXaEXg3y9E4mCNSraAT
2U1BpvSuJ4itAHh8OWMzxrdfIbyDiIpvE8nRd5HYb5PcmFmGWKdpCPUtyB+EV2tO
H/Zdjb1lFvgWQQCDiySJw6rf74HG5nbREj9TUa9ERq9IMjx/f3rAIdoeYlqJSh3D
OnztgsCDaYK7ymxNG0GpgDQdu6K5E8x6BUtN6xju2zcZmIfIxLwv5PRRUN3/n4LZ
MXZbTtVgyzxQntuv5KfRR6fdF/PXUrcHyP+7jHlmpd3OcahLFx5Z0swxd7UYNIhk
oy8UAIcXSnbjNYsTyXlE4J9fJxD60bLG2TEL5BiW/vBqCL6nlzMcXj5mkJHewXi/
/2J2ksfeEoE05+8RgIwpTEDQ7UyMUXPMclZ3LMGzn/mNGr5NqyrwThratMc/6S8z
QrkW9a+q7hq2vB8oAMf4D7eIfjOGb4zjhNi/KAgpxor5KYrpYKmMzOCSqrtyqOOn
+85j+ddCVL3f3rqxpvGFPv3OcED7mY7IxtP9YbH6xC1AMHR1TqHaVq1+0no8KmUB
Rw0yEG2ClLRTrN+Q4/MijUv0hTwMceFzCvQNG5W6xcUvVjFzzvmnnsarcoacF7Cs
qwW8nS/hM8nkmOkx6mQPShWjNyrnSkLeV2fZ6qBybriy4ivn7rQgrCeMAVOoDeZk
uohXa7VlOOHWP9Ys195WdAY1OdFexyXkXBLrjE7ykm6D3IoLZUhh5YifjPDpzqSB
OKixzYXK8Z+MPHfsS8GGI+Rmzh7UZyVvRXsCiJY1MKlRcXNvJ7sOix7h3dIi/nrY
cHtECNqLs9X3bB3xaXneHxoHrkQTMq71Bw4o67Kluqt7orfiTvmIZdZvPPFmY2fy
ymB2jwZWz2Kp+sQ65U+ahlAcLdTjYqrindEAXhKjgSn2IF4eTR3aFftKVXNf1+8J
IdHzFlu5TGp3HMXKf//f6aWpiMWyCENds28ZrQAePRgL1jWvYC278TU7oxoD8vFV
1LsnB52dfgj+yi2JlUey5+ze3cTW4VK/iMWRaNW5VCOZ6P/1RSHMgOfZuN6zkg94
QLhPC8pBpbljBoRdHLVmA8E1TEV7dc9asBlu8rJMQ5oKYkM7ciqr6W1hWbY64/Er
VyNVDX0w9EtUKSJeVJO7GeDMxfDhRFGyVIfUV8albwJcvNrWfMJJAV0UtLWcC+d0
Li6jmncMtKNbKvoWU+Elv4NUqhAtJkpBeUhvg4mqZ/nywfAICobR618mccs4DZWU
nkCGMz/lcxvOGyXjQbblixvFtUi8vyZ03DzhhgSahpCq+GfzMRXRm1NldssuYylu
2PE2Z9TQZ6oK6atPluChb2r4rCPxE11SUNGX5ckqP0bAExLQ1Q1SM2vlvc8wvT81
r+Q99HbO+8/aR6wEC9TkBBrx9zwbO0yQSiir1JqY4JYe254mBSN/ckKLppC2mC70
3FYf8BiHOe2JhYCWX5OsOvIyULY8PLbK9lNQqowCDk0+LAKKQc3wTT2XnnkuxGiT
j1uY3yWN32gpnqtAT+LuuSXdqouC6pmA0fp7AeTttg+OwbFMUr3DBmGcr/lYDz6j
m+nc1+6zK1jNfXk/EcTqOrAR9oOgh+Ph4jcBMbYZU27SAREILKSIZNLVqwhxiNcb
sZg/Iy4/KT68iUulmYBeb/0QHTA+aKnL/m+svPNT+v3+6uMDMoapfR7ElLOcd36s
ZISxvOC2rVgLz1rJ5ppYrJ4/wNpw9fbVVEkTFhrmMWLIFFknwAyVacE1SlMdkaQB
8lc1/b5il2J0ez/fpHw6/whn9shLUALgATKM+93vEbWnJ0ocd/Tt1MVlsN//v08b
DwYNRCME6V2d+gLXgHAltDLqPQk9K1x34vx44wfrRmgeZsZQiGNj9i7zUc/tcyLD
pM8zZtqLZNefuUgcS7U9g/jkppKcJ2ZwuH5VeLEc27jRlPG/4plmUBUMn9YGeyhk
y9K8RhM/V9tFRWgcZp0eKgDxOggz4sF2Zkgt15cGJnWpH6CwFk4uFpuSg+v8GOUY
fM9ry/BDZGp+AYmgH5AaQXbpvkLA168dZW+dykszQCmNDVf+S4In1EQC06vEFC6S
eMAnC4ELJaIRjy1bd45iEoqw0YRXDnSJISVjkanjP3Kc9amLKSWk55QfrM/r8BwG
g9eqI9pudV7StXGMBzNVtcNlRJTFD6SlHmwjladpGtyHUv9skcwUZ5RWdKxHVEJU
fcJvKhdnrUq+Ij/ov/QrZG8TRTgNJdjIglXRaTzGO7DDiB0SlnIjWcyqwO7W81fa
tDctMco++HRqzBe3wme46g8iPmpTl/bnqzkN/b4RveSo4osuJhowq8yfRNFlhK+F
Ayk+YQaZmibI99p83GmMq5QeOf2H2X5dVzIlOalPUUAbqhplomX3+nogRDpLaVgR
81t0U+IDnTJZLnowyu0EyPH7iBqbjvx4I38Iua4pL0c1pwVysHjeuyfAr/j4cm8e
UsfTYIkMrShOd0h3B0T8OMCyAulyJndEqR1mFIYFu3/tXl/HtirrNit4QX49ZwuQ
h/qvVFmgx4MAfbJD6S5vTP5wSK1xpfagImRARLbg3o/nm5WzrzYEnm/XPb6DeQe2
p3xF3ZlTxJuPhlKrrvIMcZlylGR3+3RHUdPKpgD4J9jhK0pqbIpqu/Lt7/jDzp8C
y/A/mgopv1vVcH+HEUKQM6+BNQwIh2QZnE+fWrQ9eAFg64/pXavv48sz34JG2UNx
7H0jEk8Pjc5CVU8tD8Z7/CBH8DmUAx7a+lFWu6yDDeRrDNF8hEUP5nZWjrowq6jP
r8Uok4b5vuopoc964nBm4J4Ui6e+/gZTBnsvR54b42SKPu27ik8hI5IF3zdhfAdU
dH8Zw4nkw239+MgBXHwhW1FgGLjWqKlTeUxv5QEyM/Av3Lqi9kJdMkShXUzriyOp
9xSQLpgQ+IhRcCdC6dcgLShAXmT8/sYKMBMAJPnF1BIjeYUJoZC5dY+9GCOc8BeF
eKRxCm7QOxw97rV/C7B4q+01D2+8xS7aEghWAibSvtAXIq9FxZ0T8A0gFRpFAcDl
jbzjRoK3yYsmvRPfWGcgRIchbCme1JqZrlFSZEcMOWPeXRHWCNooNf/YUyBeHJOc
CMMrpMdE2et0EKjlJAyoRE5lMTOFITbJmFq+N8ybNgrlo34rFeiWGQP0SPEJ09nT
kVYdT7P5ksomhoT163GDEkIbCMEGM+4IfMRr00LnqPzlVCP/y+2QLDBoKqRpf0Av
NAAjAZnx6PdK5sfBBPmE7vSJGVLqC5lBdCt6R2IvmYeAEQU7SQ//HcuntEFX3HB8
OQA16BTrzfpPVcl8jBkVKw8+auCVL3cYV1+VMFI2Jftua0/bDMDZw+uqjY+h15Yx
O9usQgoOwoZKxvYm7ZBuLICEpzwdBYrlyTimxbTJAzpVm0Vzv77VGArL3XSyHvCC
ycIXzlI1A8u/lhaFiQOvnO7wMXNjji0xuKByAhUhCMN1dXj17p4LDnUaHpbm8qx6
/aKKX8J95W1h6xCxbRI8c1xcyTcsaVjNImaXXWkWylAvM828SL0q2Zo/qfj8ngIi
0GpT5HPqSsu59Q33eea5a2Q973Z92Z1LruYQ4R9hLuyBbq7pSLbi2JHcf2gl0OMj
EOHJc5V+rsm7iz2aanirVoLfuDmzllo9NPwsLWDaEuZyjEr/C80CyVk4IgDeBu/D
CeHlyg3+DIq2UwprF1Ewas2esXdOQiWBdyJFWYF6/G8hg1cAz8XBC8bJ4P5oOlOo
fq7kK2eAAY6QnotD6wz6Sl9vBO02yonI9zjCWFNQ8aKJiIBjfF7ULeh3CD7Q5f+K
OXJiXBzFIgFYG+02b18jIq/Xhjj8asJ0jwxwqfFZkPeG0nfkv2+bFAb5TNvY4Uoq
MOe7GdRr3QzfLZ0xl4gqV2NpvWB40KQ9526zJQJ+1l5VvE5U9IYUDcpoGgVWW6fb
F4cermvkajlrBAv07pO4UWqm4PhRMUqgFuNMoh6nKV0yF4E30emlWNONw3M7i0xl
BFbgUW84f8m03zAsu9kwRjtEyqFSCJGJzbhaItl0Mv0/hBePi0d/h5Z4yAL8LztP
23s0PfDZMHcLmPiNvikSlb9JPjf0+i1EgjrOTlNwGCyc7VVlIzn29nAe2L2CaKp+
IzCDlBFx1udj+6cvWxzA9YAwAVDiZBn6MW0WeZuevjWFaKM2ajuw7P6kf4O3KNb4
doK/krcwE0D2Cay9M7PLZnAxNfoNJAtas28gmQkSIm7uhkc+phWtU5YZHKJWhcPC
F5rDZytxrNFK9AIFHAjYadH0Y+kEtMjO2Uay1Q7aL3vp6KagePbM8Wxk50m1kt8X
MEnjSuaRc2bZgjWA2FXzQkXjTzz2IO0Isdivli5Wfw4nEyDiQPYdt3gN3xXSMyjb
J52uJh1hj888twsyxzhycVaq1n7YpcxXXImaYxYISFTh/W0Z4InTSbJ2OWC17zJj
vcADYOFyM+NjqcqnDvHdpOQ+COmUQbv3G14syMFZ5CFB/BRM3DZwshEqZE0y2IPd
P0dt8ecpchWmWAG0nc/H8OTB6AzK8kb22qlTsa1VO4E1nzyxmngVwAQDmkIo1QAa
f4tcWaPYz10NlEEEc7soTdexOVpgAK0jLKi+47jp5WYYu8Zb5bnNFsy/08HA6AbR
exBzvSEfW1yLY9+TEJNT+qJsx5XHJwG4C3aubx7LyjKFhVmJFEeaaG3mEeOmq0ms
I5lEJeio/JhVkhOefvx8aC6Essyctr0RwYp71f76iufzt9uj0F6tfH2pWPc0GpBE
AYJ07hH+iCF13pErD4PXeXOG/gejYJFMTUC3QbPSXCA54Kjp0JTyUGOAAqscziHj
5PFC6HCkN0d/yX33K2U01OVZwhpxME3iMlf03+pNgXXZN7GIg/+m8AGBanbo+QBh
Cr4SzVwr6MtlL836dY045YdiEnhzUoV9g8ItVPw93vTq4bUtjx9x1JLVdxzOOa5x
+27AU4p1leuXJhnWq7ViMGNSeq97CgaunqLf/WOMzOElND+5coC0OxPwwi7S1n0z
ecKxoCMyNmaj0ZkbyEex6vqw9nXs+oYpx6CI3dDW84fb9HupjXCf8CfqTJvJtH8h
ZKZgQ41r16LqYZQeThwAM7B7GkbMHpi59JnY8lwfy6NeXcjkMqpyphdfBerjDyYt
txmcts1fM4QIZxWWyRATJ0zPe1vYHPqHYTG8CugY+CzvjlwQ/2hpf/UHVHpX5Hho
EgQeIFiGU9A6qppE9+JmXnFG0b88AAeS5GlohZEuxwjBBTpFpRtH37xsBey77vNY
ZUdUUTZUmEyL0DNrFe9GPx0kK4Jx8Tjnmpxv6n6fOJg+aWAp6cwxKkaDJl675m/V
OLno4TqhK5FVbge9JVmlArAAyjr8FbYXMfAcTrI0ebH55or1do7Da/FGVbFPKmEh
hV0vb6vBJcxDZzeySvUsI62WbeaaYYTkPKlFRlTDRtMJlDc4wN7IPOj47Bomc8t1
JDCHVP53t5mymTkuMCtHf1XhO0NmYVYOFT59+Gg5RcAv5t1VLdpCzH7/hd1A9ib2
f+WGpz53OkMjLOHjlGA41rcyWSp84bwNWsm3uYn9fqy927KEFgu1W/LSlrtBaM4C
WMOMmwoJafsoS30IiKyAMhD1fvkwIICrSLMb//EXqAy2HqKRmhTXujjDZpO0Ug3D
YfrfspADDXgMXxTWWegwIJFxbhiRx9HyUcKBkO16/R094Nbi8H9nGtB4uq2ucoa8
qi1R33dWAk5WcTUARWikYTDhu2ujTGj0QHLeLLPkiv0xO8lsQqFvxRO9n0RbVXx5
neSEYQlVgr+EhijDYzxf3zdztTIeDnruZJLEYn1ty3oMmE/QtM1oZrDDRIypWxNF
4xIjHPp8YlV59AZJHLQ/ge5/WuR4w3/J05QnRUdLiMl0R/to3Yi09y6W92pvPc9Q
eVoNLXC5Kmok6u34l+pUg46QGQdlciXKGLiZLX0hwzN0RDEhgaAuZgw9aXR3PWdc
LUyOMprnKC46aZIRLE7PWAaNJLvfma6AHqPAOX83739maD2QHxLZnGh/c9GazGih
Dfevuhk7lgoFO5+FiX2wCJRhiUVpbeRaiZnXhNzgzsXHuU0GJ0qA9lyKdZDzmcsg
opheZSrq1EhYKhgteJi5rSmx3xWuw3B266Ov2RYBozjCHgAZZfkYqUMNxYMICVbi
GfY1SebhVIRTJ8vtUDcPUDdkhp+piExISVtUoRCT9/esMu6yt7rYNsLU5wUPoZqJ
qI712z2MNTSHiEnFZy1yX4iG4Bp9Ab9CNOOH+HFqg+4FmN2Wy9iqEP3o+iqj9iti
vjZZ5zb4Th8SQXXEgdap8MIz7yx1kTG1iWkhcQWUHEJNlpUo5bsU6GEQYVFgxUdF
sKkzmllowsfJ/B40S7WJhEqGTleOH5D5ivKG7E2Ak8z/80gIHEEpAgZ6kbA67/v5
vBvrn1cSMQNJIf4CrdGQxJqlRuhZ4cU1B/0zQNoenuCm4/jh/sHq0LNNXwQwgmHS
5EhUR1JNJ/on7XNYHzsDZE5l3AvgptTBgYPK6f2cTVj18OjSOd1I97KflN++KixS
rlTjhLVAb+DcQuJA0lLfi5p8s/zGMTn5bj46HKl6IEmaQdfctCniEJdSD05wDWpf
msArjQfAnAMj4HkFJTgpt2Ncm/X+sniKPoYQKRz5jCD17genLVAFKxV1al0Yl8is
bAoFwSA5dL8WO+Ccrg6QQYziZW5ulTaqJS4EIkEIxGsc4+Rn6MqcnMM+NbGloNjH
K8D4MoK591m3I+1/snmdh7X2y75Zi1EqFyd1r83jhnEqIzaJiowgSBYPqSBWQOAW
jhrSI2xQNjyUBZoBDp+IUnr3FzwWxNkkpCkGAG4PJr8+/wz8uOlBm7B3gtS95phB
u/wIn1KJfyoh9/k+0Fgrqxv8uUNgcnxRKMT0v4zdRZ4h1WjDerOvx7Sv+IsO49be
DIZzXuDiak59Pp9CV+0HC3LVtAJNx1SQau42jglu6rNyHd0MwZjHvh3N4tAlJb/C
yPZxor4+Pu+NOzkcYXzvacH37nsE/ioqfPCY0sckTHCqlBlIjXdBC3fXdq4xGLQm
pw4GA4/njO31CplAmR6xSx3DHSj5NSQr4XtXdKrjzUm9i7bVqBefa56NP+U2MWhC
qEmDE079iVuKAsxAEhvn2PAh7cbZI8G8cSHGqDgFbKjL1fpDaULxXl35h0PpMLXe
G3y0Kyr29D8LUGa8IkmPGpE1vifGyvbSEjoxLaVa1xspwiFhGCoOC1ank7lYq1hQ
eWwdUeM9UKBnFAvGW4FZbbtvpP0U0jHRbhLPtRhW9BoA9RTHbjpRPJZ4JZHMBsRn
MCDFvQSlQ6QuBw2If8AW3WKK++hVQHNSDNQ62jjBg3G/pYNiGKCUk6gdbahEBYZ9
q5+KOyjmiiLfq7Q8eLu3N4dCcqP67hYX8ePUWMTjmXGidmilEoWZWGp582wvfq+J
A/f4oR7L5AY2pkQAQx8dxCnB6W6zaxTZkDY3yvEVZwfnBKP1kBukqYh8TAQS4X4l
kcFyvebWxsAKub8f5RrrsLVWkTDHLfaz80DpEnXvaqxU5F2TwSP+hR/YkddjTmOM
FuVM4Cj8hqu5DmxZzFUDolRuKkPIz0REDRqR7yNnoAgjVhNUxuv0lr8aWEtyL5H4
SmBbiJ2Ji/WCxzMZpMNplhet9TaymbtnOV7ukSSE9GQyZiVFvksGpuaa5/Gpaszu
VxdETd9oLXXC9ir1J3bVmlsb/9bPr2o4YLyryjoV13wN9lE78SIIpjjzC4rMFuEw
aqtCHQEfLkRjX/qLkALv43NA2pSIh1ZzTu5lJkhruOObShTP7KYnZbQJ9d4C2E5P
3PTm2vtbYaYWWZpmBKNn5FZqVKSiAEEHVsmBsX4ONj2bacKjuoEM/QD3/v2gMldX
TEcVw0xZ1fJsAlKIr4Lc7myCyoZ0pz+mF+vmfsAxr63HkTu5PCJ46OfSy70xh0QF
4E5HlfefcyA8JbXhZ3NcCKhPzTafjiIzLjc2M4QiLb9XSr0NgV9hTX8xuZUNpWzZ
2H0YA9EkowMyITEJMMQucSd/qMJHvjU1h2vdlMY5yPPNnOdgu5Pyp9nDk4IZiqRe
4cSS7lfBjmlRChKM1AybCqsWJBtYg41tNaWrbZEEe1FMOmExf12no+cubZwFzrdv
BTfl/qbOtkMYnxSLSKbY5S4qyP0CgUBjFYAiz14d+rJ5vKn82XWhfhKwJ0uVrmg1
ox8WOPMflaIDqJ7/HBqPIqZj/I50BOk7sr+iteDAnGIW4lqaYZ9m0HWZV2o4dxLy
E8AANhKHNHkVadbGTOidKk11Hshhe6u6dw32NrmhHbF5KJuh8xkua3b82JVDswkf
me27qNA/LmqOFDSqPJWeAuVlsF7gcvr3woxdhlzq/mcUrBHqk+1DdlLysQ3an2Kx
C52G2LhQTmyyKlcTvK8FfwYcuX25/E/Vtz3zUgtcNkMR0oximPQ+QEHrFPfoh6/H
4I2gG0HanoMF6Q3x+uMEhRMPt6rppaqrxZ5oxFgCFVwCn38cXLRrfkNtz40tNbV6
YA2vF6RfsC/V6zHA8tZO6JnaU5pd0xGNHzrVaOh7D3Ogf8RmHOOrHOolGpLx9EZ7
mt8S+RTK7m88o5uKSw9DMZU1/z5DovqtXjWYFcMf4C6ZfAW+EJiv6iFZ2CSoQECa
Na35nd4s41WhKdnjm7PdZyIaXUCnQmu1/jPf20TMMqjdP3i+3iMANMbDCpUIhdAO
05EjIUn/4baitVU0lf5haaoVocHaKVyzAK5wd9JyQlji4hukbp+FGldnLwt6/reZ
CeiEw59DOvM8zQm5xbaRF/fLoSnJ6G1RFVW3xKVBKss+Zz0h90Z78oa+mE5iKflk
prTzWlOxJMUAUnCwy95sFxiDb4hTcbNF/DZIoKcR6Op/cYW/GHUH6yAqQP2KK1JH
6h5MOoSaUwU7yVJ7IupG4H6qHanhrAhbjxSsUIOfQLlqEUV3H1j+ErCar4XlLUaO
T2uQHJNZ/+RWMwaK9OFQCJvGDu9Ok+Ic4GM7l6sbNJhT2+E1AjTobebFOvXApa6W
09ewjkhUXPZ9ejGoObWRue1/W50MV3kw1YWArgtiBtx3//Jvd/Yk9MrCiEiSoptM
Y8ZE4Kc87qCEAdMDHuKtw9gUjbYbQwbt3rBEZJ6NxXlATyk4MadUCdzv0coUUQQq
jJ83DpMJqna7jNdBiB8qBQgo4pkVd+S+oZOXUc+yOJRK8RfcvXPF9sfYFOhuuzLW
nfk0Blj8RrASJk2EsV/NBgNk+/UOfyECr2eET6hxWOCSWNvaGdlZYlwy/uP6ccyZ
62KWDNwMrp9WVq1kO6i3Ar1svPAQJlxfRKZaYUXY0Ce99swstT2/eJjTaJ2hI8y0
KAO9A9dE7lliKKAgnkrIaGWveQaXxW//egALWoQNqZeRZydP9wifKq0knreJXEGP
0bO4vfszCS2Cou9fIlZakInxcVvCb9a7Ctg9XEXLDavwZeBzx0dE4G37PtuXQ7al
R1D9iXJrI5uoH8J1ITuQ4mEokbqcM8qFsWhiZPGaLiA4yacoocSQNkB08kl57+dm
pvDgcowMLd4yWqvVSHyMJXF8N0cG0o3bUEc9C/GXBvldhWSCMneXK9p9RYqGuK0X
Of4+YvNrOPJgHezynPMgRyY+sqTymfhwfRhKT04wqiC0bixsT/bQPVu532bJIs7D
Hvx7DksRdwAaK7YjwU1WuOp6BJA+52lGcXrlqMJZ/scR/QpLldBgZK4L84fQZF/T
RtDEDOg+t6HIVx90jFd/0CP/WNwEReA16ujbftY2trXcq/IrbkgNTPl91Eg0e9Mq
ZYOYsu4lTla2Z7cfxAPHu8wmABGNlkcwpTIVnjWgNT6ZA0IiljVg/55jBCf267cu
xlXEcLHl4IgXLbox0mvoRygmnkzzpXPCOjZN+7mJTPgOxp8E98Fq0vgTlmAYJaiA
`protect END_PROTECTED
