`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/XSJeHIljDSDAtCcRaAAifxURuzlxayHT0T8rlGHw0NYtNVyjF75Rrcj17v+STgI
zhcIC8Odq1blnAiO9ie1kKNdz/abpMnm0EKQK7nLeBYd3rdWupsxXizUzZ76Jhdh
XIjh9WWl6MESW61Q826Ns5Kbwb/sFzzLGnvhzbGOJMq3hP0b3nucevu7m75NV6UM
2J5iw0HmtIMhRAe0LMqxCCSIwpdmafPKeZccEDgKz5ZmEWodI6nxzxw4LiZcwAUO
sGoDDBXDIO6JAGygG8FHo5j57NeLxyJdJYpRipe3jV+ezPrFPhcH6gQVdvtfpdJc
MMYAeTyEQS1WOOsDCgjqwBef/Tc/LOjKZHsc8JCPDdA5wIxfNBX5xQaD0VajSeGV
8/T/S5Qg4ba6bIq2ec8LKkQV5Xcpl5v+5Eko3e6AJ2ceWKvW3elcewsRw6kQhJwc
pAvs5AcrXmrKKls17PLMZw==
`protect END_PROTECTED
