`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
neWaP+2hep9w/LzuFdpEmZbgL5TkaJW4N2XY5ozkzoOnGJ5IN3Mez6Ik2gdhFJca
Jiy/c8uPzo4AAY2J/vMcISYbJz9AOm1OULIQQKpkdhQes7AVFGZBhEDMge4Rg1cl
cTOm4sgVkqv07/zLIEab26srT0nNYycxPHIJtZnwsiJVYBtR5kKsSubyrAjo75Dz
Skka0A+oKg7VfOsGX+bXjThfktSJArk7cTxFIHRzfbHpwkTl0ux9hAhD9z1YiFlj
zkqw3CofFhUvXSlmXu3rH2oN4AQiuD6LXBGKfC8CjPkcOKtFDj8nxQ/W82EKbaDq
1Lldk0EPu1agWLIZwk/FMrT7/ys0+quFGn4ubV7MCypKK2blXDEX2ovHepRmHghf
rzmwVuzHe8g+nM/t7N5wSm3VkHwf1oaLf3SkkJvNQA87DI0aJBcS2VK/bNmYPgvc
zxMYDAQKJm/mnzBpphx7Dj88v2DZHnte0rlms1YMRLyxXsnfxLorU+S60W4B5jKy
de6Mi9dt9E1+rhdT5c96qOZdm29eOsVbdtn3O0Q+vDGSxN+k8M2EJpzwFT1DXUTv
g3n2THodTH0CbNE6+DG7ANIKsOiYBfdrxbQ8H2GghBbBJrvukttUOyzQfLNH3qrJ
3kJnjy8ESA4P3LB+u4M93EyG8gSsuSOFKCBFT4RozzLznTrW8eeYGozTJaz2GSbY
JPS+yiez4VIMWQEyd0TqMTHiLk0MrY3lzAephF+rpvqlJUHh3y5h17LKKAo80A6b
AriF85Lf+mZOVQEAjo1FXo/1PpoZQp6std0OCd5yZnqzML2Vujb8wuViKLzr+6wS
s7qUyVajYz2Cea0VOhAXQu9lHtk+kZcIhtxeX4MgdqDx5fXrahSRXQ0ZqQ9vs68a
/RGwR9wePBsLAlfthQmyzPeGSLxVbxs/tdQUqr7eStw8yJVzGO8wotuUp3UY2b4E
`protect END_PROTECTED
