`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uVfvDoM5zwzzAon+Sk7aNEEL6SXPnMw0SIpXs3fydjTXP4eGGEx4GOssfqvOP9xO
A6Prs4T2GCuNyfDK1InmWcfs3SvYX22i2OL755WWJYiw32PD9zoWqHwbHGzRUu/j
GlB7ZXOusBKHewuFeNs/Bn3ZMpzxCHW0CE7+sd5X9V+ne41SBHyQeKTTJXrp9Ck1
2b0lrYmGu6ZBykLXtmmbBrd2qxDCfAxpduqNiUxq8+XPbj6RhFJ2CL5xSWxGv2EG
Csr3lUAjiY5Zxg9cWWJYBqbYbRJkHfibiCrwbFQm0sJNyCTpAYqu+Xc3Id//IOGH
AkzxNghsVUi+5t2ECcjdeskX+7V+X2KDN3PB1kUjHytwuKV7wTDLxSpZHDWPU4U0
vefkN46bAtjbf6J6istRM/1cENiYkdAyEVK2GtcQMZBq+t2XQrrWtfVEXkyn17ec
8yLqwwB8eg65RD9OP5xS1HIZtsFiAf6bjAHuR/IIv0VJ1X/tqtcx2QrsjAZWWfVT
lfykVZ8RbtK520lkSM+X7VhZyVJYAnON7WeT/agQV1vpaIEpLvmRd/Xihgjyv+QR
2+tNc+aL/vJCpPNMR9i/W8eQWz/C9dUief1aZJjhBR3p4IxieaWqHuWiZjOVDhCW
7CTrlWUjN4y97JUPKLKOPt2MEkm4IgAdClrRMgPHO38ItrDrwqBoyOR1YSBfW/Sx
WPG5EGcX/jAlBFeEnGR3yf5SdCJGRPmY6pSl8anj75NyrQiBJUFtB2xb5eoy46f4
F3z2KsPlCL79o1dIgfc5+mTbIZL2eiIJZUjrKdsVb41O0RNB/+uRM97AiSmjOstE
dTkFUGimhkMmkQu8Vot+ZkEnH4lYmspuzlmPvczEyPvIuFjwCO4U3MzqwcaPRE6a
USGK7lA7tq50Goox4VId53W1qMtxsSCk8OsgwdLl44a6P0Mh0ZGtP1q+XpqcqkmB
xiUQHI+/WU66IaLxcfmFJRdJrLS5tSQ7DWqCpuT2cvHCmwwt+kZ3T+3kBoh5vxUh
`protect END_PROTECTED
