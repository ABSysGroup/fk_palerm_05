`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5SvAFUHFHV2n/09Md3372VGfCxS/1AqKYMuzz6+K9t848em37tWGPAxTICRkzgtw
HYYtB6/YxbJjPJHyxYzPMPAq/mPbZoOhbP649DCzFqs+zsqeQ7FTglc3ntErMge3
l5SKde+P7qVNiQP4ANGpHEBRPgV9CuU446RZUk+qPKoCj5dv+P286timrc+Gzlln
ZohWLcW3+ulpbuuN8aqv1f4DPBgwigvtjqd+z/1Zj69Io+hm3DLPRnzIL3YxtGYp
72qZZw3UYqfsOkjv91Mx87UtTfen4hY8G3HOyb99ev1zJCL2hhsmPkjJBSX8PoPc
MxD+trs9gphGeWUC7V3TROBp8AQIDtZEE3ou8VBdFBEZQvCnDLEYl0tt8ZSYe9KM
cQmBjQ1vk7A9L3vK6sN4Qx+TN5EM0kU/Tg3ru4YgA9C5X95wfCNsgSYzWaOtwMMu
BeOx0IJePqff7gwLzPm1XetQKd/8/fPT82q7/sK81F90BpUr4zevD3KPkQmdNrfb
PMQw78IoZx9v35TT6C10C5sBSr6cJNJRLhXeGWUVuSZGB4wwJV02v0Nw3RP/ra+g
y296K0dBBrQKw7gQl3meL9+y1M3Fr1TntNYPfChE1d/GRJhoEzFX2CPA+EILjTc8
mh/kVGsMN6FgjIWp3Fhx4u1Nne+0QrKhsf8P/haL4UyPRG7Qowa8xBvCP1uzVAwa
Dk8a/5WCPNtZz3H/YPP/gQ/Xpx0FKK4f0ivBZkAkTPy4L/zXjzDVognmxiKjyQAZ
F0e1HEiZSXWmYcAvW9XmJKaLbLiZK5oRHYcT2G0o69QHsn38esDvpbRcOzhxeGkG
W0++kl37ebSS+4ats8oRxSxf4hT3oJBizoeMiooERYwYEwJ1zrLjE4X87n8sSnIw
2SV7MJ/bslyLmH+QBqxkCYK+8saoX+g+nV9xaK6vrwtMQL7QDDKig6+brGnZRSYL
Qk3dt5wOvcqxX3iCt7zfSuINg0QCyDytY876UnIRj1YPSvmREMoCEdbmpZkDB3+4
zUQylvblT+DrFB85j3bL3yr6XlTgPs9jPm3vr5YODnJpZiuOvaF5zkfXIgkWMV0a
cD1mr0XAQOmpDI40NzT0lNwGTlK4m69J6cS5vKJjalE1TPUOt/bXEAaUsEhXtCfX
0v3qPCarYxBhF5rX8qSDkifdM+pvXjYULEe14nLsH0oeYzxKmCOC7nieQlJbl2ZU
Z3q336y8c7yK7pNH693svPIv7agXl4gq42Qjm4QhbD6imkjoDLJwhlR/UKxI9OtH
dmqbvpjAQmo7CI6QCwG+Nt9dBdFXXSxQZ8Em8XJHsz0QN5MsYfXnMRZ73neVUNMS
BbLnck/J3y2l0bq6lD/p2sNNYZIjuiEG8i5oMEerVlnojK7dAkR7OEQs1gjxSLlh
mVYyaAIsTa6DMPkBa2Vo4hh9EBFv9tUet5pgqBTk9Jo1xjCULKsHZ4F2U/eqs5DE
+7HpHFtHdbbUcsgrSNpYLoVBbVmYs8iF5noU+IK4C5cA4cLzVNI3natmVNJePdPE
lRgO6fwZ7yAqv3/1SJG3SPYgFoU01o1GuMo42KJTzDMU+22TO2mktXG/6I0CBc/F
4d5/FCfWuoQb4eDKh10LQuSDW5tmkkH/ygl7uTLO9oPexdGmBaH6F1IASJKtDiV0
CNVLDsWIaPU4H6kqGjiG6ZYj76rVhqRSVlMunLsLTWIBEQ7dJ4dk7ZQeHr9wcomT
T+NeetSmcXD2tbiQb4ERm91kolD++12GbZVolsuq57Mk2TBiU91Z3qP8Ej1se1Q6
jaNIl5rj0Gd08JWICqzXQc1kZIYIFx7v7f2wesZzy6lRlv7rs6OfgZLOYTSK4tyF
In5HupdGDYBYmeCrRAHyqJd9wC7cpk94m6BymQxU3FfiXy3A8qtpdlFydpsGlmFJ
ifo87mxrrZ2ZOSC3JFU6aCqN1hE6Iv0Ow6ZVK047hFz+QEDDBsuHsMbx8hXfFGBr
P8Lh8Pxx/dGY3An9uoEQLPFmETvxW4z/+mjlEUH6rehNTWV2OnYksybuHHfu/3xI
dfY80CYe0WTWIV4AHA2Y8+I9uzW7u+d77TwZpZcyN4JIwwbslDCUWJ5+tqNQlTJr
kvBcWHGbAt8L1PZT5VzYg14bQcV5NdgjRsYKlcgm6QBRiRtTbmX63rP+KifAuE4Y
JS+wHamN+/11rNmFVeV/Y3odUcSncQZFxJsjm05mSpzO4gUI2Nt38bcAoADUIo5j
TRSORrjUl75TK2OjJ8QNxbzeqfwgcxXsWk9bkytw9fm35JMRX6ijMFopThgK/VCf
VnUq5CsOY9S0MmLC/gt0tcP3sLw49UtNJ8pQbTUCY7Uxeu3cgIvyR7cZkXE5KntM
6zotyD77yEu4V2chZvw6P9P92PzjJrQy+Eg76L8seN7t62uBCkjRr82sFL4Y0t/4
qzxOzStys8wA24exJ5RqNUjlsYsag9qr0TQuNv1FbXqNXkCvknyUkldTFlkfv5aO
Fc5KMjzTar3nhJzDhU52Bu2T7IBlndm++X4lRuNi2vcU2m8RVs1TXRHIQ/W3YLPM
FlVVvCP++jt4o55/t86KfxGg+Rg723xe2w0r/Q9PiOvsft3fJ+ncii0sVi+px0ez
7DfrUtbe7qLSBiRle8tj/vgFnpUe/YYJ0Q2JK6eyQReRXDyPQo/zZxri53EiAOh3
iOPJIL6dJrZ5/1ewyxHc42XaNv26XKpB4e1HlIFxY+Z3wfik3zNbbhPxCTmnKf3H
kWMhJld498O1IYXb07HX1k+y5nRCbyal26vSvj109PwPgBwx7RzNqtqUNCEZyi+6
+Teq4iD/4imyZRcILaZsETmaaxzGFUXnGiw7mz5xS+Py+E80HhCIgVH3esrU0+sl
QF9b6nvhlHssrUftxgb1aFSPko/mcUxr0wyjPq1sFnQcVoGA7camViUpnBEOlaK2
6Mp7e+jLydt/0JeFC3L/BfM2yfDG0YGSOTiEqMXFc8xOph9IovUzkn+utRxqDASb
XR+Zp0YrfaCbKJNy2Z+surH/k52dtVrrw7ZTXnCpebtBHv0laNwFNll/fau8f6P+
OTE/pdz8SMbIr8VaQxbhWD/O80ChJhMqJujHIMMapDrWPduDo0R1hjlPQC7oxxUC
07RrTFEsUAHc6MxFji6RkPD/aKM3L9FgeAHun+rV0WMg6BohA14sb2iXPIutChU9
2o7SXEaqn3xWC/A+4MaEKXJAW10F0ZT1QmFPRiN/WX+i50M6m9HPFwkRVExhgp9e
rq+4ymja77Aw3aiFUJN2EXRFipwwlYa7LaVuHqDqRTC/hFl0tmtmNTigOpv1j1v4
hfvwWtlJiHYQTl69Ap9WpxJdi1Ph9hk6Hr2jSJ3NCKSX63pw2HOWzOovJLnnVlII
OvCqO3AO6+fFjqzaLu1K8BYOrZ4Fet4Y270OXjejN+wt65eom7ZIPf1/u2N9lbGz
Je1ovpeb9ssPge8P9DM/ND7a2rjHddBlALxG01MtGqimJPqsyW8eq+RxI+FNWAmt
rXg+uxbuyLbzGGsem7JnJzYo/Y2tZrYsF1gmtKEKr4ymZhx+1br2YLf6bD6aGq0i
EYngtSvqPfu7EtF0N8yLULcw/mMRlXdoOCnMyTEMRjk+yVt7yBm/yNXzMUA2d+9N
i9HfR225BfBwPdIsxepp83YhskIQghzsFIwLB9jWVpZWDI8ohG2K0xqCOh03jDTo
mc9bIE7+9eaWdLpih8R/k2Gvdj0APJ23qR5c03x65mncqchvrNOkkQVrTc2Se/2T
mYf1hIrvJpB4JodmDZSDjHB8BRJgMU7IIWTiRJZ3lN5KWM+W8Mm3AroFLZ5i9dCh
5bQWoRn+V7IJqvULlfMO2JhLK1WJf2CqwWX7aP9doNnlO6daqrPw6vU43dnKZVk0
h8nZ9E+Z8QrWdAoHj643spGVLk75zoqrUfj9QBiRV5Is8aIeIpNHOIAQASlP0Def
xRz2CCsRQGjP8diztGk6lwmqMY18HoPYO6D+Gc0DXh3gDv2Lt/O163/1PrdHL/xl
6gEsxzI/o71KxZKxoE4rdtUBFnp7SnZAdxe87FwDBzATu4wLMn71zR/f/HTCcaJm
xvUPScKbzLHdptjgGO4HiBaNlEh5Q9XUpHLvW7m+bDBK6bO+C51+OQfGkZRNpudW
lUBZW10rT5tZV+iw+O9QsQX7BinXgK3MF1XDji8OruL6nTh92Ku9e4znqKNBdXxj
1d1SVKrM+ojoEB1hOD3zHSLJvuH4FBJErYTTppMCgwwp0L1LyuhByxrpDuRouHOx
X15OmKNrUm4mMcY3VgNGCKKXPIzFHN7B83YDQ5uDKSp7a8NkfRAuHkuGa2MxdLUS
tIhLN8FozDVDPeiIDpyHZN7PDvSJDeSIpPB9Y/K2ZAbdX5NpSBQR6fNkcRBntje5
PioJni3BI1fO/xLk3bXAyGIqszkBhQu+aIr7UoTcq/ImsHqCu9JiEYT8ZsxXo8bZ
TCzcKThxtVcrAN7w8G82D08/QRLUj6WX9zut50yThvi4Nc9qkhK2d3qAd4Di8ecD
76u1KCcy1c+X6bvJjpWOBo6TKyOOm5Pr/FAio4E5vCX/pQ64aeTdg2k0IXsPXJMY
m2yDIl92CHwnfmlycVmQfVM5AA67DwlCRllWvKMdtYt94lwUH3PZIdTCGF9gCYxE
Qu8RWJFSOHjEW7XFf9TeLWPeivhpMfFwNQ+EqoPRRrYzs7TNROCs3DKzHfi4/LJK
cMQeAp4iUsBSqrPQGVjBvTjg9sFRd8iD4pBXJgaZM9QrrhRqCeRZ20CoDxM9XuQ2
/DI+38FhJ4tptpmsHweKKkxlpKMMlVIKkYXpDQsOiUz1514JIw/Mog11nUz/uYOF
EGgEcl8xK35L1QkJ0Qw2PJ/mjW+WgaFn/rGGFIbfy6tCnDy/FETffhCbbQ2nM+qw
NnpWodWXXywsTPTdjc5V2knL00y97YRDkQ0/SNgITWBkulo54aJCpk37qqkK92VB
16k7bLOKTszmklXFGnG6KaUJY23d9LE0FbcXqVTRp6PbAzhEIOIVd0v9JoN1HRPQ
FUs1/Nrp2oAsbQjJreuVk6FjJFoK5OjARfvi9qFypPRid1RE4Bq7+i2SGQG3xnQ0
uZ7W3TO7i4b0rpC/xx+HcD9ISEfNigeEx5nul7YTfABdWXzJv0dGdc/O5mzlytJd
l4dafvlSenP+tOL+fQd+uobnOATZjeRnSssdjYIbYxJMQ7ZJJTpV99SXdPC+4V5S
bsKjeeDasav3MWN9Zizl0f+BgYHIEFxq7xcw1I8NjOIbaANOqdXy146T2+jb03RE
UcgC2siN62faivmWWOs1EGi6F3YS+cNjc61v38nDchCYQKuSvaW6jpra4MVa8HZz
XJJw/vooK/Gr/QvxUkIcUmEKOcIWnub6okx+edUcmiEQVq9nR09vtboaBjImyMw4
PiN1ABD62L6a3lixj4S0L3Ekilhb930Mqsq7TnS/32nR+AJfwYBQhV3V3TefW33O
Hot/mftOP1f3J/gih8P701yGBnNGdQY9siYCtHxdNoO4hk9vtQ92NVmtyXvj7OuL
rkNBbfmNBozi7NQhsTCWADVj6LlQI0JgW43eLPxLXS2LcTQBYUrPJqYttodTitU8
7paS5J+GC3SvYVGp4b17IWuU4n9pLCL/Kd/1CQTzQTa7MklsxgDp9PzgXvLdG/ng
Fq+VfkKYQ7sejhxEWgErfBlI7zqOG4OnYtC+n8BSIUpBABO48SP5MGB7d3E8+zO2
2f9yQw8Jr1SjPPOoUsUbG/rtlLyAC9DzZYkweOuAgroaqXPXP+QjDQueJzbB/a1f
lr0Z8WbGoJ2Dk8Go9R43CA==
`protect END_PROTECTED
