`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dQlOFlwsDF+fhp4BKMlAs1oN46p8My4ufqTANFTF+6qfDEUBz6hcws0X18xEhXO8
upMQu3uHPDs2vkQXSLz0JsGjLkvOA93t7zPgHI8YR0IuqkRG8nUcacod2PpbCsX0
2ZC8RdQYVyKyr6e1az8sy+j8cfWXZylkAm82ESwD30s1Zc+nvUx3rs5hJRxIS7BM
9ULfiuuZQw09g0Xi/IGxSK3qcO5fD+/pZEiuIicD8Em8FRokFW/tlwBQAToCvUvP
8MJGKzreUzGoha0cfkAU/qFPoHxaXZPOWEFYRDiWjey1/1CyQkFRzHubYs4aW+Xy
hNZ7hj4rHysUj8CM0SSP+0OJCdyrFkQNVlvP+uV5QabfDGQOfGXWsEsfwWDzBbhU
vwPXq+UNA9+tVmeX+KCLB/FAqnva2vYDhfoj/ms6z4w=
`protect END_PROTECTED
