`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ukCeJmTZRVOFJtDVImVp7cCTa12VPyFUu70Pv8UKP5RrgnwTRdk3EhjTnrjbHnMJ
tNDMhqiRBxYXXxOaqwk0kPvaZRi4xJaJ7dgjlY+aky+mHQx3cM+XrkhsZGdMMmuS
48bEc/ZWKvNaDPVLED8hKu0z5Gd7DCZ1avJ6SJlNfXjwk8BqO+pakPBArQ/nz8rY
53CYD+rQuVSPCywS1JF+lKgjlI5CfafsMrjSjIzIUgcZnStaAWVJ+juuOQP8PJoA
nESjQLQ0XQXoz5gmvUWvYSS/EP70VJX4pbBVXwwbUE6AfZSaFZL7aOGOSwEM1tKt
SyRTDrWhxZuPPIibm4bE14+UWij6KD3piincnKsgWChCDs+sXpLZmI3O1MhuRq8v
bMeYEfdUMTxftX6xSUcKY4pIYqUfRdHtuQHUjQeFz6ieaYkuSf9bYIfkAemdzo4A
6HvSvQRwmL/P94xXpMcNSA==
`protect END_PROTECTED
