`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8RtxGAHsrwSgrskK4+Ngqn+aDMkv8jCOKfMlAJ9U3NPN/J1xyV+vA1SAxr+gtn+U
A6CBdEcQJ1Fo7zYi4ypR+z4aHPOVEiNOo45TxW4gxBewpcLaD9QU5bPEU8WW6Piw
skee7PIF1TQgiJ4/mzmzSN83W/ZUBPxHyJZhO2/Bn4LcDo/LFgGtvCiid/ZaBbTt
Y7HuoOLAGa7G8QgbCA31/tLhNrplOq7DoY/upqvAvRIjiEHLkwY+juqIsaL1j8kj
C5SDSYuvfCHFYG/p+kkMqcRWWSH6SewSiVohHXUtoMWp1ESkMCSgb7W7CV1WPP77
SAiKHjip5FNUCHfeNV4JDQ==
`protect END_PROTECTED
