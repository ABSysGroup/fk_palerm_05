`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mYw0e1XxgZday2cG+IkJtAy245FmC+arzPDhfkbe1AUOIRrc8QnycpnLYu4aYQqU
XeR7xABuqlAQiM4nAAJ6T3WuSXxm7H9lcFbZSH3IOdjcYAZVeHZSelqyT2NQL934
hOIGfJsGfxU0VXl3BvLTetOz6liypAkHrn9gJ5T60ZNaJA8gJjqlFCOcmveN8PJQ
AQGqATN7oeCTcXpPIYqDJhQTEHZLN1RnjLdBH8NMGSCEELeehD2V1Kdjwq9wiAVe
K7n84/REFGfVezF4J2m098QJRaEZ/v2xcujN0URGVKcfgUN91B4w2Rc+m//wNZ4y
Pgku2efBZ9XoQHdQ+Tie2p0gmn6XxzxONzGxIioqeeDS4XNErwJXsOXEraly85DB
j1cdOY6sPJbZCQ9OnZrRwgEUNeRkgo340yKMcHzTImtsnbDL4cWZF4PHFPGaYjod
4S/LuQWxK5eV0QIEM7LCPOvyfl/BxhA+EGt3/uJdmAHW9GvprmTa8PA0LROZMiO1
Qkciknmif8X6llxcufVnrhmAkBMbFCPIEGlZmv5q12Vnp4LQ3wfOT/Gd0PCPFXMa
TLyWFX+d8hf8X5gHhgRxiCc4HhfDAQOmWRjuZw7aRyExWKSr1V25SU1Y5id0uDY3
RtAcNM/1UroAtdGANjgtxGD0FqKQJ6Jb+vTeERlRXyYJKS7i2BPmxH+K/bV+DhLw
zc6BlNVPJEvY8LVDMJfXvbxpYlt3ImFASVucTc6SOyRmJjk9nc73s0Duh0PhpGzg
IfJcSEN8ltPmPF8y7apxew==
`protect END_PROTECTED
