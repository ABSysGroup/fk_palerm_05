`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8KDjxr0oXyIyE93NlJ1W0ufZeGHq1B1B+NFFDPrG/6P6IZKGPUK1XhJdnux0DN4B
Jom0NZVh4ZOytCN+Tjk/X0ZvcgO+f9JME40BoF8RCG45YeXfkZfOrY+T9oa6iNCp
sndL62xL5UgKg2u3Nq80ajqPMz6duS9e9gN19aIz8U0OieTazVeuf7V9R9QyXavY
mXIu6Jr2RNCCsAYOPpEkTufXgtwMW+s4BrIrnwRgfbeqGcQHafY/NlLzThGqsxCQ
yYeABAzDUjPEothdWgQ4bjvm4cJ82kGwgeCVPRMfHhcs5Tj+z3O1fIl9JpvIJc7g
bhvKOx/sRz8/v9+QTU6RUU5+1jOxIxAy6il7h50zLaoWO/9UcOY4wh267t504XuL
/81b08kCK6lB9zdIIH4zS07M7bwVOJMyroI4o1OUd3aU2bJmSawT8Z3OZybFNAxU
PeOIqHb8UOQGUqTBzZnZJ/G9UMBD4HQ9k3ff9bIPMyo0kJs17bkbxiIqvu+B4lir
KhDhA+GqkEnxs2wCU/d5KmIr7F2iZ2KpSYrPbtPIXlheKIOCsor7tND7y9Wgmv8T
M2ZLtXbKm0U6pCG5xdNDo87EfpHVTglUfH8c9jV+6feuUUoM5MN4ikzAjqzW6n9H
YnWYQE8Hw7v4ANQLbGYUg/0ZZv3mo6k2bhvG+89BlcabWrCzvvHY6ZbseolAvB3Z
pco8+SUyJg90AWcRD0IlmGU6tI2h7Hy2Bu3yu/ZW6hbF50NGDHDghff/rB8ajF4s
gYVT/WHAnYETsBn6GKwqANuCIWPsqMRwm5LDfiDSjoxZNpK2qfTIEeqaSEwwTHLz
`protect END_PROTECTED
