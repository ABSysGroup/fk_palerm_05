`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1e0fWxB9m6jdL1/RMRXvVxrpq62DUD2BLDCImro6mVz8cEHaGDbuMtbx3OEC/tEj
VYkd3DFt6du/GhlnhqtBcAG2IvKnpcNuat662qZKk2ONBpogyKZGes3ZjJdSGQZN
gpTXk0vA8XXuM8liXb4w9eVhj5+qdva7C6d2JdjjSECjsxuV8mkDBawrmp7zz+P9
fgDnAcRXS5vwXFMQ6L8c0QzQPzpV+WVVAK/+MOBJOUWQ1bO6EEft3HvIeiSxkYIB
Ks4Z+MVNODfClIRqkt3uJp5z2bdsOkg00RR5cCds+K0mZ/1xEaUP4+k49uxZ1mIf
h2eHceHsOSjpKhxAxam/G0Fw6PHgJIj/ECZhkO6sD/E+bkpPEmFVGinHejFX4Opp
zEpOhOANEZJHX0HxxXy1p7sPVGgoYsQKoUVu99adgob+uG21aa3o3OpKpmT3zQ/M
N/LlmpUz0tWtrj84L+Jm3YiibgEaFGXfo4jMW05o76TjGfmzGdVQVYGVATPraFwI
Gw7ppsMFfvY5uQ+h3WgZL3Lgn4uUA8X9/Y/8tCoKGDj79yVkDimE9TNG23LjBDu2
fhOGYtMLBGzKk3fHDwT5vtHDKGOQePJ23Kmmk7YwUrammq5KgVPyWE+98zi3froe
3/9C9zLC0lbytIHbeXH8ZxVrTJ3ZEwEnwZW6bxfWbtk3lCQr4jckhIebosCjkIag
aM4T8xl7oipT3zfiD7jAmFJtH95oTxgVDEra2HrfIYxB0uoQxdyciD8P30sD/0Zb
rWLA018XxehtOY6cz7HDloc2CZZevG8pqv+BaeNHW2DAZw5tga8ouStej6pfvGrQ
SLj+icQpCuc12QxYpcVpfCdKe5UCDkYJPzcKC5ZSN3j0ZvfD+HyiK6EYKcmcXBPI
R4cMdBgxEMMAL77yKktYEp4IWkCXA3TasJJhYxoNGaMixHTxP/J6ABqf0V38ns41
C46iL7wHNPBpG/0FzSjRYJKsDA8n630U7bUW1CWHQY57sRkagbNUBUKD5n0DI6ut
+qFnhohFX2zmNLU+a7o7upgG4AEC8hepdLowndg5FTw/Z919rrnS6yDkTL/2Z96I
RBj+li4CppUo1oeaY7Uc/wJWKf8LF/6L0VPpAlaVpMXaFjwW4LJJdM5JPPkNvVvE
LNyhe199EH7wkjuHNkoa8swxAZnW90PDJHTAFDskoIp9BL1pYpftESM1NxxkHQzY
a/xiLhPdsTxCuXiWukxB5tOikW6sk6YxpuY1b4dqtwwUg/RpoiLJKTE2G1UmeMsj
/h1Dv92Jcv5qs6wnfT6E4PAFnx9pfVmtCy6/zaSWyrMuYSFE0WzSKbYWmtoNpQlV
/5ZrpEHYCscTmVnqjatw6SyweSYUCd5cSqMndj/UYl6+skS186q8Twri/WJ+F406
mjvv1EfAQaK/gr8OOwEaic8E8y/d9KbdiPxweBJj499/wEv2oTolg33xwGy/NQzG
`protect END_PROTECTED
