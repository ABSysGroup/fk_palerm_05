`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8dXm9ZzyTESnb137M0Gb3Ey19Cqm6q3MDOLppyYCdDEyg8VgJZBlk2Mt9GlCyhPV
k0LZJNTPD57YAG12pSb+D5S7Fxsiqmf1njx16lyOdL5zob5SkmBWnYI9ZV7rPmEM
HF7phqVlxMzx18pdmD6nhOCNlyoNhtqxEXWVXff9ARBFLn7tG6WZwktxHm8AurIR
Rx+YMH3w/ZVyu2OUqJhY+ge1EHS52LtTw/kQ6iEn/lxbBGQ/1FO1i8y92p7BIOGN
JDAD0be7xvaRhA0J0R6tnQ==
`protect END_PROTECTED
