`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i5Y2TzIY9acojazLbWoJKFlQ4xVyfoww9j/gsU7KLz7XpNXSrsYV1+O2G+EXiTZi
j3f4wSyvUWnhNKjkFTxMIMs7+ZlF69JkP5aGJNjVapotJdFC5FEWzuT9vF0QIEmm
lBTBvAgnIHjAVexSmxi2nT1cf4uxk71FKDf0iSp3vvk/MbNwNOkpLjXPgrsdHEVC
uP60S0gTa0fGCmjKVMYGxyVZk0/c7ppU8FaqSJxF7Uf4qjq4cyDy1ali7OoBKwWL
RbNNv6qvkOGG+PdizGdz9PGBOyxKOTjz84z5+XduM9k1XFUmbqsSiIwmPYGzLSaU
9ezSVPMHv7Ik1hDE/cRmwmTOTavKJ+9UNpyohAu9OuVZYOyu5UZTzlml4PVLM6eL
2keR7M5zIc1YY5e6NyaVyknkDAAO7sezvozwO3KR1/tSNdCf2Ezl0yHhHdNKpzQA
ODjCdLb8UtSpaZzGtzwd7lZCkdgE+ztsJbnyMsbz8ISigS/EgTzz/quz9lL6PeFS
kXOThYA9/rlVrtqMqg0OpPoDsNNc30JeMh/5c4fPP/XEnYjsJ1C5c31o77pt2FtO
YVf5X2ptj1UR4Cg/YJZ+pg+CUzQeNXcA6G2ik49sE43oeh3URC+bwvGEzZVXBTt/
sDOe3B+9iyk0/Y0BgZKayfKB8TOzFFTX1QdMXBYjncVncCJKJHg6K2oTbVDOwnP4
6F04bs/HJ7IVaoX3dMGZpypg68hfXvwG0317nznG+5uTdpXwB0yxHYhlSMCAAdrE
elklnfqcq2auva9uR59B1ZmlUEarHfoXNWu8eY1KUfcJQio/cZcBJc+RXJKhD8KS
ZrmpDNjgrvWHUuYkDMfKwyBF8SafFLwPmIc5hSTtDMBmfRHH41ZGeKTbukQXF9bM
6IuS13p1ue/WzwB7jdmgsmOa+0SEA0pIQ6biU3PfJQBbtKavcVStcIf67QJqWF6Y
ZMYipHQT3dbOGSrEFnHvY2LOVADf+wkNAnq1UZqUGtxUqYY6764qG37qYcNUGgTD
UG+ZC8OAcs7zpu9qQSY97dPVos5gp88aj+UZ0VJjNgUb64Gpv1AOHV9POT4kvov8
KF39W5GuqBAmriL90rtyWuKxeUFtRY6i5jIMNcBpaSmYksuqxJSvXiRNkpkhuJFp
aEc/j5/FKq++VPdXI0zNWXcZlFjp6k1brlob0pGn4CaBMMi6NMd3o0W9epjk4RSP
rh2x7kEdEDy0bac7ClwvBiCYbwIC2C7yq58sNVHu8Pf/KwLAtr6I9FqpSayjnT25
rDFYot2rAFcpZLmazT1O1GoItzOTpN5nr6eH09xdHkD+pO1MCZkRO9uj+PM06KMl
`protect END_PROTECTED
