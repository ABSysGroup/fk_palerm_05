`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CSxe9SFXHJoEK/eUSNNmTFbper7bMvRvmubi9w9BA4vf0hImx0rMwvfBUIDV7tP6
vhEEhcItQN41DYkeiIVHmCeks81EoA2B8uLhtHPoaI1V4roeJcuMZYH3zLZmC2qX
UNPvZ5+2woyHJ4TD7nVWMqaZhhIGOO+oJ4FNybEgQf6ege5hrnSiuzIoOro87NbI
XcSNMfVqBR8bIIqj40dIznzk6AC0Ksrpv33g8X146VMSP3YGsU2ouKiPtEnEqt4T
gNP+8PDGE/zefQ7heCrwY51xbXIJkdUS+vkjGoZqw8sEvIulL/6fOaHd7TwCep9E
KlENr7UI85SDG4ar0OfRaL9yCxmbtoMJeHcs/IBj8hN+0pqt1OTM7cqOCzAHPotW
eH/BWQ697OV6aQwn/cIX4Uuzaxq/X3eUNzUzQ5MhPYfH36PARHvzPqDu0HkSynfH
epX7NcmbgYHyhDvc3DP84CEVRPnfZk6pdt9JYkXeUcdnWcUug2jYEzBeiPdyJh7P
P+kwfLeaXYZMMxR9mXNnfPB2jpIKCxSfED5WWqeFQXrzg0s1zvqJEIaEk4R4MdCw
bYNHrVCpL9feLDJYB+Qm2Q==
`protect END_PROTECTED
