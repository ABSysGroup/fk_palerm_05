`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jDjoA3zTqgYDrmX90SbyFvchHQ+DlsaCYsnJmYcGjFvwxrKM8Q2ICNoO8G5PCxnC
qPsZcQnIeNrXHEAvdCjx4g5UJYSYs95psvKnLL49R+oivBR7HgAv1TKdd78yIE1n
9/b1ikQlrmEAkKu+IW3+b6L0s/jSLQMgD2Y4Dvi21VuJ7bwByfDH5Sj2+mMF4NXo
JQzOIRA571axMTpxk7/NX4RSykQ+iB2w5N8xukQjcu2UogGZJPzY2lO6PZoOE6wL
QTaUbkCKqlEZYFNoWytrGxSfGKq+RwR5yulTDQ2tYYkJXJWxWFZetLMRHEESCTS1
RaKurrIJ7WALHParCxcP1Wd4nCnfubny/m4JyokXgda/TMvFfn40WYkow2aq8S0a
F2Nyv7IeH+/efQcER2OIx+7rRyZ+u4gxmjHiMScrtZFDD87L0dluz7LHTYG/fzMA
yrRKpR8TBcBFv4UnqTwtpFopzslDKNGMf8wq+knMYF0nIS3ur4abPnZenuSnCpKQ
xAGHqU4959LyMsE34WUG7ZjLAghaY5LYx49k5XaoTKb4/fGpWPzu6E+nNcc0lqBT
Pr7OCSO4nR1bjhpblhXYykvAmPNEn02agrn6Wj2vGoz8Up2StXn2PkrfeDyQMnZT
nGnyf9NBFMGE89mt+/IgZwdLrSCK9jIppYe6f9VW6VRSrrUoxUnCx0SdccvxV40f
NyKQaCTcs266M69wEGuUXWcsGmR+/tqcw11oTJcVll8aU+Rlr3TPl6pl4UxHkaqe
MdCtaVVj0/LKiOt+dWB6FPyhn6/WwWkhsSnVJBY4Enik2l9YGOzp/sAjepV7QaiX
D/jLVtol5YgrWYZkF0Od9X6Sj4qAzZ8HvCkvKhPq4sk0KUtbvea6691d+7CruN6q
wHXeJfZSxNl9gyiNn159rvLhy+AmXBe82NaccDhFUFPerH1g8f3O9L0k12SGjuBf
`protect END_PROTECTED
