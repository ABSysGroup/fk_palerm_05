`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dtNjlw9WzoUSpJIL8fnLZf6J3fQdHf2dG84hrZJFEzOweMTqEbjEAQ01usSATcQ1
n77BTxLXPNh7ZPI2scfrgm2VGOwiKTJzJVzcCIuVWgzHoov+DurNQp571Jx4UxPT
/5WMmUMKrZ3pPBvYnmMDNzs2pSI3GqdnZCvaftRN6capeU4XN1FRg6BgFFeThohw
2bfP0gDGpqy17QBNNvgcHo/k2V7w9EIL64y7pUgFSaF3svf4Vjv7l30Gun5pay/4
yAxZWkQ1gqc+C5EU+U/w9bcEQ/2iwxnzCR5p5Hp5UzpcJX16mbiXyu6S+mNJeSEJ
INPiyduZmcLS9orce9ho03DF4DBDeYsr3gJMor4aXl4LY0joSP8NzbTba8XuqmKW
bAFzS+Il6gDYfruFj1WbFmvfXZsLsK8nnV7Hrxj7OOynwVIh4hMN2JvuP+mjCWqK
tac9gBQDPEL1Jj7gf+wb8BFhJQCfPrMvBTTHvGRtTR33sDCG0lB3nAl4ztYzfxZW
rR0DoNjNSQYEsCUETf6Y3LxVtOveiG2TZGQwGkjysftlOY0lMrDnYLXO6r9m/S1k
LBkola1ynPCozaQUAnFRFHGU5Kovz98V993bCrPAtAaOrATDvGioIlGP5MwrqNzt
73bN+6TJ2K39rPRyCf6AHCI8Jx6qPecXIjEriiANp0lx0xF37qz0KlLYoKm+F8E7
HOzjA8imohBMemy9V6e5dNmiI5FaC98hilhvZZMtrSh2cK+LourkFEBKDtDfFcIU
hvwnznaYlCsaPY7bI2JIV+/C93483AR5BxXNbApYzAmXsKEdTCTiv/D4LFGnU56g
forJthmWhfko8sBAHyMfj01K0cZjvxjnccdV5Y8slIjGJLlLOprsdQNKNPUmoza4
369LxueNoCZ75vSmgX+RjK2UlyiBK0bSItouUGJmb+C5y5Y0y+y8L2AqxwD8iyxw
bVcOtwrg3577AVxlRFHphdoKFKwc0OxqqtD/yz3xq46WIvnJIQ7STt5B+PkTG7e9
GijfeDt6bzJXURP+R8v0XWspuAXk94SGCg+RM2cxHsRh2mjNWrmlZkN2uA46uyKo
7O4USOTPf1QwnRnINmVB6jZDLT9WoQRJB05S5mlWBE9EaNLRP2v6TawnRVQ1Tju1
CtjQyshFFVP9/ztcroQj3VZL1Mk4fsgnkvPuHpl1u5HjMf4mWvPdQKQ3IAkscqGh
W8gAiUJzwL9HCUL2swJGYvrn3q8RtGLe0FUlC2Z2LUFKKPNYXGNBplC6mjNIB/FO
HanGtKKgQrt1Ct+TsS4KnId7bkTKDcmeZHReXf9sZXkr7q8IM5gTzJb1OIwIF6aO
WPFaz6kQrmSAS5nWgSKeFEUkXgmG9hlKNbuVpv0mX0QDqoqniuuu4HgN/Eu8OjzX
TrmRI9wvSE7qMpytFAIzeh944N0nOVhnoO9tC9dW+HWn/bRT3EcnSbQtU7IHaGTw
byFEl1avd6yxTsMQaHjORBjDJZWTdPO5fS/dis7pJFz53oEo0ZR1KXE7tnkjPTgD
cLFVFl2t0uAxM/yS9eNQQ9EKmYG23ZLgsCyPTa8I5au28Jg5lc1eLblHPBIb4u5g
sMdEhMXLKF8pxRI/70L7PxCc9pwmLq0IM8gv0AdYN817mJeFTwAAswAHRbtfXFF/
oLj2UPBoCHjcEhBxUB284orm/TJ4OKmvi2AQBdJPDHdHQF2nWBzW/wSNethzGGNd
NsWrKzpoF15wzHLBmMKf/sLuidZMejGBEGmJ+dsCalm+5OAHh0jcWRsQkghh+KTg
`protect END_PROTECTED
