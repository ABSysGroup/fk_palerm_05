`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JMo5cggWunZfvnCK/7/1//APRIUSYE2c+h3ToB3eRGJe33zmJ8mWVW1yK36P9VRC
JAugkhttaWvCkPc/v40P5yv9yEPqw4eUUWO8zT5tiLLaGS+Wi/dRwiphyxe0oz6d
ecoSmRs9ohdPlwh9uxBuJVSyu9EMaGL0k8jUkXHeKaoiNyI9UMGX0LXqcg3kujfC
k1rn4OMC+EJOdQYv6DLmsLxGpAfDP549S90VGoVzW37P9WN55qwSOUk3VhEDfZZh
maLdDvzYSLsLr9CzstqB9hw2sfEoP6+eMXoQdAiYL12qKsRdhVokQpo94sEPpBob
7v75M3pqkOpnLN2+bECFrs0LrMB8Acfk28YtWwZd0mxuZlUH4xa4hKYpdEMWLX4a
A83BGLloZWVF89YIQNnfvkgentzLU9LJylJ8MRYzw8aHNvyLdMQyY4utYsNfwBiC
PBLt5NNzsHpC+O5GKErp4p5QAl26HGuUPMXuV9NTiSY7mJw4lVoCU1Am6uQlXjsO
adLRbi6D3ve70h2lIs1Xvej0zw2gTwYdNrK4fMlBjvT6BdKXCvWKrtVsza3BhZ5Q
HclyPyxylzwCr120l7LP+Ooi8r2ZVhRelvhP839zMSfszJnjy0RFFwlPWMewa1xe
vjqB+xI/q057yokl+rxvNg==
`protect END_PROTECTED
