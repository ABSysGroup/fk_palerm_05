`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OYXFuonem3Af+lWQ5N9yHqtJjgYUlrq974x30FHOzASAHwXOfKRyLb6eHN81yxjw
bMcm1gGTOHoAbJrt73Ezqvy2vzkEOcKQdyYNAziBHhDgwSyfYoBJK5pKSRXWdiMZ
SBnvXfI1sSaQqw4977Dm0+OllzlM9Kpy77olYz+BSoAVgPZRH7e3wO9WNbLRp2ns
C2XeVKY1nq502ctnf1fqWjdEwKUmYhYwnbezoArVe1CAfQ31CR8t7hMaGGN6MftT
MWPEBr94ChlNXtMsMXUPSgJfuoZqtPoGAWm0kIg8LpjgUOXc4X64K4E7i6mflVfR
IQvleX/pMZIZ4Mf786UjG7L1zTRgY/2GNq692ZWQyA74F2kSZitDGgZQA4ZsqmQW
LpYbeB5XIVCMfmq902lWcIVzrsKDNtsW0YAbmtts8AUskUzrE4XfWB6wIgJCwBKg
faIwrmedgfe1gsUacvGXjqfVQvGG67iwOBTTYqahzEDGipTAu4cUkQ1Ww042fany
x4lyDXEgKPNE/MwqC1+iDDGS7wNd/9JvnnYqbiAy3jI=
`protect END_PROTECTED
