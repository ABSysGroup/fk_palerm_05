`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wD8OhAolXLLUKaZ/If8sF5eVECY3qw7ZP9yMczx9IklAOhEpYnpv22Ww41KyBfBg
XVatI3M9FmTFTVl5N9w6sdMGjKWcRXHMbWWYhNgLX/y2LdTY72jHkZ10yTCT/WC5
nf/MfisdbCRM+pFCRJyt31a7UaT4Ky9PbUT9HShUojgpXq38VXK7Ml7OnYAlNVd1
x9PqTc1SeZ+3GGv5UeILoS7PhPqBqE7hlsaGTqw/YyQzcCaFaHoBSeUmGYU97d5o
fGfSiwATtaXDs4bNQIU7Bbs2Nf9pk8qFYv5Wuy49xanTCHnmkVONMBuFXJgnXJQv
rLGlBfVfjes4OxbSoqTunNh0iiVnogqjV8OkHiNJK5g9zP+aIcaFRhdSPYBri6H8
pHHbx+lWG2vcGY6/SceUHHw0O9eLx4xR05RSbGxM1Qe2+yIz8yYSYNdbj3M3XZQi
Vymd8JEOO7Qt01pWZcF3jekPceY5eZCQrDOvrPMW1rsL30URsA2dbQmDI+V5HDm7
hhbWeZ75UXPBBGsLOZSbjndD+Yu7hfcBtVD+Ga8RdJwVgbulGnvgrj5a6XVQiufu
MQCWCrSomvt469thF9TXC6deoT10MJum5j1HfxR4EPqTtTe6WdKV44U0/edA/psa
jkYyXxuYc74lTWLUted37PHMrlqmBa70g5cw6Jelmn24hKbrH67Sa8qKKmtO9tkl
2wHXNZ1PYio9lToMuyVEF+wrtccUdepxqfqzJOQCYgg=
`protect END_PROTECTED
