`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V1v5RMqTr7Z9LR8xk8RxUJU1lREyh3eh8wdqbCYRO39f7ucG/T+H2FHtkJcvNSLo
eMYtmSi7Ovoh46t4giKPIttkOLCa1Wsy/lhy3yeYti9GTwbUJJlQFL8A1xjEgkRm
mj5N7G5d1eO32y5Qm/OO4/v8dZLIQuxqjnwoXz1aX6eLAhjA6EjMQPBjEjTHh+t+
iekK932FDzC9MJNCEQRLfOjVf6ufus1yAKamqwPDyRagnYq6KVTCLyvZx/A4otVr
/qGwn+Gv6ltG6U/o4Gr9o9DCtPQuVSxxriIJnqUkZXVMKSJEL+BQzUNHFwVloza/
6ewboLz0ulDToa5YLrNWSzzdhHRQMokP9wdH5S/byeWJl36wmXrARvdGNAw1780q
`protect END_PROTECTED
