`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fGZzyglA19Bs3x/7kkT3YPH6/YNlOjWeESF+QhxsHXLfJfVFEHXP27XPxRWWBUqq
1IUzYHIK26It5Us/bMB6a0mHwtC6H43cRG4hrZpfKylARsHwk/VsyJ/8z7MAmwCl
TWktt5iYmHzD/98VKSb/thdKw33/832rRb4XBsov67s+fZ9W+haLnuJm76KV0TkX
tGU4699hOaSY5AgCf3OLzCozAyygxSgeZILqIAWQRQmWFBN0V5oAL9E3tNdrj1ac
`protect END_PROTECTED
