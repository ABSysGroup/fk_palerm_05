`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IFcUax4X9nRUEwp0cxyq/9fWk9IEVJSzzSvG9yYSw1/gWGS83alKVVJSQsGUOHy6
Sjujyn+JOl3CppMQyvI1srRDVwZXVPVoNVNUCU79KSPch3nnGf1/2RSY2K5pwcJ6
yzazOqjqSc0MyzNfXFj7gFTw7VAWlm0B3LMaqk+nfErZoZ1lUZWnlcMyQBAU3RV3
+CD63QOo2zy+DAZqHz43S5GILyR9VvIdTLkzxyEXOH9LBiM0kWKqoOg6x5CL8Gt9
a2KQpZVoZPQkc8hw4XE+w9z4DzNGMAi+xJXFK7j3q+Agm3iEvSGa7wpGxaPrL2QI
fTcAmq77rvPTN5vmCblpz5nqKNKEoNnF5hXmiDxwP2Q1zNb/Y/94vEVfPeke2sJp
uIeZ3MFOjjpbHROFOF0JefL6XXKevdo3KFd50CEZGdTI8XekSphhSrecQn+ksykd
IQQUOSiGY/O3IR1SrVOBzpvaJrIpn1kMK0/4H0JaxW95fJ38MroFJItBUyOqnvzp
jG2N7SAVEEwejA7g84g6eagjhOnb0t3TR72VWiGqfhR5QH0sJjXcZKdaYcJJL5Gc
bxeh3he/LpZtEvzirv015puwbWKIMXLacpgQHgyDFtU8488gbbm/Mi0PUFW9uyJv
spN/SrEiF/CnyUmQ8bYX9uujl5KNsDiKNzj2yQnHNOXZ9B0aNzwFhXlG1CYffUE6
Y5p9jjtQN4TPEdzSz7Lk3xOXEg/rqiN3TGWqlGy6oUfh7SV1t6VoCx9lDJj2O5FO
Ns9Ax9wDqd0o/rzh4w7QCXJdwudeNwK3AS8i3ni6/qBxXxqsH8XgbgujAANn+wOf
WtbvoQ4EeTnm3e0zqHnxNp/9xS9p80ARdlv4vPMYmXARFepKFb1UPXxhT3sSIc7j
5jhYN3Nz+spCxlWPh/oKINaTISfRvaZMabJbgvttPNAM6p5+L8XxOTm6jlnOiJcD
b3/a9FGNtWY4JH0zSHdhC2yObRHvM+GPr1A9LZ6rGWiGqJ9LJmMF/Ybsz2cTJO24
KXAcCOGhWpsCLGL7KPGkq5vPFTJ+v1fPINZCdZcNsQYNqDRg2LIraaaxMq9KHjE7
9Ey46S0enFQd7f7xMvttkG5WPM31FXxG1UzPTRl7K0EvKT+435sCS0MiggmraVDE
k4UpvkWaAgRQW+0dnXBmKqdValfbI6ect3jAELzn4nosteVZy0sbu4WE1o3H2L1U
ZknH57Bg5lgjOHoN6N5twux2qTDZCVB5tKAj6m5BYIhQ3iO5U18VZYIu0GUp4d8s
+2Fbzx16vp5rYm5zvndQ5JYGOfz6ugj5RsJmXknzN8I7lWuznfZTvWrdoFyU62cj
/6QpZGULWv2AwRELCuBsQ11aJaRQuZziQ+dZPRn2ScBUn703tJGt1ffkGiYJIU2O
73TinOC8mtoqi02y4HP3x+M58J2rHvFafvmPzlYDqoJojPvUu94YX9d4UOPZb6Ty
XH5C6SKf2MB6xo0olCNIO/FT9Rj0+F0HX3hETuXcSYFvGIi3HsDYIh81r2v+RsTC
/WfS5pqcKxTmH2XPGDFEhhRbcmk3e+ypzD9E3s4YzjdgEa6KlPmf5tqg1aej4ph/
vOKaeTrB+FIhssFbd1AOTWZglECRt5GE6UPtkwEc5LxxphGRJHMUXgarC02I3vCG
H1YwjxTr+W+jdCyamDpB4rj1i94qOtuSh9uYwo0P/x+/Hhr1ofDhwU9Hq/AoyILL
O1CGeomp0p7TtpygB3saTw==
`protect END_PROTECTED
