`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MlpPQN9A9gsLZxLKcuttFh17Nno/ZGyQjOKv0o7Yiw3Vt0SOh18Z8DQfTQUPkufH
lgdIsHKST/nYtMrO+RckMs3D+Y1qZUAGe41O1v7IW2zvVNbW6xE0izQmg4bQDHR2
9g3KnJ+X/3iTCsWcgzWZgnrNFrRVOSfqilv2s+mQg0LzsU5lqiUO/TTyly8ESVJk
0vl/AfYzE7wL+Bbp7fUU6aASxMFuNBeeAhbHewQII44HqdzmAeiLLMM5ULGO5C8Q
SebzF25EGYxqpo5pgslSP4KFbGM0hhLqummZXiuMf5dSNOli2+ub3d/k9BFP8l59
dX29PuYQDCOsZsye10aR/mB3HwIHnfJSBlPabhTWMhAquZfxx2vwegIQ+FiIdNTg
NGmSAoDyIiawQ/oAJwrlNu041dvfwyg+mjVeEn4FcidrVt/bFRvE+x/oWRUBLTSz
y+qdNj/1k0Huh+bBAHp3duArHY4pP1Ucaih1kDj3YSTM8q7ov0J2zhADF8cXnpkU
c7VEt4bm+LpF/XKB80CYQebeb6LZygwsZiu9FWwrgL+eeuXQAA17D4osxYaMfbvw
g+9b5RcFg491A+0Qi6j0ZDJbv4WlLWoIG4tMbykx4yLcRlrzxQ44WtgDW9BnZPI9
ahsOuPWdLszQvgSIdQ2hXw==
`protect END_PROTECTED
