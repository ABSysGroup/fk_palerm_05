`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
StEA1bOCgBsVK6+3yVKQ25Qyg8ivxTh+Wfp12rT/j8Lt6yIm3XMmoGraMVOAo90L
rirNAiKuaIBRpoWOxLS/v33N1Y2b+ay5t6+BPD0FmxCeXaTZ2cONvbueLEehAzVb
ESAdlB9Pfos82kBms5YaB6pcOs+r/wZHKnF/rY4t7cs4LQ8Wx9B6RaelWluLUt4c
xesTSExjqaHVHhH4pl1KzKDfF2lP9ps1KMGoc9eDHC19o2KiJFsZ/SK7ZRFVxePu
2p5Vtt2lATQh+sWpIjGrvbL73NjOmqlNSrNR+vQEnfPvnRsqjG09zW3W6AFZnaZv
PlrUG40Dur1uEGpf2UEKag==
`protect END_PROTECTED
