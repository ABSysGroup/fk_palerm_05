`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TH3Um948f2XYG6HGaMHHi/XVRL1qIFP85IOoo1LT7Yb/F9jn+esg43Q6s4Q2VZxC
oYeP1zMaIy7HN2n6ptO3xuI7TYTEDbuxFhPJiC72REulPHaJFNL7ON+FOsUA/60l
oe77fBCYujgHQUOMm8naxjxPpLk+POTC2D4nC2deFM1pteEk/sS8KVdNMyHiwt2e
siFHtwY48WYG7/aWMHPeg1nqF41KTR/5WxqY0YxEWa2n4flZJhihI+FV7nMYDnMu
+aCzkdqOneG7OkW4qH10TCRdHUWOS80ZgIKjWsYuksxEyGkAINQ71HtxxOB+12mD
YvOX2s3WLttXGxJxAsxkfa6EktP70yTGaiDi+pnVW20ZGXNiI0GXzhGRP+xwXmPc
rvdqQfqMBqiuqncnIaf71L5l2sE0mW3vwS1IminY16fxHkcyTYQvUiTzEQZcyFib
blVFhEI9k9MUZ9A+KV+y3/I8b2NEhv95E09Ogg0C1wsVj5hNA8YsIF9fQcDTbp37
rHkNqw6pOEm9sllcCTA4ugPYpK8kmbXwvO27+WUbGEeHZryS/c2dri9foSu3EvYp
lYrO2FdEwVPfJKDeNBmiFkYj2aTQVQB0EOm2mYSfT+JSK4QZwlUrQfk/2jNnj2Gm
gy27UpgOvHk0JUhEhvRoWQ==
`protect END_PROTECTED
