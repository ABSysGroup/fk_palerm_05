`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3SO9DL0PgoMS73wHn0Wc2RDdZAXsLHWcS0DkMTM0B5QJjq4BUbNOM7fKFTmXzgSG
ZHMLuwoWWSrwK3he6l4vG+HitiCM2GLwlpN8WXsMjXoMQhIk2ljVj8+vYJzGB7k5
AQ+9UwXUs+Kq2DOBObo7OpzHBZo61VWyy8n1E4N8qYzS8fGJxEXjIMLO3yb4SNCH
FWFQ3ytLSMPNMxEvWiqsE2L8mcpoQo4hKpuruFk4gZifY3k0O7LCrTbMdHqdvp4d
+ueXyCOL9T82IclN1MyurBEca68vGKDHOA5qEJF3wt/VufMMEAQtio+WfYf0iyxw
7thWAIzL8avoLGaHWCiTb8xHM+him8xdTPlDTR1fUMXbQSNsdtL+nQbRDPWfStj0
jF95SmjzQLuwIgGZoZGRFcg8weedXjk7qFw790GiaHKzwnV9s+tmzkuz3qaezacJ
cN/13aaQCZBJau+9XZlgMwPwChD6LaLkFoAHY6vXa+RqzSnIi0H6mUU+XsG8IG/p
a9AVYWy464h+kC+QW5/WlBBSkrPB1y805GYyw74tGPdurNmPQESmlzz8IOlx3KRg
hjHadmx7OK1W/hKAIL4DPjdMHb1tPv9STj37gr/F16ahxH1KoCJYeaE9kEBB04V7
fII98PkV957qdHJsV6FN0UmDfKJHDyjNtsLfDZif0/pPBwyRYW0Y9kXk453Siazx
`protect END_PROTECTED
