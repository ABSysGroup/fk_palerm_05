`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mSx7Zky5hJIXlekP/jzIaRlx1P6R4kWEDI4QWGfl1bpEbOGloXYvv/UcM5n+aVxH
ypkt7gZUY8ctBqYMHmVdLHBn9+zqzbyYOV8TN/lZu3Uvn+FULjYPPNXQG/L5XMck
lxquS53alQ6Odi1GGE9CgWA/sllYU7G0oyeeaK3sr7CDTWOaQjycNyds4HFiV+0N
Iuk3H6pKU0pDmQNXv9r2jJrnoFkFSvwEclRH/M37MWg+wi7S8wssRRJfShTofVQh
tjh6E88YY+5Q9MJVmIIogruPIDDN8TOYv0UHDocuamvm6uGvINk1wtI8Jdm3/E1+
pK7F+YfrFobw0vvis6x9h3JqFDKDG/TIxrxs9qjBBtpJFhoT8w/s3RGW76BzZCLY
DixBga9a368sYDsYjuCR2h9bFT2VnjU+9GGmVbwxskqMenY9//2N9hfiKrfhP2tN
vrWQbq+C5w3NymIK9LEZnl7f6SMiEoh2jGTnr0ZVCayWKM+qoxIdL8CmksqWV0Ti
ffvtBcHN4CSVn62lQ2VM4VL6HZGnOmimuiTte7GJaSjl/qGHESHGoUKI2dpDpbx2
iKR+EbUr1N5BTgkth3O8P0LWoIeKmUb+Xbe/3ly3qedEVsHa5ngEeiIoPLjFGU9J
Xq9iwYRBxY9sW4c2bS/9Qp5VIFHgy1Huvz2C5jAasq8AzsNYfrW3TNwC7qGdiGcL
+jxVpkQT3/3+Cqdk1o0bqfGCPk4llV6MW3VDThfqba/eAxaYj4VhHTRLhvWgYgWJ
xT0u7y0mKHDERxrdmfnUHg==
`protect END_PROTECTED
