`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eWUXfgTlkdTAz1mHKPcjzAFd/cpVWrqRi/JiuAQ/udrbh3emT/UOkctIeb0IPAr3
gko0mi8xiE9cpZqAe4riD6qzQNVK93Ah09/IOiURfmDJ5lTBk4NLmrT7YKUadcyr
O3NSnBrAj0brJ7i61bwHxSkA4WknpLwpil929pxeDFO1ozR7N4AzUJak3uSTPCBR
Wm7/TEOTpncHxDkd8k7TeImQ8yl7fyk/BFP1e4AlCA38Mu2BX8zWE0X4PR+9JJAe
WMuSi2JIhZxgQ752ZBaqk8xOzwpkuwvPYbOigKbkZjwin1Mm430a8YrK0PGTN+Ud
eW1P0tXEHJlaPbJ/pRaQpCwGG9fjQ/dR5u8vtZ2/3gG7aHK02nKRIfXwyhyPXRYg
/mqVpmQ71B/LsQPdkjP3Wx6mXaVd//yGFdF7tZoqLQH1xZy2d/cDSgUpKBUoPWme
MCiqMFmOrq2LuDnopM+np2lufS3cVMgy7GsUVUrzQA/7xflmamUHRzd3Vk0F9BS6
QWvFDV5FS2vmJVMffIgD+zmcbIWTg+LGozW0H7PG1Yy51lCJKpnuwj0Ij3GGizo7
ION8F7+FzWc/Yu9ER1StqwBHC/FmBkhmgG/eMR+w3KqHG/i8mYQMwvsFRRq3l07Q
QYpYoYWk+MH/tiH1J1TURlPJPHxaYxctneVh7O3Pvlm6psxEKTKCkwnN065NNs1D
Py++zCSTwVWicz7aeuyS10qLJtcMRNPC5rBg4UTlTHIP/asA+qEWX0UZ5U0CFAFG
w4m5Fg9OmRSeVixcH3ugCQ==
`protect END_PROTECTED
