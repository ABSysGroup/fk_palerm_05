`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LfovRb9OPJHj+79Fs4YwW407tVhEKWDPR6cxCQNvJs2P71cOB6UYvPyqG7c2zsSh
yt5cMR0SZJ0yk7/zE8VHzhmPyASifZiG7/pb4iCWHsMJNEGxRpRA+xXhDOONugue
1lMTCvxgSRdN5yl6hnu3l11k9l4V75TX6TbylMS16zYIwFIGp7Ye+QDXXd/z5cDI
TDEya+8/n3zOjkm+JOkc7jxrdBByTKnT0BYjNpFpP8nr+A1i9A6iFy0XqBigWiFi
2uslGhIejom85TttGtD7sWaRort2ZjgNaTPJe/nh1yE4pRkvUPAVcbcIqw72f9Tb
8I4gfTc+9Si6LbSf1NyHhuOcmBY+Wa/RKjQP2yXsoBQze8R1z3pGfXb6BEApWJKH
ILfWuzit/NgggF5DCrmeg7YLtESLmXRTM6Co7qcc9QNnFsBe6B7/lkErjTXEebdG
Ss4wHZe+nM6xaVHI9Ly9i8Ln3YCDmk6uR7Ki0iGSvFqOyzCt9w4n1thms/jxdma8
kzyZZ+z8isnnOsQW7Z7GVHCCWUTecRa7QqSIw/+hc3C31NqsxePX/BP80vmrYRL1
naWfijwFIur0WWySUC3u3Hbx2s4X2Lrf59j92Jz55nw4oYBNZRzJ55ImDzNi5D2g
qKOniByQWjDqZ8hLESikl8TroCKlzIrvYMEd9gIxA/htQtLEeu+MgWCdHA/O/+q6
HxA0CSTAP6OsKfDUcnAeHL3pbvfWtmU1mGnu8gfZP6vbQg4uKM13ez4bNQfQGOeU
A9TeZpvqtLFdivCfkiuy80QPCvrr8KlT+FvxCwjQeQFPTLpUge9i+yuL8ZmSz1cG
E42/zlBslUNK7rB8LpOvXnqqLTPjHnpzbO2Yxr3F9sEwQ6jIx4OzBmeu8uYQPLbT
3wD7fiefFf0fEQ93W+6RDuekTUK//v0w8RaNXsUYSTuC2YKjnrwFNdh7azhyOfTa
D8Bp8QzKumUOUZbZ7aAtFJblf97xqnJyxbns/nBHOiog6MltOVMoVfm6vchwSk6N
hQyPs2tacGfN5bOKS8jqxpY23QIbhnAEL+F+RL7R/47r7+R2GmPR39k13dDJF1Jl
xz1GhJSXFilWzF0mr33mJTTWuIfCOvJg3iqX/2SzZarRvTIy6OdSQAQpAO8T6i+6
DPfTYsp7v1rB+ALxJd0gVn9CGDGesgD00qTx29IGDN0SN+4t9rSRgqbrCDKieXlS
vPaZk6aTceAM/FfOgGysMMA84zobEwjToYYnAk8zmjnVIaYbAkbXdv9rEoReFTgo
x8ZkR3rBUI/qpB9EOQZmxrh95yERa5x0HnHR+4A7RLlJUBQFjmR7NwMQnIdJeoVc
mjrJJHGxOb9gpaoXpvw1W42S9UsMVaWwbmiGYJmX//xEnpC5Haa3VaK8stofPvI/
bPHT5GJR022FhE2NpMn7NiCk0kjQMWW1ycmBLhz8AHgijjZ5Y/aa0mA9Je1Nt7no
fZDdlwg+je1JRx6rCIU3f3IohjYLQ9yYw+yKO4BQJNA0wK80ZIkrPwHCIMeT6Brr
eqi46gVSoUazFVoTabot2eKR5Zy9SSPy97UDUN5uekNWjoAahifeRjKNZdN/UsZN
S3p3/YGgzqYBbMMO0CvpsS5PvwJoTfH7D0q5F9AyJxlvl5frwRI9g8WaR1ou8esH
xLcBD58o45cJ3JQl0JEP6oaRkDKPbQcYr+rUWNfd20KCGmAChXLpxn1oVjZ4bL/S
t2aO37603cmfTGIb5JEv0Wt+OPOWs0NuOrHSW3QKnIMXc+LMZl39AAkQMF2AhW8w
3TyFvf8cBrFYb4ahWdWmcw0VOJeymY0vfVFU2xMvJU70eJC7KiPz2hLpEklC6luv
+qJn2eAcROBkxBVBf7q8rTwyTaWelNf8IictZCAt3XOa7RkDjwLOrez0mi+jXuFJ
nY8lahelWb+eUBY77l+rBM4naPLG9Oj7DtwvJrLvrSnRZpOa6zTWHhNB6YqM8Bcs
PF9ZKxucCmKWaMQg/yzI+HlXJLDXuTcmqQTiO1PtHbYXfmeFR4zIahK/33ivxI4Y
awEe0bHvG6iQQgTmoc/9MqfQUw8LP2tn9USdknMxuwQX5C5X8NRqFtcFSxMiTl4l
fXAQk+l2FdjwV6TNGN2o1vYITghsTzS9tVrwV+eZqI6NtAhV1rO5Som9Sj/jBzMU
oPG2KbezFYVWL1ogEoulYmVgMBxFrT2P1T5Gpafr+Z0SkYMQz1TpCwDUNIskxTeD
NVJQF7v/eRcBx3n9SQCfLqghz5rBQZgD/JDhUeWpXIT9qdT82a6AoVsNE7DDgJYZ
AtlcRwSNNyL/FO9IBImNw0ZIEL8o3BmzSyZoh5trsAbI+/sApqwHSYsEwG1LDijI
X02au6co6pbkWNUV6fe7IUPhuVom8Oikq8rOC357zX9y/TRM/In0+2vzm3r8rju5
rYnTpI0i3tGZmQoobo1FYMTTlOKABDKBRcYcDs7/Y801yAT1HiiBQtputzzbyd3Y
Ky3hZfbLUCJuy2DqqkHqQaLbzT1ieWick+YQoSTLOfnOXHnEp3lN1l9PAFM87zqp
EziDTBBOLkQ8FZ9vNwo3/BL8hC2iDyUsFhH7mNjQSPeUgSQCt0fIWN/XHBGhhWJX
r/7kzn4zxp4pOG0CGjrYFlxcmYZXvCL1XvnRSmmFr4okSMzSuPXm/VAAdtIdPTLx
qKNvIMPEur/oSYncWH1KSEj5VsJeTw5KNI5AWfahnrIy6qF7r+aRC2xCPxc6HkVv
BH+gwtzT5m2kpPA/dE3w3G4uLhfcj5FCRRLBrfzE8pPcxxa1dodpQ2CHzpFyCNIV
cT0oLNS7McnzCxkaSrfBw8iIDEk4MH9FE5ww0kYyOgWV+ci7FtZDufjkwxbac+xG
VdpA+MNV7UYeBk9ZOq3DYz5KJYOy30Ik6LuFjS03JnRji1QJ74i1CnJd/Omnn3uH
elNOAYohraptR0OMfsiSH/AHTHoEiFnibN0cPJ2DafZg4cjlFfteHerZMgTbGQW3
V6cN6xow6efnB/yQjUX75eKvt5NjpOTTGZ4A0eJc2aZUNuBtsQSzHZH+rJe1clgV
nVI7C9L+DM3MrK6d16R9wx8iJ6MIg2cCMLhAHJyW3Ds2F9qScvWHXmkwoF7Qc0Cy
XKchd1EZsxK152Temh/iIO8QB4b5Q4OzHO0LGvdFRqSa3j9/Ls51qrleN68xBxTD
iGU0q+sdjeObWEwRY5WeQw1BANLVuhh3OwKyB8uwrdsoEiM7x9DrjM4miA4p3tO4
S1n9lDZE7tgviIdcycLtyd6Zeg2c0X5LvGQk53AqaRl1c57V3RUApjuftLHLqPc/
Vw3FKG0BiVQToyRT28mwP/8LYDVjLHzn2gxZOCYkZY8S2dWG/DzLf3+FUeOKSvX8
su8oDqCQUzTTk9aKHUkepUOf+fHcjpeKIKXKCPMYK+wicNAOAInpQNgZrdu9NDDX
XW6eAUnRakyE4mh3JV/SdLUmOSoTqnITvrUaouUaMYRGGNqjIldxMXbbrYkR5RL5
HJwWTi4U2Y2pSfB2IlMoHWEzYzl6+YGL4FsuJ5lwQholzDQzZtYU8cAK/e5TRMxv
cVqWl1H71+qmt66tabX+RA==
`protect END_PROTECTED
