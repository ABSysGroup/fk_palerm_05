`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eiFJYi/DfIX9/FtRuu28isrFdXkjhAQU/Xiyw/oWA7Ak2po1bWC7W7tgr2oK2BBy
mwh+rp1unB0vKEnEQo70tkFzR4UagXFpTlW/36QiOHFRVFPPcRXI+nhHnalzG5PW
ucTZk3ITofyQ4Ao+VFVPrzaQgy6i0MQS9yghXHFcT1amrGBC6yGoTv0qA1mMR0zg
KxZIXsIbLXNyIT+Kixl7kDXYP6z8J4Is/uu03gu9vTRLT5i3V54/XaZNaSS0F2Z3
Gvk61DpuVk2qa1aOVwowfD4D37/XMjbLIYrUQ+0avI1AkyIduBH5+gYBw5SkMQl3
H0D9RzIreDx86kcJhagRqfZwgjDUpp+Bzl/Gj5Q/QhijrmojDouHO0tNzBTx0dAS
nD2skKZ+Q6VBD4GCY4//+DG4o0Lk7vQEebHXiMq5oVEKShjuLPQlkTZKF37h2jOu
3BjKDY1cqPV+Xm6ksGbwe8N0/8OVsdqecoI73f9lveh63WBNt1MqvrVKiIBs59vt
7lgA1OXht3CXb9qqWwJxHyw1TJKcLPd5BntanMg4hh5RQpwgub6wZ0ORX2YparK1
I0X7V0PwJIj01cSPHc+OWV47re1N6Uy32L5IER+D6UHw9NSI198+WUWqCZXdLx9J
jEuTu0BGR+u2w8bSKDkfL+Nzl2dzg4cSdTy8JDLK3mn9M2Vo+CWvvUImUrPUfI/n
BzkVafzhHKg8W8ycfoZkue8iGzA0iJXCEICtB1vYck6KPrHYWLkQg9EKj86Xm33U
vhZrq7N3Wbxg7s5H1r0M1KeAzgeQ/WdsHYvNy7ow9S6utX/Kvo1Ko/Ra9wxZW1vy
b2FIDok1dvfCWRadAhZSmEB/S4oVQioYPkmkP7XELlqEpRBL8EvKVm5ipExDAE7F
DNhOrIPqaN3rl5BRhzyayw9dcL5lKjqbtPwyOPh34oPt4QqBDJm1K/8o50AynvVY
Yrz/wpNRwHbHzWNScywQFbLc7Iu+NkkwCIOt0Ckh/wQ04po9xvXnNZk2Y/GZBP+w
/UUthnFrMoAUZIoHSUYAhMijrIbpD5M4NtJe0BT+t/g=
`protect END_PROTECTED
