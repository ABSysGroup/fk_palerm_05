`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m3qbXHutFtvh+1f/oZEVbfgJi7E2OqYmAyRalsxI5LVnlQZ2dQSAxZZSkXMz2nGK
b8IyMTs20E3YfO4b9EbEoSO2SCmakW/Hj97YTQOujzlSXrh5wajzK2nparhvWq3n
K7aBlTjVMi30ILdQts7R+olbWiBA9ruc2Szyh91Ku5Gv7DR3tuM+Rnu4tjD/SoSy
8DO8s9dnhDAybvmMiSbYd7umHDm1lEztfYLelM7ZVDcktFv7m6vurL7AlrFi3JXA
N6QT2E03wzJUim/sbrytKIhT9StnsSBlM8kCO6SNnVqbD2Xj+YgmLpzemPTgHfyI
+PSv6w7uLXwZpa7KZPBODUUqafePbVC8Gf/P+ArKa5WvPGq2vVLOZ1TuErU4ncdN
z6vRPsFKi3vrwh2wnObKFAfOFElPvMqx93ZjfhDFzX/IP8TGy+IrAJOPjBUyJ6bI
Asf4dB6srU27jMpUN625fKQbyoyI9MbaTmw84bQOTDRPo+hvaL7mKBYPpN29V1JN
Koy5leDS4MNn/5yP6K3p/A0JKUKd8E2whwBwNLTDPwt/0eHOAJctt6u/A3P3I0IQ
ua2NjC0AP2JPh5xgovB4Ane2yfxwAczbK8GBDsKg6t7yLST3qcqzlBVlz/YmpFoB
rotD92k1Zjp9V1hjyVzeSSem283xy6vwO/qnt7e5ZFN6evMWtRS2xlIrvNBwTyDE
yAqEZAC+3lz5zkD8eQeYbpAEV1CBl1qeVHpdeXS4WZUJ7VChYjlyBPMPv3IoFJrB
EAvuCcm5DbkuPWsA6MDnmBLgeW8QViPOJ7gN9Z70vZfjZdsj/kl7pQeWBErbuP2+
F0NdOJUX/Hnp/UjTxnjkpfXwAFacCI7s25nsAM5Gn/HcFsnxGtlWFNBgILsbuTgE
e0p6cvp4e9jesS0BYqkKDX9GyZR7fsKrlt0gdNmO25tnDDmNm/+bFIw0JJDESKST
DUQEA+iWm7f+baOwNFLzeMq1pLRIQV0Gilyqme/vW4QPW5IyRAhrSv5y8PnLWTsi
r0doEg1FosMrwjw9vhWZ9uM8/0yDPpEJbOo9Ot9C+D2bAhmCA40iHh0rVGcYV98E
zwrmXPYYqdCWwUxXLZCsvX8oKnKKuc6VcZCKeVFbivnSikMkV0WL1IsTrqdLzsn4
ftxZmcWPSP7D7siS2eCkaWG5TgbpqpaKEgrVDTep+EWGwzWAKpY9BdKNuaa5h76o
XaDSOK7h7uQNWtlwj1DctvAIosW9EXd1xTnPBr2CILE0t68v+MAoja/Y2tcUyyj5
tmZe9a8tBr0MVi52xd3uThkfTgGn0Ij+m1nN91pkavkaXRmmOIP9vbU/8Xrqg7BY
E/5D1k8i7QRagT8apUpEuv9njIue5F+p7vXZroxsuSpRErlNYRZBleDQVVMg/kLh
yjm2K0tolAcUn8+UUTJnb4dRbUvyP+Wbb+OQfRju82KANG30s0BzM5wlzYurkexP
SeAR4gfiXepMDYxbQBJwRyV+LyOQ+lQ//JJYOFjbDRgcAAy3heUd/qkXuS9+dKUK
lhLMmhFf0zCSfUMQaocuG594PzKDRZQgF6MJes4FrI76A26rVsjaGhjXFwtsLd5W
KGI7DTkLCTdso+mubS+d418fH7VO4/WBYmz+2+yATCEaf48X4b+UVyWmVrsoYpsg
ajV6Gx27ylLpLexIy8IDCZADyMw87enfFA33z86VWot9niyv5sCpWpLfkdJj1crP
gz8GbhCK1/nxtugYoCVFb9OE4iBVmzAN+zv3UBm7ck5GmVRBswM/5IK9gK9j52wb
eAWOsqOAec3QrfOmw0sLFZ4Sod44/2PTcfw/w4cH1s3t+n3YFuIcmbyvH+OTLpZC
45p+K7pVEwVl4Vz1NfRxl6w4w6U7rbpS1rWPTW3tN3aHZ505/Y5zZG3EJd0q4xxc
SXaP9YyN2RX6wdoZNOZk4cH0rwJ2+Wl9B+IGbZ9X1SsRt1dAqV4cxQwha9D0gifD
36ACRyU1/Ynb1l5mDDh/Pmd1I1QOSZY8vahHhNtfXDb35k9hjh6uxmSy2O2DRUJ6
TpWhYLkcmYLTd/xMkUfNjTQ4V4f+I3jXq8gYcmCUsQi6EcHAU2CMFXXVPnSEgr8P
X5dSBx//e8xHrpix/Gtn/1hefq0GcjkMukHRxVVSV08=
`protect END_PROTECTED
