`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QlbhM7C+R/oNGlELEcL0PNhYQ4JKvct5CctjRvgxZSA0+fIRFnjlQ4eWa/8ECwaH
KeWo7JeFoiKtEixtO6Ge5NfmnnIPVPxlKU/WH5c+KNWV5fwFKxdD9Hk0ObOQYtYN
f5+PmN7aIC6JF+Y9/dDAZKxvlS/oY5EqO4aiMDzqsLckwSjHcVlQI5GOVPgUKzO6
Zir8LTQ6ssDjK0WXoBBGF7PbVno/mHQ+s2wzuvT0KwOxZaHyCe2H8c9yIvUusMSh
xMtcqjAtR7dDajxNctk2mJyqF5Z0xZ1ZEB+A3KEhUsqhWaxS/uQx7Lq5N4K+nYJf
x0YPsiWuCOVJJZ0u1CSZut5ye/BY29JL/u9F2ImREXr3lUWNL/3KTERTQLZZjDGT
2EHfokSHIwvHYvVqAn92lFLIzyN0Z8h3v6jpwUIhLZYNAasBnnVyExQJyGtapvSX
1WLtEGvv+8GvbR/6aIqoGlQmW8rX/EfrMT/8VIcVtjy2CGt8Lh5XHr9vJvZqIj3J
nzNTIVdWn7Wk3Ee2HYpLFJcwjRn4xVIaaxdk7v7K5i6Ev37oJXokz99e7Rgug15S
tEkayXUMGybiPGj81wkRbzkKuODK3qXbVZKrrvH+oNOroXaSiFc6VPpSov18uT8H
O7ST2d7hLM4JPStTQo0AN2o3mFtpvnhckhfej0SeDZUKazcBMXjaromK1P0DdKd1
MSGifEdyC4YG1GompWoUh8SNS6o1WtH1VrYUFV6SMVK9TIfZ33mFxD1T19CnA5Bm
ZJ6pGYXDs8FtFEpg/D1a2Fi0HVdNtElII79Lqt0CSRY59nQH8SGzTxcRXv08HTBq
RU/mKsPR5KzMKa+zAQoAn/DPOv53s6FRHP3M74gBEgDIxNB3eRCa484mocywPMLj
GJxncATkOtDO2gNoRJHLTY69CylX1PB8kdYlNY/d7MECdeDlURmVytKptpeLX0ew
toMLXAObrw5TSCzED4kbarWvkIyMiyZFkTEk28Hui+1WK44fwzw+BvRht3CkJD8h
cpZj5JjjmEflVAtGjG/cnfaE946SsjKF0iO7c1q8Nyq5drBq1FCXVwCAUPpg4qKh
sCgCbLZ2s6RhwlFSzzOdGc6SLccStjtKVHzjDHCrQonFJUF/WrSvWy+71+IYOiWL
MrcC+EEPGQ4tX/xY5zuu2eOhIEiHuQK2pqTLjFIHQ+c+f5ETmaLV+giUiOYP1nn3
1m1PlfvF9NvU5sZPfmcgQqzFwEI/h2B1oibFf62ybLhmWtiwv9l/t0KabDMrNvM5
n4JofYf5G/7bZQj6HHkBa/Y+75DHmVWWV4sJ9lltd3Dlv8pW3fyimWn8526mzKwB
Qxq0NNGFkdkMEc94G598kYragbqlK7xTbGmtyLEjxexzTU8SM5/0wnIGYqPi4niG
UBhz3zjiqYpctB+5/SW0w2PObRCJLeIxyslywe6/aIGgDI0sOI5348ZnkT/3XyNQ
gohR5TkcRaCzFTPg/nvMbI9MxPAwcKzeF0gtXOCfZlTMjL3ZHHw+GEfjfl3vpZYu
IHUT3b9Jb91xxvrj5orOiFspPju07k2qzkpv+ppSMeHMmmLWaeVQcydXT5efGib2
IcE8fiSPr/BTPFFhYbhG8cQxJkUKV5hijKwGK1uZbvjuLAZq1Jkx7TGK8NR5kGfj
Lop2Zpf2wxtBUSuhgT8GtsUAoHDv180Mcspj2K0QHGDBZNqTHyvyLBEmusjfvrAd
E3OpkjbJfvuWOgwnaUhuySYDxQ5kSO2zh5czYsKydvwcRIA0tYAwNtY2vYtBpLYf
/5DpOLYyMlygTwqXyfhcXhsEeHAQfHeybAjvot2po6jAyEDmJkiuSIspHkRdIAKl
tQ/IxzwWqja+nwjJoLYINw==
`protect END_PROTECTED
