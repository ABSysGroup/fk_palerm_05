`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
giNl1j71sZnYOVfgajffll7l0veICmkL9AYHJE/p4zGLPHW5jKBUlVtFyna9NC8U
Fnpfv80/VMkkF/zL67Yrczc7nm9B9smqXHsmNXIOb6fBjh64K/4/ZyPvglIbqZB8
SX1ZbbQWcwh62BK87GLxJAbmwdaJqCidElFievHTqQK7aG4vaIGAAUGo+DcToJdg
a2immYS67Fps9Nt/6yDMRGEa007CHBYMdd/QHiqwvpBG2HR3ReD+GPWqGW7XxscM
9Vt5YZ1AzYUgUiV9NCKwBhQ/aS+ALJByL+lTE+qYEKVAnFB6RW9F3znzix4ks1jx
HxUlvVBnTtI31p0N0epBuoWSwZ0Di/yECI+4ZG+eYaZUm3rXMFPNXfb0zgojQ6N8
Y3iMCPo2EZaSBwAUY3vH9HfYE6ZZ0g+yFW0ZoVIxIrjY2JnVH5M1RcgAkrAWEeEj
LbqcWQF3bzDRsNqyDjNxp69JOUGTwu/DuSbio61UXIcXuh9nuF3hhrGL/LYC5Lnr
wsxQRMCozescUDC+7dhMBYtVVvHX6jqFVbHz0yvlEN06R+mvnrnCKSK1EEb0pWza
DLMZAJxhSpVt4sIfUw+14Brjg0D5bnL4/rL1CnrLh7dJ1BT4NSyRxb4C4bVqIqXs
W9jRDWuWI7GnQ4gnpt0Xjw==
`protect END_PROTECTED
