`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2wODbzye1q8X9WvaBpLUVwmfQEAcQ38RYIzFt/5ZGH9H9WC4dd/x2ZIR2SuYQosc
bZJgYQsNwlTX3Z3sGuOipuJrtG+nCTlU99JIMIC3Hl1jaWxxFDsxBQ14UPd27bjW
9WlgUsfxGdAMIyMTyQm/0sZYlm9PAGvGy9IoWob3lL5QIB3gRxiOgyfpQITye0tI
7uLMb3nLjgToqfr7Yutxecyc4LgnnV6rRMzQqwXL4c2ta7GThF0KnGvzDsoSPGvd
TLYwRYvvaNcJ6NLur3Tkb+CXQnqOXtTLNoeN59tOPDxOJc/no5rzmWgznS9jsJd8
YvDnkVcIj6PHFijvw3aV8NKO485s1MH1gouLRfHUtDotl7X8fMNJltjfYCWxgCec
Xe7NnuJBOh22iSZG1OiQHZuAG3AWN3M2z5Wn8mkUdEKNIphTJ9bCtz1FipyBSuvE
bRayz87lm4AfrOcLY7RGA9FfqIctHw6xMH/uuByhxODLnul+V9cQ6aCaAHH1zZIV
`protect END_PROTECTED
