`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bEoyXYDE5wnqiawhJcFcm/VYLvAyCLxKiWHQ8kIkgxYqMlISj6W2OLMlRZkCQ3+Q
AbddRAoTkJDpO3ofuD++i2Pdcfa3effn0XAbL2MC5m1abgkChdhlDocFnT+3yXJ+
KYTTAqhdQhGnmfFaZntmEE/poX0jBXWKU3I+fcb2whEoFMlx9VWewl+vfZdrG8/v
gAbFrD86keCiDOmgS1YLKhbhtTr6+b5C2a7QqXBk1jozOUDt8G2RVSho2eIR6yia
UCoWhYR+ZiYM3whL8XOwgxnaQC8sZ10/FRofWWYzS1Bwn+H/oUHV0LwO216gmcKa
hItrPr5Q3ou4PiJFkXmnL1W4YIsAXT2Xe4iIOv/PS0QMcl1hHI/bHri/IkQeLXL6
G96mP5FTJu9OQadbqgiNmglOvSuoLpzmeS4yQEZm7Fs=
`protect END_PROTECTED
