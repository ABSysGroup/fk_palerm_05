`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KqnE4/jZusF8lay+RIFlzoL9EpkCiS/xITeni9AN+1wD8lPnRkivv9QxYQP7zEu0
HQebEhB886aqOrhclB3x7b23btQ8QXvxntHSfGZGVElgAxeif/N6eWi5ggUNSKOn
TdHppa3Hyt6p8bT7fSjnklGM9Len0s/0nueh5pHZNCLEHhmaKnMqloCnaoSP2ajs
F7Js/WXCd4TA8eymtOwo8+bA5d56I6MJCDCOA/jKm9uVNAIUQ8bcMTaAk8A0/oil
XV8ILjh/3dgo7rRYrFZ8SCoukGiF2z1j0PECyr/w/Hi/NqsgxB+pELMlE5S+kjRp
9rfXd74JKULqi6mLDnY1Yq7fjUJSTzyqqUfjmORA3wOvPsVaOM3qDNeD98lKQatU
+QP/DiXE5LYYQpBupJw8T2gKfCbCLqQfrEORL7qQ5p4=
`protect END_PROTECTED
