`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PKRAeSC0i2YxllMBM+CspwOhX09OS+YhgnIs/DcDVdEAZlRwYrgfYyybIdxYXUUe
+UYbRCF6MVNz2M4sH7Og+1OT5koL2sxDjRaIU6FtWT0fLRfE/FCqX5lyfrRJhlHq
5wDO9iHm1mliHPJFFYxRmUPNgEzdgkUIlfWQ9u41I2urfX81uIUoFbZwuhsHTf/w
mS25pP7uw2nTCits4dqSJSMz5En5tEbrqcKN7Akl8OrHukGdbR99GdSy62BF5WpL
NnuRjUKjHakXRDHxp2xDnbiNWLDX+JqDZ5w49dAyiqlRnDZ8bX1uEkrMYjUe3Uj4
7RsdJRD84gQxOPTQPWwmyIvCKJ1IZ+bHAbylt0YSm6XxvtGpmDoXHeklQfvR3r9r
rb3gPdZWYAxDCzb93OLiBaBt3GeoCnfJYlXigZre9KouGCyP5De8D/crUZ6EvZM8
awn1gTBpCwvkjBYtWNzhVfYz81b2wdOGG+0LNVXEVRQSlKwL/bDqnbQxEUAIq1PO
bWE7D8l6oodQIrBaOOY+n73B/MY+BuVj/MuQaz6/DIB//o39byG1ufwIj54pL4EE
Cl8L93waEej6Irj2lLPGITcNIdSduIrZhEPiqOUk5b/qYjpDVERF/kaiOVwHDHfn
/Wua41u7XI6MkC7UsiHpxkvyTbIxo/1Iw+ku8eI/VlyD5jDhcpu9Ok5OeCUtwd0L
2bPfEBB2AkSfAD9W97560HPT8ZjayTrnyFaPUUb6YLm0aqOQSTXX/VdtOhviZtGR
shj4/3ievlRapKBt+SldMa26RSBH5px0vuq1T2/9TkP7ubpTG7JeuBFXLPSc6pE1
7JnIDgwvoaRnFfpAsMRpSWyPvWkswXHIy3jLevX3Y3vxr64Lx9nmQR06LkuPtnQC
j0eQH1JZ0MRdkIas4+Y6UGE41we9SWUoyzxb7BfKuCuq6HyLKVlYcEDbNRk8ATV4
0IqtazzoWz/qGOELKJU6TUbWMJP4EgpNEC4lr70rLpcl7GPkcYdA9UeUOrVg1zj/
jCKMkdk9b5u8L0XP0UaT8NlNrP/KdI/3mRgL0Y9TOOCpjOPv5sXbR/h2KqO/1Qnw
k1I8mQHEhfsexNGuu4LHXft8mATg7tcWc/mxw0F8YEIspus1dEZ7wrgrPc4Z5xK9
Jq8uJCo874k1NAWJ3f0PEs8aV8J3wXz5v13dlcPOuMB3nDZhuzEimnUr6udB6vJX
+jYXBTOpCq6bwyG3i6cSzDPUR4ivQH0FBTr0AJ8wGLSTLgOTg2ggSkcfeBhy8R/P
mIDD+/xV1k5JlGBR6OogIW0aC7RJY1t7vAAAEdNqdKBNQxN5mXU44cKhNzaFNtjd
0iMuGS1xqy/StErUWhJusKpte6GBHPQf2Sh9PSVTL0S4YbUuAncIr8jQDYdh2coH
yYpausU77wbMBja492s9t4mMKfbpC3X4ft0AdyMpYycA2zMzJFQNqmhuyHG19ToI
VZ2pFzBD4tcwzhC+R9QDXhltjce/qlJxdlJwAUDhHf8ALike5uxz49+2NjHJBx5f
luhmcVuTk8supvbfrjklmgci64rxBVfgl/yv0Hb0VJujPbXgoNaf3ylFM4vis2Jc
dZotwdErTmJpKSUqRq1zUyX/uWo6t4rSiE7nDJLPwICtOtVb6lGo0cvlIklKpvN+
cmhpf5vLigwWlvWxgQ+vUvI4T1nUal6jKxiC/RekspaTEB/oOHil02DZupOSlsKo
6jJ2jpnSEhE5qx9/SErvmIlNEvNYgYfXTMGg6QSFctm+CBHprqNqkX0hjrFIRGSw
JLDHrKYJanztWduZIGct8WMKdR1477d0SsrpoqxnNPxtv44/WzxZmVQjTOOxXS/M
NXJI/iPUUBDszmxIUlHIOOehXspjIMUiYxgdM+qBDvh09snvRS3taK+G2+qIMq7I
sA8l2l1Sa+3n5XgQbFUoeaSTleoVui4tSH4KEsHT+qmb4kTpdSA4LIeElTWQ5/GJ
nTTps1CP2bL1gK2HlUhnaEPSC/ntdRWcXNTgFHzn8+JpwgVKox4yIiNuvuhLUV/E
N0bq6azD5rvziCU3pnkc7PahpE222rS1CQyGVeTZM4kjnn3pbsdKcnWyhuDnlMFo
PNLd0RWPF+b++0kxosksMwY0t8fGfsqzIuSFpiAmtx/dIg1wBsiIBLkHmow8BAEM
8sDrOT8j27wnnKALC8phcqztboUzDPuKKf4HrguQ/aRhn5I5ga3b0UNELOyl5Ssw
1n9bpzcF7BFlse+p5JnPgk6PDdOqnlvcXf+1IYYrKJpnJ1sF2xoEGYJd18Zo8kgQ
ebehureMe+NqOkhIsPMSnCY1gd/X6z9MZOmKEKOKdIjYNb3EjQj98ny2DwbMRm1R
04A/IhEGswhWwG28xQ407D1/uKau/uCg+w7YyLHMzyQpRXupzjJMyav+i0aRZOzO
ql22fho0VP/5LWZN2+pDv5cHVrtJ58IUNGfjKkSa7+ost1wazAUgJCMiB+3G9q4R
cWtD3PPVqMTlonA6HdEJFnpDSGLlbvolzHr1uWdUfguEo+1LxgxnbWSyhiiAekCV
uYlBe1Piqtjj8AR1Y/arAU4R5oqTk9gXPPIJqV7am0fY1J0VgoR2VRal5/Mu/ZUf
7cw2Gu1RJ1sm2lPx4yK7s0jfYbcgPMohr7LgGHscTjCOJbdQZnhFpheKZnSZgdWh
PT3gpF1oBcfCWGMQ3MtTC/CAgMqMkEXN6eEYJ1K9v/dVeU2bKVMaztJRnJcz5xUU
44domLdG1US/s5pLrVjbkCAx9LuBy+Xg7Mhm4ib+LLq7h4ZWQic3gh0r3Ib+py7v
BKI4yFLANf7BmdwcMG4WqIc7St8OTl5dhmuh3FKEiuqMTx3c/VLMgJe3pm3msHoz
ItgdQrY08kUV57o16nAAVdjI1vVHe4X5BAyqbVArSOTuBkG0TAq2+YoCoWkFQzqc
KE/wOiQVI9qWC+gPXqZ4ZLatzvkI0okwwTe1FmTl0WW5VuNjjk7OtrqqzPfbmMH2
Wccpshaw3LMwyzYgYxp9or3W8zC6O/Bw5lElMTTCFQjRUfpTSchmKKNNlF4ZIp8b
ef33Df6IHT+D35ARzZ4q6EUl5JJZpZb7epb08kKIcqVP4K4u7aVwo8DlUnFXgOKJ
hQH9nqlONH4lAGAXOvFW+Td/tLgxEp5ga105efbP1MLAOTVQfZdNLrjs10KH2FLs
Ba26Xn31LqpPHgHjWO+pw9jkcOWFLSs9gbtGtaQk0lvPhhHgGMibHMS2NNdHfCl8
8yJZq26f8ux0YmwDFRDe1DXV6RdZSJOfJ+SsRqKgvyewLabE7NAQG+9HWJgrM/sf
iL96wjlI4Mq51kcqDXnnBKaYe/kP+zmD/MNUC1fzCYLjFAdQcWKuLwz122vWaphS
IKuJ5gsaTE9SLDAo76tpny8XSzr0eF9TRRBd3Dfhy5byZIG62TCt6XiKe9pTb5KE
8BD8lmTj6z6QbBo9zkvZiDiFxFyYRCzYze7KqaPoIfZyQq3EAU51vWH+G0/ufJtW
CxFMjBIrYrwE8ZZHZ4Qz9ea55m6YBRWW2E7Or6X76gVRipk1F9meiropRYdCxMtR
E34lTm3kcELF9ZiS+7CiAaxcbNDcAruPh/VBgQtJLxzO3K0SYUnDuru65eef2cc2
eGyJ0nxBHxONtDTvcL9fWrtpHDfNUuFS5KgpYpNJtlPBQucQCEaxGRYbU4dlRS06
el8odf7DBsqu4WP5lLSzeVjG9rkko50KySi5JVa+pxzAmjnurZW2rfcKqfaRxs7N
IEpVw+NjWeY1SXxnGe1HBvDILUJ2CA7CJaCwVEanTeTY/Rn/RdEW45GUgTGomrBs
TcSyET/esCptiu82x8gFrsqgkI1tfibKlkCNWFyTHgyFiTSTpDKMcAx9bE6qfbB6
fsBCfRtyDCAUaOiFxszb5Hqs/n91jm0TOrijC2HDr+dPgGI3p83OlPxHBzlpEhCL
/GvHP3r57bTtz0ZK2AcLx23kyjkam/qTAdwpfG/f0nWBbyOTHmejIF6BDh7jFJ3g
kwZOCiuMtg9xp7BTrf/tVmEiqcRBMEV8jMcj/tL0CHq6cm8pPPTrg4LmkGmKzLAK
J2YoG9wN8WvNfYtBz2moN+NQVQMi14LTxwfChkfK8rY1QZ3iqjdEhjIdvtMn1BKZ
Cmh1UGBg+DNGbPOZ+OcF7LjSW6yrK+OrquUC2Ps5OjBqLcAS1TsTXcBKzgi1eJq4
s8f+KP6lftnB/IviUuaectRhVqe6YJ9V/2kH62PT8Ki5ojsauzpEgwLh0Smro613
JBewI2KfovXlZ7v3+bWuiofhXKWIgrL4LDgMzG+zo7G0se7rO/w+zp1gDHU0OXN5
XGo9CRVZCi3CQs12gWDyDvFTlhWvi4seCcaXMH2dw6iHpELMW3vtgh6E4kO0VOa1
ucchLKJZfWZBxtJMqkycVkKxB9M8mZj9ixUd4E8+AdEStlPLQY0zhcRemyIfzrY5
yMGExH63SzzgbnXyIz0MGHHAO7eeKI2/mssDDQ3e+SDpx0gtAMaZGh6yW2pkx8Sa
P17stERV7l0GlWBV+ZHwRRNcVgEIfIt6A96JWixIiWRfE1REGdIlyWsQ62lRcWVh
7DGnYnrDCh5TLFTX+oqWV22ycDvrr+8zV0JB9uXd7vGZMu9JuK5ogdKIVjq+ELyP
RZfJn3n3Nz1E5pkOZ/fAwARql/SxW5MENTxm8z/pctnEy+Z5brCGXDpdSJ6TaZWF
RVHwwKZQUC+Ef8PeZf47BGtU5XmbQdrh8inmKpZbvyucPPvGFcg1KDlGFGoh+3dL
RmCdorMdsBJBn89XXLHTPiu013GindOFTwt11AwNqF/wTvcVVdHhNRQ+ZZael3nf
cqWC9ueYUvt7hUFAR4FrltN/zH0E4PaiiNgEej4L+/lvTCUMzMp1HIQzqcG3THR9
0FjdBchvKSZmOye2UlPubcChWp1UPCMc75pu2P/yg1xBbcUGcWVFNAs6q6TaPVx7
MQb8YWm/i+GGZ3cnCXY3Uz5OujBNY+X1WCSQ0NTfvJXvIEDfiiD4Aboed7t1BnpJ
S/xc0IY4PHfQZMzU+Tqzn1TXE07IbzDGjqs4sPCZHijjpY0yJgFYYA3HB//LkFAI
fnK/TelLDkdAb7HQIJOZSIYFILRGu+v6httxYimq/i2n5DT7ZWLyEtnS46UpV55k
OPrka4cV6gmu5Sc52ccPtXJp2mHWuF32C3hxeZZHayIN5NXc1I7pRjlVjzRzDogr
4bEkntByOvDsPZS9GpggE8m2NGXK0Hvhh3v3RigJXfzpVy7Xm37eGtCtaMoNFwPb
jD10IMTW60is8mwztg+9Nq/MNDiEibqKofhuefXkXTPOTO0DVoJCfHsFL3B7msxM
6Sxg08BmORrQc5wfnWVe5y3S7Fhn3DCd0031RPBS0pXBSZRSFox9s/9H7pb4nYqA
lt+KyjV7xgwjyDvWUcLTPr5tpNQ86H+KhPw9FIwPP4/WK2hDjquOJ2s1nk2riTDf
SIQ8DAZ3y4ZtxvqM1cEmp0CTFf5GH9xfKfVs3YljMKpjDErM9a0dOw82mGQbPf6i
9VkqHx5gpG+1E7e2jWIgdlRX7tdOWHxZB2VxRpZZkv3b6UYEaVqNxw8cmK2UdUKD
J1oMb9KHYZOy7Ay2nuJaFGuBM7E1QvseL/niBipto+dFw7oZ65hO4EQnzF13fBwY
osxxvNK99MXccRhOTXN+9JRDDT1tomEZWkqF6TTwW0dh148SURfMUnmAdWsOcITP
ctZxQ5WV5dF/suqIQhdYJpTAlX+s9N1Qu1qj85PwlVjo4v85rgEXCCtQzcnzbClo
JJMx/ctNJZISXYiLqdsZQpWgu3qRIvGsCNyxuqvKBeLq2gFEFvRPYniAb7GMUQDM
FF/ARFN8iGswSwbO1//2XhkQ+WxMBXlZq3D2Amest26xdrzmKyypgQvroNLte399
`protect END_PROTECTED
