`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jzO+E93T8yja7bWUaFvHRG8HnA30I0fT/nv8oYVJEqw4t5qdlBCyyRRf3HE/YHc2
qKgzeoafNRt5PE4b+cEwYEgckyX4r84s2BUVJPFxjW1j+Ma/GpOMZLcbEXgpulid
r5208eLdrduvtAa+Nsv41gNhMUa/eaB548ucP76tKcvyS/I/yIt1FQFJ/XaTTp+D
ygNIRPsMpyYOqwn4/0kDPRDS02lNLNm5zRtDZwfD+wAAh/r9sVJiExxIrbrCJa3r
6ufkfXGCIqjIirvyPdGRzzWbWtRl7H1uEjnkOAbOfzTg8kWF63mwNXIWgp9SbDeb
xtR4eN00bU6wq+bTLMrWAKw7IX26LyJbrovKIb7U8I3FOGFzrybQfq2tPf8wrob3
XOOhwQzcSXbQG3c+tp0uEIcKW1xSip6R97UJMRwtrC1dgNt24z2y8l+4RxzrdCiY
Jd7lmhpvEtrfFU6XsgQGDapemjBJ6mhlfxUp1Z4pSW5J9ceWVEBH5d6cpdgNjlQR
0hKBWMcdbZHGbjdEruxFjnz21tUOnZQ/a524FZOI+BL9fGITd/pXZ6XqCc9LmCzF
3j5CBV/heuxW/DGOse6StDZMSkAICRoXHi7Q92IZ6o8weyCkYkTOWD5CBAwz6Bkn
+MEIQopY0C/OKJ3RSL6Z5A==
`protect END_PROTECTED
