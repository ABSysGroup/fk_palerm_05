`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
10za+oZ5n0m7B7LgWqJPQzKzdEzyoc7esS7nwlnYncR4J4xDhSYJjzvDWnP+WvRQ
yHMijU7GVZp2K1l4Th94BQuHbIq+Fy2pb74vegNtZyx7xc3jPr6Y6Q6TneL7vK0/
ObYI4caybrE7Ev6nfnQFVgcaKdH+haKsOjdlSKe6VxAtMU1Ux4x7Tfwf1Nf97UqP
HuDEoNW0l30QVsCcdOBpn8HglsMiL8D0M8zakAqCaiq0lMzOxoGET1scMf4OOU0D
NGI3ntwE3gcYR8Qfcp0o2rOUlmG1mW6qsubSeW15EyqTS/vm6cTKX7YzpOiWYLA4
E3Z5zy442TZ4OuH3132qA3JrsiwIktvEiloN2oj5PsznHFRB99ywyx7VcaVEfGge
rxIWVyzxnpFJGyqEj877eT43xhHsxrUl40glz8H0zCuWD5syw9R+C3rX5xPd/72p
oFFxcbfyZ/RYzUqk1Ed9KFf1Pjlsz0Dpoh1+4RWHNMqrhePa7IJ/5M0zxJIrBnxu
JqrlmIJsxLPopZjUynbDvcUHhqBeysVb3kTwnpamri7XUNMjADfBzdIq5YHTIvuQ
sZEOfDS0Pe0fOEi0L6OWj+2QabXOirAIIwPm1eej2f6NGGhTxg8E2zE2/7VUTxqy
KM7gnbbzCMtnIZuuM/eJhiO5bNOP0gdAevxRAMhmKZx8GxTKImjuJLN1pSgGL5ag
82M52u4NQT4t0mfYkglvaUCiM0FO36EZLSJ6C8345L/GDKhgoCsEqDVBqgFaezq9
odkdNVT7CEo0IW3XWXsHHXOx80d0fq1CMTMINhMGkwQXD82YGKDsa45TXWWTBCZG
TZWy6XLpKuCLmuINDCA7J+HRjIpksyncbOkCoZgYdPYT4Bc+59GqcHw3Iuh6lZSG
AVLjPUnqJBqpti55TM/d+XUMEF3ljgoYr/DPJY5x4ycN3oDuarbgki3neqJsAO7e
`protect END_PROTECTED
