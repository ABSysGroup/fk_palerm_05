`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
klmwTED9hZ59HcIR+T6d5TN8yCoK9J1mkWejUhwW5p4v94Kfg3mw3FgPvuXfbrGB
iBYZs0RBKpdqavLb4udfIEMUt9CXjH/ghLqr1rM8o1Rux15b/tjokcI50d/3tzcG
tIEPgNYB7NHJbZXOBCSMy9XZpQqM9ukSYLU31QEmfjS2uljdXTE208KxyGwyFU7E
BMeFpevFVLYsMH1YqpjT34ozkRgYHYHRmtmUJeiDMBVA75+sR7WQkOLlhUstsNnJ
ddbzsxfcVX2BB0Ci5hoFdg==
`protect END_PROTECTED
