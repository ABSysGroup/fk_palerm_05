`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EAAN5Xmg/RYo3dOj2kyF+l3NQo1wvAamHsNtj7cLINd8HaP+xIMNQmtEZod9Udw9
v8+W+N5YgJoxIoqSPC90VA97cQCQV+4QAcyyGCOvCIBp5rwshx+mfjR1ACmrADzM
ZoEF2iTP4sZ561lUi/57rWPi/CLUdMfCvcNM5sXsjMM36jb0zBn2IFO7OFR/9PhR
EddlqB/ImZ7jaMqfJLB+4RiXD6XzoBihrBojxNHTD75VgHUfRmhgd3E6kb7wpmgL
VL3LcO28qPlhUwROy2WBs3/szyKT7uZDV0740VhXTm4TJvMnjfXya4xlvu/shqRD
Dr1OcK9CNYyr9UoyuzlHISP5XXNEk7AeU4OGuwSIW5bqNe/Db2fmeMsIBNezCbCl
0mnDQZo6PoLBw4BPIY2+w3GK+dUygCpCXLeYmZS13KFT1vQHq7rqtbfM425zs9Ub
/fYJmXngrW3sRXCjA8KTNXK97+nADgQwnBe4rbfMXDHNAlie1EwDEpTUkq8jbtXg
eLSjmMf4o7q4I57r2wEUA5NEjc4GlKdQFGU/f9PDtpsDrTL77tUmC4J35J74qpo8
t6pPIEWiy6fe3rPMiOwbcXoyYjzevBP1t5Rb5wBBr8o=
`protect END_PROTECTED
