`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6KFLVbWWVwVaThhl0HpmB5wPxPayypSGzuZWZsJMJugM6BhZcBH7Hx5Maa6NPXPQ
4ew2T/aLGfQwEImVkq8WTOhORoGMFZjs5OQ9j1WJaOcOMvXvmXSVAtbHATC2awP+
hwizKrD4fV4NR/6lDJ7fj8M6MpAGIRCKNpiE/wctaFrB08MsWh3er/5/VqqFYqEa
tGfLHZre4tRdA92nuhnj0zXiCWROUoCQAlvzhzn15dMfO52hzN99A7OsiOE9AqY8
nF+QDclomLbYlaYM9iVOeb1NgfCN6T8c9IC763t8b6CVXVE4viQuyZ06gjKuUoDu
8vJIPppVG1h2WAMkC2yHccbly2pFej9uLWJNyrfe7wbG/SG7lhM69YQ5RW6/SECN
RzQsR/g4+A02hAwJ7lA8BQ==
`protect END_PROTECTED
