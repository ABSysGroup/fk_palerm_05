`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A067fYID3Ho61JF2gHWDFQAKiha7i5uV177UIvanMGJTPTnRJTUz2RYiLytZARDV
BqyNRNSvWKPrrJ0KamAO54x5XX28nFYLO11IMRyEPKDqPv9bVLoG2cveey2QDGwR
6oMrOkpg0rfTFk8jICxuEcRIwZ5sBV2DqLZ5JwMU24f8nus5HPgbdJgiPV/Bflvq
lXLm1U0UjXLYK/kW+NtY7eBV2gWfFaDfQL2mT30HeCG4ywrWfWrF25C/t1hvXpXc
U2RfGfTzrmxvQBXDbXk0YkyHJWdtA3vVmSYz6EofeySD/LFFkWpbeGlr77ySJEih
mdgCi0byahroao+ZgdO0B0eMm07de8hxUASkTYZhaxwHwULGUQyD7hoXLc/JeiKC
TruM5ZCAblvzQw+C8oAvu65YLCzOwKWYp7VZFxyyQjl7AiirN0KZPSP7+r7RyRUM
D1hQnFAz7o2mdJJIcUMUy24Mj0vomVD+/r0OSDzeqqTtGJ/UFSrQwjase8mdBo8l
GPQ5reDibpINvvJFEzc1cL68Yw3NPnM1T1g7eFxlvdD6bcLBMTUPadSbfiy0OHaA
cC9RFHJGzAtsbZ7TtjFf3R3S9tgOl7fNy0AcoOQpmNRu0fn1RfkojUJQ0b9VcvpO
dSKplFMWTKmpyk9qxAcV8eFv5lH04mF+JnhpdB48jFduAZwsIqRs4rFR6W1sA72O
Hat5B7xkWcrz90vGPaAn/yGSIgO8G3Dcyo19XLKmBy861mVnYNhRykaFTNhKSrtA
An+Dyui4pqixgSS10asfFeE7VHEJEttIw6XOw/O4OKaIBktQ7E1N/Ulp9Yj5ID8c
CVEiX6VnaI2/9h11j0ujPrJ6PzZWdVGeyAMtK1+3lQavmHuFfF/4vZhqtcf+/U0H
klUTfCOhFThiorRspfEA//Vb7UiASLfqoJvRIbxiAA0stBNqr/5Xn2jqZ1+I/UId
`protect END_PROTECTED
