`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OuI7hCn0lOlZXGvwf1TpGimAB448DCb7iKcWAM4GhbnxRmVt1kFHW8ZZyrZlTXJ9
/DNuYqrL/pb3LEN9Jd+/XnrEI0uwECvewgxnaeKWmSZcu5Uq1CJPlC+pXZDcmGU2
jY27pYI0M/pG+U3XxdWfDefO1BSO6G881ZcZtdooTjESRUVNtJVc3QoTM19fc7Fx
CtuVaMna2mMSdULgaNWq8HPXdosp0zunrQ+B2aPW6Fn8YA/SjEPTkqZR1eljpAfR
QMFEays/VryOoJTwRd6KJSERFW/xKzGsj96QPwgLeRiCJIsHe7mfFz0Ez7DcASRZ
mmTppx9ElFBUKmbMFztcUPUQoXL2Yinl+w2BTn2jvZ6cLXw3Mpqg3rSMeldN2CK5
PMLTQUz9ETZjLwUSLpaUOVeoIWDLkjlQN8+5n/3LYZSwy6Nqrddi4qeIdzplSYLk
CfmjlM4HtsYV5hfQLFUgJrWWd9H+eoH4h51GeN1hgnqlLfq5Zba4Y0GZNiqyl0vk
c4XKuOjijEklZeVzhYejmB5DafEh0pIEqbVirxBscHNZvc+FRVJNnKHuizT8+epg
cpjLOESgBJPxwJ5ik09NYjqK2MTZA66qbhTd6yRh89EEAXuz18x27kw7enCxjWQB
zfGfGpzf74GioJyf8ossGRRU0p1olkLle31E1spLdmUY3iPaQxVUi2HOmoKdSWBc
H6ZOf5SbfDxEU7vdzr+ZjP2RE4+8PRdgBN+wqInnsE/rQzeWWEH0ejX6duWTgUEw
a8pcIMXxPzTaE8OiDrgbdXO/GJE91wi1zrIvMqSlldwMAzC37ENDvS2hvm2zl+RF
uCFR5/2dsDHUGUNeQIUnBqHNRB109IwuwEtk82Nb1nTKQz4b3yqHZzwmbzvlsJCl
w45fihdqSDNhpS6QDqf85A==
`protect END_PROTECTED
