`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FUy3lygkNJr+rCCgVgFoSh/x8dya+NhJ6+0UjGxlaM22MKfsZynjh4nard/zkJnE
hwfcACG4Wrgvl8FdO0Nscfz2vMh0c8OKTY1VsuxppBJUK4Fm4BKSRtowqHuReZUh
ItL2wjJQh5cb3k2uCtTivf7Oa8+Sc0ypMWpyKXPfQUZpRFh3ibh22aeow3dPsRf1
L4WLmZogvPbbn/gTQiW4RyO33g+YOTEhYk+pd5z8VW3oQiz8ejx1bpVNpUmIIiE3
VVq5gb+o9icRjlfYYsra9V6eDMtTjNsJAgS5vcq4G8xwXlSQdq6Fk1n6zRoLPfwX
uOIAigLxNCG60O0rnBy5kEpex9+EeWHLo68EuBjdZIynzW4SxFa229vyRIx1iX3l
Tea8EnYXdfC0iNAM4p58rSgMi3UKIDOpyQienXO63nkTKIS0ZUk+H73Vr9bfnC6E
bXG6Pczf6FJP/0/peYFN5feaYLzlZNADUZWwVLjkdqZkSLRdud9BnYFsyFWo3YHt
sh4Z6PogDDUKO1Ak/Jyg7Fj/tUi5o+t4rpsbCR28ht9NVUadtg/9A2SXmknZ5dbp
RAz4cu/Pjwr5Nw5j5eagDVthqknRh99WR5SOnpA107p5hubVGZZCbjGElHX4kWqV
pT5O+vLtAhPRhD2bNjU7/FhDHaYsEgvurQ7FimQzRAsyA/MBZPgTSbH+lbHmYg62
52yMz5tf7JC+Q6vVB76ISdrEMVaiKYYJWlOjCqQd+JFufa+Rz3HOcSvciwKX4xgC
mKSenoIv2OHd5rZTAUClwI4whgrfgNn+/r+QNW00goYP/YFh3m7JRu6vQVlgA3VE
gg5gQGuDYkRoc3M9aPNjBf91oJ8Rr+XvlCA4xoYjTa7QEaz9fynD8E4g+nZMvwkP
7bLkB2R+NG91ixao+DGMYAUlYbnLkkl8+mULAK5TZkum3MTZq5OOL6RhLqtWs5lA
uB/pWIM0MLIGfptNLE9bRmpVx2ntUw/QJt1wjJlfm/S4sEEwrxPoIZaJg8mwye4W
zX7bEWrCC6LzevgnTSv/LCUIn/4OQGj05n9CF0E7Y2qNpcI0GbpD+KqmSl8TuzgV
/8J0Fdyb6NF7p8/s/uTzotK/C1bTCTiz+0XIoFQDx9gjLRPgHYOFbklmK5cvu1kk
nk9Omk4NyJWvJPJXK0AXN9+cGrP2btxovLDdq6wW87jRjiedozwgonT51cySjHc2
s/EqqWdikqpt/GvsV2JmfWt5bWrS53pb8evul8hjWEE61tQqHDhR9mvztVmOdSKi
rJBeVNJip+6lM08tTWz5gvf3OesWv1YaYzrd3T1kAmMYS1cE6eGArQOJFOxEjVqN
T39kYt9EJS5gp+C2Ddf0Tw3tLjMVO1WrTOLVZXDj6o1Ou8gWEqZ6wbwart+TaTbf
7z1NDVjGVY8qhwje2OHxhhnoDRyQMUUmU12IEIIWiJ/m6YNpn47CvcRUI7GdQ3Au
8JRcvTe54IS6VectgOQh+g0tBQxIUUC/CHCMXHd1ro7X0QBjIoKU/Fna2ABFGxKX
sDiiIWMkpfqIis5CtwEDZopcRO3rCIErgJ+wCQDjPDCr/Efs1S+/zIDxsU/akwur
`protect END_PROTECTED
