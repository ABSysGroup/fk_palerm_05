`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RAWJ4d0HZq+Srk0lc3kXw0oXPU+E7Rt7mBN+Kho9sc/mtWOOjhDmuDY1cOTk9oMw
seft/zSnKTUfUfr/4Pd+V9gB/OLNGISpJqg4l/HrXtvQNoPyNXgzOsiDqXFvYjez
9Ca5ixNg0ad8y8kf3xy+DcXNWXjQY8kHtG1/OdkM/HAkwX3xLPDzYl+iXoDwZhJh
aR9gtRXvy+HExnwgxm/igZOM+heskUSZCY92tTL2ACy5RIOjYfd7V7RHC+8GMtxr
TlQxO0AT3HNxsgVvMN2xdq7wZOxhLmbUYC4/HJBYzcMo7dF8dyvJhvg80L31mfCz
ZsgskPQsTcTzyzN8YSMpwDiWufWQIIjCaF753V9rAfayeFRwwzogxlo8FS+jLIv8
jbAXBgLyxtbGJu7tfUGegbnzC3ONGnZT26bz6BooKkmDtIqz21vt+NzzGWrgwD8h
RC9JSAnUet2Viw3lR0QpsZbN5yed/VmrqdFeSaeI+Duj3x6IXVuQZYAuIHhQfJaX
0Ow3ZvWp/M+tb4oj9vyg6Xe0xFLdM5RKBxrsoF5pdbmV3hxSkbFfUNOjIzMovRQS
5lCCHLsySvpvVcDGRDk9OyAGaVXV8Xgo4c4Ll9/rMwjG5Bz4LRbtCn9ppLHaG7lY
O1Zgre9kdLUxZesxGV8FmRIYjZj+/gxn9b3abvSKVRi+uDmw6CROXiMZOLvnxwO5
cn65JiVkEOpodoMzCM1VCpBIwPpIxpEF+i/oKePA4zwG9ZfMDlcqHEqsCWk16KIR
f/utzPL5emaxd71amh1pbLLfRLELASxwtfM1ApX6Bo2NHjMWn1knwvfARhI/68O3
Q5oWYTj2ilAsHwwvaDBEysll76AIZk9aVl9vEPrAYY5+LZ1+SsXRPQDHplVCOcjE
ymJKSJwotrya4omFm9Jd7fri2JPF7Yti72XG36/qocoGHhXLwJ7CLYUIb/oUgGR2
PbHB9/ZrCNk6mQtxhRvjdRYMYJbullpkbgNL3wU8xKGX/W/iQ33s0DvoeXzfzsti
`protect END_PROTECTED
