`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FqlxE0mOMOWL6OWWp13KQG2r3Au5lL+1TlQHMxEjUUlOXfumk4lCO/H01+DW+/ZQ
+a7+BQwnXi23Rlgl2Q6xKSYSub6m8UEgkwKRokRugRgNX3PNlZThs6ucLO4jI9Xu
e79VTICW1Gqr46KOJtEwAlUUqbsVDHhUn/Tx3tBe4d1L0htaVoBBeMoPzF+LG8O4
kz4TJMvBHxyWB5m5NK0J7zUuSTYhmdc0xH/mdBfz9oPZ9nWclLRqOw0mFxGv01Zh
bmv/6gCpA/i7cPF6p0U5GjW+oipIdDLvjng1iDIWC662lGmGvN3OMENYYQzvCqv0
JkpSPdUDU8Xvidf5jUdLzKxStINjCUcJ54cC1my7bqF5csmQE9G0PmzI5r/wqiYB
1fKbMb1TCyBjENdp28aBznV40rowlJTnt8VCpxBhzKcUzjyBmQaA1QdGmWW9P4kU
`protect END_PROTECTED
