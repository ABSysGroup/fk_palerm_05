`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o/Dqn9dpq5uF3DZDGpFZKHO8p9oVwwPCCzN9HrC88kxvDrzSvlhu06eakgIWKURJ
urQyREK+AuOZaJxZDzB2fh/a0D3jWsApYciRkSuzd9fQV6wGJLBQOA/Vhvq8qcsb
N5fO4VjuI44uhZYAMTCVq2Ny9Oknv9Md1rejiwGEmKC3i3lFueLSXBbjZXG3BDDn
8OWYQE3QglVf0Vs4SGW2uv+F4RXEXEXDu9GNS66dWKzB+qbTrQpKxXqYAVWD3Lbn
wmeFni00phMUUaEc/FYrpBgEccDIQt9bw5zDZaCa8kiWF2KB3RRl3yj4cPNC14jP
zynC8oVpBlKQWdCYu8cdFerABtearq5U3Q6jY26J7dL81sOCRQu3r7RduF7/g4hz
lfe9PDwTTAjVKJSxxHb68Gxq/oVsPzXExIVCrGypRnj/9fkwhLjp29sf9YOxmOi7
ajfQ5iaqKNgnZR5//gv8Mg0wtcpAvb6uSCcoumVATVduWe4sspkkdgcN5OqWZn7P
Qg6F3WIuC0jgMH1LB+BYzkrFTy1idUmS+9UrF+3ijR201mSfg70SGaQACW0aBnRO
0tIMEHOw8nl9/n911qiz0CVThIYr1Ydlodj39G+9zlz1XVbeYJsENw6EwOZIX2VH
sUHxxKaGI3lg3pWHyrErMLY9Pkrz3eDwBJt6QTCweSztHtYgt8xzgrrD7iEXybl+
A8xPbb5pBeYc5G/OHqLvZ3SgKqxlN19+DVBwmptaiJ12DA5ngfiN5gvD7wl5nKh2
vop8ucKSJeqKIRzjXe1aSpCrGCf/AIvNRIWetb9WW1mDX1/+qtWqBMKN7wGNAQ0M
8Sho/Vm6JHbcdk72pbwferOwmxJyXk/ZRtxjXFa5eY+3ifLq5k2Sh4IU6/+2qwCd
b0g3Ag4LiEpq4mOZ2AnPmRlJKKru6A7Ye3eoP2S3x04nJUWey0IVbM1lWP18HzhB
uAdNZom63zoddLuyku0ufo6e+HYkOutOttX1TUuKkiGMuwotwo5Lg8Hwm/HoWDQP
bw/snS9ZUe9xY4lCa2pcyUFhcz4sZ5+5IqkskURcmCfSo1Z+7QiI5SgZcVLrv9Bv
a/zrekygAqWUm9NtX2MAcs7JhuSNxl6DGzXbswgYHXLN3dTtYPUAGHLam5V1dlHf
IisEbHNjsXG3RCINNp2wkFMkwwWWDWHDbNwZMsZn9e2xzc4wn5fX7Kt6HLHivQaD
DVnDBoywLm6zoZLNxP3hwRJbzC9MyxTxVnCqKcDBlfvGTTrtfvV51wY63n0R4dAe
ccO3s/dOsXvWK6AfEYP0ik2pN52jye9gfivh/9y2OFOO+qBPd3CGTgpzASrGUk54
6THq9UZbEkaFckMNVNOXdLTMA3RLlohDZDB0VzSLNIzJVSsOg7h409ZfMy5hnZPQ
LK6JtuYRB+DSO+xuffcU9xvfSMWBh/Hz8L0813/7Lx7F4rPSz7FTo6RJn+LJcd6A
c5Nmpt3DyeYILlmG8DL4lbJUIHJc8IwLyrHmXGQMWsn3Ftz5ZVuyfqg99WeYLfAu
J2NiC1ZXOiAT5wlf93nvKZbcUEhqh3Q993fBTUlzC8FScgPedTzMLjU68KZFl/ix
T+Jsk7AkYrmXMDL19cQ+mVVzwDL2fpM/DfRUrekaz5WnqwnL6xaE1piNB3AWEHBS
EMXK4hevSGmB3TzI9/Lw9gabpS69zb9z9FaKJ7Wlz/BMwAlbXZkuPDG7JZjb/Wqg
Ggtw6SDRwLd7yPsqjkoyR1gUSGEsLiCqKuSLofBci0VMbKdw9eq1deaxBZ+GoO9t
MLNMFmSlxGoFAgE4Dqt2ncfPnj/qz1RRhNCjm9zVloyFbk7kiCgKxqraSOnAuYib
2AyvJXyZozCWavUG78VxzI+jrhWxxHOQnHpNs8u2msnwv+9AYoGle8JN/2H34UfX
ntuuGz67Jd0V2GEUBb8obD0v+2fFXKNMJkiAxTpMG83qwf6hMN2km9buSLUNtmcG
PC58aLO3yIes2PuZ9VDctNpej7FcVOlth4jnv//rQex9AuxOE2g1ciQF4/8NPgLu
MgpsU+mfityTdhGHug91J184ktGizhuBbCKsc925se1uCd8LK9S3xWs937kbQdWi
ZfrECDiO92k7hA6oO5Kd8ma6uRZyvZnpxheyDiYkHqe3M4BH2TOBqpTbLJxbLXDT
zE8Q0HM3k0wPZN6Me8tvRajqW+vx0/4y6t7qkmuJ/nNaa/ABlaMP1nWQlg36cRMW
9xmnPiEevNGCMp95KvfVeslM26NcI3JuxEKISd1zCVEp3UjxlBgPaOZhm/zgz7xY
UD+qZdU3qflcl+1Xlzg4khyDyT/R1fCxgtGiOKibYVI9SBgx0yPU/lBeAMJeVDqU
OPNt5pVdJZKNzbZxUtycsYFqpFaYg18nh1Jj1mbmQ3y4xn+mxeXVKvuFysLdbFwS
eSzm025W5gfSg+V9YQYni6Trrhhb6LT5m1TZj7uHCArTLMAwRRLqqhIbcVUxvntT
RIk9xzbBn7ig8kkA4EgAAwFcsa8pRSMMwyC6TJTdN2hkAqpbVgM/DSF6wd9rr0MC
vAjytUQ+Gl2i/CoB3RH3OvIR3iENvC143T0P6P9fHHpwBkJSjM2QyaSNzae79vU4
xC2tSl26Chq0T3L663rtjRoEzLvw311KHkjdiK7Pk/rAeYHUDAZsILMH9GcNFEyF
th3P70N4rjXqvcwnoYldA9PpUAo5AtBRAhbDSDER3ItyTD0LfO3pnc+N0f/f+FJF
Zv2TGGTP1Ud0RiQXg88nIF9crYbKVaV5GVP8hVtgzvfvijmiv+Ris5OqhMQ6E0XC
jpuuG6ssEd0+D8XKfhbdn4cRwi7jd51QZUq6MbGugVf9nQCmgZKYe0tdVBTHreEl
6kLp8oN9rLB0jiuw4BzahjWvnSVTNbEScTs/jYqsfepJrBxXN+Ze+tcE133GCOX1
G1jXDN9RJrPZdXgzJ4jIIlXMb1fXpbwudWQW31uIdIc767ux4hr56EKoA+OxdaYI
ETro6m5MOTreTyWyMJ7zxDyQbKhURZnaQ2BsoFBXpeUlvfPV7QFFl0yqVD18R/o3
hf4dd2AoNdM0W9S+eZdjNxF90l0OVvQiVk7xQecquXjm4TRReS4j4wkB1FSN+i/1
XZ02PRG+yifYy/7AU9Ox8ZXhQZ2j0GF8bsYVuyhfuSc8eo5EDWnt5xs/Nt28GAMb
AoVl3bWOuJsg0B2CE1HPIu5SmJkBMZUE9x/ts6zMmejVTfa58NhG6dL8OjHO5XNP
vAt3u1+zs8h/YXVXIdHmq0j5077MdqWm/bMmwA8OKqsCcz8tJKlaM9hgqgbUJ1rq
RagAJZJExKwAUl51+lZXsz0GDzd3W+CKDXPGUHXv+t5yd+IKYUYgOU8HxGWU8nfa
w+Whqo+T43b7mJ17GZqguTnHZSOJTeam3Xubi5+JSa73YbxKlRkhyD7KBVq7Nhsl
KYju59MVCwhKMhz1thf9tnPL0ouX0qTHFOm2Q2ZhQ5hYS2uJmS9JRYhR6bIeiX4B
YAee+wXjkVfJU5spnPlWOKoVbfSL409kYQahgC9enH3rDXdgQw62nLwXBo+by7tc
YYjz94XmTX9ch6PQ/ee2WuTRMINfgtuv8D7QpXYd7Kg036nOASem0W2dsnvF3GDr
er3fZ2i0WTV+iNJGvQLBHVrFrKk7gHhYAH5lrYK7A5tcqob0QFJDl3z2W/0Va5Tl
aN9FW/fa7EBYCInGC+VQdeew5IvdrpUS/HY3BiMXMXSzZehdWnum4M9mSNXpFqee
Zt8QBIyNmWM/IDPwBCDuGcwLrUtNmdt0NqOxHWEqXXb3KU8w3ZDLFkSSLDAaWwfQ
mwiyOTpTva95p17UHb7lEp+X/8SNi0LaTWCqXgucS4yAoZcduefTaiMTNm7A680w
mqJP1weRjrumXQqOuv2LJImi9Nj9NGpfvyXrpAqo7fMSf+yrXW1ZloA3xRUaARWG
dlXMlwyw1F6xV4PyfFK7Y0owvxaW9eyb36hQ5+109OrICRTQdMRY2wNWHAP97+tD
CSbe3z3Qmu10QAe29VzkaZv+qs1Y+AcUW7AQxjnorITpkk8Ors7yidZd9gaQrx4Y
k5UrFrPxEHZ61SYGBBETaqb9osdzj1jNXYEKpRPwdwFtwCi0/9Fzj76Wa9ygSQFL
Vqy1cuvjfnNKIo5+zLPkpMM9N/BviFKCCt8HRfWrsm6ItwQFbQJBHdJ068g8fVFE
nO7y8hT0c4kKkcTk5jyxW3aF6szq8SUohDwyx5RGOUopi0ztWFZY4oxKMRPmrJl0
ACT1tSE5VzuIkiifKMsip6bPPevQ2mY4nCmGnADfdYyET9vyDa0nbj0zB0ls0uVd
7KONUi33OpsfPlTB4HrXd76ODdsQybQt4patB+OMhQFEjgTU7uYBmODaS4hs8X5i
cDkCVFbt1+6wN8Ik2ZQyjPFs8W12UtuAYiM4vWXjPFWtD0yLCYX5uQcAlsUlc/Q4
Cvx0p9n0idxQnw+S6XYyyS/nedAKFMLdHguBSZ51GhZpa1xxl/K+qfaThBRR/1uG
BHBPkACjLk9Pgl1Uxk8VnjtpEBrKLtmtlkK9CNje9mA0VaH6zpntPSspa9UW60PG
C/z55PJ7cl5jhQ0HNdR+5xg0WDBmQvqDDOF4awhtbnW4iLW9ugu8+cxg3NnTWOCu
eCt8Lo4kvrcbU0ORfKtSLJXCNC83GCKvwdV8JaXJQilZJ/2xIa6EYMXsjk/zxXe2
qRJxE+CQbAMJevZxgrbsB1OpFa1I2XKHr/IWcvtCIiyT5D10Y07Vv2s4B1KodavX
g4VaJDJjNy8kA3wH2aQcH40OJFbqbfl985OU//vGJvXVYXHl7Woy4Q4CzraWlm/D
6kFG5QK1toFpR2oZli07ry/ut0lwj1RQkn8eBTqQx/2ZcTPKBURRKovtCJ6zBLmP
4RMPtzmBNVrWGxps/Tq7w+Tvbr2qiTpNyPWCEdICoYI2US70I+1el+qxEQPq8ylp
yH90FUTcyIyqM2NI7dwW/5bN0NWzyHvsoDYo8s0q7rgAq9Ukt/kvDPessNpoQVsd
NV8owfE1LWKB9V3J1JX07CCg09z9anqbQRSz5NfVpmAnLlc3RaM1D2X41Zi+EzJt
/5b1QlPpyl1QkGKRch83qhtYa/G8Am3XfsHgT+SjiORgNX6vRiyTnt19KfekLV4p
OUOLOmRxC//RmCi2RtSnwxg5kUZntudf91qHVvu60eq329EEz6Dhg96p8Kfdr1hM
4rNvBso5gZuYXth6nu3MF2hNTpNzW5j63aZNT2y8g7VkyGwsLuPM1ogDr0Mc9z/p
6Ds66QOruXEtWRRnfgPIg3f9hwCp4C2yZcbEFU7bbxyMLfISnNp2WMPdn70guwfI
PCrO0nQ/6eubwmJ4FfEr69za632kBld65zwpX81ZUZQjxXMhhkMeIJbDZTNQ7YCD
DMpGMjNAHYGbsK5UdLE8bKjfZHN8dYVz0CB5gZO7ckYbBCmBoeNmmtZVA6l3ajaf
RVFUoeaDRR4U/XPguRSYB3O5J/KewhqvxwXkEj++idtSQCobGwv+0+wI3XDm7goG
HufQgdVM+clXzupN90W6yC0aTtz/3GP42dLXme+RfWXlut1pSVESJxHn+Llxj9xR
s4SKLdiebwV76nnqqfvj2P5n0d96SHLU/SdHzS73V0TbUQ1hDAXGcc1NH05cAdV7
ZZaPne06bAVTj58+HXvdz0vORk8ReycoFKCxcxRJnbuSljCH02krWFCf6V5Lzmvm
dlNEESvsmQ4c2RyOFlQY1tadLkwS1i9C+n8vhcrIRxW85VoZJr6uKBzY1sktXcPb
0LGu2DfFxqDMnA83lrdunN0izWkgw3CCHIA6ORs7t7ar7M2ppwFEFuuzn7C/Fm2t
EfzWSBIylGK0LNBukFKmdoTSKI06L0M8TSKktzvLDI0=
`protect END_PROTECTED
