`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UiMdOHw+NC3GeuqpMewPOusvY0kgX79o2ZyDV6G3btOnO9pyGq/v2Lz+Il/zhJJK
wQ3TYpjUSvZWCxz2G2cKceX7Bt/inPEYhRIje6ACcSPN/AzBK2aTrz4HBuHYWgxC
7aUXMCEODBy+9TN+bc2HiHxKbHmAv5mRdO5ZiJKNyif1x8xSVbQKqwJLMAIMSWtb
JywzzuJYR97pxVaXn78PO71dgrirUrpeiDSn+9bFryMt61ETbACv1298jK828R69
x1pPYt+iOdRlUTn7I5ssrVgurYIt6T3f7qXEd86fNKijmh/5UAQog60jRtLjNnwP
yHLHaYBR4QU1EVZHEEx5k9rIKYHnf4fKOxgveYvq6JzUaJ7oXnOH5pG5fujAYFNg
9YkloAJr84UV/aSit4Dj5Zg0srPtW4U+pqs0Q77v+7zjawgDus+/4lbKmqUHkINa
`protect END_PROTECTED
