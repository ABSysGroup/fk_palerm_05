`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lDAc1nZkYXhFRtcDpeNcQj+BO6JHaILO7GWsJrHACVU1k2sPiktElcocGMJIzmZi
cRsu4ZPzicgwja73EA3/fOjOWOonqVRFhuCIlLLC0Te9BWq5A1lmoahA7fpMrBkK
ZG5HnXrTgwJgduU3AqbUEoxoKdbO3ZvKqBOFKnmjB3iYaNzaF+dWpIMHvYmvvPXe
qlKlLB8i+r/MNuhjGjMnY0S8zyK4TbVW+/2PkjboTWvnWSt3qJqZL+DKx0k+utIH
CoUpgNznOBkegJkBrOSe7Povf66D6gZcTyWyG3e2rZYmmanOZOfDLxPlZxtcishu
qBgy3jTRnz7Iry8s0knJiYLonYhdBEJJAadyG7GxuFtS2a90mhonr+FbJhkOHwRf
EmVcdWhiXPV7EAuFt6a4EUTvnqtdmg8m99xD+GDzo5Rm1kAP0001kfmD+FQ6Bzzr
uO4AvAvNclJtutCjLqmvwtLx8yyRaOjPVMTHGI/SQRXINxKM0N83F7xn7fK99HV0
zecNyEQWf67+0szZrBHKfJrQ69vgnFAhf2CWH4F64CR1lKnCTxW/OQJnVECzaK9L
Zs+PvLfxTuxOofq6XpFjCoerANziI+e7UcaJArjVitY=
`protect END_PROTECTED
