`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xcz4zshpm1LZqGQpTF/hh7Sj8f2KyVj5b6Chw7HZiHkPKODGfeZ1bYPIkAv8FeqT
4NK/VQgmSQ5S0aGvAZriQblfavq39wfyhHTc2zSf0vvgSC9ud5/ZJ6OpfmAHgAVz
bbrjE7KeHIpAb96vJgLJ3EoSleYKd+m63vcwdXQO5D33FEo93dy24lPxSk6DFJB7
s6i9IvJm75DYgi86AhuP9zkX/YY99n/uGWSLwPR7Eyg2jSagS6NA0GVVfG8xgkFF
YKE63U5ZwxzUnubMyBh19f1OAybWvVbXsaQdoPqmuO9AtWafTYxFMFPeSgn+mPVO
I9bG6WCr3++pQb/nok5UPQ==
`protect END_PROTECTED
