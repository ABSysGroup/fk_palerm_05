`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ke9Q/mqnepWBmLHNsSmF9RxfZTNIK+l8q4yaF4enjL3PtI799+42TCAdR9v/d55X
RXoh593bs45Ft9JnvucTu0rltvZZBpnF5mXkwhOnvxAAwCp5eJ39WXZywxyupjT7
lAHR+R+WcFHSOplVPU+oQawnX8ZDWPguKqevLg3DKStLqCuDHRIGll7D35DI/mDW
bdXTg+W918EbuREY2sTC2MO6ZKoFm1WdoHy5nlFpWYZnzXwgsaz9MYUFMKNqYNYC
7Cy//Fs6E0U321rvhcaXWMjAxOdxmwu4RNMyzfwUT/lsacLqF+uUNtQUVyWbCdck
G1/KUt2ppJOUH/gkjpIW81oo2vsuoZ5saiFTXV4B64vW8BUwZ28sh3zl1/p/wAuv
yq6aswS0VpD0KejxBFMaUjfbXOw+q0IZj/9FRCQ8CxzmxbZBqUdtyGWhSzsO/0Dr
TB28tfaZEktQX/dpGmkswg==
`protect END_PROTECTED
