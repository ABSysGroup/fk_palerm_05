`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RrA9IY2jwGTqFDF6SUdXPe1MDfKV//DIJo90yYcULAuJAN+j36HwJGPsZVlRuO9l
AvDPYB/KFcJln0YDgMad4hEFXccTGKpFQuHnwKFa3bmSOt8n9jN/+eTarxxCtqrB
rY9NsXTvg3kQyBDKC2Jb0qTVgA51UzHEBs+++gNHmIybwu6KJnRQh8bhBxpHOjbe
Nk1/4d+jJu+KZqOImp+spA==
`protect END_PROTECTED
