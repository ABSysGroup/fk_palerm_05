`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FmzlPQpJguc0e3E48OSKHd9QelaPX4mFTM4NozrKJlqpGJ0oSkxkxJcRb1ZTNDBp
G+VgFpRfMe1A45cAw4ZD0ymfBsjODAtpoesN78kh3wf2k+uBSdlkCddno5sK2L56
U5aw+MO2vljWnGQOJEh3L34fZM10LdpsK7+yFpYhhhGjJltPR3xPkYbzD6ZhuKaT
k6ivkWfjXudsvGbF0nVvEN+8q6NcXlqq25HQr4Tzsdy3uUXHUQFDdTGCX8BvmHgS
wkIW1HNMEfsMZDaX+17HZTT7T12aI6KSd+haT8pg8z0H9ErAVXuMoq3buKPW2mtp
/6Mfy10HkV+V/OLWrnZoklZMLH6iHFFxhz4Sgzti+uvAeJCDXANP8qpNqmuaHEzj
+1nveZx92mWMwLRv8gIF3z3E1l2WOxp3QdttORATGXErsmKK1zLRngCb9T3EE1Yx
U3HOZ0fY0dZA7WT9M3/wBM375HBSez/PEs0JxPK/C/axULguYqMi5q1OPZfqcAyg
AAm0JdbEfm7mwQF+9NbUGiZCmdMNKsRhPweuPT4H+ypfGp9uCihVbN52qwSo2VJ7
14O333V+SRKe8+FI3HJyqrc4ufUDFpjpG1EokaKXLsumQd/SVzL97M9j0pxLLvDH
HcOgjF5w9XWsqcP6W/JuJziLnmFLjAYxza7dSkrn4B84i1/ajzW5ALHoBk+G7RH6
+ZF32ja1709cRXZuC62+Q94aXNNioWOua1BO+Kl4/leNo6QU3wEiia8IbOJE3UPK
Yi7KEvzk+lOKWOWnYB7/Cxqf+oCCxlBrujfdjkPZR3MKfL/lIpKUNwQN74WqBAuJ
o+VC6j4Gc5w9avFnKwC7rFefvS4wwQFrE5o3EI5PLQ+GAxcMAPUZ6+cJ7NTswxwZ
cBaKMjkD0oJi55lFToXb5ZM2Fr6Ik02VS4mHwW/65zin6GqTeTc/eqWJuRH3xkAX
3ri7P93xp3hfMTq3gnIllONsgRIrdWz7z9iZ3dlWE1LtmHbUpBBC9lRZ1++2R5W7
3JXdKvtn1QqH0GmEefC/35465RK725uUpNrR6e6tL1WfWvI7mTvdApdSFC2bLEkF
fCpctFCBBs/UijQBtbwOD7huTz2co3PxHXFghjDvCMPSWCl9Fy+dH0WcHaDo38LA
RACYFTA3DdEKrA9GQc33YNCVO9r/INgmmaUWchZlqLWtXFCL0hkllwySimgoA3xO
s8E9HcXUAQO2IO7ayc2YGez8PSHWUUzUjuyHDOYUJ1wBZ2est9Hcucw9EK4dSkxm
lWJA6l4x8TVAFO1y8ts/aZkK127HA/HvxCaGeHPH6Ubg7lbhdkFFMIwIhPouqqMG
lD3IpLmDv08TFcgQUca43rrtytLGFcRGZf9VL3FlEZGlWMPgZ89rGYebJWtBaOOM
2rC7CP/+IekInPqeYW36miAtbR5HgLWaLjRr/x8sSLyLpmL7YZSfGN657UWdbmJ9
Yi/8iv3PDgE/qLuFLUL6BG21l6C92xKhDMNqvaBbB+AQyJVRjQRH8OqgwTbf9emH
JLIPEtQiiwoSkQLewSA8+giCkvB96OBIKNtgwdRB9oKvqPNu7GjLR3ce5MepWucG
ANpimhgoAh64cGl20bmT7XkaZ2TuOUXy1kwoAKe87fPJ+RU+unSEUKlvxXQBWByT
KbJZxiTl2quGcOJaVcwSCZXOP57iP+ZRu+gO/H/WfDAkSiJRQ5mpC8quA7cl83je
4kHveAvrpR5NGS/m8KRkm1SCnmqrl1oy3IOY0ZgmqXbXb+Yr2e0URw7c8agOnmFb
8THORbTWTD/VLjD1e+eLHA74/G+VGtsrBKYBqJjOxGPoQSlPyc9kr3hvuhZSME0Q
/ILuk4e0bZ1Op5D5xTi6Ud3d2Z5Fkzeh93tqux99wzsh7KPf5VLLHu08MSUJ42N0
2Eyz7TOS5NhG36hVwOpS78oXRgE2SyKaozIcCZAjtNfUxsbxOWY+QVS0pGMGx1md
Tixp0cmrQ4J5D1g5K21/Veow9wJvTmwy2bDzq115wK7WH3QDFXHcDY5L0qL4v35r
VgKZ+Ojz/qWZfnZjJUKWClSnU370bPdx58z/cLst7zo9c6wRQMWFdARZLIFiX3/8
KRpm+GdgiFJ7UPJdyAOZWYaDKU8EDm+1Go4tTU1aI3U/MXj3DmF0WE7QVPPBDml2
t8cqV16eKGQPtuJWKjLiJeSlYRAM/RIDXg+LdOIkrbz1Ybu1bm9hkwsV1BLY9Gkm
p46s8i7Fd0FwHuZ8j2eLtZuTpPStq1wKeHeh+5W6Kej4AmHtD0K3aqGhdqRfZgJG
CZEfO9MfYWHD2dpom5vDj6aOTazg3Udno2893PhCP/MWosA5G6SnfwIgwE0Rccp1
mECp1KnQ56+rsQU2iLYK3qt6DgUULtbP1jAh/hcOGmQ342K/kSYh6Jd3qrrKKOkC
2jA5Mv11uiWdGGVaVzTdKOIyT8uRnCzSyhILK9VgocetPU/P66Jk+uC40RrSPrq/
QQjcjQgAhOoxvygDWkez5FBGwHrMX4BPgLz21bNUAVBzaznV3L9VBr+j8u5U//uh
KeNY9QErwiFh7VVmC+HNYcvHoYpH276/7riAOczaTrkVKZlNdk6CLNDNgMqhGdUl
8IKSMu8PuUOBhHKnJHUZ0vD6IVWv+JftoYlwwHjPJd9b/jdXaaEitr++1Zdfmkt/
iGzINw9VYOXZpGh9lebfrqCRx29ULKlgHazepRnF97cDxJaxiHuqZLhe1xMWJnfm
yLng/CrL5D/Hinh9cwTeDbYXC/pWSni1HS5jf7yBmvHW5mJSWmPnLA3UY/sZRABC
4cD0f/s86uAi6jMXgtPyPbYZ7zV9kjEPdW6GxB3XQppK1Icwqw94wURlBMhW09Ag
/46Kg+5Z08L3E5ET7G5MC2n+j86GqV04R/eejCYT4b57SIbdM2urk+eUpZiKIwvG
`protect END_PROTECTED
