`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3eYiguYf44cYI6Me0Umk3hz3+g8Bv/1cUaJ+DhIPI763ie2Ezz+2jd31zp+xR0Cz
EV7DgR3BrtZOzsOqno60LTxXp58362ysVb2UD63lEh4RLj/E1Ca31kyLpOjq05O3
VnpDXXLHL30/P2KYX8izJl3TkoGtinmWYQhQ8oFjxw+GL72/vN/daV/wAgsKqhOD
ZL90CwF+CQlDUA9jUu9I5xlTF6adXvnKbkfYrrzw06xeSgW7gXmVm4pTXAytDwz9
X4x7t/CmaQGDvw9hHoBd7txYl1l4UF1JCjRmtpUP61U+reaAsadeQVcOYQfI14/9
ZwPqJdlm0Mq97xZ6NV02C1OgsQBKaIKubw4xqqu21lWv9bv0I4fokM82EIcB5i7T
vy9pLlLDs2ixcn5TdGzkFFvY4sDjBxd5mL4YaFLyMkrTUTOBMasDW0bWz/FYrtCq
V3h2E90nHHJfZb48rbgHhrSe4Z/sD78fu9SrKdQFiNhIf0TO2NiZ3MG7eKMG47fT
dvh+TKiMWFHlKxOvETALQnXbGZOgJtiv5SQ4+ZWYVn4HEfXR2TDzvGS15qg/JrLV
Yq9jj/v/u2iAWx2lwOYgGz0DoeJKOtJfPeyRJ0eDMHOqnaIyg4vqLpgLNBMmhrFA
ysgwOYh/5BHuG67oCA6npw==
`protect END_PROTECTED
