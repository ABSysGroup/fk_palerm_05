`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k9s+ec8mXezEkeHSf14d0jZDNdP52tOE1fqY0MXC3BpUl6WwbFoWwsEt3dne4QdA
bSPYbQOOqUqrG6o3DVEn0Izucy5VIt4xcKDv4nr/uCSEFev5dHpfdzTXs1GDGvGO
CRr3FBuz8aG4EWL+VK7FtI5dc3su2nDNTCmy3lYqUVeN/jf9oPpmsxyyr8gymMYr
anBHrx9oTOjxE0TOkTGgvP8yHZX2IBoHh472iECAsxHDHa/+pY/YKnLwmn4ZK687
RgNRfCFB9EHmvaZpUjp7gAf2BARC0P7nR5/dKS12bIOQm/MZOCpxAI9bF47d6zH1
vTUksuY6LBKDtehArxFnmLfwrSNonJmygLMvMnpiIRn/7CwOsqi1GeZI/o4lwGEd
iKZeu8X0R8v12J0gReTKo+U3nGP3Qd/fqXg6COsBOPKkSfQhiARnrLBFCaGnQJqw
`protect END_PROTECTED
