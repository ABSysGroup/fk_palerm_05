`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kfdMRe59n8Dlr+ehWOveJFNsgmhhkG/tSc+9Bh80lSxlFM/N8QIIJxXFe6DtW5vg
FyB1+ZL3kHHRmVJaW0GyXRde9TvuwUQEtUSaxpSO4eAyZKufKpJOuV6JQCUwyaU8
6wSpbVhDYXuy3k6OJac8SMxjB7xgwWQnMiV3dKJiHANlKS4BMf0dvfYB65F8ZIY6
vfyyacmjlrZAAMXdFib9CsYft/WVE5mxno9podzNd1Q/SrRWoUOxwg01aK05lFU1
mdSOO2IAUdGal0YZPEg9/+j5oa/UqowyCQ3rLLesI9kCSx+obvreiW3Tx9SUyVJC
hO5FYJnxK5Hh/HEfiiI/q7U3Lpyej1f4Rx7dky3T7CJBtSt7wxFwawHB3qLgDc13
BuKN4Ty10LC/9ktmdHrkDH8Osc5LxYBP6erQe5ZTLem++xDAAZJSi0P9wMHH8Mey
fntH2JT32pyaBvwUTZOrOms+QSl1FP5aTr8znNxCRGZXK2UFd9IvRxGqyOnHdeAX
`protect END_PROTECTED
