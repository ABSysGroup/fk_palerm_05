`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vanPCk4vwP6/hjbhR+tY6PBW7elK538ehzof7B2+ZJFZ4uFvLA2dsJAUOXfrXgY8
QVv/Lrs68qAbtnNSq/XcmcxmgT/VW2L/eaNs230ND+pN/gcHlyE1eBLSWmGVsg3H
HveRoBdJD9+1KDsryc8U2liS3yqFoxR5wWxgqcN+MnUT3lkhUxFOL+ON8j+GEjsu
H8fOTL257zGs3pkfU18qRB4BCi9wYpMSrCctOzfhgogwDz6lv8GdsyJcbwNMwsuS
4Gjh8p/WNlMbx4BNykdYNX6+XXOXEtUq/JL8xEY7aODpKYakoZGYxMUJZBy3fng5
TLyI4TrcmSLzog33belfEJjkkFOAtdtU2/0p2Enf7yG69MQugya9muy562kKofPN
hl9ySwTZcOkb22T9UW4XozXDdb4qQggJws6jwfNH0XIP0jnEkr2YvIpIpydleG9Z
oCyLVz6H/vgiRgwWvzzMoj1toYg6G3Ltv3aP8BumsveNSdVZ8LdUSUn5PF/afhi6
4wjqLqTP+ITogGwVgPr2m2dvH8pXlc6Ju6Y5MTtTfyxK9P3crTRZtWN8zbcwxtHz
BA5cvi0nkxu8ppdh3RF+O64dY0YQ/I3kmFtaw9d5sfyqAFr/bS9eQs0vxT6/mBn7
ZSSygammO+FRvkOvdwnN3VWdMQsqtO31fk3b7MorX2fe9fmQsPzw1xw8LBbb1G+w
7N4EZrJtLdWL+c+daEorcg==
`protect END_PROTECTED
