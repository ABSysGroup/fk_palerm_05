`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YUS5rAzlbkppeynYfCqQ7oR4g4949l2UIzRLopdvIVafMopM7EcN3EHrjg/d/ogH
wiRWgi7qP77xaf1A5KEkd+Wfs65xHGslyz82hL46/q0I743wEexARgoJW8qFl5L5
8DFh2vYDAMvaCkh31acRcIZoX/GBRDRUJ5rM2hXlHaPZkWXq0ZP7/02K9UOX0rjB
oLx/nFX2B49YtGtRxHyGkWhhhvtg/0FK+5QDqYZFfXk6RtAzbK56b9Xzqu9ktsSI
0fKfBpL9Lw9SenFKzduAcXp9jIZc6PYL2qFWTlAA8Gol271IrhT+ljMDFZk8to41
DxCst6pDYVcQlMJTVDhJIP4+Vz3AYooAoUEQelLBI25k6tWgp691QxMA+R2oigtM
uiNF7rpWZGN46H6GY7rxZ5+aDVRUzYLaNW0jbT0C+vXIWcYU8Xur7ocgNT3WX1fR
xn8jQo16egVoDBrYkupskpCSCwPk2Gz0N630UHcAQDQVBw6N5t8+bNWJkG8NUu6U
xM43s2CFKe5eB6lTcvW0P/p045WfxQKgzLPqitviRcMnktdhq4kAQ5X89Wv1TP+P
VrMDvFz8zmU67o1pH8fzWVQheRzXii+qh6XgmCcRhrHJE23JMXdz1Tu3YYy+kBNI
y6nhzgfjBhUyEMSsBLHA5euKLmb6Mn0fApeUUH5tr6hotnClFw09g6/fOxrzqN8S
XKwA+dZPidb/u5bvnBMfbw==
`protect END_PROTECTED
