`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
geVl7uJRo1z7YZaZGtiHrpD19CAvk+Dq+EsUD4S3zZ+VJs5oTvLTuXXQVDEoH144
LaqvynOjrWGm8Fm0JIEH0uupeAD6A+1WneASooqwYfQXfK5KH/8AOf9Q5GPyrdPg
ffPqYZG4LfzqJzHOFcIMCTHeUqXuDN2ofAF4oQg5YxqCLU3TFjJjW9zEQkmtOJm4
ZBplnbQubpT2hwbR0xs5kmljp6qgsviOEdg7zghRLTKmMoNZ3xts7k9C0PBwCw5P
Fkly6Qz/Kg/Ay6lBIt2Hfp03ZQJOEBQ7PHsme+zQNH+JXXryTNOpkydpXKer8czt
1lst9K+wQsbvzVlHoSd4h4GETz7IkJS83FBrxYtAP/0nZDVB+2kDKyqhDSGy/Yzk
zxsgafzOqmJ+McMDCPlibFPUFQBaaC4AWGggZvdwaWRXqcitaLxKPyla12wUXwwe
z+t7PaM3OuwW83tFWyRasir6DmDScfX9XzGJW8Y9jOJY70xXPwZnZ5ZU8Iyiiukx
bfYqrN9nO3trCy+YzUFEDVsiAKdWgGaB0Mz9iRVWBagOlICsAkqvP63sshcsAyo4
x3eTRpju74Qf0GaflcLUFNXHTUFyOUkoK0B3CHIGVLdpiIBdBZr4gYvwXhzbED1x
BjgOMfq+hmseQK9OypqSZsFqXlIkTyAFSUzgywAsvjSw1ZPwoTq25pJMH5qtCAGr
9k1LK9G3NzODJAe2OMOioAt7274xjLKwXHYB4KvgLLFWx3DuHheMTFL7VtUnx61u
t0xcR1VoX/XpUIep/++8uIWr7fWWyi/eiNsIVwGD6RE=
`protect END_PROTECTED
