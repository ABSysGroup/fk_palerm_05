`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C1FfRjYPJvSNqIOi5MzZcaj0hfYf37xWMjXG/7oRBu3/uQFW08J3I8ovTOoAn/gq
hWi9lJ5kMi5iJQvqyk2VozPBY9U9tj34useUwJBfL3bRVlhg38lqBn+L2695iEfp
r5g6DSGkv4c4sdmp3pMZ2MZxtlJLPUzd79fEJp/2Z6+H3tMviTrsRSLEsjzK58Bc
UQjfNnwvoWq9R5lwOSLJNavQrpWR03a022j3ZmuDRPNBQXPk1W+T4GGZJ3BawWJf
etREPMfGMMXikut+AmPLd0SvKqHYNO1sWEWyrmXv0rkXQccfM8AwEuZDS0fD2VV4
Va1o0r287JhGz8l52vN90w==
`protect END_PROTECTED
