`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QSeD+3dMHlPL7cXOGkAdQ4zRZQ5HxGvjKb3WcuTyhs5HVKFxMZRq++TqC14kxAWf
yKfKsGh7e4zlmiHGTZznbckUCTLvuVxnRkGjVzpgWfFbGcRqZCsvuOZ8HADGKjh6
tHuT2pLwNwZ2gWHEZTilbyEvRfiLFT2+p9bB0D6m+EYw5LFFlZeiuprDXjnYc02z
VZswObkTSzqIfzTlQkArAFdvCFU1pY5KOtwXg+OzLWF9FQZa+SHhpQ5jwoICmQMu
Msgd0yii60UM9gAdlhP7hyWF7+t/YGTdgGNzU89rDPyYNiUuIOkS3mybiWbH6bDG
HH9FSdE6A5kHU0U5ie90zAnaupT0bMF8U6+bShvDujMMNJHMToAKR7OZSHkVrBan
Ly9uPjj50wfNkSEc4djbvA==
`protect END_PROTECTED
