`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H0LV6doqvAAf1oorLBncGnZ9wszSRbuF08ZgU2YiuUg7cD1GMnbozC2CgVj0D6VH
8vV+SUKaPC0jF77OGGHkjnYmV440JCx9Gwvqzhg++yZ/OlGzGoiMDgEg4dsYU7fP
PclBz13gtwNNBwX18aMr1fBRTvHa09aGXzEggJtuJOxAzVldKimNsX/pd2U4I4GJ
IUqe1EFmUlH3y0ThXeaWNrFdWCXKbKE12kOADgBCmIK7j0LmzxdesNe6YeM+VpGl
40FtOqhDwqDSsIGwjB0LXDrZWwx7aSH9jx8aaajss8zTaRuGDy7jpzaYrXGqR56w
HAfnNk8wf2wfZ95j6ju4Dxn5OJN+smmNOiphXslK7fwPOqmS8t4FLyFtrRraTFKw
bsTVoKq/gbPH3+T1Ms359LJYN9+9LKALeWsD1WuGLxOTtMqaG8SZuectKerrR/TG
kuqIwh8ENzGFBvrmKCUHblZTwCkEMdtp1FoD5AuyOJV6wnBdgpYHp+gNFJn04E94
hNJkp8yGL6LlQOtlHVXERXx2r7heupjXo3CyccS52crqE4En0/FyZQRXPF7I31eJ
TdJ3jcMptnt+V87i+2Txqb1NbUmNyzbrFhGoWZbsZvQ4YoqNTfWVvpCDFwr6cyN5
r+r3LgnrEE6TUAHLOrRg4nDbxTDJakwkmg18RxWDmDtKPVmQO1W5GuTQpAATud4L
xbhdQtfiAXkAsEMsmAQf4lBiuLvGnF5pcngH7SoDxwJRNKcM7NqgHcqUzU8Uzd+m
87FxIHqbpazDT+U6bTXN0NZCq5+32/1K2dbOQIbys48SVnM4G4iLZOtIg0NcrNGX
x3+0Dze2YzJ20l2EOJcAHnpZOEvqvhDhnzuDshsVCkrNR8ImjjivqKq0i6Wg0QvM
b5tsGFAD3Qir4sN2fu+fjiEMpCM41FJ1WVtcLj6yCrUz6myrrx7P44Nbx5jxdqt/
apeL2cl5+5U6zqUMoaVKH2KKMLyLHNjEokxpEvDzd5/zi2Bb7lL1+/WJwwhQF6Dh
SoMrBwTy/n4g90/XwTB0s0vhW3h0KP0M/nleJCnMpMvmTYjTLidCvUmpQJi5B0zU
ejhkm+jCzRpcnOuyWf0KoNSayQX/IQUiwxxRrT3eB4UP17Nc6wUMVcDibb6m8Xc+
zFGEHmF7xoKNCQvWx7IagDnFbmWd2bknZyyc1iuSxIz3EcMOZDxozDtmHa5G9O3L
VES3MNkVKayLBniCsKP7EFlFMOfMx5E08YIOhPKSF4O79Ir9OJCjFOz2uyoUeyZ7
n8O0ddQtkqtC4/0ExiVB1dqiYZISq9WRJPMF/q9Cv6qJIIoV2Lhbz7eGu634cK/w
mv+sdHSBMN3TdNS4Da9LIe9DBbuavd2U2Kwa2GjO96ZHGOyovt/ju+4xQhtOvRm0
6dB7pz9U3tmlwEaD4tEAuU/HMpBsoAgp1hTvzarRe1LHbeeT/GTfX5gLywQPoD2r
EzpPHRQ6V46VKO65i8cxyV8mSMHuLsM+U7lVpB7Qm/msAhn5X6MKW7I7wn5NNXY2
uMO2Qi1uAij0oHkNoKQNh7sfyR91T0UkLmF4+S5csIkbzykqb8pKPXNMmI4nrveo
cL6K0Gpr1LcHEQW/M3+vfNNo/UagL8mQZLNHloHK9OTxCBnwQsWxrQ2KNBufuk0A
5QnjPJ2dnkpS+itdLotek3zBhyx/WNWxWVO4VnQKWByaGfELK1vhoCNDtfk5BMIk
iFqQi6Qk61vku3iQIz0rGN7xpFHyV3pJllw7NHcQ2iDpR93zo5CElyeyK38SMtFH
W1PNWzGy/TaSCAsBFIOOzgvhrEgEJnKFkVjQ9K+u62IOf/4SQjtXM/1YLmzGDG5+
sE/8mf5bTNNyv3pTERPRgTP2j2O34SfGaJB9oShCIgjqB5IYtc/wW946PTavBwEi
3YeqdcyCRhu8cP0mynZdPs8gh1DX98XF5BHRBqYqFqWUgW1poncVoUQNC+kg+pH/
frfTopS2mAEeQ/BqrYyUlEWq9L1kXJ77GszKRGYspLLh/pPVW/NYsr5S4ppaqvV3
tc23iN7wDS/Lu1PASd6UCrrl00qcjr9uDgjoDn7PJGFvHHgJourWsFMO0KugoVeS
D+ATXg0ieB2WEpWweONC354fFqsZGSvq/xrdByCed/jhEO1SnCuO2dOfe6VirG1X
ybPM10ZFbQGQwZIMO5ndplG6nrXngrJo1sNBMWdBZaGb1RJU40CGEoXdGdl19TCE
sUkR+BW+sVjat00lPUz419Fs7ciQGPJ2+SUzpAJuIU+BkIeziONuX59YOKNTwynL
9QkEyNE0LQUuWYjtLwU7bwo3ryUAdbRWq2CxnRRdJrwZIc7cvV9sftv5redX4G0N
CjyKhrqny583Zn9adp6Um1o1LQKNge9gmvkI5GEjAs7mRP7fI0JHSB9auLMazET5
zymftVsxlQpS0XUYq3Rfsy8yXlTcHXP/hW7CKhkDyzyM05pr98pdeWXxOIprcH3Q
ra6ZAeL1ybTy48gpn5A+FIrjTo9Q+0dwh4cKf/S2YcQV/x61RhHMy2jGcle5Y9Fj
mucazlwiAWjyExmRSRsd2kmRxt8S7KE8FePQZKuhcvbBkCOIv4nr49TW6XF2I4Sd
fb6H/8qVbjgNJZD5rnUhwe7919zzjiTVHmeNyxj+pwPudT6uPCJorjprjE2We0U2
Gg+DT/5i0mlC/F81Ve3frzBoly+nwHTo1CEB0+IykJtEls1V3okNcsFR3K1HCf5x
uAQZjicjRFXydUg9S1QIkTwDgPfqUWt/nszWELTsQO6lD5A9/+sAadmjgpLtzmDt
8sFf0LdAB7UZjqbe/9IVJXksZMBYlp0dByzefkpWbVwymIfGPRvpzTyd4vYV8OPi
HsAAE3+HfZTDvpY8hrbOAJKSIdnDLXQUtqV5elZ8kHHcfpdqv9ONRadT5cpZDP11
SKPmmZueiEzRPv5cXJ+/uJZPb0hNVfPUsyu2izN3POJOYuPiUL0p9+/PzBOsZFm4
ryVYuWjnHO4OCYz5IMDwkepc9udOiAEjtd+9iXRykSBeROuCe4nHHZ1AImuOUDla
a1B1k442r7WtXvUGjW6Wycx/I5TXg5dBpAH4ZMsSdAXPZbLDqpDzBE+CpA+V7ZGX
8MkAD/rdUYLoG+ElmsTLdF8PS0RXELs4Lg9r9m/urIQFqejs8s8OIADAHu+vr2iQ
yB4XaNnYXBzJtp9REaA6yKFEA1G6Hw3KUiPQ+RpNAX8aEeqc03UMahVIuesMGCs+
3vitUEeI2NvOCRXpWtAfJR7jZbsMKofYTPp00Y4tGelzavpPDvtstDootWv+upsB
AHrLyH0edTxxOdXJiGHtOthYNoXgKhhelUqx4RfVnKlneUPrUepnWyTXyytQvgFn
7JN6smrWbhSCVJJbL/4+TdlNz2Bs8o9AGshHBeAWZMRa7R5yI7FUWtBismv8sZXQ
bCHFA06pIKdS5WiI9y+x5imc8rb2aO/KJooPQd/rgkmgkFVwBEh+wEsdT/mwgz+z
R2krYDkpnQLYFue4xvs4LUKPQrAExqUzd7KYFYqr6imdtiwkj5V/IXWTgRwq++CE
pPEe1lIF40c2FCeV/ber3oM00S2XfYVqEmW4VYR91G+wBwD/E2QfQ7oRSUdGZAau
mX0WPC9/fUMCfCd/9PPIVexQkTINMvhh7Nn5bEXPEQ4StlOp1IzgN1tLEiM/NcXd
44eTAfVIG5cq71TmA+BiCWVLe4K1h1jLgIzd3frlFwCxOguGZ+lH2xchEeVcGbjY
oJKvQbfHY9YxLWNFH32SlHhF9OaE3EjayIZ1fnGuejjZ0YcSD3MtGnM3MVWqrxOt
B4qsy42QC75D12XDQxM3JtAuCRwucRezHOMCY6BJqSCZbE5u5GtVyGzn0LZ5HpJK
ZF32f7krnZVhBZB1w4FZ54gpaJeGg2XtR0lhuXc2kKhvXuAFBpX+tl1om4QYsMQ4
EpfBan97oN3tw0w542FwgEp0rJ0uDclyAcxH00VgCPXRyFi4KPcHhtU1Bn0EZiyZ
R7avI2Y7DrhLQ7gzHlO9xakHmd7JmKXO17xgxVzkFMPAacvfV4NWaZEQ+xajU3jT
8rXnBCuf9yyfyz1gYCSFxgoTrcuKSymLQKmk2QOL0iqmPQ7ma3DL0pH9bkerK20L
DJx2KTIG7FpuNzuwPfS9p7tkMEUWsxG4g8CQQFWCqbp6R+q/ElD6NHCljnX/Yy51
bvYoCsK40486Vf7lzXWzxmQsYzA2CRQZbiQ7ipzGvxQBEovaPDIvgbdWDEcYSkaK
ItVMA21ljHExUJw12co+CxcwVRSbT1Jm/blZTTy0JGJg1TtTrvPe8uIuGeVkS+uz
WMHiEqOXjLAIpQH/gSyqK0uKVtM8Wo+GXtxq0yjPEiTssWVc1IvU4VCW+Q7iHnaH
EDhC2nTBB0twDkLz1Us5cfvyO+tosAbUKdMiPg53SRBgoAL0atNWLbp3j1fZKhk6
Tiffo3tcxgSDJxJ9G2NDksen0ESXyrFFtfDE8GN/S8jB8r1NZce0AtYDRsuNKKyV
CAdNSmU8r+0drmen2ThPi9x7HF5BNhxM+sG2QoKMIdKa8k6OIVAZz8Gc0ej1V1ak
wRh06ceCg+sYZhIzc/CXQUIK2PsuU/TJG/RuS/m4MvJMfvU5dB661bwsnLU56LQG
1ykAqdSH9zL4zIiEVSMIs335UzrWk2cviyYuvF/kZAWJFE4W4usVDqAFyv9e2UQi
WAm1mYPqwYSWUT/GQ8d6BJQzGCUHdW9+oWm9QWHYJeiyCtdTg6GI4VJUl9gXnolo
HcQ45zX1ZdyiSrqJ6AyOIjEPSOtvicPdz8fGPuB5+3yI+nB9qBzuUuo/BC6owVoN
kCvI2S2qSPeKTmTQqGH6eP+EQTzmZo5yzn6DtBUdcI5XZ65unTSJy/9WSP+B+GvI
gJ7Bk6g/iRhgnRfbcbB+h/3Cxq7XTwBDZT6rmqbAxdJJySqpS296xLlwn81vhLQb
BFZl2dFglU35+JUDzRK0+O1oLZ7INrS8Va1fvftjv+fMG1KzzxI6rRkGK6DtunD1
mKmR/NCAOubmlGtyb+CpbiE4LNBKNjuTXvktqfuKQfIC5xMtELpf1dnTBVLRMX6h
iMc/Lrsb6nxBytiDO3f8pgnAmz7pvSxV74afZ4hdCm+M/NjmWw43hu2x7xtEl9Ft
36w8AjRw0PAMCxY8P6o/9pQS5Xx272HXovRuJpZcZAWs3hO+bNepLBnzZIux+m6D
RGilt/U860tciEm/JWpz0qP5wpNqM2V0AlhIcgUcFn+b2i+gN1e3I22fX4ivI6IG
jzrRVtYuwVCLyY1AiY1QQ2GacV9NklNoDCxM/MGSOc3nZs/nYE4rHaBY45HLv4eg
Te4jTI/fdAWPbh7pdhE1k63Ge6l/OazTYX6am0/7yYBic/tvd9QU7DIUpbfxBOiy
32WSKIm+XhoAKkYpv0o5PmplYRoO9QmQx8+nQy5bCL+CXtVCXCxdX9m9XXRt0no6
jjLUjiCBj3YE7LTjuNTNCDswlFGCBQkN87hAlJevf4U4sKkdvd1fUyNNhcJpOP4+
UHV8w5pfyg76HDyyTVMPvBVyooDcaXWbZY7j+YLdKN5qdkHkHLU0HwmeppTr2WGb
rlDRursVY8RPetCbvkMcUe4H5vDaT9ArrSsrlRHlZ09okoY4LfOz00gHfiAS3e45
oHTN3a2DsUgxonUhO/Q22bWXpYREses0kskV7e7liRCm3CJ4q8GMmUjhneD7sGuR
AlFra6XN5y+mptp6kn2HonO/eqOUfPtlO6UcIUmSRIXZtWNeTXLuK6Om2WgHCs4X
HFqfKMWCbTshJEhDqE9LERzliePtW9EntwhFtRfxUomOZWXI3xmO1eF9JnOLDkDn
vaPp3xygVwEzZiG+DGDUrTJAX2IGSa7enKBPvoiaSJEvzCOwJNE63bfFymI55TNi
NXKO3O0zay5cfVMyql1WRaPPsVfM9NjCPw8oJUlUfg82zaeNzPC11R9zwOKohAQL
NGlDdHWYRFhpxtAzLHnqK4vIJCV9Fronx9pcRmWXgF9+xmPyRoKLn5FH/mHMMgqY
cVsENLY/U5b7k56A0OfkPR/9T38aCyxNGK480heWvF0oOZOIVmMpAndvkK+3uTUs
vLG5JnfVJ/AkKtXOOsXh8TGvvIigZomZ2Dmp5+pnLS8xQ0xuMfspgm+m6DS/j+iy
8rgOU+WUR8lM/wqUwlfTmUibn0O7luNwEI1IN4U/KDoAQhlJU8+TiaRQh7OHjP1s
23LSQ6oxT39xqbmTV6V1wT4G77dul4SqUKh3nz1wmihxE+kD4TgKD56n0tHjxI+8
+S/Bmdo/+xTyFBk3l0aTGaOz058eGGaN3nVDvXvFKXvW3vHh/odyOZbCDINVOTe3
f9QZRWFymqmswPzJy4OHHrVRZBYZ2g7fTnCoWk/TOd4biyXjyXI2NxrCt9/xhK2B
jESPuSDx6sGQJObUL5Ynb9KEvAsfez6TuQJLUrIzFAh7pXzhi5rNqMAQu8BVoYK9
gRCsusWWlqwzUmtPzyAnCjmPf9K/Vfqg5kCHBzvBBEiv3VHnnJVvv0MxFU9tIEaA
RNsFTScaKpypNrrjhUAI2fR63WylYO/ccpyTswerFxUBfkpc0mi8qjzcvvt+96Rt
lCWqzywEUmjfzJGVz8JO33lqAFkyPwoqoHn8NeZf+rFWwkeaHqWZsRoSgKI3bh4a
e3jLheGWx0a70Lpqtefgok3GwwEy1mMsJ+8XVBo4iSvFkW2o4O32QAukJG9pMzI2
LCjNocAtTN5WaZ9XyWxrZ7lpi1Ch7hn962rRwc0oI1fNgOOTv5wvLWmALAIOgJow
3gxCnAOpOODjJTH/cmfC3s/nkPRxhoFLqN2SgQTwApWajNvqr71q77MwSQCMWyzl
pyQwBOqjooifhhJSAaiBCNDD6C0gYZ6+Sif7ZzqwmEEKcBQH7EBxs660TWRLP6H+
cWCVn+QhyDaKisRXI494YePpBELpcKq+OClwz/pkdt+uDsXXA+gGs2sLLURlH8bh
s1LCRT/7p7/TCcPm1bmDtyHkcYHL+hmzs0IfpLvOy2xxF7BpBtpm0nxlJmDLz4R1
kbMUSEN3G5uc6VBIiGsmOBOH9J7D6GJuas3z4nD+ajY6JroMizSIVIVk0SWnBfQT
glc8w5tf6sAUEoaS/tFXAi0CVw3zNdL/m6uriXhOpkEJgnNjplXXIHmZhePoFjAq
ly1dqr/JdT3oymb2N+AIPNn8hlpXllAnq34pd8Bk0MBygwSAcegWVoLvreT9xILH
fiqX8EUceNo7hQ4BsVhscKpjmRlt3KrFHVKTqGudZWlzwgvNrfzTLD1SPMpMSfre
HcRIux+aapeMEw18lvYv1VfNpi5OOlZXHyVZDeatx3GTFMMHVslhZH2hKvpl6xOH
rrcRXt1Klb5vY65Au0Sw60qsRXZzg0D+FW8CxO/9Ye+89MCuKC0DHyFVyCfTEO18
avMGwGvBurE5Gt+7RDT8DGOurFvS4NE7s4dDMpMb/RioiuFzo9Pv1PGI8QMMRkiu
xXeYhZaSVqIQsvUHllstMCw2pJ2oryp9lhJWl70efrOKWT65DhQDW1U0aGgg7PvF
tWcMPXM6ImMO0yBJloE6NGBAvHiAkeCxoUPnoFjX9/uxd2Za//m/UwWnbyz81wOe
77j+rkFW4DnpfCwgl/eD6hAbyvp5lgo1ZeWWypUwvvmXn8BSTuJD7Hoeq+KfuVQt
xJ7yLYJRTt//pswiR7YnIS3AeQ2QvsX7g42zY1Ya07GCfhYg/l80gNGcyrkeqxkU
4SAWWuuWYOlsrjqgiznFPfMTTSOCNZL+DAQcllnofy53Qpw0MIFxPtJMUIJv47yI
MDcMdoMNL3C4FuOjAYlaObx2y2ZrkbIlasCEKGLfQg8SIWxpgOgsR1E/nXGQDT53
ep8NE7bTOrGsVONRMVjnAsgqLzxgcPNWVYAXLoi8xL5mFZ/Nrjeew5QpEuWABIJK
MGO2qkKrJgRgs2Q4/aqudcFRNFlXUdFVM3D25f9vrJ7+CR+My2JW4tnFV/t+MYMT
cpnpKi3EqfdptyWYKPaCmRvQzBxxWRAW/MEoHNI4oPd8PcXOU/pjMelu4o94R2er
OjhNKBEgDosWy23X9Arhds/WcQ/BQQ1rJG7QK69ptXyXOyyq80bVqeFUSwk8yVva
yRwubQeqQsg7RznSt7oVRQOTVhlYLb/mRuh1nWODdM1oF6yVzhkT0tqivzm+HtDq
UE/7rSL0kRs2y0GUu7VU7J4SWaFI3yMU8TiIH8dHF9y8hUdMedPHX81/pQNmqhHT
8qT5ncU65mRO6zfS3up2104bFu0N0YkcS3M7ZmF++Wk1v3IZra+eMhtFZgOCCNkw
7M0pVKqT8o6XU/50keAI4eymJCp5mJr1o2173OwfKqa4PIjot5x8kqzT2Op2PgZE
lOh4lMwk9PIrgRAS9biiUtiYftydMTdiIEKqc2oBHJ18IXAqT+pT1p5C+ZtkFgCv
2IIKjerkIrVCh9FPbU51c0pHMKT4hozXmPtqbN7xQoJIKpUtWFTktnfndc6mveMc
qMOTHnVTr4NOvLkLHEpaTW8cyduzhIWm5fq96W+1C6474tTz9JldL1glD7e3C+KD
9OvLFKBHlr1CuAIbgleJhEsL8U5fqLRoLtd8Z/XiN/QLXddUEBatzHYFQAROqqIu
zx6jAB8FDZs+VwXIyO/4Qb/zb9eLUBU/2yZTC8K20plhCGREJ3pK7YNzZNH3HXFv
oYqO+oLjSe9INt87Vt5j4GcAJfxej65SWAO0HnQ3Fnc1L+Vv/bjlzHPGw4I/foZm
pjWPDx71W0PQ03Xm78qAXKo4fHhyaZSnc4+L4dRfOiYuo7+t3ObpKKAFV7Ntw371
hsC6HShsk7HJA85/x5Q9OfzVp2Eu+DhYMChv+XbJ5T1BlNAgdgUfm+Tu89JXQrVQ
gQ4eDM5m8PjCM311jwthhHgPrk/2msJejzUcwKMluhIFTmQmp1p3Dt9IGswa/OUS
jA7T9M1BWIQgPrPrLqwuCXI3K3n+aWMv8APfWyXYa0Czr5fvSKPOyG6goajOOh7M
JVyegSaw1mkWccP1DXS4vKFUCsYCjmJo3IUmCT50nN/nGfXC7OS6i5Lk/+UYuRUr
COIBiA4FJFIAf0isNHafVzobpnvVXRaSQS2hbz75kBCRkXWdwXQcy0sMA9Zoc6U5
Nj2NTxyz5C7uglKqPISlweZ6p2H01ZkZRUvClSRjv7Q5blzdT+BiMM+cWhLIPkZb
hLgsMZeu6Mex2yTy78jCPdGMrzFVBZn5HSs3JsFN3MM+Z/xJrbPxLXlAmeu4vCmV
cZChfe1HPkP9lEubzfPdGa7QvxgQoL+tU0dMW9vWjA7t/bYIQyqJrJJ39km//xlL
A6XpCxa6pcartj1Rwju77QyA3JDi5iaUFe59ilSZJiS7xKL6LBGB9Zru5G/uFcH1
4QtiXsCodK6bOdvg55phfNiLt0T4FjA3wmrX8u5HWPk8CpxaGetkQAAxQqcZUVE1
WscTSqQ51FuzEsqUvI0i/labPgh2bWU05WmJShPg/skFB/ckEFKLUGMuG0OFId7j
8QRViqZc0yRWBLG32Gzt8aGrxCZwJfPqFT4DzfZbNPmV1e0jBvOty4GUXQt2XMbs
xZ4UbguJQIL0LkcfOSvJZgGCcasIgNc3sAXUgAEAGR8rUvIknmSdMGEieGnaXwng
Wum+Ox4XtFBs70v93HsbQYMdQPoJSHk8GER+qv608VeeWWGdoJCJpzEoo6FbDCv4
GNU6YeF5IyhnOL4d3EHC1QWtiML8cE/9jqyLDmObtaNGFEjZZGb9Kp/ZXdV5p9Zs
OynhxjH+XMnQxorFgzsmhOOhXbk44WZtjzqAFMYTnFj9ExYtm+RW+tal5cB4j1lm
K+1azXYCoT/KVXGh3Mjyl9tL5dgvPXi5gzjYySSVW/L5WqtSPNaW9CTK5BdBU0vE
qx9TmzuE/aAvMqckbsdZ3QukiDfPUIR6BTIbLpx5eIksaYYguXFiMyu28beyWjgm
QhOs10F56XBiK3Jd2az/2CoxOgzGi4AOOMuCjcMqGQLruot8eN0SgVK4s9Rf9/Li
ZD9mSbTo6MGvNOAhHRUI7QMVg2QRBiqd/kQzrOMd/55KwGwybE2tpM/Aj0YIKwf2
dXB9xnTmRPltqZ/9CIbTy8fDkf1DEiMZTddiLqsgL853iqpGA2OCIK61jgb7elh4
0KOkIN8uBf5XbBsbdOx4gcfK7SgA0KI9mk2LZrFuthzmq666K2zbyC/adfSEhcX/
7HgbR/NjJXuj0QNG2byQ4za0l1bQDTe+N1UcUuHmCaWZ/pDrqbo/6wOwe1KiGwp1
dltV9w8NXkTZ4+Dd53sIYD7TX1sHwDk0QAq8PgTJQpvL5PMXgvNW6YRiO08u1AlV
5z0+4jIMUQmTbev2HQxcEKN/MA5zsgsMsjFqXViTYoKEFi/2yEpMWDTHcreTYj6K
waaM9MdiBkv1zY4PjFTlZ3knS8ikYDcYc1nSzfAp2FxwqH3Iwr83HykpI7CfdmFr
qB1Oo3kXoXFlEWUv3DtEckS91Fm5uSSCtIvdTKH7XB1DXCMMZ1pdoa7+OuZcQeuU
Q3h0kWQ73VmfeNjk6ho7AoCSGZLd9Rewf/3Cd6XvuJmdoyN6yr671Os6DlVENdhu
nlCWroohFwHNMEGISq0OFav8n5Ex3PBzOgeFZjSMYQOj0i7Qk9K8x30mTO9gPHSp
H6Snbe+o5sgch0eZuytxK1uOf6cq4qTV45+FhC7s2iKaTcMh8dCZTSMtwtRFmKI0
DfPOhh1VdvblQJktrEolMfUTEUFKctDrWsh85TlsPy7JA/CMd9q8Pps4/eDwcPVz
vcf+6eI6jqv6EZ19AtkKT3PtPDKdeYTIRvSDkZtpuQZK8sOBep/K6eADeteG7J1m
xMGoAs0dNftPbkmsaY/kbGqR2UbEi1j9c6gB2WV+40lutyFW1K67a/e4SP4rfB0T
j+uw65BQmbyAPMUHk+jA80HAoZONbpAK3Q3WV+cqWfWs7sJfnB37LzH6tECq6akP
S0fpbVChUI4xyJvLc4K/UFpQ9ukv1myBAlKDZBWub/xMK7u0p6xajkQJskFuUBPr
H4LV4iR4HZIJhukSnltzjKDB64yI4RyadjahyMTsDC0hTN7EMF+Oy3ZJYbaIa8ge
dVGfcoM27WZDVLi44m8Axv52wJLAByQgRAU36iynN31jUlNV8+QR+aquPvJvX50q
RKbcDprbpaonXYV31AaPZfbNWLdpl5jkyXoE4cFbKNIKi+xYAIM4aOFhcOYUxox3
q4ZiVIgD1vWumlajMwomHbjgu2FcwCPZr1mLwgb+SFAmfExeTnukvTIeZwZaRXw0
S9/HXVvziEfdybyiESTunAwAk+WtOVZjRwb3tDA+8/iEIZXVBIzklWta1VHjtpxk
H9f/4aXrQK0od6YIIlZaa1fuzafbS1k4EGWMZzee/rBTQvURVC0JFNiXRtfk0FWp
sZyryQFB0b+nWeY8AryFP911vNy7U9UGicEOLGdST3jVzdRygW4b9UJuPyZv1/cZ
+mMR4NDsWASe1G14TKE0CX2E9HTlWpe3+Q075XBI8wckPeNj2S6SmKnqy3Gez9tC
3LnFLIQEVyzT0jbOUHEvFHPdDJEGsejxNW85r7yrjxIDftpAKqOF0x5QkGSQUivc
TXv7RwD2v4Kf7Ljj+BFMbG2a8B9UAUXTH6PTT9o6RzjL9+bOWAdPBZU5y2m8uIYh
ztbnJblrLHQu9BMZ1k7hqs2ruBFoQWHqKkont28dxGE0FNiaAqyER494qQCQj4DR
2uma3mYRYTCd9iqDzzUeuNQjwBRVA8w+qzVNqceUyshlusb2+Gn+2pcyW+iG1RTS
h9ikbA1n+jPwpgJjCAOsK1XoG5f1/s34pRwCyOxYLpTJ7ms489al3hiB1fHFH+oU
tcS3G+49WXVrkcqh2PvEURrLWCBCraEX50WWz6Vkh7/kPVY41QPhTyfEdlhi0sxg
Ym5q3uQ1Jaj2cyFYWVmY3FjA2DNF3nWMPVI2rCSV0hiCKB4y7f8Cuh+1GO9S1qz7
jgzZLDW3sgodOj42+DLYTu4JO1iY7BO8YdMsbQg8LBPjVEixOdFvxYSbQkgmBx9A
g5HYbHyiKUeposNE40S/J7F0k1OIKk4izuADKoc9mtJdTq/ssELo3RTWtCOAvt1b
1RTublXmdcMwZDgNY0OJ2jOVq6n7BmyQipAIuXghEp75cVKDZ9QHzqJUlTlKNdxt
qEzNG5AbBzDUVLmS7d0GFZAXfk0Y5hrvi5ZePN4i6ctJ4VERBEzdRUZBahKIUyF2
2+AEM0UIfhWiC7oj/vivsf0sASM+zHbc76eH4wS7WxgLFZYGJ4Jtln0o4em82aqm
M4CNXbsXWtc0QGXx5byLSuG4YlQeMWK7ARTUm0K8GCerf9qW92MpTyPRqRHlHsHQ
87+wpsc/ZdPj184R2330GLdtY+zTtJv3oZxQ0MzRgdWPHnt2WKKNi4VrPUxALdiw
GRCQp6reu23PHSSEFOMS7Vc92tFFMPDWk5rn1dOYMepGpYX9cirNMyXMjYpo9rYl
F40tg6mraWU4rRXIuyFxomLTIUdQjATrZ0ioNngJFzS7PIWStMzXimWbJ1s7H+ph
yBiFLaJ+mBWqePzcweDuSWeNA4Gr4O1qTDFs5YJHDTJfl3tS0cTdci/XPJKmX7eC
Y0mqubJy9lujW789fOUciw/YHLviA/xxv4ImPJ26wfxVl2zKeem8ytzJM0Bhr5vw
9GKr452hB5UFoYnrgzUMGtGL2Ov1Mfgf0P6R0prMz4GeBgcYNtN/+7WQc33VL4ez
BexT8yS5DeU/Im0bP1rHsS7AQSIZnkFzQy26IySCkLtoFNoUHFiDlJ7u8Orn5M+b
b+L553ziCmxYcgSr3086dRZ5MH6rrlB3FZrwIp/CsdhBZ1j+lt5vCBeYJjkvpoTn
tAG2xa5A5JUwNif5zTwtemsMB+WJaB4iZrOpc0h4DtSjw+6j9f+SE8KLJF0LyyWH
W8fXeZkF2wzGrcPunohsPeAqJgo7aNi3gOp0hMrKpxY42/rI7sWDuBzSTBjC6h8e
VoEG7/1q1WadaRMSVvi9HK/ohmYSy/JMAOMBrzsJijaLU0j/RSc1w+qS9+jL7DTY
tk18XU/rMysRxClQC8b4KkjbDfK2nZYhg5xotfd7pum/mbGPh2SyBvMdjNHJtFmu
xKFgh4EFqxt14QvmxBz3jhkXpU5nxhTyHXp/p9++x4++WPprkIpAvcxwm61ODPgv
WPvjUsL2TIlyA+4JoSzHwmoSw1JRPTgwzxFy6/n/PaOUgYB9d5ulmItZkSvwU6wf
srF2Ggbsx0nlNa5b/AFQfLJwotvzpbpehwY17zW8NT4R2FBOLVPm3ET9mpa22/Ye
8YoRcbIhtfiijkzKbPHWP3l/xE+3ad8hS4AdmTxOH5CYd+KTS+OuZqTZP30iLcl8
HJsLYpl/3famY577OLiLXNMpdqHFrTGBHf59GK0W0kL5JczZgtNLcSWCVl30etzd
0G/8yh7A+0CXG4mo00VOuLDRHugS+vRFk10Yfuqe4WRrEiNeQqVJqlwJhtzMVOYi
eglUnvMunVSEpOoEuZBsf9BYuymym2Vsb/+WaLJwVZu4IBMoaGZ3FFYqhTD28TZH
hPOyMNIzt2y+w55vcalEZfh0yv11iBxEzEj6ssPg3U9rp6Np3xIJ0ZE/2lI+HG/a
J2UEYwDPz4Z2kPT0csLl+3mBw4ngIphCiCCwij49fXGtAd3l6M4w1raLbkUgeCGR
bmygg7IpbyPeS/xUtF2Op6sSxl6QkOH+gQ38fBeyJO3I8GNxP1TozJsaGkvxbV5M
D5qfBcvnvWDyIH8kpnh2g8owS3O4FZE7ohM4QzS8OKfjyIAFH9bWUOSmtMNe1vTZ
o9XFvPETN/y1RyWGSp6/e7DF7TKqu37YQTsh6LgQfMAZmoIJUSgGiLPQrIetzG7e
PJBB9lEkNVJ96XgY2iJLY2my7BD33dzU4Jmk6KnfxNnQFtMw8B+npCwRo8dBXYg1
1axtpdja4+I+sqS/L2Ikt7zqK92Nvq3WXOIpxpj1+6IPJrZ4X+sknNCCwAfI7XFS
ayKwERE8hytMURrgx9jFgmVDacOJQl78ZPKlVvcPUY2xFK7lZVmnKh0WW0/Os28Z
m4FFc3A0go0J8xuNovZPcd8G3G+dcOn27gCiiAm32JzanvceJH+3psIORnlcvEc1
j4N2+0NGtXWUrQbTbjFRmWVkip4aMOSebEozoMqT3w+uF8+Vh6KU0sGwBQXDKHMv
IYdtlY8GfQ5TROyDqbSWhfBO8qZbvhvCtlRQxYrWrBeA0Jw/arqw2Ddm2weqFZ5g
eOU8a5hb/glX8zszVdoC1M+0zKCs+yYqMAwMdamTJFPDSOywtdzqPYOy5LwJDuCo
ZyDEfYlq5HPaUVJ/fTJkOkgm4XQ983KMjkJtn3JE735KAZ8C5P+rkvAzWdb9MTbC
Y9k1RLPk5LA+a7RE+8wquNQm1Ru1F6u/qh1FpnfDuHLw4+yqPCP32DPrMqF194yr
jQUEWgoaKBRWikNt3sASQbHUg+Co9L5ucrII/SLRqMYpMtPH4rJ5PwbxI3yR8Q1j
4YsoREDb22LctVBxyKUry5uYUEIApSdn2baNPVEJjox7fTAdOmoLno3EwyWkEVi4
zeK7BeGUKPvXJludZgafvacaXqH8RsQoD1i1ar4fVj2LH27pN+TTO0YnIk1bKoIg
zFrPA/zu8a+KC2DL5thLgtqku+HLrCKga4qkHLTgx/GBik1UcRuKm18R3D2EpJ8+
OMgvIKTFnaTmJXSkyctrNNDtXG5sSm+SRUhcAmPJTUW5uC2BcZH+aCCxm5TL+0Vs
zJIWkkx1l1LXael2TP4VwPFIMzY21CyWRTXAA7qN5zGMWqygE9M9dmbf5cHL8ajH
RwUVvTY36IxaW7I1VWilHpsBiNE21rZ9ioqp5IePfYK4WYQRqfLVTYaD+CwFkCo+
Gc2HoPiBDH6Wie49nrvjveDSt9oxZxYT81gSqKclLz9rdGnABunswSBqEtzu73i2
4yORCPHb6ax5HMIi9uYAWUPiXsjXoG/e24p8jC1do+xPo/csh22LovqXaPVN4jsf
ZhyOhI0lYPnhdKaD8uY2mCMV9dP6xDJrh7weJbVB4GwIX09k6OzRnkInIYVNQ4JB
URaPLkeXOrhAqczaP3KVJ9G7oo62jxh1MnZXLd1+TZPrCdBVt/6ii3ob3WA5Sazi
TelT5R+DpZvIuNjetZkqEFDu9L3vDSw2hrPX1yJDTB7/qG4o1YlP5mBohxho60TJ
A2VQ1bOf3sbxdQ+Qv4OqqL4q2VNg3DDxsp9ioGTlPbeAR5tj9wUstudNPsgsHPz1
F05mZw3fD1lNt9oj3Ep+YBjYJLXC3vUaI+zLkWTIeFvMKqSHfhcFuJ6tkjH/2pB7
BV6U6b0hKVYP+xBDhml7tbDSCLFFBBdWj8kYdG537jfuc8iY1ZizTOH3t0YCg6FF
DLNGQCZq5kFMkZYnKLCbHsIhNpcQfrMV9YCjCTUe7u3fXOOnVjnn0HHiQwQBdC3H
ion8yRFO4HjLRbzXDGU/VJ/IrLIcdy0we7lkP0y4IrJ8SMBkxJ+Y8ar0MiMPuVEM
OYAs0ti5nbTPuxSssPWz6zg8LjI9MS10/bBw3zriowGFiixEkYj2g5r45/2s76de
frjzgLinK54iC55xSNFvyRumw76oWCcLnEyW44+ychSzd/Dz80VgZJBYv0HcZqVP
+aLzpuyZJ1syqdln+v3PL9WciS/x7fIIGInllkaanckQUzu1SE9oQUQ2F3KQhDaj
Fm6ni2HyBvqZdFjkeY3kRqo/SIwkOfjs4aI6dKhGmv88J+97u0R/ScRzeNoFC1C5
K7Zg9wnvPpOMI18Tm2T1Mhe3LL9I4XUXSWSxu+8UuSwVVLjp/dDKkWRHF8P7W3Iz
qtVcG2ypajSxcBTRYYRdDRZXFWJmO/qNveTBvw7ckkjCf2Xpm/azYaP3bXdzGVOo
eqC2GJOD+cQfxMqAJcrYK2HbZlrVSbGFib1F6n6VekZYyVpN2B9v2nBhCHNWOar/
tOsE50dFceAb+4i90zTAg/QPfJdcuGqALXXl8FVpUDetwOIy1gm2TTaZbbSIFF4j
+neRYzM26DRXFKbc+5i+JpDN/npps9nJZsLT5aKmojQSGlN1T4Gg2aQAKFgITLfQ
WtCavKbbQKl9Jxyv1nE6/qFP4r1ZCjXOoOT7C+yP7BTAXyETVy0XfX7T2r0AwpPi
MtpjSENHR6kBNIwRb1qhuAm+x9gX7946nER4Lqfrd+nsZMWgvPhGnBDrj5s6pWix
GrhXqPCkBJKv1EgWuAAKH9w3kGdicTVm0dMvVC6/hCC5gsx2E0tDpWY4HGKVlU0H
pAXcWaXpdmOC+mXeUXmSRsQqI0oktVRkbBpi6b5ARA4+Z4AJqjPL0y+OMlmRf2Dj
4AmCIeZel6pi4ESFA69yKAmDBS3jdxi6GLXFqNIjvSyT5yr2+G/4eAtJGDTiJSjL
9cZTTecWVkM0kM4z2WHBI1YCrP02+rkIEipunrkWmHYz8KhVwSMZipqualxwDe4J
achTylgpuLpkZSy4s3V8srCuZiN/s2iwlEzWfq+udV2Gj0t/D45/WP63PKrTZKaU
4QNGDpueGubKOfMFwlCD+b/rhP95qHDCO5AjeZkbqB8w13S45HtTDfgARiZAI3us
1mvZ7SA6bnlV7YQWF033QSkjInLqi+9Gtq/dhnaJF4kpMiPCyDeS7W3U5gd7759v
iJ+Mkyq/Lbfa5Rxtwy5/0xyYB3EKYfn8eFic0iov5sVVXV37Ds3KKsAFWvdCVYfv
leZ0IBINAEjRgg/4Uw05LraBdGC/cbB9i8rglwU9/xmVoNkR+kkvVxb0EVKVruS3
c3VR+pB3YMEJZ6EvtROD6VrGQpkmF3LrGN0o9V6SW0Y5kJtW5TVjOQSgmOZ+AgEB
Nu0m/jzkADPXc5RPfR1r2jwgpWCfIgBe4FRR7wUkzTD7qBg9obmh6XGwAftm9COG
ZTksuphRDsRB0YCbm4b4OOFtzkk9IZ+PFeSN2igTXRVezzySaeXj+mthX2WVwfI1
mW+feu/h9T9N819e+wiX9r1gVDLK6aF+U1Zfbxjgq7QEN7Xhw1eB8hIlWQQbgPKz
Y2LFT/83nlZNt6/lnbLz97Dny/4Y38lhk0AOBD8xm49GTLbqWqKWtv4ltFHA7s3Y
BkXS9Y6r/R2N2sUybApW5dp3Lwhf7PP7/H9wPhRJjt+d/AKfFchuMQYKe/nT9oue
ZDyPGU+8IJM+0AUFwcW5HQ8FTTTZP4Y6hfdxB/J2Kd5tlka6oBYxrCnzQ7Ra/MFq
xj8X7ImdiZ+xqsT40pg4LvRMk7l+PzXK/QxkzZNE3yT44ER2Nppe/QL/+37l4+4i
9/3Sl+7j1BH6eQqOWzwlQFyK4cfgeFkDZImhf8s3TC+GHYB28Cpix5G/ZdjjO4YD
Y7vLxHYRi4OnP5oWPIm0WKe4qEsvbYsBr484qE6+AD+5IRDqAdNT+hdWux/o0GS2
nEkcXwZAjaXyKICkm32OPak1FbhyQRWSAKZRbWrqF+Jetr8zxFSKT3p+Gi8c1xr1
FM09G9c3TtcKdR1zLW/bjq83DAzPjkAupKssrNK/lWPJrLEbQrFUKTQ3rBCXRikI
ZU+69bL7E7AMXqGacjgkYdw8i3J/I8xL1clAlge1vOOst/5WB7Efoq8lnRRDbuxp
uLkQLNd8mXJzhV4R33zZmuFUYKGiUbZ5ERZM+cNB6XGofuce76sNuOLWoy3iyCET
lAmL1HCgJLHkER7KpVJqnCP3kswLQQ29qGh9jtW9MMelFwLe0F39j9afNUF5QG3I
VOaP9YqCHgRPXR5r7Xvha2MFaacu0fQna1s9jIelhgEkEGapFAVfQcwvXud7D/M2
4QSikXNLa0qFT6yQD0LCwdzCNIFb/rewlVx2KoL3DLebP1oG9qci6LiPfviRxBHs
bziGjLI4L25RnGSFHWirnJTPKL4MEwmyufvnC0nR8+HGDALs2sgX6FcWj/3RX53n
3vQ1Z+lMlEauRV9B1JcnTWxL2Tu4UnPsrPBYkmSDv58jrnnt91szfIX69PfWaaEC
EkW9xlHcluIy0R/aOTUJlzkkgo9yI8fpdxpNd3q1MFUrXooHShj2mXgTikeWTj11
NZGEKd0R5QgORxm+Sy8MXhzRzupxSplir9zFanBlJc1gjnu8wjbDNAkEZxwZ16QE
nupIJU/aFkAbBnLUbzA4cS0bwFY7uVRx+unZLF2sBxzIHqBPQgCGW/dL0yfL5i96
YKr3YU6EJ4uHNkKX7vWpYV62cTOvlyICr0rsR1VbbZhs9eu/HrPt8VycUie4dGk6
Z+hX1jYkFxZg4jk+LhLuIaLF2pmT6K8s9bG1JclU2jeuP7WLJe2Is13LTzt3DBnQ
QiLpL4EDLMpLDlHuuMZi9dwDV+DqTM1Ci3bgIeUldH9EsBLTCr+H1cPOTvaoyyzq
2Rp9h9Av/g9C26fH4Xl7vVo3IGhE+afcJuVWyeRY8rMCPzb0oAEoeM/+MGJBjWfC
GZ+8qINggOBxq4/O3AqeICRsEM5iSRhaeyLXTsifuMq1stgh8K0EAsddOvnvWr8q
oqSLDFUrn6miQiQgk9R6NcIwUUobhZdeI8XIeGa5tdvNNevIWSgfM52u5MVJPk3Q
2Xfrs49geeZ+iEPqxuC/YrPUOi39gNLuToNxP+V25WXLUfPRZtprree4MZQFT7qE
/L1CpQMhBWEfmVbz1QgHXbeKdXGyFSfhBRjHKUJICY7gn4S31HJuC2YLuGBmSeBC
dwFqDqgHewoj78orZjGZ7FS/TFXVN2C/ZtKg6/8e7wP8ADn1ulxH0jSBJi2lkGkB
lywTAZz8Cs+ASn51V5HvY+KybdVqdrhsUK4Kqd4dwgYCaxoAPi3ab0fE33lKXccM
4jQMaS8srL9quj1trCtsRtEqAXAH1GxrtwH5SLeVk1FbMB5wjgM67IvgKGsg+0Qy
bAZQDaqFoISndHXAEU+xM7jfvZOl40me889MMmk0Q1+aDrBLeBMVAO+DrgKixSEo
3+lQJ1UlZFTvVXAtYz3o5Dq10HDXgJZSdsITJOZ9N+GSCY7BciovZQHwfERQtWF7
i1sqKjoQ9nQctLOfoDK4iD2TYkRQlNaSzH63ER7NBMC2v/mvqV8g6DfKgl69F6C0
uOdiDuprUSOBE9WwtxVi2kTeZpkH7M67ZMT+nsVuRunVm13rsk8+vUuztjAQFvmW
4rlN657mbLdzWZ5wlD3rKDu8cUGfRbmgmwg21LO4s4Wm0/GHv1b7s/cDT6+CaTQv
dm/7eDuZjcZK1JH6LRoN/Aer8z/TOFhhz0akmMxUHxa2ibJsTH8atlHJhHt7Xo/U
HastliDh7JCsxSbQl34BWPGeBlhjwIITjBdMMJKzEnxytU8W9CaGUV48GQO+95Kf
xUqNRYQjGDgB4uwOWntvtAdbLEy9Sbzq78erGRsLvbWW3s7TxPq6HXhGT2S9k0UP
vplhRnrJc97fBZQitiUmqs/2+2a2f2hxTHsIjCEZb+kYuLa0IndZh/Sq9nv05sGc
DfWsEew38ik0nM1d13KhIgjOYuh31wZ9w1MspIv2IN9PCXlGtaaDPrGkatXIDqY7
a/HjoDNL9kZf6WlRr9ndPxjI/ddWKDII+upsfcGlm6lhVhcvj8o6x8u9pN2shRZI
HKxe7MaBs62KG9WkffQkhu4O5cq1KOii75H1Ud1CIOAx0v34zoS3Dx0n83ptWKn2
rdo0Ck4KNdA3NWmE5GMTTadJep2RlV6hobikQKU08Dj2S9x7uT2rz+cT7kcI+ieZ
ma55j1RA0QPnLhxm1+IWKWy0JmvqMF6EVwIfqobiQgc1h8ZZVxNYqjEnZCzdBKay
PZF1GQNV+yN4Ar43FTcCrcl6Yk31hFYRNU0NsyeUx2KN0Apwirv/dC3AAfpitIXJ
wrWlKhy4VssSEUGefEoW+OJ7AUUTXIaOJg7+Fz5GTssh32krYVQv1vkijyFz4Wf2
Syrisy6eAL6hOmTlRwyo4aT4bscGQ2G7/GQwxEQHDFmJQjXAIT/bKUBwENLZy33D
QGCL6AKDUUNBARpuJcjZnP0m5I4d1hYZlOv+48IHMG5alzpiysfHIYdKiBM4DmGd
WyLtTgkI+iWYb+Lxy+9Olbg6he5BzdspFgnGmu7zMmrojPqzwXPXSy0wWwtzfZ5Y
TaaZbFavJbf3FxJAPrVbHgfWy4SEpVLdWR2BU6mnV+A3fn2By8pK7bQ5962WXR88
FAbNAXeAOMHVWv0Dsi795Sxn3zb/MWLKeEp51R5sRaj9aRCzwkkh4YFhpwFH1pCF
TPi9+zsFwz1Ei3dt+GNF1SflPUGO6lyNZsQv6m6Q/YgrLk+6qnqbidb1e+0YASNz
c2hiAvRyNLpkHSYOiwe+PCuXzSkheIPDheZ+SqxxMtvWnnAxMMr2w29q5vLK/TL5
FM6K8GO+oWJrtnUmgxyKFo1uqPSDJb8uVxIpKFr/a42In7JJp8AtWNFgAscbRbVn
+ChCODVxneURVL0Zc5/aY/kFwAQTDyHWS+Ddria3o1Um5aHPNRPN2iFiskhesWTz
KuqAJktQBzOBN0ERoQhEc/gDUQyazlVy7zOhDCmP/H8FSFzinZMd7e+ITscJ/aF0
6HRHVFQzIFR7Bc9NBFtAZJtnoyPikIj20ropwrza4JcwQNu9rTq7oNlbrLv1ezUG
Ab2WcFtZOZmcErQu4DAXEPlDW5n1tCA+i2uWfl9uAIZUhH5Xu3FkJHnMNwcXygZp
F7VC+qP/9be/M4l3Xn9TQbFxLr3S18qaVP0onNHS0K/LexkarK1yiwx5cYJIG8PE
3eI2iXFXIw5+0Bbx7Ni5qNkBr/P5bLFz+ihasmp1ecG9ZVBeiJrPzhKiYhwb7Gc8
8Vca9aNQEm4v46iOQj17FHsUvwEnfbGQhDFNO+N/IHrMLzUKqNitbkN0556o/P8b
Uf+VFfPCJab+4CpsvLahwBNn56RnkSerc1HhDM/UPqr1savvQal/Hvn4HOTv3lia
yKTJ/LA+7wYMt3eha4M/zUIUYlUmqy8kBCMvpAl2+viWHVSmWq6u+XT6N0leuTPy
QH9l5etdN/ZEBfdNeQAhmzYncJQTBfRLKTMGswEJ1NxN9qDG3SHTijZ2YMJzYMoT
+vjNrL9Ig9ztpDFRdWqLV+R6Y6+5Qo/osImr3gahtLziNuTGFg2QwGm39IWu3Ng6
JL6oD0twYSgzJeNu4FnjHTp6lpJ3wr4GzQv6aN2x4gKB2mqQSBfeOmNl4Vy6yZ53
n5qNXlvxniqBcuORCfr2TrVFG6Zjh0ydNuJx8SXa67CSjCxsTmep+ViCxDiQpyd0
JDJDBJQKaDkcq1X9/5XluHoy01V+kkXtRWr8pSjhKjp4QY/xzey0JL2q37/8LkdU
aAMIdjKUAYDt7c7o1YzxOLj42IzcDgRTClZSa4LMD3as2jxE9LW3L+1Tx9WMH70V
jn+d9HyMDpwXemfQnGkaujPI6IRQK57WiLLfl6JVmm7zYHkk8c8iwzFoZpBp+0gL
aX/hmkBFB43wht5yY6NJuNg79WtpXRvN4vJ7VFAFIyw02aIX7v8VjKQyvB4Q773U
kGZBEf3B9pwcJUEMRFcgJEbBvQ4BoPZ/mniwR2MdTJejEU3CagD9l7TCVYc5SPkT
c6h4ZW6KxNzc6exjfvZIoSGmvEi2EkPB0fPkFmgDZBvZDo4ud/ln/JJEfD+lO32C
037mRZ8o97lPvP2hukoJSpApmAGOL2URiYIZyLMp50FzuJPR7MTxhY3JXKXfSpao
JGi7ngm35Wqr06xkewoAGiuTtnWc4dq1IvDE7L2z/BpLu2mBqXocqBjLybK107sZ
72tLOMFV7+c+EhhuFGdpbzEG/iN0Ugh/vENR1Zrp+XUzv91QDlqaPtaZs1j+kSlj
OzJb5FElRAH0ybTu68rHAWgQt9Dd8MqIdI7IchpdnYYL4c4DtQ60unl3S1++u54o
e3eHICfSn+EuU6yPWhtWbQGkch72Hqe8mCPF64MVv47ZphMS7Qe+MlmCpRJ2ZFE7
xTp31VPwQRJIjyYeqRLrn23+j0gfPAlYKxuWNmfV/heTXhW7v6wB9uFveqi+20HC
zsaLjsacvriiOHdfx8IhHCRvQ1emvolx/N7RXxZQGh/L+Bapda/eXICk+8M7fx5C
Yh09+vshoP8nJN4J0jsUe1p8arXZux0WOKiwrTi5NlkoL13PEBTNyuzI70quzx5u
NRLOYelfIqP9kvy2wMMF97w+dqZfE8/tOmdBxxD3LJM9mOjrj1AOxUC8PlavDKDL
hwNIHbswCxdSHaHguqvS1P0RjLwzb/l67H5wJTUqXR1ZXvcThqqKkCnbtPUHBvTc
ZXaBs1tfyk5yz7g2cuMl2xDXHfePXaluAWMP37HOClXR/YXXvI62dd1HUWvRVXNr
Bn53FB9SPp0XR7pHY0lZ2DE0puzLYUWf6b4p0yjI099JJ3QVl58esKyhJPJzNYgz
/dxQQouxhTmF77YaJtyz5nF0A74cvoy2FYQx8raK6YlzkJyMx/93pAk4sVGfuN8e
kXxijQf+aEMUHn6nqwM3SkHmtYZ/gFI9hCzRkyWoHaBNfoaSXjC+HmlPIIhrhbBL
TpmBemNCNY15H6kV0sZYmEgQj6Ee+dmqTnOZLhcBbvIrEN9Daw/rhFd/1Yoa88yl
G3UOaBnG4vq6I5EFNwOU6zT4HEIZxmt/CBx1Zg1+BjmwGhp9W7xEA8X2wqEgeNWw
i9qTvHiCbQiWuY/edU2L3DnO9H7clzz8GLEK5Yspvef6fnNEys/2K+Oe2IXu/dQ5
qgApUFQSrzsw7ex9ns3xc1u6bbtnI3MVvtSRZCEASjPDAKafm4gDJyuS58WkGQfs
QELHo2X/xw4+N1RCvLDqQDOZkqv2XVptbZ8eKVXxpE48ar1WqPcUkOYbH+t4Lobx
ztBwX4KOpoTlLHa7EdQYsT7//rz4PFAwhVGiC3ufUNv/q/cLF2Do0y4w1H0jaPVj
YtQbLHjCjKw+BhDvjpcOy9nkl7UC25d/LVUOLaFkSGBlKW8FHm6nRy6BWPaIcMvW
aR4mJwbgjWhsplfvEpBTaZ+dJ2IikVZ2cF4ARzizBfCKXPMME5iFfFiUL007qsYq
X0ycicDQPfB/unzHQyckE39oMhcUp0nD9OV1QEAf5cZ1bNPgrD3+qoaxmKi3pAd/
iKBCpqQAOeQOtqgvKvzagDZpCqF3PyYc9/QIAtEcAn74+g4Qkezxy+/UQhvDvhEc
g7QscefVOFqtVpisTDZ+OXa3A0eBEmgZw/3lSVgL3rK7iaIzLfJcoyL2B4o8qsGE
NT2DRIBqlVBKzSO8mF2/TB5JMBqsExN3FOt9Z0qymjtyKE9lyK9IQCc2fJwYYIg5
UYfN0JyXfHpxUxSquCQPMXMg4f5sIWpg6WPA78wEna2YVgdujBmwG3yHtF7LIjX6
MiZ/1MqGY8ZkgKbZgUxE2qJ/vYySMGj+pRxuzT8nSaC7qNEDXEZZQL1L26G4Tg7j
/r/gRJK+ofyeFU3PIdg/x/fZQCiH6WUYV/dSBcRVdaU36jU3eSOxZyyIKro+W2y3
5uaFRpQe3wbmWUuLHn4V9zJcxhsGlM6Q9zydI4U5n75/7zuWA6G+5Cnb+H3XIld7
qQqc/1njnl4/DvkrgDKiVRt68UKfDA7Ji15W7U+jo80xq7TnYGIA5PJC75AAoGrr
x9ynfYB7m/hNyIfYm0Rtyl5dSxqWvtdeZB67taGLfK4plp6xwgnXtdneAwevuVeg
o39saglCLvCCZ8eaiwgV1xHS3e4qD71NoJzMDC4iY5+xDPhj7OBw4EhtTLi+X5ea
io4atOLj6uuNRJlE7o+6bzZhMWA2dnWF5N3n3b8mFEg51GbZBglDivyntJWpyuFL
tluYE3cok6Ve2mdungIqwl37l1XgYPdVQgjPEea/aAaGY55f87C/h2wUVT2njmyz
MYSgQqv30ulMpGb+WfdeostJqqpVWT9NgM8Jjxi3e6nFoJR86slFl2+duhimSF74
LyohsuE4qIhZX3eMUok0zOi8kDXbXzcIWWJnasLaAD+ttFcXU6HII3TtgYmMryen
cFGQJ8t95gZyMmcJUa2BkC/u+EOcI+ZgYpK6ojR8KZ4Ij5SOtrOfZuk5cqJ67BnP
GK0SeBVGquLQYLJkF1fmIY+yZnZ7lmD1RW2BYlt+VeZ/q8I1fUR3nyNet7Aka4ct
yms1Hm2P+U3+JNsJHv1Xfww7FWjk7PZ7ak0xdZhxFXLZrrzKNaT6mj6YVhhcaKd8
TMc+cDJXK/r9jgD1goyyoLMuvJ3k5RDPVIBHR0788D3hETwh+fRysX1hqw28ALrQ
3o8jf2aPqqG9e3Bjja3QG79V2kX/Sb68p9RVdmjKfwN2q0/cX6gtodGZETn9AyAL
VhhD3XCzYQln0vEaB4NFG/36+HX99Q49Tr6Z4y5/ZHI909Tl2+0fSChS3y0yQiHq
b3kI9GPESxnNAJXDp7zorhdbiaIrkMnd9UnFSKErgRzOsHjaXdXfGrskgGImR0el
7WnZGEuS6jtjmau/vlWVoZhew21HdGHvfvDhvCbts2tkFwrbROVOkt3SUggZm8Qe
+uMf1B3Ds4MgYlNS+29Ej0hQEbIS0ibkAi1oO3zMd/kMAVrncXZH9a2k2t9j00Gy
lX2XnVztuR9XqONU/yaBZzsniRkg7PFHB16VMq2/TDEZjK2IGgAIJULWKVFmICPR
INwrfybls3Wf9Ic5XMm6m303vBqPMf9/1PxSSXYNMcdEcOEu3fmQnSuadnKxpYmK
pXPi1S2f5qoPqnvmqU0lNV74yJ1ggF4q+Rel1mkA9umSRl6NxM6FnXorUyzDiVKu
+ezgRzJoO3avXzJXowL+9xWqYXQ53dxKwknEX2xxqVR3LGGhcZoilX9oMXkoMFvs
X7zm3jGfJ2MjzQUg4MSBlZLNzUrg+O12CGtMLjyv9zhcje0miu+/+0VzHUCRNNKg
ASpu6gMFTSp88IQ4ElZaIsMNEgfc9HNAW2e8KAWntON4EoHUtq2hqzLGDh4nuy9X
PUrWO2OwwEe3xkXO7Z15bury56KtyBKqKEHe/fw7ExYCEeAlht+u2iX27I8MxFEL
WJjcQYlZZQaa/ZpiRgRVTqoDUG+3G3OVNwxWrMjkq4IpqiGAX/8F5EfGPTVBBFi5
kNSB9qdixVFdbBncirb6BDtyPr72l+JUT5kTiWdt7FAb0Y/IYKcabbDdoU0mZTz4
nWo6ED7seAuYsuJMcHjiQEKvnntO8Rlnr+NSOc8WpgWir9Z43SzLnVbnbSt/JdGY
UOBDWoD0pi7isbs+0ueomxk7nI1ojIW6QyaNQJmt1szYV5Q0jI/z8shWe73Cj9Td
UBHsj7g5NnwPeThRxWzAjGhK7gJW84W9+cpkFHEj4jyNXapkuCDUwUWyuJppUh0I
BZCjOghJAaDyiKHnhF0ICzIx5Z/I15/pbpoKacbIyjcAdcmkREY7FmVXNfrgmsp1
M4rSYiYvwyMcSGDiT+ZcViffBktnwPEYY2fjQ4ISb/CjE3ENhHqE7yrBnpjl038V
wxufc2Grnc7ZXYdNg48vGElvrIJbNC0L8OunrIwdDKbbp+Wszs2rYDDLcAZ5bR85
ncp2SAlhIc9QcyOc8rb1q1Nggt2QrZk/Zj9CsXd1pyH8HT0E4R+wUuxQc5/Zs9nH
j+2ht2NzAkcOCf16CZODjIct08BIEK73n6Jte3XezPIx63FycB4s7MwE2L9jFZ4M
ManwGjjyPdUb0dk8ROHPIQ+EPp/SAn1UkYwi7WqRHzHTVSmbwulwWvM4KX2mtCjO
iULWatGSZqiDgg2DDscvoorkUr6OZ8gCz0i9nCjsN1JFyL/G6oELgj3DikLqy7Sc
IhFw0HaG9HTnPOfB0BwpwuFUCXlQfJxSRZ5K4c1QaP3rEk7/X5J0ajm2akPPyETZ
T63XTLbiW+2Y7Xo9EPq1ltSCckMdosvxGu0dq2enw1cRihe5eR4nO49LdpQTB1QJ
j2qBntBidz5pytHa/LoZx3gKoaZqE8Pm13PRWpLmXGG7VGgOsu1OcS23bYBm1zQB
FtEwFvQuFu0JTocCRoAZ5A2VcSXrTazdEPYMrVfDlRZWS0iHAYI867bda/cjtuTk
HBCvbu7DPwfasmFOv2QtRhQIJZWceGMNURjMZlowHitHzfbmMmWDeYvbrg+7Hx0r
H1IBx4IoT2MxmuYA9JFJ6a8kmLT1rSa+X3aj9GySopMz4/JuuTAUoo6hDVVAHk+n
gErx2yK3GVib77LWzbWDr5rUxwgpcvQ9BpTUH6SQfhr188j0qeCp8HB45f2j+IsK
gomFyPYWXEvmZja+tjY/ykJsCjQeY145gR+9KL7sJzpk3G7ObVJM/Q3+Pzk/rmYZ
Wa1yj445wMHtjUDKd+xUr2zhwLwyb8xAb4E8qCim59LN4ttkdn8iER1ssrhfZVou
WQVbvsxhu7+wN6le8eiq3fKwakZnDGXN/33AQSLs5NaYFzFGK6lTM6SqQ1xzCM6x
SneolPp7dq4U1uBZrY5irQc5KFlIBXc44dd2Hyd4N0k+qogq1OJpUH/595a2ijbE
1UcEoX9QRL7QJyELWlxPVa7yE7Za0CaVFS+2Kh2DCQPO2OwhA6T4Hg40yet2mA75
CcYv+GMF+Le7g8UP5XKKKOlMvBB3H4S6rTiir1/9PhQFUgUn7EbGHEbkqEV09yjX
N2lZIcdcvkrUVGHGNFIfzNsbDuZNG1X4gdixRgwedxQ8/p5SWyYCnkD1363RK63J
RTtnInQDR/f/AbyO0HWsLuevwFIJZIWl3FaGXN7TVvgY0u20dz5EJX7z2eyGHK/b
EW72AIRzmenceedsu1yOOYlJxKnqr3KsdsAT8MBUsDmPqxpXBuF0aTECh+BKmTgX
IE8isUgyPRlVVGBxdU2I3bCDUlROgKrLX4LORr6+a4VXMT4tlAKBHwVUVy3GKtYU
f3KCqkvR+IsKhuci6jhZWH7l0TXA9zjKLZqFOzPJRN4/9Xa5cr9lkDlvEmDDEKIl
UEYnGD9ybp4rcrZxAn6PcAerrpvNzfnlMGX9q38j2SidMLonqMbT3EFPFiErIJ47
dq8cmDLOoW3GmHKsDmxX0FSm3e621XsES8wlQNJOLSxg0vY2OAJPBgftyxL4St4f
/awoyhmh1Kj4kHdpTkdSbG8FgrJWxW/bl4SZ7VKg9qjNY0iGb9lvGAM4QnHjbxPY
bxBGCkVdNqbigBcftEqoGMkk1hiJCFzJbzJkvQ6V1wmj7R27KLk/bZjvd7iMCvb+
y8jFR3h6O97G51Bl2amwNjGI5Wtbk6Qa1QbfejaeJ1BZ3WdCjNtEklsRHtA1bdqp
qxzItKAuLu66gvNBtNBfi0jmeYCPBO8+nvvRJdSHpZ+/jre3j57Sa6MYOURid2KJ
Y5nuRUVONhF/y5liofPd8elVtH4pIgONAb0lKAe8l09VZOsGucEf9lQ/Z1/vN0Q1
5TGdWdPj8Kj36SDznw16alZvbV2sZACxyikPf8TTtBAAhIxopAPoovSLYCwRCXEH
DOokC2PsfaGVthbfrd2SBWQtchm1KRRXV7jtCaMOiM/nZ1xHixoj7hoaR9+02YBC
qPTyq2XsDrXFrZwMMoQ4Yve0FM8EHNvpm+VIlJabnv7PnFPgjgGGKl+7c922QlIu
CwZ0qUs07dD5v0fBBM0qt2nZTYRiGB4JfcJ9QyLdnmgW0lK2+2bWI60lnkzAKCUx
xRPZ0wCxy4sNP+X2bsNqD9VSILMsc2iQsJ0hvO6kYHKbXYFZL4rD+zx2idMA0Li7
6xezcaISL4kWltkN11FzafYCo7GZnq5SObTH+3EEOfig1vgDZVNiSPeZie5Em3uN
0VGll40slEc6nYeYpnnmqA==
`protect END_PROTECTED
