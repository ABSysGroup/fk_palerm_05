`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KCB9YgekXPdc+PKB8U0XXQOa7C78DFHOqQwXhsixBYsYcrt1vhK7rb2s5YHI2jOn
LEnZMBV1nENSpLYECp82ws4sis0eV0ZFSuoRmSgPQbqOqKtIVi9taxl9NHluNaGO
Fhbo3SBqx+M3NS0jTEyOIKAkfdChNxW1FBPCohxfZhJ6KFZBOCM49viiMeL6mfi1
HPWJFxy4x8S68XrCUeK8qxLndV28XDW3BzLzTbd4IqBCNtMSl8GLkKPV4Lu0YS6P
ausYF1V9Mw8O/ZRVE1cBWR6AZcmGw5KqZl8lgpLBH17cmfuzD7L8DZAaO58OrTfT
MOojRKSReVTRJxmorUoTI8KqiF/8NXzZR4Sv9Qz6YFI/lwC/EPRzSHPV0J8ooy1c
Fl9tqQiSfAjvqb7HMFJjt6lhEi8QMRaOop8YGERViLs=
`protect END_PROTECTED
