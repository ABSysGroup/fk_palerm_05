`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZHmgDFo/RWC9QwYaMDkOibB2faCxA9Er+WfWy1ZvyksTom09zd1D3qRQlROkGaAj
Zh2ZKYyyt7nzxjPeRGt/WRyElsbwKrmCrBxbkOwON6s5Lxdq8BIvnGwv4QaURHIb
FJq4iJU5kX3QrFkaKtWiex8FiKuA2sQGuGUIaDW2LbXGn5OPnl3mbZdBRhNebgx9
FnHqkhLg6Iw73IoCpOpcyocOOYyvNyXz2czOR7QG6P8sVRWdGeMxburAOtb+JgT2
BZ/hPDpDFN0mfS2sGsOOOg==
`protect END_PROTECTED
