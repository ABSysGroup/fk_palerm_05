`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oePKTjOrJF2AyELCrWnh2L9nMShE+7/T8/6KN3NxUrG2ektGdB0i9SljT7HJokUf
ZktCN97emGTOLjSEoxHvb4sn4rcZlhqZoQXjIKYa1NofAqJzjeh6LHO3beiaYgeo
wvWlvOJmBqkkvuQcrsDuRo3OwoaamIdyYq8qvN47uScs1cpycKopet37kUM7CnZd
/eGXiNB7CWQYYPcIT5vcd+lWxmjbv4sj5kU2WGOpFB/bb79kap6UYkXM2tXbaYzM
CNLr9icb0yCUvA+tOVS4MYxo9ewqZLR9p6x3vGS2uemp/PfVd1JW1HjySdY2FQyC
46NVNKliSC6hvGVGtz5jYR0QgQlwhGvDPc8tbXpiH0Zm0Va+y8uitt5LEbieIQKo
cvQU3LWciX8/g7xXmkO6xptvpwK4aUifyt5TT8Bo/gFoyqhz+I27FS0U/je80fXb
gm6AUlauKxdoFX50tRsuvdj/JTNSe+AZTyFAk3VU9DuANiDVKS0F15lYCZkuHeaz
jy6GVJxLAlMxPhp4xq1CdbBIw1gwvvo7tuwRRg10lyo6mCc9l0HCE/z2YEcDNpbk
HZ6hxCZyg3SbFwmwkRa+IG5/tCXQUr5N/zJTSHfOcQQkIyRfD1vH536meOUy6B/c
UWLSMaBpPY1h7+49KjjENQeFPg3wKDHZHAl7wiHyB8oJrYGeLRebsg67x5+vE2lp
rAEU2nKSwC6NPoY8ZtqjJIRlNgruCu2DKYzApwQkbOEcQXGuoif4DVhdsWge6crC
tl/YASeICuPRTHM2fal2oeMfI5JL399VZdUMpsJvz4kfsPPUqVSdBVK3iTmKT5Lb
8/cPbCquR9Ic4r2Dofzb5ae3PqfJ7dH22JZGhK0f5udbU01zzhHIJEXh1I2UxSV4
/fcArq5rGwsBPGYlo9RP64nX/xfBvk5vD5svIi4bprFL+6lCVA8LzBJWE10CtblE
PMEURRZjp6BcIWbuBH6yERYqv5U1WZ6MEn03akxSweOj0xK4JzzzCeU8Wizj4uiu
VU0h+eUJ+hsvy34j/tdwSk0EOF5ZpqSyV65K+nvFUvdcZ8JvaQ34h6A+nw6bzDBv
PtEAzJkhq9y/lu9rFGLLPoKp8zueCbYs5SXEvi0nBumyjZ2DD9mIuDczSObkPXEg
IbwLBGHBA7WQv1dyFbZf/DQlwk3+0AjMb7PXqnUFZyYpfTZjvkFD8XUJxWFftCHG
VBQ4VTwVApacR/rgMZiw9ntc5zTQOfMnAYVQeHAIPd0gFODXL2Oq/fJ35Q0hcc04
1ppm4KiTnk9BCABthAPSLyU4zf+e4mWxIpHqRlBwekOaVGRP1DUMp7Hctpg2Cn0Z
EVF0mF6oioVLGvYKaG1qWDAw2ZhOC6fTrAGS8f9HJ/9VHPWnv30DFknw9CRUxwpk
wYDGAUR9btrFvINlcLchZ0i1jb6kfwUIf3lT33Ze3/R1qPkA3xYIKNBB3hSYOC/r
7U2F5P3BSAC45jzUzxUwFzWeKY9Hkzh/uJrjbOnA/jkM2HoFR7wgHHoPegmbr9ki
vouuRKkWEQ3ZBTnBYDsA/NNGfGycJTnnwbVKVqMK4qfuKZAS2J8FSg1lH2a2I3zJ
MO0dOAdHlmnjQpB7xqVttuLWJaN/rZnBEX9ClgarJEa+PDLp5U7CiyfiPqazdDY8
lHd282EU1kUdfBSQWnssd23xP1A1hUKnkxVQeCdyMDGI8rXSFAM3WvHifYABei7N
N3fdPiVbjD9xHZhiHUj6Tn55C05KpE11RGs9QFDbAsREbjuawxe5ooWvrjkctnol
F52hD0mIpUzC55iejk0Q/5kLUe0Ea93Oqg8Joc1HMM298C409+qiCKWOxSK4RaOk
wSIW8yM8Jpo+nfX6oqvEi2Nqt9J/NSsTRRyOTRoD5pagYC7RpHgYlZfdoTsd2Yi6
K7flG1AKrZVnOnmjTu1Gesx8tKrB0isKZs2BTo2Pr8uCuLzCxR3O9xnG8FRRhQuR
ijfi/Lh8hbXApaDLE0oi9yy/e7j9CEoyL0D2zg2a0V4TRRi7QPOMQpNJVBJqWQTz
izzdK5RDup9gKcXu8dEGvpUjMMd4lgE32wKCDLK9ls3ndc/OxwpgtvpgpR2bvNBe
2E5oKB0BhExBwKG+UW3iP8Yt6E6HYY/WxgT386j1Oi8hUpJc8JJVMN06bCQGLV4t
YBa1AgtSsDX/iMWiADS5GvidBCtDTMG0JzUuLt+/1dwBeFXW38WiDZWNZEFHU0yq
lV4xDbYjut4W8YKzy9thyltilgLXQp3uPuBoF8dReSHnHjvYinN+W2SE4+465kiH
rrTRQljgEJ4W54OiXRbxkDKv1ekPaObertxWhFz+jeaqonknL5iHzfUONt3Qsp4u
b9nK4Y33wNVOD7UObhP5UyAAydnjtTbcxWck9IY/gftRbKZWmMfjaL5ouT43gX6F
mZwRntvtHr5VO/n3dYAQJIB8yFNWemoY0Tl7CHd3H72BQr2vsGUBNBpUYRIb9IXj
AuKOa43mP75MywFIwkWgy4csxo5jugW1hK8it68oq3PX2OgBfBOKZh6Wf6nyZVPc
sERBPurweD1OwH7C9jjbFz3vG0kAxN67orbhGlpDhsIPjAAtzKJVNQYrMeFkaIiP
AIVnB4mARX1XbO8V155ipW/T0QPmgUeryiVT0HQqEfohMJPSfhzS9EuIXjjJXiEu
oGK6WXkbDVW1Cuj8ESLxxyHDdKvM3Uh1ygnNGmJZ4PaZdesI7BGwc0sa4QhhX98k
K6s+ZsPD7BHm5gjoStlcyAwM8fqlWusQs09RHQlafn5JVAS13f4kvaY/wq5aBCug
uPdP4k8JSM5Lqbz/JjFpxUVup4IT6knDFs6F/zkAUDWKAxHHpAlPx9JK2jfrdEui
s/LvfA5C1VEqpLSl++yF8I/AoL35sdiYa5e/9RfU5DamAk0IVv0KUx4abYwcof+x
jfGKCG873H33gBU+NhKANPAszrlWSrbmVR+bi5J3URBr9sbgZcYa41tps4yUnQNn
XqvV10/+IbP7lLriIITQPQjwxGSEDR+oD7r28TErxXyxorIY+PXIG/lerEGJoK88
SRYj87xXXCrASn9dafP3Pq8rUru3Zokfg3MpEcmVJCERUbj6zuszpUZf6NkX3Z67
N13a+4AZcFHNu6geSAsoUCV9EFPjUwCH+XH5LYzl+HwHEai19KYWoJNG3j4jkKHJ
LdOC+Nv99Zht2nWbIL9hWoQa/NLktmgNxMll9b3V+rbIap1KPF6dKJYqeEW9l/Y9
UNuQ1in4Dg/LLcwk8cWkTDYhzW/bVh886En7DT5yjFoT70JXt64pcR8y7JzUv+dX
6paxcf7zPrq8FaUfH5JxCLj3yuXW0a+eNda75zdQoKrjdcutSl8AlqiiYy8bxGC1
jJ9rhEk8/lE9cebLhejRfyxvGc3COBItn2mTX6CIE2xO7IQSxyQ+XuTytWTCucND
KVhrBNASTJg7jn75IZ4GhUosP2CdyZdfiD3GdC3BJ7uh6R19vn5GT0R0dYhTLO6u
KbPfRfyZ0SA2+wCm00YdkJTWsxSol1dTBdRho01jhmOi4DWhY/3NhTJlTiOQZQi1
MuPRszyHShl1D/9UjSZAQtMD+jxXaZAR7vWBFRcZrn5UDp7o2caD1N1oEJkD9KQG
0nbDOPljqb2fzK327Bvcgz+3Mm/zndlTegOfabRLA3eOCTDEYN+ubTkMkGhDC6MW
+qF26ScCqHWV9us4kmRnwEuuxFW7RG8FtEa3CzGoaHAChMDHULHGDrtq5MmWVUHR
vaJjs0e1yaNZg8kv/mq2mzPvNeEFlnhVuavc91pbY8UFraEsxLaAZ4mLdXtwFWjS
x47jaMfpwG/v6cTOOM3Ew1vApLrupHjgEhfnF704tG00B87YJRENzP11Ww2DJsFn
vIKOCVpLKXhFgMlvXAE7FO/nDwm26FTBwaBLEimL3X5EfO8t59xrUUVmGUqbe8mE
n/aXyQOqnFuHZ7bhFzdxTREJtxRI6iQ8Gbsm9DG0fP20uDTi+c4mvAagRvPqS58Y
ytQbUvCm1f/cZ/6rmYDuI0RzSYFVIxkcA+1rNaJ0KsC7P7yV633iwAvp7L65s/4e
CxOOZyvwINDUJQ33VmcqxU72XvdQp3VC8uuNRGLBF4qGUegoOeko+O9RdxAxsqNE
5eYrKaATS025D7YTSdZSt+2zXVA4qKIXdrst24yBiCipqG7UpbAQlbJiSj38UxKQ
wpg5xv8LTxGIanu7fNMlH49Ag/XxYQndXmy6PWMPl0aU09X5uAcMEeiznHc1xhOw
8RzH8TJUrGVwdBuxj8q0ok4//rSmIJygDwPpx3H5ntChTcePF2wfMR5FvCMNT2Zu
h/z9KdddX5WGB7vhGlX/IJ/+rW/H19L/0FB8zXI9gJpKtWPr/W6JWx93sM5hkBQd
X83aLdwzoHnRApMnMvlMIF9mTY2QumCzysnIthFSmDWNzeOVVACDKfF/HPYx3n3e
OLsOeqYEysK+i6ijr5nG6jxhNm0EenQOb4Pip7GDCN+dZTaYMXzP439SmkokIEkv
8qD/DvRVzd+lN/QmKIVk4znWfLQhzFpj6RweEpA9S3jKwAo+5NNar56wJyp3R924
IC11hcrHnMyQale2uZ/KJD6/NTWe3ASUhIFe3ttYLbrBN5diwqNvbwIfGpWv3+Y6
puygh1CMGxkCuKP6Nwb7QQ==
`protect END_PROTECTED
