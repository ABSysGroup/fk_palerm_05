`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8TrvLHYSZ3dvjYPX/7LrM07f2uOWSbOSk0e1JWcnFFxFHz9Lf4M6k7lsD8HHFXKH
6SHQyJ7pGB5CeKc4+sElt58lGs40eJMWvuQC9/CEyU9ulsFWQNvhxECTVZEjFXLC
f48hZoldyg4VjJrMoIUg1kH5y4PcQK/F8KuXqObfPH4EERTI7lwcHXlC/ins1n5g
XRXHyxYvs1KhIiniwBsCnMK8yTYqjGrNdq13sbYYugZ7CZf0VBLhB20DDq8+CrZY
elvxM7HqwVgu1h38fYC1RhqLfY/O8F/DxkLPmFRm/e2y+hA6CmAgTxP4hNwSfdFs
oso3/HPw9BXzfcVk2Sey7ingEdVtV0JC9enq0jRpW9UxsKcH7Hc+hHW+HzxRGn9b
sQEw0LgYKmKmxUf5qrNEFKUGNTkGA6SlO0UUSdeWeIY2D5evA3T2OuuQ9wubcdy9
`protect END_PROTECTED
