`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g6Q6qL+RZkn6cHRFpxF1yv8QmIompqmWAriGEDjiQ4BcCE/kjyMzK4bt4Cna/exG
d3iEolSpYgfrbTW7X6prhm++8dZzffOqdTrqXFdiEFJzj2cvwpdUzSGAAp8PGpTh
Ja5vy4MKcjMDzHkQGBy2tTk++ryCbcYoNRza4wMzEKzudwe+unylAnjFk+vOwyBk
pEdu3cZDyE5gWI0AMEwmH6xL83mqGyQa2yWA4UCGTk6e5ybXa4vME1W6NCtzNfeU
gX5vzLaqE/JHEd7XoIHZ1uODIukL+AaefhWwxGt2Mm6z0tIOt2O3QsNtrIlOpgZD
Vxgb+syK07nOdeLoxaPXcxaeac0uVGVk0T/6pts35vpN2J9YE14AzKWm2W8ZcGgS
0NFdjRcmsdBvNuePJwdPaOu+rvITB75D32IxlglSEgMbTvf2wuIE2qc7in5i7yoZ
eHTSLjT3g5yaOHAPgdzOgnQRCcsNZCZlxyv3of9WuCKWJ5stNwORtV2L2acpE6cy
+s+vhL/84CZZnErEMD05onXJu0pLcngpDYFvRT9IY6EjboHK9rzRYb2Oqv8UPaDr
ODH8epimBOXqm9L4MKkyOCOmcOVRrT4sZAhIU31KiZFe4ioH7sTz7Med7StGzMMx
ZlJplAyo7Dzm9I7V/RvbzibZIxO5Jvd6BV4uKWDCMVpookOBGJxmT7AWlZS1AxDa
GmEV684Xs+mUyQ4HM3UF9d5VRsYxMyf4SiJi7wRzPb4TA6Gi0Gi3HdseLhETOre0
ku9BfXwFC8t3Ci12mtg0aed9d77eO9Pq4yxVR/lMyqoGGoEpiS5lCYpAZSd+7jW4
NzkQSNwGa8WaN3YduL44ZtbC83RpMef5NtZYxW+45va/zr/o2uKuUtXDoN19P8TM
cJk3ZENI3cV/Kgn8PVWC3YhiCEzJkfi8Q89GGKS52xqb2gOxL/PFy5T9RzZ2tvFM
sJeutcd47/1fopWSpDutijK1Qov47lzQpM57ZYABbs9sQzfvL8bWPvTWpRApVoTr
vZJOR+dPBfuO/Pu12HSMr/zIq8ez3u2BG6ytdhnxx5L3q5Nih/cp0wLgIz/kfI5G
8l6M39mu+ZWTOKICeOE2bAk94DCYF1Gyd3pPN6BU7qISUcdIiyQEs/kmOWqH2if4
TyQEjaNvSOfBh659BNCA/3c1XcXg9vYmFD6q26SQVYPvc0s7edBlo8MnChQZAQ11
qtdb7w34sNMI6BMvAX1EAXSxH+KW+YRl/PvwFhrfqlverHeo0Dw8uRiw4jojec3Q
npS0FcYsxN62KOMeKbcyjX+GtfKGGszkg2FY3U76i4tSyWWoNJxrpn7EAcJH0jhC
TOX0aBKQpiuHf96l5ZqsFfdbwDMQ2PCcvyf0CugjJ58ZiN7iwYsNUJAPZpidy/hw
/mtnSh255FUMPaeUYTJS89xG3o6HRIhy3az9uGzJz8iRZNTrHyUZZq6fX/PZCfWI
czhGzaATpfJku4fw5IRsD+2aEGr0dSlUa3nCStElWtaBdqsijOuBTQggUmOhDuav
Uq/+3KVYnjism3i1i79MYqzw+2f5XqcDaSwuX5eLIZk8olYBBOkTqA3OO2EMBUZL
KUbA3RYlaS2t2wDp98baq5XQ5bw80+yIP2RHRGIBGu1IMji478/lchEwVAVUgxI0
7ujMnpRTpy02GPSqHMQ6wN265zFA0kxPK/56bEkBziJxpdr3EFi5BplQfzjqUX9L
IAaqrUJIwS1GR4sKDzKSKKuyki/M+1+Z1LXSeVrXAuFxQG0YbcUHsaBFMZonXa/y
3uknBHSgkDXapdZ7Tjfe/NCKMB2JWuTCoJPC61sJjJe1LRsPduo9I3IJmfoHV37K
RR4vqiZneSW2FOf4Y7cEPnFxiFXB7ljQ9oGj/M3At7xKyuH8hxzkhikM9fY0Cw6u
CvpY//L0eLKfIZAfznI1kP30KpBJyg0v36TVzO7kiwyCKFYU57kj11BeFWBOGvRF
sCBwTuuRG4b5G9KgcHiJN+E22uoWFftRQ+tyXN2o9OGbGD8saqY5CSxCwnS7IhQW
hdnKi4QDVPws5WhlUqJhmaVTdTZreg/wuuy+IT5TGJg=
`protect END_PROTECTED
