`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lKVvoVOpwu5DgK61vm3oyLxNuMcQpJ4oH9ZyKCZmb1n1IGlOsH4r1fLQ2fERswvw
Dy5vt9iH/Ru7TZz7ov9BAgvfEGPAb8XVUrZlwLIC2KP25t4R30c43g6vYYIcRAdq
Z9nMOJxeQYlNbF6W+Q2UE5B7hUrmefuyD645q5YphyPd3pt+IpWpImi9U00QdVPa
OU09Npdng8wR4BirNbOI6zExqYcR4wLxbbo3h8i+jPKFRtOhou7aUbKfE0dFDCmM
+bSpLX8KE8wNlgCBfupbs5CqLoyZbhkdm8EXiaepDZU=
`protect END_PROTECTED
