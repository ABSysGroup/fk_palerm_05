`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lexFfYEnvwPa0QusaJyQH3wcxkR0vw/W76UdGl0ArVzamyAvVVmr4PPjFA7YyCdk
FHqTBqZGj2d3VtGGXbxqRtnUUJDwVjnCpCOcyGDsuhE5vnoIHofO7YcJtAl4J6lC
/lvhNtsWaPUcINIk3gvE+sICUcHzzhDdevx2Fz9sZ8GizXu7aeHFBL5GlBcViQ6d
BxhKhy3N/kg/U67GE/elPHsSj2Hw0xrSs7fowbvnc4C84P/YZDgN2YVbqk2OhLvY
xGOs0cWXyhwCcBEQdWtPC0zpS+nmD79FuVDHY/2eayvd5zIYR+53PDxsDi+N/Zig
8KFwFaSpagyUSQuuTxtcLOc7MTKPLDoMCpzbpJJlm9POgLbjWJ8d7wlAxc6Quz81
dXA2e57DPF4bCnDRAjus/lD1TWAfaidsHxCf4Bj9pWTWWGY/wDuOKDCMV6Y8ZJUW
WYbe++nDOR+IEjaRT+6ukU/PJRT97DcUpQ/r97tL6fSOSCw/mpgsa4yU2gRiurRw
JQFlKl2ZKEFFanWLz7Yjjx2MKX6NSHwNuNAoo6sN85hO5kENhBjDRqnr1yP5wriW
x1bOvNy6z5Rbc39pvDdKlw==
`protect END_PROTECTED
