`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+yYVgdE7Hp1fmwC8tOtgLSgocVfwNVfLURwSU62zjjNWyZvP4Tf8lKjTFBkodDy7
WXEXYWlYIUmKkLCInYx5pXqmBtyspRjSdEicF170phSJYLEK1tVIa8K24JqHH4Cr
YIPMM8xj2eTMpXoqHCRZnTwHamau9/A84UZBykz6EVAFx1wxeRcI1FZCWbHiv5un
QUcDRnxfSMVKwBi9xe+rZBMzDFvuGn0WTW9fu/dU9OdysiRTIRf8pKeXuB+NsCIT
nnG7MOMQXDIWp+D37K2j8IbUlJAYmYm2n/caCSty740iXws9pvPYVtqLisGdZpUu
eD8xiaTf+OrGKLGHl6MvTQ==
`protect END_PROTECTED
