`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DvcJ2jEd/579B+0CinFPVD3QPqPr1baZ1GH0GhGS478Ipc32nAlIdI62t/3DAD0N
tyti4ZVZK0ogEkhi3o7ZPCx2NI/OgErn/HnKg8E2njIyKeBd3hWh9k/H3Oq2mDvd
V2llVjo/zRyEPmboK1igMnvSLpHjUd+KSelXZ7ZnQ4fQeCmNXxhfmkUpVcItCVkZ
ctrNPzRHg2IBPAntfGsRCxtbRETAUmVNdHjOE9/d4ngMLyga6kK+lEiBwFv4+5J3
LMGjTsfq6UOP1qGAnE35x8RI0TyM8vJ1Jb7LsjtT9zUjnro+euSoVPPLQMz3kzjh
Jo0z1+p2xoaRX6BGSD0ha7XGyBnknb1vlSh/xWKTf9EdXFmLomB4dfJePgYeuzwp
lR613UvoYSjy96xqxySbtEicsM5nGRn1RzbYwOR+d4Hecz3ziqbATACSt5Bz3H7C
fYvXXGeA8dyCQ+QDboSHUr4LZ2PF8Hr5lLxPowstUFsmbeunexTn1WJe5/3yq2HM
y/GumF+E/uScyrsXeJ0auf/lN/veMNDZh+zJ/ap8xTSowSI+N6LH/Torln4c4hOh
irP3j6dV8RN5GurF/Eh+NARJ4ZD+rSS0GD8SfHzb7K8B7SEWM7uo845WrY8tS6XM
mtIdd9SNzpzGPjtd4V/q/bLaywiRGm29jncMmV5iDQwgPaDEGXOLMut1aD8ox3oA
Anw2CkWzikH3DoOqq+vIs/Cxi3xaSs4kUO0CyX8VzZhn4MmOYVoMHi3EXI2yhvom
LLCiGLkjpt5kwqqQdB3GMphgSv7BkPcXj7HFrf1/8qOyHZviBsrbDrBC1308ddUj
Btjb9DtKD58Cjdjp8lAY5Fg4FsgN49e8123Cn5i9WRxC7btMVAMEQGbABjyeguLk
byRc69yWmXio7zj4irB183Ny3qGiQZB6Q0pYSn8QY9Xl3ss5QoyL+tXuReszRqhe
iHUyNZ2VD3YAPmzFbTYVZJiXGXULQ6PoQpUAiVdT+5lYBy8z2Sff3HWwoe8c9p8s
1eysFJdFeohghjOis15UGTjBX/gQbgAhWD6LxWfqSFCcyGc16TOzT32suhRQubmW
ysyh4P38C6uxPMxVAymIX38U+H+AMAMOuziESGnKTCMQUR+lANgJBnrt9AIVzikP
2P9DV1GEunOxTt09v48O4lSojIYM3tAK7MsvJEiAGoYkKSz/XWcRT92nAJxG6/go
dqZ8ZaaUKMs8IMu6//SxKMJVKoYA2oBigSLRvS4irySlpPaimn2Paa7nAf9G6MOx
yFBlw9EpwUB1iJ9pV7bxhcY3f5CqMcds44nXZZnPW4SUF70v81zm3fdq7atcl9U1
VeIWuPHiJvtH2issozt8zHD00pKfbHLSEOiTUnWmW+BTYilRXKfadNf2swpjOxG+
lJC6w1h3o1ses/zzRxYPJK5KCnDrEHMmqVK8cKZk37lerFy4CedoC4Zij2MkdLLx
JggVQtVgH+e0MYWMRGahafTIwJ667V7Ud+VfqJadDxr7nJz7N0DHFw0Ogx/VxScm
a8eRmdvlrsegtgGeNbnHZJqmQnPW7Weo9fCcxcnp/pzD7B7kJiVBeVmQsU6xzvZ5
0taStuTisNrNGwIZkbRywEpdHUiNZrx8VW83Au27dmo8D8CADUak9K5Cjv3ZmhjK
3J/4X9zclPS4aULaRptNZCKdVABDxOmQ+ILdO1Vg/nmlJXseoBTF8J0JYhK8qeuD
eUdSJ/4WAnvIba2rGtIjWDABrJKfXi0Y1vfkWChJ23/PNX8fCGFxcTXJmJsF2brB
QxHDMFxqan6ZYJ69YLHvEwKAVbZPH31RwgnSDlccpI5Vv3H2CC8AoZrBpcZz29kA
7VClZe+tV/D69Utv4Dxsvq7kqB9FL/X+fV537Spt/vyTzrCEIgooVwGsibxvRHsS
U4/8yURSeWeBJeyvarsqlmiHsWT7mMrpURsy8CjgWu/dkfa3nANTmJwTicfyNcVE
wh4oVIZcmQs1iHV9fH7R1cLp62aDr9KPZzbXUi/DnB6TihyI+AvyP2GBsmWhhq1O
UHL1bCDXx+Pp3tHjmbYqzN1Xh9JA59rVrlgUgru1i2GT+ZWiiRkR/wKFiu9q1ZcM
2TXvxTXa0SGlRbemGxhCyZ/otVF0SD9BN8cAbqH6qlTX2m4wm5rmx4StNmQiH7E4
tfK5+kdvYEz55qPzQfPSyfJpfwuylMwyV3JZmcmmRLEdV0nPtGmBVENS6+qBZBuo
CkDX+M4o+3+aTmSeQLlpAlqeYb1J930EvWEAZJcSRz+tQLhc586ukM9W7prfzD/d
jpRwQ0GDu3uiIvRG4/WCPwOIGzu7c//hieB8wz7TSHw=
`protect END_PROTECTED
