`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NRgd6xELcd7z9ktXlpiOgFfczxs3UtSGWxfmPH43MB/f3DdB9WqgPL3vPm2gSXvf
0Kmdynx+qMEZr7LN7OkQCn4upgk/5EXjfz410WvJOZkBIWey3Snj0qF28YGhlkLr
covq5BaXhiX2a+/vmFvRHH99eC3KaUk5mv4WSxnd7Y2b2NycKeSjOIMbmwvjCj1R
wQzRotDvm0gdWQp2ArYews6Aup128xNKVSW9ErV+nX2VfqliW+tRkHz9nBmzWciR
pQnQe7FV44Vh1rvfbW4CYWaPGyUtI/tEFsxMH57b+QP6O+dcn4KY26ij4OmTnt9j
6TJQ/S2s5TFpl8wGNB+FxRuBkgiwp+Te6mVS+lB567YsNkKJIkohT0KR+DNaRkXt
purna1L2u8WJa7yAGfZuKXVZu7cZCZNqEjYvVRzGQsXR1KqWxz3im7aLsWcvCrZQ
UKNDPFfrGyvgJN82ZWiNb8nsikKpux1jB59WJTJB8i6MmJsr4SdlzhyQYaLSiYmt
MeJguKd3b12uMpO1IsOV+MesI8A76Vr80Y6V5kaIMw8fY2HbC4Uni9c7eLdITeL3
SR3oydD/It+Nu4BTGbNe6A==
`protect END_PROTECTED
