`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mYiDE+Qhzb/IkesvbpcRyVg4n4pVXmwIFVN/Eqh8wNIH9WzRhmQlVsAvTrf1Bnj9
EcomBrXSj0npS79opIz9RRbD+XUg9Enhs0Rx0VXz/iFoOT2YMLOJeQygZSpiTVBn
aydf0iLY71xQNNLyYM1w1swIND9iH41Y7TOol7JMLRInxQUou1nDVfE7xBKFUmRK
gZ9Oe09PglwOQGP8hpaJGjAs3IBD94ZcqpJEIJhSXOpB+xjkJaV4uIDlbhgk/8Q1
J58TAilQXyelAiqZbsq4jT4dbYuQmzig+2EkD+pRCbCCIQKWLSipszwwkqxuvhAs
Y6aADO6gLcpr8NSZJmcllEjqnVOzniM225ytIohINllSyhXoeDsJRSjjHKN84qhB
QlxnVqVMgRN2FyVXOOIPz62dnwuP2yF6BjI28mTopyk=
`protect END_PROTECTED
