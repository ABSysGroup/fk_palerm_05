`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zDOH8H2uqwiScffMazI1uQvSOvxTl4vFdiXq3qZkHcmQgxNE8jY+GBCl07c8Ta1Z
fOONxSAMGqIBeRdXG3TJPdpamGUWNZrk0UgUeLuW72eYPa3gTUel3S7mCxUshrEv
I6U1+/+ZaIG/o2D7sLn8C6CdCNHRZU5aoqE6IispwRPvidFE4Whfdm6nNh1zZgUE
QBP+lonkpPbwQjtTGtHbGuvREQqneX1qCL3QYd5pkff+df49UMiegqXeFgQCmcWx
Ot3RpqC3WcVWF9JHz6Jf9OghOsll5hDceuIE2Z3OFzgK3L2etuzhLsfO4O49emnw
HWZNW3ad5AJ4/zjYfD62Nu6VEkVtJ/nrq7XcPFCHdrwMucaWLZ9cFyP+zQd8cZZT
5vHHQtzrbJLbMer+Cjey6hfM/2NlBRBdS8v6z1AOvqx0du2U14PMhCahMhzMBK8o
lHS8TLIXyJRzDILn5xW9EWF0txIe5DSi/FFEhKNv3bdX2qHjwHSPuPp2Q4L3l69r
9N6rjXWCtu7i8hkS+nXwwyR5skki0MgOHkm6dFTlfHwBghaV6ahzi6LWo4I87Ypk
zP3Q+NduElypqUbogfdEr82zifIUFQAUGY669GCtfsyVicrsWiyWVMyXIlP88tRh
HUiBwcfbsxjTxrlphY0swzvuU1VlGLwaEVnuKeumxS1pFQhhu6qz42qjqBNmpJZs
`protect END_PROTECTED
