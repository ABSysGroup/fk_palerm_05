`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AAOrcWry6SqbkhlHdkp3nP1MnhnsxBPVcQTBHZfxoBwSogHr2VBJohhiedr7FULK
q2mBkRsSlwsSzGRPUIeD4tiez3yc+rYQI1Bh++K9Ej4ee+nmnbjsMkhiJHGxuvIl
Ch187Sswh20KOiQjD24DYWnIXfKDn9WMXjnXziL7YuXkW22ScosnE46t8ZWS6rKp
sFaJEg8NOVgk9G8gjwCH43r5Jp8B+fQvgo0HsDblP/mEfYpYDORuub0jwwJ4vtJ3
GPjt18NzlGwo1SFviVmKaA==
`protect END_PROTECTED
