`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BvFCOOmS9lgLZsgD5K4JgBvo1jGhP0HaAzelpRctx9cnSWTxzR+fz2Tgutl24s27
lLZ6mtSRp1kKfgEmT2qesSvnhloNMJf7N5h3StegehmokIpqWkm+iisTeP3H68LG
+en8wWV4SefTKilBuhwvKTsrFlGbKn35NKTo9lkbQZYEp3O5VCqCSPy1vhz/U0ka
/sXH/UIkdy76zip4v9ASmXNnOrhY5Qr18CNLDYpIpAkyxJB7p2TvH18zbSeNNSVr
Bug0RI+y4+374Uf/cRO6A+UGgsW2i0U0cxd0DOlQ1CEDyyk9fjQf4WvswyxnQAth
jTBBW0YMuHB8Ovf8URSMJyDlzBie9/hSQKXk2PpXYYVmxDZvp9cRwf8ZgMn29okD
YT3yvmqe9prF7qTmvYtWa6TtALmNs45EB15mp9uTZp0=
`protect END_PROTECTED
