`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
knmIjSFBEMjR35CPmoTKWcHDTKJbzj1YlARD/nwEgL+1aOq/MBYarnF0PHnK81DW
i7lK+DRt0GwUqMhMdFBr+EuBa7LHIL0gido9Ihck1WjpSpUy8V6nQF94AMrgip0+
bpdnjt0h8xZKzdAttM4zWDYYRheEmLKd9xqRrOegD89pLyLfoAIC6S0WHhmubgYp
O2b3l8gwcLwMjyvTeRn5icZHLagRapAPFtz0kXviPoG26rWP4hvIu0KivBMTBL83
WmX3qOLs/h5BosS4G1XlroOdwkfnonL0yBInhqFxUnnl8xigSnIllE+dhlFtBeSc
F9En83l9UV8D+PSYAHOfG2V0nmQF9tWT2/Nz9oYeWuDkZu41GSPyXmsBVZQ19AbT
+Us6zr45f/wfwpbVNh8k5Nq/npB9MOKYWNpcqgbMM0eTzWDRbK5veUviolE1n0uM
FRJuC/bOc+Df39a5oDe3ktzCwacyIwzztm9Ditk6gPE=
`protect END_PROTECTED
