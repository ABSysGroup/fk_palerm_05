`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EQMCstYtaRGgwDR50NZy55Qm/kBohvC5jJzcaZrJ/eGYZHLo75o7j8OcAGNfVUTK
vJsK9Ca2o2ojhIPFlrEljy6RIext0AJ7AhEeCCqjaCBWOP8ECkL8moMRPv5E74IB
hfyGCzFOFNOVNGOFIvBi98GnYAGj8mwJvsdUxkE36aP9d1n+0jD5SWS0RwwN67q4
2M6JVQzxCFQNI7L9zfSM9lsVfygjFDm5Rvphf4ydLTXsy+1DTpbBiYeWsy4rR0VM
2ZZek8SMF6sAw6IRMrAYg5DGz3UyfEEpxQ9C/3Al5O73ggPilgtPflEjNXF1dE8r
j0l8JCHYrrKFImXM7n1/YKiSgeVTu1yHwP5w6tvOpuU6wOHgQuRre533U4uNrlXT
O5PhSA7kZ/Sz/QgEJV+r8NYht1g/A3f0kcxeKkq1O3GFeDPqYZ5QyrjR5nliWtEl
qn0edkzJrcHReTaEIGKEXSYBoiG36z+5Vnbx/QgRI1hhOSQ91l7qtX/593pGqSQg
WLa4d4spqN5ESkixXobGo65hqee4HpWbFNGy2mATp6r/4ot6IMiiwSQ3fXTAOkTI
DSpjSYL/NaRlj9DElTxHGl6vsr+UZKEargmJGxyoCMwAm0Bgq7hvgmuClWf+G/E+
2AaP9n4FdFikTOh7vB7uK9tRxPLWzfDR6wwhcCCF0uVnLIOh9NsXRSr28naR14vt
`protect END_PROTECTED
