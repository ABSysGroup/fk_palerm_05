`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W7+lmxCUQAnb7TCUxblqvyBafkQw1eP0y0KnYPB19+Gtshj/AaTM0rlWcXU06IaY
Jx21M/TBJhZ8lW2zvm3+B3uac9AxDqgR8xSHkTnaAnEPCGpTws4Srp7m6GCQ76Pr
jS2YXVNfjKMvXhzomJW2Gw3J0apY6KIGIGpUqKDvP7HNjRuDGxCbtHBKyfCsxMFt
vOHAMoIvF9JO77lqvu/xI0qpuWAQ2a97/aKa7A9dSD5tIDCV5yht/GroNvxZMikU
0wXlmubvDWZzj9eAR4K+X6xPCuvYy5KBLcC/1IzAc2utviZasTsWPAHD4Cm9yZEr
LO/K8EpxxjMcZluEJseKsCREgiLkYJrwgm+6p10Iew+orvcoNHe/9ABAoS0vGWA4
1VbEWRxaRAL26pjIYDnG2+YIpblhK1sFHghyCBPdV+VOee6DcEXWSDdvEqojGeRb
m77hZMc9y7OHmbgzWYRHyxHXsk1SLoowFdmVkNjSjWj1FtDjcJ9blgoTuB2OHJx7
jNx/ITYSDxft1RR7Xrfmn/C/VzJOFTjztQuQdHlMc4XNCGxbKX6d0vu7H7XdRoGM
q5pAptKwm2Nnk50FHBwwD/m3PvVfqVqHeFiZ9GWdh841phKozZzfvHGRRM5FnScD
DtLF9Ti1Sclky8kD+DJTwcoOpj8ceUJ5+BJeWBKI+YI5DFL+YVmrHD8uHlAuDCXV
Kw01dWUa9WFfrqWgg+zT4GNa5JjNN+SdjkOsRwuddsKIhD2taC7Fppkz+Nio9Bhg
F6rzNid9XiyOZoRuwJ/FZHs5prWujwxBBaH+DKSzmOLL2kPxuGqEpN9i6nBGXqcY
sJS5ZLcZjw39+yTexGn5hQR9k0k5UatBxEo6Flkuo7tGacn/X8X8J5PzV3Jb1n73
n7sESC3JXU3Ay/+LpZpqT2HEQvTPqaKZzaN7jbcS5MQJKG+kDgJF3J9e5JrPh6iZ
9n83bsQZomyod2H2BX4F9a/eNr99xMXSSqmKPDAMZ8JBW6PItVs+vgGvFC+PJMaQ
Wpl7amYmE9gCcvgOP6YzvfXZwPgfTNwmcmQNjWPqwZlAHuYLLbLn3DFWZw4T5ie4
rVNCGWERW7f4BzlS2JnvwycTPMl7M5Wiq+59wDvP8Jo=
`protect END_PROTECTED
