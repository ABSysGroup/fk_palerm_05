`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T991GLrezVpctmRgHNC4MPH6+QigLWNj0h0L227b01f+vxKOJMTFaLldY+bYL/X2
+v/1h3FLHvR/t4qvv8yTq9DcdFPrYtlbQ6NxfcxCtjjKw8kbDk8Y5xoYOC1uljof
T5JWfBN1X8uAOZeWtGDH+Gtv1znwtBR+Ji10nYU1jfIVKwXlXetmy/Qtv3nRcp/O
JiAVC2XDYQjihqq3zQJRpb+6DkbFywcGERhgfcCbDwIUiCdkuYdS+s+g2zzR3PCJ
n2+HkXJUxmbhRW2f7XsPieg4GcMu1rr2EGAJX4Bm2zXfQv+8Cg1BgdKpQmUBvVTy
qa5goTjgKAvblK4X2c/osT+RK8QNbADUk073KqGAEhB8RX/DPEFmfW3tBCdioPb6
1Qhf4i1soSJ8ZPzINj6WLXHV+pJJWbbZslLSq+hNQdH4eY/MOW0P3MShALC7OPUp
`protect END_PROTECTED
