`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZysJlAJz9KDHcZeasBUBNZJ4w/3+/ZkJ5EA+BKqK+pHgaJWroh0SzmPtmTy7ZWYH
ViU+0JqFcI16esP1d5jPmlNWhFkmUPY1aVdnsFUsSL14DIqh1UdYjHblGcii2CTH
GMFhP+bJfyo6v/KuOzExC4vt9SeNjiuA8Gue6Z+PEQkZ2XT8TNqdNC9o3Pux1+FA
mDUmLETaSCngFJaDstKZL/apywSANzhfo7lHptiAVWiBVBfVUQJRrTITVgMnOXl9
Vhhm26DSeD3A1z+gYDHTle4gtyKCbEUnpcyWF6SWvTZDHAQViOgcFP11nwbZKMHC
sa14X/dCwyqgU9FshnS85Ldyru35q2fvLplref4dsk1q9PM00xVo9LdfapvWDBvi
XMxrnUFFAhyv9svpzNLzLuUf86f4fUyOonvv/bDWiBkHBYTjNPivdtF2ImX7JbSd
Pj+ritcPvP0pQXRTHpEhmZ/ku8MwDKTj/mw3KlM7O5Di+2rZz6rqnMBye41pZnD4
BSG+714uSBGuIrNTbg6JMY3+KBYQtT+otYGyjvJQFr4n2VM3jthmjSZhL3c1Fkp2
RvbWabogbDutIvmgO/TzDMqPgQgI8TcFzWTc/RPd/xEfmWCx3wA3dU11Bx0P2E2C
GM0LH2vJHhQto4amJBS3n/xVXWDlfWfw9BMVWFW+tyR5CZJzPnsaC4RT2eF45fTh
4F1B2fEonyts+JPMgejG6PBpmlDxnkQHFN/Bv/Jkv0CyCI4cy+g1GppF9xkIYulD
AEhV6kqWz01OsEEgOfuWaA3gw/f81DglGcbUUcfDb5LskF7xvNQa6MvoC6Fv7Xs7
QzI58XxXlfUlT+wk2V4OPxjK+5fh3ilQ/Sgi0rqqqbrLUDUzdrxYAXZdbpPTgEFW
BnxpPEEvln6Uc2DXywUokMqsNlRs9zpe7lhhBQHfIuu1QdhrkoSNOOUUqMsEj16j
zEt6+nN1AH5VjkbJaRgyN11vEW27wD5APqXHrZnpOG3hnaTdUkSdvXc6TjJOKcXh
tbZV60mnSCbjcVjxNjlWhjvllIWc0LSdEmAT6MTsTcAZCBt7N7TLKD7wlev7RZ0W
IN4tDmngbC5IDRqu2aKdnwxcX5v2EfwaWr3K2tIhS79MQT+B8ZjJ2yojkTH+amO2
NgLm3gVDCRnxFgDDjh3vN4CgaYKcyXjFdifEq/4kxN5umOO48YCAGEg8lagbv9tx
WImRsSGC9ydIpgEIcsw/MUPXg8c8etF2Ee5e8SA2rmrhm6kqWxSZnP2A05AHz5Xc
kz+fR6c0iLWcsL46qeOGEZ33jPl6hacnSThUy36k89wHYiwgk95fi0orsq2kQkYm
gl+ejUPlS5/pUCG7UTYdKDBflj/CGXyuckSXcoUmfLbxmKjQoFeQZQQNorvrW9Rv
/mg+9NGjMfVW5c4XLSEGafVxAe7ETGRArOUapsuVWe10VcvJMcqk4f7uLMoU9+Pf
piRmZ/nRb5I7bwXBsD1b28r3+KZHPKRekiVqqnAr4/xvO1Q1qplRR9TdaXjQCiF+
qUASJKs1UvGaCXkC6LFYN6H3jGspcNV1PE0T5yBer/5Xhs5MCS8p8orSyT0I4T0J
15xvU1t2vLMLzkrzdY+HC/xe8vvHdJqXT/tzOYcTDh6S0x533p60Gq2T0oV7AZZ0
aBDZBlqlmsJ8Ho4Tjt63KGjNbf9YYNVBz24jLS2aE1ojKpIKfNjmglhpj7/uJKwK
1ddDJYw+Esw9VRSCtei0dM4jgj4U+L1JqtnGReG+50AkzIWSgNmaCEzkviXEs/9E
kL67c3YlywtpjoZ+HIwQjLCzs8GwIUl+SkRPHPMjB3Qp2YmfzyseJMnGEt6cENyc
F/DycGvhW1zoGIFiazc31bHtbxg5GSwckDbpjjISpErdQWKqF9MpXzOfOAbeU2cj
78fRvf3F8ea0ye009TX+0S9m8Rf1cWiZcwvVupT3KjJi3fX+uWTfFszW/7HS79GX
785kbI8lzPQdvhV3830o8QoY7sAeCuCsloyZbYYAUZwSx4Pf5kSswIdflgueCXEM
EGQtRNNl6JE5ep3e4F4YizskQfeoEHCGQNdRhWTsMHGIsXV54ku2xBq2elJrlQQt
1uWKAWmpE6gccrM9LFVwJcswyVfvTx/PkrbzTdmf0Q2T8e3Uyor6A3Rrs055SAhC
a5usYkYDzimdN+pPYcmaw5hTA/8TCpzsS9mZ+jlHPeheIzH+KD5U5FgeKB3c+Heb
h2ZRKluPItaFL6x4eFAmqeEPPVUPWyB4B8IYiKZTmFq6QB5GwPc8sLRvHwjSxQx7
pZl41L2C0aCmhow/TZCdUK7ImSxUTuooYABky+0tsvgfGpxLlRmiRiUtbzImWzTf
VZhb7lU4SEcQ+S0TpiRUtbdnZ1Rgp8LVu34JNbbOeQNvbjNurYUlBx22H+eGIUwq
zxLrXMOgSh+DrG0I1Zlot92rIc3dfH70sFihk4qnWaFv9CWoEBuUl/Qzy0g6dJh2
UIw3a6uky+etphsBV52U9qDjleLfvunAL2eNhb3cCrvQ2DSDgp6xXcQB1oThnxq5
xBb33hDdz8JFyKclVxZF2a5aSN2t0txb3BVuwNWiPIdZlB07q3XWGGU/jtf2QA5f
/FyciNl4WJUM56VDwlg1vTHAzJtu4jC22Lmn4ofXTrDFeCSoo/esorl30KNkcqDr
zK3IXQCsujlLY+VwRy+IIooew7Rlu33hdg8tKsM9d8LDGJoplTulhLHD96SOgPMw
NtmzKz2PnMmNao1sjtnvvkTnnLtvTokolTC6JtYk6ZQZbG2TKPIl0Qvxwht4md2/
pKWuotqBkbUbQGzGvpcw/QNeZQvdPQElf1CaSih8zBKwfciCW+m9/i9+/Rf6PAdo
6/I6XULQIWFZieWlAyC+7gfpk3u3wy+Uilt/EodaNhHI2OSpD6RyoimS76T7d7kb
3mOaoX/NunBjG9dzAKoaJxYL4DpiNjRF+noLFjsyA7uSMqqvmcPy9RUXK8OkiloU
5ITwpjGg6MSYDh3q2SMgW7qZnikg+mcUP20YrnLQV5DZz5nhFPpqK1HIgIsbUeaM
0U2dQFEPCPXgF7900lWbdNQSVSLoO6jVwDYDYREe946LTUpPCb4KbPAVHpCtBWz6
oI1DA26gctnVnq1EWgRRsDra4oes2qgekYlQP88uaK4STjIE47u56nnrPMRSERzx
aIGRtws6fwIAaYfbRcbAAkKGm1SLLsvxSWkuext2HoICmZVu8Tv55/bRmP2WtOzi
l4RY/NsByAVz75c7YGjGDlTHezNJ1xkXbv2m4GrXOeT1ABBLdtRpSRezk/q62hXc
oSKW2MQqsl/Fajd9vpVMFZg6Y9QtbfHWh69B9DsT73hn8QgaWgqjbNF/vI2AjktM
ZZt9yLhTFDBaTEXj2N9EZxnzw66nPtxHx+5MOqgBo4syE2rNX26JKbzkJyen60Dx
04lk/NRANZrSZkdkczX2qeJmmApCsQr9NhJ4CDBMosXSZp5AcbVzi7AF3w08FUL9
/l0lx7gzn2/vM6qWx4Lwq+0fGhnBXK+sLwpXf5ODzSQYs0Vxu9sJs8Opdld9fxoL
XIFxJp2HWg6TY44pdluM0W3Yj5ockQsNJ+x7yqLdq1jP9Wcyafyse6UtFwU+1Jcn
QovIoXhagrokuCm1srHaox+V58mT9aHalMQYotR0RNaI1bTcdY7VXyZdttJ5haSV
JvDiT5drHHIJfzHJaDMaju1VP89FZvqALGFYy8NPRGc0NgxmWJ3ADXno7fMdjutk
+3aquhlnRxZ3KdkcUhw+AYy2xaEsqnwnIVVp7GidGXpXvuvKF7s/Xa4KIkxCSd5Q
GCCYEaVxQOuFw4K5glLjIrMKmwrZOu02YTLmZJh7Kgd6y0uf99Mk6ZMdiHBypWXI
yOof85Ebo8UHZDcuT2VCwUN6tmabyoq3RLD9VacRPc5gf/MJ3znDlDVYWUjwagin
pjy3dU0f60iLcu9CQcU1y8I0UQ6WYjYpApyenjkXDmq20bWxO2dEzsgHMmdBEOKt
Eq8x/G3rP8PWJu9uQ0+SzQeZvz9oOJ06SYj50ENBnlxKGUVxKsdv+iIrWPFlBEww
LlpiNI7iR7sm5f337x/ms25ECj0JKKzVfXYbjfbsnnrIA7eKgAE8Ci2Zrtmon5Il
oPPDlj6spthgwLTcWv3QdQaf6dfTqCjIPsc1SHb05PWrIFttyJ6KCpUm6L70fkhp
DsMkXFYNinWB9Q27tL3lRUy5ke9rPW+tDQqMbxyql9J3oYq0UJ0Xhmydh3Aw6Ses
o3ePMDBmuAKAGtAcyq8XDl7RpvxLObPaTBH331bEv6I9lMaMmVck8irVB+YTBBJ9
49IdJF9RxNakY3v/kOWITf2GpPbum5y8gxBLxW4PbhyRI3WMF9+RIvVYO8NDOYn8
VZ0eYCAKG3LPDrUNp55mGwFa6eeNsfKR3lACOYdXIyGnu8c/pRTtA1176mcoLR+h
2Dlvskdv1Z+X2Se5I+ot1u5bBcIDv6cTqzTGBK4xhKxYOCYV23AQkbzV/qzNgt50
T/RnmeIhGs3hiHhU2EEh1yfuXtlwcH9G/dKoxgSCRgC3wrukUnsqFEx5VKrIsdqi
EcSv6OBGXxggXjgaC/K1mh0zoJEHyGD8LBM34quAyorrfd/wDrjWOvp2pf9tefgM
0DPu4P32VZAWmieTWyXr9rZ8zCuiyXWhm7G0dvT5QEkJ46PsoMeo8I7sJLeaaqxU
nT9LZLXCTvLmBLD9EpesnNSx9Mbb8Pe8G0iKHlUjGT3MV8YApn27TQl1WnfMHbI7
aKH1VsZPPyg1e4KNGP11rvQdjbfE0HlGOs8hlmEt/TEjU28rrdrGkfTYB0oi6efx
FrljKqMSyNyiWtlM7U0fwB3E5EclYIXUkX961zWF4ltxlQDlPEwwFUXBMEXjc1p0
Uyv1isuvA+6mBqKmY8aZermgtuTpsLSy/557crEgK13tDMu5xS04xuUemRtnaFav
DbxVUmKbGlg/swidGwk4d38cPfm7CFvCFfDRwS6KjPyvMd3MUwFWWRzk2ZUOfw1+
pThp3HE4q8Hv6MW0dHbd75qjk8HOHdqI4k2C1Eg33Md2OcyvSnqY2KehIaLRbGqY
ql1h+kbLxJ1ijivHjQoI+mccHrV4XzscSBgidE1+V5lKWwau7UXSvWC/dLZvUwCA
60MlVVuWkeBv2CJVUP3pEmyo3D4VVoLRtLKunyUcLaoqrpuEOibfmkuGKkllqJ52
+xmB58XoTyEGd1gqZKCu4niSR7goqd0lMwGY+H5XQA+6qlpywETTQB7BJ1Wr9l7P
4E2N7pD/7pUmd/oC6nEyFgJqh426v9sccEIWDklu8ssN4qbmxGTz8YZtulOWSHM3
coRKOSYtM5ExFilSrYnz5krIvCeqlekUGI1YJmMY2Pj6lh7UaUXUrnNNNpyc9wL2
qLWVpgvuELw7NQXRlE9sVdHjA34pif7T3X98TBfNLpM0Uqr/7MvZSU0D+3U7xqst
ngbs5hWjJMkPosiVw8uT1uC7iWuxwQG/97YIQFIzSXbJCWPJLNrgajCI+mcdO63u
QijR/CbH++/EWnZHNyS3ztMrKSKl2GuWUUoAaZQoQa/GblxA9z27sCZNiDnpwX/H
n+KpPVWt2r816Z3Xfprz9Ei/agdmLm0dOdtvYp1gNL5m/X4gxGqmL46uI587wizx
fXOmHG0LY1Bvb2QYls/plczmSTIZd4rXVCO7/PBO+3SBUxb0b7NrcZoFFyd9fhwG
DV0VbSC5l6hMYfkGQTRxgFMelUB+wcgMGd52LqldJ5zqlKSiyAlmyHwS4Cz++vC7
M/d/SQDUNEvEz83b8LO4rEMOJb8leRC0uK2G+drIGj2Y+ZzhI6eIt37lrL/C6sDz
9nNBrvymZzpxQKddr8bo7twnXrWFwMyXGsil201o6NohXB4dgg+YPdb/6y0sy7ph
gjo5skUcF5CQxF6oPK/3j0MSN2SqgduO6HRMRyW6GFza+greVeLDGVI4HGKT75d8
WHUCD9CbXrOSCa701pUXIJLyJetYfoluDnySNFix+fwFMU23uoKmYogVYr4xTb8k
UlVMFtgyPxDPwEhwfZeW7CBV6NsUGWHQhv/qo/9EQQQSAmVrgFkriR+CPAY2/4e/
/f1rd2vCcAtLg1BTVuZ3IVF+bSJs9e3zLaVybwI0nxm6z3tggRA5oArqB8SKue5i
EW5/u8YJfQAbNKL931YLX4PkQ7PyGKe+vx4qyz4klNCOUnTmTYq0asVrhrx7GtKU
1fsiwDzJ41+TLumlRU5vOCHK096o8UNzlTZtBKSCPzXIs2sJy3Nx6ra0vLR9jTGw
OKBVyeE1jZd/QcVPzGobol+r3BWylTxs3ohqaf+qi45Wi8NxRrbjfMB1K3lhZSe5
aBmhJx2YXIbclmaMPGAogIMb8Z3l+xxB5YhiLsHCO9I02QQKqyPeA/6eEUk2OTJw
deZWC6kqRcvz7dpQJL3DSdQGZS+I3CkVW+khL3oWzzxxM2FYpK6zziWaiMBEM6yO
cPzdulgtZXeAheW5AgNdxbzY1smIBJdK2A1wlGvRWZvqe/Gp7gUTb4/jE4s53hMb
jMl8sQtAP70ZNSE8daCkirztIhwxdwJNhik+SDy2v6aJa4Tlq+lGlkuDDfLW9UBH
51c5LS3q1K5ue14xgb7Of/Mv7jxWotn68LuGSefTSn3UPuJHXY9m+WdSJzHOIjL1
IN2d4pQbjTtvbOmdIrl2zlE0t5qejyafuW3ohSiKn1oMXLppo17dwTKNUSUFK2bc
91uEl4/Gc88tG/buKyzZ6anky6FLVm6a8+UJ4VZHxaFnDFzc+qsIqid9d2GOsI05
ZYRYdJplNOduckSRg8GA9Ff7R3o/4SEs2Jml+j/a5xstHIf+5Qitj7FI9mvqFg4X
mO5oA16PxvpmnjzCQdbQL8KecKNJfIICBecyEmkDKBUa0hY6aBlFBwYYDCUOeSxs
SE13zF6T9wFv9LAgtzx5sRA7gcIZov9Z5kBS4mWsKoEXMBjwwaEQdK1iJLdlLNmg
nfkIeCeh2VzhflsMu3ZpAILZ8dH7grZdNOaxx4MGREzjvqufuBW9gAzhAW/DuMXU
Vd9Ae6gzW/o6tTYPO2EShYMLwg0hp83p1kwAienIW+p1kl+9L58L8TBaB/QgacWo
RiUM14kYUbty2VE8+MqGiBn+c0MkTHz3DH/2RLWZpWCFC5hTRDRe9Tsl5b+u3W3G
lgDp3tlRTnkvsr7VAk5+fYUSDegvQkBjoTvsBGlm/Q4thoj3tM0n4z0toRMy7ipl
2SVW1nXJkpY03sF9Fj9GqHL667WIqaLoIrE+smnCyV9Q++J93ploCXyMSA/eJV67
CA2xbz9YRhhgybEklk8b0HBxv01/mCt5p7GPXQPC9E7FHNQnudfLaVmgTiEcWHcF
/X3hAjFd7+Di0Z7022MSrl3/PoN1rrYGonJmJybZIvFklgwamjeU2QJyrH2Nkt2L
ELAMdlo4b1V3epzOZsdDkkgXCh/a3SkU2I3UdLIrdNGp7nPxqRQ8UylokaxW3BuU
1f8jo6VipcKH2dEleEqnHJ8CBVeNMsmXdU2b1Z3sLx1SZXg31TYXaObfDEx7JgvM
Wo6ChKlWUcjNg2VqTnUAZDD4lKT3zDroOCobNFh19Wj2vuihLQSKcG3QDTMOZvaa
tiUP2wPujvJzrFdA7ffulNOK1aVo26nW2jaY8ljmsyDstg/1ZXm5+995pHiuj7wb
MXHwernakOtscSrQ1OVX6W+KvAH0SghTutCZql0OLM8iBXEQYP8KX9UhOCySKfG3
dOOycpsE8PS9dPRTlrFAzjxc6I8gKRvRvapA8P8U+K3Vc5dbR97H0nL4SJol9osY
XonWGOo44PDUlIG3zEsziL+2C8T218qSnJQkw7E5nCMWaVpmZvlC7wCOJ4b0XFWQ
zb4jv6sLE/H8VLdGbwN/ctHJ7kN56AtpJ8K0/f7dgTwsa2LqfWgNNqAHeYM/8i4S
4HFqUCYrFV2mOekgegQdJkN0oTabIpN/cP4Mb80CA72pLTwzXH3svWoD7stmD9TL
Rz6HUv/mumh5dIg1kNJhq719tqTcDWuptM7V+xupvzRHLVKQjDIG98PsOURAb7wF
urBAGfVJLtq27/M/UPKQhImY9Zfbu1MxX23kY7fmVx82BMs/KiC55yU+8+CW8WGQ
pnBLdGpJW01otJSEt6cGX9xfaww6nRF//2QHZm3PgTxFVtFOE+QJngW8XqTYhBOc
O9VU6Cb4GoTx0mhCNU1KOm/BNIjGZNTs2cTQcXJz9pa58hpt23RpaMUef0fZAQL/
aogWMdFvPHbd0GC0QFVrXDiQUPaadm5O5pQIDJNMbP9ashSr01tSnhmuuDQe09iP
lLuIHS9rX2ROdPALPCqin4NbfBZktL8xBZ28qoDqnaGwKdl8Geo/BpcCEfbMwafe
+jWDbZFKA1rgdzgmvpgX/eG5HrNN448PKP9L7Zm5M9MGF2Dz5oUe8ii7EUHobjLh
pH2MhePXILFK/jn4/yH433Q4GTruIAUmyP8JMUQAYaOkLnHQ0101SW9WqV9xM222
Y5lT/fGoQg8FPeqoupQ98qYiYhn93ZThW9Q3mOVbGw1Or2glrlhScvWYU9MBRRAO
vDjwKexFLquaN6f3GL3MZpjPeQl4+9ajZHLiALrZh80oXwLIgQp6an40KQxsmTMM
MG2raJEdFI7sCyT7Z1BVRKvpFzx0r+gtjHaXJMN0grxzjIrjQeruUA1rjY0G8i88
7mD/DIq3NxUwdaN13bz+VFPQRM0cxBE7yY4KZwfpnjASJSPWuO7r8Bacf/S+8iei
lMJAnt2vOVjmyQB4sdN2q6IFu8qH+zbTrU1KYhcZT1RPADPbMHRbJw/0KJsU4H7u
lQ4x35G5f2AgnvXtHVKi/JGpHthzNO+0UvolDroTvv1RA3Vs2jKS9c20JXSp24cF
QZZr+xq/+KFssVQrzr43I/yOb9RhcshOdMek8Jk/pNs9k0aey5I3bFETpBY7PK/5
IwRM2Dwfp6NiU1JabarkItqnR9eWgNUUE9QtzbanseWVoFCarM/LzYJ8BK0YxbTL
MIp8YHf16uOuTPFefVIyf9Z5ODn1YCV9ke9zsTcA2T1qbjuli76LYnB048403s3I
7E+X0eznFY8J6im/8EY5Og//Z2qOy9k3iFlvrr6qRIozuwQAWLUB7aO4b0MMsXdp
DJ81qza/DLf6/NxsDikX5dThK3nCph4WH7gW+6OokWD6OwPTniwvWUbW+hD4nBFV
iZ4H1chV9q44BWDVZV4iEsWp8APu2zCsVrxYkoWaWf/4fklkvkRbLCJkCoyGQt6L
zTk0niQ2ngxDG6ryE1w5aeVLeSCxRws5sfjQqRhQzGts29zEGNyM6vb6b1fJnds7
RNuWnJnD0bbaPwNVnEXOudJFtvd8L7BVIgVwDb0klHTnD4WLEKFGBqrAiLhqDEpK
LvhvBY9GqV+5vaeanWyz00Ocqp4IsTK3NGa33nriKDUVBsJWkOgqIseDrDCn019X
sNvudtZYGzXs0/xogEV4EeWfFCzcwfBWaIRUTZriCF4QjvH3ozGQlEpQV6SOs35A
4pnQdOR8Cr188Duxx3Ujbl2K254PXriYL4xICOeIBbbpVxodYDZkNEaw/IWtdmCx
zi5WEx4Ky45DOK9kAEDjjFz+umw2lpSZT2FHWmlI4vY2oVe7zKiGhTU7qGuUsQ2o
/8TZkUdzqQIA7Oqbid2SD2eSUGg/Nzyh7MZugde17MwH360YWQBBOJIDdDhwxEtG
cm0A5X15aA/iBBNQg2CR10fVHQmRmgK7AVFjGF++XS+49Brwv1JXlQvOwO3rPKcS
leSMntWWKUka8PfRu0AzRJpemSAUeCJU5u/DS5CS+Mnn+Kq4RWtU45+ev2UywGkp
ntmAk9QfkmSX5aAjDgkYHofcXGVZt90M4Sk9Edcq/DJNgJMyHZlwqk1v5REspVeL
tC9YWDntTh7oIfPYcShzwo4DJjTo69YRu+aRSTCrNSK4S1ApERJZ8dkXniMqzRT+
yJ9uD65lV/5+Xo0bmc/fC45agI4z7Z/Ik89DmMHAO2L25wS6+BxFXcD7m8SQdNnp
TIRU1Q8LUS0cOuVC8L3QOSwNuNhHBtFNP9BWhFTMJ266uSZt+5X29DgdwM5saQMU
bC0dkrxAGg4luOpzCkmR1E8OKVelV/UX8xjQ364Sqy7v18RWTxVbDlZdtYKRaWuD
EkcGrs3BNIMT8bv4PnxtjhgWFLw/SvAN705mLSDIDLAd5+ZLeNT+wqaRcGOMBpQJ
QhaGflxYODHytw+tGy1kc7pYxtjlQORhTaIYLdSI3FYTzZq9LSyU/kJL5zaWfUpR
6U4keprsMBj7h3z1xSLSYq/IYAFphWhraAq4Icumciwsjooy8qkICA+IDNalmJMs
CrExCR1+97KPPy+iSmQCpiT++tn4EJEgWIlTsBUmZz6roWRuH/sQqUgYvy2yUZUB
xldOoykuS3KtXVP6KJyryoh46xK+BPFzAv6r0Ab/dBVeMxAZn7FsyJr40q/kPHxS
Rq2aqpgKw9qYydKSAAgM272RQivIWs36A7H79Fj4YIJAPg+ul+HCjvtWjmorGFJ2
sadWc5Fn7dP28GoPppJGwbiwWGoncVgffi6+xNMgbFt9PjP2Iqmt29Sfta3G5TAT
RMzYw7g71z457J/pEAGsKaUtxgh0Rconi5CvAdjFgIhgOBFxg8DUAYp1keGqqyJF
BqIHbJgTbeQtQUfwfdrbGQYYM6UBRU0ZKhDOKs/nTeS6cpuaESJRQHXApIKYftvY
5gzaFFNMUA482+V/mW3MkZXq7QooO4TYlJsxQfqUMdn1pk9rzus0o6MrcL3tCsxJ
Q9ZJVNVJ/ZwUS+tOjvjjHYiGlMlNFY0pu0hqhed/dfFmTMprhfTJPNe5XpZVlcf3
kxHJFtJP4KtqNJOk/lU2NdfkuBdYxU0U8VwO9u0h2ZM1Ve73Gy2f7m4CQJXikWo2
L/VwFX+sXlTsp2y/TiuZiP5e5VAL3FzAq1ZGbCTXFs+4QiPV79m5aBOjmPhWI0zZ
swSydyJREUndxEdnRdqZgH+U/Dnna+tM7Pt+VWRWuVe7wPpku8D7C9oyIOo5qvgw
TsCDbRkx/WcFKxUHSFBoGeEsNTkSSXnVRFyUytDV4ILdPuq/du7CBoT+ilTZLyZH
TIsjs89vlOqYtIM4ROqXZRmMcxAQvWWIef3PvDqL/Uwbkk7bjURPhVfc7nZ+yZdM
tuN9XdW45p+tRt92vTdwnnPD1BAZV82RH1IdbTe57tlukIPtFHeuqR8baya8YOlm
r7vNZtAeJSybIIeIbO4vMFrbrFMP72o0rhx6yt1piugEx7Ml7WNPu1Y5i9QR5Oos
Ppw9f/qdpDsXRf5Dtge3PfB/nq6qpFGAa+9zIYSpPkAVu7ZPm46GuTGny5e3KUtM
MZMmvaDBPuhGlm99PRBXBot66ggJQz94mMOr4jDamchsV4Se5PE+UkeZ1oPRS7C6
TLxki9mnPTpj4odfdGG69WFLYjbF/t8h9pdW+h3UZOjuGenda90EOwBpt8NI8ljZ
JWQtLEWmsJtuJEVnHFLTRBrteOROhV3uEBw2skfeSsldfkVY+m9HCsg/e8x6RQ6j
xosc2nRL0JT9cnBhRwTAiNtFGO7zjocSmNqke9XVK2MjJC4C0N+suHOYlHDUagOV
TBQ7LfgO3n7nG5JJpwqIgrR/kmVGRWnXyXylKqsXicZS4cWcWJBRovCxZ/GgJW1a
yzOMbTMrQcWN+sHmBwJLN9qAAAr3wSITfHGL+s9tCjhkbWPuWKYbBCYX385SjesG
WjsDTH0EPP9+85JnZ2KIde+PIcitGwqdRxPtw/43DeMg7r6acfz03z9uu0W/5tOA
cO6xZLWncaXWPxfbRovm2dYXNAG3JtJm5M9486HJY0BElqpusD1WIY4ESse/ihJP
cpQZTX7LA/gF4Y97nk5WwFwt0DcNk4D/iqxKphyQuttWZb3ZMq9ecDLivHuJHj/i
HlpC7iZM/1kj1UwjVoUARV03fOBPjG9uU4PFefhifhEjoM0DP+yPMLKnl/29XdS/
l85rQxbzgPGmJJ6obuHgZTFJFDsrX5LBI04E3Hfa2DZHeIvvmCgiVecMu6xlFCMU
MufhjodY56JPELsKMEXW7uXt9ggrP0dWsbRfSB2WD+ldwuLE8Hi1bE08oGAZY7On
PDvTS/ZVVv8k5D1CUcW8QUSqHPS+MP8s4RFsTze6BM591Y7uOP+QyBSOWJxyyEIw
+iVTuKvqPjDwjKhqhtKtiy9Jta+nG6tm1jtUUEx58lhI6GeTN6LF95yZswJ9aANV
KjX74tzEgLnx9fhtktegsXjmNPMrzedkKY8XGn2+Py7BoZFSDcItjVJiv4+LzIYH
G2Dvl057W8hfvUVJGkjnCXK2VP7UyN/kQ7JgvYvakNeutpsDYF60vg3I7ohUbKic
oBtJ6nfjE7JW86vHC2P8H41hKN/e8EwpxOJrjHXHTn0zqxqvM1O7qdb6gUmphLSw
E3KPT/nd9u2ZhtKS7JS3LfdGWnvCM1MYxYGDQhUQbWu/IW/SyWK+RZNuLzPRE7Hl
UHOHQBYTxtk+9tn23QkQ4GPytgY8lEXP94vt63v29DTLm1vQCCvFaVgnJFCEIYZ+
UslvmFemIykf333ZT3XIZps6+ZvEVPIymEGLGbHtCPILO8/K0TgOxwmAODGZMCU6
yNideA5+DD2274Sc7s0Gi7YPdrazv0jvHDfmFfuFlE1ZoPJupbbj5FIYdlW82x6B
abBpXj/D4g7bny2A/2WI9g7cc+nqDbdrbUYCPnjYk6HRk4NqNXgqrXZV4ZTNFJO/
2wlG59ii5pRq4Q2Onk2T0LEqT8Q/xFNkSXmUHb49inlWWzoOprdUUyZTR+jByQ3A
dIu4TT5Lb6WqZRMSy36Unptl6CVlYXNfzlB9EDKb6cgxSc7Hj6Vr0zKEn0QH3y1/
BxNGotfYfugOeF6WcIUyUiE7zEhifM0KmpeKdC2I49MTLpRfKWoAi0XPaal4MyKa
j6hF+iHegN90YpJGa0REg+ndn2j0hCuud767MvHEDgTVlyTETZbRycQcruPVg3kq
gP+QKx0JMEaEiXJPWhkfytQPxb5TBYqREeIX4Kzo4BTecTigzIBdde266pYXV2rg
tx6i5dCweq9RdU6u3YFBOYXfPDxfkC+4ENB07aANkeeteX6PtsF+ORYgr4cpgkVO
6cwC9pFz3zSTsR7R2g4cKqFIOlk/GZCQQ/vkGTYGYc95tE9uJ+KS0cFsaziXi8Ch
xn85K5lJTeLpupGRHwxrkMmS338Vu+XXfnQ09xlNh1FVEE+5w6l+Tq+WALL0wkAM
np3cq63FyGaFFDzTYrMaFFyr7fPhK4RrhslwEIUmoEj5HsrpBWSnZ/2glBvcgFoa
sNmuIagt2nqQRHa6Bj3ZrYDYdZOte0RCg1QkswSxZfIkGLbIK1x3b0g08RMbcOEd
KVrBNCbxvY1S8n5NLRtIlOpcs4sJ/qvpRtRRMSS8X1tuZ1M4zPlAkfjRRgLm5ZiU
E8Wjo3YWA2oOQfQ5gSkPyvJ6bXrNcXCzwza/C98Q/XZ4GBrRxZdICN0SzhZ38KFM
QspRDiCJZgqLoHQ2d0tEBVcCkON9OzFcmPaWTs3VabQdtGFbVF0sNarVv6Zjm7Z+
+Okl36zdybWhjVlDK7yWmwQirHRVZtXJB1mG2VrY5QXbGjLN3tKKNf6FtdN8tgvX
7exK9Ec1M7nuLGQBJJ3zJotAtmt9Qg9sVnISRnR3X/1cSt1ijL0MtUYNw8b5Ea3F
iqm0z0A9FS8R4iLa4NJpE9V2H50oiCMqyZEoif5peVh6oIuKqGPDJRjtA8YPzb0v
6Bj4SGVVb+R/E7L1YDsgB7L8g/SQ+rolEIzJAnuhM4Ez3sOuZr+zk1s7G/s25mzN
zgAE1Yt14qxkIQOPCH5/oDuavsJl7g+rqNy3C23lPmra4urrQGbcStSNbaZE6l/O
VbvF47wcsWsEeCUrP2TDYRMAo2ztkZiEJ8W0cC3wCU2dqJ5+sWCRbLo9p0tQOU6d
OtGRHNQAlu6osr+B8XQgIKpRm3/LcbzhntFZ3XZ1sImJHsy0VnJCaHvhovs/2izL
OQoS0PJmrim1TYk2gKItl2t2UUjsupXboTFVeSDLN4RDCCfagM41J259CfYXhLq9
VROHFWVJ04Cz4Xi3/2TBgp9HSd0dKP0uLzbt6cTiY1gq+PKbintn/Hn+ec1hDgvd
mAuvZGKJSszYA4SIh/DGj59R6fRkr7Em/Dj89Ih8aL1UmFuC+THQwSVD3350H+rc
yDUGbznFcStuCgqDE7aNO7Z+Ukh1Ny7oYRpKDRDuCBTBNem8kNMslKvBTrgMmwLu
t2tgubbSxHFEA47W70azgoJCKHQMddVxQ+0SGJ2j9/enK3T3wu4he/DEYlj7aNC1
vykzFhlZXpy3jhbWAVUk8MO+IftxM1UkSCtyG51E9WfcExBuoj62r0GYBq5fFImY
zm3HOG9xqjrurHG1jB43hffpUjACBrnI7XvmgOt89CRhuKQXg7cZmvUG615QV9No
VFiIUDuxXRkPJMZJGsaOSHSyLMYXZi7eUOihyj9a/1uVRb6XZfUt0Q1U35b3Dgs9
g0tWdYZ3va9gHjD/EnbWoiC+wijbaCSAAvvCn67R3WqoPawns9P0ba3GPIBv50Yk
RlcUx0cn9TfaLqpl6K5/si0ALj1pDWVdHGUpdyeDXq31Z+QnQsYVW+OQ58E4h4rj
0QWP/a9crPHCMev0e+nUIgbXv+cLUC44LEi5eAa8WpUINc8Hp1yC2qfgmaz/lBWu
VPm7Qt1zI2PbcydyOp/jZ25IUyvQqtnvA+Sg2qHmdRTjjnv1V+VqInhNBlN9fAiE
jIWsvz6LY1r4d08L/y+vCpHzrLj3Z5tIIvRV3hoza/R+UHDb51BKfjcp6ZQF5LM1
QHLibjXIzLerHPoGOrPR9UGe+HqXAVi2UEi2U7ZyybO4a00RzD6avLWmliPJQNNA
WL1n6lUBCbNZWEw7W0EjQXO382Niu8SDm4ObQLxsb7+OScViSoq4gkjl1rQb6n0z
UfHM7SIuFJ+NEjkvP5GDhG3BWBSJtr3u6vOgCVRzS5kadmCMu8+jipfRkcQR5o1l
FpPf7Uzm7ZVoDSjS6W/gVTauSIP/myhqGjpJXJaumGdCd8MpxZ5Gh348/i4Lni2z
nDNA4VsHfOiLgYstJOo9gcEX7UvmhFXSznja/IMjxbdeRKVRO5Xh8CKEHJt599s8
uaSzCfhydBGG7SxRvyKJdAlivZrf/ANZDaP+WSMANb37ZzeGZ2ON65X60j6UOFpl
nFQj012S5TLdLROSMv9E+YKRJ8Mja0IzEFKGXXFlnnt51HlLejb4GiNTUhYfOmnf
4BWId6eECckJlvwJfxb60bPjUhOw7C6vPIWX1mTuo72BLDDsh/9lDklMsNz8nTHD
yvXYoLF+bjEODjaQ5MqEJklvT+iedKd838Yc2PzaukNn6XRaOub1n5QHi/1KX+Ww
vygEvatVo3RqR4jJPxfEESuILN6AFY+qBvLibs4d8e3Z8p63E76DcKy5clZfR+JE
NVJVdlh49aD5SD96s2JHZ2xxwI7CbtFUg7ZrVdvUwN30+TZFCUuvUCZ2hURtGrWa
xwPP+3GHvVqqoVyROe4diQinVwMWJV6JLPG/Vs9RCAXvrc9SoS7IkHr/AUQpKXwG
AhkNMnbOXmROHOO7/hLbQYplZtE2eajTofZLbu+ICYzYVP4/PYlVC0Btxt9BwKAh
gVr3+mIiGFk7YxJfOxgeNNVoS8XgVq106JiYpmxGN7MXDkudeLzURFzYzpY5+HZY
OVqoBA+iX+xbrl4k6AbpTujlXCSzxE+ciiKYe3bjeedqU1BMvjgz0bdXXM+tVDQn
anBS7H0864FLOiQbXEPJelyIDn3UbmCeqT+Ood2b6FOFO6JLJ8JwDJHjv5XTwLVa
h0OAunBajg/AZ3Nmk88wytZJr1c85RGSqdwOAExHzIDCPozhX04EvEqOzRN4gFnO
y6nImk7p6dlA+2hPBFstd4io9sScMdBJ7/DzO7/Ic4ggb9OC4j5LVyCPs0+B1bGV
uZqg76oXGDr9C3d3AJwsQZl5Ah5Wf3xRi8PCcG5EUnurzzDVKPVQZRSOy502yFzn
2nnpOCwjHFMYvk6ArsvFRLKK8urll575MLoqtDjD8g5SDVN578qxaLerMU+/8/l9
mc0UEx6xE8H3JVGMea8WlabnNcNu201aYCOhb6oKKa1mfSUFNxC/gdP2x+IPPNhG
Y85hiHenDerbckzhUe/PUOy2Mzvc8UbERQMWQWp3q87SKGFYivatAdj7ZYUn6YbU
bugTMok0Q/qcyr/jOIJB70RNms6fXfKQ2Vse2sXTddjwtLig0z7rPJNB5PlJzZ6+
rc2kqmAvJjN1y+lJ4kcEmAqXE71fGEMSopdkabRadVgrJvFmzGHIBwfPOKzwZ7XZ
XrK32wewNDdPmLRB+hASFwKqBRQiovkAX1N2LdMyk8RD+LflQo8ti2wnuC0k+wND
kOpFIhFTzRQAEsF6kZZS3mg0XDbPoE/eizZHs/fOVMMDvmuiu2AT75CfvsL3xpa2
MXxT6hC42L72SEQhg89Dk89kvHEaygkW0qDF1FJVJBnJEsTuZ34o3LnK8FezSWAg
B1vCJglahK3SH86dSf2g9/EP8GUQ6qSHPCiNA3g9+Q/4PX61nvl1jcqjCx7xiW1z
KqT7kW3C96LllZiuoxx3k50u1amjhXfY580yH3ZdZYVzsI3afg2x7xgfLeyS37lW
Z6VmYcBebcnglNoMFxGOGqhr9XWnE/NDlTq+WIk826i2wdN/bWXYEk0lHFw/RfMu
bsDGVYwKrjOtT04HsrZJJJIR7PHt4/3W5vypRleP+YbdMBDgbcSoaELhayGE6puG
lsLIVTi6O0oP76jBmLFSxTLVPr7C3nUEeTNZ0XN4WohX0SJVGDmRm8914L0lMgs0
TDlLOQhRyrfH97PXql5RMIci5qFDUWORgw8zi/mIv6uCApU0NwudL5e49oa2F6wb
cDIGDdu5K1ITwPgHqooDCyZlXiFT4pluvBznZ2EqWVrsMQjpZ6qfxI+vA132uAey
FA2edMr/PoieIWfzzpofU89mZfE7pY5eobgV1lsBRD0vc1Nzc47RSycau+n2PkmT
aa0E0xY/L/511vaJvb5OAynuDu4Qm1eGGXuH8d3FlrrQ6i4GtZi53MJ37LEwObvX
AlObp1qCQ4H/en4ZK6EplGHtpfEDtu9dpnfXUE0mvvT62yO+OB1IF/Tz01YVekGb
sT5/lRltZvS9A/CxFnr+ewh34kfFB/IVXbOkPmTZZMTFiaJR3B1aKsPYO+cNt9kq
Qs4EgqhdoWGSKtkM77vRsIseEn9PWKffg0qgZ5Mc2xD9H4A/ropsJMOqx8A8QleP
xsOmzq2pcu8Xx8r3KwMoAQyAVk3VeDbxo/XnsGabNEE0wgs+c1o6oILKqdeJYZuf
Uzv75IxdjVzE+1N2G3GgX+p4bPmgdB3ZLzeLRj7o892yb6U3gXvjnaFaZ72anzBH
9EkKZfvi3sQSWsKhwV+FiHyE5BGwJ+gb7+r/0M25uMbc6Jgga5Obh+aDApb3u7jy
DkNt3iy6di9UsvwMVgbYf3nLI+Qa1Z7KMhSOZZqiiyYy5HxBv0S1pXR1C4WTImRW
FO8/Q/FmQD7KGv2qS/xm+7beyWf/DKsOn4CLrFuW5Cq4SsaVqwC3WeqGWazesS2S
MTUzTDeQgHjvLPf8y5KYZYDz2pyygrJuBfeDjFsd68V/VNJqz7YHaolyvKe0k3Nf
ou2CHsZUsEwwYH2lxfe4TLA+25H2Zfj0SqRNXn5zhxNi6YqFAsohdEDHBLBNbVzf
9zr6A8ASIQWM6Vn8ip7sIipxg4UpYKQX+EiUaEdqxbahCvRQ0kezVJejyANKMLom
wN2aVLdN1GihwLhrt7i+U9mAQDiLO1alDgD1hsSZASPoqMo9B74cuSkL8vuRjyT1
zrBsZ8g71LQoKZTEUTVUqVe8ovBj3sITlw0B1jClz9xqgVV8GWTOeTRIj60kLYi5
aRSn8+o08P6z2M/2pTsu3E9TbMeLfQTg/HpoN8J3/hw4mWToq/mtuk5lH+bIHWqc
//ZHN8pEGsHIBQx0RjoVvKgjnqDv/afAQTBihe5XALXZi3o+dRyR+R82FZxxGv6C
wYclV5pAOx+33+ATlb4WtuhGiPdaCdE4AvDktZZ2hQ/a09UgsjrXjOzMCXaQWsFg
g20W8Ue801XtY7Nlbb29xGyud5lMhlt8cIjF+X3EiWQU8Ra4N6PbbnNyEO0+GsDS
B/XdWjCRc4IX9gerANPdJDSF3v/Mi8GQkmGUuqUzyIL+3qwu6F/VwT7NtDvcWoSn
QIdxbAilh3Kkvy0bzn0JqCLEWIkN97gShat9w8mOjUcjwhGgl4Br74Xnq3bXUklE
H0x+M+1dQO9oVFJI540mb969iZpcY0MC0hRw+s0+MEcT6Z2T8FN6fSdnqLZUS4bf
1XkIgs7N/Di1AhwUOlw8hoOu67IgbRQXaU+A2ydlvxnIxqpqrqGRACF3+ZYM6o41
zlUGtedz2aeexJy3fqlfJ9optUsvPE4oMMFjR7O+h8eTuwWgU6hzdZoQxtZja2+u
U852Z/24Cymez9Og+jUeAJ4jy1Zbz1y/WnIi7lIjvOobUbn5HRMWxGBeDE6qUImh
svb60tTUJ8bqEXZXm9MyhtRfGL1T75cgQKJvGKp30ZTI2G+D6i8nipn6D5/bJ8TU
Ul2jNxAS0eSlEjAzSI5MtVmtBy+ZhBZGfbJAXcm2PJwmf3kCi4UsogIUnuNcC3aY
mVTdPM8/GAcEhUuvFPFtkQQEyoazDCt+W+dL/qZ9FNsRbXIEXe8PfJsddrc409+t
Ldqb61OxRjBcj0GeEE4grhYInqDmOacPcK7kdgKh9BpwjTV9qql3ZhFxMy75pFwb
N0ycz4Uv994qCbsGvV0sziiTqzqZa0xe4kSSjZbPVU/wJOqY6ycmxpV6TBVXNeBJ
StFjkbntN4C6017F5oGFPZ4zp7U5zVigoIJL/w3Oedp0yDL/E0TRVNF9hC2kXlfk
D6g1J4y5bB+mmtKiU9hlh/6Plnt8jxLol/m2CSn70ftZZ3nebdia5VY4UY7mpfja
gJQfYt+18OTAb8y4yxBfG1DtvArbMSd2iQSW165QO7no/btGq1bhz7QZ5M5RuvI5
5Fkx5/grkC+s5PvyNH6vUKVDysy3FVmiB+L+hGctcziR+B15UYftph9YM/tfdggg
QkeG2TIlvluXM8JBgNXbqoHydDDlQVYcv4zQrT3eRRRsSulPXb2CZ/c96R5oxJ/z
iBCKWod4NEQbnUzFsmv4xIlI9RNZOQEDk11F4nNZW5ja5PiZ9Bhd3UNTj0LOrUhr
T/RpBY+wNEnziN6pjxH2Jb7jpwmH4DxVyqQoXU/fWENHR3G/NSHzcG1pDAb2W6c/
tvpcsI95CtQnw6/J6cctJWQGPX7gJJTBdMkUGmi8RggQ+G/3FxBQ9YY5KAPiTtf0
mtcr2C37VmTxUDaM4ZxZmBmJSbGd7ovc0+egf68Ybof0o++XycbQQ1Pl9x/DMOf2
RvWKgpXM5S7v4sR1SUpSDlgT8Dsnp2xeSAFbZfpCb1mLM4CLocT2zsCjvXbijHdP
h3hcO9hYTNcgEh6+UJfHLKn0GyUow0IVmmXTT0EV6IYIOoiQKeSiXOR3KewVKrSl
Dcyqcl3S4tZyHUnuoyUizXp/Xd7wRWnKww0WhlGbzVHsO554wbIungOwJs/BxDdT
IOEXC5stwy6DWQQiS8Q4xT1gTx7R7Guql6qoeKEIWmwF/n6Is9kUNydB9iT4EmEo
Knrsp6l9ZIAB7KBG1mxFdZL//XIvUiceDjSTuPqc/YUSWOcovFtDxkJcq2QfsnLW
5LxbD5/4BFBnkNbrsFbExiEFqDWJJR2uUc4x/Q4FdHr+j3SDwMdSKJaoVdMN3cKo
LGmruBNwl5VSS4Ezj/9kge3kS0WsrLIe77cO9niw//gyOxQSRD7dGsq/Avde5J0I
Ejv+2Ub4ieUOhYCZ6xzuVbBi09mWmof/4PFicXezvJh7vBs/ALmWNewtKrKSV1z2
4RgfettWlfQpsxdQNvAuJ9v8l7kfgK8RFLUnC+LiyGOx/5zXKq5p1dMtrg4ONZPU
+sV9Htnb+ZtS9xPK/2tY+HPa9mla+xlgUc8E9IoII8dVmOouMdwlVWc/+GfOUrL9
GsMG6jDFUazaXKujkVa68WDvD9wRf+TsNfyKFQbr0Lp6uXfMj/AZfEuRBMscYWpa
hulyo7EoNqlxkLYTx+9+coBBp/6hiZOOhXGClh/8ZS89/CZkwH689Uju8pZ5J1v/
ka/cnDgIdrEW9ha1qryOrK0MpnflalWZSwiewLnM5T8F3upIgIXsFlLFjBtkC+Ds
snPEAghrbwvpND/yLh+xpDb2pm7RHZZRevME5pqrkxZEyek8jrskhHWUT9k2oEXD
kQ7ZUprf+jy+fz16tJg+SMA6WluTO5/obSl5IibkUZBH1kaRynk1CPRmEYz0fS1p
Cy5wP7XcunjI9HhPYrZngqCQEUotGv8gtgQudtfYokTBXOvq6oEv/KHDemZEbpEu
FqywXBoHmrau03J30NvG9zB5XhwqHf24aMrqfgwYzlND4QrWGTwvsh8jy9THqNsu
NRCa4DaIWp8qET7wh/NCk9zDVqj2Rma1kSleotW2dnw01LtYRcqy68LkLvkz6ee7
YaruaV8hsh93ngHzzNlTQ79c20VI18AcIGKkpB1RD80K5Y1szZ18gANJ2GvseYwr
BSi1URK9UGhllveBd0V4X5lAP2wvoENryx1RbTWW0UhgNgi201Z+hkFl1kGFTOU/
e2iTRFp7Cff1XRuFO7DBmrFSToJ3zdR130mE4SCTSvpm52ap6IxDdux9RSZu4vye
GJ8eN4k/KCiWDVVK/Od+3wC4n8bHLiDswTfJpxAbOn/hMzx9CYO5BQr++HKTYpZK
CP2VNMZn5aCSN7BY74tH/obw8n+y6Twwwepyj2HegXxEIghQfoweRIfglcY2Fl5m
Tpv4m9GWc8UJuNzcrvjKWLhp8aVlMeQf5jaFrF6nef+/TDMeYist5p3Wsk2tEfco
LeXBEUuS3ql4s1OdSmRV/9LTZ3c45gYgUTOc/Ry7JZ6jkGeKgYFoZMH9xAnl0jlL
eIar5IcryHLMQ9sZge1g596YTa4ndtWlS4DXIPL2rcSZdQqdXWoxQBYplB41CV0b
dDkPrtPpOQxzOwq+DFCdTZiIb2t0lpsl8gtZAgTt5axz0WWHMQrIYuJxuzB6FsMW
q3YhuBuxS/IvFLOFeSB7OI4p9PyEmd7/QYQGl1eiL4EmKrkGG+xI7KKQhe2v7yjL
bu8L92cSe67/hJuMjuF+r1B1MmA7h3ekwkhQ4Rfv1DkJhO3ADepAHXpUme7IpRJ9
XY2nfGhK0mYpOmZ0P/UIBjo9m93tVkqFF9TwtSVjIsn7jfAVRhXJFfPphp7CSMPr
mRglNdl4tSKixW2yZhXB4IQAwfonos4ma0uqaxNPxX54nw0VxS/hMSSevHJYVaE8
2jKs9CDC4lljpPu5eRq3VL9GKD+hbrhpcXX95mOC5myze5fnb4PZMTJbFKzGNaxT
RRkEym6nR1S1EobekWbBh9yLvv/2hBdsGY7VpXKugj1MFh50atk6MO51aTePvgRM
Ifbm26jmTfBYzYLh/yiRTHO/+uw6gUAkS0n1P6kgQYQmgVNvoJsRZl7wYqKlTRHh
D6nVPNKd2BY5vUhqklpL+jUmgMyNffxuAnEzkv8Ht5kJUhU5rQ3KPp3E0I3giRa5
qn13WmYc8xKTSVug5+r0jBxBMe2El7C7YMb7DSZbLnI48h8HF2K19tDTdEmZbZH+
0ZEovFd0CVnQVKBIsXBNey8G+cEHOJBRgEOEDVO2NL33X1+ri8ysjyMT6LwKifAd
UC9Fnz4WLFq6zqkgVk+R3okqqWZLAZCJntT2lvSdc5F9hBD4+OLGu74FHwbkny/f
yHYxkqJFP5r8LHVNOK11UfvYkt8esoCtEr2sCT2jTlmoa5FvMD25unn7hvArKjWl
YPKOHnvq/Nm1fN98K34pni1nUuqhjIenBnaH9pvrY8I7IVO6yWxCnN081GIlIdhO
X3ZAc/HoiA9gSytiUX7Pec4dq2V6+ivzIJUmzdX4rXjJj68UHT6hkf6UV8W8N5Zo
vwyi/a+GmLg9pBlXsy3unEwJ1OA6D9kSGSiNzrgiWPekyEfP7A3YLsD+9JfTtMwX
0aHjH6E/xMLzzg8hBraDdd2Zfn0tzBtz+YKuVy52PAf13PpRSrXpPuTv1ubP4UPS
NqzYNmbXSswr7hv/dscREVmhXcN0BFXZVmJgT0KNwhqP7YtDTfE2mWeylasMBpMm
Wb0kzzU3G4Euxu8q/8Lj4j9LC6vTripHlbYtiuQ7OaJVz9JU9zgyrRc4gQgkdVnF
mZTcp6pfG73y8kQVLoMfG4s3t++vjlNnmhFr+JYhtPZCxkZBA6Zna/On/GQfhu6/
AEvFmtbteNjd/vrAMdtpT4A+afRhXMMljLsceBHfQttsRAOnicL20olIZ8JNhYML
S3j9JHatvoSB9sbdwhf0mb7/HXqYaYE/gzBl+oVHmkHUaNP9KkoWPS/CwofPMZfG
wPfoFyFdy8XaCIrLtOa2r+aHg5AaOKeGBq0NL9o/JGTlECXJ6vQ17p6UfyRNiVZU
ATIoz61Ht/GfyOFVlmBx+jz0TGpLx3xEMQaR3GvEdBSmIUqPs6uizwgvBnj/5jwp
hKSlCOi8E5ktH7QjUN5hq7u5gWLUkQj2lZ6xfWE4Di/4RlBz+hXxUraTi5ss1H2Q
I/GyQZp507VpFOvV0+/J5AmZMgMZDKoCggtnd2nqYKftdh6PtogpetA3YOY47Fvl
KFee18CEeWE6NZANzY6PVIm/xr74KyUVEysNvJmOswCIYTAMk1+qoNGmPDjXajP2
XuXZYy6GDc/K+4+jEFekJJirRcE7t5ExMno/5sqJy0OCCYyquJgr8rOj69Mf3uF7
ELBBNjld7cJa2ag2X2Xlwb6bWHO1ZoeJVVo28RoTaIf1rZOGcLxBpkCEBSt5NKGg
v3ICDCyLth5mbcrri5nFvcjlDmissApumI7+HHnY6wVw8evooTz2fSi117czAiU0
6olQJ938g539FlH5ulIabdt9u4GKtde8DOcKA1tXf65sE/moMbdOu92r3gGXXe8x
zmsF6eKT/mRGEejYwuswS1ZY85fUnOehCx76r78aP7jZw/ZN6C9LQFIje7N2akI8
7IovC4MS2oZbkk3jGyM3Rs3m4exFRivUm7W/PcDE9vooTEZtKHwqBOzJY5OMpGp7
domZjgcinMcO1lB75IMo86lE38JNEm1eJ0qYXiZ2c5Xg153fnpxOBXNFk0rKRW3T
q46kx59Ae93Ul1n6VwhFVLj0Q8t6HMEq2whUd/R0WOb49Wv+c+AnfOh/cHS6pQpT
ca9KtKCNZPxO0aXQugymFOl3t9HoT/V3Br90weOkt+bZJH3LU3WNUvZF7UwmNq25
9qXEFMV4eY+soarSWh5XLTq857JfpB3BNmfiQ8k5VVh5C1SL6hSRv9q8xPBjoWhb
AWkkb6/jIEBAchOMuqpbpFolQLsKvibJHj5//X0hW/tVWJ3Zt+uoHwmslWBsrJvt
VQtCOQpohR6L0ApBMSDB+whwkgH0j1kClZDyyNLaEpYOkMDbNTyT8LSIAES9+tWM
Ojrxk6OMTDawOCMCIQeBfThtK8H6RPuIye9gd3n+bmDt7mw5H74mvGu0tTxh/aWj
BIBVzVDMdPfqVSiRsgb++YtHKoVA89YDOI/BVo0TFyV/vu9g3RdObqee85RxysqC
dpE7NAjZM6BmkiNLkOb0Fpryg1fByZgLm+0cDNvZfCEcDb8SpyHEVSrcSe/ldWlA
rHa2c1hFMPAwteSCfhgmgTjzfUHUb7p4ck++GGM0ux4QTVPh5SGCGXc5mIBVbX5s
Ak9J0OZqRyQx63QCVy8D48rznoUsBpVvWavKsHseRNxCrKQBt4mY4p89omqZoeeE
dHae/0mu97Abg/fzWrJ+eQsg8unxWnhVtFjS0py/93ZCCQ8rf/vPu3h8tATV2I6u
BiuXa2DyZjHv8vB9Szq30rbdQgM38G0UU9gQIyfG1jsHSn3QxVpWZ6oSB1t46pGm
wvWYtmVXL/L4fOQ/me32RcoCLHWtFN0YrRV/DhsT/fmbK96fUT4rzND09kccMjHO
5XoK5pBXlyjhyfwujodvR5XgUF54OqOmn+Vl53gL56VncjeBFz63Fk7/5Kpk8P8P
ns/8Fnzdpv+Oi2JXBOsZjBdqgZ9SB5dJF+MhhxepoenKmWo5rpWXTZYkEJQWAGRg
SKUgRRE8s9osuMMW8tvN83wXwR+bf8D5l8z7+32SPS0WqFMJnLTNdk35IohJuvL4
tR09cwezc7qsZX/oHcoiJVYsCAPDbrTblmxRHliAxeLhkgWzxrCkgEIPQAUoBFVH
FYhC/zgmkw9daYPkFmvWuw+c68G+jWMGkJWAXwQopy2hXPApaBGxhebL4mK5ExnX
V6CyM8KRnw0/mtOmREyAyXDxyHzpUQMFKtFaQApDBSoZusrtGk3oDRyJYRa/zn9n
qG1WfDzncVYLIR58vpG8PCaVbE971nEEPhRKqZ/Wlcsgd4acJLMywMacGyDyQYUL
Z8fLhOxR2qNQ8qxB8H/pJMXd360oEkrVEJGNvpZtBUtwHHba/H6OugDuXva4odhL
RszEk/oYnryRYwqfcDD3aZZs9Y2DNajqwiI99IiooieN0Bs6BOCIdsh4eJf9fwIA
Y2hfQJiD9ON13Dg2b94mOJ/zwUS6lTW3MeUr0NgipFt6HU5KyXJA9yDktwYRmPpC
qC6R9TpItnXgrRMLS0YfcM2k6IAHf+DwkCwitwze/Wp7J0uk3LBnHIcwNUX/IKf1
VeRYjbG4VMWhslDx2qrYDcCaAgekPkXiJjwrepShvwYvBnatyH7t6dezRDQYYqcO
XgtPsZAPR/Z/o4ekjfcN4JhYEqHY17Yr9F8PayfNs5KGy77RInklLBxALwcIQNKn
F1Pwxc0yD7WSvkz5SXuFc8h3s8x5gmGgvtaJ7Wqhp0H79QbY9i2Pji2vPCnmQQDO
usnKXH4OnUORiWRtmEpQL+2b9rKWA3OWMPYdnB+lFWAvlr3k5hGqXHkLFiyQVm6B
ElZdXKRnx6lUl0SWkc1mbPra6/AgifJ73D0QCbCjQPgpAFLyxs+YIVYviGYrgQDU
PY1+ezUgEKu2MLPyLj/7Z4oDQl8j93qbA4PyqCqkLnrbmizR0T3PhCdu308HOSfx
ZGPe9VXazN5ui2lOTLc03BS7qfe6cc+D/cqgD5FsMdedE/R/zgSDAoqH6lsd/TvD
5U5dWT57IH7aXjJQ7utHxJ8JcDB7bEXxOfqW1gzLNnZE6SmAkTVLXhYm/NpQu1j7
P1lY0i/rOud77DUN9ajh9sL5z2bmngPueRmHDscNvfcnOOu3mI3Q0PR6ZzyNrgea
YCm8h+WgsMQe1qz/lVvFZFTvdeb3EtLUY2jQsBI7TTvyIJSxStHEM4UWS9IabdT6
ESc5FctAOh2IFZOeT0Nan10f2rMnKz2ukL81llMxKWMHLoEi1hMKGMxry8cOAV09
P6/Td9vRWHuUoiUabJTfQiPLUxQWIJ2klScg444XM7bNvTJxcgwfFlZKMEXbMAtV
U23lIFnvDrGxVMOttx60cZpJBJmbAHQvrlnDneRjKzG7+B/RQJshQwWbTFY+z0X0
cx2O02Rns5QqwB85NmxzTObnZ3s9bmwgy2hnP695kWUQ28RYxRD1EsQjfawSlj0Z
GP4zSYM+gz4yOUAqIABJlDtXKysgxlM1mUHWj+cVJLdLlJ15logUFMHC63iegBLp
noLmkVGKXaMJlJgmEwaiDh54l3w1cHWxPpxuSIbHilbZtQGi4TVx8PXItER7dRNn
vK01QBZ2Gtgf0pkIiOzOiKX76tE6uS02XLY4rWNvnnSBtaVyFm4i95BxHSRAFODF
5jwBT9vSLoa87OmW8uYfq6rzJ40PIUWEt0HwCMSOlse/tLvL6z6XBIecPUue2iZr
9ZY2sCyH8YFdK/Iv7Q+q637tBvzOyQzklrcQHGe9+Z6A7myiVJIbvtAcJZa60sxC
DX554qmODkfdd9HxBVczKtdejVcYs5nC4nuyp13Sri1EMzEd79LVDV4+lWr26keb
Wn1U601DvIAl7ToXClGzPZzSKQYxW6fp07ztLa029M8VupyjoLpghv/1MMIYVoD2
yP1ofD6TBmsvmegl0yamPlziCm3GuKmW+3rAUpYtXTkc60T3n7yvzugZ3v6fmYZ6
zZKK3NyE0uufvOw8fWbL8LwtK2eZtYzVnL3UElnDsVg7H+UU2iiocgxTKUxuY74c
NR50Ro6+yAmML5pO9cC3RQSGzplTTaany4cNLwnmBc2gUTwKTJfjfxoVvuEUq+bc
iqWFgf9x+s5SbQfSjMs0qNNzi/qfBSN86uBmuekvtHPB37wKOj+rbUquVmOtQMLJ
IE70lzPJ7mEzZ/ARW2lOs/Lhh0srUDPYhvSb67Efk6XciUhjTjmYT6/E/uAF82ys
mmi2aDbUVt0ocuXXAkc8rmfOi68oPOf+JKFJgu2Zm66GvQFXb/YcGTBpfrkIwzta
caw4AKTBbSJlgo8Y7ve+SBPAATXwylGsfA/8nsc6bHEH9iFcwWHkovLq9ItWIE+c
ayCjuXxkmI/HOMOxNkr6vFrwhzGetRZpQyN9fyNZzevz/wQ9KbKLcmOhSqjv0+zC
bOHXMQakcRwQJ1FkKZRIaCO/yp9eJh5hZDHgg+Oov4vobY+dGlDjDsyVs9Sd3It/
PxZ7HMkcxWPrP1XtNtdr4JAL5ygTNlY21F/GTHy6MGTbAfLfdsWdWQgEoD1KhXNs
MTP4GY/ejIAeZxkKx/fo/AXACqfZSI24w/PyoYJQ+7ridLBNmQppSKBoLEd7/4v5
VvAJJTN1Ar96ztCwXNlZH7LLyXwBZQiw1BH6jQmYilrVMplzSzaU6Cz9e8uAiCJh
TW9QmLdC3ZVNHxdojMMfjjvRm/KFM62XU89TBrAzlni/J0AM5r0LkAzBU2gIR7Ds
xrw0pnToO/lksEFrbQ/lBXfJnmswjGAGLyMGXLEFVFjRYbQv0VrsQfDkkcVqOYRp
eJwLK/4Cxmd+NL2s+5fRLBbLT9rrOuKlfDHSemv2Rb83oYvUf8DF3Z0h4eiOuaX9
2bwX1/vUrWjqUjiV3PGAzUSiWidwa4MQ5cFksNE7gIpuS5EZyokVWAY2mURBmeGi
mJRHQdgMjx+pV1qLp9XNb1+5IbMb3vGpl3YjcNjtzicBSpf4W9EyUGnXunwA/cJ/
qbrRQbVH6/dC/VksvTAOwnaZxzw+hB8BwVy1y2AVtZf+xdre+AkoMCKenPfcJ8f1
jlRTWy9RWFsdewOcCP4nYUlPw2TVHudc4UhzAkZ0D4NABJsyflPHF1cOO0f6mv4W
zE0ppukD+Cn11LfgMdnZG10AxziTXIrQ/AZHgzt5ogvw2BYLZdQi5ObwPiObE+V6
QRGIvLOnwESsSNd2+NljtyLu4e6HOyl1LtP/pjx+yVqRXDOJQS3tvTfIc5tfiJcC
nz5/5oxXy9AKDx3F/2flBUR+aMH6+CMg84iJqUV66TrZaa1k4DOgp9Zs0WJcFnDV
yt/OUSctqh7cIpcYG2irAnTa6bnwSsoQXgYsXIs3Aw7F3lWqiFuYTacjpkpMR/N4
Dk7lhrjapIuYa8FESC1UyxhdvcAH9/NqWxq44eWNiwIOkCuCmhseMOctmSqKtO1X
S/oBHy2fH8UrXfwqd6i3tTrhMjP6Sf+Xefj07+LNtmoPjWtBiicsDq3nlMrhZkVt
QZ6HMpkfp9VnICiRgMH/ODLFUxTzypm0RGg4ip1s1Yp1Po/L7wxat2FqgegBPAwK
bZRaoChdqUPeXMl6347Mt6jR0nIzAr6E6uAcrua4FfAuT6gdm4nejyqI8GsrGxwd
KdiZ3y2BXtljTikEHVEMcB8X7YGeB1ghbSXbv778SkHaDh62dLFp6UwLruJ7C2oI
qO1rMsJBVv4H9xCvbXlTRCMox9h2qVHX9oVfv0sA2xyEaeTr0lDJGkPTIOIuNgcz
wNxMZ6+7l7MVjbPMS+cjutX0SM3L9lukkxHkbYJw0FYUJzbI0tzz1LcIS1zVDBFQ
vevPO7rYWgikPTQ+Hc5BlfXGIRtslYFF7TIiJ5XIdNkcZNNo2rMlXAFjCuBlG5Rg
/NZNxUh9xfT8PwVH8/tfF2i5gj8xQuyiM5JsPXmXZ5JMRIiyj3ymZl7PPYb1ryjY
hvxwppYAx9P3pbr0WKZmdmdAblRWg691TMX6QwaObdSar5V2BPB4BjC67PHa0WvY
4iyeZ5sQS7wBV/158OQ+9Z+415QTHLu7pRAr0Gh3CQ0lSdWSlG83Sb+7fBvJLCge
jv4SO54Lt6J80d9ZTwMe/3H9qQt5MyG0j8Mp1NdEThYsxgdjjSFY6cNkT+3k3Tmo
wU+if1pt8egZgVBFm6ohGfXC2zR5NGEZDC+4agase2KBv9TFstT/E6Zg5bjT3++p
ALWbSeFzmXSbqot1Md1kMlK5OvKphlBvVKHN11642OsH4DRQ+FiIxDnfF5Dsyr5v
czQjfMQZjghlTl0LgLljkavUoRekkfcgFjhYxFX4ucJIQD9VdwsW0NkxlA5XUU3A
F0SHAD0ddIlzqLSGEIdY2WXBuDL7vE7inDqSjkpmcTgOyiObnDzc6qh3kHjr0R3/
KpoFwHeiU1AhrTVZa7DZ/T51Z4HwrUmi8y6sWVb21exlhXwyd0ymJOk6+dEoY5uw
CaAJoApGEbzOezSKLK/f+EDZtt6J1GQ/adl0NlyjBKMG6r22QLsnZAC8sA2X99JD
+jVRa6kmPfOmUtyxc5fN7dhXxSm6zyEc/j9Q+KGmjZh6EizZSJipHMJeiQTjAatJ
kpzPW3EsgvDs5WGjZ+0PjZE5DaBMOCj64woT/U3QIRemqrKTA+paPPyFIJrn2o27
Segn2ZCmMR8kI6XYVii+L2ENFaagsOEA5S1AFUw3PfOFE1Lwq3EURv1ht380tQVt
BsVhJLNLbjefVMsMseSFQqUPyPY00kkaEPe9yv/F/fS8fqqSXi6Lu8060IrDljGV
AUNMXg/nrQ6T9dYj4bjoDp/rL0hvHe5mQOxJo0t31p7ZhE16DFdGPjR1LWW2dzLD
/OmuAL9vOM/SwhONpE1/Cc2WYUBBU9W3m3oX6q2pnqmQVlJfPP8Mu6zU52WStiQC
TS+SAZGRd1eryHOl+4DiJDkAx0nMKjoJMEHq6A9pxhxjGk+JzcYfgnOhpBEuR25Q
bClXhgjKqVhUr+ci9vFDfGYnmJW2EOhXGtETv7YsknRhry+xTwh03ZYoC17CWir/
QowPWSJUhOPXSK9wMONtbG8nWpsIOmJIswPIRMj2q6t9RYt6kKbp1ESdf28WelUm
/mP+5D77z6dHwpdsd2IhLPOICvLzd0NUSEibAGSHN5trSaL4gHbHRIY7eWlVbgxM
o+Buy3WzFApToKo4cxbm/6zwsmAHPd7DrRp89PbUdE2rbTntmSxjiLeDwWEeVYKb
hO0/3YlwKw1nZLKx4lawvaBWCWph7wMYtRlEmbSLk8HCAf0Hps8ZM5f2Rig6nqHV
3bjQhqErxy8eRC3uJSnDYOLypSKo4Mofp0h3eKPRn7mY6KG7JPdbAIbeEYJ9bKAD
L740L5jLFZqmWwxkxiMUq6eoO4amjf+hrZz8E0F83gGw/jhAXfOSNEISXeGPVjoe
ouLhN2chG9IPgjKGqE0fYTqIa3eBaD4iwcOOLdcgBS/ahGo/IlNfTWRNoEogHow6
fMqk28eHsWLQ9m/X3SDQa75KICwXSGCquzhoAGhCZmMSA+mbiojT2rXSDgW4R5qF
ROsKyJvsjidHXG+ULesMS27VvthgfhnsyHWQfAwTeoEI+6hwDxzcGxsL6ITy+kPC
YynqTeYGAXrrs2HkVl/qQ/D4yvYSyvvAidxNL3Lr6qD/4BqiZ3aMie5zWv79U01B
jQvdq7Y6XGDhGCimqhsrYlLKJ/F5kIvmtcEa6ArM8bYSp8Fz8e7SVmAt/Dekff/7
83zEyUlis3wJKCz4WX7guGv6wWxywptIt6mUm60CngPWEye1SYgFWLqDYpeMBBrl
Owc1Qqzl9JFyrNtAckaUyDrQfeNIRHglg0sNR4n8rwDcAyvew0YSw9ZCSPvVgMdP
absj39LOV0Q7R0eJpOCAFGug95Lfxct8bBX8oZvs0Ux8LIJo5Jjzq4a9ljuzFhYe
qpkfREw4RFKRgOaJZcJV6WlV7BN+GubNFX2fAbuNDC+ivo3F+xOP7Uk4If5+TsUM
Msy18w2Ft3PSxaRxps6zVNkfF+vLJXst6njHB1UWcjl9Pa4oDO1Z9bI46QbtaJm3
4Yv2AYBgVG8Urva9AEOr3f5+1qsEygD7QdJ22Q6wsEIxHbcUCVbcH/XzsrSOCQPe
3M/Xoskz2bL4C5Xf2wkq1V+zFnr5Lmccnl98YleUa4elqKQDOkNbsq2I2XZgwjdS
3JBk9HJd8OyZ/84muEi+sluOORSERkeTl4rOqSlt/35klC929lzUzF649W0DIvsU
iPpokPXJQh/By/fKQq40VDBAwqFTAMVatXG/DnYyNat3fA4cqALrKYUqpD7ga+ok
EB/RTM3ICa3I3/sn0D9jB2NvMYWOjg6YJrBMHsn1//Fc0OHTiGYKcyJ8+TP0REU/
78qFzuuhqab0z5dP6t/kp06B0nS+cphiF9hwGHwdEJ+RApmrL9d8ywbaYbbJ3/5H
Clr6aeubVRTSFf9jjWlgwFWaotPdK7NO27vyvxMOVdCyJB26clFK0aHsIb/ElbqL
uLghziEoDhTJAb6Juy8EE6LJDPRB0FU9/6WEIvH7Y/cS5n0Z0JaakBM/CM1RwHo4
zmATv28UxM7yqAVa50U6mX/49GXDH1l4oL8n7zsDhr3B0cWmvmHd9wAeMmzD+Hqm
KWXMro3P5So1bTikHh98dxgE7PzxJITsBJl4ySD1Br6k9GX3C9yX0PjlDXguiQnL
uArz57bhckG3AbH3F7YsimWpxQvEJnzFRk/o5pworXwmdRfwfRmQ1ZwnqMJDqd9F
aIwDfDyuJkKVI9EnGjelPJLtywWCNkj/sobNMlmXGLSHUr1n3mL5Dx0vuEDiPjck
l+V4fsT3XfaOHTvv6CccdOYuvf1qeE2OpqOuPwl7dMseZkMet2qsBhwBebXJSC9t
UUEt7WM0evPX7dE06E3yej7bXBd6bnmiBVgaOzxU4DhK/6D4eCx+7j3jVcaMjt6e
SkNx56ddwpnW4HZb1MCwln44h5N2OpcqGWARuC41PerXqIUOEXxbZ7A3a2ClQJ7C
sQq9qaxOgRHb8wXW8G2Mb0dxGkGMxMmVSPmqm6WayuRw+tLFnYgkp3AkTcZc9mxT
l5x9S2vYsMKVTb29lmhHb+R1ZS0F0mDGW+SoYTHBya/z9/lwPxhgEhrudoh7hm2s
CmkVlYXwegd+rHHws1yeVv9aPufpWmdtrAmErmbsY4fhlQ3WCJXqQImIBd+bYAdh
BhFFzS+yDQAnAzcyjoh8swQ1uaiwRakR5WJJThiMhyAyfo/jboWiCcXw+tS+CbRu
4W1BdWX2ANmzSih5Yb9LGlEFTtlfNDslMeLVtjjy6OKoi26TUZFq3+BCN1+dTmBI
2buqAb+5wB0lABgnTcdfSOTP8c0GOui7rzn2fQOzfFe/42A/KBz9Ock8VPMPSKln
/aknSc4tuIJDD/QdlGlcNSxQcVG/Xy5ktmkfCqsKdT8l1JcD2VBfL1C2Qg/rhHFg
zWDw0g7bWO6UnF4rUX7wqd0U3qojtg7/zQGX1rGfr5K/cJ4mjWZQDx42Uk5W9Q/e
gY8mD4+gn60xdJrtIP4E3SfhXykkox0eVEwBpXMR6SFS0OeTNfgE9JgNV5bPrLPW
YmISbS+unmZtAsGR6gv4PHitAZDftR3Vp8485x8hHWASOcXO6An3NcMR17Pb6pxI
wTgQWUV4M3w+y1eIlB5ABZjBWSfzNZ1FzhtUByFP2FTWENJGRxjenQFOYmxwxtBq
JOFiilOL4KF1JaTdtgiOmdzcdcDJVTYHgPDGGWYeynelQbOt+/NfmXh9FRGrEsrE
iEF6pcZaZ4f/HkTnk/AAevvsg634Is7Soq7LkXQuEDeTMHlG8oGLTOaFNWjbD2Xd
ncHp16kPgBu4wKiXxywqcXqIl+bEdiQi3PmmMSfEKb5B3VBK658Yi5EuwI9yUwlF
B9mPJtrVWipZWUC4qTMDM628bYsRZns1KRMzLFabe76tm4QuOWp0MmsQCimYo0Ln
qzLrMkMH6GP+uRtGgSMVF6WsJE96jh5H36LMD0hqSyZfJe/U9t5X741MJey6drET
8LXcaceeks7cfCN03trFnJNXddcafmB7b5gNDjbaoMFT8N5+ha1EsM4Q6jNyKKpf
RJNN5ixjlJ9Rs/zNYs4Z1972QCTjTkmAlibwj74G6FsrQMcWR5pbljtGBoAKhKsI
nNZyU+rlVl35OBil2IC82+IgAG0HoSq81X3/67nx5V1s3oM02NFL2WhwSLlM3LT1
GQa+tdrBaT3KptsE88iGlscbnOJ+CPl4ytoyg8Xtr2pJ1SnYQ101ZNm0Kck43xAE
GW1/b7z10MgQFdiDl8jqiEQ8fdthtwuRyi8+ElpsiOTbKdITe/91CVxcJ/Ugd6i2
Ene8QfjYM9L5qljZo0MjGeiyYdC2yP49FLYbEtq0KfRKi+bmsmHDUaj3RYQzgXM0
w+USIhbGCEVSLecyZ1trWxCDDniq5gLneYaXlLvdqwHEs/0hfbJolQR7Usze2vBY
gseWLTfW11VislwkZMYFRzHiaMlsyxUM8NvS4k/TqIh7by7wDzOppkAbWv8uy6Dk
mvF9xY0faGDJRKMhDper4YMjm5VxR5AfVFYe1udhpTBMwoEMNwhq54Xuq2VZPr8H
LLL+zm54ejHOw3IjY6crd3njHERPWssm7C1OVV5HX6qhe7Cl0A+rMJqpKJz/iZgO
W1eZcgOJ2d/bk1wkXkPaftZAdG579ckkX0uFj2EL6LwjUwTClQCV/HOCPsHMw7aL
dxDVusD+cpgxO5BMgmR3k7yed1szHnFmW+cHP4JlT5TF4f82wjrwJNPD2SjwbPiV
60+K5u8S23gay+8O6pXPWyVBArWKp7ygGQQmXBzn07YFdL+xMApumLEZsz+PUgvR
Vc+Le6Subf9TGMNVK77NUsvD5Iktu3z9xGr7Ka6sFjF545Ksa+A9qB0Op8sUJ/h1
gWRhfU8y3PwjuyacSDogCMVz27GJN0YXg6TJy6mhVP5s3glYyjW/aWOJwRpLx8gg
ZVt7h13qsbQZVl4JBKDFSg+4kH5w4ksuEjvDHBGl+IEF5YTOcZDpzzle0Aib2NVg
/F+GYPjxkYnY6W02JqTeeRkWlnqTSBoIbQpvsTH88aDkT8tOAwz0PvbDwMtE7GQA
1dLwcMpIuWjyno0fwlt5v7jy0pzOI9WRupmDDdKLrSarV5VDUzaTP8pfHh7uZctZ
yF5q/xMGaMjI1kSnmWiFsbaeCCZbnFhzTZ9zW/HWKcGffoAjis/C7QC+nmzwEjVq
wQvSeyqZif7ghukpdDJ0TIDr26SKcvu2PCheKXfH7F89qdr6iFXI7nwXL1QTSjjQ
WlKksQ1VBJKGqxlGFQLx58yBWitUKjnsu3Uvr8eeGeHb9s0yRWFZCnqV+skfL3jQ
TqU1fuhx9QKRQaM9qeg88YlBpza7PkKnSZZERmHqXtQtnvaGWorNn2o7vSdXY2O4
sCNPh4htjT1M+eaQtn2w/g5yRxo/S6YQIPLXRdinEJMTCudji7yKoxjsMBykD9Ft
qU+ZuHavA/pNedlfxkMAcPPZL4NsmPMdvAaSS6bvvEUXYcEUBt6Ld99hP4FHCJSi
ToLTnfZBbfGQ20RphKyfZUv/3m1XgqI9gaHAV+/hHo8U+X2o8zybm+ugikiBKOM7
cH+U62wGjvXSFiMfhoJPRr2pFB4nBI2ODDVT6QUzze6hv5clakQnGtAxdBuPXBUW
oZTkrXDiGaMoxmG2DB6A9wjLBvAM307ZP4sIlOthgwJ19NkyBlFKZ4QsUcyb5YiF
0BjwE/bLai5Q8fkbva0fBprHyjEN37gV5ClOFRmwzcjMZ5soPPYahgHrs0S5f1IK
f5NEmqgyzgGfSfs3X8UOwrXb6yINpV9kQLijrpUCCTb2t/xZUxqDnpCnfV2pKMwo
juMzO6TpOUjRfKmvSBVLnxYHTFqWLc+GRxjUhsiR10FdyXDfyAKlDHDAqkayMTYD
onACjqJdHIPZoUoXppe8jrhSXHoF3GX1cvdNHdk9riZA4TW0iDU09kyBkZl/Zfvg
r+3LlOz154NAmuNWhIgDS4mWtkINljVh07DDPyYnIbXZ58bgipUozSdzfZfxyyeQ
1zpwNLP08+NuZgobrnJAdfi7+Fn3SRmGMEZ7DGlm0JP1WOHGftQLx1FC2ew/78jx
/NzFVWklxZslTgoeAtfpK77m6SfdMRqWp8JB6FE74d1QNeKWQoJvsXSvU5bfv+hv
0Q0vmkf1YviE08lLrVmCgl758Xt0ewEphjS/6Hh15bGz5gtzITZ5Q+yTE3/+N9AT
7yXak+dhUgI+dtHX730ebIgTOXH8UKRn5zufErx95szntyJfKaC1sPZ1geV/vdXe
ajvpK/Us0DJezo/mgiUQ3iy8Ys9zsIweui2o+/joJ0IiIHHLbdU8JmHz5tkD9TFz
CVM3FtcOVlHQHX9jJyBqHCb8iGZTEllx908s34ek00LSmIZjUcaNVQKJhUbfxtl8
jrJ4bnNO0+5atUNY97oNmt8EEnkSSLB4qGzlyub5tH2I12mMfWo+CDs8UGGTpyHw
SJ3flFNmcW+5WexmmkTjUbApOmEvXWBxgoLv47YAz9UHXHHKnGEdhyI88I2V2QN2
kGzMkBFhzdG3kseV8GUPA/dO796Bh4a79x30Gk0dMUrR3EPnTlX4Snl8ryBf7iyD
pdLtXT+r5R6lnrRFgAcTGbg96Rg8IuTAYVA6SSvF6quESkUxOkfzrAmNwSIjigsv
JAqXKPDp0K1RNk+7zX7BF8/6nuWrMxzigHfp+mDCFPHuGcTwZvEoO8OYC3eDQ88b
iJ/h56JlA9zD500yqJyucJV/x+umYJ8LY2VKIA74u9iqFpgddKJxEi7B/ZP8tVyc
5cpYyMIAkT5Ic/MO2kVOgf818Uofg1ksdLnVhahgWmPINKdtzuHKnsx/z7h93HfO
vyPl2NU4NCj/WzlzMQdDGlQ8tWj+2TUhR/k+mUjqKAU9ifMRd9WqpaYF8kv4xzV6
ywMOHMTCQ9jGAyMy0lOLVjq8kQQEO8KmwDfh1pBx4dAFlJXTxtozPqNz2wSMiJaT
L4El4ZxyMlY5nZkBhiWuIE0O7dn1QztCjF5jAzLB0xUIa1TRBG12JmmiY/TlZJ/Y
iSKEUf6tY3xeey9rWRYYzTFa/fMg+8TwH2fmFrgMm1LajObfdIcRsSgx12LrBLfo
TjZQygWYTSeGr8KM8XeAwQm2ty2VDPX9pFlwXYaeX0sBFTjT7q5Fk3+v0uqVXFw+
PTpnQfuPZg4AE3uxYRTCEi9xipXxoZ65ExEJGajK4926vxFuHXmKPTznr0KWZTuU
21I+mDEPwqnO228xUZoROC8zVTjg7PfZ4SgQzwh25LLoywCTqVCvEO4Q97JaYpHK
RyxiCZ/tnUhRT36PIt1mArwE7LsQIj+8erNp3EZakv4xKmiPPB1wxhDhyjn8GSmK
Mh+F6RY90smUiPGCubTOv64jJPWqJRH4ER2IZfhnSzXxfj8qwB/mosJO+Da7+FmB
FVkrMDItKjc7bfs6Efr4ETHh99wHV2VKLNxuFBj4grvA9lLZaG3BLd9cy6qW7ejI
KurN18vJSM0k/5kfHHpD88RR7Fv+xRokq3LSIncp/Sc4oo4pFNrFGOcHNhQ0HHIN
DhfPWRh72PuShHfDfO370AGWFNGjaj02ApgWpiOSrvSwA2kdACeFX4ZTma5Gj6cI
675yWLgcWjivYYaES8J/xWbDlivgXPcSL+kLfumhcILcke9g6I+r0m3T3sjIe9RS
U2bVTCynHL4lzDAnvgRvpRWGm0iSBFgU9D8IYfuBKq4yJEhF54Hv2xTV47FIcSPR
+ZfoTyzcaaBROE1uI2B/jXFF1Wk8VKML65omUutdsG1fWFu7dz/sgwy7k6rMygEn
fDQS5jXfYaL2WGGltbvgzoj7BNHL1F0YfPy9uGefkVeEnoLqZxExcwzlPqAvabs3
Gxyw0VBGuMEIxAlI6hagQjY0iQ0PhVQoZJ/RXfDgg9Rl6HvmcRnBnEJkmeDufL+I
9vUgHHHtQiXda8Z0UdNF6j7SPpy16ZlH1640zUp0uhvLJ+bRI2pVzYxfeqEsy3Zh
xFG1vmJLQA4B+BxDZuvsXi9GEtpSYMz1gBNJaL1siOF9RW7cF8jMpC3+vvPQ3ody
0MZaJaCAQX5UrZAkEfZWHOpoTal1NIQon9rK68Xxh0It+FFQ+sM773lmqgOP8rWL
ccHLO+wEGDip+lTdqjZzWdoTo6XRq6aDRal3O9RwxWLTswCN5C3EKhOYr8Tnt5Xy
AAJ3yZGFVchTnqD/NK++zMCyx43W8qbzdwLcX5sehykR3tg+jL0yR3Gs90Vzmr2/
b/BrDNszXrEK2X2gcuTY30BeHM/YhkZGKRIXDJ7AVjIsZeOs5/9f/tNM8gyO+3KV
o0G/KAZEGEi8DbVIgeggI11VZEQ58CE1a5IjFtnZZOPJFS08+WUkV7hlAKWZEL8E
ZBw58IUGBnUhmNJMZ/NBoSDAZbRg70ughEPvxu5dxPKmyhaIHBG6P0TJcDo9VAHx
y8E9gcdfjTeEJZa9YwK7Vqq2efthzkOz0LhMX1DVOhuuGcGWeqLvgEoV5qrCYI6o
4CicGUmNFWL/oDAcWeYxYSFA7oLREtlPlqMkWnd8w/nBYXi/RxQHqowE4C317TtL
LfAU7FkCFieu4nvu70eV0vpK8jaAoZZ7wpqWrhHefgYSIGjC/oigHM6my5z7ub0m
dCkqd+8a2xyQJRw3uMhFEf8vibKvBRmE3ZXwaMUcun7VdymZgyh9DEKp6fccZ2JZ
H934OETuSzYDT8YmUVJGh9lP7vkcahsJx6KkP0qkl9XkOQlXu2IdZg2AbotgjTKp
CeQ28pgJFh+Is5hAdegF0cQX3t1bl5Xz8F0cAPBotBvUAQBN/Pm16AWxq9PV1a7/
ZUVtMJlOkYVNqDl7zxiXXYSlvI+mwBm626Rb1dGOYs+eXjzuLmgvoxKaUaaPJDw3
vYK09DaDaE+MQsXuVW9aYxzbpxDDCfrHuWciNTFtKuwxTmfhJWLhzGwAiH4yd6ec
vO42rs/87z3EkcGhVvKQ+lmCZtSZRneTa3lpb23efbRe4AyaBQf0mJQULbRlbQ4Z
sXdmC2vxCpgq/BptiPN1eABbLU1nxxkDlIkd4txyEIOaExjLkojpNVK7IVDe/8jm
YeNqwStS4lfZuRl5k0HS1SLJ0fxTuhBTXyNUu5TieJmunLbl7tG+QQ09dmvMVqlE
tclnbMQlzTW+tsy7lohRvhIQtHGzd7LGz0evhYb/SuKb//m2MB0wbfGrVl7RxIYo
CzqHQJuqyx9+0ORRyAWYQyeFqQuEl8DLzrscf2zzUKA97L49dEwcSQ/0IU5tJ1dA
m2r+TmWtsnRg2P7mmuGXk4Tcjhvh5+RcSGjiQKf83mVYR9K+4qVXe+3jd8JmMKF/
/4RgUVqE80osPtSBHamcFwaP07SCnERYgG2z6teZre7wkf6lQn49h5On66Af+mFK
AvqyOGnIlo2doc/3yW6jbW+P0h3K/rK4xnyPA/NnG7Rj9yDRQo32EG0rOfqAC1Wj
ruDwK6jW0v3kkxFKW6a8waYyBJYcmLqP8H/rmWlEEdSqiLKRWTMTbj5Jtghf5T82
YQBB2clyPwPbON/sVHNB9GjH5al+aVa5y5UdCYbMaXhSui/TTyatlpa+8HxORpdj
6ZCqdzhxXs7L2iOMgfrXB0Rk2XmttxpYoM6l4OqUh8q/JiU+y/vE7GCMPFEE5/+f
IYmGG5z2GjmDIgq16dmrXq3iYPNIqgmPJ+Or7UsHyJoZGExgwyfcqVYDSm+35O6t
tkA91I+UwE/dBEdDlejBKuFfhxocuHh99c57EsqwC2yHLRQ/BFDwrjfxy/um/IMD
ENFgliRCzArQLF6UmCYgJK/SGRWaol6wUaYKCI9Ru2pjX4Tp4MumZ8VRB32l3MN6
lHZHpwSn6y89t2zTGLBhFE9psP7MKrgvm4ogq02eD4HGu7maalNfGy1DNz1ubKgh
bX48VZdfxc0+vbrnRDbl2UVVxZpjTQOxMs0whOnovk0pTuKARetOhuMLOmmTw7UF
Z4DLp8RvDX49ecYgoPMA4scYk4ShN73qGoUN9b8OZykgYE+U44ce448bJcBy5eHK
cIrf0YB2yWg8xenN42nyqKwLl92xPbzyMcm7/OeNoHtzHy4gTYgCFwvh0BHbIF7+
2Lr+Cy+96udh0dXWlLkIIYWZUULuxX9ML3WyiT0Z8Y7L8kDsqeCyh9tkbR9ae5/n
xYVqunzEi79+FsbLrdNOQBqOAU68+M68/GzMVvQZHTDcXe5KdOW8sjFkeMeVYYGV
JD7RFZg93kOTQuyzucvtYuDmUrrD1SVzwHycOLHU92W03PM9pUR+z80kQK8Gxd7p
2GYMPWqe3nzVW11klw6DZWa/W99/QSy5OuTXKNbIypc4kVLj52+93krPjj3IiJhI
lEcy6UiieE/raNHOceee5CUL5CU5gQdl5KKNW9DWbDEM/TnmHe2s2a02mSDolIfk
rjf6AJSkYP8LSkjGZEK/rf9It8UN14tVNLJDFAqylKGGpgY1DLnV32fnZZqmymgK
F/uF4UcvASST9RCZ1heODK3psXmjAo2fnXBsd41Mx4hd7rGBmnYz3ssJFbVyv+Hm
`protect END_PROTECTED
