`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mf2WucFFzm1OP6Z5KaelWjdIWIvzN9yFcwtwWcMoL7AxqdGPRj5tginyoLDosEsY
Ax6W/hP40/pPpwrMLhy/hyiENnr1UqUbwGU7VZyI4RKmN82GdJAxeoj/jcjZxcYV
4jSVScTGzBeUqoiJcGvjfhoLdtpJmz+UAyEZPT5eUJGGhSQf+L1mg/7xdwEJ317n
3/g0xQ43hUOzNN+4RfSmNlrmpkb7yZxMaPho1/0yq6HLzxYDTE/RPUd7XTLiGQ7O
QhhVMeWN3TyNovntAm1U51FkRJYYCv9A3noz00IgdMYu4Rbl65Fa1wJUWIqvgsj+
GfmhQ8bRqKNpzwd3Yal1G3+JfT6xQmzmjNrHkJ5JEpO90r2tQwomB5+m+zdR8zyv
T+tG4mpjPJYpjyLvMLrcx/Yvm99+nTsCWhR/pFLGfZzsyTkD1UGy7tkG0c8iTNl+
mV/CF/tHu74GjZsQ/WBGJZR7PlIieq14BQZeaf1CMgUvY1ZdrTCqgbqYj5alOQGr
jTkTr99RWxMWK0VmSeIeiQnfcbXRjp/Lhm0sq7b++Bo3f/JKFWJAgVaDC6pTGyk0
OgBpcSyhV1enH3l6ocy6Y508/WsgT07LO8sd3BHWalpw3nUJICCTzHTeHZUHZ2fD
88ubRWhlcD0VXsxHcVWW9nA2MMG4wlOtAtDbY5NVTnJv7zy570WgnVgU3HxAWQrR
Zzivgw70r6f8XRNuMTXXioEThot4FnDfqaL6CrAYQQ6xMfmwqp9v61PsqKpSGcGd
D1yBEMDqDXU8nDjLTX0Mv2YO2iMIEl0Jf5MTrrWnCaAktDbOpYvtI+5J18odyup3
YQLZvtA1EYXlokUIk4e+UV47n611ZJb8j6c3oezF92dWvXub0xQOIBdSUovV7yTj
V+4a9R+m0BZ2xIvcBVNw9k/Xxct19I4FAhN8a8CUo4L8dJklbfKxhtOdtCwswlPS
kSDiu0lY/eiLNLs+EXWngYVo/rVQOmIa9wX5+NR/a78RRsDae5pd9WXezoAepWn2
uy3xsCqNjcWzGdhM+efch9E0eiwc71KJ3WF9vgQVN3mFpA+143Jfq8mBRsiKlRGe
KVZKq2hW1wvaEOsjjoAevUBeNzLbiYSt/rY/1M/TR6WT/DywCF7TCqHRUhEK2f9X
KVMRaj0tIB3wCnwxQAVcEJw7R6CRkZx+TP6V4M3IJcXBVxp+4TbG9MUfrhYNQ82E
8b28Xf+rI/2eP/iEWcdgdhs83CqjeN/azxhj3QhvBy/8IC86rde1P51VA4Bo8JxH
hutCFqVaJ+9s1eL425jcsGAT+hph5+PzaQ2HPcEEhxL0AfXrvbb8MXEUsMQ8lRt8
qBWHpjuLsmkk7n2KDt+G8j+9yulsfc9T5NXrf0gHjsVCfXc5M/QUGfLf8aT8qft0
+wc/kQ8LYeDofP8mq5Zh8ee96gmyMIs7hcme5GoiFnfkKTW+oajMpJlZNhTyUBaF
wPHc0WBzyP8+YNxyF2E7dhFuX/YcT23UrPUrtAFLCb+AxScr5zv/7TythywEzgnU
Mu5jpzIDmUDpJtKFnYo1zGpKStm7xz8pAtWe3Z3FqgxfBSewiFrMVg1QpPLyoxEn
`protect END_PROTECTED
