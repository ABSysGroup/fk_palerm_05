`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XTQCHziYljlMjTgXh9yutkJXoKRQFjnyy17LDmUsDwUd5hELO485QWsAA9DquU9T
YgboEAXCQWlIh8s/++ILgytcWkihb8Uyj3eywWmPttVXz767/BMLfXwArcIC66A6
ZJ1MRFcLrsoHTKjqUSxKh4176AVq/vx58ep6pKVxaRt87frNvgTEgO9wcMumnUmb
hO4afYn8/0RZj/NJ7uoUC3Krw/6Wn24bvLHktCIcoU0vEQSYytBdMgAkWQbStrXE
4Y31Kw9neS2LDEGd78lm+dSaNW1udzL2GJegpVjilf2KgO+FtoNdcUAQc/LoAmma
`protect END_PROTECTED
