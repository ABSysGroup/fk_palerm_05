`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PROXSaNzU7wRgsBgcqt/kLZqVTurZX11+w5FTNxew/zLttyYCOp/sI5m8YL3eyZj
5RtyfvTy19xPO4SZaSDvz8ANDwXq9kHwRNJ2sHcI13OusxWb5+H2iM5/Mv3rF0BM
+jU5GYAooXcFaFKDVM93aYOHKZAsj0RF5eNBluejB8iDmPqxa4G5V7Hv4fvAabec
w68vdHi6d8oGj3KCF3lJH3brg+zSlOjqBSRr+NXlCwxGrTsMApf3h71es7TXPhfy
nbnrvus/EeWAIMsbvq5QjJd2KFqP35I97hd5aRG9XlxA9x1WTKmEj9eEeljPLynv
w07aqOjiCErilHyDuFELVBorhbG3mbQTdo+buMZUItt8h/95yqjGJSneAu8xuxWM
EAc9Nx0JOGGJZc1nvj0IsPlr9qDjtYYodZ6eF9/UJ0GvOMhC0nMzzc4R1Hu5RaNL
GOOD494WXDBYPfLRmz78dO5/kK13xMWDPKxfZPkHaD/4MJXAbgpOEOwjADqKtINn
GjaccAeRAz6nub1lDlufYPHw0WQGFBuOGP1oGO8hrD1q7Mg8xM3JGMTwNuq9uuMb
/r8Qxp0R2VHB862WHgUNbmYPI9RArL+vYc+CMaXkmfk3gfCeA5bJcV0q3s4Zilef
8siFEbauwQbbe/upSDwRBA==
`protect END_PROTECTED
