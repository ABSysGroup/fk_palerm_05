`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VjMOMGl2Qj0fJWW5qksFzfPnyhUMs3/7PfF1NzWXppM88mYxjliamMcOhm2x3Tt6
o2+TPHgvxmd+5my0oa17dGU+Si/WNwq3AbGD0B4bVDCmq0WTf4UdDNNJhpWJRCRc
BqXsopjTIXLJIA2cvjcanLkF6oMbsSWf/21tu9C2nvsEToJxemIcZVkticscYYRG
QtKyHPAD+Qc0AlDD89WXt0O/SQlYx71JKJ06bC8xMGf92oQkSAB2i8qsPw5aM1Bo
z/yrU6sQXZkt+2ayvra9jbOWsc9PsYNlWEuCjEtfOsQ=
`protect END_PROTECTED
