`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LSYmpPGc3vIHVuIZ0vZfW/n80WhD+vshw9f8c3p1jjks2j6RSMtZLF5RIN1zwqiq
r/jVlbJ0vU+pprfbUaFLehCiDGhz7O85rItZ+4XfADFMGvkTawwLFkPalw6Eidu4
auGqxeKwFm3OTPKYPhtJamjNo1WJBlb4JpaB8cx3Mlh9RtEHdRP3xyon5bC89BD9
EzvX+IlLSpByS7+OIp4BDI7/KD+4sv5D8wb69MIabvQDBiRrcvaQyaWcaw7JEwDs
JxPzJXn0nx2sxPT3YojQAt2YmlEX6SQPxl2nz9oBo/gmFhWAk+3EoIS/+q825bKm
tVX0ixy/00yBwNMc4DmBnMxlEmVn0bKTwKDr+obPXwuAk8vg2EOfcXapr55K0ht0
dq3zaQK6ajkZK6tZVweiAp3jvdkXBqVieFOWTvwDBGIoCDOC6BOLg/4A6kAiu2TG
EZy5/YTk83h4bYgvKiJKB5KpB7RB3rdFQEQE+QAZEvcbeav4e33djJ+xbDgCg7I6
mlwlH7cG/M5h+HUaBUI9pvNfadfyFe3b8RVq9Tqh/JCvLbDXZxYspxdB4+aHU1rp
HYys2/jNaV08ZMn1rOgVDjxO27w8rEaMiaA/H5TSEygxALVH8IiuJDi1KxBcRN1c
rPH4j/8qeIN5lub5egJaBBL/zHSreLReKY6yMcv3LgRN2Q4LdaVZR5cEkXXAxy8x
08LpN+uUHBPOSrrW6sUNbmPqWApQc21+WDefZA/cBaUTDimbM/gOVx37hBAYQOER
`protect END_PROTECTED
