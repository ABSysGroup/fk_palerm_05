`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K41RtgOadSh3Tn2KwqQedxOE2Js04ChJB0yo/qW8BOZs0oDNpkJnrfvxXp6iXeyI
eWDYYki7aWfUzlnuU5pIjPlad0pIugizWCQehwzN7YemOP7DBp9Gpu/DnuoQGgXH
AmhR7LbiiFWnNEAelxM86VB+bzzWPUAsEzlmy+fDvPWLrQ5rBWfE4dE0n8e/lGOI
OyXoqV93mED7nhUJMdtvv48+7QAOecfGq61IvXWcJoqJ9lmD25tfexZpG5q8Gk7y
HFM6piGwxVjrlDAC1Sl+ljsInxjQXKRDi7LERAeRTC/tFDDkxnP5XwXptZovYsEl
iLpM9oa0oFO/8rHqka+JryTKpyyXK3kEDqh1TTwkUpC5vKY1Aiz4t3hAkQ7xRbuE
glfud/43542XH/9z61Cm6G5msv04c1uC5kEuFSZ5ZjeciJZyBjRWz4qkUFD/ccRf
wdfY1BX7aBq3MkEAyYcvNdSm3aZQur6vr0jxsakL+Y9RR5cdazhzdsO669VYvR9S
YVphufEVjFvbFtZyhLvgDMwZIru3D7ns40QfY0Wp/5GruSvHrqwX/MHHxC4ywlkG
0B1+nfQSbdKEEToYLrtNUEy3MgPxjrL8EAbeXylLti8outhCsWed0Lver/Xy4hgi
IFuI81Fm8gogGRminEmw0acjHOnbQaSoeXwYLcVmz/f1rnlPRu7ZEgiei3vPWKUa
`protect END_PROTECTED
