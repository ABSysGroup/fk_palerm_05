`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KqjHaGBrvg1peWHq+qnLpmNU0Y/iQumQS7L+CMC4yGaplWs6m0p482vPWQCHBHqK
qABXo27X6nmvNZcqyD481oWF0lxZOYnBK8yPo9ryqFP9W6/j2Q2a1Yw0LotRvWLv
/l9ZgOQD6JBfr8QL5JBrmdnph6WbWTkn4AnLzHieEqxsEWY4zTJRAFu09isyn6jq
+Ec0j6JspthpslKxzxWGJ/vVZlWuwQ1lBmoM8z3+2p2c1+yiLGLo9hhXChD6lA6D
Ndvz+cEIU8PwfLPGkLYkqCbHKxez4TKNHJIBkexHcegWcAAMFxjN1pXEQK4HEhsS
j0qOlbAUqCkkvLq292o3NW+zL1107AVRsopZDrDX29ia8TlQKzSzZ/00zkLcSxTH
LA36QRrCicR8D8tFMbk5C5YasFARdfRv+BJ16Hmyx1ehj2+6w5dMl69hI4NrZKk8
n5k8VoyWGP5LC079h6RYiySFGortViJ4hn2/TimwJuZUXQK6UWLlqO+trwBCwVqt
deozixhgOp/LaeRbgucg6hiRHr2kBbt1odacJY1hFbSqmHgNa2xdQ4dscuxYn7hA
Qy1uq5GezYSRwRFXjx6SlgwzXribrs4v0W/m2DlY9K0IE1C3pZoHK+WBUNLf8Bdw
K+XXMLfgsS8YATlbDV0UE44dp7iaQRHmhVZ/lqInbuZsKw/ebcS8g4g+ijg+P/Px
vMGKimZn07pYpshCdkJSm9IgXEZJGojaReonHOpz9I3sfnBiKJENDknll+ZmpGbg
iLZLQWmYZP+Sc5FAfEYOMfruKoMQUQT61kvZngR8rOuFo2LYS/u69YTHp9o+p9i9
tdwCmPrLf9i1GUxs8JsHEiTBadycikPnkiNNXbELChxcuBr+g7ZO6v231uaZBza0
0oiWFoNUSNxaZeNpUHE/MqRDa9VyO305NZjuH2cvSd4WloeAQLcUybDcN4T2Klja
KFFFW9AXdrugMiNEDdLWhYcnrzw7ZHMgqmunqM9OgUBNRQGblQDu22pxFJmWzW6r
aBJigIq/MirbvF6iQXi9NqyHfhpKW+56uUquWcUgUP45TVkBVp8kaEcvtw7DaMnP
e7MFsCbiPaKagfe2avjFlcqW7RRNdQZwIzh5KHQHVouDvj2q+XOiSyiyurMPpXQD
xGylYoOc4TRF4Kz7W3CdZsoEGAZ1ipQywX+fC7c8nw9PRlGzUi61MOKzSlYknKWY
iOGlW7jIARp5PeUHVgjP5RWMFGwjoY/hZ0SO1+sqSNJCxBbRzc8CfAM3Ky86yqC+
WbF5r32nfSzXMY8NCJPPrnGAvWKBLJjadsmCkZga6yRpYEQ9TDqowARVAhaKuSyv
kUKBhGC+q1WmW3XEcyKcBfjsSIWNs3HogGQ2hC+cvxf7T3JZnRpLQtCW/SvtEnfl
eEnzl/Y4lOV14rfyFPt3zCcEyHKeIV6q6aMWwVpqt7oRIhxB3Wtmct2R+S2Qbgah
2S9C+iBEVCEh3OQEMCLXwcTQzZljNUKWNpPuoGmmfWgwfcpVpYGqzm70c9FJ3CHX
/5CpI/7Pr3xy70WsQ5iZuF4kk9EOx3nNAwBrATd42dfbvfYlUsE+VyjSKhRFJIg4
`protect END_PROTECTED
