`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0E63rqW9ylcyq5UioEOFgITv48l2hmbt/tmCLXYpsAWbt8Fm8xHnI3Gua1UCrbDD
VtuqcYtTsOYcpAcRDlpsVokHBd9dSrFxcRhZ9wr2Fsu4slYeNI1rlAATsCvBMmaU
W6331FJFYAdrh1bc77iZNgIPXHJW78mPJUiv509sq8htO5kkR2vde5/QZmCmWe32
0mIArCnCuQkk66WnL81Z3beevBJoO1x7pUkDko3GsOxXwa66nQq1LPe/L+BFQ7Jz
FooR7DJvwvjhuvT6ZUZA4Tb7SI4u69p0x3LROmQfptXBsneGvZ2uh0fh88fE50JW
UF0tiuKX2xCZ+ATE04DnSfcdsRyM5+M2jd8MWJFswFtGo/+rMMDW9eMRL/+KsGin
`protect END_PROTECTED
