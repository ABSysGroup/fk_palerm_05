`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GjwVQxFGvU04u+LYQLF90f9Bdp+h050UT0TZPU1lwSJsTuRFTMRncTyaOtF425cL
P0f01Ri5bR5+KTXNUzNLx3a9QXch872miHT9J+eZZA31VvJvMaEKgEA8KfQASJKr
xiZrRJslmRYJHEWvVImokNqocT40HxFdKF/B2HcBHEtBEC1nWYR81NY0Ra+12shs
HaaCiQkzshLY4LE7mHIrBVnXEo8MN/7F1owNVg9oveUlC04maZz1fRuIq4a445mJ
Cjp182JbWIO9s07oYz+alFhmWWnH3oZsfcFJQBNxnwX/oE+H/Xqqk+Mo2RNhOeAQ
MZXnCXz/EoPu8SdAuK/2XLx+GIEJHLHUR3S4NwEkt9NrW6Og0EEHsedVb8zQ/83n
s2cHpFjuyBEiyPgxQvf9BJ2sHFc80Y3qfG9ELF4wSsK+Nrwa9Qevuwh1NV7gmPH/
gDCdYvgvkMJwKhXSeMcNVIrQIJEmQr1QSYxdEmNsniCcbPRWLfMtREDyQaezIvnQ
bkuEybqyDGDqba0UzoN/vYK2JqJYhoTtjzqVqRK2yq2nDZgpEwQMbQvKkuBgard9
8XBx1sRO3seeMxVJpxnTCSavUxw42N3F2nM24oB/cNTdFxzBFEOPeHNny98A374Q
wa940VoqLbbzXNp7fncDA6dLMpCPOrLGGwarptidNTZs46CMfikqRDxu7pjF+be7
6wAY4MjvXJORGC3jHT7bKMOPYgNcxhITB2hElG9Sb5u48rWzP0oPGIgbQeJ2A4ra
vFYCAuA9X7tePZM+hdkhJNiGxmpCgIByjDBoocEDoy+qolnm9VZPJ0YoR14wPNkH
NMtaxDorsWYPXVEDJbUuXDkvDUIuuH9JYxrXx5Hd/PM2qwxsjIvtNb8Oz7YH/XmN
yYgY1OtNeLAs+eeMWXtcNl7ZcoDMncYfGFRdtG19ioB5siS+M6JEMyfLjpwcb21+
obB3hfIkqXNYANfrueqHmW0H8qkji2nYKhNhRg5yJFK5g4ucK0P67lqOhCnZ8qEh
ouSBNGRf+lvbFQV+TJSMrPIQbo/K7E/O0e8uID+PLIEo1EYSdoGF55qkHsWMGiq5
qfgvb0tUMI8quPf4nJIBNxgmbXWRlnIAhiYv/aHzIoPMGKCUs64kCYkssdGnp6/s
rDZf2z6lEGIqAXBpjEHUH2D1ebuLThiXf21kDqzOSkjSjFgM2zmsb9MnA/WXwgp5
GGlWsgi/JCpeL5/xkFukUIo7HZzPC4elD6dnpcFNlS4BiiNPb0/64eiOerss3poO
Te9sT+bCIFLjmrqv5y6h2L6HsokDT4YOAnvLuHkKRmkHwwhqDVTN0rMsQXrlsVPm
cnAV5eVcX49p/K2P6OxoBmSEgv9KGfQ5Rhe7wHW4uwKI/RZndi2DEi4QM/avZXZh
3y8vQtWkjllKa8fgL7ZmwaLXijM8LEpwwl9zlFHhBK1TC2xuGpttlhdW9ynxvwXQ
IBtFu5GIaTKtQclG4nehn3w3K4VrPn3vcn4mzzKZBiz4fSqN5JukygPq7W0C7BCm
JqzcfQUZzV+H4enbwFr36Cc5MY3sS5qdCbJ4+IgYXZVCPjDxfQg8Y8RE9gU0UPJ0
vBDydZKsY7pW0t/8wmaKQyjXILN7JEzzGGUchXCcoWJSVLpMG6gNPCoJpmt3K0dt
6YCQol2ghNOyV9X8Tfc5HJAjUSGhZ00+UhB+7msg9wd79O2aNRPi2DurtMO0efgG
0BmeA9DBPYHyW+//MHBjgRV5txBe9ZPMKEuAM2xSMAEkFpwth5hbskciWloWZb9N
esDK5hI1FgX9YvDMK0Yk8wYMbdUvBXaqp9DsN6O2q0GiRQmdXLy13fLSKMXACB/G
qdH4nQjVbx3jd1ep3xI60jCYu3V3wgj5uP8+hLCUAs5Npx3DCoN2j7EgqLfl+if5
amRENQk51F01WanjLsAaKA==
`protect END_PROTECTED
