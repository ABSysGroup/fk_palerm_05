`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ubcoXwiTGRe+1Vk1Ml+o1sdy/9/iEQjGY79nXsZba1rcHE6yy3G4Ihp3W6tri4U
sn12GyNXZgkIWqAn8ydetH9yII3CVYkoNpcwfQqGUc6BA3W+OqDCK41/KGy78c+R
RC1MC7M2aZFuZOAtcA1XtGmgdFQh4KJbgW9mt/M6hNp4R2g8Xm7CnDVmEsTQS3wr
keTAFAjSKos3AO1+L404QU37u03ubdlQ/ZKUJwh1d7na4bP5dXMiVjsMzQeMXTZK
hwUD4cRPppVY8KFmjU1J55gQa9taKBmSmN9ZWScF0OoNW5RAYw6qb+V4D374z5ok
pNu3OEOWWpOpcw36q/eK+A==
`protect END_PROTECTED
