`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z3FJQNBXOiiwxrhcdFjKi69P0WMHOG7sze1kMAr2OchpXG3dgKxk+eDzy9juorm0
CBuV+78RKvC9rUTXJX04Qar2Bv42kX+LdU8cVXjZFVawFndqam/PtbZxTbo9eNl/
j6541uGdQOy/Vp+/F6nD0dt/eVPCsAWPmNcGO1kwJhC+gaPTFfhw9FUZ95lNpD1h
oapSt6tCVTU/tyvvbRuE7Ffg13Z6H+s8CZcZyEQRqLPLGKWtaiv0sn3EjVH3zh2Z
HyEkvtS0YiTOEDJLVdQaddC5ehIaTxeRnhzM8SVqE5hfaWft3ImoKKqrWz5/a6qT
esktN4H2+KJgG+C5GUdC6dzKPwleeXiVCmtUyoksLik3DTylmus2dj2j5kQwnjKk
h09NjT9PDrUTMD8ISpQD36t9IZ2TBG1MfdGr7qmUdVPWAhjFTu/j7p/GvRg3yUYT
tT6RvlMScoplTXMu2Z1eNeyOt3qhBOq4MD7P/6BNG2CpRK7CQatH0NL+Skz8ng+L
JlwTA15MZoGUu0DF/C3X2WmOCopNkZUuR34lAkap6szI592bQpB8erb28GH277ob
ueswIWecngoCOaprdpdqQyrqoncOAXMeSAGqtO30dnQfyzPrH+wOAV8845zQzbzv
s9d1hb46AJ5JaRKKTutRmqbT8vBnBZr/cF4YrgkwrN19rym2EUZ7HAXo9VYU/uPL
KgLNTI2QUrMOL8Xs41FUk9/z9mVTvbVUPItgqX2dmuLaf3Fe4Z3cuOF4e2xCi+XE
MU9Xq+0XlR7JVFVunZ35C4YH8ESlXciKh5Ug8SS2NdFR1KBeIKWq5qjBk4htSQZP
97iIrLxBxNAkYN7RXVfG961C3Y8ECuS5v41MRlhyUa2M1ZpjnIHpm3WdFNOfDOOX
PliHhu1C6T8Dh+i2Sf6Wnzv/38Vg+tEvrQLZO2Iv6mmHHOGQsofUy9/CcrHM0QJu
/3/1PATkxpRmxIPsPPRqOPvV2QfFY+8a3RP/ksoxw3U4QBBukFaMFbu4sRYpET4o
0/S1dtLr+sSWH5CdJ/EclzUq+LFBA5hNA+BNhJ7quzlkew0pQ13DgFf0YX0q+4c4
NhpmkJ4D0kppF89q9mKLqrh6aZTUc39PgxipJuSWiEZm67f0zSvO4vp+7bq4O991
23kVIWgf5/AYsqSyPF2ZjOXSrPK8TFiNtPbN8pacHNL6/GxozfcPXAUynfIrxm1C
eSNhM1WVBinp8g8W0ewFpAvlY2Nzr5G1CEtGD51s8ur5Ftqn+YOZBkUPnPMiNUml
`protect END_PROTECTED
