`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uYDzrRD0vTM6B7h1O94YlxK1annDbNqVD1korupZbM/6ihJ54qLg+seVF75/+dF/
gvZ1NRw/WwfMi3JTQQe9OxQA5hQow9zNvTrk0ZZgkhqr5iAqOSi40St47QrWAkUa
fcTUa6afIHfStD8kIHKIe4S3zpcd94CiQTyrsb5MlGpABEhJphIM1iqPOQhK3HEx
3J0MkdxRW6xLElbzuSoOznK5264RfcKd4Xkx/vN2rHm+Z0LaPU/y+sjuUgt7A6YF
NWxVUHJxmkMihF4FeyBFxtLSz50uPGhl8N7lie+/DtBfVj1/iUuiwZBF23vLbUGQ
Si9W/P9giDxFi5X4biMrS6mO3wEM0TTswNMdFq2cRu8XIIWFWPiRbHgRFQFRZUaO
OEyBCbWoFxpNbGdwrmOBS/Vb56D2+GHn+FHwirSgPCBxkTlOTd3Sopq0C0m5yuQd
TgTxmbcO76dZZZPphexT+tph5RS2RIMhZqtdV7N5azDPUiyfITt0G9HC+zgS2Vk6
idMcwQoA4TfeA+2YNoY7c057ELHQrcVAnBbPzSAAYF6rt6B9GgYMrglIDOsCTkiG
oZNb2IqYtf3V4XygwgTmW5KTDiyFgfjsdWM/koCPdy+E3wIoJiSzDGvyAcZ1JcR3
rPMuYLv73gNdQQwfs0/dxKAj5O6eQbDpoLFggTSnJZdMJCbHeX9JQKNWD3sRp1Zy
stwi7YTbPUwvEyy7iXWaJLOzrAxJMh0aVXr3zRcwqies1Vua7zCwaYvmzmcRpY5H
tNtlRPCiGSeYOThVRzXECQKjNpJ5QFW/KvawepbsZk3+8pMnnPCER3VS0uubiqyT
Mjj4mR/2DdQj1fzILr9dt782paVDq3MO8KPcpZ0yPm3MfR6rsKwgSibY0RT402l+
fopZpfAb0mlCEqqB1b7Mb7ITuW4ZohRBPq3TBU/cBhIVYB7vld4nmyY1P6RUmIwV
OxJMqUVqdH9i81DGeGfnZg7awUBpcTBBJa8vNgS5u1L82fqv8jCzd1aixKRfgVv2
B5P7edMcqocZlb93Wx/6Q+LC4X547mmFV2x750Ak53UWBbb7NQzRcbh6mqFF76PU
WOt7tEYLDOrYYSCjMsatwk/ktjxXVmaeklEvcg8UZ2m5SfZzi3dxqjPxNs8vLmoq
MYfKHgkTBE72V2Xq6UcwqzkeWN+CL1YE4lJ5E2w80hAXltr+2kJRiGbQh4I0z3oa
kTM7pxMucCaqM7M39ZsIyEAHUrWdiqiFvmkGpvi8NimJcvq1HIMYPliJ5aAGzHro
8iine88Zte8rRkuiSiYFLkOGrznjTcbi6EryOgCv19t/uV9qrIDMZZmZbB1CyW4w
stWy210iwqWQNXgcTzliOMYpLAQJPEwqH/RSt19BR54F3OBJCwF+e+z0Xh304aNa
6JEln6gpuMQcAoIdTbOKsv66HGdmHfm+qiOYWDJRedXqiRQL9QMuZCV2pMOzpj4y
znCj0mL4jsp3TSmNTlBUTmsoucmaZUoPIKBY5gnourBmiiEeIbkUxhnz6aTneVVW
n1XGDdJ7knYm3ib6PniXNitbBNm4IOcPGFSIg18+yz8wH5SB1PFDQyNnFFxSR+rG
z1ym7r+a5c/qRFscUuxA6k9GH7XQnE5ruQOZ3ExAbz8uS3VID/h9G6/hK0HXWBtB
GnhNWn+fOoMktdRjPSzKiTCPQbp8/thzLNBQRJZe190TJmJCNC2QkHftgV5wvxwp
SnyCAvb1E7FC8ePnzvu8LJxNzl1Ob8ND0PS9Go3FHXTbFuJhrDbM9OmFgJRMeU07
Zo0RJC9C/ia9e1tHV5Up0hlPN3Uw+oXN15asc1mzSwn1AmBWFrEhLCxOIc+tJgXM
3RIaMYBf9t0RRouQ2mXIZygjevwmgmp83aavGTvdLI6rNy6tfNibnAcA9BkfEkfs
1EiaDL9yZ//V/uozdvYQvs3RgF1DqeH+VIL9gKhUMUj2vop3Vc1JfdinuAdkVQjc
5YdbXqhkm28yL+9zEqqzSRsVxWh07/gy+XazMi1C9u79sGZZ7Qr64ioEw/kSKXyA
O49pzZgnxjOyQRmeovR6BOs3zTLOy3py5FJjSQYPdgNhjkd5V/CfWySNeSlSkzmH
Q4FTtLP197FhZlPxtM2tI8jvEenVsm7Z+aVf5sMCkEjFoGEI2WRqxky4TgYuvd3z
WmAvmX+luqG0Esoix4ZlwxQ5F02GjPzZtVAe9SNhiV9baQTe20ZfDNC1JQqbjBxq
2PP9LRze5Guzm2ZZUg9CQQKWyvoj/jUwP3DiVpWj1zFYsKsfcGorLA+x1TNW4Pjp
+jqsSzVraiCT1NT/nNOE97rek4cCvCghmmyTOBJ2e+qVaT9es8O+xlaT+PoT1t+r
AY+Z5jTucFab6TMzHVES/qjZud833XT869ncEAS+FyXNTDg30jfWTJYL7i3JONla
yYq8+DYBYfQvEa2EcuaT+9Fxo6JrxHG9E6nYUuhEOqBTgs5HKQnPoVSBnWJqYCxn
EU7Zu+6G0zIXR68QnN0YHfUDiL5V5lZ3xYSRk0mU2vB7Kv7Vj8RHVE/s9hAZxZxl
eYTN0t2PqxY8REDrFFRLzfC+qfnxdmmXYt+Pjh2r/AxAXtNLmRYRUcfhNS0XhqjS
+0qjAHvzJot1bJ2Hct5DoEyiYPY6vMeIYKN92p/EKwALboy0rj1x0dkYPWbuddqC
wfAQ40m0eApunxanu2a7wmW2fJgXUDtx66MQkwXFhTKb0NnLrcNyngukh+PgcdcC
phI4EKNdyCaHxarPCSFGsZVwbfgRdmqa9LUpqXFVbxU+VJdeo/oDXkVz9327sY87
8zb2HLQhoQ/mivpSVAIqS+ejdAapmpwHi/onWM2p+qxfO1b39qNt942A4frYC1rm
6hrFpVkHB+OVzsFV9LC8R7TYBTQRmAflmgdMWpyi/0fVl0QZG+DdJs55raRYNkWh
F4pyglr5l2NaaF8fOzTXhMLUtI/9uMUPKvH2DtHYjVeCL95Rp+jNnGXpVNH3eXZJ
luxla+aoGYgCxyQtlXndhzsJ/Nm/qUO/Hbf5BIid0h80o4rA7xf05zh2hJHMtYEn
wlqMugbmT24xOJB0D0h5cjpudcB5Mcv4tqfWbTz4b/XdWEyceqQ7go9Brtfr4msD
v092PkR0cYSkA2gnapPs2QDbpnarmY+ZaNUjC5eYBU15rm2YDGI2wl2DOS/bFi4i
1Od4gIMDtQIbTvEIMJOJNjDZhEo2H3SQtOFF/1PuOIXpCPDAeg8N89sDz9vnoUch
poLdSCDXgm3aGaaaKKyr9z1PEA/9UyAQQjx5t7skfD4vsozPVDnYJKqKOHxs0tZQ
lHpvkZauc58X4+eh1EOI4ztfTnc56AAcz6/PPqT7/TAJHbVy3IfQuCXu5Sbl5FSB
gLAj9UEkjPkVawIrbe59q4WralV+sNIa8SdmlCeLecmyL41zqE8CeTbVnJN+PfOr
Y+tbVFJdcebwzb4+gZDawZXltTy+3gPGuvs6JyrWVMhMuIDv49y5HcRd/Z1zkuJq
EbWWkiqcGyS7k2lae4HmSwO3F1i8kzIVyBnx1msdDQlgPIBxg7M7x7Xe76ahbTF7
IMhdrBTa7g1NflqaO5nEF42HTV+Y/SdKlUW0/yiipiCih90M17keCmWnE2TzsYuy
Vjg0+EBhelfu2WnNOncSxhkbHL93DORFHdIQGWvcdkZbb6nBlygt1go8WzFUrlSg
SG41l2S0s9Zbw6kIhutL6kg4tQIyOb5kUO+tF3/mJGVVddS+ITxxZEqO/Q/+sKpM
n+YDpTylBZLQlVX9j3kxP0ARSLjX4qPuIHraEbWIja9jl6OzYBOC4D0jan57SIuy
qjeNV2MV70L9fAYvoaxxqKaljfkZA85J+sYW092/V4hc5PEo9Q+knigNu/PT4U5k
qVub3K7hdXKyfAJm5zwHmILu0SyYfD1LmuMfbZpi6vFZW6D4gaKm40QPLfnpYqXo
oyYoisLXY6AO5CIZffvAjTT61orQbcTSxjkvQ9XbQ6s=
`protect END_PROTECTED
