`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SjOF8mXGSA8J+DBZRzwnHJ3DparUhZmG7UCWPjI3FNCIrc08gT6PLocuJ2j27SQ4
NXtCR33eS6fFR1R5w7saM+TFLEVnQ9Rxr0wold4GUwlHkUX8+WfaphneEG9dxznH
TFZ8Xg9GVXyWf7i32Ah3MsUvL28SBUwxvgj1A5YDLp/ouBB2jmCuEbQfnwKmUy1O
pUHgYMlhJvP2NJXH7bcKpO5raIxXWPGXdDWcwMVyG+Vks+IZd17Lq65ILjK62EDw
wABJfgjpMurNLpzyEU8HtBViZph1UWAxL0/iTnlu8sUkDH79rZp0DoOY0FWsoSKY
bKbaMH5ORvmXQ4Sfq8Scc/2taid5OWLmO/hXW+wi79tOYQt7tIDJIjkD3Kwb6vs+
GmTbGx9gi3se2n2/qGT1AnbE7IwePUUExb82okAa7YiYy3YtMDq/E2ZSf59o4CFH
y1Lr+M1eYO9G/aaH2s71nQROR0SmBM9Tu/YU662D4RjWvLSaSlx+upaGyeB47d5b
VD5mpc8h97a0fJmxKRWvZIOCekZOv5cHpIV8PlfOREECIuiDsopQDR6B44EXWHFt
DEuirtLlny6ycENsLAzUkfa4tyTuCj/KWuhggzK5AX3hA2lI11ia9CU50va8ceE0
Zmw2dbgSGKGxh8peqwD+26MzQvLGtiexU6J7qdSnSFSvtZKDwW2pJN+J4n2jStJx
u5sMFQ/AgtESR42rauUKXw==
`protect END_PROTECTED
