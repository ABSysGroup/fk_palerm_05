`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+jSFhsTS83KsbsoMJ1hrSIgB/fYbY173gXCp6DtC/ne6zGCWkh9Z5lpF4ClwxkS0
W3eNh9VhG4ZVFy0uF0kDjr6OMAsPNWeDusxR5rN39otMZEOYGQ2LI74ZbjM/iRWT
BRKqKIeJ8rKdN1pO78tpbr5+0nqyZ+CCS1T2tFAitFFnA+DNvbl3pbpNY60hoyAu
G07S2wP2Y5KgIkcYXa9iqb7/FdNr2QFCer5pnLRRHN8yFk7BaKCKZnbpwt8oc5hQ
RwkNIlNyVNlOlo6+EaImiWzDkPrAVgKJjFboyMI199cOSdwjvnUPOJO0AaWc+ll3
44cL/wCiNClnmROlK7L3DhNqRpWKqnoXS7aEF6jkVNjiD5QYxJNUnCap5fWububg
PAG8zdRyXqqTxxc/X0xojOvKSetPJaa+Pku3p5jyul2mLPqZVO93Mntv4RraGvSD
8bcrCGWWxnZzuHSeMMjvRJu1Hi6o/O9hb0B/ihOFJI+5HmnkyB2utoZZuiSMFMRK
H+EcXTaVJ1TAxRn4WAaM0URP0wYgtqj2mjrQpIfxBjS0yvAysDWMNkkm7JyXZxG9
Rj1hxQsHrzSL9o+qPPruKNE9AzYD0u7zj1wXKlAUWksUMfP7+5vQ9qXqrRhf13/R
qFwTn6ctXJP/79VN2wChP2vPU7HIkKFxDwKm8CqJDN6zWIqXR5tLmMkMaXX0kFuR
`protect END_PROTECTED
