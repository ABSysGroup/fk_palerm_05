`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CW5QdLXP0eq9vdz7nrybmtWPm5Yf3o2JQYMqigFNZ9YEiDX/4KZxfh25p9bJkLBp
6FTJ8ZLMSAzX9bVbNEQtNwu4502s24Ru29fwvHREt0MKQPtU3oEFwdI339z4ehyj
QpW1PSL8JmTgNyjVpoFpmUDjJj/e9G/CTS0krpRbVNj95cYjl5JYS1ynp2z2krT2
pbfYRZxvz+FooDdfGrxupCyugbavfC8c4Z4DJR41LPl3HCdIyBjkc0dVOTrcdm1k
ERtEmWNx0fpCKHhTpgEUjFnJI5eWEuzvYbef2sYlBNdNrpiQcpcKbU6CHaNDH0sH
K3xvdsNFTuza/hGS4mJ+BG+y5URfmv9zQfkvaWxnSSIg4Weq6ZD2YacAHv1zFJ6s
p5zqRmQkxDzLLC2uda2SZA==
`protect END_PROTECTED
