`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
roycPysCvYTl4qEhVaZdNIt8Uu642ib+2S8EwRh04vStM+BU0kMvZiQTeBFDglVi
GzKpAm8uesllnWX6s7nfyNcPiOHsWJArtlJeuEFQs6kCDyy9uDo37aHXPuQSydOY
419kBbzAXr6YOeJAiEs1mxVXWxYiuJpJ9YARXOHuMmjJNwQ+iO3kCieiEVU/lId5
5wBxKy5u7fcBq/FXyt2tMemxDZ/zq4M4cE390OLouwUtohOC6nHoEztF7WecWOXW
Qwp0ClWe9KILrUjiJG/jd3/EWyACNvU7HhigMpUXvJRCf5L9f5CyACCQKZ6LAw4l
IzylCvYNY98JFfS/vua5jVqkgJEpduXXeS2b6bsIgFKcEPYjNEQzQV/VvnjLdV7J
bSvAyAyu9J49iyCw3U1U1y8wt6PTjhUZMivODjozPN4DR7M5vbpdvkiRLO8341hY
FbznlN64IH4+ZYP75gI1V9gPrpaZyHdf3CePLdnrtyRtK+KFOBd/0vHDqo6quMPQ
4hB8RoK4Ar4AzwWvheSn36D1wYnIz+x3oU2ivbfWLzF2NH/GQS26NEwjyZmrDTGE
Lhh5HMok5zimpRQH8qzMzZ4G9AF+p5wZihXoPLMaQu9ujX0CLweKjQ9JtSvz9tKj
iXf9c9RPLXrWLR8Nm6eXmB6VOVP+h5aBNw39KxwdtsYfzvaxjXBIwIAwmaRCAJoh
byup96MtNHQsJ1ExoM7+Vmp0lS1IVTumbXerm7lE7cn/JT2SPyIXO27cO1FsrJOP
mIVSE2nGsYhTtQl0hFlEccFL0wIyXdKt7XlUUR7+shr8UWAAF13CGIs2qN9XIgY5
lT8Lm52B47N45CaArcdGmk0oXlxVwHglFMrp59M1BZdSdPlf/bQUY7LSRXbJ22Xb
+0FDPZTVeEZf8HpeaVg0K5gz3CX00khQ+6LbMbpWrl7JYenAJ0ShMe3VjNYbiVQm
IQa0GvgoB4ct5Bfb1mnzvFdswrYAF1yXYOn2CfAW+/CsMCPbOFHcHKsp5A5qq3kQ
InbeQzotbbhuUTg2z3c5lhlPMucT8RyKxMqnUFmSJCTSD7vxRVc+ookMCMIFeVqg
9kHh22QFUuvMexYraBLrlZ6ovZkapS0mNR2VD6q3vTL9sAGTF+qPC0DdDERYdBaF
XcQtI/iFgraYb+cmy5aOH9PFTMNzN7K/WOcBQtf6qRepeVCB/Elgzf79FGAMS1p2
lonJBdABHw+mBGGoBPRoSPGFxZtuRPlOg9LAXFR99F9+A60ZWAvcpcYTyLw0axDM
UxP+Pbf86IJ5h5ovX0X/+PsOKYwp5vokP0C67Yqy7wvr6fU8ClrdTNo8VkWm21tz
UTkjcj8sA31HPcGe6qTqz8SZmkJ///xwNqUSc8NxbdydRk2Y3D2nbQFp5a8toG1s
kNlkWJ7q+abjR8iQGYIRWqrvbE8bzaDIVNkkUkFWs9czDlapEdwM+6Xlbzy4krAs
mxD8eCv8KH0OohKyzkbSrHL87VEGo+bwnogmLvyZYE73Ij/aAaSAxgpNIVZByLzT
k2HekzhcycoIE3Hm8fE8zloYfrgbmorBpMh0nTqIv62HIbCuEPsIqakU5k2fNlWH
N9K56aOSFeCHIM/93IHJXG99xavyP7KsfFh8n/avB6xZy4R9YnVnVA1uu/2wk9eR
sPeRMFRkJ2LGgtYB2E4LTvzw6GH2VkvqcpkYh5CkTTVHzCy4OjNxU+mLT1ZB6WcX
DWjWmCZkqZOtB2SSRH6ZuP2lb8GiRP+1mM93Evq0JoUTFd3h5eRU8OkVeC/8rvIo
8sZnRpwM07oiyX3yU4F/w0lnjSY4Ujh4wyCLvNZaDvMkGRI64MnMHo2CPEdWSaSh
YKRxllBAxQuWnd3g/bscpVBKDEyZpGe9guFmQxJwwwj5VG8ZgxP8/mio3mt6Hcf+
IMIi0n2mAphBgoohT7gxpEeQm9NQmHsdY0qlFN9ISiaQKJoTLiDJQEqLrQlfDhr9
Jyr+xcsCqJV3ny3FSBU7nwaOwaMfha8OGMyFtSCmTTMNcwP9qo79gKLDx53axAtV
wJtaljt9Eekc6rLWJQRWfu3TLlYxt+xLooGcHSwyxHqrvJ/t/eOtIFG6Imspq3P5
PxSppWVxDWQyx/7RVhcURgCyeQORsa/9ETrmJJm9f2lfEozUijuA+omO3krDUI16
RvXffOb3LWZhrUn8DEbF94sZHKoBMgew6MBHKgvJ5LgBvmDi2Pciq6G0oRNZLtQc
tvW0ha+spsArJMyOcRN9t4GdgLFimwtgK3zCep7T3rn9wEgRSxCDzmaBsbe7qRa7
EKB3ylZDnpFqFYYbcKjPlkZm/mI6iUyG3r6NuRnqRGAywob22HTbXhPJYmcfBrFQ
PiOEiCsPqK3dXdYC6fXYVOsZYPB88dOkTQy9eC9ubMfKR3+kclefMk63SXJ4nAE2
FX2G7WFiKVi9a9iObcX7zYD+byOU6btceV16zhnoMcGDUb4B/8gYxtFCMcayZi+x
QB0JOsWQwf17BKUx3A+LTj59EB6tCX2RSixSwIe9HFc=
`protect END_PROTECTED
