`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
533r4kOUjP/HaHI/476MB/T/bL00cq9vpO6xHr7BpoojNKJM2e2AsZq66hY7TtAf
Y9t7EOBMGRC53fF1IzaPayod3z0YM4cMPi2rMEgcHwUK0X4Lj09rQehLlFkKgEHk
Izn2ix+kj06F1LvrXNVcvAss/3sNF4C81iZPh5iRK1ct+IYQut5QtfCy+czHXOvR
S5vGrE4JLpdf8DXaZqvcIOnoaIS0ztGNexPp8fjxgI0pRN38dv08VFU/GGqY9Rnu
UrM6khGb5RP3BA1qnIRX8Xj2taCaPhmaTULGsfgAQTzAHvh+yf6SmPt/qdWwBzPv
1Ejq0Jiexp2+DxnbRqHesw==
`protect END_PROTECTED
