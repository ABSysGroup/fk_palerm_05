`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
alr9D1GEtjUqsA7TUHkhsAZUMLLvcw7e9j+f0FZQYz9fdXUV5Mx6ohVsETKCjPgk
lPZIW2FaArGyGvaryhANhpy51TfpRVAuFHUY8mpeWY/ed1OmU2B/+3oJhiNedfz/
hRll1/ovFWUgykRej2ZHvM7gaxejQJmzNDVU5sL0SVeQEwhdL6hsAQOLnEOgN7w5
05fIFIdn6jO8zAeeRq5fMGEDLmkD3ahQNgKwossAUBEm+zHbjY3KvGGV4hes+V4w
1FoRkFlMudQ15V4fKdIQFQ==
`protect END_PROTECTED
