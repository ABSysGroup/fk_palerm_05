`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wg1IELgYlADuzqPH6E3mnZ3GT0kd7ZWRCEsVQKd0z9EBmL0Vv+JNNU21vaSCx6D5
UlKXMF3SAXjRuBjiZWfM2AVKcCelIsyc+9ViegRpGdczIFa0yWLsa1OxsQN6uHde
q0eBnJV07dEhI3BQr3BY6XRemgOOw+acubqackyH3kquCFI3O5yy0xNtxxyqyShy
8yzIoLH2Q7XKA9SK0kNmqP/fdOvA5IsPfrif9jYV9nTfqSsfdj8SeSBa80MM8WOd
N/0GYnYq0Jr+X8feVyITKFbdhDLEfzyjUQSzjCi1MZYJ+rYMMRtuoUVEpU2dk8r3
Yz8Pz0YjYUFpVHxzQ8CMKDI7w4Y/9NYsPzDTKcfoSIfRkTUb3lP09MzBCWdyNtFK
RW6mOQ0F7vquXEa0p5DXopYAUwOLQqnO0JDB1cecFXaD91L3Mxo0e2On0yR5giZ3
LrKXeY/UhXjJJ47cZvh/ckYKPjlZKmuont69NfHqOOaFuzX1YUEH01UJ3U6/qWQe
RzSpAbL/QbfmhJy59de4PO0Q5ShdoQLa2ojgGI+DjVTdZ5yomAHiUkmtVGshsxFU
uYFQABK5KlHBT24RnmTktqecIks0YR1pHhjxvjHCybBgT6C1Do+eFUQ2pNyznQPF
caLvGE1E2D2Jt0Np+3vMoYmTLxWvnBi6jlRuJwo8jJcHsxsWlNRHAjXPedUY1IeS
8Qmej913gRNJscn9dyhYjFH0O7PMwQxsuIG9WaH3tHXYyHsZjmlmfRdOC2jalcLH
AxeD3puusC3Vn0a0XHTD9BvcYRbtc02CuL0d/QrPYH4bQJPxNNV1Ai4D+OFNOL5U
xnywJVAA6dnXZoYvhZA9Th4Cndz2b4wi15O4P3ZP2ac=
`protect END_PROTECTED
