`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AR4bpoXS4Xsky6DaF7NHArpoVMRy2ppy2p5iLjhJsZAijrWRepBKcPpu7PCsTFY7
RXDu8gqEr1RND4QH1b32/oIO/dlkQ1wNh51PYNbYGtD32F35ZRPEqsMKuQRQVhqe
qeWlO6sIsWp2Iak/gcEQWo+MqdXN8mTI3+tzmqYOq2lWS57GrJyrJXGASqmDHxcV
M6AjA9myyVq5AAZwgBQwERo01lbVUP2Yx/IpnPRuIbjw4ty+M7ykOrrlUrtnp5B0
ycwsR3d7fO/Z+Gkahdt6BsgyGBJsQ9dyWDuxxg4VbndT1NoMasQM/ze0NfNVgUfC
smBTabtrhrT7vcQ/QAZnq7d2NQz7cDLJYw18Tjngtcg=
`protect END_PROTECTED
