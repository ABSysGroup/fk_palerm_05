`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bL4TzDDG9ML5rEzRAD4Jy2YYPqpQmzFl6Hd8pL2EboBBV0evj8fzl+1iVEIeANkd
R0H7NeyVw/Wvn6HHjJldW8nh21VYE5LMtmLflNWGIyM2HrQ/Vg7u2ZNzAcwRpwl5
LzJ9/n+tbPSPUNKyXj4HJXbmRC4p22qq/DoECgq7+mEMPclCzD6DrwLWIZYwyMCB
LptkYnDbkHduiQXfRbB7LSkwtNIXhSCyPQhGCTZ6X71CoeJ9d9PdlC84A2OeMBww
4FeYIkVTjxPnUYKF2kesYynK0Yhm0vN/ibNP964M7PVVmfR7vzthMl336GnI6RVa
Rl+lV1rPS4jGNfp8casj3ykVkQGb2jUGJAU0YEa0YxJGVrP2AdPHXDoNWGLDCTN6
HBbRmBWlPMxcnVYJioy4Sz9eK65v3oHm0KOS0Nz9qZ6HLaxyDDpVZcGf/qwnC1eE
IEPtCfUV/21SINT5Wt0KzHIMn5fjh4DtoAGlsjlJ0rG2hOXBwiFKk/WPZKnvD0Tj
A+32Apcx4WMbcKn3FZKis5FAHnSI7DwFhawNPZunAnEEGjWKmP+owFMx+QSpC4Ux
htzOLTwF+L9Ch3W+HT7Y7YBJS9+cOsnblJwpNCa6RSbcwbyUdYGLbnE3e28lHu7S
WzOPuxIDkrI7HT8cK9seFrUndb+yuvO1wFfB9+xYJoJLvwtXW3zsfMC7P6r8rq6N
TdS3ID9BBBIIH3LeVpCxyxSvFpE1+eodYZNfP1KqLxSmD5TKFoBCZMP07ezpZZwj
k3t2YowVOpplxsOy48SjRXLAbSHSMILoWW/s0AJJ3eYhP1pLean33s/iGAEgxuLt
CzMan0Qt196/GpRY5XiHjlH1mNNhtpHP/GpVZ5L+t2SvXnQQEbNcwlIjFrV8Nag+
ApSwTXykHKJrYnEvUPw9I0vgdZTUwWXyE1UwVoCKaGWi7MYi+8ZrKuPPiCySFl2l
/YqlfYz9LR/V5pd5JNq5cI4PXYNxdRkB9D4IsJR4tKs4wpIlLscVPLJ/J0/ffCWS
+oxfZIHabqgqtwJBb2bi17hbZ+XzX2ZZseiHXkzxlD3arKEPf+Dw84Vjl/AxG7XB
0tGxh3GCxAI+DeIOozqzjRq/6wWbh0ge365A4womJOJvVCC9TJyPdPLHwiiKBm8x
qciHJJVhgNFvbtmmiHeQkc5T5pPjccePKEZMHN5cK6e3E9cUcDLp+vMwwIg75B14
MWf2cEgWTZWfWa3Y0W+DJI101ZloIhmkakw/fRHP38YdTntq73XAYsqCH2gZqFnm
DM7GdL/E96owFUOAeVJ6uR0YKLsv+9F56FQAsmfJjRh1MBuWx392orPooJ2VHVrV
w7pnreeJUTA5ySK6j5Bs8S8PiBpno/eAkceY9x56jGRcmqHQhJhS1IiQ8+MQpSbG
RE3EqUdm/wGBhCLw3r1Og0SxS1+bzQRuNuUt+WAGlFtM4QZ3Jukl5wqFGeX22SlK
7uOUN2jCsozSU5YM5TKpNcMqBDR+WXIEv9ATp5wus8XjliJg3lzq3BxaUF7PXgDy
kpMbrGDzd0TYFFCdgNvBB/E3PFzk32JzzzmVyrNYMMSqP+a2j+brYNGDF564VKEJ
L4IxqUyLnFp3oyJqQZLYm2mTsrK10d3/X9unsH00Kjqn3TUmK2P9fizti8RW+K+i
NJBrOmO9oK+VTI/0g39bpwqniNiRQP//M7I54UxkeTQdhckrm9fwmkY5cw4CBfKe
oDsfNy3GWAbh5O1dJCPr26IB5rjFaCrxKGeS0ss+3FptaiPjP5rhlWUZ6UVaQYGR
SNx7It1zDGN5LAkYJ2JU29AeFYt+WCtcJ4iNxjB0gDbmGBMiqfs3DZ637XfYyhvG
lJd2yPhqxinIMiqLUlivfNMvUI774czwvgJKb8zvyhqc0CLsBnzWK2n4y29EwrIo
/kQZ0Y+Sgrq05/J3wG81mBbUdHHHu6hrcF2PN23MMFaRolzhY/6hmFyZ4Wke8/IT
98GzGGVz0PoDsk+GRghEnLebdqrUINelS+T+jQSgR6OKLtbnAgAmxYt68s3r5fPS
8m6UXimgr4KbGboqMzQ9rtcrxEN8ctv4QRKqREBVYTfwEfzdY3lRYP1XzASb6YQe
Hkj4JZM1aPo/VEE4OZM8HjQ2jXQ7oXQ4AXVsqEoKvBr09QFVE/ivWc/wgdTEbxtb
C4c8xsiLZDWJuM7okr5nduxY+X1gYy3JqyjIjW7s/albuKRWQtIcYMSiohvFaXDB
xJYcmpF0LmUfD4+F1Hw3dh2I8J0aamVbWu3IgPbFF+k70EhH8ymUmp3vEmchtO1F
gilsfoyV4YWsflyx7IodiL4ePgnCwagqOkST1RSK/JkHV2R1AJFgkhzsTTzoigio
yacqtnt/BkYzRY8iAOH+XQVfa5rZ1zgm6zZpWdReJmsSt8XXoIcsFGxqhIxFHSoy
1cNuSMa5GDm52mX5F5pTMm9V+AP2wP+r7yTyqbtaWO2KNzc6Qodnwh6kB52tcEvH
XkN8jWFNjJkpKUYHE6Jw0ic0r1JrzJ/yXiGJR33ryaS+DCPybAUJfYxxvyGgr8Yz
4Tau7RPiFGYaBoqHIqQsLeoHZ6Q3JVPmfBgfeSzC8+bgyHB6elpw/BB6tvy+N6FL
QULce21UJLDw2J1QHYtDwKExpGMDNEa5oqg5pfuU0YMzP9Sa/+8ckQzJgcMFf1BX
7ojWMoCt/1FRikqgPyhrdgSEG0r0ztlgxUMqW1RSksE5EM7YZnelBOzzQDBjXOqQ
MBkvPhj7pC9wmTCwFBtErB0pC1/ZuMMi0yKMpMbP29BmxP78W+SeUV8Tq5LpX5QI
ylTH1ekdaONmMEMILwPP79LTednhYgX+gSkxr5Aqc7EstvKwfe5VdzXkdAV4dHyI
b8TVFwW9LpSwdvln2d2+Ng1oct1lrgwjmLNhqGdtlxRGWz5UbdHcPfbV2DTjkdDQ
7u5eYjC5qAJXOpkS2B6MDudrY4Sc65pPW8cp2Imxdvj0sSFuyfPSrNI7ymg/NezZ
8XSA6FdZj3Sl/ShQ4pk4OBlBw9Wc3LX32wmZb1trz6+Fjba6mJQWl9PtJlp0SfZF
nrTE/QR1e8Hm4+kPdbUDGUSML1LZH+482K2MKxjYE8sqqQmGEHx+q740exoY0gOm
htDyIHA/h33rH75B2RPO7nyutjkcXoi8G7qEnj2ANKtViMbAm7ELJ5318kCk3BEj
ri6EeoncMVdbL1guZh+hXs9YNeHbbSreenlz0QH/HWQEQL94ujmI5GiavPyZnSEL
hKtR/xROk/Pw+qOVFaO8zJkyK6gz6pCWCy5PStvq5HBtm6vhjiUAKX2J5ASaldtC
3uHp2AAae342UyC98HNvPUjSQ8PdpwKL0LHATFQJffDNXS92297wHmzvHyyCiw0B
woWrdJs0b0UFi7wf7MhZqnLqZtnwsjV2Avlc5vZy4gRYOYGpMn460nuKZuhkMlZL
HcG+Ot6QmavhKufCN0QskQhTOheis4Jkjvu2oxHTXvYD0tq7InP0lAN7n0Pu7sP+
IywR1NPLpYx/thG8TdoZd7fzRz//oK3c73qpMRXJjl3qq9BrT0G0HFgz4+3K+Kl8
Lo9SPubbBXDU7Wq3OmEBZCo61Zz9lXa+BIixGwd5sw298mI6bntjwRoAyRLMcgfn
MRMwbkyplYcooAvgPO7Qor6BiXm9k1IIesGL5Y0wya9dZ82zR2gc5MX6HLxLHvYx
YJKg52SRZmp25aR+T0gZPfOHEmk91jMLi9hI2kNjBRlgeJEiCdawC/s81SnZ2xqL
i4skVrBix03US16K9Xs97LIObPVd8xZ/SNUq2rkDIO2wlNIiPjxaL1pjVgJr8sI1
swh/0Fktn0+gGyoZIspxmqkSWGdPQ9PV2snnmGz+/Iq8flHs8lqssDvpSTJrPYxw
ggfBON5R6lgrKQvpin4v8nPo71LXu6rfRHufm3LE9ABayUHqcX49QnZP87aLZgNm
kGz7bnebr2cW/9Ti3J3IhPYnOO6jYPtjnpsfDp061wTl9yAhLAynQuCdpEctWe5l
uj/M2g5oWfbKNk80qwq0oQyl9a4tLWMU0k8BF6Hxnyoirmv1/QQ0ry5BrDN1S2T0
7L/YQ+zFyCvqnZLP3zRChpCYclocKo5ySabmRGD1peraa8R4+q6P/bAmxfc7xoy1
DKKGdyPADDq2JzZ/TCfwYuYj2YqS5D9bQ3Iam5AlY/nhiANiePKTr40IqIM/YPLJ
ZSnnTNCuPJ+c9X2yqDUeIdyHwZOEM9ujIV1/U3bBXAyGBtx7eTmDrC2Fh0s2HNtd
y8Q8EDd+ItzFsetsqYj1WekN0VhjxE9dxsPdQHHX96EDmFRjesMPhcu+nz4HHhGu
YVxNz/SaQtCMwta02W8cC9v5U3tBj4T4oN8I1kOxelaMBnp4WFzASd/Z1p4UfOeW
MLqPRNwLZemlS9oc6fSUvbFHxqYuxkKl8Cpy+ydWr4Y=
`protect END_PROTECTED
