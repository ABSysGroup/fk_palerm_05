`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pXzjNNDDPckMo76l+dbeExCzCYStRovyppEPl9z51TnRDnV7EBxyAZ+YUCsHVMHG
5CJXcE+T4nsdFsKoIAYepgko48cL3emvuy5Jq0Av+eohgTBvd10kx3luD3B+sbJS
nkTbLeQaxPGt2hM8W+eIVjNAPRwH1+hmdLkHZNJ/LbhP9BvdeMnq2PB64mmXu7on
fGC2qefw3il2VTkM87qIbMYjgzPnNQvsnXM32EfcEUnWevqc/3JSeXN8+p2DB/Av
7b7MsoQTdXgujahwI0DBdvagNzRoZrPDhIIhUyRja4a8u84umdZlsmsLbk5awz6O
GLUuJMxDAauiVVwdn+NTf+kIQUTM2FP1j580oLi9hoaZHskOdoI3Cpb/GDkXyep7
qEDX08Cqqkotiv+rb/GKFLfpTDQOrYcs7JbHESGw56uwClZ8a+9AZ7lOFx6Luev2
DlLbN5G1kH5rna2+OpnkhQlZRGUQi5Pzy2fNXqiNCSGXX3z4hrCOOeSy2lLYAdeA
OAO6Kc1r8+0UMWWrPylxqRbPaewfb8hc6RhR9lRCTMgS7OXWwtiUsJ8Vp7Jwp2ZO
PqZPHx6a0I5D3LtVplgyESv0j5loRXiOxeINifT6LCOxUroKobktdxX5FDPzDNe2
1K/wVjgLU9nPuIi7zEFvBoXjEisnCU9V/7b042i0I6bhr2ZoEfHHoThfOt5N6W/H
qylTgICSM2w1zUY4KpUZg8fBCqkyGq8rRqbidEa04HKs46O+TNpGjCWIW5LeMBBj
d79EgWdQerFRqrPtEDhTu39MLbYOhIyI1S7UjsTQ4GXnn8HZlDFNKu1F7ImPhzsy
ziB9nqwCCrMpv85TTO+74ndtFYIMoDumvFAYVCnInLz6FuUm7HBqLZK34mM1h46p
PPzDETWZKTT4VWpE9U6wLackt7UpIjeBsdv+EVI91Rw0lQNkPE5sQIGFEAQjpMLn
h8hbWOh2LjpUKKFsUvxzQbLGzP9FZqsAJqcL/+8uKAqbvc+1tJSVhtPpt2n0xrtr
8LpswQxqRvAq4h3ulsXMff4ieLU+whJ658bYsFfnAwQsiSy44iw7Tr0rpyqrICcI
h14gMYsirmm8fWpPZ9MvbYY+UHJK2PZw6+n3imDdkjW8Bo8uSLpRkLxg3+Ym7bit
RFb/2uVsvsCsxXkPFQzUIp1VzaJD6MD6bGWqXJMOGb+CwrwK7U+l+nlLOCq+4jaS
Hk1ENZHFO+KazryNFpPrx+u++dyGq5Xr39dCIsKNk+tRqloe2XaBnBFawhl83il7
1938OSCFKlThWkfBpeW1ABoFr5FpP0ctHkOf7Mxc8j90k0OjF3br0lDRYItWwOJi
yxZG3NSD/GbCNJVfMJY4lyVRLoT5//dlIhQqOp9czbFNU7d0+RgJjDghDIyKTHLR
jC5YUALHSlf0rLuYzfitWw/shOj2v3Waac1uwRk8jlumgVrEjCXTOSsx/h+Av7i2
097KMNwcAKzAcChv0MoLvYQ47lERK+C2SyZvCvhgs7KOlT+L9nPmVn8POaYUWgnj
0gdUBIfIkD0OTweF6eOtN+m7wRCWv9j5UD2bKdudw73oV6Vr+2ReCJXXUHEQhJ0J
4efvFq0Pf8/Z/EwBwEeWv49XyG/af4xLRwlqk+I35NzEyeA9EWash0W7FUctZno3
usmMVXFQNedMwFplD5MGxw==
`protect END_PROTECTED
