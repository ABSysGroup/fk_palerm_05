`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G53rUFNT+2BDB6Y0rZVOw7pgntqEzvkMuTS5VgFxsbRuhmtTQRKOKcWhrxR2mHEu
7yXNyFHlJFPpIRc3kGrFYmbvHs2b7SOTEVb0jJT0gcqoakN3HGNhgOqiK3gn/6eh
l84MEYS66/bnx2PuwreK9D44FYztm/qwNHwI/ON5ILje/3BGI7sBj3SP/cohvJwb
uPhMS4N06GJm0rD0gG7Vn6a/m4RaKE9vydqohLtDaPPjuONirX8n0PRJ68UE+l2b
E7EQjqkV/INU4SMde/0x8fGLksUYnUxIW7Bp8StUXMFDiw2Kkz3ExWSB/tJkxhpq
poZXr70o+7wbgp2Qi+1O0+HESEA9CINcjyZ9YkHd0B8hpDxq1b/G/zOSz9EIyCis
HEHlf0r3XSwTy0KNXNtjSk3P1zytyn/gZxobC2BDgq0dn2ncuBPrZ7LP8EbPzaD7
`protect END_PROTECTED
