`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vqbAnTNstNULW43FqwCpzX3oo+qLVoSHrm+redEbbvyG57Nq80YFjYMWHvfolr9q
+oRZaWzjf9j0wCva/xgUPW8iOJJldhQ0i2RJJ3YG9AMX6BoFNyt8ZF0w1R4UFOhB
QQsnW7UDvtKyyjD7efECPFhNo+1OPPPc6HXweZz6OKV1uE2s6Nhb1FM64mA43sJS
Mf1dTVK8hlHd1rkumA0OvehHRjn1dAqAlmOKQa5dhRyTd8eL83cdy/whlALhh0oS
PcfaCjqaw5NukENvufiQDhTLEsS6Jl6jcjw/FPvgJ6g/F3Se4nh3RbCeFSO6Tff2
NxJ6+xT5NQ4mL9fMUddM1gFfV2dXJVVrLCVRbRmmfCHmmsq1h+5wd71ByvMXw8xt
r2x2mIHrWN+P9UKtEnMQT9o3RkOpU9JFpipZQVsAC6U6RJxuJ5/FBkmKbPbZCJ6b
`protect END_PROTECTED
