`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g5Bd/yjmjsSDX9jqrxHuvS6itXjIY59IWPIO7wOLNEQF53PdS0X/UoiMUafLYM+c
tVDQvSjD7QnVP5w3tQYY0FPMUFLxFNgUJB7jB18jcrdylS9ASoYQDxdeiDpIvwvQ
YGjZOE2BHeK1ek1NWVdZ5wMx/fZfW7B7KjB6/O1tnp94V00Zqm1gB7G14R3U7SzT
OR/I2e9dCyTDEGt3KMg2dJt++ArEbYSOSC/AxfKdkA0iWmtJLwY0lhP/cZ2ZsZAJ
52/a5D1IPoXdiy3AmvHjFnORICS2mrzvWk/CIqOXGGp86K1s0nycexcIzuYuEAxq
w11wWsbprtX17mSphHIjFgIdONxMHzfjDsYVjCrCYtejSHblNzPgN7faNrpPZYIe
smpqLMKFz7Iv38wnuowE39wGKw4UYZlaMQLFrIqaHBOdinKHtPgDml1aRkUs/7tu
f3WBl9XxSoEj3e4LzchNoid1OQLgYE0so7YjOuX59Tt420VMn01GSbhDRdI9k51i
Oo9tenQn6hLDLZC8CIbaK+fTsm4+jlfYLr5LpDW/BnlRBlt9+JWl9hWRNQakyhSR
010dGlF3+xs8IhKcoMOgVE3yILDZ1b+u24ofq4iiSf8TFf1gUTPRfX3/obhILoEB
MAJxKD63TlyUsh8g/GIUUNYOwuQQcFzGntPM3xZeK/xWJVQ6EZ3fdg0CFaIvuiV3
XhFATnHSfcI/1JMqwAxfZow9pl5RuZDdmgv5kOyS4nuE/807L/Cupnzm+m4ZJQ4D
3B3Z9qtGVZekT3DGsDnK8Q==
`protect END_PROTECTED
