`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x1LhmwbgxAxx4LKzR3OcxlFoOzr1+ukBFJGajOk/UeSV5f/3wh/3BwSa3tJdmXu/
RJoVHap3sWY8p3xipca3BhHfIABLWhK7odomamJJgaTHq2UiewoSpM7fFtg+8zot
1qjwCeN3Vltv8/xfAZSD9IYR7R/OEuWCdLTMu4YenE9meAHY9S9n3FGTthIkB+tv
DtWeOfVTCAJkuSfBunwBtEUJM/TeoK/tHfdQQJ2Te/Fy5KC2vf8Iuu0ZH7zxUD/3
i+61ZJ5BSceBtXmcS3utrud/E0sVVLX+U5V0V1vqEwVSZ0uzof6OlmH+iI4gTaQr
d0wunSnZXaIzPfUU4dorR8uZb92ZeVdy12Hx8OSrhQsQlzkmuBbwKKweuZ5dbv/3
+k2GK4sKXx9F9H7BGMek76qJvBSxhPLR3qe/W2XS1X9QYRxfFFCmILtDsSVE0rvM
oKh/l6U196KL3rBh+pXG8YcmlRZXoDqpOAxBUNGgkoPQiE5Nbcv9ymBrkj+ZXYen
tc6Psuy5Z2UTRq2cp4XoKvC0msjwsecbiK07AZySY08W1s7ZeJS9IronXzC80PXU
1azkatHUSDwhn6hm2SwZwcW1c29yicffAe12aDVh1/9rnhvfwZL7qWRPl1SnjidN
/agiWRTR6kUvpiAz4DnhowfhLeAz1IzcF0kS8fAUDBrU+u7mJJ0PRUvlncO5crWT
/8RjSpTidQdfILrxDwVx6r6TLVHm53+kx47zyD+XCjKr/w73VBPrtd0ZBQfqMWIh
cMsdTz1N/s748x0CZaU4FZ+C52NezYETWH+zRqFwM/lT1W5C9z3LR+N2pKH1ETxH
q1gxn8Im5vvUypQ+Yw7l2IhIN9UAhd3he+smbD7zaOWRlKKT/RoI2vqL1I8qTL/r
yGBQtIfqLwpzNt1e3VDnXq5sIW4in28sES0DQkwC+b7RIw+86RFHjUNdD9xpT9sk
9L8SzWYhY9aTuF9eBQyZARmihZpNKYTQG0KUWOgTkYqESAPyPEu0/QZ01HAf80vh
GxYAC/R79UdGX9+8uyfuB1b55bZ9JoJfAu2gL04mHaGbYYphrycxdSWiGHZdK2y8
JrCm5MIuUtdZMHgR1H3GROmbnrSODGbD7De0LtQO1CfTDqhkoRDPcqVhydsFQTYy
wMaRAYmdNP87UQMP3T1VF70R1Q61b80edF4JuI2xN8KMGxoFfleoM9MolA+Um/eM
v65kSZcsNEiDejbDtGa9ol3UxcA5tNserbIFAxAnYoEicF85kM7Tll5RVUbOYt+L
6LF8a+aOBOxCqzzU/y5zp9clKGmmYGNJrH8FaPzf7cgPauTJtUCx+gaz2SYVg+ob
gF/R3naZG8PKLDgj4gtD0qtgBEkv0Yiiz9o38fWSzRyIPV4FqUSv0jmEjKUOMBAp
+sXZtzlK4S1E5JWGnF1bYQ5Ch0vWFhCa4VnMiBSDeZ2Yau/iEgvr9Gu3l51x5rF/
EmuneulE0UWWp3EbxzJm/zIjX9lOeNWf4YOCfyEjjN6OPC8O9H/c+U7nRz6Z96i9
cK1nzcGXy3kgTKKfNCzWq1PUdZ+AttEbRUOchoiaDrgPMNuvIpypknPuDaVFye6z
JZUOylyAKlEzEMrHogtM2YPaDywmw9+wJ3KPcL3+Yy+x17WKbgvK3CFyLFVkbW5Y
5XEbq/CLo3xrytGASXWluSgAUrNi/39Sukju03RBV00TfNiPr5Is8rCZDoe7BjDo
dcfnqrYLaSBBCS2q1U8hnUdBbfgHDj3/oCDooauuhBgFyfb9pEQibtBONT+LSsQF
1ItPLXqRcygwqKIS5hfDKblblruNolPwOlPFACsWjG3Iu10Xwl6zSaDIaaKSpcvk
7l+YanVrHahmrp0p5i9XyhGDPUVfBeFcgAIets6D5ybHqcyoz2LsXxuUc5p8/CYc
V87dxemCfa3AdqzQsvcRjquKojimUPpjJwJ+3DmHHI4CetN0BRkzswOvJRv9BXU2
XW8eNFNRFZwRoRWTUU0gmw15Wj7cxoebyFN+5C0iK5acGbr/Z+rQbEeDEzjqSbo8
5oVRMLPDL/vKrZpzKsyEgXGgLsm5nVrYDvvmi4+0hfE7AiQADbpRKHUDCEJgj855
SAgeRexbxz2DNsc1Kudf0eQsg4XHd1i3VQobNBP3TIVAiIflJFSPau0Hwl2xOdBs
mqnpqchPH/aO/dkcXIfIORebW0ziUd9E/StZGs87AcrB/+YP3LRJXsDS7U6cCu9b
mMRNDFDWhO1g7daRbFvKV3jgHN+qvaC/DThC9niFP2bGYrHsoLKj/YA1nAIfX0gW
UYYkXbYVfUdKrqYW2N6If9XC8YIWIbtjcRgrotP0cVZ4yR5lmeEs51IDGBWb6lhx
yfXCPVyEKaNz90TPfFRqtZH5i6dgPgu+QPsxk5sQQq0E0ITFQxQGSuQmNIlNpiG3
`protect END_PROTECTED
