`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b+7KUZQ1kX8/21BpgTyrTGVQA+h5EWozSNlL31HW8pSTOrO04a/WaDicq3+K+v2b
ofu/RlIzzjYvbeeAPiY1vEXC9vzyHTrjL0vKGRMJUKxS4hissyFtVWhW5nZlTCy/
eln4CYOtiRzACIeVKSjCSDleTb9bTYCDOJlTb4LN7FKduZRwlEwPX7zm0E3yLdCt
4aE+PfuKbR9fRW3OP7OSqTnHkr41nmKE6AHBljFSQQt6os0Nur2JQBOala+0X2wC
Ws+kYmKjIOcTQZmUE6L/zsDrcjRAfKyJHpXcyRscq+Zab37KqidpZNCdeQEYVN0W
PqEm5ppnK5dGhP1knlxOR3Jjk8cJrF9xSEAhOqq/sq36bDUwlsTuEHC6fEPMCObU
`protect END_PROTECTED
