`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
REcHhZ07Yu8qNTQKBgNslEp0nNGnsefYfqy8wGd02j5u1I9QtTO5C9rnH6ZHh+bE
A2UBEsmT+9yBtp8ilOZSULQXIFMfvZ8pEAbOpZa8q+5cvTyGLyQaxarO7eoypaXZ
nDmhM/h8t5Ld9AZknencVPiSEuerDHet1oR3vQ6C70DWoSzTaBMBXjXiIi0A4jqf
ODNx2xooIt90o/EJD/7zQkfuUcKeT2vbwRbDdjxvZWtpshnJZcrC0Zm/Nm46Zcm7
EeD3NcV/ULzdy122MBb7y6HnBKSo1sOGtCwew5LQXv02EJ6g2MH+mRmAUGn3CodW
K/SlfH6szA8Dd9r4PdrCRFNIvem1cDvHjvL5ZCL4ywjpaBvkAm9giUxwsYd/V8AB
L10jF4f/pdicyhk2fiKkk/woy+MmHHLM/aNfur8fGfHQR/Dxvfy4DbggwVabSy/8
7hMIn2IusRyotYCH2CSXvHzSM/XbihAhJEugv602C02PGZloqm/3564eajVsMUmN
uJKtig6QJulewvqi7FMm1CLwax15+NL5ZROJf5AZUqz7VGL2rQJ1PHqA0S0byD3p
/X3d55NgCohExon43R2mLUgZ3pJ+W41KyxXoXAZwBfM=
`protect END_PROTECTED
