`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LTfjQP9uULKCrYMGfZfCFaArgTWvn5+DlykULsgd0uNOpAC7upRy6H+jaLdX2S0D
Xb2z2ICvvUODppKQbHVgHAfnUvt+1x8Dohf7eEeM/fd+DKS4EPVJdl5E8gbC5ZER
JpN4YrU0Zvk7vDa+u2BlYUVDYOZ/E/d2UXIxxWC6JXbr4n/QjPueX6Lke0F4KnlI
5hoHGUEtabL6FmmduvGzKccNM4fD2oLvbobjHRFU1Au85Y0m3t5MHLw9+AQQVzUk
gPnxj1dfaYocX66qJQTZVdqma1ZJN8X/ttHaCFR1lim7q4CMiOZkGaJQDx5LD8XO
BbMvfSmP0bVmQt3rcq3SBUBH4nilj0w2PWTSz+QbVUoNzcO2+thHCYRpeK/7iJnS
LOxChhgZNu64cA3cZiSjvBETPOcBu4K/fpb0wEyQNCY=
`protect END_PROTECTED
