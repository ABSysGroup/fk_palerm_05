`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mjgWYURtNtUc8xHl1Df3ZvhOa218OYZmeVXN/XkJcWJ1mZV5lgJRQFVIu4+7mT9M
gRyW/udVDX81+Ia54mkHnB8Xq8486zYSb8pqu8JG2/1NKsYWit/NtSp2xCRBQRwQ
mJCe0IeXKmvdWu+fjw6fVzYWI82F3kKhAp2uPPgHwOnBloDhMcRyvvPTIqxM/KZd
slUL4392udQGkvZR8jCTYsBEXG55/kKtS3C9JMTWf0lJQg/zWvnL12oqyyEnh6SW
sVODKVjzHIIo9n1a8Yt1UIrXBhLS9LRSv/hK6gyr5H5BcW21omuf2rZ9ukjbAbDo
nQR1si4pedfk88m1baa8nMQrQUPp4qgmlZ6ThscrAm3XPSUdsn6y0mT13Cfr2vVI
bSI8nImpt/1NfVeNylQ/El+XIYgaBsSZIPk+r03apDPxHtCSQpls8pWw2SAXfz7S
2GlCckjri6bBFaLHwMKylrZV/+hj5261iG1XAcslwaUkmvPjOMy0DYdRNzISKyie
E6Lx+rYzOQFZLGMqY1iGGRmlG3Fw6CR9qj1MPp+5j+4=
`protect END_PROTECTED
