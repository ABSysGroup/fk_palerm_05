`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VX5lpSEylzN9hDdgyslMPQuIRio3WOZEpVhE906flbKEIWi8lobeZ8w4+Lb1Vm9b
WZFhPBLWyL47e9wyGACcYJfbBYQPlrPsmJqWlDYPkJ36tC+hB2NSlbj2qLRQAHDU
BdIuBGsLDD062qhOh/cghnC0TvqH0Yujm4veMRPgAtGRzV+eUL17kiHKHxarjUFw
JQKJtPAfE1iaox6XTUsXuAwq8Z9qKQ1esz1nfyG/9Rafjs8pGEAS+XS91/mqd2wy
4z7Zh7laLXWYivaIDDASS0ljgSHbwKCVNuuij8LuW++BMkQJXzEimdsmaCHOaX7t
71Fo6MF0mXIrW7X5FrW9oBEsXj0EC6FLG1GS8FvQK8MNETrikjVLEcMJmO7eU0sZ
/TqmdffNGhnnCNSAH7xcibLFI4qUQ4/J1QDh5LntG9Za4lxsR2hsJdXGZPcDdha1
CQHceJ9NgJ4EnDTtBeqiGxNrTjDY9hsaeZMjA1iogQQGGBQ84d2dqiynxhvtvdCE
`protect END_PROTECTED
