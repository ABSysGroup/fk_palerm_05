`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ns7B+U4Zs3NgVqczw9P/ZZnn4VeKXW9D4K/QZf0VDTZ9n/EJZ2TwAyP2fKC/zR+E
4ymHTbVUVJbBUx2KM3Ajym3EocN++j3qUNfMS4eTMW8eKmzVt0wYjSdPgxkGB7NT
WndtPkqCgHPpQg9gWmYcgHi81RFpAoZNMltypi0L97+EEwAuLpH4yYI7q7scjBOV
EvtQn1EQV8BVW6q1VN9vsjjcE/Pjb+sRMSj9IP1XMV+HqtEq68Pm1zsBBTRr8fmU
VS/JWtMHDaX4msrm9ZhKIRlHwbCyB2Jm+IO2W9A6BskFPVbdAsej/XKj7tjX/h4A
ErJ19nWsO2Az/iYumPN06S6IbRKtOYzQxeOmFKcR46ejcmvIdzByXwiAMDCfDsGu
1Jj1Kdcvw9Bbtn8gLRbOM/Nlo7WUF1ueMUcMu+w+a79CsB/f+PfTQEBRLz2wHAGW
UriPuSNk+Ao0+zSXTQu4DZuTtM13FpFGj3xSIhJt2Sok3s7fSVrZtHYXQhkTxLDf
Eq9tp47BlOepntieQ1CC0VPn+/d6iyamgvpdWmFcAhZjOrKaEtyP7F4QT4i/NbdZ
80DCiEIwBuCKID9TLpsSLOm6fjSn1VZDLoxfGT5HIzeX6nVyjbJetc2ey5qJobpu
I3lVUGQ+nI0WjIOMyYOxTw==
`protect END_PROTECTED
