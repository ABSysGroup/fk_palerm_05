`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7yLw+n0GYi5WnDEWY34G29atZ0bhNZdn4MGUkLPinBauREP4IjHVV8fmife42R78
BWkDJLP+xQNtuDpjQhoLT9RnFLjks76rzMtrxfhn6Vq0NTg7KNRcvSJeSuqsZgef
8PvLcHaWOB3fRnMUjKWo6flFiiA48u0NUA1/3tIjoTvl+Kd5A2fPhdNICoaQW6s1
j9I1QYWj+0vy9fDjnYajc4KCIpaoIHd3cDIEvQQplU21FUhBLhOLWpJtaaKqlxVm
mD4iPqMWlZqXAf4dWo3hWDE66Ndy5JS2g85xN292zQ9uVZaftYUqQ04O9OUSRTjE
TjLe7te47YOUibbq1dmKioZ5aBzdaODft6AitdRJNb3LpKntPd9m1xmkTscq2gqm
OIlW3tHXDi5syzF/eGNy3YEeKt8qAB5LGo9mtwXJ9mHQCEktSVpA+ox2RGhAo3S1
SxeY4tZlkH+Y8JEi70btaXSibgGYsJamsddiJh/2G74slr879ps3C2iEYMWLIo4l
iD6sSWWYgjsi+kLSrUSqf5ncho6yMCShYje/iPDi2JjM83OIExDJ3a3yKp9cui1e
jEfrH9Ise019CPn9egoxMNL3rGFhJzfwIcduA2Kss1RboweqM5LQ1sHnpf6NHlsC
fNrgeEQNPT1ykvjsvZ8o8Q==
`protect END_PROTECTED
