`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ULQQuF9lJ27hIBexKonzHmImp9Huv7tbQ6E+HasTtAfDMAnlztAo6VJpz94nSaWB
l0MP4qNfbqDcUYAVagMPVYVIU0tufO+1JByGmLqsKplL9c7ZDESAsuvHENSmtByF
AGA/wm3kI/zNuQ0lwx8EwQbJFJWYGiMerl7WeydjHUCRRAt4HbOQ/o5DRRzVffYi
wsy7EVECMIuOy6sC1pEvU4GKP79aHQHQLfHeOJXjJ5p/rX/ZnnuIK8800ZTpg07J
FJ41WpxMT05vNjmXan3giKOMOR41NuUpL0j7RALaXEQcmjcrJW5REMqRku8c6hZO
sdUm2CylEjWBIkKs23Ra2mIGHXUEx8jesyQyUcNN6kxXlpJU8zv6ToiTuptxP+PW
btV3p58+rQmNFXvYiTDpHq8W8ym9hO01xKD6uAzj6Ys=
`protect END_PROTECTED
