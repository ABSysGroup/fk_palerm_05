`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MG31BxR9r5Qiso0bL5saHOC/FrMspOxkDMFAC9P93N33jFnayje5lPGY7GZBsI6C
nywFduc8lqL3KwFhTY2f/s0QYC63zvMQZJq73f64UQOlyWc9H1VgHC5XdeBBQlhQ
FiyyfhiSKvCgLlKkKcbjh2Zjv4esMsW93Icjc8BNJhxByHBH5ictjBrKwQ3nK5ne
ENdnEgmHQwjgLLvTz9Duu4vuNG+KQR2TTniZPgnJQerZMU5vzn8rSR5v9RTpFr6f
ptOC4VKFJa9oO9a6La58+khudd9yzPfNWP0+7MSXFujsAX4S56c/VwYvD2Y/qewR
QJjpJV2TkaWB2xQazxklDRCajx6SFLm7Cn5fJMxPMcV6S/VCSq3wzDsmfnY1O4Dm
ZMAClTlR2l1qyTxFXyY3gStkYPJOS/Ob6APrnmjVnwN2zEH3MdMM50TtST/Ij8SM
TEkTfL3EcGSCOFGqVXlIQWCAMgdO0wYjSfD0i9AV/OP1uEsfC/4L2LKvTzZYfk8c
`protect END_PROTECTED
