`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s/zcKXtJOb7uH5xlGBXUA1tdbU/yVQIDeEu4z7sEZq+nhJ1huJLjxrWWg5rSUikR
cNMnsjTj4Ya2YuOYuKsHH6KdCTJntySaiVCx6fNynkxGX8gbPmjR/R+y3IipkjV/
NBxN93CchAVTlxDTjvDJJRROqYS9l1CctqwkbdlKThlg5Squ925tUn2ZjgaCOri8
O9ftv+nALQma3UIq4EC645Bd6BJg9P9DqRV+1hHHMMKF6694PdJnrbMuBzW+HSKg
xx1CnOwwgDZ+gffARtLW40iGuiG0lAn10g89MVX7UjHP6O8eDe4VgXzZdRSrONut
mU/qseoAAjdAdZ4l1z96Pk1Y0Wm8n/ZL9jJixB//8q5TN09tz+AP4ogmge2sSWiw
avu5aTyPXXujb2RGqn1wSNxZiqMB0fWnOjEKzpldbUbfyo+Ug2QT5Ro03bptbzhk
4XAhodKVKkBTMJXfRL79fFUxPPKkUACNIPgTTclAABf2vgawV1mVMqdzRoOI87N9
mkULHqiJqm3cF07PNQ8E7mbv3UIUTk16yH0RXWkA9sRPjGbWGmKWQBMFM3ZU4ErI
L+TKtqBVkJzBf16itxJ/NXciKW+Si2a7lW08HIwFf/PM/1O2GMj0pst+W38WAf42
SeGHLSti33W99t9hVmog83yhfu/WMZ7yBth337lwtxiQEPpke080BU1TbrdJv5s7
`protect END_PROTECTED
