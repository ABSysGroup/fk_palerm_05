`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nG2+MX0CxI1reIyXHZ6bPqmr2P1spjDUJJQv/tUBubWZ7bbz8ACtie5vT22oxMup
oChnP0FA4BWRPBcqtiPi+Y0pJ60DvMSsOndvrNrLRnNNWHscfArS+gQQ9lH80tn9
OCxalFSX4FWvtx4huhVPqy0eQspj7MmUT/EI3Cdovrk2ynp05OfPIltovnJdsuMx
fmCCLud7sklE+qbzMUwu5UEntI7OhOYpECsEe/zeWO9RFXuLt0USFtvjQI95PhF9
HAfeasbfWTDHmcjg/IwxCLarqefkeKf3rmBYiwkGbWlafEMuJU0xNM/njZiqaF1x
MERjyf750ozQL+MJmsi0qxq9OpvQPW9EftT47OMkzqolI2eFXkfy5Z0J9it35bAO
Dxy5bfkbonyWx4P/w7+Ykzb0k9sSklCMqOGgGcaex5W1u7HQ5z1I7HdrDTOl159L
8U7MXWmdRyLntfW2jC9xifARXzkoO2socaOUa5YoAcGN50rPVhfERWy5gQ7/iooY
NVIaTSvEAvMKHRNTZcTUDeshsqXp3c30ffRStJvdSGMu3caKLgz1EP76SzEuqh+Y
VhCGmksbpZIYOITLZETqByWiFip9+isEWKwxe4s2VezVkNvCPWCpbHbP5BGKmF+2
4vCRbx0DMWLHjOu2eWN5qkAY8O4M9SeDNsnufe0hUN0k6MItBLs8oIoUIINbPwEh
U4ph+zfiUYaqfcRgb+lZM2o+N1BYSX2c52c5OwVgnqwoffvWdKaFULXOCdzNw7RC
uN3wJwJcpvrmPpCWaA43WWlo0u4pnR63ZuTzPN9jYbLHkSGqALFSKVSPvZvbKLxi
Wkuu6/pzZD2d/FS/bTvMK5Vew+DyJ8oQ1I0AJDrprTsQ5JxbPSoog8ojui2A01aH
gT37I5jxHznUXkI/MFzLNgDttZVNisUzI/ssg5j4DwH1n7oav7U0s51e8UkEktFU
GchWPIMtxcW0cMZk7HAgZqVezBcxZnGtLexoQ4mLSIkFqwg1wuWsJ35dANhRNEST
VR50zRz3CHV3rfKR0h595nCFraCcls0AtyQIzpOaip89XKS3xv3toziZDSFdXV9+
eso1OXfnPiyatnckd1d1SPDjTZDcM3u2sQ7bzKQg/Nc/yj9iIFpID6wiO3iALHK9
/VCXgpJGK1wLk/8/cLhHZdbTHYWMI9bSnZfPmipzD+02nnpmJbGm1tvcX5PFH7S+
EZ/Z9nWcLV0D2B3VDM/NJAEVc/0DAxS4Xip+aho5TbWcMbF58HfiWBkkfpy15dFy
B/dNmb06l401wFPgL4Wc2eLyjnOh+WOvCRv6LRlaYXbl6L8PMoG17FM43kQCbQsg
AzRtxFcw0EiC3unqopdm5Xs+oxS2miIbfdG3CtUtjutJoSyse85/nyoguJCmoxFV
gqBjLoFzIs4BIaa9+MEGaJ8baZHvrN+f5Dw+3uK7509I/JYHUOl8xK/csQglqYt4
TQ/zw/CwR/6J5EqslhxEIrVdjlZb/vJZnTNaSKzl+tDCwrojNYPZdq1VC/WPjFOD
Ob32YithVOWQ5r3xCq3p7xRLx3Y0fa8z8HyJYLTHfERtGphvCAvU7dvt+oNh0P1q
iKRu7V35Yg4dqEzQS2nrv2K0V/lKGv7QhgznGeuBS59TlMt69dJi5EWgfssuDqzz
z3a6K/twLBKonxh4kXqY5WGo/2cwhgyv75uEz+Zm9izd6BT2OiitQea+GBcprdO2
1+SFTmfturYQi+W7tfLAGdr+Eo7Ph6yblRhMGuS5jGKjCTyNYfKXHiCgLeEGnej8
lhXc5NnfWzn3z9bfHqRS04AEO6XFnlK8ObBV2RWVviSq4gtaaqSFryipqV2rFGPK
1t0q4mEr55APQGYakPLcl4LSCctBltdJJ/+0jz+TRp36OysmW+yUcyAxYhXveC3T
dTSljB44y3mQ4z8zS6TonSB4RLkyEwxnIooPPH1tHHFljKTIWYM2UYpNAWZ+9Kbs
iTe2E1gebJiGRmLJLirK3MSmbaN6R6chIXfHyc7YZfoK9d/zSjxqw+uVgcgOjQPf
FsAcSNOc57z+6LI37Nb2/yNdSSOlCX8zTix245VPlU3xlXh3NO0/K6wh7jfcV2Om
WeETjkblJqyKPV2ORF06Z952pXDwvJd5N2tP4LDZ4WwvA2pJYbh5eImcMet3wO4h
fYfdD8VJQUmXEggoM1FM7UMjAD3l/rDi86zs/mIXheFTr2L7RybsgkNVNdaYAlcz
iYSRX69VPD6/q3qgVgFI0yZY05Jo3PSpvBxny/0TBiaPSzQF8ZFS8Gl7chDDkneb
Y6Yigq7kZVXoQCIzX5SrxgJuftJvfQwLwU7Soa/IX+z4061JAQW0O0AQLIObQ5uG
1AaJQuzcfJQn7/kt0edt3Hu8H2s2JWt8Rpg2Bd/x3/RvTK0i4atqVcAW+9cLDE/5
1ioXn+klVBTl+7OEtoYPoFaDFpTl9Xv+IHwYFwOQeftVCv3Sq77xOPYlkCZ7MalQ
b6gUF/ygUK1wYaOApWgLDEwJ8Q2WFpQB4CP4FkqH5LzOCoD0aZ6o9BN3TlhEQN75
3OfKzLvul9wXlZsS456dFsZ5e3PtuH1qnGQ/3LBZx2XAaqhOXJijiCZ5AuY/9fuL
rp+BDrg2fX2QHzm1muCHm3/GzjirjoGzhEF2ChiU/fJue5UNcjhVMKXloIc5WnX5
ijYVCCe1QCE8SeNdmac5Ejg6XCj9PlFwLqew5ZL16TcOw90bWLNhWMNilq9NKRwL
u858yIuA5cn7LnJxSrZEhpuJtVF2Hnba2bSRrSYn2I9HZMro06MHdBv1RxqTbJbU
teASk8wAomzAxjRujhB0EpU9hW5n4D/ggQkME2D5Jb+YeOLqsLE5GPsISsCwad7v
Ws5OL695y+Vwnvy10p3PR3bRluI4rzYtcHsmqPzsh3kc1kMvDkmOifqcewjmkRPw
M/xbOgKc+8I7tMjdd3Bxw/Y5lXc1kLT5JYJ7d2chucR9Xy+FhdZo4wz/7TFYdT5O
WC8GQ0rbSxKl2qOKQPfa0sTMP8TI+PAqpeiLEE4/E8UixPULKIEpp9hhGiBdVwJy
coYStAPW8XlBU8fKrJ4iZpkn8FjcmDiDSHEunzcn8B8EWkgi0AZtIZ+CmUvLn2YY
j2J38a77kvPiTyqVZ20U65GtJsSCxoN1ih2oJEZTN8qd//94UhUoZXNFXq9dZCTk
hK56XatsKm9e76U46O4OSrSKGKeweAYRUERiktVWOVEHkVszj3SouOEGhM2YzMEo
b0XxHKu3amjVVMAXfeTzPyAICijW69rITfOo6gyfZKgI+vrZgmVJ+P1tiKdkdnpP
fBt6eWjSd7zDOy/zbUTknAyOvfFKcQo/pz5NftTL1ShrKcj/YPPWSbA8owRDO1qM
3GUfA2Jb29ZUKvHXW8ivFGidyuvhbuSV8TUxFeyfgBuIVs56VU1OqMqCwnWYIFcY
ctlcny+APsDbbmyMUO7F2i/TkLywVqzL0Ii1ba03CQ5ZPZqan+Q/qb+mOpAgwesy
tqj6jMdETTLqMNszfIRviOmrPCyY9W8r6NUYHEJB2ebMLa1OPnixRidnw3xOfGxw
0I9JB/JSdLNb7knG4ZSFT92JMVKZibHMyOXQ7I3onyqXW+ihPOro3ClO/uRPl26G
V0nMvgc3CZtHEju5qhw8EYATh8tNKqkTbOMoeSKvEt2mmmMW5Scazka5bJ91ZfR1
mmFY8bkqRmjrnhI0YIE8Phx5pLvU1MwtmIPKyOeaJkV3osoS8GmCB9bp+/Qm94EU
jEuDD9oBfYYSA5EUnGdoXYmFWyn2AvMJSsAwDP+OO1ELkBVjf7SXvdNxETmQWv89
Ia1TyDN3ellxfpe8pLKkANnCRjky6siOBg1twAJzvlxeA+oKu5+DF3jo9f1JEj4N
3WgMUxFrW5VEcKSE7WW5y3C4+h3EVoXs6usX86zZDFP62fHfXnvFvLS+0JpQt1S5
Ypd0N+PE+GAylYD02uB5AeF9KMreRKES9FqxxiXk53rJd9ai3z3Az7anDobo7Do3
BsaTw9jPK8kUFi5NU+NfBI0j31qhV1B05qbvfJu+p/bpzy4uM6TLZi51tGMzmObP
3ymUR0i9Ngu1FdFLpMJdB+RMBC2YaYH3+XSyt0Hf6K+8FxX+rhZnZsq+PrV72K4M
/4QtgenrbZ0ansgoDxIdc8+zPSuyPdx1we526/V/XVefaz2bx7yf4sWebven+6Ly
/jmkJlnKydueIzjfmBZYS7uAuKfD4UjiklPPjDBzYKhWrqgxDA2j5HR6WKsw/fei
fKyZ1Me7RXj5q09YTImPCCYnArkDp7u0dyIz9ALhbKiAPc1MsQ5+sEw/EzQNLLWd
3U/xWDxf/nPSZpr1YzDQ3v/YBKzBas+0y4KnM/5XcR8CZI+1W92dZxiNUIh7t2hz
m4Ne6CgEp4ZsO+RF63WevnaGQcFb38DQbCAX+yfAyuVCwkGRbTASVuQLZOWUYO/F
7rNISFDeFbPY4T/DAOD0Y89vd7SLZFx6o3ag2dhaaU8HmjeBr3dTj7A1bgl5MmBL
HgT+xJdRcWa/Q9Z4bs4z4m53CH9bEhJFEtBrod2T151s2FvtuhEuJ+Dnv1jDGfpS
ao84YGHT1q1LFHwvkwzoeJrD27tfmNa2TQEfvXVpmZnm+TEqK/Wi1t+1kBQBZ9Vz
mv2xHZuHHfs+XotrjR5/5UcDA1qXS75O0L9A8pneI4hj/u84sos449tjRWfOe6Np
5/mSLVu+mlDSIb9vY7LZv/JRtf/jb5hEVHUaSDNTGMOsKjLoKaBSkIIOPaeZ7WZk
2t1Dn3dasDckSWWecXLTMXZpBUcKqX3LjP7vYp3s+klZcylHBOE+w0qEDJubaEgw
2XI2O19jSqX6M/baUSZkLy/Jgtkt8J+z4BDtlZjR6kP/IV32qdgTVa++hS/DP3k3
hB6DZIEgftJ3FgXztsihHMtQhFYI8WJdvyaLMIThse9XwhbcV+3ECx4xUOOnhOfU
jllpMv+E+eTV5qPd4dPF9RkDbmiN9TTzfllazKJxwXjmFW1jo8ESM9/heZEekjAj
SB8jyvNJZosb7wEg4aBzbsFK0wI9iCibjr8WK5+KO/h1BWG5s4fW545q7edwUQk1
v0RQHbij98blCwrGMlBjummLCYYSA8ocQmNv1XNOwGOSiJAoZNow0slUFl+NE0RU
Cqz5x5MG13KvuSH6I2l1sap3h+mxQvpCwP9n2MydyBksOmPiR9eF23nNOuHInokC
IHFNCS/bF+J1iugFc/qcElJLkZdG7l3BcvrEK70vFzwybhyEdZABlc2zr+excFRE
G2+GUZVO8T9xlWcab5BWJMGgF4rUkrUuQgvV96ZnFL/4OLIJ4AcuqcW6KIcbwEY0
nCKa6HvYUzVB1BGVHaAhXCKkZIP+I8adJ52Ur8I4pb6uyuI+VtdrKJYrEmKHqZoM
7BX9HLCqlmd3BrhPXiRvv+R2OaK8E9Gq5OLg8w5rWl8twx7WearA+klTNnruc3tj
US6WZs/pWPjm28pk3t3A0aL+1M2zhLwBy1CVmH4uIU2gWyyfwxlu+/L1PXSvHUBG
AR36Ag7bl4nTETJfm3h6phCpbhwgAE7hHE0IjmcsVcpI4JdO7xnGW4+JDTlrJp3l
PrLYUFhVCcavnwbn7mr458PQ+qxz4MCLosrnq4kd2is8eEGJb7W9hPnGY65pB4xX
9t0cahDY/iADjgQsAjedwMAJBk/bLB3bqR0kfNerH0DAw56bDOhtIKsFt6GOyeMO
mSMtSe/F65ZLjEpRpBUrpyWgOMXyL1TMF30lxn1SZ5Wpgb1cQIN1Ii/2asA5ElmO
1tkKtlr++x+lFexyBqWHyD0q8VmZ86plOY7SWZtKMAbGrO5IYwAOZ6cicR4B2UfE
S7p856VZEc+lgbdfAZLiCTSEkwxL6DxSNa7ua0Hhros=
`protect END_PROTECTED
