`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V/PgZv6dYPX/VQrU/TZHkXxCZOaF8YqVfI8BYAPr0WMV2dou5Eau+2iS4dpW5ufJ
BN2pANDV3DY3smj41efKBet4Y3WtxvOEyR2Y69xk0UwKLXJMVe+L7q7L0UtkZZwX
tDrjNjl5p4LPmtD/zo5KfKIdN2WGuAQ+q7RKYcH5tEBbV3Z3l7HqzMX9iBKShe4r
WTXGoHMS1hDF2pvTXqm4p7/6ihWotJqfWdhqx1QI+AjclrAl5VtgRKH/tm/SFZbc
/8PgBysDdnQq1E5KFUebu4fnv/ncaol7XrstiM31IvwYnzBffG2IWfzF213WMo38
Kk7oRD4vhJKR+QDPUJWTcCjwCULc5Di9Wy3YYnoUPnczZrly7obyqyW+znt+QOMo
8QUKJF2io41pMFjH44tzTC1IqdTxsn9y2IWh0gUHHnW+bJmHs/T0ClYmfZgVe30y
WxYpRCby2qQnNcDygkd/tdNyt00X8+3JFZOQBwK/woQmZtiK/V1mSOsvLzWSMqzX
OKais/jbvZPN3gN+/7JQlsuYRgyOz3CQRq6S+Da7ERwkCZKSsVcVfWQIApjfU+R5
VDuvmGqDpm+DJCo554uR/jzMmyUepHr67imCsjSqYzXWkDfjCOOSvS/uGfGctkFh
`protect END_PROTECTED
