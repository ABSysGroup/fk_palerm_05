`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SsNlb77uV+UGFUYxqg9aIWEqtAl1/wtx1xXCGf3T7NJLORNyj3DNuE9gIOLCuubK
Y16uKUp3sBD8BadxFgPbIzcdW+A2M2qI6OqjqeB9kp/27qofq6h5F2XBOKloARVl
7fVB14kellDXQlC9bZwerq7F8bAsIHdXhZR+OupTHVWjPpo6Uz3p8o8tT5P6lAel
mAmB+vmhhtPLj+H2eYE5Ibl8ev5hQvDk+rloQkGpL8Ye+nWcc5qMEyioB/CF4wPK
uPmuGl2En16t9mfHPeACsQ==
`protect END_PROTECTED
