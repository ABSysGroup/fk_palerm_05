`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D8QRz0zXtwq0oIZc0JojRih0IPMmTSppFdTVW4P3/yG41mOFR6JbDZRAhJe3ALBF
8D9PSqF8+0nDDHqVu76iSt8gAWvER4CnaQV879gUATqeRMKJOaE/ZLVNpFeZ+iei
kbA9dfsI5KklyafYnhHZ06r71tmQHuh++M6iBuhLosT3N0vc6OhCMdh92Sks42nQ
ghvwKw+TfLie76oXULCMA5g9eXAs6supG1wy8qgncP9asHxtC1Cp/j1GMrzc8wOf
TugJkZP94g5tDu1IvRyRxph0RUzUDUSZNhLq3V99kZuW2PxsjBuHodgVnuOZe5nm
7/DBMZLOv2wLQ20WukyHiN4qJ5Y/VhuqwCVpxHrfds0YTqCkmF9wFyqysWX5Qos4
XkndBuWnWjDMYGqtwUU3BSmeFkC8jwCB7D9zCAzuwPm7PbIERaNAq1zlqbGicoN0
A2lHnHniWahjf9kmvi2cnOg87jgUpjRul2mcGnv8kSKfe+f4pO/tU8G+8CrsCa2d
IxG9GwXCci+8kHQjsHn2IQ==
`protect END_PROTECTED
