`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LKv8SjtufFl5gHljCzQNnM+Klhxj9gtg6+FmhZQS2DhRfs6rLUCd5xv2QcNlt509
l0F0Lxl7MfgT2Ni5EyKaenzOPZlnUnK89wjgeUdTHjBs/75pqNKlL7AzYLPvRG14
m+UJc4mWGFlPnVK0eQQu4amsDcfWAJG2T47u8MSv6jy2ORUmmbNu0X60QJP7KlUD
Hn1rGqfN2WLkWwSNAX0ogNJaMi7Q7LTSMz7OOSzfcxEAgbYDdO2xsAdw/lHZSqRv
2OYA71zYYtTPE5PMG03Jssjo2B1kd5r2hBbs1S70tk8pyU3+k4mi2urKIJAsoGmu
MrBhTNpmEVzCd4h0RVjRBVcSHDAjCAZRuw1x482cQQrArOw9YsHyR6vGqqqrpyEb
Y6sVVbJAn3oISmeOSu6STSO0DH6rIYh7/IB+3yylEp9/Ch+8c5wQ06sDYPsBXI66
gMrFBl+X77brz+6Mh+FrSwghnb4L6SpxK36/yHEqX15bY5gF9208G0K3ZFEssOWa
0oaiVPILzhQR0lQQ4jCUDpl/DyrcskhHoNU4TS1IAzrmVXc5xfYX5nTPbHhwgXrD
Ul0gt2P0kpIQekzhYKvCykCh4V7zT21YP/16Zr9JzspfvGIbSgPf4yfUM7OmiZJA
UEHiJocxhH98aEPcMfB4cmw0IID83srFNjLQXR23F7Uwy6a0rud43eE6Rw3umI6h
jUowcBo+VHBJGnGiJ1Mgx3f/QTJliGA48FRtN/a7yJ31Rak9MxVqcfvdjdV0gjqB
/6sjtB7nqRSujfZve3daBnXqbGlLXQi88PheLdMF7V3LdzJsDxPrySWg/rWxwlkX
eZOFOt5ALWLAPbZjFqx7oqxdEN0fw0ecCXXuVKbImz7y3KWYGr6CHKkkNAQ3WZJN
RQh1V54/g+CLBRp9rAGWv19ItmJimyI082Yhi/VvNLJ0iSQpCfKQTV3wBnYc0k/S
BAaDnwm4VJb6nL2PdgDGLVb+QbpM2s2gjv+vxhsumCLs1QXy4Vd00DRsAqnyEWoU
xfKYva3X+X529363njq6Fi/pAKAbI55akf0HL+bv10vKJ4Fxxyq6b4NQsPBFrvFL
TXIs6JizmrTarmVOQrufTClRRS7O/14wBHXF6vyjEl5CHQ7SJVEy2fa+4hdsvPwv
D95tDWOl3FNfiaTBYnCoX9YRTDsU0sKdV6hix2pJr3gHyk39GM3wn0Lo7ycAafk5
0Do2lQdThvKxuLjWkXNtQWTJ0rCOeUL1STOkGCXdN/Wvm40v8S8WNPUxItKlbZ4F
YdUfjrhPPmBKzzuXkX+d4ud+HtaFpVzC0wwtyd6GSpom3SF/azDyOkMFVK8U9Lkf
0Gp5/56rXXQAPMbUEXa2HqaXi/8ulLV1Sd+E4vSUq9BqaKMBU81O8l7Zk/UccdWL
HTLbvBZUrasDHRabXzV/HyjWHBcMwc7zGMBgxltDjxEB4x/lLDOLlmtkwXnjHpnX
cok7nyif8WTAOa0inGM63MU4mzFjYC+bmc5DpFafqm6fPGuK5bYLQirqSTohNzsL
GvexssmDLYtpLehexV/UJuGJxwF1ImM0FdKaClYiuDpTlyld6IOdoT6D3hH14ypz
P9hCifBBzgBqpilBgCiFpHRZCryZ3zC7/Ha9rgnpu7nNOLW45Z7QIvRWhNGVyT64
oyNuVBX9wav2Gp5azm9G+AxA4/3Q2zz4jqjw0d31YVQCikx0Cj21rnwOopaAiIB4
wQxY2/yKiG7QRiYV+URMWUR/W+/BWoz207vMbUVwOoOx4JULqZQJTGYVrdPu3+qT
3aP5z/IgtMKu7f/MwpqVnL/Xay6gTJYiYyO9s9sQaVS/tarA9ZZRfn8/HVBdgi5P
e1hFuXgwKDSdeDXIWnzDvbExpL82MfVp4B8bw1DX5E4L+xpmMYYrNJpAdHMGxZEz
YcTeNruntLp+BFGmM5QkTeNEjKqPj3HOQ6FVhZ+JD57FYKU0v5GzKQeHR59znRdQ
2Kh5QVx8SdcXPzm2VAuLQ6HfLeQO46AHJUv28iaI0IJL9kubOb7lLq/GNuWS3uJU
q1ssqWQCe6PrPKxCf4RwLS8kersK/FFStx9D5ZY3lALGXK9kxkhLkmMXsDWc02eo
/aucN6k9kAFH7NPPHLi+mbOMHfoa2huPsut95KkdG5SEntEGYp9IadRDE/k6npg8
gKOOdFJDtyydNbbQsKyj1rRQkhBcfNDuGn7xmxIRy9b2yJvixV5qlxeZ2sXpXQrg
ntcdmDz3IC7WPYmzv+Y46AWf5nx2ecQMD0cdn6wutu0panCc7SIAnhhHoOdOAQIq
uwnXGOJRxXsQHc3mBfCEZCRQnd8L6uPZJkjpv2E9n0uNCxY8o3c6Vp7d7EWMKdzk
RTCvRsBgf/zU29LHyS+z1batbJxrT3E/9OfWp5+suzc6ABinQ16XQ3Vk4JvfmJ3G
YQCQhhzT3xHiPE/TChGuxNZQbNWNHxh/zKmC8luOXfEtL0QlvRkB6oo8GP0vEmZ+
ZLB879ziPrP4VkBtAUJDGwJQrLIfbLkkflACGE6hI8pn2Uy4Cs8r9hMKj6NpQoFe
R0jKgRItbJswpOE3yBEX0AgT8UezCB0AaIkgKusisQZfhz0AyZDnuWwicmV5RGcC
DkPZKW94dFeWpIcBaN/DRQwmliYb5NS9z8bOtYFrDrV5poFjiwANR5oxXKd1pbV6
XOWkLwESmzh0upAZW5w+lY5jFLBObSdqCH7S0AqqzkP5ByQ5Uliy3rGpz8WLBETj
vowvajqRTV3osv48VtWQWssW3+91ybaqMS9dMl7n6n/F6JGsA3fsA5/p2XEw9UDa
oZm87EnDtVvA1wgGh4bGeDBGRU9NcFp+05o4RXWCn86UOgBHvKmWdWdM3bEALwd1
UH/P5n+mH8qDrW+/CqaijFlH2uWjVb1SNqmC62EcHWcS+SUnKbyug9WRHTvRS+sG
aM1izAvcL8LHtT6d9W7+tlilqCf8zAnZqQ+s7YPTRLmHkETwOERRMQdmFe8sg/Pw
HKk+3cQizqDr5rYcLudL/WFc6OQIPlJPlJCABFpSx/VXDVjzThCwRg+ZifraXoM5
33n36n+4Hcl6QGyBFgQEdAkNkPGmv+uT4EW1KcW7d26T0rKGxK2mUfxJaOnmRAZI
q3EiIX9afFZqq1BQ4syWniNmjaD9B0An5CxC43p+UTv4ywNi9oigO9sMiX8bzuEQ
Y8exU2oQ9wmrtFhtXOHBeRnQtnuWA+JVLcYO4o/VRYS/lHkV0blIhhzc4lKA+UFL
WEhpGQDGmolk9dp5Qe6CVdAOKjPg/ylJHd4Y2YH80UF9wznKy3upBHXpnGTaKg+X
pR+dJ7fEtdy1Z8W4vqeMFENJOap56vPIB+bKKNsEo1ABcS+i5SivesCuXUAvcCmm
v3SlaFV+4/EsTbs7/A9NiuBCScgO8bZ9z97JfhiLFoK0qFJ0rOo0WZv7KSrjWdeR
obpz/jzvT8/YuJ5eHLYx56gXsAKM+O9MGt4IGgN20liO85PlhMk7n013VbyXL0WT
3kuFrbnmd/HShVRo1tHiy1wpB981NzIZhWqSvk7R9zJ20/eT9NatlOYUz8+imZ4q
nIYyX4hU9iR4Nrk4UvNQTVxXBy/b2uF6V0K8Ds84J9N385hDZZO82R0pGNnUecKA
gHdlWqrPYo9TlRy24Fxt8RRktJXNe4SeK5ARHZ+bijiY2/JO3UdzGqzS/ExB2Aqz
w4jx74M1k9HU20Sl1bjgimmdvwE5ek7xumUHl5g9F6TAE1lU8k2S7hISJRDHLfWj
99X1SOZ5Mz8zsJcbN1JATK9NDPy8G2fbdnB7I4NwIUNiMjjsroqTno6M1jxUge5B
vGNc09t3Py2o8hCwAQo/KHXy58Ff3zixOljjA/6QRxSckD5J0i/cuRfnkv3LPtlt
pSLzeOJLC5EsarUXEI9wmT5M+bHP472DybdjARRJxuoSu0DOC+jT9LbVM6kHvXvb
3kKM7VAyEkuk5+AP29mBKeIJL9VwZ/BzYLiq+WAVVPMlwUpa6ntJKx/FhgCABU1F
F2XkubOJ6sOJgBa69J+shKI1T728YS66rTxH2JaX446ipUv4Z7rp3CK33LRyZ5BU
swJljhpCmXgOrRP4sKXWRTmE+OXZBH0xjGq3n9OtydTa6+xTkbb+Mh0ZPP7IpqHC
B9SLY6Il2OmLRwKrpRHaL8VaC8NUFI6ZfCJr1fAyRxAtbykH14MXIQpQYCZsB7A9
vdRewyykvqlP9BEhvRS9P2Qm7vNhqe+ZWYMx6HXMfJ8KedWCfQ7fC2pD1LNgkd2P
zp2T6Z1uPrJaDqeKTWn72ugJCoeTFXn9tmMdN1eCmKmaeaiY3y8ibf1dZkTMr1Ny
1/CMoOm6SACtq2c9u7s5ZWC9YDk7NHEQmaMKaCxOPKUqD7x5QA7dJLTisvXDyjka
vlt+vGQjhOzWGCdDM7EUo01dYcCb0YKR9qh5PwiGq9And56QktEXm4bIzKMtQTsC
UzTzzypO2yWJxVzZT4HX5TXns6mLXrTQO/OcgXevb46G0Ljw68sH2+ocsXBYTJZC
9K+ejX3pJL3y+wff71w2MosRaSJ6nWHGPntqsG+k04hZgFlDcTDKMCbgiNSK+7Cj
bIngxr6pVzvycaeQoh4CP7hzYNXHvfdw6+PzwI4QAb5upka8m56y5kiOdx6DAgpd
nIKU7lG+EXEojy7a3m06p/jtprK6imZyMgIts4QHoEkBjJ5i0P1ROi3h3ace7K5R
g85xK8/tsRft9A/D9BhO6W5MeyP9OF+Dfpy/vKAXoR3WKuFWkhaoFaA+7tK74MaS
nALhuJVCWuUHpoTWHvJ8hpu4W6ZcpDcc17rAT2ZGxy2atkqEZL1AlBzcBXlFnIOP
jHLXP+MT3OFBdZ/FJV6TGg4V1bqI4Y95PjaNgkE7/v4ynJIdZdlbr6u0yvHCsqMk
oKLRN/S9QCVHCbR/pmSH5uFYFF0Krc3/92rNAPzp4VGgk0q105aToehZch8nX+fD
PIos0Zs6kKVtgCTOAPZbZ+NEZrPw5QidAMLz74Pxyyvc54/UwGAtv3eBUsjkAC36
8n8hDa2J6ri4dPAj1udtyQERpLGJyQth/Y7ORpYs6mpTS8yWj5Vc3QCrXY7Uolg6
18flokBxU8xaBWaXjCkv7vpR+TFMeV5HW7XAUDF3qn3WEggxRosHWJP2tDBkEtH2
nljA+9z3T9XkiTBoPgdFyNtPQBuGrb6SZGcSJhZEjOoSdmnWubX7B1YG3dQQzrjV
B/+rS6diMIAHHsa4+1Co+gA43YM+8r+N5Vb4otagCF3AMse+pmOtVHgQjCFfXsKq
0ejvpK3fhCrryNP1buoEsMeGOQwVYBergDKprh2SmvH6Je3mWHCqAvcKoB7pkTaX
MOiMSnPvUpdTkwup6fcDIRyUdj2LBIgpZETKeXQOFWGdhrDgafbq2/Ptrx/zf/pN
VXg6fPdYVRwD8V6+bn6LAag5diveg0E/eS9iS2pR8b8gnHYS3r5vFyH/8AtNqeNn
qfknDnVjtBAk4ohyilAq0Je19Eowbw/w4QILxG2Iw8nIUGHhZKD9Hsazj6oDCcmQ
XFFPm8Q3JyvQioeCuFPQYVwZZsKTIxekalWA7bmWaWNtMbwL78JFbKBdoLM30V1U
Hc5GWDTBnf8Zi13ci2r82vzU38HJeqfesgM15laLUrzDL/PccDpxES3eEdKSsoa7
KEcJvQGPDWNa8egLsC+T7B/hGz7uUZIZ6sZzptCs05j0wDjwWk3TiefKP68peDgN
gMoeD3IfEiIb5Ns+zR7kxBOFKC1/hKfSnUChxPFTS2P/sosrl90Rk/1TXvdoTpo4
YP84C3HVa+c9xxCLJSA3HLnQrco5hcIKaCIKEbQvnH/Fy3fpjBNlPTfBNX3uNjG5
LCfHSr0ZDj3HMNtKfRT+LvBeCtMgrBNtIsj+gGWwEq4xRHZDAoD45/AIMLbDiOD9
55P3zY4vfA47cBplzbVp26ncNsvQ+Hleu4NU5T6/kG8ZxRiv1GXwFDZ8RYtWbJGa
Nota8+0It99LdOKFdSaHkKs2BKd5pvUpghNQOYcGfPqw6O/TQDHvJfGTnNbOmaml
GSvJ4tr+6hmeRqwMmjacwYc/UTcDFX60PFU6BgjcKnAWEF1M/046wTeStJdDLrXr
TfBMfEtYVmq8uQ8oZ0cidDUjHgh2HDkL2PG+WqFHmyNy/m0L7dRWc0LlUAgLVLXw
5K1p+F083WC/DgDbFnP2Uh6r1qxDzuefPd+PJEJIhEqpoHcr5C2Qus/lUQ1T/9yo
1JC7aur9joKPH131UCIIwXcNIidqx461MIPnf/g2u0kRL9RxUTdG+jTVRj9iHQWZ
QCMNLdv5DAeTfbTfRvY78lGha+DO/YyvvqlOXm8MmSjqYgYEN9bDy1K4Yy+IWrHG
DpFnfcFyAB1Oy3KcXC81kCki6JsqhP6wB12PnrouSOnuNtnWQiMSQUqeA6rSAxJp
fOcbTColvqIiGWsWX4Cuz7rNhjU08zXBefPfp3g/HMqQHAz/NXLO5XXTPNd4AJgQ
SIXDB4IQ6Xb4MzGZDPGmzYBL3jF963VTXL/O1VohXD/aQb7VI0wzs7DEPyx/Iwi9
pngRVsAB+Dz9k9bWIPr/K3cR/xBicd9LfuzkAXoOdyUGJcaqLzOAhKp1bHids35a
betMRu2Gpw30YZhGe8NrHCzBVT5x3u+4oxmjENcsbPh4QX1Th4IE9xgNEhI95sti
SzVG+BziTu7iR+fRKIEsemrXAA2mqq61b288sBbGnoEwUKKY0ke4Kf8VDp3wcFxy
4HpbsZ3YUqpJDhKZ/pZoXDDEqT3jqizqTkhAWIPwZLm+nE6o1Z1KuEO6MZgW+j4Q
2kHjaLReAx9tR2awGsCWwtz20j50trFHgkY5swrEl86utjKlAvfp5wYu3LOhc2AJ
QY/NDflsMGd/Vshz70EPyDbUU1fS9+WRMubI7BJO6KOicwfGh5uf3IObOM7QvFjE
MuXzXQ3UxyJWQbBu84chTF8wXUq9ygOmQUbskzGrcW27gcxMM4/eWExC+Vr44Uap
NbIMUVkcPdQbrLnsMmYyruFListqUJs8d94QXTHBZPQnZw9YfGYmBrRcHxU9sR22
QQDmQKAR+RjBXGU8SgGsOrIQO3GHoAdartmFFN/jEQcMIbxIxKoukeragzNPXOEm
NUCxbK5KR+FYRGlOJ0E2Z9Pi7iKfG0/5IVsOWuq99QLYz8+ReXH4TBplQuBGNQUg
eDl4fnrfFYbLi3InzEI7epib8QuvXpybRoTKWjvle1b8U1DThqB+fhiOn+YE3VYj
cZD1LgCpb8/srVYGRkvdgqONAuj/XVOW3BZrpISfBiCYvF5eZGxwVyetWTJzhKzN
RDQR2ZJmyXjPNp5+lJcI987zoiqCv++rN3oBD/jINpylOY3HJLe1i0TybRhnLuRT
j+o9Se6tH547z0djuAWN3ruD3azjocfLUPacyKo6jAIXz2XotL+AofHyaDY9qRxH
xcwr33YcRAYI4oe3XzVGcjZc1Hs+FKfSBg4YvfAFqAl8cowUq3L9UAED8eGFHus2
5uE2Ii9AX0PbjbqD22EpeFENFOd3Ek+zLqwQdr2YZpsiuMd68R8UVopSvlzA+NPC
nVsrHUuF9B+SygjmKMnBKgnKGLPX4N8NouVpncDwfVxjoskQ6pvzCcii1wRD/2SP
AJJVeTYkxGjCtK49RAH+Ny21fWMpRiDUJF7HsE9mVVW+VU+cApdPcCltX3oTyu+9
by5EomcsAn8n2c4Fgztej5ctQspkYl0Wt2I7MgtKqo9PA4Vq4RnehO3QaDUgzOdR
n/+SCpd9QI2JdVJglW3mcHrc2Jq4vSSNYLznyt+zLnnW8OU/1jXK4yDSQd3cyUvL
wQch+1C6DscFTGegvJqJpuqPVA74vga5pfGc0Cc8gu+/oEdE64HJckeGKhOYbB90
jULx+BBydjQpKzAzOyYynZ+qWjPd01Eh6cpD75nkEG3U/2zDI2oZ1DqH/QmMpNRv
kV4Ra+hJsDCAD6h19mAw1JFFC6/6b5pwHE5q5XnnXDmARmLE2FV7qKAIp+1aXtHp
fUJh2rUSwOelFMGVyYtJcfkQ0JM/0+zda6inf1FEY8Kx49Px7wJhmqpV+n04mCVc
+CJNDYJgDhYRGwd4c2w278C7OXu01M5cs8qVSQUpAsm1gIiAJS1plusYxZGZG/xH
70kRgJEqUWKIUdCCCjUMDBYoMhghIxOY2LYMGnP/w6Mb1RoArfAhayiTO5sWUavg
2CiiPaRSTw67zB7YfT5/4G7QZO+MPVao7YHTcFcmD22N4HQtZVG/Y59K0wqpF5CS
P37R6BuJ6IhILIK95EVRnhGgrDflB20jSio6aedlfRDNc6rX6gcOClV83/H/lNC5
EESzaISWXk9VtqDggHRnzLhMjwkp/kWBnWDp9o0YmZOlocm2FR0pzy4CnxcFu7V3
y20NoxT0vs5bGlw458yuCHTqrtg/BXbvVVyVrmr6+uJkkMA7Q2c0Vz7eeb7d5c/m
TXDwfUGwlZyJIII7yDhG+pd58Nf3Nxa1b/OWB8UE3gRvqzH8nXwOufW55oMtawKf
MRx21hbuzlvbGyqRK+mDV4W9KOToQkY8IqOKMEoQNznM7YTNUUmSsZGORT/3FrjG
ZvOg8nh+uuAZAhb0ftT0WVwTs6b2bc2xNSWuVYduzSYQp+P5wfrijx3QNzFfEl14
QNEHJtkKx9GqoZnqXxHUGSuo4BMYyadR72EOkP5s7vAj8/aG84On/OjzGQJQv4KV
lxwo5tIOC3mzCP6qOmX3qYJNJ/kFP4oZDGDp9z+sTSTCwPzGaGNc6SdWPjP7C1Sf
yDlRdrVc931yBOU5QkO/lpBS1CaDyAw0y7jVIERqfrLOE4IWQ54LPOvh3p3GOdks
m5/j07RJe20a6HgGug2gAoyN7A/mUUxiElgcQxYLHKurfSMpoaaF5Nby7lf5Bbu4
YrC2uxd4r5wy6nC54UWxJitXq+/LzJcH2r6V//NMghYSRP3Vd1u6q/zimE2GAtZc
ZXaLvVS71pQkX7WTKSNaz2lJmavVZX9LxtQ0ICOgeP0E3pICWyQqHbs+tq1VZjz7
fePx9/dcbznkJ/HIOEcvGdj+ZBZzgj0WZbSEJhk+ZMTnsa6PoIflFZn0LyVjVlCn
3ZyAMHoid4ANBYs9qeEXd7g+pRP/7+r5YT1Lh97pkVS0wIWWaQl+Ka60kkSpULNZ
yGzy0iYIyEn0hdtNk4x6073DAkMkE8ru9vcFcOShicJ/NYk0XmpZMjUks9oLFqd+
XJMnXfbGVgS+GBNoQU2J2x/AgsOi698tFRaHvc5LBkqMWymJsxK8AZdJxDOf+jUb
dqM9NIVPrnEl3IcjZkY/wYf9vwiaGhohEwISiLPCULKX3MmrHu04NEBMXo+Oku5j
KdcjiLm5nv1+z9zpHQ5oH8/4e0Y+ot+zjNrPq2O+8m4tAccm03Jw5AHMe0vanS11
gcnCaIbqpvo/Y0Ig9uXbDfOThGYVA/w43yFXcASJXjYV1RiKhkK+BDc7irGcZTQs
oysnN9Jrppmc34E1mfm2ObHBYpqM+L7+BjW66+ad0AwzTuJ0TnR/7+TVvIYK8k94
5NQoZ31u1ayU1xjYzIDCY/BiCbbDLatkCz5n3ur3QSvhe2tq9TdC7Zp/ml9xy4wB
/RidJZhlCdwSzdrpuqCI104TfK/YPe25eq5v77/1Ka//xFcuXx5x5E6vWkvT+K6I
JaMHZdCVesnOWyYLu0DrGFdosU8g3HTZhYOzMfl/QINA88eXfY79QEm47aYwhQQ9
J2Gg47zIKs4ihRD8xjOaR5vZwUWzgAn7Ei3PHP2zEXrVi0yI4OkFQyWZNWRhrpHx
ZGsgjdhck+WHDC10oVDA3RTCnHwxVwI1p+ur1TaWlJo9p6BHquaFfjf4ptVpoKLZ
MtbC3XPX4pBKuqfdvxwbzQtnmk7fhRmgXHyKtNJKd2nSt4aDCqyRI17bJSXJGNbR
6TF/rucnBsHcTlPcN3UIE5vjPW0EPjTIYVFafmGklj+b3nRp57pS0bdWIRfF8nvz
ivEJp1ZqLMTqumq/K8hZdae3ziIdPlo1zFnkQ+zztpV+3ystHtBv1kAnAgBZs7to
IacZjZexGTKT9JSN0evs55LBSrIT8zOmFwHndzTz+4aZrgOD1/7Wz0VtoGk08rZy
+JShfQUns1Z1nVTlecGHPG/HwXaJ74VSsniKmQXZnBGlpSAq1gHG/ICVY2m+VF8h
c+vj08v847BFw6uPgNWXARFEAsFvMLYLC6eLh4NgBK73dZTbMUrKG4xnqEVEJXux
ev/v7tA3icyx71h3SKl0Cui3qLxUJq38aBn6Lqiq7MFZ/pvcP4L7ltAlddR7Svye
eQ7kbCkQdaAk53wAMRFvNAt0Ko6YsYdCXmRl8cvMNXJEJMO6/C+HNL4URZP1ID65
Pd0Q7S/wlVnXYZL1czUOYBlqFLYrKS4E4I2EObXcDShB6MNgiWGcAmLe94sPIqd8
aj5Rgap4avcG16K4eNRksiU2OFqWrd+nNSWQvTnxCPH90l9BxRHQKK8rOyOQx0LR
a2vhBd0WrfeyeQ8kffohNamqKUHk2833BW1+KKvVanNwZWsPO1C3vs5b4OVwyeFA
Sy6IPw4wTbR9TC5hyuOaoorX00HuCd2/JNQxmgivcbqFLqjS/vxuqgb2QjQJV6T1
4Tf8in5YFNjR/9mYCD73RUTgxa1GQXsIGjEHvVI3UxyGSstJNfbSrNgDW8ZEKTej
Pz/kh9L/M3BsS2YWRsF9G30vIG1f+uD16hLWuzwUF/NDHvg3RS+zTVhXfN4sWdCH
rMdHAgYe7dQPCJgwbZWmp/9nVgICaTckoBkaRtEhnqz31OzvDK5UL1Qq4qZIctdU
oGJRKmJmkG8HO/VCPITIhhDURnnh8AzpNeVn654B9wqhaDQTFT0e1nh1MjH7Ienu
Vl6rbHNECfoYu5Azbu1B9LTm28CT+1bWHA/Pxdvzb3DSDAS3qwksXEZlC1s4xqpz
eAy2RpoNaKEZGJk2TwV1r9CXYF3FHNvWKUV97MjtsgGhQB0DEGEGStWDByFPMDfw
++G6Jem09ZYf1JLT3U0letW4e9KAvvTVwxaAd3rmRYRewsqP1f4hUm6hFdAI5UQj
mMkvnGGE7dBeI5z/aZr1VxgY+chz662R7CvW70w62Y+8SYPy6RqADX6Nguz8vmx5
gzmG2N8OamKGZZJVokodYj3ayKIV2VWNF+i3/CgQqI3/0wtKx5yxspxS74E6V59w
UE5ioYksYvZpyVwzScASgl6d0k2hIyQtROqQVhwupjm/qclfKySuN7O3ZfBDb+O1
mUgVYo4NeZJi2LQMwuF3BQxkOGQ6OWhYSppoykXgNSpbOpaSHRFwv7/XV+zmr6Rl
82+QMKBA12Sg2sqjKsJJcsgdXDp6w41MrLDN2gprDwCbnBE0X6G/k1zCTX+RYNZ3
wFfUKiBb6Kv1bSPNyEvwEKDrD9JRLQk5tNTMMk7iWjaeA5faUYoWzR7wYOezkIs0
CaPnDbOxpjcFElY4fkB1iB+e+7/wpklpf1e4gT3wekloQUnKUuNwqHklTy4I21/y
NM7lvEwpy4QwxvO9ExXQpyGKiN4r7LvMUD5hyRPWIh0jKIV3Hasnq5aQfSOQc9Z4
jzcYGkOey8fgvk7gqcqlKe9pYqrce5sblesZfaTVAedhpeW0jJCSglr8zzI5d0r9
DtZbfiXvu2cVuTtJQr5PvdjSLG/mocV8bgYdsXbV9e50jq7OMjzlRNkGsoTSb9BA
bENIAbHPMHxRH6ovc3/V1PztkTqqYaP5Si+XAYpTu7pnuExF0T0yEr5Ptvr08yna
1vKOhW0wtigckamRCRVb2zDs58/h0wkbSJFJT5j+esvjYYjLV52KwE12pOD579vF
VAEoHsGeGTuJcjn+ZU5gbzuqpfocyUmQqjsDF05B+EyEfbLHumh14VtdXPIxl9xN
0B59RlSXcAEzMAXWHUkWbldnwZYhbpil5y9OYZUL4Eu9XDfiRdkMuiGI3E2JmuUt
WzxwKc1xNC4tRszcHBmyn9C3ZaGZ8gB4OgODace2HjdsU8GNmW1dvBBRQyZPLXWM
4wW81aNzuTVng8vyNRN8h2IqqhyNVpyJ3bD5F87F1lV972l8oMrnUP9Xh0ROKZeu
Dk8oealDXaydR1J9RqIgU5HGeiSSClM9Qb0kiS+8nW88IdUUBRWhfNPq+pHbUGA+
KCNBFeJydGMNERrnVXAJVVM6+VaZ5w16xZPwj+CNB0en9oZGfQ2p3ERuDIPdKMTi
wIXjDBTRqMS4XEeB22QKBYT0FLMWn7Y8K6XisKYq4w/Z6QUjUK+D4hEnbXXK7yv1
Xq4owEBkSJkLWf+oh6+7Z6VE5s33QpdKyjki12pTe9wt+PQsRlXlccrIn4Bb0fY4
Xlg5dBu8HGUJVrXIZh+3c9whJPQQlYA01UuHa7y6RemsrKRiRDqrf1WQJQsfoeCO
TT2ApGXR2DCarIWWxop0ws7aNySd0PY3kfWrcTw0rxAZmiUCU4TOfa/5L2rR6Q9J
ZCQPqBmts7E6IY/Ka/CU9dcTh4fUegMNV26Q5tD+jFuZFQUtA0RJHWN7Jpvh6tYK
4LhoVO91GLlXhfnMTqIEoN0kGip5DhsU5Z5t+UnULZ0rGlPfSHGje6ErrYa2tzYy
J+zPU4fkXNzEhDYBCACD0tJDuUPESnK06TlPDd65NvhVRLozqAXQJ+WGS0RIcVeo
UWKXjzD3EOLKIYJc1l4Jsw2kiO3U9VqaEbtDKT7PjTWBX+lMNytfGN8v/4unvfkU
4ysX7IOubbtpX+ztjjOHri9Y8iShtmkS53YvDBmw0lgxLz/4jYEJ0ECf7hfo4cok
FDNdDB/WOFT9Cdf4t0Ba13Vs+Q/FmR07uXeBbZkdcDt9S6pKb0A4Tx7yqrDCGoLw
RCKDnEjiQm+q9qfMyCizCTi2MI6GBleJXAVmHL51bNLE1wj4DUQ9lMYfvtuwFSkX
LZPHPwSB6GoQrDEql0WjLkiPQgFo04pDwzVYotDn7o49p2mXrTBIIqs8+qYnrChu
Y9aGcjPJVCHqO5H6SoCsMSj4tc/lMBsM7UiQrlsmDXyLxOw1zuwrxIlg1DxwcLp2
xea96pXgb5f42Bl2KLzLr+vXFwWhEn9aCygfg1gliCzaim1oJHrnUYyyEsEUvLzs
HggX/3uqQVfRTrt8IND25uchxLhtSJgg8Nhja/q4I99MUT//W/QRfrx/y2clPJz2
aZ49wvyTjYXFJDvsIVaJ3sqJHKE10AmZR1/+9I1cQOVsYakEVqHYrlC4yLzLpZtZ
UZR032NYQdrBuP2xi9FUC0tk1I0nfvxTkDWrq/c+TLzu29RksroRudVinqttMcMc
AcqDJUVKwAsWHVYKtjmuwhM/wkdsx+9DPZDyzC5NvHARBJEG5PJvNUsLAUZ0t3FU
uxQHjrctfgvzUi+SABMYtx6VdUg5vTMmSlyRluIB8dDxAMv/iE3F1WpSScQxi+dE
5tI0AS3XGz4XRw3o+Vupw73B8470CxUqMLVCm/MN2HSvp9+EqJPscfqwU5Kz2fQA
4zXIiG874JdbPwlHaP1AJVmt9PBOfsvPMpefhh8FFIBX0wUKDF5CMquifb2OaPw2
4dzb5R1yanjV4RX8AOLf82BvBwYqXjauEQbwo4RtplwnWJgdsEIKojBTmWjedlkm
WLvV4EKTH+W3gOJis9Cj25WLaKLfaYKjP2K3LpuGhQLRRJ8L0FyainM3gI41jjB7
bAc74S/rJVxulxTqTwztnMtDVoRwrCQkcEwMlc4wD/WmMLwkVey2AgT5J58u+oKW
UeL7xwmnE9huzeD9QPnBexJFHHiOpMApr5b3AfAbT05z32jCAAiw4y7v6DFZ54Rh
5pXnKzl1j/b9wOIrkrzlywd/JuR+7gUp4Msvb+JcHYqgsYtH4d06jKQq+VCV7Khq
yR/1OMGvCYpHTf+g49Np2cBxtRJSf4ekqj5TA01WAHAjQDE1MYy7oHK9oZz5nGNj
QpebEIn3ekUSJVgGdbDGgJd+PNTjPIJ8RhNfGzLg9u8TM42zHPdPz68tlp9Zvx8S
gzmw2X5S7H0OcOGg4yGDzgK/0EnfPGB3bk0q0JEdUD+WaBPSJh0ItA6kDVbEeT3I
bTVNr3K2H6cyg2rJnBeWNQX/8EA8FCZrn6xxcRRQHmKaJNbqqPLdlkhe5/+Qb8r1
YdpaoxxFZX/ljuMPXBfoH93yw8Sujul39Q1YVTJDQQ6bvlMVd9V2v9RwuH8y/Mvp
2AY0I34MlkMTqn6Rb6+sH1yk7W48yrrnYPGdhM9yJ3LbgmnGb3p+w3j+15WT3/mM
Y0maWeTDrcxnWnAGjBtlceSOkzfNFzKQNfIVqh3sZc8AhRVP35Q4MfVrvdWk1aHZ
NoV24pPkDQctFcUR9Al+QACzpo1+2KxGm8FzQ+lwoGfG/qvX/eScFYmfulm4jPZO
UFDyZtA+DzjGR2wXDmdgfESTHHaJ4rvCknWD0aS4Rm84PukdR+olSRaVPBeyAgVg
1XhrM6zO8mybQQqfhCUBke0dLMIxVghql/QHO1yVf7sXrJfHJAbAOJc/c49gHDi9
YkP/EiOsEoWdkTf4N5NPafE8vh8qZ0AaqZjzeC7xUN3yvM30rbw7LCmKfk0qpCtD
/XQzBWBp38y0ZfQADDerMVchRooY+1jtK7sHp/WX5aNx5xA31/KC5c9czOLf+LiZ
f10l/CskPtEkqhJgTQyxSwF0aG4w6NmrvTWTtpGu/2SDExJB9HCEo85BPDT0qufT
ASl4u7fGSXIhuLzw+A7DUszhkhk5XQtZwJLJf5fakTU1RHd3wLFkNiWyeFsjL7Df
jqAaptXxQzX4wAwW2ivHDNKx/Tg1bGZN+lb9IjSwstUKLY4btP+vJYvg1sHg0Jdx
lQalnS2tGC1kwH45YNn7SsCnvUJYXRWc6dvdzPSNksuhVRNoxCIyhUhBJvQpRmPS
3AIDgSean5Sq+0ZGu9e1UPc55tgvRd7OHLrwZvJxd6MrhhuFmZxVAHoc+bcPXk+y
TS521n4xdmnZJUMl65bCvkAmHBwoYQGtsykonLjIXAHQow3i+e0LWfQMwoNLZAt2
UzmZT8M3aIriP2MAollsoQFg0sORwFpWMQSN9JJiawEFs1fj1acObQZh6MKGjsKK
4QQjic88JjfwZakH4+jjmu8cyBSjWyX8edOEWwfNa4v2Lup1kHC+PDyozLvCR0qp
kNTW8bS0Lc1UOxISx9NUfF4LGzs1kMXgZ2zWNjUxzJrMgrveZq7fXRP6skrUC6+e
BTU/z6glMU15l+YK2s3U6srmOOOlNcIR7Sm9PuZpZ//rzoFXVcU3NMs5YQwkNwsk
W25rsm+dPqu0hC8rNluoAgE+5auK9wrT4yXGoOESvlg6qhX5qiqU3PSI2LGDZumK
I0sH1MIhKGR9PGaNl4nl0/BqtA0LLParKWH3Y0jpV9ugITSfh4eOs0DDPnm1VVoX
z9DnkAbcGijLzHupDeydMdgx636C9+q6fMBFuj1Bdz6dj5XxFvqkTkSbghSXkTLa
JGqYgLiU0W5jvPb0vRnv1plAgAcahtPQEn8gJ7RZQyuJxU5KSxYHY6fMMvAeKCiA
qC89FqGEaaGCFNB6tOdEiLIWAm6KknOH9UCG7RdR62OO+WiIIYueg48NFktBm5jz
ZgmHyISzpMKKxbS9uAnISz7JdlKa/iWILmKePuGCvR52GbgTJ8bJCHnN8V+Ki+zL
koR3l9GYTzn4pAhfLCltRqjXwqqbq7V2B2+zoLKZ7yEzWbl6JJHXNi+k0TmKnG7s
/1c55Q8yjhlN8TsryzlxjqefYDY6OGs7EmoRHfFoNE8kOWKbmDsPd+ISRKjeJIRx
bxS8Hw4LJIxgX9gsb6f1buw2Xl9kYZd06H5MOcD/sq0KyhgjdXej5d2jQ06lZWKa
xyE7V9M/Te+q79z8B/eNgHAUo6vNAFuaMpg/yXZU6yn6vs0BZJhbr2oG4qfBBAy9
mkwo8vfrDtGn80J8WaaRNNELkq6eWKNEEl4XeAE02rhvOXloeaAyNZ6dggJRr0Lc
99zb+eJykTy48QIZW8hyIj4aIH1YPObtHNykr5rxWYMZSKXXzpknAJHmFc8XlhIh
fwMSoE8Xd9hmn2VXm94o9H2HJH/Ch5/aMq9fObJsGL/ixk68tLOk65DCDqfZbY6U
2zgTGfBfqiifoLchBQcrz/YgAPjBhu7dZIkFmNc7xmJKk18xLFKFP4obedOKC5VN
6i8OUCtWDrMoHscweGlg+clo34oykMp3B5W7sIWjNn+JjfbPn/bCJcLZ/GcOrsXF
e22UOQZzlBT/AOmrwszbk3axsTDuhlpAUnvZZchUUpLQk2JBH1gpP8q+bKhvfwBH
OQidRBlTAN+mrFVRYCmH6Yn1VeawU8sjJHJ6emINoT/jfhM/786a5ivwT6Bak0Yl
53KY1c6LhISfMu93NLIcP+1XfxkJziz4IzqiabT4dvnpsxLDFBlw8sDRfi/ETKBn
81ivJQjjzaZE+xlzsPP9xTJuzO+mS7KzHA26brnAfRP9wYYaLj9dp7M7I2PqacN6
szPuEzvH50MV3v2B3+jadVXVsAfJjGE1r5beksr1rbxPpbRR7RvJDuQ2fp2xGQVH
f1kuciAmii1MpVaU+4wzIC8QSq5luP5HkLB9/VdQfAhK0OXkwyi40EHRbr41vxh2
ooIWPYB7AT2rzpBTOG9msiQDC7Pxgk3g14GLML0/Nv0Rf3EU0G0N2ERiv2Id9Vv0
E7/cZsGxDhqlwLvPzrt4td/l2i1eDwh6gQRMBi9LK9RGm7mDfCLedrQeYd8QXI9G
o09lje3b+cIMr+rleNoFXrA1rnNjmxiukKIga+Dj0sawIt6bHQr+qYmWltgDD3wo
BjbIjIXayRM1Rq942GF8dLWSBH864QvXXa4tM94BI97Eel1NRSNAnt1ul5ntCuO6
nOIOhi+aYcT8Ij15sSbojeVJ/naFa+7hT+evWOOvVvI9TIWyG+13xh9c+CYV/tZY
pAdzBuFKSEttUrFjCVgK3ejS3qlPIPij9+iIO+z4Z3lLVSkevno+y4JZKUwhezDO
7f0SmfKbm6XeCaNWBriyGGTFEKwTYyzvW9MVsq4DleM6ntJRJ3OQUIQaqU3eDymM
OwQXToQD8p9aAflPF0/5mj3nFJKvSFNWJ8EqZH3ELmt7H6koOEvv17LDb+cVEH5F
Wc+uKXOWWk07668t6+ZFp5yOOs/xdUeAJ7SPKC3/xwurHPSAfx6gDTiWB5L2V3Ng
3U8axPnEEp6aeCup9ScE+/03P2M/wW9vtR6BW1Kd5KSO6bW/hU5NO4/c/62PstUr
8Shoq2E+Ku9uuiLvx6+eQ0M3fabs29ZUpRcCrqx/nTJDghAk7IkEnTNDuO1Z+PHY
+9RIUzAnwYPQU5DEAITbow/5j8D9WdwVmt3JjhTrolOO1Pfq0t52r+mA1oCpu+Fe
xy/sfcujc4DfKkZ6/dCraB0ZFmLF0VDUoiDKD/Xbk8kUjju0H1naWh6hFRyvoX45
BlG0W3OgM1FQZmp5eizyXzka4pLb+6LC2pJIce609/w0Fo5el9du45ood1ytjnb/
GSjpsQ/ivU9JWg6y9YuKaKbpVL5Ge145AGjWVDmAfH47+/G+HJzC3yicS83LES01
qV7r7mZ2kPef5u9bUytwVwFNuROLCYctEW5kqGv5EZaoFuXpFBs91RE0kbNrrHkv
KYhOLwshvEbJURj7ff3lxm1ywfXu//mEBiU9YnvzFKnmMcQ4nC96rfAZHi5zd6j6
WXmvHYleGcbwKem1YfcQPO1alaGlbYbycp0pvEwzaJoa7PSxgtWMaMPC4ER2KLxd
fR/xtxTpAxbpIHNfqxHmUlWHDc0eNpWo6JdKbs0BAldY5S4qRaGiHwvLcjVxlFmZ
yqWMphViXJ39EUPmIAT/53zk6TXMFutA0LTDpTXloS7mlqOHk/YVXpz++bhyXats
NDpKDSUWl4xD9LvVpKN7UwwchGXr5oquFmIpvcyfzoCR3yPpHVcLjTzPZluheSUz
Qo8VNu5dpOfmdUbgm1YfHQJHSx8pj/4MJBpo2Ly3luUR1rGWFMdvSmMQsbgt2bPp
jFfXKX6UPYED3fO+Ee+NywTUFuKKlm3mwa73bgH/nYXgWjtc6gt4JHvKZOnMn4WE
Cz6BppDQ2vjt+CjYEgwUlJUUeAaKtHsGI6AfdAturUyNLaHV2foyN7FVBQijcWYI
r7jTX0Sl45eYO8ZsqyfY7G63Muz0R5TIRsy9HMeRxnC/4+X8WG0FinUUq6oZzflS
fGtaKx0+SF2B53ybfG4rK9ZeFPrOG2VhmbudzOYhakM+TpOIphCazcWFFVf6KVMf
ggfSOQ11UfzhWheCvCYvqNzcr6eDjh8qDgJNLXXEBdwmaySRFZTy/A6f51ntJ2Se
nQsKzVBBPcpxQZJydSZbJgdY0eD8RMJhqXy9EnWPWGJLYxw9mMEFqnfbh7wK4bW6
rYwk2D5E+E7D88wA8fgpF2gm3wkUDMobk4vxgf1+hNhFU0hj54Z7uzNhPV8hWAJI
xhLKgINtEHEh4w/ZNoepP0R9PeKjcP7C+GZvKXFaBUDm7JZI5mLezHXLFK8LTt1c
PtXFFe28MsCgip33Wesh3+7vD5lof/eyAZirmxAAV5bS9O7swIXbTaQvVnCPbu9Z
c9SXHf2FqCC1m0dbd+YFYj0lD1nkKqTX6QZp96kU1Bxwx91GmRfxX7PdTEfXu96O
mvNjszJkdH8Ir7Knl4LokfMpZgEP9vO/y3HfdMgu+xEH9E8mAlCYLlpmnwYO+5FG
oWkYL8pLbyL8hfDu2Urq4fdVDg9f6JVmdv3OYF5Js6Q4tkQelspaaoZli/M1Itrv
UuHsdaK1WdF6TaDpi1NshF23FswJqQg7mNwX60ZHNAu9HQdTKpiujQaKXN4ynOnr
uFNAit3BiVLEdXff0i+RYNF8aSTpmE1pbedcSydxKjTeR+yaiHLXlEIutWPC381H
pRZOm2nlZRf2vSinz7PtYDOH+tOfPcDczkKX/flzI6oFbxsftGipRy4MiRnA8J31
EVaSm8tO//7rlnDWBoVIHtDCjnxd2MP+03qpca4cz78hDRxCgVPpGPPoloxCaMrn
TEcSzrDjLQdsIT09QkYev3Vedge6/+njqrEbfx+WNSJBppHoB9HMYiBShhDyBOpx
sfptXdhNotCe5SG1ClhvQ5yIXsKJ4NVz4asshjtJet/7Cl1zFp7jF0Ws23DOHFio
TdqCKSq8CQ803x+eAJki2WfYoHCkRPG7gTWPMrYSNPCE2cOuHSYWRdfsW2yOVk3x
dkBySzmkqF2QZ9vrNtGV64gQreb4CCqtNHQWiU3Bz/botcwqVlx7voB9E386KuQJ
e8xWkPZbjF3q7cm9Xw81n1oMdnmm/2rtTXL7Tr/DxZV3JhHTAM6G7D21GxnpOQCN
zqiZJsHqn/z6dKd/sKzvgKZWQkolihxlyxb+EBeNdeIIuvL1T2xhIRVmIuu7bHIH
6PaH9H6J+st/vPeFH1FqY0UOCNzciq05VCEC8hLsdE0vgJXadCkSX6a0Nf+cJrWs
8tOnanQGHf3fUbzeSCX84qLBUxRKcTJSSmyVYWfVei7ztYrDm0waYC92wxaLAthW
4YJsfxCB66DMtiqr0kNhf1XDh+4c6rQkkBScEJkMrRWuLSOy7a08mqqH0ZLksYxP
ZgwcuEakdOv99s9SRJOaw9k4V2n8ZqE9r1KZvhfBBtZM8Zo/I52XyDP7H5qxk95E
3ESw/9U/AwiHEXG4Y2/7qq/9rQUV0FODBIQiUpsiPY8xLpoLgM4lMiVLogzD0y7G
QZQmgrWFpSPQ8DTRz1qEgvkZ7E2KyY619OJdCqdLGK26WQkNwsHVvbkF8bLfgWzt
vgptjOYNK0p57h9MBNm30B2lvHUfSJEtk3+PdLf/k129ES9fGXodi/pD5ekA8El8
bzWHKIjpKzYxtHOUqBqSdh6gIBwKQqURzIqu3L6YAE0qyPz6vaPGZM1mh7+SuCp4
slp+1H7AncA0zwOmkzm3n4fiuJX1z1B5sEVZ3MY7Kszr34BlE3xX2V+5KzQmrWuj
r9cZke3cOWXjkMB4Is6wbwZni8IyC5PUBFUjno7S43DIT6XA9BypwgrIaf/PmeEB
4GIPAxBYM48Et2+p44pNrwtFSRboY31F7uc0cTLFH18eQ8EqvbeLSzJj7G0Rgo+I
4iE6o/M8+oxKiu2VaeuDj6RTRCaXNdOJ2XnWRNLjrdYZXDP+NpH0XAerU/24eNOb
3x+PopMFVvoq7tia1Dxujn5+/5la5QCRZ1ngczcgNwBydm4DaH0pdaphgvPgiW86
gCzPv4q3MisL17MS7jVFZoF0F5kmY/ehKpMTho5rZA3TKaXyvcAevVK+mPCW6xzS
WXikqU4uOANRkRxb8nEnC71jf+kW+LNHrg74uUBVK+ymOIhbVknhbuQNA52j0biy
NVJp3HyBAAsCtHxvGQeSr6z2ytCJBCvjZ9L0ylVDiV7oEU9zrwaIqT5DahvibUbK
Ssli/c7xGJuAZYQrsamRa40bYJX7m6BJKtrem52Zm4nXx9PlDTL5hAKE/w5fN1Eh
J17J5DTZCuBP506lrlB0W9PeNT5ZOocofM7UvzvucDfQDkxnf0YNsBfYbCEJg2Rq
oZrsPp8HwExWt9S5/RD1p4QFzRo8y+/BQSoFMGzUyZtpq8TXXkrTG+niTjZ/4ea3
wlhbyTLGiR9VycGr9QS6KVGr1M9p1ld9ak+ndtpFKTGPqq1EsjFW+qcgt0FuDiUK
c1I3yxm8BVjOR0pRDA/2RJ9kiO6ZuqM1LFx+ybP4whAeOvI6t7BWE6eESHGu5BwY
PfrgWWkdlEClhKHlHCyBF8ZkwmWu0NAp97hPjrTXD7eiYoXA4iLB/a8U9hwI2tVw
Rb8721TrEpQsodfSNZwDeNShNPaGAlN/O4kd1hoAszzHgKXlt8gL9LL44nmyd0Pt
QuBP+uVVVRuSjP1ZYejiPRwWkBNi6VjIN/63uPmgklSS4Y8kN2UQLElS2s1qaiqx
zKfD5cvGgre+qM2uQicEuxML+in+80YnuUUKhrFt2eOJRCl6F/664W43GwMwYg4g
fr62f6yQ5zQX5AY2WN6TRnrULtNb8bKbb8qXe4Zfg16/NCV/cXct3TyFA4gBAB4p
c+HdHDhf5etBpSI2gCvhkCPTM0YhGoAbH3szDMjAThwFmTPtLGUEdkBQyWbZMIhz
JEKpoexSPOtS0hJBLj38MhEAqmRRpIEKu5vOmM/HWgQEaID5lLLisPiZh6m+DL4u
wXFYojCj1dONEyYwpWFsN9g3ouGLOM856jf9xxuRB7Avqi1Ij8C6CrPswn1GoeCA
bVHTVm7f4NHXKNwkxd/XjIZEQJ1jAZn4yKhfR1eWuaYBGTP8WETSwC/WzHMJzucn
shMrACd9I7H4FtHt4ALB/PwSttvIzwu+c/+89PPbMAsTdwGwDoIIABe781ROx5Rm
7TWq1BCBO/WxV/rr6oeM9f6ICr5Vv0oAiLOYvWKXfoP9+ewDzcK0Vb5Z3E88f5j8
6yJHYHxhzLBEVEQf6Otd6I+A8vxt3FL2Kt+4pk9B36n3peOQqsyzyEd3U3L/rnKQ
dZmjQHFWFgU3CkN7TEK94y/rXF9vf42l+V7tkNqlCGgcYkSRBLzQpzNm1WtaLQ6d
CKDjcUcJ49ixHVQK55bzNZf+c8UQqkLFnrGipZ2eMccrhHMDIoNVif9TU8/Cr/4a
LvbbaXCAKVDogaRHyY8AB8LLhk4asp6UFiG6Cj6ti8+NXg1ugGS6AgxktH9aa473
NzBHkuw+YQhvs42gg5wFSPmGdOxzdM/4BRRKN2F+KHD2wU9QXnZ7BKl8uLuSt6n0
EW8koIYasZ+2g1cwnyOxzEs1xgRl00Ri9I5TGKAgCZb2Vx1eNQeJ/FdED7e5AsHn
rnfU3tRbVC0D/6JNOAO1evpCrmlMXs+AcB8winIM0R7/y1iFsnwDOXn6TpTZhO3+
fY/GLApaRHbwEgKx8jfireSVXMYlr9PkBhNdVmTt5813NX2om1QaMQVO8b8dv6sb
3yn2iVMWQM1wyLoXO2U2jmXV3wGZrquURRPXUYMoNHdXfRoiCXkD09L9/8wJofoC
MRd1HANID79GGoiR3KbAkxZ6XLr2Fey0iN7EohJqx9VYzTisITRN9Ihsv6OlONQd
wPAZ5Hcz2767XVHQYsCaEgWW5f7NLwfe8zeDmJeml7+W/KHHj6mCZ+K27y2xzpgv
8yHcccbkxnblwyl/5k/cFjjR3N1Uhoggx6GXnNYv2zamUpfDBteENUIOUIDP90bF
eHEqTwMet7EvjT7qtdN5jLmxyFvGUudxp24T43Y6W6R3R2YVkQSF37mji7eORYm0
FcasQS178OgQH6/Apk9wKF5hk2tvZwPVZhKvU2J540p4o/H57VJuUMojHtYp3o68
SbXBiNMPO3+054J9TRJU9O3N89dcfe65pYWkH75BAqcOkJXNbTzd+JA4Y7E5cPrS
/TUPFS7bSStv9FFsBtAAdcEImD9YKXrBruzmMtac3womEkix024VFi4bOHW45R6m
dGUJ36eaMbioInjLGILmMR+5yYuic/oXgcq2TppC0enqvHKTfU0wvFZ0v7UwSB1a
kfvi7ZI81j8b1qQDzkfA69frJuZh9y/Cz/3FJrIdn0Cz4GbBgTbjBApCZEedHIl1
fKFD5zb/78YrOQCGKimOT7wovE2M5OotT4OydQlN61+GWXl9Y14Hoiv3bTkc8b/i
fNHiuS+dCZDMjXeeJ0LyuriYmI/2gS/V6xPT3rgkV1YC66b2UKaoQ31N21X/YXu8
MMg0iDexFimBRhlY3c5M/Ev9D5j4el/OgKCe/mrAuaNO/zXg0D4tATq90WQzSLAd
S7ps0kcpgp6sBkuFCaLbBubgIkjV7nMuvmX1lPovarGv8lgOEpobuIUHFZvp6o6H
qwYlOvXxzU4hmdUp+jTTVRJ8ze2SWPXTVa9ghtRcnuGVbm1kNo4Y7nlrKCtHBexn
ekBoH6bvMM6ZQ7HFvU7+QObogT5P0uAU7TGAPvbmx1a74wT5dE5RLYOLjowEf4gf
grVUC6Wfzm6qMXhjfOgjMVMhnRFmhl3lRKdsYUGtylFjaiOvoHpro9v4MhIkRJ5l
qg+pDc3uMvg2IkLHCqG62zkIod7N5Y/pykoAfCUyZjpZfr9m+4hoctTxn7Z6GLkm
o/yNuJPp32zgH7rMtHJiAgO6ZcqRUlfrkWAkGV2+O0r1xNPsME4zuvSSq/kuKGf0
frlPCRjWsxWhP6Fjo8M6ZA1Q22pISvJJ6H2IIqVnWbf6o8E7b9yv8S5Txz6pOx10
aAuviaGjF105ZMLJa53bQlEE3wmBqpS+KNH6jtuyGfAYZXNfDdTD0Q+dzR+j//pE
ZkNguYimqcONKiIvzX81XPtSsW6rPNeWvtBeEmWlnNdLfSsnJZY5hmJio+ieyjzO
qphuCZLMTwKm9NQ0z/gAUyRvlw7cZN06XeJLYJ3m2V6DqtcpuA4HeaGVDJNfQms+
x9IBd2AxDnZl+qqLdElW3KOEspp2M8a1cQUyt8TV1Z5ItpciX/jf8m1HfmlIHfVq
zDyrXon+cgPXpWg/WOq9Kn2bCAyZ87kb7+9nYdjK29R0E6kTtf8719RNaiL83h7E
UiDi/0rcXq3p7aZqEBUWpglXO1CrZ66aW9U0dYIyAnnDvkZEd3vjwnsr88x8TT5U
9lPxmGm91rLetlMJcfKnU+4tGL3kDastlwdHw4eIxY/5ho0nGG/OBnAUoY47h8Rz
31x3+JrnzsRpmL4CVl//HnuaZ/iEvWUI+kYJTKRpyYpdWrmb6r//q2O7X/8xhwLW
geu7XeOxFHMzs2mojmXdTHwrIQAj2Z5K6oWFGWWBNPWWkXaJc1iv8QIy1dSiBOAZ
riE9OSLZfu/Xz0kdAera6XxxjTli7VhTyc0qaiOxEIpfjkPzms/HlZU6duxBWDUs
WM6bkQwLEhxaevOLtGETlsh7EubCudn0KA91B6VLW/qaeiaToqNc4PNaKZ8B7/Gl
F/DgzJnaHaDTziEGclVR5qEUVBoERm0VQotKl1GG8FcB8cUVAIg3V+MsicyKYTZE
kcbuz47EVaRt/LJnqGojftJKUB3vmt5sS+mt5gf/Wcy7Rs/nEW/sL+5Mni7qDK6B
wTQ/UlHwoQu3huq3sH0zbMZtCERCcIlMeikybvUjevB/MJ8DIJ1q8YjtfNfofjqn
jqJVvQk9YT2NhGT/fPo6XgTGU/mJwCTqD53Cf5zlmC6UTK1LScmGjlRX6oA72WoP
uYE9qp6SEYPoHFtltzf5zE4RXGaniorA9frU5rpBNp1AB9AwfamPJ1Ug/vyvRI5b
gMEd5Lv9W49PCmx7B+7Ryy3S6b0J4/Wz4BRgsk3KMdIQMo55Iea5L+XAOkg2KZPO
YVc6E/pPFZcLUq9ZtAWL6FBc/qavxDfhv9y+B6kPhmvAD7NM7jW0I97GQbDxH8fG
hRVlcloDJe6sCvrZRy5lTZY50wdkAzzWwhY6ovp4zNdaMEoN6JLwZOoZbCGinrnJ
UeBfuDLOTElxQ3Qroafaj7biMJGGVx+gtXlFmw0GmE0yV9JEgOb7aSYDAN/IkkmG
RWjLP8JD6jCNCeUB+TkDxqodbOm7iXpJafUiKx2wiqwAYk6B79zVAWLyRvVgmowW
4pF0gwiz+DMJtxcxTAlCZ7rgBTk6oXLPdoGZLT827lqZ77vMq6YcoQ3GhVMC70kr
PE1GXjBgasZAmFBYEzxWmG01ghpVOSFbyd9pDmX3Wj5IIO6eOBu0+gp5AKqWGQ73
vO5+fxb4tJ/9scI4l3lSfB2zx8woEAf6KlfoFsdL2AfXusPVbOtr6SiaVaSdaEb9
IXOOzGh0qXm+X2VynvXosKnTOsM3V95iyVquKMhU/2jtAQAwNX5X1c1bJ3t1p1/m
A0MkU2yI8MyNDFPArTZTdgQ1uzmIDOLMqzHESKpo+tkxL1+M33uKmOTYaOI8W8Kr
MtzFZkJIXD7QJM7M4N+ZzZnAHa5O4HnZTHfAgsFrKyqcSOtJrzSibJuO/IduVYAL
AOMPgr6J8Pq3USsorNkABd01hvcnUWbM+lFZqBPsOI6FbyY8S2UmsN5JYTtBdxH4
XctTVcc+ymCVUhvps++DoXlDZftDu6PvEzyuXKUmzjo+Ui/oHFDtQuYPy0LAIFsE
DSqhjguOdo/bISIFAcW3OlvCSu2tpSRHQ0yBmfTuSkHXGxk10BVPazmS2SUCmMdh
xTOQXgAV9ynURAUk7X2cPW08T6dpxKc79pCnRCT7p+K7we9CmwB05l/AusqF1fa9
t4+mviCSSHVFsPoeAYAj2YXZWIBggYc2Grgd3XgM9jpT2tMTXqOuZMh5rh03Ys/4
JJyf/+ylCqtGEUBKwOFgx4EdJr/L8me0ZmkI2Lnsj51V7OW+6jbrCcI1fPt2/4nH
EiDsYDIMfOUn+9kfoxQ28B5ohWg4e9mlfrw2AtE2tOtvVpAxNlag/AtYxOg34mjA
7j82y7jEe55hkgcBWqJ16Io/PYNTT++vo2kDOoOici1TP2BrgiGF+my17AP3XtAV
I3Bh1xgxAgGHsmbuE4JvQumUoYIEHALfAv+hdD2W827za3w1RFp3pqdg0vsf3Oa7
j7Eo0sMPXhpkEsElVbcFIuR8d01KvO7Q3EZveP3oFrg686UlXpQULi3bZHqgFJp9
MNTrYGwcsskxGkHC+1+RmYXmIYA/fAkN4hMSAE5cd+4O04aOLDQNOEkclTaW6nUC
qHS/qHnI7xmL4sm7OIxUzD7I3qfSx+OsIqoGdUet5yMrIAiva3Mj8gC9zGMQ6CY/
0cvO0OvUGefmlfbQO4U6QSgCXi1JlDF/Qa1YjZuttg7f+ZJxMSG7BPytZ+0obrfT
eWVW0ITOc9YQPl0svJh7NGCglI1t6Dv+iwN4foBBUtizW6yvTS94uexII+23j/qv
gLvxO1iyIP7L7kg38v1sPLZe3OVFxxS7uOSb/Oc3XWKIEox8pt05kKXC9cfoS7qX
qv1SJuo0xlZHfAAY/IKZ+bFQ8VcZtTItX4MKv/0/bdylCIucMJF1SXx6+xt9/yZv
ymqkwwc9Agc1G9flCBo1hgZzYHNsU9XPPUhUHD6NxlTGoR1FXLx8bnTsfWVuS4wg
sSDSnHcinFLaGQEH6wfqPlcL48JdZEKPsc6LcJGjPMyz7zn/cx5zYkUG3GRdQHtk
vxNBVwTFzGdc/yBDxVeQCBBwd61phShYN8MLNcsGrMNuDWsKZMih7Js7KNgo0Umb
ZCMdaDw3BJpNWNK3XRtuotBh45mpHYiTecJFlulVv9WZPQ9Dyf8OAx3rqw5UeDK0
yTKDChlSy61NqkDipSAsO6n9VFBgq0u/cmW5VvYfw7cyQZpdAKw487IAL/zS2osl
waC5PqzP7Tzi/Rm4mt4qqtCJOvplYQ4lVxF4TIIPhppgirYpS+Z0xXK7jzKZ+Y5s
TvTowUShEJM4aP0pzSGa5+Tdw1MZG1K7WcDzZk9SOnDxu6ZjW1IXmq3EbTc14Omp
DQLbAfz25CXuFQGITxGpQ8ldPI+9sQzFZltW+q+bLshz1KgmICNQTyzAk5+fCMOL
uzdGYQDh0A+7mhxCPXUSaZDisrZ83JSJyQOT2ZAdOExZcVybzuTcppcFUeJbaA4N
xam0mHBicnMOtD8yIGzIdLJ+1m1q5JrecdliRJpxvIUa5rtZCSyHpq8aCiu33USn
5K/GcNtmFvzeMAYf76KZAUqdMVbPFPqMikVZxbAFMAKJdGYHi+tLjZHZmPDGUJZA
FlZidH7KmOthTqYehIo0HdhLgsg6+CpgfNxtmD10vrjVwEQBWj9FxMty72KwTmY0
oZPXT9X1kGjp6qCNB0GoXhWOdySqf98TjjYA20G3paAUZOg2AtiC646ZGVkvI0Vc
XhL6qOGZoJ/5cot1aUC6DqjCkE5qjHeQ7iYSNMyFB2pGOiLpSiZJXgmGJ/+bcEOU
O0cq+3QLrbTFHZR7PBX/s0ik+SAoHA7qAVBIyOF3zRhPkgH+naFI24BSQh6yO861
nIx2dkNCboxy9Sk+e1uVCxI6f2wlSFrVggE4Tk5PSb/lLV7gzbjDFAqXzxp/wL/0
11YdxprU3wMQzF3b3cC5CMJUD6rpoP78hvQuVblxYpIIzOtuqCqhCNdkNv/W7UI6
aZuPx67B0V/jbU1m+TnOYWStbeBQFJvR3aco3HHFqH0+zSilhQGO900g0QQp4xiY
JL4Onwt2UpJvJR52/Ef2CUOvM5haD+kjHt9Xu+ueyPZnQHDps5jr7acZtOUIV4dM
cXe2WeA7ozlvwMDLmkepWfNnBUt5Hq18kALmkIZvVUi+4Ya/Him3FkmdlB4Of4TF
HL6RvgNd7D5B3lVGD5yJuVtEyYmx6DO8hfLL/NOUF+m+ONTfwjWb7zqhHLTMQ9/W
ILBkPopeKCanVW1N64ci0DmJXHw9e6dSxVP3vKAZqKLUd42UdNkLMHcrEH4VPMkh
eRX2oKnllCYfnVYOyvmsqL//b1V0Zal1Fc3Q35jJSojGO8zr2VsTzavCIabPwk+w
HhIRO1xKpvEmjNwK8R1gHFPLMd1ausQJPAvFzKA+0VoRCrdQZXsDJpC8LrBGfv2R
oPmrmAh0BpN8HjAYcuE4Sc22ut607zzF+hlA35U6GDWbey9KP0d9MhiJZvGd+w38
Meb+UMddADo83JFsRE0BMvDwycXFe9+ENpisrL09tVfGbfuEFRiZ5OK1JZPqqpCz
wkl4j/pLiuHmz+XrbhgzyZMf/dOBIJ8GQchnQLbcKDczceZ2qtLBviOXlLXxmo8K
SL6kuc65IALvuUydHCwxyw6O7rEBkyP0zB+ICkDrpsPl4duSrrB/HOqv2wwJeMfo
apUKlbOdEXkz8KGnMwGPxr953yz7llWR3hocusEzA31yr0IBiy42gZfMzfcT19bW
CiFHV4E+m3ef//Wq0+v05sZE2AIgo6AXgyJZMe2wotB3pxmCGD3bOvO757tMsouc
lvfrZf9e9y8AlXTpi78/VKnCePZS5CNKkSJ5KRiObRJSSqLqp3kRe4OmLNw4uXlM
boEofw2FIr333NzCWHWfImiMGMu6i1d+4LabNN5A0R4HI/z5Jyn91UpCj506AEpM
XdD8VG6SQV/OJoE15M4C8tfcAXA+VQHFpRjSksPLhYJPF1anNxvQehp47eQxdPvO
axwJTRKiPpmhiRhh+OrXnHr1ZS4lFZPIPZhwg00ULmdDW6U+8HDvx+2EMbgHNN7G
cV8ZwJ9WIUo6nL/23g8QXxMTRd01ZS+L54X5TAbcpm9R1bKg4Hxy0Gc/8OO/9tRx
sfRlAOG1y8Z5vrql5yvFL+AJNoACVt9zfIEEmbC8H2qPERK22rq1geJSGe2T6SHa
J+14rwjq8JOUSTtnJ/L4anvkFIJI9lFvYALZSSPsNjSNVA/EO/uN7aec7vM54AtW
zot1U/YhJkymL40ScsI0zzybgr0rJODWhmxXd4cu/9U0apI1CKmgyK2PcacdaZdC
Kwg29EJICk9OLD+Yp6v0I55j7a6BP5HEnR3s6IlZj2hjJUf2ol10OqjVlCMYPBnO
Rei13NsO3bc60TVge9wnA1UhvfJcjTLjOfdZaNH8To6gxJi5RppAKkPzMjrJNSZB
1kRftaDZ5IfGscE7Wz2KnxfXmkFBZmpTDkUPpVQZlnCuKzT+o2or3LbpfNmC/F4K
pV5G7VB+FBSvKKk5tm8F87LlHqU4f3Wcdujn6EIuBAFhhQKm1g8WgUXliMBGsCbJ
7P27lHFhqeSYg9PLucEHWP3skLg6M7yjuHpWlagws+nSrWkcoZdEpqLttLwStSEp
h+UjoKBgG2Dh+cWCgZvQL3ZRz3KW6SLDiIU1SmEWfb8+j7eX50y+jaMqOVZpw0IT
zYWK2v3iyTbPviAir40yGSBlajY6HheiEOc3XV0XaKrjZ+jp5vMWysXHM1Q3PfSJ
KnhMV2YS81EeZJjesAT31CjTeQNvkf+lWVU+O3ixg5+oxy3UNYklKbSDZZt9HkGY
tfehej3DUt9rFRuocoZewXMgKzjGjQPessgyV+LZTjCb52FoVrkAwMqfVhm1CTKQ
B4d9Pjq1Q86Aza0gxBe5EsIoVjEmcp4Xyxp/jo0ALyqBjsA+/aRJ0VUDaa4ko6N8
9ZhEeGKvL3BYKkUIk7DbV8ghZ/hJUGac2SL17Qsp7od1cxvLxvg9+anrEeyInliY
AWzVr6VHa3UdB4wikWgfef5r0NvdpwEHSK7zkvAVZ5YPKMkgPuqw9oOxZ0fxLIVu
XT4s40aEuCeucunAH2IA1KFOdbFcxawW6MP1X8hEtjFqY2RN26lB+pMhThuk4OE4
mwkwCMYEmyYF2HRCl0e0w8enfxI9wi67loaMEmCTlCuoHI3ZyREznlCLlpqDK8+M
TRkIDtf6IpHz86cwJKKDLNd+g0TEf2sI4YujI1GxXoR/pPiGgbUnZRX9ZtlYyuZk
EGolhaY7iell2NnHMCWp9eJ4RR4RHYDE4SrPXnwH+Wyml0yVDPEDvCuEtRDOSKJM
xSWI0Kg5IqFI7y/iBnOBqIe8yeGCWwjIDW+QYsQ5Ly9npBYz9cMofIrUQZbZrr8i
8gUUKStN/u+Q8FS5RLmITcWzUUrGD09m3ICP1fB23/SQBmOKn3RmLtas07k/nr0h
6G+fZgaf2rF2gRe7cL1JMAlHI7/CWF/TXdQnJZWg0gPysuIglf6TyP7QtBKjo6D4
XSxo1S/f2dwz3xhiqzd5wDLoonaqVzk3ezn4kK+nGzekVSeu2LZSTy9DKKCGzKKz
exNTp7bWbjOpmDYImQWsbVNoB5ItMUThBHfo33oP99QudtlqPrKAPwf8NsTprL51
oI7yn0WJinG6oVloaDjT1T+Z5WxiHhaCpmalHMIvsivKdDMChwdQzNYK5ulBX/IE
M56VkdWYnLQWyjnOrYIeA2nPAuwhmxiUijcTFR6XObIZOw7VDpN3ehBhVgfR3Fh7
npbVZM4hjzQebw/XPaq2EFq4/MHA8PJelEENmIIZ+6waQlFbI6mSlOcV3Ln0IWzw
3l52nnFawA7PuzYHd4zd4De78lu25XN6aii/mFetDtE40uvDdlp6/H2mX0LCstl2
MnQgZTDxx72iI13Idc08GK183HXP8WFpVtoQCT/B/e6XvYUBpLOxPbacoDTT6LPV
1sIklx38yN/mfnUEqvpmmpeN/CihSDEJkoy2EhfA9kYLzJTryCDnD37orZwP4eHu
pMMYHxv8hPROjMb2fJ3ZOckqhvZDxnfzmYwDAdo3mQp+Twr4JUIUIv3myGJhz2Nj
nIAZM1FEJuOQ2BdEo+9cMVAHrlHAn/OXicwuF/w5jm/BbJkzGx1oDKJ1f2TBxjv8
tDftDN6LZUba0SSFjL+G3T+Z4lMjqlqF8yJW9Oe7LoxYwywZ/g0QvM8rM9aYRc+I
GYQIBTI2VZHTRSjRJBMu971NAsn+u1OBNU1tmQ4MZwxyF3qoB6QMR/VxdLmSsN5u
yAY8Ks2CG52pA2JW67mY/h5cppcRiY5f3oxWGCxl+Qo9Mvesu4DYsUnOKKBZKn98
8Oy7uaFi7CScObwL6ppJac0zFg8SUAcHK7ck6hYv7oHQLDkkcV93L8akNm5GgJv5
Hsn9oGaS/t0WQllafdQUnrSe16E1rlY2st6bkTX9iSV+efZBDrcImP9sy6X1M7SC
wb0lKDvo+XCNpr2KQZAjKckIZzH02nraWUI9NifJeEP5YGFRqT2VcHwMJ2Gu/p9J
ZSEg90xSWLNjHXwvx+U9N1VdLbwlHZgAOXZlsI6j17bfEQdVuFiK8ECV6UDE8JAy
6v1/qg2i31mzZYbvJmWWuYRGYY3X4+e0d02xGLlY7muGNqI9NF/xvR+/IwPNnGAY
0HLqiMUBjSKslW49gyMpO8e9QkO/vhSHeP3qVKpuotrxXp8I3TdVQbM7dE4Zakqw
J+4bxaaBdurygpgVn3PIjSLJT+0PMDUcIDpdBoeZdJn0rN8C05dSUv/t4DPLVOGC
HoAktBtSU6CdF9NlS54WcYZm3xkVbCcy3qrKILWu+hR+T+HFqFAUxVEVg7Ss3nwr
KdGCHX33kqozZxjGkSyrGGCW1s/M4+nsRDhk36CVn1a4+kueLwuLZK/8NrUGaUkN
wreHzhjTEdLMCTxbhPfSaN81NULdH1xV/H5L9eZwollJku8e18tBJ6RgyeSUVwzL
dFKrG29t9nQV5rWIr2S3033O88JUGgODDNAl2ewMjFZoVwJfFYdywZ+IdFHSp/w6
rE6cE6QQHYstKESCUzxAFcWJe0O4EjqnEydK+Nv22gOmDK5PVM4eIqraDlqXvikk
3wMgupUyZUoOrsZmGEWfWSGOEOp2kbJRpXNtCsDXkYpsvb8gRhS1FeL0LbD2wea1
sfu6R+e08UynmN1S6PjhKBLzYrMj7oOnDXuDaNXEIlI18Il1JGWOLbt3SSjxUn6P
avZpzp33qkZAuFjht66ABc0ZWErAici7Em7Jy9OQooU0VCWpp9Szg5Ou33ha91/A
YKjQeTLw3CbbwZTZWeiDQ1Hzj1wJW7ScMD6gdQoJzZ5ivEAii2EtDKnIaNH09LTC
acd3d08RptXEGhPEQkCoU/5KDBo2HRlg44nmmCE1FmGS7Yz/RaxC5YPL7732xVn0
H520oELlBX/T5Knxoj4BEE0MKyKiscWLGO1tZ2M+DrS0i3/TSZ7szQadw9J/jhaE
evkJ3mNPu34jqZuBjTM3uOW4P2e+A8Z04bUtFBCiJ87169uoPf88YfCUQRdb8/wa
XC22j+AgdCxUdhYX0rS0u3zFFucpKA0/q5tB7N9QokzAR7EC3snKarFx9iIkqEc7
aMmujrIvbbMEeHCu6/9D1FkRDf+11S0FIIQgfxBGJ9gwOr43WGfBds6PmslU9lGO
yuPiIb4d54n8nJF9syN6luVdYPY49CHHuMNd0PdYYwxF+a9tlb5LOqiWNYaI41Vo
DpNgUmDBNm3KOskoZRBFFpD1y0R8J6CDzvKEKal2u7sTrBO/VPFtPqdw5WQ5QhEu
Hb7HnZ4rP7EngEKJB2NJ9Egb6ic7CMeOIvK53tXnO9413oxxsmOqwr0s61Y26W/9
VuDKOdqCqQoHfBdg1T44tOC7PwuLM33FRSxG+3BWzK6aVhop+on9/S38wogqg502
RJKm/ojS8gPIrxV66NMj6P8AA+Sm9ee6RP6GkZt6rtJQIx+t+8v3/OuejPK8CYIj
WUJi+DNkvYGsjl3iUQnCrnQeYbFOkpdTsPPIRyBgzP/QAD0YsLNQlFVlvm9PB7Xk
WNM6/779aRtwsj+EM0WlmE63rBtD3z0foD2IbBpj3guRUXxY2T01J0syzj7JF5PP
diwFzKz7M/AvwNj0V61ae6E3u9mG0LeUSuB0WAey0DAwU69UYeRcJp1CdQDMgriu
qZNRNk3qoSlH2XS449cam0FRSoz0oW9UN8wsaWAK7slMY6qCo7yxYCLZSfunGzYW
8gzE6QwWKy37W7mNoDjF0Ft7nFheoGEZHb20Xf9RjzZRQufXYU8xfZo4LwJykm+5
Q9CWlHOfrvAKOqHbJ29Agyi/JcvHdslS0sSXf6Ny85owJy5lE8xeqRFBbEkW4ZeI
oC1IM4uZchlyRIZxD4CP9jWF/cuoFiutHHfvlii+/Pq9SV1OnQbYCQkO5k2bBm3L
JpYIedo6NBV+ukY0BdQXyAOrzRm6nPxqJk5UFbtIhlsCpmhwiJOGLJL+l1P8f9S9
Az93EDG1jKyg7sWssapu22wiuFhK9OS7AqOmvZGf0JsmNivoNlKMSzaaWmUnI+46
tZroYldRkWY1Jp5Zh0pFDkthfVdm9qUGpHRTau//61kXfOaeutF6ZEEGnjqA8Lwh
SxbFqJd2a0iDhoV1oDlZG+sCxkzWO9dXKBXMk9nrBfupm9fJdAqsjsMkDTU2mHCy
3n8YUclc1G1qizJk2PZRriFth+vtU68PGHt6NQbS73t6OqRNGCB6Srl2Nrmv9eR2
EAlqJIUkuhaFxd3JxahItxJp+na7YOGS4jjASi/jL2Bz67lRRVSaXfFW5x3bel7k
0q6VDllDWPGFbzCbSEeuOkq0cnn5+u/3ExGHzcWK8xQNDNKB23K2p6YgzEtMsYBj
ZRkLi97U1gci3qG++KRNmQ6ZQEPW9DRB66HK2UCJVfwYqSAyLhytu2zTRRB79lwc
87qEe8JdNMemNjRVvY9FkKzI5nzJaLHY4OLuiEAnB2uJ17N9v/r+QnSZN0vA08YA
EkMjImhzpzLcG1IPT4SfCYJV/1+PpF5NY0TFHl74RkMP5meAJ2QVViMERDLGldlg
yJWyMkXE/viNlswqY0xIKfGuRdGxv6XQEPkS3bLEs2rF3ETyr46nG5URO6jb+y28
AA/8wP/SPu4uR5mHlL12Xbqlfn6QHFGCEVRfTAY1R7wssnqTaXdaFTP2fqBUaw0C
1TuWc+z74yIydQ95Ip6P1mekwk1MkyMNZPJO54CSQ42q8lCPMM2h3SAhrF2jSFFh
lZ17lEmdeuyE6+qA3KgwjI011cvAuLvLoznqTOTpWw0BKg/OrRpR67U8tlM4iDrK
Odd3DV245lOaeGL0SIuk4ZvJrp46+BN4dim2tboecSLZqSjmrf29oSNN7Zz5MHxo
muLoP3l3Iytaqkhs8Qr21feVXaYMtzWGSnyxz+xRbST3onIXrS9W6NhJ821Iood8
5/LO4P7S4jLkjrO+TBNOWcHddh59+jeiBYmCFi+R2YNbIapb2OZE/o0fFff0HpMn
i3RrcfkmmAXPJlEjjfRLcQfdJr3i0KwrrEPi1BzPzsKnLhgeq4tTifmzeqan4M5I
LoHhpN1NUv6+hKwH8pqoKqcNjKNbaM+02ImnmIj7QiAYn4P3Mvp9xG/ql2CyYAqn
AA9KbwxSydPUc4gN7n6dE0F/Ht0UEUKwMRckGJyHEi1yaSTjGI5u3fmrNC1lf8ed
vwOYaiY3VM7QBbOpkvjM3WZYFsRC5FdQDbHYdnpB9rvm85F2/KX11ECwY5uAmUW+
W2kim/nwYk1roARvhvpKrCECZ5a2yjOwjqGHMeFK2optNP+DCKLielNszcQ3zojO
hlCp8OXvk7xkwcy3NE5EiiMplBqwWHg1FeYfRJ0K474PAvoZi+Ua0jNHbjOPV5i/
aE9/dedPOEnHl+skoqo1ebRaisZ8kAZBoSKI4kxefojHn68oUq1BjyL15vjZPoas
qm5AIIRs8uYrphMwxCRXrm6KqDKPmY5DojGzzrE6XxZucKbMdiQEbyT9pNovWFT7
OScOe/Gi43EMK2XO5gmiQ4fp7S5dVPBU3+U8Og4Y7lIVD8eJGIYh5Y+5EC75td22
8vs77WiPm4Y5CEQadBCIerKKeIi00ruu5sgjjojVb+mMdYXajaOCc22cNbg1RHFX
O7XWoWZxyemM2m1T6T2CGeTWKq0VgtIl9DxwX3OTk3iCGHvN0oyPIgy7hoBhuZ4s
EKibFIuZizIt2k39/C3RoVJt2BovCdAyvMgVdZotmedA+2//z9fViahf2CpFiDil
3j2CbiVMbDZVthBmD+U+iM7s7GIWkYpi0zjBhdfFdXPtHM/oXmFeuQ8eL0fen4/p
49ySMw/oGdmVo3ZGfyFWy6/ud9ABTp7nKnIXUVj87AONe2XBZbo+iRi8sLi2hk6o
LFj055aDmEFHJxoASwUxejHWWC4Z8sk9DvmOX8DmUnA9GA9qcRcR9+MrBAk1muic
yB1ubbIQAknvDplxCnq4DiaZTMFdSkgC6sxyYylrG9gG09BNqSBME/Eh+3/DC8Mz
FArxsBe2GkYVq3L6KsFMuBC+nn6Dx2HT52Tw3yWK6Eg1RhM2sfiJv+qcmFBm5Sfv
8vvWzCJK/lsLqwt71UZzU3pSiCPKhxsKv4Bqia1tZpL8EMJtOLTM99ofpNmCg9y8
owM/K6lEBD0Ej4wMukSkKBtW6ZYz1ldaIuKE0d4OVH0WP/11UHotj4AmTmPy5Adk
T0zwC3767sy8YXpJnJ2rbWA+FFr5tg+WrC6jxqZwLNyShMQ6wmOxiW/2SUe9CxEj
kyBXqbvlYEmw9067dHu9HFfXmmglNxwO7hXbJF28uzzHHHTOraWJK9GBD0apvRvq
2V/iVlRx9inoZZPSVT+DwApvh+SY3A2PMp2tN6DmC0kmOgR43Vu2ISqpMQWhGUhe
usLskiS7qyrEocGris3R6O0AB78Nb59fqzz0+t6lDOcumA7OkxrX56UfKGWGHX6e
mwYKGvadmWH45e4uTsiJGKeuet/WmZR/QfBzWIY8T+AT7wdYsJJu1boHPVsqVsFx
o6gBqFfdLjdLoFbFecxQfY2wkev9Az5cNu/oHxjIZG2KL9XH2brut1QVpmWxVU5r
VCbDS1jm0VjymUAEzKcRnXODurzjVzCgMmM/u2H/PoW7nR1mIWNMm6glDMvLv+al
LR1hzzEBrQmSCepW/TlwgrH7LyL0hMbzSrrClyIpN4rdvcdD8EoM2F1kLM1/02DE
rsS9+GSzWzOc/CQdSbpvWw1B7Bhyhq6+PpQOsGwFcCFOrpzDGWSHtyCbNIJVpT9U
y+Am2NtZ4WpoXlz9RD706Yq0r5UpeO6g+Zwl/YxP7Spvu2u1yXW5dxD5nS8keRTx
sk5mmqRqiFZw/reupZ2v2Y8Fxb0aGCwuSRu7DDR8uKun5GcEyc3J1fj8d0GXu46A
bzf9O853ZDkdxfO/XEoMkeSphAONwZLzLzplZoAhntVse0GnRh3Z7hp8D1CgWR7l
tfIjv1FX1mh0pccOoyvKALfoG+r2ZeLawuQ0aCbHZwGIzyv7lJ7tCBz7POTope7a
9cvfqTtJyn/MJcWduASgKD4zfQ2rsGbzym9tdVNgCCqxR5gb4oY3nZ2HwEqBOeD/
fHuse11Czaynzt9+upOteReZoGj94XW82PWSbq+p4OxPtVWz9XCriyhBUUR2SRpj
GDGtwGNepbq6lPgTmPMEPIamj1uw8SNPyMmvplxJz191iOuMyGukWCftazcAo+7X
pE8qb3DvLTDUjLLDgF3aPX//BHY/A3os5cJ02GUi8vRaRXj0bQTfD0R79QfcIMbu
svyoQodIrMMH8aNnW/383uXVnvz8OtdEJ3uQDcyaR45MaF5DgY1bDlJDVI4xIaMl
uvtTGGK1W6RtusoT/HreQS3fZcMryqvD3hdNqR8+Ab7XOBZQsUrJnd1H5NR6I1/V
ICaoFMkDkiU3cFz3c8g9Po4EBC0jHdahseCcuYMMb+e2WVBfg5IVHFvOS+6en95i
iWvikRsWleql9MXOBldHXek4Snc9ZP63e4s9XC47ODd/kuMIackY72FDBq2MBQGH
y7QC28/v/7R7JFwVFWX4i4P3HMuTJdFjE2r0slIBc7SOoH0eVchbB/B9+ip3PyAi
P/b3EBDkjoX0Yu73pV1AGFTFdoKVITWHkfpQjEPBN2Z3fSmr2eojwZIO1AnGmf6q
4aSQ5u/pwnAqyCPnylQlOecy8jAu1uCDaGuoREFnTwfkPtAS/KrgaEqelqqIlwtJ
H+q8O8EU/jE+xU1o/5EIGdAVFWcRXItS3++6CWeo9KZ8VfM2LTXeXbXu1MkNzHW0
yej0Fn/tgRLian3/2w7nZ2OVIKcavRHpovTiGUQYKpCDeyHDJjRViQq3OyX6fEEP
A4EChxPxtTXhdSoTdC/0kuj/eS3PIZZMJEfHwiNEvylEBC5d8xbQIEkJ95gxuPoC
sk7grIU2GhStNpHzcZ8JqICImr8bpjFjubR1wlAQPCbsBodboxKG8i0AD0KCwFVa
3u3bVlw0RuXlFQrX+ayG+GD773MBCusnNFqgzP4Sx602edqPKsEddxbGLxz0Ww9d
K/ZJSf2luTK9eCfLTPkFJiVU4WebfNEmhToeS0T+08bb1nma2OTMzldvs+76girH
VK/vh37XgnjCqnJ1+iIrzFp0sHHNGO/Q2DmU+O6RV84vsBh3uLD7/CPf6JGxWFlq
jpOxZXp5Agoz3VIZBZyfji6uEdytqnNYyrfFIOdql1COltMyJSvteGsG70lA9/qd
OMdvdPwL4dacZaJHBt45rP5JAGgHyqT0gIFxXOr1jqQ1Gd2vDL0A8ecqwT4Uk1iB
1++ztGNkTLL5kdb0UOtAMQqjj5tTH81FIZwCuCsBZf4qbQ2uomyqKIpxn+zqFL8H
noabR2dhW1o0WzCe5w7EBZBtlBkciyo2JGbo4R63GugILPefkQnFNCZBw12jL8K/
SHFgrH0QghBiH4YbZQSN32EcAG+GLfvSsUqHjTjaigaq5391Mx8/CmiWYCoPKMDT
JqhlYyWC8qVOg2aDfLFRo2x7q5m5K+PNMs7Q3zUGYvlw0GFX6CUI70XLKGfjC7JP
qdp2HlgEvgD9T8p5KCp9LP/NsU2NVGRV9712FjH7E2IgQIQ0PjIifxpqTu1Po2Ux
bg+p/2T7s8XsYl4Nlc/LUvlOQgDhqia9zmzJ/Gng6+ZOsUpPqEFt0PCb0pVu0lJl
U60ofvhU6yHIh5VDjkZDoKJzMOb9iPJZqWMHaN6dOtOM7kPZtlBwJqn2pqutUgcL
ycQtY0ziu3FRXGH8m3w1O+EO77Q9YlF2waHCri4NywRLyNLeS3U9Cy0S3VBRYrXa
KLbeVqjnXN3IVkyYQiqrJ81dlebI+e1WXtrZrwZfN8fE7kdq+iJ6aDbSGRU2ugf1
wqmwHh1KeuWfQD1Slwq1CvZSJSPvUe/hQVGRix6Jd7t9Fbwdgr+8ckh5bGJhiAB8
Dd2qUTtt94AKTHzYlLytUDgdqDlgJWuiErcm12LMV6O/X7aSXnbbkCI/s3NDLlAg
mXI7w/NrTd6dqAukecQcA832EM8ZxY4StO4Orj0FmFbWdE+HXHWvKX7151W5aqGS
XgzcWynnoLsvOySJIDLLBcsaTn/MHrQbDArHSle1uDY7+7F0PpOTYVvGf254elYW
2hnhlwUiYV4jiRdr1NxEbrit4xQQgsf3cD5ggkZPdOsjWu8Ig1SMLz6kRXumJDkE
fOzd3gsBSrplxDvBapf0VWE8hjLtaE7V4bcDqB7B0C426JBDkyP41YRXoH0W9x/M
qc7NyAWEmISEUEbjqYDxWtTQx+gfyQyz/dgPjd83qjfeg1zxHYo68hZOipqCl7nB
Ldti63XN/S+qmW29vK6Q0WiYT3A5JxVdaxwehHmnNq5o1R3FDN2ChiwKPGGXMqXb
NJilkua28eY/H08awY4cIWvP9IlW1QOsHpNlxbHXaRey19hqMX/CzB1b7ymSHHjm
JhE17+H/kMyR1kmKIxklxCkGY/tjr4RyA40F//iJNQXgfCmz42fJr3NIgnng9u0S
eSGE0E0NAPeYuc18dpBe48tPspnSL9PbEgd9fyTDu3x8XRezEI25yu2G/QOeir+P
XPt0xb2OwMTxRL0hAkhFbkQwsIGNsy7oIz7gP6OOCcOWoC+LCuEo4R5O+c3/Edml
bvYBlozqzt5jWKpvwHBOYj4HtvJzNoJxnABTSOUUr9IDJshpHMS+Ij3H+u11w5N6
qLBHolAlKub3lJATtHldk6Up9lHArevDw6YJjp3MXSNqaYsfB8rquN8j4XuauCY9
xvz+S+Ip+ZewsQxJmHxb3WHZD+NPqkK1OxLPGp9R1I1o9aiqlaVBq9YDdQR71IU+
t6dvXPEEQVKupgzu5o9H3vM8MCyw9IYjSysIKpp0sWoN1tJF8yALOCBuvlM1DtN+
nCxmOdmYdw0O1EP/8tVTK0Hy3jAgIPB/Gs6YSAiPgMQy28mdtgmrcVm2qzwUvBes
9a900MHPfigw16+YcS+eIcl2UQpXobv3FEGs6PKfOYxfDb1Cvg6s68jl4kZaLBUH
+XAkuJC6RlzWjoCHFYP5FGh02FWy19zvpq1r39/Z6+a5FLXBePmxKRkH5vhlcKeM
scGZpsP+/BKnWQLJEG9iAFUdO4agWGbFNqwCXQG+7Jcmn/lDkbjuUAPwlnV/AdOy
Y35z0eezy3+qcDRAYxNYTR/uMKgqMqcbuFezSSjWI3zQWr6MsgsrRGI857mHuHfb
jHe2dkE71w6bomtOZ6C/qm5kGh+heVbE45e1w62c3DEsaqb03Vx7dZjgTKRJqenQ
9U3HB97bzFNmR/AYgdJqztUcM6rUyq5OPaZZZI84Oa9RQP9hPHoFuRMy93Qho58D
UpLg6rEgUEobn0k5BsSm0rh3ARFPA1CpVWbUdETj4l7vYPBoLIYAQ+84cuesmetn
P2FplgyA/N2O/dBHEwfiwBqix/FYvLvi7XzKJCij2BLt/T2ONM95etqNSudyfclT
DwQQRf/z+xdKjTF8Aldram3jMSuEbI2ivKG0S5B4rkRExLEUbgKFn1uv1r1IeQMt
eTwrbfTl4hKHi6jza5jl8ZyzQZsw2BsWBdSDsF0YlgpP5jJ+Hs/WUkDIcJPnoKLA
FTIh2tJgML9ZGuj3e3R4y//73xgL4KfjdwbMxJk9nM5Nlm2qlZafYGykPp95MIDC
8LvOXiT7rc8lleAfAc6qQklz9PUO7+JxPgyiXs0Ywx/HhBq2ELa8IEL0MqRWwwz4
xzt3117KequhNkoDSDtEp/CRegictQnjbNiNyab6t695hOg1BOS5CTuVVDeC167q
15LLFtbmHOb/VYobyIYNZD9KDjA6Np8N4v87fVjoOd70VeJcj8Yarz9aN0Gc0y0B
On+sqlrT+8F4CuhSa5yBS3IuR9S4SXjpAlGaP+Pc86n35lM4EhdWvEblBb/LO5iv
D+E2IToT9e3njCITzmhMhgKOXVG+93WYO9lxttb81yVvSGZN2Oi9wRywSE+8+3yD
aVXpgzCEtrPh7cjWK3/JMCLmc6CFdcl37xnx7VGwD8FeYhsy6gCbVOYzVT1DC73T
I+aD3dzzO25p4qbjtsv06sh4qpAZfl1bCDBrJLEKAGWjowO3WEhzPCufa8h0V5Sm
iyAqxLtbzUAL+BRIYKLfPk3YWq1rOh1VFA9+P7tzEN4LEKTwofYfMkcNcbjtBPoW
uZUBzgyAs+74wwC5e9D9++CPH9gqPba1XSD32McviGi1Nl4Zb9juHexc8KIxTIrc
2lFMt76hx9YYnRFGwejNT0aFVTYrG2gEGyrKNBQufyeqmPyueJ+eATfk2Rjzb7Bo
hwlW2XNarJ8fwcRw746YiRy/TfSrrKhZmRM5euVPMqmXMgu1QdsG9+ZANhi+Eepu
X9wx4sE2e7Xn/dcfP3mxmI9l4aT42IcWWBBj9orNxpHHG+htBuYcRATIsMr/MzXp
fglU7qh710mMI7n5X4QhZlsSjc4zu57emkNWgZi1dqqvdbaC29IDVCS+S8gHU6VJ
pYd2XQ50h1fGkKBg0pDGXCu8qk0hGdK0IlQi5HjEeb1SBtk91fAfNK8qQb66q6BM
rzkeBZ46kfoRW/BusZV4Oh7SK1+J/y4xJLatl8GXGB0GauuOorOZb/AF927UXtVv
Fpz7vgdQ8pn52LU/HbNPh9h4qQeWYVwHM3oSfiJTTJNa5AbW1ka0NpdS5xIh0/BM
wPWytx8ixca0gkCeU+zsmUhqK5vdysUM4WGwocZg7PEf0NonoZKsJfYXC1VBnJnP
QvVB7P6BgR67y4ODoWGHOQXMdQ09wuDLH5Yp+5yDX8TbfpouPr+HB6s6qoHItS4E
SnlOtpfnqhhQTOCeuKxRKTOwymY5dPbWw8IxVjwx70mrxrG4GJrOjWXs8SP/P+u7
KNLsUC9d9iuC+uKCi5wKtEDsJH3KlC0zcKOZYUqlzv78CTnBAXFbDcv96mi5KnMf
cxFLtc1E2Q8248xYSaExaCB+SUqunrV4S2mFqigaHCPZClmQco4G1WqovFtaPggS
0oU0o8JY1N6ltYCadn+2FN7SlkTczkJbAlu98SiHOGLCtqd+EWcHnMXYDZTKa9LZ
LTc5EXlYPaDy4mHI2aBM6N6aPZNWN7TOOXQyRvNVeF/Cvx4j522mtJKzWNTDCdae
a9/tOxKTeXFH3IFTZKlsvGyoqy0eQ8rq4f9F8nyl5Sl6X76uiXtvYQbZsqZ/wHsy
/FJD1fD7BcGlrgCB6QCWVKby19WqV/xZcOzaiCL8QjrECQGxJgVcfROKj7mHSLFj
37rDQqTDtadhLawXiHzcf6ziG0R9GcJfQ6jfnRGRFL7p0PivG5ddLPv2ctp8J+oO
F7XCbk6QbGWZBMRzH8f3zuU0oEB1VdXyhzNx28v9C9q2j397polMg3f0UHTkmBco
ozu7Ab+iEJBcJfNuwwWEw5mdzEWerBuzKpXWlxCdfxaP4P3rRvs1ZEnzzjFP+Y5w
NoAmWBQRD8UJIlGibjxPHXR7JRPOCCkv/w/I88JD0HjK3DF+Zco6fzow4dRcUQf/
xLs3BLjItU3dJ/cLa9jS3TWVCD/jp1VLNbZIXixq3TeK5MfmiIdeb7iNHBQV4FlH
sS918z9Y/43soFVlEVHlrs86Fi/BpNrDnLVC/a5jXNu83D6JpqqUhteCBSVFO8xo
WGFgwHoKYBMaeVVKLovcYB+mILiMHLmuXOHJjZRlY9k79cmdk7t7/hWxzu151dZZ
slc7kGnpQG/g9Vmmx958z05r/FIla7hsEUtay2yVRy25oeXIK88aPMZ5trDSrExz
wAGOFqrteTtUyl4Ak8RvIcfy0fN3ZV2uVwIFeL/T0Ts0iSa+baWy0lDz8lipBIdK
Gjv4VoiKLH6VMhZt61s3ET/m9Ewuf376slr9FtrpJGrAln3TUfwTHFXvvzeTw/Gb
oikT4BWFqVtHQrjCHUle1HXgsIkTQBnqzkUw/OdGnsVk+31AuUpubqmt4r04FMV1
cJojjs3BSsF4/5ySq93hXSgzINdHOYHG62sOz3/GRMd3dHafed1Zr/VGspW3HKz8
vjuX1ksJAKhIMj6PlV1FDyHGzF+8ickDbJoNLtHg+kYoYDecMMcCAs9Js0QJDNFZ
ix/7VdsxxVVU5V0AwPlzn5dyc6TMFyJUgGMTkks04dP9Ay53UEpWrkMCGb12ZBLw
L+LyrFRwrxCK6PpCEcANsM2Ji2zPmlcLN15GkpCK3IhOMpJVcjI132FMob1CHYJI
qDdIRZWzdKc3N+fvxMz1FStm5O0PWR+Devy6xeWv0YcrSIC/z+27w91Z/XHZluep
LSehZKp0u1oA3tKV6TRF9H+xFbI8oBkE9wUSxZcp2rnZdHU3PsrcH76ndEAtTJnp
TlpgIwBoVukjIlszbjf5BAgqKX3AYcqbs3Fo7oxPp1TQIsjoK+PwxGd1miNXyWEb
Q7CZqfrGKFGWd4LcznkZrI4N0To7KtCM62QZivL3SYyWGcSJYwQ/hos9sfvt7ffL
jN0KtMlB7p8kwGANZmEAV4bDRtRdOGKdmko0SLjMZbGPm+3y/Vyzr4WbyMgAV1KZ
pN2+n4c54NXYD7sRYE2zRqWm8GgwMES9fQCY1dJz70Oawsuqsy68iQw9/brbi83z
7yoK89wBgkH9X4Oe6xGEZ3sOKQKV7HmVnvCKIGzmSRElWi7JfzivtF3DgGYm4Epb
o0Tr5HHJ/gIpM5Lh99SF25j8X7X5HtpkVIUg4cfNOqj0kNkFbDJFJWb67UaEgikQ
oOezZI7tqG+gXRcJhEPo4XyloVYVJoo3U9TQLAezqMVLi2mMwLsK5JbVh8kDOMZw
8XHNURngisRtV7PGGBIFjxZbZSFAZEDDcUNXehACIefqNzvinS2JfFQRHK/JUa+I
qv2d+mDjewXY+G/4n20O1rqr3I02YYotHhxvpbwiDGTwtoZRQpsUpu1fr2EOt46x
Pp3uQYmqiirCPLM1PzAHbhtOe/DBPYEqF8/slqWVonkBoFchxaXzZ7g5jvtg597Z
bX79bh+pFcIpwR0cPvhOLjmLGFR2XzD7ZuvRlvSr5fa+iv7mMRlNhUJAVj7SaFYY
4CapIA2EakV9MMvyB9fJZjrws2SK88hOx3JTbinuhlyGFh6akxXJ32WiCrzmjkes
JwTQEsdd6O42dBAfP/UW/LLtbfae3ldnRYQUDmGjGZns4Sqlaf3WgIwtFPxyTFjg
di5MxjRrDpXt5c3fsAxhYtN6IGoPMsqB/sa5XOBvhmNaIoL6cKuMafP/ubR6lAd5
uIYutXRcZS1XX4b6fSVsVrnVAzZQOu8RFMUps5PFxPVzcFS7Ks+VhXDJxVtLctSd
i5mRrDML3D8lOjYSR+fPW4i8oz0ok9Ai7yPcYNVyLa0tkfhI108MJGX9+Q23o/IA
VChAA2f47CqI71ItNmM5m7kArTx4l9Nmqp7GSlFDG3tvIBVY6UZNAaMBMnnlq8hZ
oQE6NjoR0wrtglS+ZIPghFagKMY44pjYgo0BaDCxmSUCoeLf9gkL4eQfmE6GHxBz
DWBHctbNQnKFtO4eBUgKI0xR253v9UuIT/BWf279nfuxwBfLrW7of2EO7ML4PR/S
5MeszoRFbJWB0yl50u5TJrvzHY5YN1R1Z2PMZTHYkq95vNmljOYv2J8Tuf3PUaGg
bMG/1JnUYqM59kcqUmzCUh1RZTsQ4mWhSavtyx/oDdc5f5mJaX3V9QAo4rm5Xlxo
Az/wPXVO/5wbiy2j8lvOLCSU0BDvm9JrUBD/cvmJaRxCXzH5KgE4G/cazY9/O544
BIoTx58R5W4y4FwRsr3GUzHeTlf0VJZ9g5lSAeAX0ROosBD4GejA0Edb2ohoEv3W
CXxwlhK9M5TsipwvB2MbNL/IK2ao12eu090hkKiNwf0/Dmr7CcOTdHj9+i2J0oG3
fm/p0xIFqkGChiXvu3glCK2wv0/0yv0BH9lywMesDNt93HUWhe6nw2zG7SMoyINC
2D1U8KtEYULUzViibCHXHkZBX0bYWPTOzLurycP9WeHDuVVxZPSTc45ibdt9Ej0+
SGARaRzz/+dGUlrF5qQE62uIHL0SnHX4rZBYX1Yk0wVoerRHjeWpWSEOzspO1cGD
j+Mc/BbKLc6uls1CHYVIuBxnt/1h8aElUdbEbGYrf0wE/6mxDLHz6kOV7edhnGl3
SfRrL7WShPtuvFj/+XyqITFZuiAt611ze8YvDEPVNfeJqcRyqqIFDjJw/hi/6pdS
rGqG+ue265QpdEfv9LYJymr97CsFblAdwDsT7XHAcgbngAt3657nghbt/Wni7IrF
z7QZXP1lsgtcmf0zocwmwMzf2BTltpm3qVu3Mvy+itgxY77x8cfrAAbUnK4/FzO2
DC4hQcYB9A54JwuY5NgsdYnnpMpKuILX3OqRRGv6dXpqCoWaDmDJh100wyUWQL6Q
i0whcNckLlDAKVTn8dMKomh/xDZ4v7Z1oTbS3OiWICl5Uf1VgNGGwraiBUP3CEHK
SyCczVFG/7U89gU08NNgf+KziNYm3VToBaH63FQIR0BTBDnPpQM0WiNmSPocqDIu
sx5tZgJUR+218WsmfRET/8qE5Tk1wh2O+YHYCVo/3Q9oCXu+XLiOtfPHvZGs0RlV
406d5g7IHQgffaEq4wpJain2TXmDyq3o5H8fAI8WcVj6V9jJmEhkg5XK1jf5UJAh
GDsah4llNaBMyPh2EF+kbZffnuz/AiD2UHkKd1ZZo3BHxyChZ7/EglhT3A9d7dRg
XbtDfkcnE5AJhUuE3SMfSdHrH2l2KlZye3WZ46VDPKQkWsQXEIcwZlVEbCAawQsD
/KL9FVmqyFxLa3KIke+IivyXI+Y1iiGNr/A99ef/bduQ2F2OTTKLXbm2BXYmGs9Y
VK3WV3/2orPNU3f00KqXsgekNUOn8yHcKkvu6TwkzxdorucuFKmCMgBNyuAa0EFz
SAusYVmn89tWPrXYcFtbVVwAiwJ/kz8WrfhCCxT1/dnzP3Onp3AagFdycw/SzUsV
gSUrKkD1+hx2Mgk03mr/m2De7bwqmAGBHkDy8BwhybatUx8mNN34scKmQRgxlBym
U3GRb+un+WKEYdRLZ7KROF9Vhr9tFLn4VY0vWh6dh2G1Y9TeJfj6ZAc5pg0Lxbf9
Ppr+qTP6kkwaUs2ExLY20nLpPPgqr8BRbm8qTET/Vlcq+mlj1fXccEVGWMMM4FUt
jgnDZu36HVFW2bph7NWyJNn1BzIauvHuX7g3JRPFi5HJQhkbfFMiwrDva/Z7h1Yy
8Qx6SomWBBYrS+mdeoUXcY6v04Cu5XmuclDjvdDGc7fjLcZD9DGgFaWlF3gw3YH1
H+w0R9hbeOd9+g1NovQuqifgAgRddVyFuBTD59wRUrIV5cNMr917jzGqqBBMUUjY
vXPjMPHC4hf/+pNT5zQnQYH8nRnX4GtMtS/N/1Fvo/sdncV6m4h2I8f7oqTOpLe6
bVrp5ouzx/geipU2xX3aZghKUMSxSLTwwZSS6URZmeFdDRKpan7uyn/qWpbAUZv5
1DhLKD9mY2SQT4K5IyK8lpV9cYm+h0cIP3QSpAJNpzRLXLJBfbp3nqsE742gU+wS
9WJbS0qGQwqk40wJJUZUyfpNnxr260lqKraDZfIJ1nRDACrDUcEQgQQYqNJWtgKa
KSVpOvGKPNadY4byAO8ZDl9mhYhHe3Qn/SHWcUow1VgUNsPvoYMWXSPPiPpflasU
M40NgyEbyX0WH9WfT/VzohuG3m3UD12QRjLbE13pJeTRbUIf1dMDrSIr56aOq3VY
SOIhhBkqtgB/XzeL0LitjKmI0KTap1ToTa4h/LfjwL4kI37NSwBituOQnn8F5xvk
FH61aJLos7PCjThn+0luGls/Y/FzcOP5r0Wo+zEzOyhaVTLesXruaEto1TFua0Tv
GNI+P3ojpRngJg8iWWBR1OKL2tCk3vXfCymV0Dix2mH/CQ2fRI5O3K3YAxN/6EWb
YGXqAOD7RPOtUNcNWJHHkCQdzB0mFUGFyfVtEFI+zithk1YRrUTAqLe533WPXfn7
Hui08aYDs13gdmAuS7LFBtws3bk0G6PQ2pGX8PPojXcU1s/GFItU1/8gzD9Ec8PE
ppVuMPgtCgPcl+ocb8+odG5aaZH+1drrNFhbVp4ke5WfldIs4CsJEOAUNcCE/leN
nWdNQis8mXDnEO+CpvnofZt7sXzfiCDUuV1WvwVhxA5Ae8AxgmtLw6Wdy1JTGfQ0
Z6i9nXyTosRWZJTXrGGM5hPbbDF9dMjdCeytIzYNM7p2ashkFOAQHhFGSrWYlgyc
aj0KxAN5DQiMd4CwEp4R/4qoQMCWYbbiKAYhRxON4qDPiBgZZJ5UtHk0MsZoWqqu
5zZxoGWDq2HGsWv1cqf33Tto4o5tFR/Ir9OX5NukosmVQcA2uuSpYcdW9PwKI6yL
jGqoLCHaeiqqVYEaPA/gJ+E/hJURe2MJpW5N3uaQmKWEBCLuEWRAXJTL1WdGgvRM
5LoySK/rCbTfmB+YHf93rBQ1UDcpkm8/6bC7Y1jsmkRQVq95EfBCAUyoyJbw1W3v
RYhyuLnIlylnW5J+YByWeH/qXXnJiRzGpscoCLVeNGJuPjsL2hNoOd2WxrCi3WzQ
fAmTd+nnW93Q/eWJM9qMFb54/ID/gXgZ8HiO0XEZyNtrPT2UE/7zDpsdhWDNs5W+
oYiUZHKYJEaCUqhsIDZvGkKm528eiObeiS6tkg2U7qz4uuOLHJomqX4Oq9vjfzsE
J4OievpF+tiJigv9vyh0DCViy98Ax+PwhNQcrG21TsFbWGVpkHpnxJm0bcNXH/VO
cj9mF9sRm4ffwSmjuk/Bl2/5+U9vlT43MQw/loNQ6ZwWdTvqX9e7DhJ+56GzjbMQ
zGqOOTZleKdJuQjaGIILOsyVysRVe4bdAZjhv7gfemGqDZGNqRA6uMpkezKkNQdc
qGAQCeufE4bTiPdoYnkWfZJhpapiMqQrgqTs2kZ9pRa+KM9XDXhD48KBFKTz07w9
pwkg0PFpUd+DW6nsb5Dc8hMkRN8njzkUJlsIgjGw3xO1WdCgsMdKxsuedqwQ6+BP
RnioWh/A9G/UnCCWCfsENF3YK3nJMl3UAIJLtZuYs8DcZRYkVuOSeOzGH7TW0IO0
sjS1eRB4YVd/rBzqp7hze/nK3pB292FRLdT1tE82ic3PvAbn1tvBFVvHvHRbD6x2
OG7l03hjLDpkxM66Vyw7rwPJxzknF8io+M6VcAmIVd9pXNWPgRwEU90yR4mulsL/
4FdP72FQ+9uT1bBJ2Y95ePa3se56VUQtJYqQSFyiHBoYGsqALJ5GB/KsMBhaM+Fm
e1l2vibJhDD74l927szz+NCrU+aGfSk07a6pX+fnsW4Xyk3fJHHOZerc8scQjp7F
XCmxM+nJ9/eLSb2e633zGz8jd/+xEGqVoo+yQFyzakLxxm8Y53zQzZ4u5ci5B0J7
DgPKEav8T4D86ztpKuHeTdtMoyzGMpFfUNe6d0hvCdkB/bYeCTC3+YZUtLmADC7V
HKid4TbIF0frMaiS27Ffce/Tah4O+3/DpV8eK/tsXtTX2k1I1LeSxUYoRCuLl7My
YPj8htu5V9RAgE6A9tgMv+gGWATbZWyXsEGn9MyHTxbgNuOhGqBA3E7DytWgaaB2
PnYFiPEeNHfT9+QpU0I9FUnDN7/HQyWxNlrh0D/n/GyRK8T9Yjtvtd+ElkWGgdKk
KpYN9iYn4aSsEizI0KHUJsHkQUfiBl+psESQ3QUAWeVkRjMmukZVmiAvYsSy7/Ck
B4B2UOtL32eONZGpTRVsg5uztNdYo8YOtHvKWehk9G+sPZ7Ql0cVRMdiJ9RCZrvS
8JajbxjqmAEbZK/Kmr1RNDUZO0IVOud9WiFlxWw4S8oSngE22PpVt13xCdNkTtpP
KE3u+d3czMShz0XmwwjXj9TrSIgVH334Gu70zJpE3kvCrk4WvLO0/dwNtT1XcZKN
jDDsc+Yz4x3nU3YShw0eENiNd0B+V2SzBYDypcaKlfAQqHfSeDOcEh72+5SbxXUZ
LLhzWlS8c5+5SkbnL6FGyZGYwqCL1/oDgZNw5CA57iaQM/nrwnJ8bdnZbt2nt92K
zOZX3UoS9GyAAxU4eWyxt28AwG4yv6OYAwcDHmyl4qnnk+/4PLHVNCteF6qd04/7
aRZdpgpg8QNSNsivJiNnl56Vy844j3fpNqpJxLM3CVRjFLL0nPPkSu4gFMsDVO8c
cNHvlAIhA4wBSaHUP8sC9QDt8fi2KMeOCZMV04Zawru1KtrLkZOeoOQUI7RntSLe
E/Bssk7P+4GeRql43lVTDELAX3Coczc3xGAzO7EHQmtWLN+60RT+FZqMlfuO1Mx7
s0bQ3P+wl4zHe4NVnq/LEi08/F3uima9lhXfkLf1sEEGTQtDpgnl26wLk9eMvNAq
o1ROrw7QgYVIReLiJ+8zlkGNo7GUAKhmiqGjWHFILUoXeeSpjycUN7K/KTPiR3lK
HOKNWB0UvVdTAj60ZdrgTFlF5QuNxFZN+ztgAkmjSu5+GGpCEwvQPrx2/001UIDd
GPeeZLSxVhk9qPOqhoqz3q4fBIonF8tSJizHC6igt4ce3/0jDnZdXT/qvM0zzt4h
`protect END_PROTECTED
