`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0M9hq/Qv4C5lLcE0Yz+tuud78cYKpV9gh80RwDsd4JGFUQwJp7RqH+/IWp8eYGWG
nzne/AUW2yqZf2qklmfx6PgAj30zj17KPqqsm5L5+DqWp0vlv/UGy5K8o2FUX31Y
f8lMbZ76mAoPDGEuwBlMaNmHqDkuddZWfzjd+gjvyTgNrIUG/sklpHJBuJHOL0uX
8RCkp+VmTJIxRS2+ht1PtNYLxjjI+Dxla71AjVEuHpsp+vSZC9fXacqJo2rpDjVl
q2LvZkq8NJ2Y758zk+0aw3EJBJxjGwrJPa7ciDXIuqvdKhLso57qHcNz8eOdijTY
URzdzD3IQpKl3pLmsrIah1T6aQQs3CT+NKNzsKq1RQaMd9LJIUKdAzyyHdlA7ArC
cb1dzRa9SwDBdJS5GG+uGavfdrzRrTivA84iuzfN7ZmOEvZhkZD4+aUzgMmz80vH
i0BZbiI8gMCgvjFINgSEynbAZYqNDyCOXl2YzXWmZOQGd22YrOdtpPbJ15PDj+6/
t+TnzIlx/L5lMwA/XgICdOlN0XxBzfZdDfOp6Q2NiHL8wF/Wj8/FMvjP1QBEQS0X
EW4ED0Tk2SmLZLITJ3S209YTKWLRTLNnWckn3rQdIRguWLT3592d2or2a1xLWMKt
BsiBzmDn2d1wsnm31tftzYucnZ8LJ5YXRNa3RoWNa4abnhqZMSbE9FPuiBYqG9y/
UEUzhb69RfC9p2mfigpWM621E2cTXDQXUpTjoSucVAeWxE+ElahR2PtblcOd+1Ja
zm2vZ5JaG7Q5Zjj4Ns68vFljHdNdVthUGpowv1AU9guL3ga6aaPPuHQeVxl+o3jT
h2eLZwq9B/Ovx7wf163yqkfzgkE2p6y2mrjx4hASm1U7HSBOfz/SlTNhSi9WRGk2
AhB2t88atXRMnA4dMD0e0rm1syXtdfamPFs+bV2L3hVdwjZiGvBmylfs0C0ZtpfT
`protect END_PROTECTED
