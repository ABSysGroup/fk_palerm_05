`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a36BYuAi5+60z348t5s7N5hZsGXr9+Dg71d3NwpzqjuXsLQ//Ypoj7J53n/L8E6R
8rDTt/7kZjKFuYz0gpqQL0lhn63eYRC02p/a6nTQcYfakHkhlGNBi2BkACxF3xeP
zRHK5Qq3yUpp9colO0nySzQ+7fAI0+5pPkk+DelDggyvqUlfc8kMKFhQSMUrFv41
J4Y6EuWCrDZfhIL8Fy09Kx1eBbjW9fdyAGTM9dMAN9VNvziro6kKRXzORewJwQEv
JX1GA7EfEnd5XS2Cs5G17g==
`protect END_PROTECTED
