`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m/gudMfncX1R3n+pifWHgGnZ1+9H9oCm1uBLP2YmbtFRNgm4AzVMD5XKASF8LnZC
K6AUIu82VG/Ne39Ah6rCmIyGCTFxaT+DLN2z4E9ljCQ0eNkdLsEKPiawcJB8iqi3
wo24jrzHspk5fIRL7jpdNNpT71OssMWnAc+41OudPgbbvDyKCgt0qHaAZGE6PVYr
wHGiBQihqxQcissF3HVmmbw6XtruPtGEz/uMbaUyDB94VbymthbrN4rccanv4TPJ
QCtbjK8I5iq6n9pyzUBa6pmTRLyIpuz2/nqdgH5dA7lER3TBRdimzSonGieu6yFe
rAYbVdsPgxuZU8iF7w9JH2IWMwAgp6dq0PAWH2x98/Chjm0VUaCwx0GedBDSuW2K
2ius2f0gPXTBXniVWUbyyG3SK0VG6r086/QtsixsrD1qwHbKUHyXoH95jYF8SwAR
vjE1Mq6UMTzVvcbGk4O36/qP0EaeNvdebFYbI7s5y0uIxMEan6+u5IYNvd651Zwk
C35sksbpZ8YzhYKOTRAy4LbC+zEVQlIX8+YLiW6BpeU43ULXH2I8gg7gGa5Ciuu7
sG5/xzPRX7rClggG55TbZM8OpNsHFw7e6oXJhJKIkBUMt2xUpIOj5TJV7IOunIdC
5UVcehEDtC2+Gf55xhPgtL3GLMa4X6/KQR2PAFzhC8tY7jjP3qMydpABYrVQWnMm
IHO0ptIp9h8eKp+xrFGb78DvBrZFAjKjNz7++yAi6rZ+IqbWTC04iTD0TQO5qnr6
V6BmuZVDvQgLVpICwjJEvF3n4mVh9YYNULcriOKFCQC4mWaXXh7Jzdq6AGdt5mb9
U7J89RNxElwXqFJf+87508SzDjkMohqsHq4M7dXGAH2KIctxIn77tVY/nJrFtXg1
qlsXUwNWN5wldVGdKDaZKiQfbGGreLJdQYtdD2IURb4Cqfj4UFD4gTgjt677dWel
uN4HZsqtvwdRvKjPO0gzsvffLFEqpHom+N8nTf7rN8mrQCF1rJV37LvsgK0DmJHw
RncKmtnGdMZlt2dMOa+YRN7DimQWIRqbqDmfbvDnqrIHayntwjXZxAwb8Z9MJvrJ
nIHezrmH925RkLWKR46dLCXB40FFrkvDRcmL5RPZSor6TPtIKgAsMJZhRJL2wmyR
amZT4GAVrAZu4P6f58AqiDW10mYYecZXTZoL34LWZm/miM0sUBN5FehViicAQmVE
NGj7OBMwbh72tU548s6Bo8+LH3VM5RLXMujABnhMdnnKyvvvUBmZ/kKQwvP70YRg
UyhYwuUQYjjloSg9y6i2/q+mn8ULRSBYM79HxUjMOrC55BUvbPeoulQSXvInaPHv
j4zodaGu1t3YhZNKfJHGDo4O9GVBczNbI5liKMa6N5c8/YZGRdawSg4Ywu/UKZV7
mb+MJqFwPzZu2nFk56WC953lmGrVCTKbEQuuLB8kV54KK6KD3/h2wTAN7JYAx6P0
udPyMLc8zjQYNhz4kI/vfW6P5L6FEgt2w6VTYglVe89pIQelvEM+gK65+tTwfuM4
Hy6H+3VvHIoxHmeKa5KczjnRCMUc0EaJhxH9i91MuMioS4/owQbskQdKcIDdrzix
lpJPon51tzSlgfwQM7tvvOxlcAb3g6YIXfoIjmQLl9MtEgec1WCqA9/Y3+ehWdsQ
rvQdkHfgKmvk/vmEl+Th4vtBJEsZsKk77bc12SNz5sBH8FonO4hUNeNDMX3jjUc5
hMLcjVZkPsC9m4AUzU0XuDIuYPqKjMwUnU35BRYcOQe6zX6CWdLiRe16Kbf2n6od
PQaTsbHYYEY7rIjHkb5VdUmGH9YhWXFTPs+M74mxTEgnpz5Hg6UwYejTkFzfoh6D
ZScyfVhxnqFDc93vFZq881njn5HxoMP8JZ+gTf6JdsON5KIYeMVa63hWISPmVWlk
bmCsOXGvupu3U5cUVyLdvhS4pdBAvokGupxWfgMLdws6XQ4RuVSLFeiMgi2LchPH
1kDZPPyxaF3tpm95suBqaNp4IU0EyNA8AW6cTBpZBkikIWIaTgBv+leU8IOIJcH4
5hmft7tIDMPrXkSpVmbeyrM0Qag//ZO3bnKR26On1XLF0wexe0EpuKQggHxN/38x
v4xzJU+JS7R0GZavUNv/Oi1pR/KNjnjiMcJL5SONaq7dqrhC9KeJAeubyK8N1BfK
8b0LJJxUJZ1x38SQh0JzhbVVUmet5VzTZkz1vLx2vQ8kHl/tpXwSKR/bt7CUVvfX
St10fQW5eLHEiUHhDEHhmyZI6V+ldNVBOcw+1v8YDiag9+GGK4sVFM5oiqvTRu7a
6/B71c6fKxnpy5CnlGNtwMIGVFSsmU1Gev7TCzFUtSOqDMEdBV6XF912bUFODrhU
laFvlNIA1mg9qq180XRclE7UilRWxgyuC9dFIMog73JyNnc5u3WeMCy5+kT8dOsG
+9nl6hnKKebG8UDny7qDQsx+3w0ZKSnfcBCS6ABEGy+jNml74nnbBkn6qfo3aFlH
QXTY8ExBcDxWVdRXjfFsyTdCUocIw92U3FNex+j5JNz0B1PW3itkRlWs3n8KC9um
flk/G7m9RVZIs3U6Lzv3Dmkg/ZIB9fybw9PIHaPPdojTbC8LoQXyMCa5Hm2ekHMs
qrZqQPx6u8ygW1m5tx7ut4NgTwCVkZ+aQXvR2AMNQGZGOR9C/eqgvCgdMg3thG2i
P8XDH5bKquibUUQJAI9apewdDq2etuTWauGNEaeHTmAiUYZzfZAIMR/eIAxZbpaH
LTtKC1DtKtWbvehFzhlUACYK66rBjVj/SQi/aDMzGNyhgJVYktwhj99AMOjyYjJY
xoWphqrXRQ8nw/ywbB1ndQXh7VG5EaAzxnQDHd3EWqs6TTU+qffbwIsA32hMgUqL
csCv8NZFAL3Wo3DavtEtMIFLLmwvUFZgFMonzu9y8Wybl4c9f1tJ1iz0e8YK3/d2
XyeM2paVJqpQ8igjsjnUIO4hTJ/Ib2I6ljeDBzPtAcRFlLbqEhQkKRItxPdWjJxK
B+JSvQguFJQn6UkFKhze5fbAb9yQ5Gt7/DVQapdbwKc=
`protect END_PROTECTED
