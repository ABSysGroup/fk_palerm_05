`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MiWWtRa/54SO5dHJvRoiN0itkM9EpKWXKk6UeQSTxOj9uO1RFHvWDrT8730S4p8y
WVoBSGl6vERWHcdcg4wzWBoygXqKtiCUCwTNA5sAqXuS9kiKEy8+bjWGTFg5JLoZ
Uq0QpY6/7Jw8JNsrq2xXZ4gOvYL3WF1vFw4e6uNo8jSfp2V4DsVdsjf5XTYjJX2A
13PCvgAfwdN8YFQDveAtudlrmzH3DBs1Rp5UkbiikHo5cQ2usdM8R23EJVU3X0bF
5j+jL/3pJyvc+3ojpMPWyfQxW1w9+5bYnvjdcxQHkaC46J154hwUe3yO3oLcwMQa
phorV28anQdS3Taw39MtniLWo7pXBzc0PhtLZNiPBo4TEhUiB4alrdVSymm7oKiM
kWVJzjAEYk0pT2yC5XZGaMJKdNThTq0P0O7wHRsVVFY=
`protect END_PROTECTED
