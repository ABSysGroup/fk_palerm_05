`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yuxJPW/zrMqQVZ1Xb/OVwPPo/hvjPAyAlO2jwQEM/GTNSaVgU8zemMrjNKwom1hq
KIzd7Y902gg5BUXI15YtKI7j5Yw4oMj3cnJC1LTPkm99IkFgREYXyxmpfH4zATaj
QoM5PWYjaGGeFPxBnS1ixVcjZYfurMvqdmBMdgBxvv3vzWYwtpaghfnJP87ksCvp
q/mtSK424Y24YFLOTVxqzWIzGKK6KQRBg6KrqUKgDiT8W0TBOBdcHRKfWgtj6lz8
zut/ezmhYAjIBmzZSvTcTKM8mXOJLygekJLGtVtLzhSRVkAi5tIs8ahPYHYmqxVD
CZ6Tdurk2wkBj0jV08EXdKMRo0HopSlZ74at4fzlwBAeOZJ5htVw4qzTEvSWdBxy
lOKNpN0875LmRHMafcslnWzkSb5CNLzJC2ip6+RexQl9JGP9WftdGwO3Q7nM3wzY
`protect END_PROTECTED
