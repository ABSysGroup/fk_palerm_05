`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VHDHIc51rCeBlsmJ2bPhZ+izqIniJ5RCKJQk+3XH2FJnM+kzVFlvK3watDsPRRcV
5pX+1DULfUqOpsbNTBCVdyAGajApXJG1E2N7PERwpU+2Fcjf4DTxIWk2wSljd66U
5l7lgjv2g35WPdDRcqq69baKzUuYug4v1nRcOYpqNyxd4NZBqg1uvE24ktpTmqzL
Ogs4o5oQAmCY/GwzpCZljXd8T3qsPRBIuFjA1GnM55oNL2XBMFKDM/LHnjyJ/3P/
fRavYAP2q9PP4yfECH2/ofSdLs6ffEtGwBSa+6aGXI3ncyCqLAJ6iNg5pnk+7Ut/
CzBr5U1/sK3oDIrjKZE0X4+FE9EAwJ1jUzQXW5ZOCpYDfXQZDJyxK31buLtJdVHR
g6BPUO/WGkuM4HfJZP/tbHysLMVhz7hutXVfDAm5Sxlbaqni8LRuL3s59SPi0w7T
FSobo6BFdxQO/RsRMPKaYLQf4BgoATWST129VbyqDOuVoXcWrzoDfftKumWEr2ZQ
j+EGrUetu1UKnmxND8hhMV+FImIyvVrGMO+27tmM10RYaDUA1MTeTZIAtMsc3s2T
VVQhto5N82HrhCPLkHT4ICtTpp5WLjopFil6VYWtjFC/IVMmCr+8KJ1dQXxs8qqS
jYyfZp9D1msHOTD9lvCaRsRZs/+eevprVrVtudXAON5ZuTkC+tSHhw0j/tuovhH3
HBdi151H4Ncj5dPw6yoV5w==
`protect END_PROTECTED
