`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1r8UOj+jXIiQrHG6av2mvCyJIoQNfSw533T5eHjZaYfoaiGUpQpMu2DLucQK4O56
+c+JV0hcc+NgUSYWi9w9ZHvhzTft3w3HpeoaCQecwe6jJXGRSJsEBV2GF79VBpJ/
NmrKSYpjQreW7yGDpN6sgE/j0PGFYIBmx3daKNT5fh2Sn4Ul0ac3KAyjxTfTbLS4
QBEOnhtv+4KSJjN2bYn8uWGpD2s9TJrzY+HXABTu8Dzel5DKOqPxLQ34lfoz/Srn
JTZIaNfNUm8iQPtUDJF7lQ6t1YxYh0wyHSrcCQ9J1oxV3RF4eS++yx9s4hBr728U
203vPoUBEs/cReRiTbqb1rjNG6ex0RmWTVpG+pYj6h0qOGKIkFHlPSCPBb5J0+fn
6wEEL+r+wNb4N8GqzHfluBAMpkMSyTm3YZjAH83nYL9dxhAt++yLOfYsK8FYZpjY
IlHPgQw4/AQRM2uOoE7NPGwOzc7/xzV2d7VhCHzqgGMwYGOpU6Isb50aFlWNyTPH
FGb1RWkXUXtItF8C1t7g3agivqO7M7c1hrdq5Z7sqDVO51AHE84HCr58sW5s+22n
bqz3A46bt6HK1X8ZSqXwz3DtLnwurlijSblaNXjj/B5SBzAGgSNAj9iAH1PlkYbY
Fjrf6tkySFz+xJlLPy/0LbJpYPIIhgrbU7fi+rh7pJRXBuPWn6qdrUU7ccBp3IVG
MWwR9dbPW8wnP/ZJB/wIswMnhrcx+Ay3WQgAD34+5rEZ5DppspUKnaB/6nyivkqe
oIs5d1w3jhiLwGBPJB+7umTudRbcv6cZrS1WqakA43fs1PnhKyeuI/eaq+MqNjhR
ODOQfb+hHuucxEoFxFQdOWKzhVkgLSevbHgrm47xArzFe+AO3EZEOKqVstQsUJS5
DROfmlfSFUWhMub+2ku8SoTPgZM245eqU+hKxJ/sNljeGCaKWRSLpq2OBlRnSonp
e1aQNkHCcqZRxaZFxJZin7QDTbuTeq3UPsFmBS3L7zM/KYPvy2krUjYOEbDZg1zl
CNtY5RYOVHx7UHc4Lq9937zMVV2ToyGbP6r3PYYRmdYTl116nGT1C5jI9s9ptKSJ
AztpX1F5aULARn9N5DZcddokRNQ3eAlD0Botgoc+ATe7NlZnurPoD32QgM262NVz
xMhYrKWqImP+E3ptYRG1rfJbSp/znOMFUR9utZDA4HJ9jdvYb5+wSJ5hsEyIXCSv
iTPPhoxHimTJEmzs9iDNb6cqTwNJtrwVnQZVdRPc0916bib1rdspJJ5wL9R+72Q0
kgf5wpV7lTdJLh2ijZ15tC3V6bypmeg3FZZFoRJrWgEaaG7rT5IMi8QzAnADeNin
yZPbAKjSJFqcxCVyQFHI37bUrVLFI6DDA4Tr3di/qUH2nSXukWguBbCAg5GFVbG/
2qKGNEneFaEtWfSILTzYG/kn/ZoD9bF8VjBllw9SSW9T1hTg8Kyl+quPpeYXJxwN
VmW9mmNkTd2JXLcn0MT3RaiGH85A65ohx8O9u+P15aVNOBxNMY7mvUc+ysC5kCIH
MopXTd4NrpskwdCL+6SwwPGIaaxo5ZYcQ2gqwRZUViy/UDO5ye9KfB1zQkVkXOGH
Tnh6dia+FkMOcjvpdztMyz3lct18ljH51SNfJvQ521jE6iu+wwWXVZuNjtJMt19o
vvreFkaC3U0TIIOBmMSoiuyWhC2FV4jnMiXYfe2i1/S7uRW21lhsYqEJiQ/rgXgX
CTvrhw+bn/eGLeJ7Wx0t0We7xHZZ/DW3MEWyjNiYeiHCJmjZWK64cDo46kf+vusc
PfJ9YgSXboNlWKk7FKf1MNh/Izzjsxg0ZpHHt+l2zoyqX+9lgB5S9K1trreh6kH2
oeMi+cU8/XiDUrtU6JZlbA==
`protect END_PROTECTED
