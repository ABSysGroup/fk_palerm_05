`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zB/Yvb9ILXTUhB95SLa2zxgQmA1SZtEIiAORm7CE87SD3ITV1x2A4z3p3trsf37q
ioMFv6GLTkF+WTcsgX+rMAgv0DrQ8bO7Jr+Se4wHpkQ1cggfh8qfFZxNmAY8PQSL
FKOYp62VwNHEmaGays45yRsWyrSBuYP33pKQaFvdxuQ7y9gEW84LYiLV1biG6A5R
Tr8wGHpgWrIvKP0qDbOuuZ3SfDrJi392e1oui0RJljAmRgjQPO56FjDvC/71eyWo
vQ/nU0h1w69kOGQfll0mePeSGknH7mMBtVZjvZAKh2WFaOKAv2XU/uuG+OvmvdnM
dVBk2Jcdy1Jrz9gS49uJJHR6egbpIS0WxUy1WsNCtHLYQbHSorsHt6qznKM+CfeC
77En7vI9y42Lm0z0fC4+ElcC6iEW2jCQLBLGIDFucExpnY/70LbrEQ9IzX+n49Y9
3K8sFUiPNXEvmrjuy+WN6uBMPbr82sPajSgbAzu6jKv3JeWCpzABHu0B1jS/iGVH
wMS++qfzazd3/Mjrg/L6xVhyvR6oVwf/C96f0bWRfvnGMvSo9cwrW1w788RXEu55
BJg1YHwt13FzaprvPpm8vYC4ffvnDxGQ4WfX7hGAFkSvaxjyEKYkVeSdVpz0nTcK
8Nj3PlxYxSSe50d1eyslaxzf3m1JgrtZcVCs7yyPSIC1Q0NzzLNAG9Oe3/1kef5p
AvExuqG7WkBmjT02ahP1b3PB/yFFYrKfTwvTtkg/H2KOOBPacCV+lQJ/hTuqFuvx
JgaHSvEQRvs86pDYWTJs5X5wtwaELRxu5WmhccLkEfGLA7tWE9mjcaksPuQviD39
p6JspgKlM9VLVOwivIwZRKvjAP/n1Ms9cbXfThWI6ncYWTGzsx8YxvAWp24w1zET
+vuQxhQalL5IMZ9cgl18Irj5tsrOmnYJZG5P7iTCgJZA59Su0skEXQstMI3XKWHd
2CRC6iOfeYrDcx72r8AMPTT0kI5KTTd4rQKjGbsN70gwG3UU8bTFtMiL+dst3PSs
qht0GMfvvU6LWYVN7TU5fG+4CW4nFI/KzSTs11JgKMYircfWPT3HDWl4tK+lNOco
Yjw5XoAacL7KtnblDIhaZ+PU2sxY1FRz+m/0gvJj3ypLUlwbxs/05vgC/rFKhaQC
+gP0CZFof4OQnHGQ4LdmX7DrOMW/fZyg1DdZpCjuWB14omyfWNDYrOHM7VBgcDuj
G9PG++pcaw6boaEhcq83Rh5HOrd4CMkKTA0B/MWy7UdUt16G26Z0OET+JMwXZVjo
UE4GkFn9qRNfLYKU5ILZZIAtH7zkrMDlDj1ND2i9895hUPWZ9v60ygNfzSa3ux3e
DwjmCwrbDyiKVz4UiCyzSx2T20NnqokDxsJp/RSkoJGEL07sTgBvP94/pNQZZeg/
OlZ7YAUr0YiDNI0p2P6urD+ihp/UST7KHw3Vxo6OOf6kPrnkNFdsUnXb82by5KAk
uA9Vs2U4npLWbSbXBbwrvtYoxoPW91FnBJ8n0ACfUsUFKP1+xHphIXmEuaB7aGbS
+uY3HzmwhVrf2JQaqwyxMJNYF98eIIvFlzZnJbDIK9tPZRBy7MEnpIAXLRTa2U64
5SeW9ziJjyGqozgcBMZMI3O7RejCTD89P3tqcMg7z9USM6TOB99qbIlso8t/yaKf
RfqPbaInSkyt5L0CINmbrl9KY4UwmbfYNpAkbgPEydAldguEOzcTnnfjTwyw4gAK
YHPJe/gSI8uh51MklgaRZZ0VDaMlsSyDscBV1tvUyRTHJOt84NiTSbuKAW0vTn0e
wpG4LJmsoUAT0dpZxRkQUP/hsusWwXPTChLb3LFbMCOkOH+qb7s+RM7Ds0HzZopy
zopQCYzCva1H5bR136AGKRaTtAJrWVmtQ4+7t1bF3vh/3zU3cAPOTZP1zUnjAPKM
aQoj/HD8FdFIBPFG/AuGo1PhlJ9Gfi97Q0HFlLMkADrkJiYAqxct9Zmc2hAK+n9k
jdgkCBK3W/fxmHq+IbnljVED0qz4AwY4Kx58b9+i/oURzwkqw4jaqUu9++e6Rgtw
nGAHL2UqM9ZIdDKUM6FR1OKxu3vU3/gtQiMiw027sCjHBxj6wk6pKFrOgLHL8G8L
tkIJciyjZnGhvv+V5ys6D/tpUkE0t1Jiy2quj+7OPOMoFZl+OFqAEfrFdfBhQUvC
+RjhsZb+xFbEssj+6dkrkviiPrIBquTtYcVKjAXmsaKliUBY0eRXlfPkEyl5hZHB
Wq/rlHc6v8tVWyc4AkNN5DCnOW6Yh28twTUHfZccYTp37Fel+dv2jxoz5MS9YmpE
lSQcwTUKwGZ7JUOdV/pD8szMTE42Sl9m1t228oMqcLdyZz4BhXTSQmWBt+PfsXvz
L0qrsRBIHAMQNNznw9l3c26Qj5XztKddi8iSAnEBruVCaKNLqyVc9tTh40RM54zJ
Y/nOhqsS49Qn3M1RlqFOsKS1YlraV/JoQV8uy6/0xOYBFz2yzimj+3sfgjwaESKb
1bK6XRTIDD9QP9vyy/PSZDAxEzo1RsiJS/Je7ddEirYTSy9kU4dHWIx40lMAK5Rz
BBPxtjpbBzB43WgODEYBvo82BnBON5r/E+yBc+w0BsZLfGtGhKAeo07NrdGEUO9/
d1IB2gzTPEbbUb/7/hKVoNqPJB8eUHUIlhdsOrt+waektH+3jVKtFwMcXuJJQ1eI
f8yvEPQyaKNHBvUkDEG0WGS2MOY4KT9C3sJqNaFdra/haweLTd6YamjhGHlC5Q4E
CWMnkdEaVguul3lcv0/C1pxnpsjqHqo0sGM6F3p/qBlpPKoXeDB7WH7q5qapuz4h
MjVXlApPOXPsgxktL8MZPPoDfIfjlMwkf9iVzhihV5y94pWKj464d8uUT6vA7c1o
E4TxIi2y0BdQiha+S4fXq/I65E9Lcgc3N6E3t3iCd+HfflQ/iJQyCxl4ubX/Qy4g
7825jzpn6rus+rIstlPpR9lJn+7BUZV5GT0D+/LQhhcL4vgR8YIPW9zo5ZpGOan1
7UW9Jg+73GZGgN8/GugbvX8iH+/c3PZQ+V3xTIYqORBIPhidqdvJS1ss/zt7rP6k
0Kq2u4Xi1VPsG+WE3cREc0C23z2XOetUIN30OaKPj3wnqfTkpJq0lMgbT5THYW5l
T2BChEMWG61k+0PBTvj3XEWwOL4j70W1wJwtOUfElDNBfNxHHuoRaDIwX1RRmboG
8u6L4FO3g9LfSwe0qSF2Ax6UzOVCMDdaxLJ4EzX/Mr1iV8bjMK2Bs285H05/Ot0B
kiCDB0WdMuegL8PrVW4jiMz1E6ebrr59mR2n3ynMVOMCHq5CRAOuA1lrM6s09JLf
/2x8V8g54UqIIZfxzPSx49d+/XbP1VtL7izx/lFMClm6UCPBn2Ife0YGgFDpyQK2
ZDiC/eK2WJxBa/xaTD8GN40BgZZL7w2hpXmloXc+rqY4Egol0cLqJDmRDckOs+y/
sglNXlnYAjYlGIRz8qF7Q8zzClrFsr8Xdbuf6nsfnARt1oEP04olujXmq032Anda
4oJS8ZGEdFDAV2kJwuEG7q/Tslp14zx5td5xluYsXFdiqyMYZ5iq6rPGmiXA/O8G
Ot5HRfGelaz3urQyCAyCeSCYkhnLv/SJ9piuycvFfqWoS5UslwvVR4lrGOLlrO2L
DLFPnVL3igQK4Yh+r10KS6vy5D9KPRiP8JBO/8ibarNf2rX0bgAQ8Wd/6t4yy98R
v9DYvASYyqm3ijS/V0FBt8nTnJmWYGoziqetgyYG7Nub9cbRGqXBVyZ/bDFKvZuS
RsMx/dKTEyAr0aISJ31tsHfw9le14j5zY08HzTiPKGDws7rkLk6tfuwY3BwN5KX2
5ba43UOtSWnNdRjXNeTj8BimtEGRPS4GcY77VSbVCWAkma2XVwx4oI76xhdytbu9
hEXjDqT/U1WaRLnuWonpQKTkKgWhcTS1fhecTEnrYk8AIt5+mZaQy3Z1GfUhBVh0
JTM16bAyIo859Qu/HK5+YHpmfGpgcnOaD3JEOw443y2mYqaQQaIVNJTr53YQw38c
cYSNsmqEuI0pczmyL1YIzQoMjnKHORmU6CftIJHRCQJWUlRShmpIParJ7WaqN5Ep
64WVA8sVO+xVHHJlY7uLJibAOV5q0+N2Uvv1gjlZPwoxSR9zEyaYPrntqz2+qy2y
kfNT9Ag2ZT7gjtxoKYTnP+rMx2ntBlV0WSiIxf1QNpF9p+ow1fdpZrmew9Sjc+92
cxrglNx6UHUTRj5AvENQc9VQPlb6xrgccEfmfBfRnPyt3zmKboUTxT+/gYA7ZMUQ
qXVG/YTHO7QMgRz5mdByWOyKPRm7mHoUukAoh9wY8xrhp+pPMfCGCAjMMmEKKR5N
Ee2Sc6Tzcql0jFCR6uDietGqvRBHbTn06wmWytGwU+wCkgxY3UiBF2dGGsZO9tUh
mdESwumgu++L86zCxi8sYhww8ixO/q4OwmIFFqt3gM29LRl0DCyPJ7SjCyAFQVRc
aD0bbWf1Oeci1r1WSJMsv7jr2nTp5iudt9ue7/Wh5M6ZKT0qig/cCp5Ffu+KcIHo
xwDz2ziGXA0Be2vlhHuuzCnzGhdW1c0ORqZDP5QLMa3N3WrvdGbez7yeIu+fuTcB
R7DjrEGDFWSXiWNgfwke3PRiY+NdxpdZZ4IxshLlAwT1bNzxBCymN01AyMCIZhb/
z/rdRYbv7RA1WpFE4ViOD109CeRbOmN/wi9V0k8lIrZiSr7ds68QCNSi6zkbbUDA
SCICXL9fcfgobUveoWJw7TO3yfsPLCr6C8cFWm5kmnYlw9Q7pQOkB/DYh4CQnpG1
OOPyVVk5qfBrtdC6r5RLtJI8PJuccHePhe63Z52xplNvT8VPxJe6OYcuEUpaZOdW
i8qF6c0ETeZl98ZhdBtciAAY7QKj37K6rqfLS2UmqpzmM6V/KvfJpVixNFnRfN3P
OiAwQUJuUn7XwD3SMOWEgFn5e5vrXxyfvTC+K8MawCgI84EeEK2RpdbkQQCxWCvJ
yaAxULNJgHZik6B3gcErAonjaVSK7qlsO5v7ZRoA7kcJR/CWgAL4LeHn4f0ZbLAX
9FvA7Y6eUykV03ZJLhkStaivzwbKW5nK4KpIVXM7vPPn6eXPI8qy44cFKZeQNnTk
2cDFHZenY04h4/Hj8fuCEVCI2+By0Vkxefy4ApUu9r8LiJfUfFYIRCT8DA0ZAVui
Uh1XoO661Hgr46q4DSxcRpwr/5sEmXhiWoQAKjqER+JtJABBngB2IYPGrSfwu5Al
0BxQKh5daRe9QxEAgiu4rXzHlpG4zmz1Z+6Xh55D7tgaJmL68w/kpbQU3jTp1fut
IW/D4O+7OmFuf5RzXcmCfzB6wCgezCYll3K8y6wsrqwrglMtNFtVu4GCrJJqgymU
bSEccULdBr+8W0LW2UPR200Qq+PXlr+uFMQbomNVwj9Jdo2ImAzlvT2ZbUrAZOOv
ZMA0Vrk+DpBYEQizAHimi5O7dZvwA3w01V3L5OVM+wdFgvSgOvIp/qYr2LAKBmCZ
Rs8L2VAQOdrLeg+T/NL5AYCE3mRvQ27erzWeGig9BCUePOT2hFoED8a2kV/6Wv9T
Gz0VZd31SVRv4BZu0dYgzLa9Cx/1qaxFwGZZvXz8FsfnnEXwgdtpVr1k8Jb4RQGh
8tlBIE2Jw4snhx90cd4jfyEBJ/VQLtH+z+bCG1/zO4FMgrg27LWsgW24mTo5nT7t
4qA6Vl1xTuzCTDWOMIGplTJ4LYW+VuFteWlTGE1FCYWeGqjqMCMwzLQSP/iDEiZF
Vz1MwI3KpyNNBQZytl7Qd1WneXs63BBp6vOS+c7r0ei3EiMUa1LdwqwyaAEB8qNm
8lhUsHiFY2docE+cq7ge8OfjhF6D0G0kIIyBUQC/wYCow1cu830rA6ltVwskY/Ny
RdtntjQodqhLRYmv2zhVCB5vgy638M6fsIv5WTb/RAUfv87pDOIySQoloLvIlCFN
+0lITKrEjVMlP96pIyKCEU5bWXb+w5cuC+ZWVYh83ar5I1HbiN6c4kMjURBUxfx1
sW1Hj+pDcpaEq5UKTmD/EEN7ERGjKUojIGxcUfccOVfKvJmquESTCjLOucK+ueC6
hmtiHZnBCm28rbyb5dTS9cmOrFBo3dX6iPOhxaqdYU53ZTvGS7Waf3H3cntOTaGm
5sYXCkyuhixW01HyYRc1p+gfS76DELuU+xtwsm09MyXbioVsz6/4ph4DRHq/b5Um
L1rQU9NqF0jxHh4xGr2lYwwKFLg4R8oRqEKLZ3ZG2OmJ/oWlHPPxao8w4Iy3POl4
M1V6uyJoGcxn/TOCzbsOSFJo2qDgBF0EMR2Ahvyb3xANJR9sVbX6QaAiIbm3H50R
Nu/xP1i3YlvAV0C7wi8TLvsQ1VtG7sjz+BugxGT6udZF093USTxMQOrvKbeRgO70
RvQgHsNFSzX1tuftU+TmAKkstcNZFjsrJm6CFcP4mSwezCxCSD8QQb+2Y+3IcjTG
h1AW8rJilmckZgyja714mrIrBgre+y9NEACvu2wKYtSWQlnfp0E5jVoedeiBXOmL
fhx69QzDh393z1hTjtkRUeo7P0tzi4cEXActMerT2pmH2OoUyoozsq16oUNQu8HR
YmPeE88nreLusmrhg1CqAFtrbL+Bdixyt6XRdGkJ+WyGeDAiMQZQDbS6A44pFpqv
UAO0kt3sM9Jj2BxWxM+o5gcNKFa1IdlkwLV1qGR1rxibWmUXcgl541/44rpiNZkb
cwk4eA4xS8lg0XRxDbmzYpVL6smmShkUbAR7uQGSS8nxAbED6wsdH5lw8Atr9JxT
diT6tCLnCn5zAgyNQWzJGcHLbnctyASONPJ7NURa2v/AChjJnTbVFyXw2pjbOuSG
xAbacUI5V48FPKc7JWYxFs/e+eXCe9+/0VN92TXt3McfUIYeBW32riymRk+kosmN
GcYL15ic3yBvQx52+2iyhXTMpw+aWUslL2vIddU2/N2k0iaOABYyvmc9OPQ2raRa
tClxXOcmUzyyC3Zt78YHwLW54hGszbgmt484eEy9WAZXhqNOFbH2RPJx/oDjpJZG
jResAKfBYEXv5aITUBDy6MjPm5Rj5q09eHdQRLp7q1mUlyZzk2ndtmasxlbdl0e3
oqRZ1ii+D5EADVBgddzTGX2p1t7NsoB/dsvxlAOOdWFGXPcofOchSQJ5mD/nVU70
4t+oSqO5c2AaMcE6J9zOPA4VlxAO8QQ87UUIfZsp75+VdYDTW1pCfmSFmfPrGmjo
h78Re3G0x0Cqvklj5fXx6dC5DCkk/7SuP5e4edb2IieOIaSq9Z0QOaT7lTZOZY8T
9id+TPgt/enBDTmYeBTU6A0YeRom8FSJq882C+UuuvSZDfm06MuSCnpJubDJdv1S
KyTwStxLiG4apY9xJS9dJt5bsuK3ucBTyOR5XRFOiDCgmGg0t9VHnnH6nYEt/6+A
///4VNIjK6fRbj9h/UsxzYe5ljiREotX54Iw6o7RsiBocKlabdHIaBiVTX0YLQDa
4fwViLw4XBPJcK13KWIwsXMRaMsD+YSujs5F6TpqnOmFRJPplld6V+UeNEyZAPPv
ywFGSWcPGqu/ay6Sy/HfKZui4WssnXuGlnL4EEpohFCtsJCTPyGfS4+7moEZrY+9
PElvVU0tCG1Ye6nEM0vg5DSQB7XFrV+sCJcGt3f5rw+HZD9VsRUvmL28Z/8w1wgF
i8qjEMVBceU8DN5LxHmvfTnq/G6u/dN3493mKgjC/GAyHRb2+UGk81+CTwXjhj50
WmeNeNHObuimQUiUlrm92e9Z3oFPGRF4cRfgopG60isCrV7Ctn5mA1Ugnfx6XKZi
54GWtc9EQyOc/ubVH615nXCRCyD7vOb4UC9Cu5VmFIlA5EGoLOhFrsFja1O2auX6
UaWyNX5qutHH8CI8T6ra3gIfufCAyVTH5qWjoZ02l6l4Hgi5G5Qm5zmoiAq7HeMW
g50Yc4bbolmaxW12IaIXZkjKLqw8FULiLvttS2mvemvyaOQ8WdNPKiEQnW0R2+Br
jgc5GCSQsFoVxE4hYZkmksUCWxCDDTshx3tnl11qzMickNN+qDFbirXmN4hhc2pY
X6V0w3kW3e/uo4ZJ9jdmdRtX6nTQoy7r2838DFfVYJeyOQIC5cPFzQVLx2eyYEMT
1iA2+sAFEuJnN1OoDCDXePwkx8yWw51S3x45YFrf97wWWyxHQRBSH3OQpvtAPK0k
L41kNOWX5pkddG+ulbOejIiS71DyyR8QPhVE7FPK0UgHR4WNmy2QK6zUu3YAutQo
G2eahUogKhNzxBTLTbPYu/iEW76b+qfnE0QIjfsiuTDJnD/+oOsrYqjv0bgq6rwo
uR/DtDPnVI5Yxc4xhwF4Oo48HCcC6mT4GzBnD0La7QGqiaq5WmHc0Ehz0ED1jVa+
MhUKEDrkE+K3RCy6FP5VkJZP6aSKUHcwhMqSPvpJ82m5Ekt4qrVcaxdDIfAqC9hl
sP4MM3FUael7Io5Ofd9OlednCq0IN7PY91G+Nf11cGcm9W+Dau3dByX+cncaGwEx
l/xysoEnpzmxIKjkcwIMHrJW6rMUK7bGZE80a2NU/Cqo/o5h2nYEOtvQZvYxT7+l
3ETZoE9WTqX8DQNMkDWyHLIE8c5fo62azu42F4mf61smg4rNj+3efN5FwcfKxJMn
HmzChuPkzAoNJsB/8Fc/RW/LyPh/WVmpt9dU7HJe4HfUi/ynvcELAchy1YbVP1/d
TsITKHAxU3ptxGEssxq+U0Mk4HUSWKGkAFGLirQkUjVPLTCEczqR4yXpWSuzrA0p
eoW3rQPv5KG6Gdh9lz3TcPWyRfNY3Kw3kpTtrxtk1ToOEes+kntZbbrmFiTYRz3L
laAJpY5LhRbVw3cV7b1GBOAWkk1ajP8U7oNhq8JgqrXy9dIZ/ruS9m+8Qt9IFE0I
QS7KBBrkQ3jZI/fg/c+XL0IwF+3EfClmDHwJSJ+etQhvRdNmcrcZbwu8U45jmDzt
GQd//BjfWR7Y9XxtpOAge3EJ/fqv0h+Uv6BKJQM4/77uTTVE3Q9lsJ2LUuRsZVtF
14QG54Rc2/3U11uKNV9bkaMVewngO5ScABGBh0ynGBVZXAGs8WCZczhCYTl0vjrc
qGOzfwfIvmmpBEflbsOtQ72qHQyIOY+uZDvz6tm/CpYMaLBFhoMf1rHHmD+YOFYr
AlviR8bzjVHpRWi+BpEg9ErD4RDbnWxMEMKNKVxW5RQIlbKSFKE5b+fND/sevVAT
ULVBb3e3MJQKRJ0T59rULjeCl2g5ddAyjPLmLdQQxcA9j7aNOzmcgTslypSki6C6
OraJGUlrGkMeZc5meJmhjrYADMwSvsdlTpcqvB66EdnwFkXM1fMGsQxuCM6V7GS7
Gjzi5P2cnAV1W4Py+/wyUU1AFj2hUqZQFsq7u4NucU0PWMOP1Zl7jsGLwXSLpqOg
vq2zZe9ULBUFbNpC8Vd8bP1wf0OF3SR+C/6BXr41J8XRYEX7oXXFk8EOLmRsWI1v
QPKhOwSrmszep1bfl4x0GocMCoPe50m5qoIcsKUj/vL3h8AiO/rHXOZBseoLCkNt
cWMsGvSBq7Y7pilQ/9ZXzjxmzfUudMOsODpqlUCE33v9aeuSWFPU79H4c6/22itL
Hs7EBk927rcBW0ij4fmJEbjqa5jepSdRC9QNWGnotojiX2kmFnReZrqJtgCWBh1A
tFcJK+pTONeYVqsFXXAMezcXbVvSpLy1e6ptjK3SkpBsr/Xfc1afPwNhxo0VFhN2
W2Ces9G9sE5zairiy0iBOfTL0ohoizorq01leiqlAcMAD+1Q0CThSC7s/V0FqOyY
QXs01T+N6kg7s+JhqUqjnohx1Ah3Ice+BjVLh1ZokJHwtRg84fm0EqXlfMo1mJvW
JwTFiZ0BPGa93knKU2r2HHK3sHm0le34WCDa7fUbRJ+2FMBKjZe/OqukQWnkUnyg
iJM1dlt1N5HKJWRpkAt9cWOTzUMk733OELM6Z7RxveJtTO9Xblu5icQlEzAmbQoq
uFQ9K0bDQ15+Ozm1BFdfAi0H1QhGgMhgNibjFsXaoAH8eZyOw4YDvUT1/ZF/Wofp
BvP29runnp/r9+IV7u7dExfzK69UkonjUt0jTCwmuxp50TsAIHVEscIIs6F2S6AO
7SzDq+FsNFmO4qf//vcHBGVu7CmieeETa0mekAsdgHl20+Sd+tgHyR/cRKOvSGb6
X793i6CUzGrFS3/afkbFbQ5Lq1L7Ul8tqmX45PzbJYsgcMNVxSK7SP3yJ+Oxa/NE
RfRmRK7k3dZn/lRfFXYf4JWzCozmlu5y3MwU2dyJh+tYavCoD1vBCyyt8EgmPNdX
wK++BAhn+t8Bc8McXAinqguPeN2STSkIZE1jWy5VdUgMcr266xmelg0YtoQtAfDx
lktfHlhRSS3knA3NkI17HJOVK6ozOaW9EH0226cCMbVgDuaHCYzRPD3KmZaH07oz
TQZdVpWCknGn60E+MVotq6rG6JSPDQ173yJOgfnyZe7fVgpJPp8Hwa7muW5oicAV
jAR6zUsYjNJSPMIFHDt+x8yoy4OTVETSWRkfzS945WgaKyHpHYL74ACb9t1aUsl9
rysFW7FQJHkhthv1UakX79v0n30qwxhKLCRV0+3xMX8FalV6xYGsg8ut4jtzqyJo
a5m5gqU3hyKzKOdyZWmxmeesy4wlJLVYK92s+lbepdvFb/mcqWjFCvIj7z4waTzo
wloK07Nf4foEE060mcmpFOT5QD+9R2judtqGG27sbn/cHZZX5j18Zs6wNJsg/w11
3LFv7tZe7Uov9sAGm5WWG/31O/6DdjIifVTkArxv9OqclmTSu0cFHYrFGWKdOfxJ
ks51UZV8QUdFD2zOfquoC0FXBA9CwFBsVnL+YQ+5itR38BgvxVEn+auMcaoEv8Pb
r6E7dcnPAd7+vpV3RTBW6/OvOb1NJk0L6dAc2FX34YRB+61nwkIdYNWoOjMlWRMe
zUXrZYH5McA0PnU6nUoGmviDqJXC3+7FySIwhuoCJX4WxjAcg7AYZJFbAICiiawQ
XzJUUn/7DZSBbgfP6dma8ptoLVTQ9+oZ9qWurA1gOlI6nNIqIn82EMQWpQOJA4ED
XqB+ddIpyzqtkFb7DW6XkQ5dm3K70kDPX13aA1NGTXwjcveFCweDVkrgdWst2s/N
3rX+ecZ3Sk1aPzNtB7TeifOS7q82J5IjtwbEbBaMrYyAxOEfDSbYLFWEKhi3amDk
WoseUNWwbFVBxTozSzJXeStkiUsgywWALNcLY/wUBY5HcgA1jwuC/sIqSAXCqP8/
hqbeqXoZfT5Ty9HYyJd5nDyaygOq6Yyhyixe9G1h0hZdAZwzeqrvfWWCw7P2ERLU
+7E72v0wJqi+ISXiZPQGL28IiM7D+Xd0Is2s1so2PzwgPpY+/07UX5xWH6Xm6Vve
X0Bnptz36+anSDz/M/4ce8DLhQbH5TqYKY7r6cMB6NcX/rPewzSQjUjZEz1dHhgJ
SXoJox2Spcn4r2scu+Plw1M2SX4Buc1r/8ZKu1us+kp2RNu/sS//bwFf+Yx37VIm
GU0wd+oC4qsVXZm9m5pb6PGww8DoySZEvgqnp8Uge789MY9fr8E/gZxKZlJc2Iff
gXjM2drr/nEHXoOwf8K+902NUYucQblBUOnXe9UD1F1w1qwmd7OtuqJBKN6bGEt4
cHLY/uDphFxUOWISu8QG10Yg4b7RguGMHMXTmXLE4ChyxmY3yPlTHoyRDv1PH3yx
i84r5MNf1WAaenunOOGczUa0I1lab9Yczi/D+VajgvLIQgdA4EDZIiZFc4vrb9SA
MvZxyfkZ0zntzv5r69KJmcDnaPb7sZHuO87enVIhMnozy4cJDBWXcVvGcJZ2i5PH
BdNIarAJmWR02QSBtcbjsN21CZN9Uw85apMaj41gG5ztUv0nOePG31cadqV2GsKC
2Y3o7pnqDRxdFcnW0waUakp9lGW0rV/SPFAkijfG5xf5Ot0vf9Yl9RlcKQG7a25R
qcBiTtCb8UHHYF4u+3DqnYpWjDT0/IK68U90rUj8bd3uTUMlLZPjbEZozk1trZbj
9cqhtg4a6h4TPCUksAmcFyDH72TW4/2xbEWvRzfvUJ8eHpbwejkVt3jrtUZ3BWI3
XmqTbHBafLP0+kEWYiE9EGE07fEG4f4ZA6xqNsYpK3qdkRS913yms6JG46EPQzfg
jaIIy7fq6oCPVjrPft76za/MbWEaFn2i3hk4uce1aJLe8V6Ul8KjsfUhFkzLNNNj
lebA6x8ckJjWKVCH/Y/q9e0C8gDhl/a8dNcdEEZoIOr9U15g5rKSPXFxxBprebN8
YgPA2tmq/fqgdHGNb5ozzfFBr9C9MkbGBT+YSNT/2AOwAEJ+uEwEMjqcBajDQZso
X6ZO61AsIWRiWY2XK7yhieT2C+o71qtH92mUpU2PzR5YUwmizWNfNLCK+utE6q2F
yRDQIjY2WJz902cXahoYeokF9rXE3JbNZdewJ/P4MVgqWfw3yj++p20IU+f3O5C0
/tH9iL1LYaSqYNcSVE1CcnS9FjZhi8Ur0Q+6IMSRlRBKOdhd0SKQ421RvezbXaUw
wQV9Z1apcJmeXFxi0Wrg29WVzpJcfTRAUkXsDoASEJ4EA2hKN+0kIFMq1bbjrVUi
nK+F5yjekOiHv15tmwhzgTAt3eO+UsKRPsUd/gYaNnQ1+oGvnTsBNZJI/aqVKiEU
1oSG7W6cKfhQezUdWzIWNUceWYLSZgtc6oe+2T7LqSN/aRLI2/DfOTkDIAtpwiNH
4U6fbt5Ol/9w2J8fyame/AjnLB3qCnPhCGP88YCRKOajq/OnEo9RA7BdjVeoViQm
uHf6Jk0dPUSYMh8PrlVBP2zHNMwvFbs02y6jCwyaKR9bR3S8DCVFEn2MBeKAVYGG
TKid0+EF7l2XPau+Y4McoupFwAdcbw1yQKtHqHb8eODjjDxn0ghlP5w/rw3d7qiq
6W/UCS1UfO/p75e2yukHzagIQQfrj3yDlS6pOL3eW3XjWc7HL9deZN+m8Flxaw0R
2YUO6CSxp3oIm/T4PtCx9RL+6Dy71JmmDp8NaNKC6NsX2oEdNGsGUL1hN+D0ceCe
FmTb7lTRq6utJNVlNWN7oMkLbAbMu9hoFQvDey+IyMdfZ4Zyk+tb9jVfRU1loKmq
szykSC7Vohnlf+EIemFropA6EyjOVkF7YOMHSb2IIbresIt2ExqquuiXxC9umfy2
VPHlOaYkcecjhtBKjmwYs75xtUwH0lyOtdzX+DHbvWs01SA50b/Cx3AKSXzkXQZa
vcjyVwpvEQyLQPaghCVioaqDZmrGQloZe2JXp31Ek0e60eE8ktPUiZPrucuxRUQl
wCUoVzR76uyE31YjrV2/Ry3JBO07Agx8S5dew6oFMhWp6TAnyaxqydTy6NVR07Pb
iwKmZBDuq23Tup/z+DmRInObLNThRhAPUFzwhk4B27dIFE10wVL+3KsjfuEMkC3G
kOs3TLe8YyQj28wBcxRdP5fsLLwPaaJ4/9fmB3COfERaemOv8GylvQURmI36t/zf
tOA+YoKxv2hTpo5sEV6Cys5S6qAPSnemAY+y1wPr0pVIOpYI1XiNaFpisNwM/ege
lrzmrnACWRFGpnxvOOPMUGedQ4J3TrTLpzJKtRKBNeXwmqD0wGTELao2oz9Elid/
AAyFN/GFVRFiVer/1tJlg3DhSfI4PSe3aebMMqlbLoX0uHXYcj9MymOTrqf326Mf
JBIfC7cugHYNaC22hVx/PIjnCKT7kN65+LGwZHJ0P8A0gJGuj3f8Slhs2LQQ17A0
xEWvGUxphEDIk/UIY4IMuRIZ9/FP+rrnrlvQkW4M2NyiJa9XogKZDNlr19gCqC7k
TdN+wGyPyH5gecl9bigb9LOLvFVsyMnwojluMY0XE7amgh6qk2Wp51LDgMnfF2TA
+/XbGVv4oCNvElTuAtZeTUFB7lHpsaNoWg0dEugDlyuHVjdSwvP7jM0DOM4o2xIf
jqwmMo7Cqd8RUhonaHghacjX6w0YOSldLSNAPls3WFgKl26XAN+U1z1GUdNkvSJK
JeNiYAFXdHFxx9gwg+VSv8rA+/402BrOoZH8BCvWlmXzlAONQTDdh0wTiT4VKcSF
R8J1zee31pLaYfuuThzUjQBceIgIjg7q9iODddZe5pwK8VvotJtmOzdB7HCrIFsJ
2p+azTid+3MM4HzPjWx8V+cIUOzKNJ+FAVAoYO1RZ22IZMxfrP6BQEgZhQgi2v1s
z3wv2bkS066SBAFdAqoN7uSQdZVF2Rx2qFQvD2J7Gf2C6L+YTZ5J7Fe+1ZFuY8aE
smg+rLFUOzM3jIM1oxtlZkK1E1Y7mn+sfPyKaN6hWI9YtCRYWacRFOLLUplh9L4s
9gGug+8ZDTVM/ngFLDdbt5LOHy7xeVdWfCa5FFFuYVB9hEQG6zwkh7RdB0VtCBVO
OBOinVKIXVUchOq5U04JKhVYvVtySiU4XfcYgE2x9ei903x8yBhpdQ2Z7W+GvLJ9
q8IDBP92c0W3cDyiC4VF2Notbe5gwYE5PNEeAxzd8yTfrwDZOk+2WRsBkhjso+wD
8U4WKZBvzSMxWOPgW+8M03Xj5ApSDnaC9I2cYrlqYrGGkSPAQjOZtoXgwYl/rn0G
t9B3I8COTZmJbABD9arxPdxVtq0WU8ZY9E7EpCYpIvg2kxbyQCokV1vYhgSIHhYA
ZkQp1PKS+RRuqf8oBQPeHc3mE3AwD83aW8bfutmYhYxVHsxjNzr36EmQsjix9IMp
kJNVDzKpwjwbWHC0zeXFjoU79ea6AX8wcr+WBopajieKXTcb4IXJhIPNaZtf3Zu5
tYEvj31QuIkFtAYyxldjhvPcN7hvCdJezA8IL3BI1+RbPp+T9tE9iOXVF1rJdtyi
21kBd9G9opJwQ7O/TIHZsaHTVkrZ7/39kQw0BmUGZbFmEQNbX6ekUjkbNM4w0ENk
GoObTjCHmKlD2PM0jkivXj2geNohLXc0J5u3WFiS8VkZM4mbC58fF36AhA9rOcPP
WV7m5+r9g9VKloSzdFJ3oHyvWyMMOwzU9iTPXaosuehRsbWsbeuJEJvLVBTzrb4O
y/jU0od4c4TNcuGv8sq1JPjBBEybgH2k+mWnFdshBwKxS2sWxzPHlNdpGRWhwWhG
GEdhVmmD+JCpGiv42Nruc2Q1Z8883edKvb3kS4gxcO8Gqyj1f4eslmVC0EIrKbdo
6uMH8foZFSH6DEYUfFlYMr58c6xASqLm3r/GkA+mwtqqNxjTOLMD41vLzyEnF8X0
MGeuXASPTYtV9caZVPeCincFqlP+35XkOqxaSNk5MOQ6P1Jce5se1UTMAxlZmcrS
AMHwGBGY09I3phKFFvPZXnxeSqyRMIwMz1KGHxDPAzFUTp9ufXq7iJKfZRxa+cDz
1b5xcz2ovo8MJQC6fpByE/ps1u7Y0nd5uT9Yo3UiQpR1XuvybpgBOdV4acpXoKHN
DFyNkPh3KS2wfynCZAQzf8KshGFieyAwHprY4IijJAEncNPQVI1mhPH+LpLZtTok
CCz6nfgnTZjoLjJXFrdwYJ+udz3q657hixJ2UTCxU2lDFkB/O51hyaQdg5TYc7Fm
Vzn7k3o7dZowhoj5Fx8+LmectEzgS2ktDLKso8P/1h8e6F+4wSVCDa5l4mxAQXN3
5q9xma3qTMfWGIIwSQwsRMX1WVoQ+WcprLg/3M2efmDRXE/+5HevSsFCwfgaxfCq
N+HdvYHPnOq7kXe8MVxcvjF2o1Y6I4zvSHzJvTZ0G7UFCCxGsKkYing1QT71LeTw
jzf6Eg1VpIpxANbm07MlSiyxKBf9fs4b/oajK5xo4avadv/o3djyRFd+j5Ian1+f
qlogcpLbhf0lIWTWRt9WldJOPKi3PRyGIehpiI59LUmnBODiVwee4BqFDL2QxN4i
G6MKFp9qvgZQm60Xi9cYtJkX3MD5GGZjvU/6tLk34LXnrtql/5L8Zf3a3KUfKN9U
rPAdnozo19pjGv+ZiSnWPKp+kJhcC9VvelamBB/fHHoc8F5JPR3ZqV/BRG+L/VSO
wVBQkRagLPq3PzAhVXNTADNHOFu5LNEIRNNFG8UMJnEHQ9f32sUkfuRKIlNYBlVQ
Ak/nfpd5GWmoYFtP6+xlJffzEeT2JttqwHIpAqXefcmyHXFT6jtBpiLbAW5tWwBM
vKd1ulEj7z3T272kjsrN2fCUCiKHffInY6SyxVEpqKmSkX1/8Sj+NkSg38slzxcA
N9DoNmiqLx0eLgf3qiOs6y4W4izEmz5b/a1Xz/ycaW/5vnwikhUWX0N23FBHfgNb
WWlLVuE4z+Dl98HGgk57Goji+5GF6ZPbsAwg9pv1/2fTZh39pDeSrJNTt7Zi1LXY
wyv6LX4aa3soLd3uC+kr6utV5SNHZddYXnr4hk/wOyiO+QtZm0Q47V85BVVz8Hw1
z2gLZcjRuoXzlGJOokG7JJvpCnhnMvia/i5IMEHMVDhwXlK/qP8hO82zdP1xywDv
rAharkErOWofYiT27E+Cn7kiu9+VnsR+on6Os7IP+vvS1ybgvjNUYLK5JO9fdXLs
H2y5wGfxAStnwgwOFrmXJM9xIrDEJgdLsmAckpJKBmsqeAagcFmcjbookL29oXQ1
TA/mc1dX70IxvDSggJA32a3XwctEFkV31xlFm+SANYQsMLaHHKeGet1scw7X6iU0
2N6kM+YC9k3KtZF6XqjkFWNflZ0jwzb8WMLKvQPP8Ff5krCgWmszEPab8Si3+Y7D
YwZq3QmndppE0eIPB021PwmX6AoCiMhp4yEPk+/ylw5GG3B5ckDnW6J4gyAArZAx
44fm4ddjvD4d73yDDZe2F0TpgQS+NTSRECP4PqWy18r+vanb2WJhAh4IXwZp5qqx
UOVYg/XRGmNmmq6fSRQsgTEOJR12/nbj7w9Eyuj/pPJql+Kvm125aJeGGU4/If6A
6c1IxItPNtfJNg3BSkrtZ9FfXRK/UOp4PUlw3GXxqJnK3PV2GQWpeqKXyQcrAoIZ
okNOD3UcCK1yWCku1XWKq5M0xBvcfSRwuPuUWu0fqHayyxbxvd51K5W7GLTJStNZ
WJlCYyyRZRvAd7sNigZb4HHQgAMO+HhQkgly4EWnNAeZY7tVPxgPhH2PGZue2xUk
Ji69tPIr+TCQMu3ERhJBPvnOygLfimOwxHvZkw77jQh9SFVQ0pUbSmgjiixKVBy+
bjEj7MYKfKaV9R6GHbRG5vIGeIvs67nh9YMqUgnyCwgRhzANzN1RkwoHaRgwUUaw
ZF5eGcHLMv30GTRK9EkHCsRBbJq9dg5PFLoA/rjRDXKbrehobTDvqp2mbfbcYcDm
4dRYM7Grp7mvgeESbHza9/0/a4twMvMKz0BJ42sPEq8hfc3kAdqMQHQbDj4Gobh3
L1kHrL1m5FA12gZcNnT0Md0P3vO34bLz5kp+HWQk9TEOD1bYhIfz82cQDSLBoufv
+38jpYWNgB8fCo5XTmErgiM9MW7+ziKTHXvJKEuB/b70Z75WP99G7I8RqnMZx5nM
9J+vujrzD+suwssQDuesEngSHAP9Hm45kqZ/i+U5OVJEu9/VreG25s/+1boES6JB
vdjWBVjO2qTyfisjCqcYu+e9cTcOlkb9ImMNJv/9sW20PRPCi3fi2aeZBtwisvUR
1i8Tg9chu4YywXAa45jIi88iK91v1RcmhHmpxtRfU/0Va5YNcfyHiOhjvN+tzPT8
KFmFo7KMR30/36N7+dPOuAXLVEs17wJA0XQc+zb+B3Vd2eydRv7OugTy2VQGglhF
fnZpL32Xrw3iOU2L5l2aFAGGYKZvLdtxb/tLXOmtSLMR5ks1cDz2Vgp4n8JVLEth
oxClE1VpUHjZjvia/w8ZYZg5XhwdJfrk2G4vvEavV5Ts1h4vFfxgRO2wvGBB+yUS
wrcGv4qfqgiE+JsHKefHOiPrAGhbcM6mn+BOQs3ql+fLmU0L4XNpRFFQFIeRTrQF
HOPTFT5ABL+wCIQ+2cDnubmbch5o6896EaWksqoAyPRHg8KbDwmf0L8PXPqNHEbx
xCz7/wZuYf+Bp439V/2vrYOM8iVXDKdSV/3PCpa8ld6nw58gVQqqI9pbK7h2VwVn
pPkufFN6hskwYQMIZoz2yKYwKbpDhYrJ02HKGMfCQ7LddnYVGjvPHt+X8MMUCtgL
Q0EaXErOAFhl5ExRW2VBFl473bsWM2l43Y9cA7UFOpewTX4/Tv3Q7xBdCdFz5MBl
SRoYg6xQ2d5op2GgrjSXJh5eP9kASp7z5pAeHG3IdtIZ/MF9w1cHnXXoJjqYm1YK
G+ylxbmyg/aG5EzqjqUgT5DnQMkxdtXB2l1SDCKqOFfjxp2kvQSud0midw4kFfOd
gGsFz87t3zp+/y9kSeNOwXfwbTFpXEM5+Skz2i8yhOR7bZHn8XiliUwGQZRXuzad
tWY9BU9NrCaR4ADbW5R7Vp5IKgUZ34JsbHK9CVoLfYGXUFk3lr6nHuqXCssmxq6H
o9cNQk1pmVC9H9alZ9fP+IxlGrfou/wad8DhfMVArkOJMtLmYyb1c4q5WtoSk5iA
ldpmOF3CS9TMvs7p0QbaXX7lLWg2v8FbeC0DdQVEsogLdyFYRSZkw0PfGs5l2A2C
QXviy3Y0iDu39eDAgBc+TxaDdK+R2xw/lyMsBfEqdLPK4I31pN0LuMKEASPRs/aU
GyRd0WrmHtV3RZxqsRW0eMuNDW8IApd8JrRzaPmR7lgkF7+9jAecFL0zmSh3V2jd
V60h2jW+kPNS28yifhJYrsM7eMBev63ssDG443XNlGBsh9AAO/IPPRELkvRvxK5G
79ng6/4p6ulgWiaMI9e/MimTEZLv3F2+ySvhie+qVGgA627xpptfOTthHqxgEkY/
R556L9rJ93ZYdCvIxzwJejXozR4UgNiqJP88FqgqnO+j3u1x5MMRi2cf9FeJXRIq
9aUzgkKYV9JCCIbg9+4srp7WB8DNCvZX5C0A2b8kakVL2oaO8bXJNurzm73Ha0Ot
vs5rroZzeDhxOX8sM6CS2L9khQSwPGQILnKPumlJHBfoSP/er8MIIgpFKFbnSq08
nT7yKWbY7plGROqcJQSvkGPexovWsaxINgrJLGE1XvnNiep5XEnCZR14M8Qq5vv0
uvuoHuzGiHggQGpJAcvLAvYbnlpEF+9QXqH90SKAizy63Lmdk4KNZ4DDcvOdRB6/
UnwGu53Q15S9ZdD6IldJsxW5a1iklXu0fqUnhL/ygjPqQBgwJtlqT0B3xOHCpoZ6
Eksfba17KK1mz2qze4iaVvb0RfElyogmnbZ6cylEMZHF1YiSWX6fyuBxmv88KTJ8
Amt10/fp0IqpRy9CXILyAPnOqeGAbyVEy5eFAxKCP0CW29W0ZmZrFnAdKECWHrqd
uyWr+9Dgck6kQykdzHKNiT9Rp/8TPVm/99jDxnLlfedGJmhWXR8fkuFoDllEavOf
VuovzqR8Wmi34pGo0LcMLWzMqmMAxeq1IE0btmIfMIaw3UCyZj0S43l1yc13s91J
tuxYj2eORdVpen2mioXLGVCUKDBnyljmNrksHvqyVy5T1CD/4kKIJkP4t1Q4fv4g
weSx+NJFB20q7HIZpm6kpGO1IkN5DUGE80hjmcj2xhNrRt5zjlKKVOsBFjtEbeiZ
LQETZoZJ8DYQYx/LPeBf3QJUR9QjB9shB8BYupHL9GApf6dFJZ/FJt2Qa8sHKVSl
ocPs/0TEQFhHEIhw6YfFPnznX2yVAuDxRbXP/FzbQhc7g1Qjys/K2CixjUx+5xmQ
h0gON8yY/0sbvnAMgqKznCCP1cJQnyQk8PdxykBmINMpJRaRQmZnxnkf3YyP4FO9
Cpl8Sh6JqFDAQbGyNgRm8U9rnrwuZocnZ/v/GXO3yDIb8ajSoktTJLKq99fwFWSX
v1r3u86VNjbzDosnLXQrds87FnvTYa0KKz71U/gsuk/zpja/2GBHGm4AMmMFWMNg
g9czjxUpTbfV/tVk0Y404gdz9X1ziSWBAJQ8A4G9oAN+3ZRB3tGdugm/0mrizNXf
WDqlvBQtljdP3+0+DH6o4uoJWsO9ClZItNrAf7+uY707YSz6bIZT2tzFpKYHj6Kd
bFt4D7EiuJl+ROo0q89k+nKQPo6DOa9hT/4kjJbl9CcxwJaHq1nr9rUjQQbaHXqS
ZQfLHNFF4O3pO3e5hwXdv/A5TqUqm8U77T2lWeFWKvI1zsIRvGOKZk/disn40yah
SH5UtQRLcd3AiowhfJMjQMm1CLC1zywWXYs+HML/Hd5XRHczUPKtepbPK4ryqlbg
9TygQ5Z2mKEnHeBsykRRKpqpB05IZptpcPw1tc6jH2gvmNKm2rOcXuBWhiemXLYV
eFvrMxaypSqgDIV4ygzfk09HIS+AwmaZtz73SXcq6kGEWlrJx3CFVfjRuywmEGZs
cDoIc6a1XGWki4yC/P0EyScVOFckRTNxk1lrNwaJaUwiJYcR2fnE1P5oOJkvep+e
h/ZOD1l2ZfmdV+t7X4xNJA9FDoolfTZyWOBn14xIje41iYDkwDc4ZkCFrcHVjWZ6
2Ll1vTHrcuG2/3oxAqk0QOCOtj9SBUPRB+95+Z4gwiuZW1eOi0IP7jiXjIdEV5kW
sgxt0S09zMOEz6NyCs6sKGdFb6yehNsbZqIoh/KPKUUDOVzCHqe5x5Q+ox2kpKgQ
TIJdkA24ll/O+GIhkTEcMHhzlvOABre3wThke1vp7x4KP3kv24oBMl4zQ+kli23K
cMFgpcXf1FCDQd+UajJzlDYgTPLZJQ3WhBfzZVy73FfATOk2b5sBahpddZftcWCN
ojhnQXodNVC+0R2oljYE1rRhhEWDOHavpSEE1+8icGF3kxqTzJc1zsR0L9Oc5DBX
xy8q3cix5WKxpAv4cquet4TzghQiRqKL6Nfj+nusoPbCqpkja0omCLIelVxXUVGi
Hp089jgGI+yUAHR1j0RzKbCV52DHApA/cTEAzrp9zVv3WanJxaKXVvoHMAWTIZ/7
DG4kgg6yj3Ul5tXzVBwIKZF1eG8cCfBmeECXbytB45lj+brmZirdih8g6fEZ8OIp
+nzAIOpGvoCBYwj5J4QITF+iKIFvqtGvRcL5A/tE+BsgePweGCvUcc8XziSLoJHr
r6aaFHWumRRFS9XMAqgWmQp0xblGWGn7CUH+f6610Vb6rOtw0FBi1+2nQov5Tgef
u8odh72wK9TmNBIOMgfKPq3iDsRzbd9XF0z6pETQoR37knPz0SuVEWsMMpGIFGnK
oh1tOH+g4+g/6r3oYemN/GbHGuoE1uO2ivUCmUopiKoCrtq6Cq7VCr44+2DrrKwt
nG+3Brr/7ADLPN+0UiWzcQVq8BoyIamEPQk7wQ9nWK0bs8nuzr9Z1ZYjoxo4XNnP
SG2ZPkIBE3LLdKVZN7XUv9TzB62PutSP/hcuGpLA/j3ENPDRMicrUwAlzIbpzjhW
25qM1arKUtlH+Mxd8pHIsPoaQIZdSqTGrDqD2DtzJUqfNBlt7oTL/XOw6NtcIAxV
fviuBd7ID7GdUEKqZM3bUMyv02GmET/4pi67eAhoEEQmV3PMEYJoFkjInNHYwLd6
OLVtmcAiK2/R7rlJ8BiOgzRInx09tvjm5uxFxFJUjULHaLz+FTaqXbrtsd9mO90B
3/ANp6Nj6u6+Dyl2J2DrdBll4pJKS2sgKpfI2WODao5mF9YLpeeA2qd3V1L81/G9
+mLQZHDK6uDi7nd5sSx09MyXnUoZQzgu2OIQayMzc+htOTTz6H367omm/O97zqD6
O5IQmVwMxbVZO8Hr9edqXscxbbkj+YfwwTWIQ9tVsXuQKFw3tIKoUar6JTC+9Lmt
Yxa7c7JYvK6ejIAJE7mGLLUHAJEanuH+drS47QJS0UJpANCpA/4lmZlfn+T3lDYj
98pK+o20a0UBea6Ck8h7f2efYpIklfycIVnR9CENEtHgoo/3bXH8m8skjFDNM6c+
sI3nQSnkc2UXqucMh/Fm5LLKSzy9Nx+g1VuowEnGP9Zoe8D9RPUJOAgQ3ZbisQiU
D49ixHzScD56iW2XkRTXwrOCaXNgAC6wB2PPoFYjHYTXfYFm1e7q9fYKh3+Bh6rc
b2U4A8ru9FndsxU3jkMBwYsy6r9VWcPmflxPkj+WLfz5hl9qOlYCH3K+zgVT8RmT
fe1HOjZfMQxbD4mVCv65cA6aWL/9hFwdVBQudhiHCUD1cfl+/xpjCjvHt2XLPNoE
h4Lm6XtWUiOgo81yNYKFG8w9mYZR0fv0Q26uCgUUybOEjlTQQOQdroZPm9AHAabP
QzDGIUJPmVv3p3H3q1u0ARiH2ZT8y3yteuhhe+vEnu0OlTGN1L9mlXZuIkteWNTA
P1td9LYWRkdUyMPFLBhdFdJWGdjKCrZ19cGUYQFQFrc1ZHl6+DLGUd5kP75mZAZS
RlHAjIQXJ2uu/F6UcJ8LtXCJFGCpBo+PxKt99MR2NGaxgjQvIQ0FX6Q6qcJyq8eZ
pJ4FffkgC6tFtQ8b9COQW3M1cbtZM8pD/0tNGwu5vzy9GN0dcF1nEiAW115yU9Ob
cSDSPZuYrOe5Z3D8Tn3hfkOKt2w3Pr0EctHGjw3nyuT1hhT0o7xGOkWh5A38AWOk
70y1qibsaW2BRAj3WJENwF862PJCqr6Z+rTnytxGMCuJURKj+5Szqp2VJ/051GfF
rx9yFPTpeW5OEhaEMCRsh0jIZ3LCGGJ0IIZBL0DxmUPe5+Efcx8d3kkEBzqav2wm
MSL8EisiFCZ7cXThfCPVAJyu/Rn5/duhjgDQd1jcyd5078NreQVbFQS4G1r/W9ys
7Snkvz68chHJ3B+/fq5MbEeQj9skGMVhidWlztamPI4CuAkGRuFK0oHUMlRB+GaE
NkfJzW0LLZN+51WCS7294lf08K0Dx3ExEYazFJJKNyte83KVNCe2raRKpCQhQ2Uw
xNy7THXCPrWk4I4hEwwGra+HY6hH0YmN6YCS36JtXkB6Fy4GdJrBv/J8qCf6q9fH
FdX28vXSF5cq1AF9vmGk1XthblaJ3ePcYrFA6U5fQ1plr0FKYXDLHxhwLf8Ghxar
VAOtdkHhO5mEuFW4d0+qgRPX8bampYQYUm6TgUWUailV1YmzUPnyR8TfM/l0nMVf
5POUPiMXOtXPrJ30BZrThVcaua5ve0qI+9KzMYNlQEkFCQ8Z+USPn9EQGHx1+Ne2
6s8KHfgvvLHbBhyqCvhHM9Y2g37q0pEk+5QGc3XNC3nJxGjpecDlNozzq2KQm6zu
HF4dcA4IiRlksyibeLzY2E85zQCnNBI38Hm4SeJfTJGCMKm5rO2tt2nfBlVbCZKP
wEmBnOCi0cuAQoxv0wSuchZxEM6aw8yHrlxVNXBzjeH9kPEMbdmVR+XxGYJ6snLj
B3eXcZhxqRcqUJicQRjxIVbBgwLLt+VXOSy3LsiXyur5km3UKbQPr0H0j65ZPkCl
95pQ5Ro3r05KwqfJ4DISV8zcMcyx0WTlypeItq7o7zOfFWqSC1S9pbRr9bPN6kh7
5eXFoiJul05a70gN4RN0jGKMqpO2QaAqGQL2KybYXgcUj0EOWhNp5/5pyQfsv1xR
hSh/dk68PxLrFX6h/upki9VLLzdH0QqYbUa5QRsaCiXNsVSYidKHkgvIb5hpa2c7
EkTLmuh5K9Nt64v4KwuRrdjUCnr0oNPLXAQ4sEr3iEDrpKqL6QR3EEFXuJQe4noj
VuhNCgEZwp0bELaLtsfaLDdgQZ44nbdNfdiuCKKf/FUac8+fDtYwNPGN02z1Zvmq
W+Ygzlom3/JBpRJ+ieFLZePHrmDmNGU3FyuUpu/6FwcwE9A0rIXh/AC2U6GrDPfc
Cr8fgQHN8rkGEmxSaRsujdI+AMMZUGnFyZsJV87A0uezT9tgNrxTyjmQpAE2CUgL
Fx3VUWtv83makQcesNhuiM1B/8hN8msrA9LuszzR1OJ66vnXW88mYOEDUqU8goZC
Ket5jterCw8n3YqJFPDHx6f3yDgdCLAFxmYcz+Z/42T6fgpmwQbBv4K1RXKmgcPG
Hwm1Ru437jGUBnoFe8xn1QRs7iiw8L6onYwYFQVfOv5+0rlYtDMbUtvFRMpiuScI
avAmjTXCh0psAGpyGG35Udt37PVPlur3nxWrE6eQfLqBT1woypYEBXUIy1tDcct/
OgR86YIWUcXpTs7V7Nrros1d72RUfFSVVnVEtEoNF56kV3GohWv7ZLTobDZ70Zpa
Nqld8bV1z3YvAY5MzwCXUfwHIF0GCrgsL2I29zgnoDDlBJzbZ/x2eOodgPfQ0TEC
p8vmKBpcDtS3GT6STQpuTd2JD/ZGlpjbTUUk45CMGW2g82tSMPUyWaT5gIah6NSU
t05LAREcDQmBGX8my0IQY5A1ahO11aZjL8kNiKT7zXXDKlXlDdjbQ6y2H752bIxs
ET6M7Xkb0kQY0S2Y8OYn7nFiqlhgXp6LIbeLNad42nkyfnlozNKmVyt36tXwHnhN
6pM6rbrQG4+Ck4aK2Qj+5jQGiE+YyPiaNmQm1I+ksDBUOXY0Veq62FxyvpUMLV0R
L9K2KKSOvg8CRtFwhWmGh6V127/MaAfEKLCi5nrKpkHCzHUdYASVEyfED+STlE0r
iacdwzapskzgvy7EPdWBJypyOmXWNDLAoouv7MGh7EILMpwYgOo1m4D3nBwpwEyl
Nz4px/kOcbK1ExiWMUbWgVPIQALgzZ2YHMSgYoe/wJRkSYlCR7bDZl97gvQB/+X0
+MalwfFXVUCP8w/jRBLuH5vLPDWQw5VFlG3V83WsX4DszV7q8zAGKgBC7xdQTh2x
Po6FEI1bR966EIGESvG5RImnLL3LlK5gPWpM2R0H/6nmyQSc+Sy7Kn/WqEBHYtZ2
8UwawJp1T7pTUDXoqVyOtC0tJWb+W229KZRZr6+wCITJf5uJfcG826uCw6DVuOqF
9nFiF8gqoyKfIyBsIJNz7e+rUtNq9NYC2g3kQeWcnwP5+vuVWw0JrcMPDFK822W7
Kd4hL5xJpbqO+O6DjbKHVoFB6yCDuO8Wg64lDeCrNQrajDkQupYZyTfeedvoVPgh
UzSDF04TiPVZyKUPP/SBo6/SfZcTvvkXRHnhmH9z6vdtBM+ZSx4QZ1xP9aOfSAa0
9vwIXoe7gKWrZiKwOWJZQe+eB+PBPpJPly1ma0GX37HLIynpopayjqifQabApvAy
rvWWsBdUY8M/25lKahHaGA+gmGqZ8hC6trYpD1oIY8jf3Khry9BDGHXe4hKkzgcV
dvTACq7w+xP0tUmjqnE9xlfagyyQU84/x1W0VZ1f64gFjHk2uDpmzMZV3Ir7Kyxi
mpNXmQw77POdHfx8k2SA8WIzIExzVXRYxYi8WbIKXVjpfGDX0thP6V5RPFTvin5R
bUtAPGS5zkCs1fSN9ilSXuv+BZEgy/W/yEzVTZVYml4spbKvkCtTNeWsydIgkcJY
rT/blnIUblgPLY7i1XuMEcvIagDUuV8ArFDEpXLzsGNtPO2y2UFK2p7lqIn3ItsJ
CGrIWtuWpF2eWwB03bIe8XrLFTJkvbK5U0FtTuIWIid7RDtZwi7qSXMeH+QoFZ3Y
A034FN+0g9WFC4/LlnamNnqnP9DHc0EDX1gNAE/RYtGB4xmFx/YRbvr6rwBpFSJu
Clv6fneYY9pmVZnpzX9JDiwsT3XawDPch3P3NiNna30ih1hsFztM3CtX0s9ToKk7
GLVRxURh711p2yNYuXImrRQ9PDmFg65i8cg6tgsNxjWWzxNdwwMJAzNqmg608hYz
dlGbhLLZvmpRnOGoKK49jTegsjUBgW4bPWHieLZR3Lt6wogX3VvS8oa64Gt9n9nD
zySr34+itYmpaVBcEu0V0Z4ZlNTPXcbeGAr2+d5dDtPTdQGvt0mZibgIPf22G0Rg
UWa20HHx9Oji4aIF4UUVC2pjdDu4/etjkSAlY4qu/+4+t9b6va0ajLc15SVv53yM
4SnGDOh4V7uvc3p2T4HN0k3NAULqqqWUr+QctCV/heix78/PGI1yH3gKYMD+S1+x
xPA1dkdfO9gegiIqjB1H+ApOi/X5wqXddya/84bOsoXzJDU9rC3I7tWIwwtFmFun
kY7vD1IRYse0gIOuY0coSzWPIDP7dEYx+qCy+WV/eXIx2yF70FDbSR/Wf6utfspr
N3TeWW+Ww/g1mFzfz9+ywNp9J+eTsCY4A5ayEiZvrYozWml2O/0b5PlTHwrk/GeE
tMa3dv5f6pLUB7WfbuTaXyNecjz6QHaU9GUbPvMyGdoi/S1VNWYLlSWqOrc+SYGV
RIK3/h5C/wHlxfafxeFISmkx7RUKFQz+ERmDaTmSX0LHtU2RlSEjFdMSoi4QyoZ8
6i14QZvyylACE9O9jP2r4rrS6JZwiUebevfdr+yusIdz3AFeL3g2m1pPSpTH+TvT
Wclf4Bn1g/8IBUZGUnQyQhPNu+sMrqTbLayCM67QiiBGzqIua42+MA3P3EDcd83z
fMnfdCsJWs2LE02DHZIARWXR00xJ1qJolvHwCAkh0LwzMJna3y00Kqb7QFWqsqkF
1iY20euHaG9S3WNKvHBa4b1dpfMZsmuf1CI7Ez2nwz9t/EmVTYHkzRYI888al2hs
F3nCF5CtDkblm/PKdeorMMio/rBRIdW4DxkTWNzBfIP6a1aaMGfEGJnX/3hp5pjl
6T1O+A9yiIDWR0dHOQHnKMIn5h7oECeO/bP9UVH5LuEQD/qHVebFblFTZaSbSz7/
`protect END_PROTECTED
