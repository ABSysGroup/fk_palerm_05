`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WKa3M84BEZ/2QbfW9H4l52dFTM189Q3sYsPEE8wNwc9afYcuLSCeKN8fE6PIhF1B
i36n059IEU/tYqKFfPhBtBI/uHwcexq2VNXotKE1A/v3Xr3Pbzc5fgPj1qi9UsJS
3xi7kEouU0SGNOPwRTWTQntYPv7Nw5zbZ0PdzI6gafo/TwgWwOsZmqRpYpOjrfrk
KinUZnKe9HRvqKo2mZq8jKNFFSS3FB0mbMYegNlvfJEbHCptz5yKnhjEp6rrXeNI
zknRP5dkSpMaY4TGlI9lkhNAEmbzD5OYxj/bhfuLiLNLou4m0i91XVvTbV6UenDu
Salx8JuxIY6urq4NPPPj2ATojkUWCgtaIfdLZP7NBPXJt7O2SJ7Svr6LACGrUqWD
bh4xHAhwIoPwUBe0VhNkKNrwZ7KJF2JRdLAnm589U7OAUFm2Ui2bJVnQjadSZ5Z5
r37o8tYy3exAU1A9AFjqWkaP8B9o1DruFhJpqBMk4xNXPUIGyMfz7zO4dJTX9PmW
0QRrmcIQHS0wgKl4j0M846jLKT7vF1VlEE6X1lKePplHsBRraP2peKkRe2bz9+Q0
IbHllHFEtxRY8hnweGS/QA35mXUfhvOHeOWPxhKwt9geyX1DEREfENwAMV6+P6mk
rkRSXREdHLplJC5rkpdOgVMr8uTj2tDHLANJVY4Xr2GAju6IZBsR39Yv/flUVnkk
RLoLfS3vG+hn4CkCioZJ6xkYHh4AdFGfsaD654NEE+9uJil/wMsN6NFL74/Z+vRY
L6pk5Qm6JfGsdF55rOYjbxcPPKQ3sE7majhW862RS6dlzJxGtGDtL2+WbcsH82YG
MdcSm9l7CWL/2Tmg8Z/yIJ4PRi3cSu61cSETvBKdmcrKA6bOGMrtbQC7uIixB2gw
725fUOjQFMsSlv24YDYaRCXktMQagI1kPw2cEHdYnXhfNyyy7ecdJmPldMBtMJac
Y+ECaDiVfwPZGkOzNhPhuVIPc7mqCsFo/c4ceUPtg8SSHxXV9oY6zccbF1r2+LQw
W34rne23FVTxii/hWtBrbZTtBR+mthcfUP4yfRKSTIVeco7FV5+08JnasJz9fJ/6
65p4AdNcKZnvRQQ15Patd7aQeX4fycLqkOWeVZiV2o/CqU21UpzBEE/XH5997S5U
G12EVevnjJS6dR57pLXoT7imx0O5vhK8ylxRUHkRsDeAn6xly8BLH5xa8g7tmIeo
sz6Mlh20qm/TpU3yhLuf1nhDiVx8k5M+OOS1JVgFpExP/SLZGd+WkARsxyCQ1/71
5AYDWJo9fmI2mvx2mtoN9Pl1L5YUoz8tp7RBWpwMSBYsN9ubWjoiMgONpg1Xf2/b
eIEHQVCwFFNo06v58fubeAhWSAwjjl4oQR1ABsZaecD+jxcz81iYB50res7kPbHy
9p9Ko9wBYVSMMfV9PH5F2bYC+lwvOOSiBPeqgND+Oqtb+v1vEsqYK5K1/AiU1SBs
Pt2hPW43HGfKhpKloPYmWc8bHQarLStMkBH8coUQCE7A371ZKHOIF7bx/VwJUVbb
tfYWL83uLDjd07C+wPQCvoMhNkDFj1jLR+t3gypdHNRsjRc/crNUNHMx1pY+WoSZ
2skYzP8T35/mF13VqI+erSDMsgf5sJUuS5/Qw4tqL5p13xcy17TeF0fQOT5+PFKi
`protect END_PROTECTED
