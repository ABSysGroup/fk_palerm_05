`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uUR7gbct/pSqF4WCoaS8X3UWiXsiXWCGP6lseqwGNPZy+fMlbj6hcXt0WPOmdWpt
/rsuxv6cywjuo7lHIsGeRm7GzSsaCODaOrEts2dH/1D//iPKVrP/TqAibfmieZmG
6gnY8Li3RGx+QhKZTN9cGTgjn+UZSSow+Ai1/BzV720I/oR9JVnCwiHVC2NVzV9E
svG0b058BY3dakSPKwJsbPBRmRYKuiB8QM0kuHUYpAKujKD87nqHZ0JSjG79PNKT
15Y9N6WOgZM/dLZ9ZVspgKXRqVZ8hXUxjJ868jGinNGFvnvUrXi3SREFoSR4p4cS
KcNpOhJw87qTJVyIgn3BLTwp1YlyiJwT9xy3xxkHqioKd2VqMv6I6LKzXug8opsE
A569T0mhEhF3Xul/0E+8Si4t6rmiJXTNIuKXJOAQ8bsNHgR/USe8UUR6ANIr/hiE
QpHVjw9MXmJz5TLfgUZYD7kUlU1PedbyweSUnFoejfaSXYobQjPuGXtJbDwXJ/mY
nonC+VM8bqck2SdLT/2h7WpwOX4LIX0LZajQbW7chBKRke/hN9vA4gSPGrbVk2mn
MpL4+0YQUyiJLuw8sbGQe91Kg91ZEpgW1xd01dlq41/Yqx1orz3uC/Ma91XUJSLh
mItYUVc8rN9jTIVTVpNHOlj465YwgCa5GTF8juJdMFihRlh0ICpPUIXCQzGRDE0D
eGmMF3qxWZx/L686/Eco+7txh99fmqhqLZ1uvetyEerTCHSPBIme+z33jx3WK13Y
2tiVyz9TAAibkURtGdC6SQ==
`protect END_PROTECTED
