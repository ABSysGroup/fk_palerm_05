`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1jw+NSstbrKOatcFfQumziA3L5clpLK/j4vYsFPldEJ8E35/DYoLwV9Gzpe85iCg
UTRyiW/39kQB1IWUU6AA4k8pTZziAMRGh7niPGIrsN/WQeaXMyvG6+znErJPuHDn
1q7hlN2dXhfF2pjDo1f+eXHCEuyfjACFx4mNcDK5Oft9P2fX8BjvPN/uYPrPdvru
odPpT6yCuTYe7U8ty+Ff2JFqrbE7xooWjyB0pT8RAGmMhFe4mbkUmnxS7NYrWnER
`protect END_PROTECTED
