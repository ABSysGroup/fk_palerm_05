`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T8BbWfiTcgJW0+05JcL4Ptjrz19aonlXFIzXVf61fZjKCfYKPB7I2C8FV4XIcy2n
KKn+G3XBG7kNMWgK/lfAQOGp31xOLfinbeWR+vV1LpfAaAKMkSZaGCnjA48kZzex
tBYGLne1cbT4HfShCr/JOk54mFKlyVxWDMd/251sa7QSjQdv18SrWEzdBaTW7SEm
3eM1gT8sbMhlmW+D2wMl7nY+nyk9VoNCxgnxaGOL4trTVjNpp1cWsjc8u2O2aiSy
fPuiLAouDLF4EpuliOmKxEPBsNe9uBjw2t9oRaPvpVRp9YJO4UMYEOSiqwNi3xGQ
eewPvfCjNqk3MKmOsc6ISggFjgTt/RonugZ8mDg1RQoDtImUhFZAg6BlWBLfag1c
RmwIkB8eMPH8J7jBKkG27NnIKjMdG8zHUDalviNIzIPZPUaYeJbxIbfLVQWH/9/Y
V4ACmVSjXtbOykclBfBrdI8wASYdt7AszHxEJvm3VaQaVMRfj8eOCbTcJ3Or3nFx
Si90DRKP2EvfJFhFXaOke05MzQ+BEItk/UH8muCujuxvvDe8Oy4/qKHd7yHWHfUB
APT9NhJPNqYekKICvA1mpRMec/WVdw1ypobhQoL/z6h9IBYngJwMYDeAUrmIHwqe
kqyhZkN6eVRv/h12K6Wje1Vq0G5ScLlUaRoYq34GJRbRyK/PJT6Se0886eMfobHX
lhfpjvMWlEQDbxFU4+iIljhvittbhPNSFQMTO0pow19G0L5eJeqfBd0ojLnaWXai
gvFS7cZToRgRUjEPDurEZFbpy+yRBGvPhaTQOlUihCAucZ3OEC8sqkeWcGkUtjGO
57QvPmORZy58rlmnoZeEOW8d3Toojywv/PM1LEyZOBQlr1pwgxyMHmxLiblnt9lI
qxj2INb3++O9dD8jnGIF2nKjj3sOUSLS40lT5X4mhWeX+F8gM839hM1lTABHxa0K
NXReE1U07ishBNK9iylnabuTPjoOrFN+tot1zwfGfDiWk3jhDEs7BOJvF3YVBrv+
oUDDSFNg++TG4w4ES5lEmxqJhILPV7oAraFT3QXm0ZbbsikAYzRrZjFAtvTFd+ce
pVVKJyApbrnJYAVBRMytG7akCLakf9d+jj3GTlZEB6rTDLpw6EkJaKgySivAPhaB
TPQ0hsBoV/jDB4F5hCyVRw==
`protect END_PROTECTED
