`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uJM6AfTepFLF+SyfXEezy3P18SXLd0f3RzaXeHUUjWkFvnDNdXBB5Vv08Poge5eF
ShlxhN3OAtQMsodKeOoGCgAi5rOdo1ztngaBcc4bjtTN9DsHlnTmSPfa5eoq9EeI
3T93onxyUYRvw52/q04XNadLclDnQJBCLV5oDsePhbZjqBWVlOkELhKKHXaROXMI
KywjkdtkHvTuBhMfRY2vtaFvVVvCitJiMavsQbtvLzvg5W2DRHZqYScmWKDIH+Uj
QXm98TA4ZAJ8LzKGdgoJdGnIyn1/X8kS0ZJjZ4KzwL49p5a6TJBvCOYjQk7Dvw16
eQFdjOGhujJgriBbc/Ky51S3HaOj/Fkd29GvlkiLDfMF14Rt0iRVvr23Fu4q6tRS
DJGefJxvwL/NgQ0n9W1sWaqncL1ZwEmb/0aE4gxGTtM=
`protect END_PROTECTED
