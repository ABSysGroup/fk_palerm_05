`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
baPNNIXL7j3DE8TuXGiMQ7+Zzc9+xCAqnwGn//4CuAs4VcT5JEEEzfwYMJ0QliyG
jqXfjOI0+qk6KuHqUjM8tulKGD8mY+nbN5jAHMWjxjoHf3qABtkmYo5Aqge4nNn8
FPmPQGR8eRfO9cC9oQeCEbGT8tdqqCX6sqWv3uEZ04mpZvqeYr/vqncMTljorvzp
2Ezo/WzcCOhh6E2Nk/5TI/+pkauvXudZ+exSzJkWP9c92Rj0j1S/pj9vyWQ2AL2b
75QodxnuGPIqAMTyy2n5jJS0o1bqJyHo+eNrAjW26ZlmnoluOWuEC3qN2MmvdfhX
8reJp2unz9z3uDvemqNs9zfSMHK4wYFmw5KtChSzD7L3hraRjNxbHdd/hZTf927S
tkzg/7J3PwpS4OOwUe7kfTxGexxDI8izN53ngyMq0pnjAnZE+SNRtZGcGcCmPZRb
9zMH7HpXnzlXEXRfOyYWZGgNvMhx1L51qAaWm2ryaAijPxjHvCyEf3iWk1R3IC2i
xA+WBeZQMoM9hHoQAzja3dhBjP0nKhHNsixUQQEf9LX7W4K0h+E6y6zj7evZqsqN
7O4OBRHdEt805OIzIhSQitvJDNBh2EJgQXbox7PJRStXZ19jHluq+MerQPcJwYyF
FiQY1EiFpoV2wJbw3SzZ1u1cDWfKsk4TJdmeWAn8sH3iQ7+4rZg9FQ6MutxlXIO3
Kr71qTEX6kdh3k5u+Pd0AJlw6x5F7H90HU7g+nJ64IjVyswHODUNF0Rkt+tQN8HD
PdLYynMhnvYx/h30HuJSyHGvwHJYQuIzpIsyGAlW4npKz1PfaMEgLI/28OE/RHGH
3paFDP3VeA1zjhFIUPnT9Vs7KJpxRfVh1saQk95XdvGV7dT6LGnxVfDBR1TgmXhZ
5ImF/NuAc6apMcKLVpoelS0zt269zhO0Snj7icRPgoy4HyIiuvmaKoUwgGFlsokG
wiNrnSUi/Jri29jaqdP+PEYoHhq7hb/jZ/jfIbnUZJejEJXV3Og9R5qmoHYSQFVX
tx4rIzJMkAo1nbebFEQp7myGtEknid4n6Dxfkkg6omscL2C1vBkqvjeyivYfGjgC
STr67ie3GbkghJGSHE5vly1sdQ77LO/AAiNbzc3MyajjJVjTYj3Li3v4jN6hRfpf
wBIzhI/cYsROYrKK3bgHzbXlkmbkyGOTGZlYWLT/Is3ATOgFMeP6n9xYQWg7q8mb
jPqdUbR+XJ14CESg/rtSPlyv3FGjY1kLX3sdiJTu/jxswJcArewvUyvZ7Nhc7UYz
YqMGxmQtRqV3Ya4egYh9lT1V9boez0rwIoBKvpZp43S/7I7KqT/VOSwPAvFDtmOc
yWbr7LChkH4NDaV+sn9PB1OxSpjPPKly46AG+ztRKVKOPkky+9/is0GWPhnh313S
deNOPkUCrvzsidsDp78u3tL2Ic0ncAFj1CI1Reqk+DqUbcJ3OyaYBq+42iqxA2a8
JzdixYmow6LHMVgM8VX6fjv8i+gnpI+66vnfqA6COzEMVRcCMoCAbzhDkghXQVGs
SMOD9gPPV+AFSIYLJQ+HGXR8vuRoNRK8zr6VQMWJIufIeBA2C6n3y8whorzBBBTl
KFts87uOyokKNF50VJBT3iRGMDGyhNWASHgx3j74s8GKeNHe2VL2U/Veb1gWQZhA
Qk25PbDviXlHdYjSbJV65wZArl2KjP6DNmsT5Xjml0cUe7XEwdjCzbIoTZmBNDyG
VdIWrRFikjBSPRGW0FQw68uei48sQbfw5FW1RNtAHbiSYZqTUtRJ/gSUpJqZzThF
ZF6lrHU9WD8a67YTFPWPdFUp14+m/ioyF5OohZRg6IDYxfym2K9XsubQgTQNy/9P
MhFwi8yvPxKFJKdPyTOnpPff5JakJgmWoSUg7lFrIvR5qihfQP5/hWkTjp7JwwQ5
56tr2qpcVRwvrTr8SoI5osIc2l5j1JzouBKgLudlD8YeYdIynoGtcslrdeBPhLsc
1oER6xU7s2tmI/rwQvZGK0V3zyYHoCE/eltNawuYq1t8Zj45u3yPBFXxyBA0uppA
XEVYv6DSYsBm/UHMlKDDEr7x7aiEU2sBMS7yXj3wCn85mYQSnO6V0eW9Zmw4eymy
QNxa2OT6PUAHunXgGtqWVYfDN+1fjhz/e8L6RllpTN5TX3BySyA/TtFhcKlI0mAq
C4TWyciqUE9PJ8yQN67a8+i9n9H7vFzkx9BoaQiuJzn6S4huwc+lc+GjX2yE04Jz
G0ePJaFxE0tGIMcnba+jQYVwB2xL+zprRtjX1GbTQfRyyJiL9ebIx/xK2+Z64xNT
SBXFSwYq5LDMqLdxW3WBgEI3X3rbB6GcF842k8OIrnCMvHPHWLKHef+4rQkPHCXF
HMmmOKxMo4rNEvfhIknCLKv0crROGdHGirgqZnovC0pGa3GgYnd+uotmrALNjA95
W9FUKkL96dQoHoCB6Z4AdUBh8M4z+nhycfeZlhjP2tcPb1NVhx/++SCF0hkKvZQZ
hW5BC8h1gVMpqP6j6NBtZfyWINM/y4nHSpMDWO6IMQ57HXvfPtneV5QKfvyzWP1J
XUwCbStbePbe3dW9vLIxzzALibBz0v+3tQPof76BO3vrpO8wWG0PnV7B63Uy9h4C
V8Nb5gof3+DOmzSD0ex3xqsio74iy7ztm6m2gOCCH5riN0FYGrD2UM8XAhE7MZNm
EpWlC+8PAbZZF+7rmZYWkbVVm4s95IQbk7VFmNRyOIC/PAIyvwFMN/4Eezww3pSv
FvLQawjrmN0Ye4M5C8VmUs0kV3D10ihzhA+J59n0xKg3b2TCxGNBPw/ZCvkbVzio
VPdhPtnd1syE0UHDPnHSBU8IrH3MWL9ZkBeAENwnmFMaoClEZG7m1H2kUCJFcQm+
BSaZ11GZDxcdht3VUJx6oJ2Wfb1UZoPSUlFb0z0gPP2/A5WOprbJXQJY5RTI7r4J
Ia5mqmV87OLuFLUKOXMVqDwqI+MH4NyGu+tAt9brPVBNjpZWXMW9iewepIE0mEN4
vRQW8N83Edz99u67DkwndVIZKogISAl1YoxeV/RZtDOT7IyUGG50ZSB48j0kWzwc
/M+9j/OaSC2wfd4KxVZRIKP8A/F7rhn3V7EEfx1GJm5zCXMmjWowvYB+R+kSv4FZ
P9pqaTxXMnE+rghVLy6Kd0wJEOG/cILOOoVrc6aaGoSDbe3cfB/840gjrtSdqIhS
EyuIiurhpthFhgVJRliHXz2iDFp0RdG4PfqRYvYdpgsPpSFlZ4b1Gz9izLFYxM92
mJUXsMo9rfUEK2QL4QymH4DRq7XJpnSdIFr+ucLFM/gHjz4XqhWhcxYbD+nTK8/X
ctRLCRRnYDQ4lKSCQQoN/sAIS9Pc7AH8z4pGfw/rm+O74MSxplrraCO89pe/V4L2
A4QCErJviTQwnEE/GkggzAa43Ft14tc/bLtlXvzGOv2fo7etFqscAOHPfGvtOUsD
WLQIanw5oxK5jSE7Hd6pTM17WV1e3hIOcSlFGwYx4iUeHGhY2PLK41IEFe0Daq5V
/T9himqJEtLw7hFl1QV1SmWd7807ck8Ymq/2rS4jTn66D/yGrR2ESlSANKZjj6X0
Okd9gFHanBjceomq3NjonhbupBsA0kBQwBMIu04VWipQYxPLt9TTFyST58h73EM5
hfefFeB2UsHCI5hbR56iHOkC0NP8iT1wsbc/NquYHiId8Kb/+3UvYHQ+Gh8Xo8TM
kDoV0F+EIWgOQI6vPDkV56S6pkthr5ZCBhID/LB6SSS2iVTsRKsPbsDi6MFEMjvl
4ZH9UfGxwik7ei0iIAtw5+ShfDWDg89k90fOtPKmL2YhlUZJfLXjaTKoXGFg+Xkc
AU60Uusj52EXBTxIZOQJK+ihzjohkrJZuQUxG50K/rS1Koe9e2oQM8pWtvI4t/sA
CEcyFyci92WW/6INpnMv+ilIlOtnu7G+7cVRocVFTaOsaAi+TJWGl5M6Bwy0boWf
xF0SXcuYgBQmSXp7/KgVY3Kw1ODUStEoJPKyH8WrEBCiPZuM+55V2uoavc411rmx
/FS9n9Rgg/w+WK79LkB3UZPCiNUIK7xluaZM7Yl8MowyZZQx6Itto19KZ+NVaC1e
lWCARa49aFfpa1K3dk6cdG4TSdhjhVTMyGHuXygBISNzuhIymxw6m+h5wDS+VrrU
JP93s4xqTM7lKE/r9Qs/dbySnPaVXiNtdG6u3fcBzAE1nEwGXk8VzuxDPSqcjqpN
UMrkbE+7XcOTfHdc6W3zQuZZiVVdqeH2dX3ukQuCaCDh7j+Im3chz7vJaacNyWdE
kVeRA9lEy60JEqGrzuId1Hp+tNXBfwFpe12YIIPTrncIk8mUOSfzT0Xn8BjAYhN4
ffHPJCC5qbtofv0QE0PQaimslaMsG9UnN2dahNpgpld+x5LYCKl1wOurbzTzAUOR
Cwi0oacEtop9NLUAU9uSdD6bENiynOf8wOEgxgxRdworE7HwDQjwiiNdZ0tZNYHv
+2sLcFGriNCEq2v63Jf+d+QE7JOSqnvj63iSZmEGqMKXUxYit1GthWp30lsiz1NG
VbeQh9Y5xOyRQGaY9pfwhy3YesYKnMsQwt2MjUipiYIlA1aNQaq0XJgEpOM/EiUR
u+xXMrVnY6/0fefG9AsxYoG7XmMOd2lfvPaN9xx9OZ5RPQe6YplzhtN9sRqjsNYF
azmuFplhwfGvDGfFSU3B2t7Rwgp/DS9d+HaEC40cU8CXV/o0+wx2G5L16p3uklQD
VBlHzR3+qWg52bKfNDDO8UhMDtY77KtVPWgjCeSLUpRGaNEuHQKYtxKptVdmx9Kc
/jM/swEYIolkUycaYUEEOe1JpWSJhXENNVFwSWrRrFI0jFuXvxIbSXoxULlXZWPD
cQhBIAQIkvuLKtFrUgcFnIu4HTKu3pjDDeoYKYio1ZwImgTrqcGd6JuznbDofkfV
lcgGXyC8H8EZwbi9GkewXthTcSjDcLnLB4IiSCNzMKoPQAl8PyJn2L3M6UMNqa1M
n0GJvpVoEsmvqNf3XLzcr1U3NTGWabntZNc2uqCT/c4gJYkdJwykemsOxsWUGzyQ
HFP+is6Dzkkjpb+h1hayKsUfqpbqKydYTbGu80kR01d1fYRFidfJWH9ZXqcLQzHL
6NkjQ1uZqc1cTrydVwJVHlEN6UsgoKHiflcft2X1pmIVz1icKvvOnMXzrppIMp4e
jQuV9SuHMzylxZJEQAq3NAz//3/XOiwxg0NJrwaX+FPXUk6JSO0UEwiKFxBa6EpY
vwqsgCqcfBtXCBowhtlcubcF/7GatQrlQ7IZfZLIXhRskylyNPUdp6PXYxIXqk8E
TDywSi0mw/yiZXlT6N4cuOrlkxmSLZcIX6bt2k6s/vkZP+DnWdZfRYkVIBi9cu3X
+JDTUsG/xdIXEelCuHpBDC7CrraROKZOtFRHryT5xpUPk122ciZ0GW/YLb9Yflwl
S8508QQFlLguf+SRB3XALUZg9FfW0UnqNfqo9zj7ib2Teee+pVgbzUgMf2FvgzhA
ffNdivkkN7dyyYHHQmAf/ObDShFJOW9kHjw2NNXCDS6Vs19E667dkY2nUFjSOyUq
tOs31Y9/aXGCjHygFRmha1IHIRZznDyR4fmVAUVU2CNcsQaqxTv2Zng2MCCtT3K0
85U0d8tgUCdc7zPg8ivp+T0hdtAwGzKNweBcdmTXmRhJebilUQbg5KOOPjkQHppJ
XfL1o6TIoAyNbaE1WhkD4xNizN59Eua4Bt2KyaK9MXUCnHFkdOlPBwt0cKf38DEF
`protect END_PROTECTED
