`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GNAa7se9O29dfF5F9C620c57dZy7bfo3eZ/RUu6iW37pfmQbI0C9Va/euYAlQLkI
mrRNP1a/KJ7aV+v8nmk10+QkEsdC2acnsSAapISw+8jxELaK+L1PDb4p5KDFujLp
Wqer1iiYnAcdhYc+4rpwAoB0sRSaImVQsqNFyX/PR54IQ6MYV5oY3F1s+Z3Jr5NT
OZDX20LnYxU3l4msobQnHxcvUWS1e0MiIN7iusnCBszxLD7568D7hO6vSZYalVbo
uMsswqfyjMC6N52MfPjGlS8HZhz4balPbFfFSGH1tnXthsv4L9KT7yLvpvCi/MFW
jdcc2FBdlCwaCHlvRfFRIUde3iJXfkoj1HlrpnMgdAHfndrhOG28/RIZo99PzOuH
aQukBQ9SWA/PVErw8VM5dSc7v1ThMykR3mpr8820+h2t+WJzE4iorM+da/2v4sM2
mG2i3u090tcwZYJ5LOtmAP1zjrIKiP5EwJm7il7gelN8L8EUw6BIEDC2RbzR6pz3
qTZEZmeyaFxrulUoOBNxfPYqyXyRbBFTOzBZnYpi9Y7bDHvfUKPj3A+X7mLAIg7O
pMiE4wb1yP+/ksKGtikVwmXi6ymzwsp63J95G26YtYol2EO8/vFWqSK+XuWiA0pd
1TkyIrOJNuoTxoc8EWQuK1cfk6EUmc9izDqj4jQDQUMu/qlir3i06P6/yVzJlE2X
B8r/7lSkVPb5L66yVnc+zgYt1u58cd0PYaoRZxS1wGFlQ/nfvxLwjzWXlrcYMSrS
Re3dmnyL8q2qk3bZ0xbTKilbRWfqb829HPRZKpNon/TzVuc2aQeLBSOx7e+82YA1
aeolaWnN6b6baAfWPYJuJuQhFkMk2RmmvrnffwTZ5lhu8NPx+jCnEDLSj1oIFku7
`protect END_PROTECTED
