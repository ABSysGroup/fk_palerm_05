`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5JxYwHFb40PFaWfFoZ4EQ9lKE5RkWxTq2DKqP8jfazJlY4hWdfYyO+OIOPwySD4T
RzXWF3gazji2RhCk7/mego+x6NrbBzEgx8QQni8zkFnyqmyhrR35GcktgMkrqOdU
hS312ZExfIAZJtJEQayfKSYNp/ycWygfdS+m0bQm6GGP63kxIP4LK6ieydbfHU9h
XpPhfr0EIKfN+B89nQ8tKGJ/r2ca8eFufq2bcV6pzJ34cMe+TZxFIl0Ax3jHQsUZ
GLW0zD58SOL2N87vbI/UY/CG+F2KsL8wK2RkJmbB+Uli6tdFQX4z1DDGnlc0qd2d
MqpBqNgAvbig8C7HxEhdlspVYwVC9PMN5TVw+y6OnAin9uv3j4zULVBGlTCa9T+0
502iIU2FGn/kPOKVII5BOh14g6mKCClB2MMr1qx+QjNm+mB5ziT9GmjJUxvo1olA
/EhU+4dnb+fc+x0TibNmvWcH+XDmzUuyNKWy/UPVpvikDVIcqwmkLrG89Dcw0K2W
9IKu2fyCnD0YAs2u/J0FYk1IuKxcSGr5bl700tGyYztZ5y9ErRRUTLFrv0GSID19
/hPVdsyF4Ns9IAiOzscLwkmhrszlY6+fJ53fgYIBuCQoiIIX1DdcA3uiANsM2XZI
s8CW91x10wWwuVBVYn4u9AIrui0rzin3+1u9t603LkXMFbLxXzhDNqm3VXGdtKTK
7YJpcGc71SZaK7JQb3VM5THQe4s2KnkE2NVTtRrGASNdBn5eyRGB6bCuYiTjJEvL
2E8VweYyBbPRnpdB/yDapQG61AAad1zOG4oo7CGGm2t5wsCtFHfQrbdMybtMKaxh
eypdrruF9ZyH02vmuUTh/AFVOQEZJp4smKhYELJ6htTZ9EWq77R4F6ywixJABODP
8jXPZ0fT8fm267VGyrqYhqMVWQcKXLAnBAxDsLP+L8WKURPisjxaM4ALFBxQdilv
6mHO45CW/hAFQUPan4piZHRNOieurH76MrrxYgDLq9j5B2SYNPbtlz5XEpLO/Dfu
y6siObj/ClupAz+CXfiF8Zc9Nm9jB1WFPEXbnKmxGsJK23+BNlX7gA/SuRXZ0tbq
AXwauSXMjmeD3ugUQQQ8DstDxVsXiLQEr7pHO5jibwejFeTst8kZfyM8X8uMbe+6
ZoGJKwPwO96W98OvuEttPYWE3oWEs9Jq4fRMbVSE8j3nsZ8RLpRNzMeZu/MTQmJC
cEKnVgWwUd5a54bpDvgcns+vb1iU8K0Gv30s30IUso6MgENPzOI9O5LbCi2bv/U7
7/hzsf4reXcBOina0wLUhDZqyQAYYwuqsYl2+HYe1EH4lZar4v6S6YnN4jGA1S+Y
3OtdXNurBoAiKV26R9x2V5yfGkv8eNKAL8sGisYCM3A/HxnLpDtdBON1bq7xo1AG
aCHqvMxMcWrFIFuOJKpLImF0LHtYpXjwf4bnwv1Kr9bbSa/LmbBjZZrDpe3RdzYZ
fjOKsHSsPk0S/F7KfyvgPk6ppkm2CJM4qhFze7TgDJSRW4lUcN6r6qzFEhRVkdQ9
u8QOJ6WTxrPF1y2SUrSCaedih7tgCcTS8zWJ+9AjOJkgwsmc3rjc7YWzZu3Bxz9b
A5GGhbPEHVz+jeqCA1zcdmxz5CDuJH4IrOzKM8ucnsSpYVSSb+cjFsUnHwDWvb18
Vdy61gR4cW+NSrE6ZMDiz8Un7kRx2Wtm+Q1cVzaZgyQYGCVYu0QfQWgQ6Hb+qFg0
03dSRowvFc+C1+Wjjs2ImmKO5PrUakknG9jv7Kka/rAltc3WhXOed0scM6IoDM/4
9KNNzvFrZ2H8mCTqXiJYdTKhsCY5UCr/0JmGwxR0tOwpgEWgRJULjIBo+QrM9eGI
KvPCnE1BFAKkswW7z35uUCuXf1YaVfR2au7/RHGs/BmGOqe3RAuUp1DqJZhJ/5Ff
lhxSzgyWqT4xJ9gpxsHRPVTvoPY4QJ58A4SRiR2uVptdBN0pxsJJbOm/6fDWmLC8
`protect END_PROTECTED
