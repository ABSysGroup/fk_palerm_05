`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Un9l4yUkk3yojgq5iB6VYQW7A2gKlSJ26cwDNM+UnLxFLs2k2TiO+7ZpHYAAXt9m
GlF4ftZsNM6qwzI8w09xWNVNBklqdswsfPxdZ04QpIbfw7Tsmw+j+nH8sVU4STvG
vH6S8mo93vgpz6hE0DagU6OEqT99FGjM84fv+sZvSaOB3TameOCWMgD8TK0xAGPI
5f8qQBrEsKfoFmR/Eg8Ep/n52pv4ECK0MUvdGLa3QyTQuFSJ+1ARbv3x7yuH/9fg
g6Ldk2RI5ChDWUg+dy1ivzhYs4CKAJZp+OUfnkf0bkPe9XMzsTkze7Wrb/lh8VYQ
18S/WQJ+57/S/dfqqnBkhoIGJj3XXG/p2o+9qtm1qMssm8WX2/YZZ7/KGkuHHbrz
kZLJjjft/j1uiDPJcDJ+bsbz5t7TCZ/1c9MfNiHaT1kTDKeY1mjckS6uqQe72CO/
XnFHPnHM3VK0vbvBND0Fxu7hulQrG4x4ianMDejusAY=
`protect END_PROTECTED
