`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u2BTiKWIW0X1KAxJr3qrC0ikeYgu7SksJzdu2GgNCSqFViYMOd5qP7xfM2Is8eQl
VdY+GyQArtCZVrq68mgwkTkCH1qOmbN9EnFKeq6UGlvfeBhRKzyCbHKcWGYsJG9d
DJJOOEnYV+v614pFPfsP7BMs8ctAnzrqzKZe3V/vajOibrA2MTp1KO3Rv0HxWizb
tyTqJmQ2hGIhVz79uKeWZMGoKzZD3j4UFzUegZePFbVmkWIYQlFCTK1ENOJbMAb8
B62kEfXJZozBUxdfYLWOlW72FBWXTdK8sm+h9Cxvgb2TwW35bz8XdhqzoRmNfEw7
QtjXks/CtEULTv90OfRaTf+Q9bvu4+7fEom8XtCdAAgGCMB/UZK8cbz6FMDE7mLj
31Hkh1jvlHrcLPMC80X1wg==
`protect END_PROTECTED
