`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
riF5thRDRyCmUsn52Cdyu9c/ss7Zpsac6/HPVDFas2wpyHMpN1dOZIJIiYzIUVSp
lPol3/L0/B+eBz2Z+r+4jJKitj8UoG3n2AL84rrniGxNeyyUIjd94jREWcLyPW/+
UGbQLMcvL7t5doWoZaj/sAXX3yB3lEz4BUeAI6PQ6Rtblfii22czeRber6xR//bd
nbP4EbFdtyza3Dhs4viGMLZ+n1CxXc2gemn7xiu1KIRaSGV09ZrfZesGjI+Nz9bo
obNJKjNDyAdagd5bVpuBjK3YNPG3PFWaO6Zr8w423eraC5YMXY+R/XTAhpMEAy2Y
`protect END_PROTECTED
