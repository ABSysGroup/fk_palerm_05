`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dHC7g7nTj6wR/tnYYbrIAueJedcvlpksassLx4TKmWiED4uZYfcN+S2ACJ6mRSzN
55qWgcanzWezdNr8sfxJ+Q1B53Z4KXWnxQ00Ck2MI0LcyuqkO3SmimKsD0168av4
IbmcQ5wPHaHBQ4+2gHc3XyOhtDFYCrsNOw0PG+9w6wKSH6emok0t9KLvF6xrLdqA
BP/agBA3oy7z84+l/TBCyKeJhjxW+4Zy5jvrkzw5yfRIiDyKbBi8N01MAhhWmKY5
7Ab/vNUyV6P9/LxPHoCFYdaYdywPbru9mpiegu/IkYH+EugIxzY6a8m2iEsluKlW
7zQmdRGJjBjQV7j0Ww4eeSNb0GQFgTwgamWLOEmBMDKsxR4+WxY38TvSzBm1rirk
6fC41/xv+K/bdhEX6AQJWqoKy2YRwZDIqM1xYM32lgtFMhu3WGKZpab7JUBsysvv
ocZNh9qNgH80uzHVJIzdRtwA7ZcUQ8984SzY4RyQCob0sDtu+JSXaN5MHHbRBUO8
5Ub35EcLZBG/OTAQOMlES+jF8pPgEKzdcxOsxU8/U4oTkrl5aiCr4qWB33ZmO00w
f3b1eqs+jcZrC8w9xdqE4IxwNoagoKQFQNQA9I+Kw+2ijFiy8HI/Ye6G6Pm9ymbB
bgt4VNaXJmwgAnLT6NAa2bxMWJjetFxngK4v0if9+Ty7EJNbYIxWw2mRqUzCTM2/
m97DYaG3/odWZMkzPhtApf5JWDxeXBdilBZfFCOzZ8BP5NePXw8nnHXOVV3kf83J
UaFBgIFAsAJn2seTNNN2kXgNFu3qWY9lLUboONfgB0FOfttdkSlnz31jcyP+ZllQ
NtUrph/VXvR960+3BRYSDVnGXgFdz1fBkuw5mVADiNkUpi4LjJHfzZkkR5HyEyt2
9tcZyM3P+FrgF67ol5iN40sFwv7djwu3XFsJOSvBSK227g9fRLA9BNAUtOaKassI
gYq+Rpwjg5Sa2FC9Z9TXldgt/KKsjzcRct5JMjS95LWZ2VlKZ1HsijJec80nkGBJ
4wI42+9C0lGqTB56MIv1OLQMpkNTCOHIyM10bUH3TFe8XR5DrPKZwv4NfPGlJBTt
JSBr60aLNHv9r4jOlZZFjC2kozpsIYWuPMcWEDLajHut0s99m0Wpab+O5t1S+rB6
ai7TckvpRMlZLeCkgydTWAfURUPW4bJWvu5jI167XWcBaeK6Jw1k0CPK2iJg5Ajn
YJIl7zIeh2TV//P/DgvMZw==
`protect END_PROTECTED
