`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
psGurzidTcLXDHAAz8rPAyXpDqtB7eaqW3yU6s2lh9YIUMfXf6XwDdFg88aKLSG4
n25Ld59CfAfTs1iQAIe7aKGtSDq6+MedywfQryXFZPlZ8ObROcufmYnUgBHMN/Op
TKhhnpTu32N3nI/4sP1BXZZNXvdzJhQpdyv96/WKmK/cfTpZrQIS7bw3++PbuXDv
+dJA6FvEHBCtB+oTTQX1AvpkBXlgsh/a2G+UvFOwAK/WzHtQUQaeXlZs/TvA90R8
5qCfSJEHxbJfgLFsXeXQ9OqKR324H0f0ERCQh9fOtQ1KGWzMwVb36FMKPp6Sv+kq
WfQ6gqIqQ5cAbkqdyJIygI7ZlUc4kRiKskOIAVOmb/6r9Axzaor1KsLaT7+2ndmn
QizgGX8QLXS9bPf1l2eGSW7quAk6Qs47kLnzYTJroxFqFsS8oXon2Yoom0pKFDDX
`protect END_PROTECTED
