`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
73TPgjHz1eGDDMdNW9E8stF5c2Qw/xzxqhxIOJWLjOw/YwQJDJdf/gFLp53avqJG
/7fqcMmGmI37tfsxmG9RiCyweHX5GojXvEuH+vDprpXknDcw16+dZ+mx+xbefgzF
rlhOwhf8gDrqu2gqXqYvimz7u3HvLdmd3VkBhy97+2hFNY3BWbep+i4qcl86l9Tl
glMzM6yRfsdSfi/ygSGukC3LuzQuwK2jeOi8CGKHKZQsT/utNLHMwK7cCrI9tr6g
gWEGKbgAvPTjUYv+UQQhkaQa5HqcZi5KupX9W7HtatwiyHXT0gPpz+mQxnvAUWPF
R2R5zxIk3Ix+GL8saw0u1fJs9SLgY8TGLwX9mogfx4irMjzuncuIn3NwjedY/s+i
FQIwj7C+d23d7CmA/8r8ruts0PFWP+po7KG+V61tYOFslEbw5apbfDtQASOJLoiF
UXQIf89g4p6inDZOVHmuDHPtm2Bcd3TsulP3pVJreAyGYojdB7rihjiMJ/R/3S+q
xkL4760tq7tqH1ETH8hYv0Q1m85IRGrpvSSFyAIU3WkUaVwiUvvkk8fi1/zzu3aN
JKJQ4eUHL75j4qB+ydAmgEkAhin/sm0AmNyLN//tu3MBLkKjz7oTbibbFym/dsMr
jxmc77MwlFX1Y9YGfWoBmXVzAOk2dKfCs4Wt4J2DdOKvvRuHG16Bo9bGWbJUsDbG
7AXQq1Cj1AcnFEmvvmxPQQA3QumQindtA7zNdMGbOMMbFehNomRaxvfo9SJJeeQn
fKgT/hnFxtSK9cAg391i795waTyCQftuD+sz2ZUeuFqCyJefnklGfPveC1Yw9lOo
hL2XK25NskaPPHtqMxvVzkNWfho7SaqpQK4hqaD3Ahz4C457RSt98pqVb6WEQMgL
MfbCVF1Fbpavv6AJkW0FVNvH5AJX4ZYgRBBIZs5F/4CgYfw9uZpI7mGeAGHZ21PW
xC/biDXnaU0SWH0KQto7iqtNLYY2nCHNiupWjAYd67XPGzxRN+lXOlWjPprTXTtl
HHjE0JdouplgE2ovHYRkbUI1sxhcnlbuWMGRys7xaKr0lxRjBVxXU56INSdO1gXg
dud1K9IIQhhY404MyRAkgM55KNyCSn7bkgcQz9i6Dx9PE4HWbK7cWgTT+X24wv7J
4iRkoZEQp6nB8SiztXNgqYYgtz5oSgYBnvkMHXJ7RUQB9QDPCkVzskbWNTcmPB2l
NqGJ8TuECNuDclBo4Mpn0DPCWcUhvCUj9JK9Ilqi1xDfH+349T+iY5NUCX62UKWI
DyQbrogT0ajA+pEfoOYFScLSFgQh8BkDIY1ehVBXq+CA9jhdz3l5M8GE2H49nYer
ssRocGeTYnUcOVXMvMSSVCO92uA0nxn83vFd0kMjpPKHDomtDOqQ/3DcNw8f3087
mUQYyd8Gl2TbkfidvfuuM/GOvqVIzjBLwuXyc3+sCRJy8qxx4NqlCi28nANmGVll
c/dbYbFSNq3OzFhasP2y6SENDwaCOOst5ZD/UVIHSFq0FHbHQNrF+mDalM4cdVXo
D7uECfWEeMS+iFhdtU40cy684Gh2KCylxFKcR8827WM6/V2+DJm5XMh7fBVhCw96
S3WCpqKXgIqK5rk2C9qJOua3xnYbxckY4oCQi9tDlvfO5K1roVK8H77B4BeytrQm
diGreT0XWGDMkLBIBfyxKgcGpA9n8GtKmLmxdqKeH1alwG8zgfqV1nAQDXCcmoea
jfFDhEY0glays/mFw89wwaPa4YYtx7LdpAhXF6ZKN/l1zZgF7fXsayBuZDVNT2+E
U0UKcChCN8ugfkEm4idsP/bKgRdNuaTfLRw6xCvEMBmTR6ixS5vY5egCkZOm8nXL
Qdvk8IXQgXfd0dkOTdCYpt9fNhgdmK/1UYmPj3Dg2X6gI7N9GrmnUX/Ak4BgjLlH
y9AeaRpW/LMvDAJHyesJHOe9Zg6DyX5yGLzz8xc7rqxYeo6sVZqKxzmclvZ9GpA0
51ZNDHrxvc2iA/aXRU4wzW34awdjQkaKOyaiBvKIoDPNOVa4Ngvki4pKlbTjyrRU
lmgjTuOc7q4ysMoDbc/stGq38097s1MkWkcXXzLfAsyerCR14HUq11Sie1jDxeFf
6wmfd501jUQ5SxEuLCyFW/UOsd0rHylB99JYW9GK0Z65zGFOiOta54e3Ab3w5BxL
bg3Y+3KtyI+cWmhlFD0GPtDJZUmqz2U1yrUiqrhD2XRrlJo9hMSsq/+8vPcU0rWp
`protect END_PROTECTED
