`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bzs8LBC02gbIEKR62aoPMBZq5sfuCbJ+EZyLHof1HcsKh524GRVCkzJMvLVbqYVj
nCYl50CVCKX9s3Xaf7/ZYjPH/Vj59xQV+8uQFUQnO92g0u9IgkaA6hAcVO4GMnDz
jYdzjh6j9biepZwHSTVN8xAdJQ2fecTSSPP92U9Y8BzNOC65khfPae7ki9eOY3LJ
27TXA1ynTH+ta3UJ0LeAUWD2vTInrGmxQdOS47zSYKtX87Eou2CJnY4nXLOU3MqK
rxsvTaR9RMgthgTSLT8rSR4LvI1M6siHPcRt4OWIlyIosutQQl+8dYQ/f3GFzIcA
8edQzAkefyy6D6XgXogolpPVQjwzYhsWzDaCiiiIOZTmPnz8HBGETcpBv04OE5qM
2TLPLIqfNZwwFXv1EkQsYeT7Coss7Zsfl8p4eDZnN+ndVU3ft0AcHIQcTF+WGLeG
d28A84xxOVoy5O5hmGmBWo5wr5qsiYlkOy1o1L4/WNmIczMWKNm0ni2k663PVqAV
f2jkWvPztiM1Nlr+1U1iRx0DqCi9Ibcms8+GJuL4hjOT0PdLfdO6PSx9fsY882qK
YmRuwKaEHarODJZFFTnj4Q==
`protect END_PROTECTED
