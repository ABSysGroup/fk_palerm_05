`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tWRrw9mUHJFQebOouVq41OxJU84g5QXQtuPoXxCAdjM57TqpiTaCKhfWyzIwXTI7
GW0CdLiGpNmljpEcZA2j4Qry1Izh/cLdiY7F0BLkHKiidC706eZ326stK2p8/NOK
HFUTw8N97+TssU2+9D/tPKpnbN7wuTiND4bNeXRIKIOvEmGs4mc98PVBvBdvKW32
tLXyqUcHf/bjghqiyGrgOtN654prQwjJ9Ibf536UD6VAVU0UFoL27WRYRLZZq9lk
NoaLC5KqgUzVZPaLTyzRTwiY1LwrQv2rP7CWlXkmkca+229WNI6vs5V0ONt9+xIS
AJ/qc1zjdATxLd8KLRpUeY6vg8PmBtjQEC4PR6YspI1y/ruZemTHfRJ6Ggqn/3G5
XBA5qqLDkC1Tsih9OfIMDQ==
`protect END_PROTECTED
