`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bETDs0kFgsOMRJfhGNRzqod6neYmsXk5ojx8SPPjRhlV2WbM0CxGBdt88rfW0AXA
DwGjhGWdmXU3gaiOa2Z3fxCFPpT/Rdpy3E54lZj3OixlXq4Zw+MKWNSUkgs3+zBg
XVLFZ2uXFZzAtv01Er8d41wZVr130DB3ULSojDn+4CVbhMRFYffqsnsQkSMpeHIl
gk9rUJ6xlWXUcFbeYD3qhVTpWhSYYuAYgv9TvKnOZjs2Aq3BmLZMHMVDcBbFx2eX
+xVc6js/HCpRYdXDK2XSqgeGX/hMU30yO0sU2gYsYbA1DguXLzoQLyr/esgomh5Z
c5wblLQmW3oqEBxWz3SVJp/GwrxhIENpd7F7mEsIaANHfBpQube1dz7Jto4IWAHB
DLPxQ9uFLdQUsexwaDT091baLxlgWX9zuptMtNPuERP9q38fLnEbNi5+NmwI3fPg
6YrWZQRhVgF21SKa461bUS7hiTrUQBBT8w+ZMJWEJqFjtPxcRQZvPMMicnPpWOO4
6XfUSYZ+mExV1ZVWEuJSvy+OiUlVhephdqJyLIyDZ2LNmH0vWdGNJJPbAsqW2obt
Sio7GempJ+oeA3eXLv3jnDzhlZCRJuWh8JtTakkdEv2gT/7Mibq34Ri3XLMWTWD6
a+KowdxidSxVrleCTKozvbLLMDuWWATroAIPQtR0ev1uafSkdK2gNqDJEtswcsha
9T1XvpjeHXh2ImqYnWb6Yq9FoGgDwICplCo/e7leHktx7Ds4jwN69HWLSViezGcB
DWL/xf0rpoPJ6/Rk5Mt5tcFQdUIUqILZwiEf+AdMWindZhVsqI6Xdm5e7BqSugys
JKgzbF9fs2avvjQv4nemQxayypdSgtgjbg3NF8w+pDcnmdE8R24yMo617Jp8gQoU
EZ6nLsHuLUpNuUPAUqkVOWFlXebMkjLIIbHzR2+tMeN4AXcJFJZ3UiLl0KVM0TVC
g4uxasM96d324lr3LpSM7iCR6XuINT/OpyXY5Am3IQC6aMj392PNtsW3IMRBZX7U
5b19V1UjWapvrLgT3NR/Uf/P5TGrFN8NM57Dv7RCKdIKhffTxfBsK0DIgnh+Ez93
6ugIpenNANjrAw4MS2ynvqJgiwu4wqP/xFNE/fmTpphySyVDW2+CUYlg6017AZ8O
01h8MgjLGYNmPkpPeheFyVmeqUtbhMGDOJg5yhvyLuQupYkBur5lrdZ+vT68k7g2
CsG/5rNJByZkR4B6VeXtj3gjOn/rpLpVVwXXcmu4DNKHUOqoJhsBHeItsS3TxFxk
kuPYxjlx/0eqnKsxyOJf1/w9/Vt8f1mtSTZIG015L7KIk5il/dgtdznpObQJAKrx
bmkcoC2s2tRHFW7osJFowNBMnZdI3uM6v8SWUHrcP3e5EEeF7HHaKP5vUlEaI9AG
5wSLzGIwnteIZgIO4VnCTNegs27d+sGsnixMRTKmOQhWC0m6F3VULmQIJMv+X1QR
Tf15HgJZjyEz7SjVluPG5w6tqrtQhtncW4X4xIfUKz/je91dxXi/DNdUD7cHO9t4
DtojXTz+Z8c8mTrgfX2f4rVBlIV+RXfB0gd7clG7lrvkABqezsHqqctS+qTOq9BW
2wM8lyuqc/85V1on/O3LwxLdLb8V/+ae61GrYzbiz6ok+JqvEqSpOJIfLF/7x16q
0vKAByA1J9gJ0twGe9AyUvd1uLxLFB6yUPlJH86CqByWPmkS92tBtaTTWkC5ISZ4
ofFqP73kZDLtuF9Inxq8wgyool7w9JJZjaIp/VgLv6H2Wovn4k/yUd8fOpjqrMWP
xjhGIuBukAa1lHldp9RdPQtJ0e0sXNm4TjYGTHzobQXDllAd+QfnNwav/QKyBjQi
OqQehesCQdW4swfuB9dW2UJ7edcBXPK0fIvvlu710DfNLUomg/k0zYl0Smgo2091
lH6ep2k2YfIMVZx3C53eS/yJDBVoPAeGjf5eH/nXVIW4Fu3xWa22katso5IOjkwB
OgB1FVUJaGM10up8NcbccANKsTK/1CjhGNI+WcyFOpycgjFUH1G72vPUFIRy+e+Q
0z12owNfD7i5FA/hGaj7Bmeb6nSxhxTRm2aXPm7iXWhJME6UyXguweyaKr+reOQp
kRjZzXGu8UA60nwlzCWytspJKMbFGlSvi87nly7cociYcY9wYvIyB7QLskXKgf0J
8quzyEKoXm5uigL/yg6XVy7VPXKZRTAXzfJMmawt2VcYozV44bd/7hNFnYJlLL7A
z0jB1YZ8TyEvRCAbs9eU8CnQFxIBPC+rkEG5h+HJOPefDqsGgvalgPVbKCoZslm1
aufTDQ56X5CoUzuWhDwV9dQ1SPTAclzgkgQtUHhZkMit5k7DOvyRjjiJoId0WwJH
qpmJORzT1s5IM/IKL6+DtlsCGbt2sWMknFhkzS8/ZLnqpCm1IDUJUYvj9nyDCvuu
uktCUHCw397BcewbxLc9GxBWxfmZAqDezpp6OxWU80ipVVTjmAgYmVmRqKJju2vP
jAO/kNC6ph3233dITBulANGv4VeFZDGiDiDt+ocr80EK7RhonfcGtENe4VdDiGw6
vk360iUys/tPlEY0fajd4/+9tceGAbQB02LIvO0wybHFzsYJ61Mqt6qCkCI8tCbu
h7vtBf4NlcHOt07+iQYFb8aDYblt+lC2Oot7qVn+GTIcc76BZrpAp/R+aNy70Spi
tAStQcGODcQIUoLsCNcceTO806L/J/+v1FMplYBhDujN00c7nxq/HSKwIvu71OjF
J4LBJZbSgzxZXRGBjs3y0ZowATi/FAF/gCFymqVinJkYHMF7i2tbNO8NnwkqA24X
8PUYaxiBLb5FDJMdM81vfHiS8K4QEupx5hhfSDQmhyT4vpjNg01JIr6vaJCfFNFz
3FIOTECc1BnecDiztw1UPEgJ3RP00I4+9QS+yVBBrFPI1EJoxfrCjXKmFdH0X+i1
0D59tyAQqQ94VsGRQZ0byLiqWES3Xz8aIY6wrOmU+gtHe1lLDSqOyFqk/baA++Bo
vJRlu6Afww9VGDzt6JqU3j0sYblPa7vHW3kYNrfaHVoqHNDPU+lLpLanQ6XOn8jN
uTBrqlpstgF/vfeQaKQEddw4K7pDEx2ryF3iUC93ahTJ1s2qrgPIOFp0daeH25bZ
H/G9pkU4I4KnnV4bFiK4MT7V4+7RD446sRqH7EOW2VshbbJfvyGQ6KZ2F5NW80m9
Xm04jGyiQGERaKFejNpa9APlhb7wav0H1Zg8xmT1GhOymH47RGSH5COV2N4ai6Lf
2h4tdtLEfNsgPlq6Id0waeplKbYvl4uGPh59Zkxv2BYdet1Sh+qltFJ1TqUIh4p0
2FCLMtA/VVeaeIWohglxS4TO4ehs8gWXta/m67n/R+Hd13d9E+QnUiTQfaLIYteT
v9SM6BwxawOzlqCEpFR1C1JiCFsc9Api+6YN0BRJICm9g7s9DU39IQkf0cuVDQ2G
/6bS3rBn3zptxxlhEOqPvuMT7ROIfcXI4hM0HlCyVaKKn0PAm0BOh802FT9LKW4y
vt7yzkD7IP8oQnvj56X0aMiP0kiDtE9uILkk9VgQh2DB12Mo7him8OwZkInkjMv2
xASI3Tj+d0SPB6h70HGT3TFK29As8nIP1J+pylUBhwhx6KQDcGvazzawVgyQIzON
yyvOEm/bDWRAjxP8V7B0CUDesDQejWkLRD2habmTbc93pXplxZFW0uacTeBcYMgw
5rdLLPGO2HiDJFEOPx4R4vFgg0izG4ZEmt80wGt6kMuKt1/a8rCkGN3Y3OxegIVX
ynHv3+z4sMnNOwoYLJFRhmYYThtg+pRrwAXQMpqkl3rHXuSewHYMeqMg8SyJmbXb
jYM0/CypemF4/q+xUwoe056qbRTlXgBHK5W4Ek28IaJ8hJ+FHzmG79CMYYkFXZT0
HEG8leHgXmUh+E2NY6lNGRiJSDA9vQE5FueMbRNCzsYMj9nCKZ/IJ7I0QOZD7zpe
sbGAjvCcYgnPHCprSDOeYkXf33XAAfldVu+dpwN4ykrbfQ1N+atjCDI8Nwc5JHPQ
Qkd1mqo/4mYNZh8fAHxyZPCSIWzG6UPMIMToJThAjoxNMOmEA8jRTAlv6x21Zfrh
CZhsL91gCLHDHFiNK+7aY0Si+194UDUiMQARFV42kDwy9loXhYxskgqhpz6NUvFa
K7HtoVahQLFAa7+qN0pz4JzPgKGrAw4F646Jd8oqvn4mqlcYD0BZgdtwZu6tJMxd
oG4dROAJI6OZEuddErTdHb+s6jdHhJU8XzRvCNrR5zXVoXcZ6i7nsVp6pIoW8CeB
dg7ru23GyMrMcYsAt0JVdzlG5YxtEMznu4y8tKwES7fbTxRR8geCWG8Vyqzp9uk5
oO0HkNaapiKd1jcyYKVWkGXzWIPO/saddpxbI8jp1ZUu/4lhmXVrHcFkhLzeRlJE
h7I6eevFWA8HiF2PnIAxqXqotPxSAtpOlGa6FL1TJdZtz9V7hInWq9L5RTn39mgt
mzELcNGDWlEaQDS6mqIYrkcyAF/d+L26d8TI0nogrXD0w7i58aZpENM4+3hu1alA
KFoDWfojjVTy2JWIJMfxdJwlBBqVyvKtaPdvxkbT9AR3vO9GCdivfFN8CajJJBOa
FyITg8nGW+2tqCWRzV00GOa11RZ4TvDb7CTKNqmXDKc3ImUAffUlwgA/W2VTznzH
5Gp50GanM7Cc4SrqugVvWV7Tp2lLW16pPy2d3GJLekua+TYniaofaQryBicWA4Jh
Qa6F8yyR0JvFU+o4b1OdbzrY0JHDGOnspKdt8DTpg2dnaCfHCychCVMvmLAIaLXW
mShrbJzjXBCXquZuOphzSNejP2r0h4EovOiY9LhEXkpCyZ+Clav/H4YkaM/ACnZN
VvoI86aIHjzg840ehrKgH5Oa/7srDCk6uFd38vBhlPejmnMPMhZd1vf5H6WH/IQP
tV1PSMf1sjqNblhCfEKMz6gpsA8fbBdNcNAA7d4DuwsGh8pe4+qbiYXanbzG9Pm5
SRn/mdThQ6Z+OJWLvzQYxKeE4K5A64Ljp0fdqsXxwqZQMx+z62mvRXO5nKpnzmHF
epraXpY2dRH9FWENtlsBrm9C3c4AgeXYtHE29TUD+jIzXaETvWTgetxt/oqRMuFE
gJetwLpfGZo5UvGC5Yb2Iru/P0S1/6fa+aUk4wyD6t5kzY306mYUJ9/fAF+G3pBf
/Txmv5ycSOxEsQlwWU8DI4VTG72RkHMnNifQ7DFAI6DxZzfs28BrhX2a/35k25oM
UtycpeDRS0Ycxl1Wj1207LBfg5k1Alvj7hWt3Db2qUaHpIGjRfyqLcos4aVW/QVQ
l24Mh7zgDoeaAQ+OX0m6G2r4IHDAPUdaUfGxtRRv+rsZgOHVbTy77L5MupwQT0Hc
JXp9ODKteOAecdQXjmTU/auumJerrdHtEJxrm7jD/9AxXP3wfGMiMGOJfftEMDMZ
NY4xwfUj6hAwPSeOzHK98lcataoyqRSPy0QOKHtbi25EChnrab4PDvh0VWprS9qB
5NZoTAWMG+huuC4tR5Y6xvBGgOBVBIRZXqKGCj9KfSBrRthyJ6rGMnuS789lpuOV
bfN7AE3QrvIXgQZhyaA+ec2xZKgA3yUx3sz+6I1GS21rqQWvmCPLY+wAQfky2M2M
iEJ+4/tnebltc1WxFMfZzMymact20Y+EVZ3JodBfLxLbl276JSNeKZ6CA9vmd0hQ
22V+7rX5RbBU4f09VaTCnmQdFTAbknDom2Ni4gA6wB127jJYfi6Eidc55MsgyTFA
cEgUqL85zVv8+geSqYbtxUwLm/9/2+Iey/hE7a06/gRawWJECW/849vpdmbVE3yi
+A6qThLHPf3ReBv5s8aSLIwDSkwq4V9qOHjkfi4McaOppStCTYGai69wWRORHcWP
U5TKrQh2eP3NxxXHjJL3oXi3TDK3YJ0sSjiDLYvqrJFDYBsscz59iLnt2sSAFMqc
5A2QpyRL3qAqmSrDGvKTUlsv/1i/JEkiFlmepFv9E5fuyiccRIo+0nxMHUFrv7qw
TQQwitvycwF+xE6SuKX6ln7w1BWGo6WuSYvi79vm90zsu9chB5NAdXasnUACZCvJ
IJl9nh04/o97A/x0MBbTaTEKSwmHK/mkWEsfyDsqCWbBsfiqo2yNm480xA6U9eWm
Sn3DqZECiMFZgGgrPSGjOe/H9nm+XXm7ue5LmmclTtBO30Fc28kWjaJUK8kc5ZUI
kYQLl1WAdsXxvYyswkmhRa14/0JK+kGcraSHCacOvun9U2I8cKR5YhgY2uPV9zZS
MUtvmPYttBPpdfLjMysez8lxolVo1nWuI3GOkCtRa2Yxw/lhAidG7phog9udUIJP
oxCa3x5qBY7nKtijuEPmGnwuYw7NuGEVUQgyP/YzEQ7qIwVWzNioYUXfvnnrN7pZ
7s1L0fABp0u7Zbe2kuJyT/lOSK4mZE+N1Dk+0Am9ICdPuz9zny9uEXyL/gna8sjm
xeFaDGJDJneUzMGoxHvCdGFPkR61ALDSd/zKRcdqssgPGU0Iz0vagg9nbsfuTMZE
0sOmKPztl93JYJz6Q9mRc5P3I2FtKQrYymaEGJVpMGF0QbPmkDU/BFkzxmQeg4jI
fO/LdJQCwj7iQRzVC4btCakH3LiwkWD4Bjh2on0XZNymal34jXQyHXCqSDK24wvw
uJ21ww7X6rv+TELTlKqN4y9yNBWY1zGOS26SSP+/WDtVXjba7/t1rVWpIkMypnIN
8ElMrwRvU6iHm58Fxhbi9pwLB2Cb4zwdAA4iIKC89FZItrnDRCmeL3q5wrtV+pLi
fW8PHLjnHU71aTPKJMG7HFwgPskSauhvJh/7yY76NannB9WpPpHje81jVzQhJrNr
jhKio3Q0erG09xltND3tx5TXgtze4x9yXZ6FUiibyOzHHLrNOHqm+kewHE86lDLp
N0zPrPF74GKfZ2qelW84uOg2/4uM35cFbSdXMQmgID6Qg8ksAqnNYNMRMjGe3B2k
CuQdyxS79Jx7lComuzR5+xq9PCzcIARi7fpKKI0WUs4GEilYzq0bXMZglme85F6q
tj9X23AkJa64Q0fv9gEWuT0ai0xTd6w1BQtxKoAjaMEVA9n4UMmvtIq07Qhvf2G4
nudDwdVV5yvoiV+jUgBvm03E4xN1X/b98GnPLQYjR2/1WJyES/17cG7HmMXG17ts
SjRV66VZ/WYUW/qZlve/LdBG0Hx2ZkLC92WqpuUI5XVCULr5S/2sQTbdBI4nOzau
UuFAzlzR38M053o2DPeNKm6v90X0Mda7QLrpYAaAvpn06Htuheb6CLYyKobnKHkh
9FlZJkxy/MsNmP/EeWU7QtfHeFq1O0i/xrdkBwGhFQIJhpaKQ3i6/HyIgu2CWu2x
dXMwJ02kVzBHKR5/IuLEdvZdkQ38dZX5YrEpwDUzTbGi7axpaGiwXHQpoqRQjpKn
5LghwrmBJzTqA1dV8w8AoHJoenhS3JNY/cHs9b4QPFQmLG8qy/BQWtDIJDM3Xljn
XayCV9hqFJbNAZtCsvLu94fE7j4zwosorSLt8vibVT3pIjBMvGIBOJo6i84YyhXv
gQckH8L2mPk5awrT2bKsf+RWqDjsLAVuRD37sxYQS+o8+szRIHntzWsQ6ZDPBc0p
CmKT9XEMHp/QT5EDWhvkGplNypv1JrSReiCvhhBpOvhdcCPMtGcg9VgmOAETMqnz
+PWcipbEliPhwKS+/IrAvwwHsDg9cFbLdBygI7kV6aOxQJvXmSZ6lwmT0H7hXDof
Fa0jUWdIuVoBszpHjsWIL75CfF2kQu/MPRaNIBahFVxvB1U3QW6qrkfnt538BQqV
jq30HHwgZrPM/cgFsH3y02lMldt9OF3/fHyirfQ3bOUjE7GYn5N43Lbam0MPJjCo
quUwJjpYQNRGcbgihJeGgrezWnrZXpWpyV12z4659U4H4x1vBMYQZiGGF3Cyfb8r
qZtWka+8LMoIjqBnhAIOT3jsa2SSics/iSyu+5Fz28mpSNRJuDqZs3fGdWY5R8Ov
PjjWotFEL3622BsowzZvJ0yFrkWQG6MAw8dvgc/ffdb7YAY6o2Du+6pEqTukN83J
oJhXGVZHy35apaDPBhTpUrUhQET9WlaF1SoLFGdJSHZsNApVf6MUhbz7BbBhdT9x
94kDCjvJrFFygg+Epwfwsl16FhEO12dsGJVOX3hVzt9DJi7UjXqzw36pXXiad5vw
mCvxXyOWYkUYbKbsSgJ74kaGGXWiJXV71hj2V1Z6Cpd8eO20FTd3mfpx/WNkUwA+
HIXHTgNiyHQYytAbM4OyoifR4uEgHtrGl7xOQvkUnUveL7uYK0f5DcG+WCYAGW84
ne0qRYV5piSyENAqHOGzb96jK6y8ZSRBjxWq13lSQwFWX5NEBAQvyze5Lkg1woAr
VAGkB4/ormJbAM0ISZdKhL8dgBqbgSQc5bK912Z2NdvVbKyn6hhHD04GFUJ/y5ZY
7I7o1foToqvMSKgyr8LVyIX4E1OOVzgZ11Bu5yKgrziOZ6n2RXUNvq5dkn4RRHFN
AiUnPCUeV7AgBFo1kkvw0ZS3Rk2HbdPS0h0DaxgcyHjM6l7+84SS6t8SKTdhhe2W
u7At7zjuTvOv9OKC0AT35uONNkxipEdpUPrhZTV/hssBvxlv6CICYIin0/fGIkS4
BCRGZmna6QrRZnnFXQat7RooO6I/0B89JD06QpISxhmJQm241pP6fHBErYSbWEjH
oUC6G2W9hrrer+d3uG7Lw2Reet6r2eVJpwHqFHa68e1teL8uTAD5AkBZ/2HjScB3
3p546kW3XjnR+4r7aiI8zCUjKHQ2wYpnwNx5ih0gF3DLSugisXwN0yAPkcrFZv7w
Lx8XQUCFVpRstuq2FsSWVFw5soDSumdFQavnjWodiSoFPeZX196pYszx0lO5zPk8
gKpgmA3r21zoQxZ0stHcDL6Y1OHYAB3UsEmdp3pdhqigKiRXa+o8XJB2qcJnLD91
FOJx3wwvjGpjB0SnqCZkwFHAIVP/umAEh1N+S/3WefVE28tzoF/TtD5MODWfRWKY
f06PiEYrJ5kmDiOGxDWi8TklGI6XNL8dbmhmlUmWjQ1jycDCZrN9459QTyrADlVW
PZLPD82azMl2tfqSrRCV1qGmL1cCRaDq3+6nQ2079dws8p2xIXarzbR97vnPnDyB
bNCwovc7N8p2YQvu5UjZcWrKLOegddg5W8Rxc0CCMX3YS+In24mqaCLK2IcH5Ucp
Iuc58UkwNtdMjvLYjB/23CuS204Ua0GUqajVxUWhQYNjnPBlcap0ds4Ut0p8URPj
Um90S+0Z5pu0n2JdbWXFxlKLjIFonZatKRNXibgyjK6dHXXSC/vHjQClS1lWC3dO
ggO+uim/oiqLGLnb2Li8uMgbA7Izi+NZeRjol4yLxWLVzqkZD33tBDU4RLLDTAuD
oxjy6U5faD49ZvxkfXVmIlS3gG4DoS7Nend8shskB8mTVTCOAbIdpthr1L5KTkvd
d7vM+s8LpHjPd1Ypnr3U6PyhH6Mw4v5ZWaZ7QtCGFpOeX3HZ5tldW6tJdmuhV9C9
0P1XAs8qJG2A3oQ1QokduBzRSPw7IFT7zLauP8MOaUrXMvH8lp+CsT97vwtUouNg
79DnpqW+CxbarvpKSRBv3dvqrrqsExegNeQum9SFUfdWzdFyQjlBvZpQGDpumcWP
x4yhYEUGIBgHQ12wLPL0xGzYTkS4XUBSEQx/T86iaLqrzOpqCYHIQXF6e+UM6Wio
/AbpFktMU1QrSQEthKCud1ZPvg4kAaKo0Eb2bUQaDS9IVcM0eIj463BB9JC2tMJD
S6H1J0u5Vf+mtdu4LKAaNbtUgQmm+m28VAFk22WzfuOTBy8rFgWMpEC0dVGYZtiL
gAtVLG3wIKnGpWburg4FElNxQetO97BqwNi29ikCL0/gMHyU1ll6D8HOo7q6H7iW
VwJbs7EFLF2kor8L405RRi5KHpirg2RcalkpXZRjgRueS570bY0fyCg/Xx+hO5YF
bYo1qYBKJD/suacXLW3h3eUscoRmvLhYdsy7hNKLpfpNUcbaaeLdY98WZoPzP5Gm
ZIOjEcWirNzR0OWCoxkT5vHNRBpCrf73ZICWRfmaK1Z/4eEqlkE8SFNFuCofs5Z2
+SLps/zpBmDpQvJUwp1aznyWfG5Kg0ZOJaYmV3w0BU87u/Ja4d+s/WlhjdboKrpk
qJg5fE78CHfN57R5MrtYCsesTi2D3Ow+LGloB4/viMfp42vTzwLwfaznJ/xoZXyS
pHjF25g2jTSL80OWff21qxDuirwIoG6SJENRWqryEO3QwvVA+a3jEWZBdYnCDsTg
NI6YfPH1jptn++jrRTPr4No9CvOm2Up7OmCagUKe01ZG+2KI8uoGZWG+MVEwTRfK
b4p4INfZHVXvhfTamK+5rhontsIA48woTJBnEjAdTOi0hVglbeDYR/47INhszMA3
mTMCRa0+abTEFClqEUWPCuGvRNQQlio22Xf5PjQoEm7ENcMzfKkR9DknjJYQafYS
3JZX4oTgTZ1k4qnRnFxlrsHly2Q0iV/52VE29HKfJhoec70jHfvM9+yIuJRlbeaE
dpm88TavgtxpkTm9gkyNE39r+mnJSqTsXOi5avI2G0KUEea8f24QKUSZpN8syBs/
eqegtK28zUvbD+loE3f16zs0cNPy7g/RNuzziw817xg/CVU+3F+sj/6gEPvfWxse
SLEGkP0gu44KIW78U7ChzOA3AqB+HQct5n8VhzBYk9Adav7Y2x+3wrnYLdJp7OVT
QJPtzueQgAp4dURe2kHu/SPjTJ1Z3X5ouj9PFExeMH5VMG85BsKVI4ZXVNta0gTW
QCsJR/aSgcQXwXjWL9JX3exOgiwZv3oO4Al4nPSP9Z2zK6pV5CK/Oh49zWvX5ipQ
FMXm6tYJ5iiLwjQZfBQlbzcRat/j37TiEYlQXDoUoYO//gdD0qfqbxxAdEprgYzk
SLBgyNcJ8yIXQpDVou6zlpFKDOJMaQatdccmK+zze6y5F5ZjXfjo0a5jQV0K+IOm
Bq3NbJRKbyH1pJF/lAenjrttcFtYsluSHJu7YDM0/kC7ecpjx3SR49z2bi0+Mt/Y
4Ajd8UNfQjIeoQFRY/ffut+G3VrNiCAp7KPAMRE6MGgKLMgvxx/sR+O5INFihS1H
JntLpXLYB9VcBu2uceB4NKSHspuYNJWzV/bzr8FjiBG8TfQg5wXZxz2XtFb9yeqX
OMyJrLEW3tspZjkAJ1izcIez0u3TN+ETunSBzpZfZu7Tv5bXqqkWt1OZooG2vz6c
N+LAMZgRCyD1fTqqc3+2S04c/2Lht9TvFfCVswm7v/bay6DXkBukjGzcMWkmWaAg
Avyh1lY17w1y3U35/sKdHj0+EOUv2VPyTKhvr5DQukOYuVKeOwUj7FiL1hgX2LrN
65UwhYHWUVwv83lHlPYHxzYaozReD4wxtPX07zbIhkdi9UXz7tTGqJxQ2EpHQH62
0VvXsm84GVyaa/Z5p6NvH9eDHxd4qJjrzwwaVCRzrnO5GnXjJmzyC8MOZI4GFVlE
oSNqjYk/EJm6Rnae2eUIcOiPP57HwpWK1eVJLafiDf0EGlyk90l85UUIDt4wI8Ie
vVo2MjbAQP6mKPa6/nUoX4Vq4R6uAAa6cMvMd7K1QZKn1V6ANByi84WnmuYYH3fs
t//lzZ9qvErrkD7bYs3Yl9bD60Rpo/1wX3R297Pm5GE09q6tasPkF8pFR4ysWPTi
HOVj1jIDXW9qiXZsmzsFpmekiGj/8O7yRRbD0LmldTlRwAB+E+hwT3Mj9L6Z3xGe
yFQoNdjosc5pABF6VXTc7aJ4qzvDmcpxv8wbBTCdV2GB+EUKOtTOpElpwiLiNSCK
uwddjUnrQ1qxJeGuHHeE/iCK6YcgVAm5cmFrscbkfwDGsFYKbKgnj8mvUVts4+ij
mcD46TxKHM7+hLzGoJmbvD7juTlXu1Ttf9XTYxQR5onr9qIH0sGE4d5ccHPGRZSU
CEPSLRF7Fbhw9ssGqqJ2v5qTYTPU8gcS/DNujsT6QcWOswfN8te1dNyF67FUiLb5
35RI9GdAuN1eS1oYkmj2zIGc6t4zWF4i4qewC+oM/lxpM+XYz3Z08AM7tauzQYXt
EZW24YVc9CJBQRSYHlYFJ3IBdWt4wswBAVKaLTvWpbqW1S2KBKI9EHoCitMZ1eEL
Z1iKLJHdQnE4kzaldefn4DGbmN0Gd7pHYWag+V3lQVw61A+/v9rACg69erUAldC8
+jX0r0tE45uyQ8Gb3ZSKIqFE0WqR8hmevhzCrbdNivAyR8K12OVRDR+cgVEl0sho
DyCsYfKH864auW7ExaqdP3Apc43UTh6cd0gwC4fXmKbeBKy1ge1MSZlR6mW+NlU9
JyDXh9TdKPwMYo1MI7LkeumZgfYT4941zB6YY/2nn4flnXPUajPwMUBEqrzb7UfW
5sXjenJ18uHBoyrHQk2+He9+MI+SkS8hFA4NT+bv2AwSbJgKl/XerP71UAxP8nQV
vdK2Uh1kNubyixYmiZKUU8dJz+kGNxlPNL0NFx9NBVAnVUD02YHO+2IIp8tXdsZ3
lzaWwqbBanm3vnHMc6NTVBN67FTrd3dwqmCm/P+NViNBa5AMqXOXaheo0Nni1Lfi
VVH9QlBS0oDP9x0VjJ5yNadgPunan6HyNeclmcq+VnI+32/L4KKh2fSJsCnt3VvD
JhmlUi/NKG5hhCpJLnMQQz0B0726uQPCqZ5xZ5/EG9d2bI4LXPUgUyIIBateic9F
DPaxy05i+xEuiJCafBFKBYE8yCmIpI4jTFOTdJk4ltHTYldbQW8Yo1y0ZmE5czL6
TPG6e6o8FiCDKAKOpAMNrgwmLyZz13Fk181SHIYvnOpgrGr50WmWcoujMj7+EVtb
zO4nx/wBFim6l2Lo1uiISbJiGfpA7a3Mel42ARe5blCO4NlNBKd1iJQ0mRQ6hU6T
cI1zVrGvqYDyz7dfk7mmaaxEByK//pnn6AZF6ceOgScoE5zhfPSnS2kL9ZnC0VN+
Ed0TOpxK3ouefhg/29rayj+GQqtU50fFUVAariI/UTtp5O4noShgpMvzYFVCdJQQ
D5ZTkPKGEJcvF7Y1CuDLNelBG2ZAfMJFufgDu26jPb+NhN7ntdoI1sLEMIuGQLSc
E7XqlJrirxgCMEwnfGu5zfLBlpZ0yPTsYzDsvUxDxh6qK0ryY7kRMqeIfS3sePVG
jrC2++KtCU/66AyxGdzEnhwCovAkyQvoeEbPiYYy6Wq2jih/rl+biW7A9ViT73O7
SBKXKiSrgv5yzAZskhr+HSreJbkJ1D+YzRwxoJletR6tas79Nuc1pu1aOJqWMBrP
1t/k7SfWL4hqroxAOAVvrNepeZFW75CcKs0uf99C5okQcEyr8z89Cd75LbA7f0fc
dOA3z31ffnUinDuXWgP68aZR6IE6gCqEy/Hh2IipvqcTvwMK90BJrfps5r3GvgnB
lLi0Oq4tUdgyks2TKr43c9bZCZOu4vM9xniggY9yawvAuDHZFFs5ITkwaIVBwOvj
5J3QZYK8W0cK6Q/0owEAwQgy+6o/nX4gokosipozVeG89DcUXjXMMdDRB23bOTi7
ObJlXyNkUBv+bEKQLItNPTzVQZfkmfQswGZvH81WR+j+FhCNHcTQrV0JOEG6LR6D
9xym1/ti+Z0gDL0pkqHb1gmxi/L6H4aYFC86/iJX4EhYkU/lAcPXzK107gu/9mZL
WWD1aKKWcskSehZNrnVZ7Uhmdy6PzAKacFpOLocxCeE9xopz3eP6AzWxbexfCW2v
9Wb/m7Tx92yKvqM7hfU3scU93Hh8Q4v2/Af+LJdoBLltEdLM0aXNbbtynBiUtA9D
if75oVS653Ssz+PggqxFkzv36JPyiuQhW7Pf9BQX0+y8XGKIn5CG6TYfD/62FIcK
hazqN6JwK/JcD0020SvFQoC28FAYP2HMWhsLsesxOycaNu8URMPvg0KZcHd6kA6W
euPaeK7uDTERb10OuWqgokw1LzKsNz75gTL3vI16+emAuscWTEH93aYNE05uIhrA
kHHDBGTs56c/6uemzVfY+N1gCBDZ7FHnDj3WOfIwXpvDvLhM6NnppEKfxzUNCl7H
MB8OqDcTsHKzVGDAiXVAH63rdFf6vMYEmj7DRAhjQ5PBE5bcJ86PeJdofib7zIhM
0U9vV0xRiJIyMAahqR9GBXPW/HPL5B0MFi5NsTmWBj9RrjJNXW7YfR0VUGiNqy/u
5KJG3Jp2unNamE49JS83TCjzZASqdlq+iXpEeJi0SNYvg2NL/y8FJYtZfwGFXGuF
iZ5ZC1P0zqhJdBCz+e3Mrm2TcKpBZgZwvjhuAfz/0CvztMMoYejt7UyXYW+WCeow
/2l4NgYM+OqNmzD9iEZ84mZ/iVS5GY9Q7sraw1NsBQmumtpbzAly5l42QdlkSrt9
A/phloul7z8ZGFVK9R34nYQDIOlAYXc5ySU6FrtUqmmaf2e7l9laUvbVCFkxxPda
IWM8Kb9iUw9KD56KkP19zdJEmAvXncOlg19n0Sk+7hFODiYYiHpY2f5FWYFqzqkx
iNBYNyZnm/N8hpfvcEPya1QWXc5/nVv9vCg4xfcv+qGngyn5QaNBchBFPMyFca66
6bcMUZkW9PK4XBo1Wwz/o+PqnkXUDb0pHhN4oi/Hy8vk2m6UzV7fHPjXAGF69wzC
RO2CEetREd7xX+uTWa6k9DA0aFk03a1RI3HFt+sGT/5R6hLHtaJsd+8BkUNgjAGr
kBvfh8NaUkoAbaQxNpTRLfh1uqSChFycsC9xxO6jmipMYm58C4gOPhkkfaUgqkid
Vkm/r5DV334LLC4TYFrUKemWk0A+fyuQSmTLJEsrCh66E6VgdHCGLcJ6lWWmh2MK
J1c8osyWyD2EMTDdHwCsCbtNnalCg1cVQgoMZZTBU/ouhS/x78/oI70K23nqzz+o
yCcPp5apZLf3JsUiVih3d4JcMNtvDgpvynVaQxpbCwe4OeE08NypcsSyRdkxh+HK
aoqBRqIEoUpL0TqDRbbIcejwFGizuJWZNzu+KnNO5MtW7+IzMShReP6mL98oHAbE
IuqohYZiHoD1GF7EfQrYW25CRS3RQqkJVo24+vYMbd3gF5gJiZ6ybmquvtDeFUIc
xa7/7CmV1Uu8TEBA+ejSu0fKvrHoOZvg1qlyrOetrB6/STS+28hAPIAMHUhd6GQr
SqpZcYlY5+0qTFwNkhdFxXykEf/XWJgPxVls0OK5fl8tczYgZX1gKZqFKNWMmWW8
fe7N907Vu8kniAXy1X6EdjVFM9wyHlppDlRJ84/SK3585g7Eo36rRhxuSDbJUYG/
o+MzHfUY+i7Vb13O1lQl1cbjNh+dXq1DdnioBSoWN/SOOOgCNmci0EAW2ePwDHIo
ONJv6Lwkpdm0pMcD+JkTeqM3xJVvUjX7cF9DRAFVD/cCjYA/Rbdyif5C2p/aGitw
mJ9CbC21qWIWEB4wXpjjOqML8TDsggSUytvdjoIV+MOPX0tNsc01btf2u6LeoMFg
2NkQSevExOEwJc32DUpOxOlMTjnwteORfuHkWXDhUzIyIm+qVaVb9KEZNBhOFpgo
oU0NLdMiveyNcVqAJDI16uMpq+bwrogpj12sEnLYMP/zEMr+78rLpeHiWMcHavnI
oFFyyPZug6NlxmFZbabaYAHuUmwlSPTuNXZtPmMyjfEPGqsvK/mLroyjfWeYtpf7
khxcPFK/HWDRGvlAPWbI8EpNzAUlrVUO/Z+IRQ2jvnoQk9CKoQ9MMyJJSvsoaddf
wmlcUozRbUSma6jYlzy1B6M2HNBxO2sSERARyfkkfdDYwp1V0k+un2T/2/WbnMMj
00yxLqzIWQUGfWIsBQ3Z5CTs0f2KB05o+L8dPMOLAKeHASJfDwVVxbLacW8W+eF3
Rw6HGCyJygVc7XByhgYJMBwLzJliKchZIChySgwi63tK1oIHv6OFHuJa7OigiL3P
bRM6iZ+L6Uwc2XTAXASFdfN2bPFrfYFNkhJKr3hnJKp22DMzvn8bTUogTSaZ2PKZ
lxNnfEK6VdbPlyUV1bbf7rySlODfazbRBebHhz95XieUHRxol9q+zjETfXjTs5Jl
luf6vKqJXx4WnjZTmrcDLcvKF4wNwUutHaWv2BrlkAYtwiYEnQka+maXTc4O9a8l
2zrq1KOqQuQjg9aEaUkJLifqoEHnIM9rAqiKBNirmkgWyHtCwPTBzs/sPQUxv0EY
TsdOqeUcfrNTi+kZQWeQN6yjz2KVUB1Povg0Sc5ongqRGzEcz9+OMO+8Raq5iOXR
hZncCUU6vleSfl8HREMcLCRgdaonlQffsi3/HxXycWjLzGLTmeqCbsh6ImvyOx1u
U8Q+30LZbKwsdC3x6ZLLNiKNK9PqnW32X7Wy/Qde/PUYFA/IXm3ISLSF7EtQM5Ov
/7PhavwyqE5lyPv+gU9tFw1+jtxBH/5F0dTeZBCURArtI1w6qkqRJYuQeBJVAtqt
OFqmuj7+AMLQ/GipmnYUiOWsux4qBXZmB0oh+Tw6xIc++TqE/91iGpbaW5CesVUc
k1BzJciPzgfUo+hAiQzJZlfvwNMdg/LZ0lFgtte5+NFjV8wy9u/99yBN0G3W3Aik
SzaZSZ/sU1VO9fV59R+k0Qj0b01e3FpdSR3Nxey1zCe+tcoUVzI6xY/yHU2v2CgU
2leHBXQ9WWiBHe4svvMzwYMhM8whsnGW6LqsNCMpV3463kgx7oHdWrb3QDBUPTW5
dVZ3V1DbmiHucqV9TVb6rSZ2wilIFHbeguJEeoBTKkCpdVLUocJlhc20BYsFLT/K
sYqc1M0vFsKMmkCQJ51O2vc6WA1wevSHwy367FizaRL934qAn9RoDItUx83rzZpI
90pYAXyDIf5fM8GqqrAotPrCC6b7T7G2rZbwrsTiINVeHVhQTvEbhbpmBiKorE01
/6KfSGQaVFgvSGPaHbuC1CUISFSRsQdQFUnL1k/uTKG7Xjmi46voy4f+kjWcYSKv
mz8TJwNDoh1v/j2CbsgwSg8yduHv8ssS2Ye3hEQq84eNzUNc2gVyV0jbjsON+zKu
gc/Mf56/LkJg09dfUEYuPERvIgq6QygXWysV4mUHGGLBMx/rtZ4lrPRmIGHMHbw7
Nwm4QdiuMKwJ+rzJLENW9ceBuyR9v+MISXdmmOynBI1aL2iGpxiFJPEoasXKBHLF
4FTjcHiHwCXgzTfjT9smrjwVX+fZHMuphg6bl0U6sx8NomPsl8ni3SUZzvd6t4og
01c+hQlHEhZfMaG4BxlyY+zbdiKh02JCXvsudoHHJMZtGABAs+5+anDIzHpRf1ZJ
5jWaRba4K+uEqOpN177gynT1hVdW3R+eY2fE8aSr1gcVXpEb7Ks5yTi3myI4syaA
VxgWhQFJOdT2c1Fb3DVo62sdgIEaXMi20g+WBqMNt+doAs8zn7cmjDpJ9azC88zz
f4i9byOtD7DtpFe/coUqNPOl8bE37KHIsiDOE/aQfbgYj4mv1uP002Ztm3PZKLr8
Fn2v9YCR7mCRHVNRx9iVYVpdXwrazWi5o6T/ZZD1uoMuHNZG/HWu1CNK9iH/VweC
d8pR5X1vccc04bctPhONfWr7PrNEL9gLFo4OwfRHmoE578AvFj2R8LvumRxpcb+L
UCGn60r6oBPW2LWd0XT7n/5dstErvlDSiT/zFKzLGlOUVOdmZqERGekZFdnkpJpl
UNNgEX/4IomRy0yKrPQigZHQpIKUq2z837sVDjl8zba4LkALSO8XuEJxKw8NO5P8
E/8MjXNqhCKn64+RDWSdufHEufpxPSqQ0eZ53QlhXxZ/+BpVjUUy6ddgQ5pb0XOG
5RVtRZcDqfdkI01kKdp0UD5kcuHkd/lp5g8bmqBOJWA0kMKwLTPdgxLNmYceaMZe
NRkVJ2LD/jmLKmLqkh8Jgt9WDZOmNiE+cxSKiSes5SwrEqlzAALMaHCXVXlF5lNB
jLDkgTCcUSeZ/gSV1cKOHYXxYZSZTW9zyPssR79nj9Eouz9y/0SZR6MDOvCqfstl
QPx4aiCzjSNCPxBnbwiDyrVQ8Eq7k9lXe4Jl0eYPRINXoleuWr3y079GEA0tEzss
GOJRV/UWFb9TkN5CqAwe4TYTTXz0vU/aYmST5tjNk37dZrMJof29RIw5ua7flbkt
AyPDqteaPtTKCjM28uGjZNGwhHUMRYfakMX+CburLAOnUxC4cJe8f6ds7YP+K3GV
DtjJW6zJytvQNwh1XEYvbfmoXQPJ+tdR/1khxzxT3OhbjhqvKFlV3WlREm3NGzc3
xcWTCWmFVnkbz7FjFmmPe+3AkAC5Rrk3Rx/XQ4ynkA3yTiCM56BA+P6RH+/yvq3i
smld+K4FC3l0uFC40Svxm/gBvN3kFw9htD5Cb1OfpEkqJj83Ui5uHi3h2Nnv/5/P
YRWaCGBPmEV8uf71MbRu6tW7Bw1JTssD04Qi/qPDrTJPSwgLSD3pLnHZO1LTW/D9
1PAmqHwiiLV10RmtySwD44QfHHUJWzzG6Xpk27/fEb6jIZYOVi1ptAoPNMrnDEki
SJRWhDzIsLjalvJZr2e3lTw9iGJNfs+lCDz7L7uq5tEZPnvK/GbA0xNsCz7jesJh
rcEyQNiRIF5vomHkD5btcCtATrXvFrCs4n7Z5FT/GiwVjcVBLxpi2N420wtgS1BA
vE1cIeTtfo6FSxck1ihTrka58RAWwCcMSCf+/M7gBtlTcLCDYj4DQ87hxU35FtDk
MKQyOrMeKDP/rLKTPAK4NobyFJUIC2q3j0YZon31fqGNJOD+eaLuMxWlZy5ea7UR
4VF8odVMEH5G3u1MVnrF4Q+4kpgf1+dEA+VLr5NRia8N4QlGCbDw5n8wt4ND2hDW
ccO5vNvhQFo+3XXvB3mvU7yrMMpa8v1Txb4IECWQJpk5J4JmpcWFocTBQkN8vs62
A7BbJEZ8uWAa5fIE2qo4wjRnTDQc31iGYzWvX91DPsBLE7dylRn3V5v+IhRBo36t
KOJyS1xV6h9hsvi8MiOsIFSD7v7v1ygukRP58nuJTtL51EPh35ikMMoeTMM73pmK
Zxw9tj/jWpOEUZ30Xa0AHIeTLdUzILvLbR3Q+DVqvqXdpqxQuc4WW1b4yBC63gcX
3HTIvID+GD1hr7NAqpOh65r4QsaNlrne5AdX9jcn+u8g3q0SPwBN2dwTq3vtMUwK
ecqPN1gE5uHI+Kz5KKZ9dqGRbCX6LlFdqhQAKHhLjpuEMjVkcNogRh2L/JCaE+IX
9JWUbScC8tey5sYVg4uwm0REAI7j8HkjtoznhONP09CEvChgmNmQajhsySUpMvdf
64sgqav5uIElctFtJkTOG+WGthJ2DSNK71HnL3eSL4wYgJ5mKJZYW2v+Y99Tr5n1
clkatizMH4wF3QcLaUA2vmWGAgZ3kW1pvjjoP6OrqF3sRy+X01CR6RGlV61as3tM
xTdau4Kr5GkS11CgyilTGD2XHSxnXhPb42P/oU4WfQjDM9zQQQrG5eh+rYvcuJ8V
x0d89j9rQL89Lin7dZOIe+G5Mvzgm6B+rbPp62PJqO8mc/p4S+5yrPKXJ6cjCh2c
bGoTv1xS7/wTAMfg79u8eDrJ391g0lmWhgi6IQqkYpQrkXRSNfI1obmbBGG6iT8l
1jnthRHm/NHCYXZYsobtmpfTOh0KBYvScJjZazXMYE43FCjOtDyaQUdkQy09zRmB
FWa/Ur5W6bUv+5xqMi1KJG++zILRIa8CHS2tRAHG8GTWWTWYQ1DLCb4W9Ftwq96m
ZVmUuoIEVUCBccBlnrlPbOiSWEkcNZb0B43Ar2FwPrsiJpZoRS1PAUoZO4htRWi2
K/cRptQvKmVsx1cXs3iLxtPRahCFom1FI89CnYIapd6TuQXlJwFV9HJ/901md//G
dXP8Nt82bPg0I/IT8H36Q1TzbT+LpUWB4DjxTNF+F6qaOg3TmKfOkGxGnvkCgSSZ
dMkZYiitzkC8XrJU1s+gOFZaKhtZUhkdPMDAo1tiqXqvJVeF56VURJz6cQnAp8CZ
iBn7HH9rfiN0gd6ELLhQJQVzy0VNUVb1Dx3xJP682SQFW26prk6ZUiB9OksOoJuC
jMmHzDBWx/ZFYe1KoqFS9rUMMH5wDXRZ85zzPtL/yiyo+ofWJY7abZ3BEUS6naW7
5xeUOwmChVXnEn+XYozHly2cSHqh6E8R0aL2dsgbP4AeuLEr+wQFtozK9ZHEVNe8
osEHBdNVrdKp3YJOP0gYz9LzCVdJFGYL2aqjWIAXIQnS8Ec0H5Lt3U0aXjVs/Q/q
Y13tLl7hznrrfppA6sRxrN7AblvN6YDUq53xYvt3i7CLibVWMHTEusYi0Vf/xM7K
aEKRTV4DFDOpUMVT9ZbFaeLurwvPF2zlsw+g/Zgon++t+rkvaO6R+6oGixMn+HxL
Syr97fZSW/jgAsTjAWreMW4eWhLCGUP/2G6gJnDIs0N1oAkpxLJCZ9PS/LwBW3uz
4GjaOqL1Sr+FvdQ7uJgiEyiybeHB5sGwcxWDMzK4cAJGVPBVqM673Dn2+u2CGc2d
0aw+Ad+C9TDvGaaFWFEx1l24QffVZ5vbJ7rf/H3KoC3t6ZhiqUaB/hMnu14H+j3B
qVARE0cSyWzHvakPUXc8/7D3X/xAfJ+zl5njDNfOzYiGM0/v5zV6mVEk6OlSwczg
NUf6dzozGne9iHlO2DDPF0wjpY1FtecjD9lLuLfERYgUhnLNJa736rLv9NbWYDIe
HkNC7KMk0NVfAxBXCT/bJG/JWzLqBFdNr2B6eG4bbMscCnF1PlO3RAEuntDltPIz
WrAjAqqIil48QWDh5chg2uQi6fgEj3IVfI3bbAK8S6HF2EuY52Y3giIcJ41k+RkY
+m4zjEAurxanixlrXaS+wuaPI419f0LuoqgcQKycOEks3S9ModbbSitdOOfuKPCx
iYH7EGNzcGwIEyV4GeYc14LC5Ja1+TjYumJawh9UYgbKRBrv9xczFtooal2G8Q8v
CUZPlbfZ3SKzyb/Efr+AbuOARudgpu6vvjmG6jijX6jsad9WN5qrezx2pREyUIeO
qSN21ouMoeKuHVrOO6R9ypmWrqRWffiaIrhCBhp+VbA1ZIardkJlbGwnBzZC/hkL
JV3p0TiCH3ZGgOa6llVvuPQnCqTvclTD059JFXlkm1a12mbLYMCG6rTjb7MnSPnf
YBH9t+Gh69kh/ouiERLdL+M4bPAbPtM8io48aa5z1k6aHnVdvSj510DEdzPFTlEO
lhsnrsF83xuCLpMa/BZiII818x4t9eeyPpqUKbRpgMddMEtunNWC2zqSP7BtZxLA
QUq6rZ6JMtBQV6ONnZQ8CSbxtZH/PkwAgenX+lNyfV95Lt0ems8m4mHCmHFUpA6B
o/6fNxUN+AUG4Ymep2PjCr1pUQ0LuSiXnz2XXu0QfT7GzssDD+R/d59H3NX1uibI
ZgdgPISfe66MdO2Jmg/+VP1H/pwGEZPeEtGnmdl8ZYMY9EQW9gqeoVIlvA4k43Mi
Lk6aGwWLgFYpwC82J1oJP6I8dRBLjuDuglicotFtxwwnAA2IC0yY10whFm2BJ3GF
c+p5L6xJCnpXrHgjo1yAUlnm9iWrS0Fwajd+qPeihI8TleetKUzvc9UyrDbMVER0
+7/QaQGBEVzYb1eNXSjYwqS9NmaFStmoiXY4WJQInZH1i9nrevnScDgBsfX+aQ43
nCttQ+4/e8pav5sUtHfPfNLees9X+bKfIctHgEI6jCcheC68kpWjMK9bZLIXWxW4
r6ff5ZypDckyc2Lz+rI/d1IqlBHrdsFGXsGzm5hvSrl6tL1ZSHAoLQzfCwWR5iTz
HG9Q98IR5nMRWwcBFZc1E4a0c7CIP7StH1wNZxkqFvgvYprJkxaR6uco31Kl/Yzz
tbF8irRONWh8IHRObogV1LSTMSljYqgVmkWMmAtLCNNp6UDhrIG70JnXCsKZ4xl2
6ndyhIqQH7nBMIV6oLm3trK66ECpzPNbRKS2av8QD1iASzSHND0vDMi42Thqz7k0
bR9xEogSVY8Wjxgvxp21qeqS3hw85/jMvqM6lClhLq6JAgebqygFNuzNfWWIJet5
bMuWzyq95SqvF3yrlSyvdOONT/aQC9vQ5w1hmHi+e4MSq3jNGhZChQKC/eD40KsC
UJv32XmPt9DllPtERJAfkzYtmbXloPAwtLXpDCHxxWhvlcTZznUESFygDZWAW9sR
AZRSLO2fvlnJxtsI3AQ9ueM0Ikd+Z0zzJQfBhNy6bcfr9JVXc9T8CBsdDjtpO++w
oGAkK0MEw7hCq+zdtTb6gysPeycuwgHyPm07CQud0hPzUK1bKsPEqW5QWl7RYsT/
Tm9gJl18XKugdlViiKby/vaiF5jSipIljbm9gXTcvJL+d+PplfVyrKoXNvZ5NSVS
yA7TpRT9pzBH0++5Tz15hWW30sLW/0YpQgqJO2BblEn43HF4XNeEpp52Huf3tVAf
F+aupypaSOp4qBP4vTREYrnsCziqBvoUGkGTZhgpP2VzRfn35H483LWuVaZ87OUL
CAB4OMMnkrm3OSKKjZaOXpqyGhuJ/yTk5+gtovGhBqwR63Yr6+qEGFpDXapioGK8
5vz8ePu5/pWRslSelqWVrrySxFQRIWAOSxl8+v71ijqWfTI6j3cUghDX2PrzpES1
j6y8VfJYEMbnt4EgPsy+vNXM0t8A4yN2cbkII0RqY/A0/+ou35ONG6y+g2+GNxl6
py8SQSaq1DFNfVXys52K21/Ek5ev9g8RIwqAU33CZo7INlHsVsoSTAYacIB2Z6Se
DoLDz1LyRlLcWMm3nK6CJcmvhGVAd9JOtQ1V4vxn0KWSa6WKWJQdHG/mqngJqbVQ
IFrQ33UUaL2BbBy59T1pllYgu78ZA+5ko7LrgOXlnZmjeVWidAlw2NU8nfXyhXpw
EUm+M5Bldu9Hcr5MP3iZeYFrUqCrVOrcRuSjobxNnZda/2p0Jrw7bdklSYpjWcMY
1Wkp74bGCQnvDB7yjaycOerh6MmWhg0HsmJZv5Ga8JL4XEZY+C9IpYCiz6j0oGH4
BqNLHCBNf+X02rRBF35Ikw/Oy5oovFR6B7YSC3SZmPHay1Flk8nUWtP9BqSytWQE
009bjdz+zNFJ/py2rRG05xeOLMoH21de+LweZ8a8sIP548QOEFuLQXLMvncZzCCY
yRLyoWC9dW/gtmnOTZltVITBA8/jynd/MrGh0gJHorq9nrY+jI1tzGNm+DNRyxPf
rN7FLOVPFUaqCgcH0kDx2eyww5unwcvdDdEVOficVRcNimetd4ikr7fjLhqrXFZ8
N+bhPFR7i+npUbLTu72tuW6/YPHo9wROoxZ3XhRykI388QSVEiEuIJksC5cyvK9n
03kpTfSl3e8zmh+kcz/pi/fH65dKjPK5lzSb6kgH+Cm4jBmxr7e3d1CMj4gDKx8A
0jrvLnOBmnCEMb+MPVrdmEkT8PXMmMVi57hD0uxrbmA268P6iL8WbguC5W6G+4Sc
7hZmKx7R73a0/UGo9wCCLvUSDMrlQssdWCMucLt2USZOWEZrV4o+z5/oC2pdKVMr
Iyr+dEnOUDxM0mPnywIf+rb2n7nzP7E2T8FsX3bj87qtQYoWhe1tYy7IugQgT8fI
T0QhbUfXa7y5dTv4U+MJRrUyi71AwSQdUjSyLnifdlHS7UmBf1oIqiN0iuA1qONr
/MtLd+zSa3jK3jOZAVW86hm5AwERwmPm8hluaYqTaenyUXQeBy+EL/dj2Tbnk42n
USUqObnGjTnSd7dqK0ADJfPWL3lOLVtF/uLEc+6sZ54ijsouga/wefRAcPT2VcpN
k3CUHhNcye9SV1U+fO+DvxdBQ6faWZoPT+syrNullf9HNqc/X5Y1dsY6eW7xDzKG
uXozhNm5CUioKNf0ujsNn1PsMAFBCT9ApICpIrQIklmYgt9nsmiKgMaDo2EaC/Sq
Y3wL7F1pSnDl4m487lwj5h6JqzntrQVNZpmtnG9PHbBckC01W3qnR1ldOFS0ccY9
aso4EiF91qnx95sRhm6tQyaAdWPCJ6tRowhxJ2avMAA0xzg5MQ7PATd3sax/9vHI
jBPVpr0pNDFJACXmHpDHWbto7/v60l3tRRSAjE4tmN3eY6CyKZ+UBTxBvchHoNo1
U3gcmkwvvE6BGQwkNGelVRStcQT8RYJyd8CjG55VpYQyOleyR6XDghvmRN1z4dzA
2/1/NZcnxsSDSYuD0MgZ+SLLXmNB3WGu2OjmlGOCdi3JQ4FoC4ceFDK3HpII8pSF
wHHwi3lryQ0eQeeDFjXY1euL5vlDsIjqCBnqMjLpqDdjPkljrSFXi3x2x+mqBf9f
MBJlajEFLfrJbxAEIua/Yl2G/VuCAq6M5rjQU9/X3fWjHP0NAU74S8W968w1Lo1c
QIYcXnQhCkp9jxvwfTlpvYjHkhjgwPU2zemhRejVCkL39dZGzQ4vmsj9pkx37x50
HfIURPrhnf6YXn0XbRCRfL1iMa7JhB9EBCdvoIcqMiYgetaTuvVrID6a38zAJ6ST
NY2lf+uAbqWJB0udQpXaYpGdMBe9Kli1KJC5wKf9EMLHuiuDIQLLvztTXT2s6VRQ
0sHbVkdu3YS7aurBZHFZrJNRONrj1BPiuHIxtrzh7310/6Rjm14EO9+s/HdVr7sH
zpzY2lNkJuFxmqAv01GmaGkVfXAzPzXtPdUdf9a8u0uHtJLee6wclddW/Czdsen+
+24Kh+bE0Km2xkzulWOWX6jVd+ikVOe7IOS9pNdV0C26gRxlnRSW5BJCK4RwTcoI
fIqPyrpAfJZhnU8gbSLFdedB4IJO817n79ZfVuzQypp4YEI9KowisgbIU1mKNsm4
8EUTLVyVfbqdGRln90qiPkfDxsrhRUAB3EKy7M8+6vCu7j0I0/rJRWCoPnKzxylj
XIZ6r4i5h5ywc8HlKxX3oOQHbh1E4Kgyj2i5yqUhQUjG4Y81Z0Fo7UQ+NWqV8amK
zNFHNU3w6/9A6cpc4fdN5BxBFWhxHdfcmVOG1jSnKqooB83ydg6mongp9tD4RMEQ
a6Nn4KVedDoVWU5AUD9+4QVavOL8QUogLeZJHev/bmcUJ2e6Hl5eWbq2bPgLSTig
LNx3DNrlrI+H34j7E3LyBjwAQrDUU326gaLbwwUGmEzFCh1PMPXz0J/OE/W1zRSb
C656IPi6XYutsLCfH5Llv0WRoZYJQy+txo/vC6CVnEckSU9GPupQux7pidkUn2D5
leLSzqbzF6OtNQhTlKptJcMFPX5eNBVaRWWu/+A5rShHcWfwteOXRlKTUX0d+Gb0
tGv7LkH6nBW569PjiSXxGKaR5P/MVzbo/HW9s0b1iUpyBuTHRD5LRcE0egGmrXS7
G1TkLeiHYmWExABDNPoUzPP0TFGORRhls4LN0og4rBKe6UZs+Vm5HbjLbjvuwhx7
vdFvA2IOxPkE8DKHkFhu11JRRMJBuPo+IT53p9UQe27Vu47SZf+wIC1acHpkwMnb
DqcUNDtHh+j/TI0LLYnmHm6q6z6B2sIjODyDq4K0OWKXe3G1aJRQZaDPuximojOR
i3Yl9irW3+01CNOcH20v3z3e5M+ydhfRrVgccL71wnVunRq8w7DQUg0K4HxhtqA8
uKbnyTjTTN7J1Q4EbWPwM3auT97GM81NuJmRP1uVTAlxZNVasktGY9PJc7FeIPu7
3k9bEzXefV2SYMktpynS726W3FPt7yzhvNx52YEm6Weh5faHgGtb9NXBCCqkDPO2
MvDwld8cwdaAi8V7VW3CM2XhbqhmB56nVJ9IKPkHz1mcPVO0v7itojy8hqTFhZb1
2z4B74Iu5aCKD+YCM/KC7EnDLogBGPJcAxBSLRf9bSv/RPDGG4Bm3daK6/kU12eK
X2xz4JxsKC17e6Z8IhxBandL7aQFbIhg6zYEogp8jnE32OQWCSAx6jHCzVXz2/Gd
8+bsIaSQgC/JUTRyHztGXwM2XYGdzktFOH02d3F5hgYUP59qo2k9cyOazXN4xVEa
9sYzagCElV9J88tEvNUffQHa7YK5B5BdFV/xrjO7Aylk+ExnINlF55CopAKlURnM
1flaS22TYFz+bNvkHqEgzj0LCKLEXOMaF+8VfLnU0vY+tH9HhPx99zVyIXT1iQZY
hg4CJuOZIv5zas7mNAaPoN8oqLaBCpk8Ut4aFYGJZ6WkSUi7wL4me5EYvmlfjBgW
Lpmop/pSrvaM2nq8oAGWXPSQeDt9eOZo9jUWPJGmPk4pXrhwm0ousvjf6incSAXJ
UmpU9vwZPAsZHiUyZKJBKJ39wqM56HiMxkBLMdl0xfhREcFsiWtA60eGmHCfBOlH
R4RmPBhQenh97xdUwc4Yp2VBiTCphgUyC0KzTMuTJ2f4Cme4eFaBaMCUdjqTE4vI
zo4dwGFUldQ+MlU3TN9zfw1XSSpuWShYxQgrXhS8WqIdqUM7wPM2CpVR9w2Wh58R
u5ZSL3OaAaDpKUw3a7dY64hMfIerL531sLvTeGmUW7rSZNDLNr0d2Rsbel1ejo30
BzgIP2Lm5pzQokrt8AwkU+PL1XSyWr7yVCkpmNbakxHDB9vTMW3kyG78+VA0yH9j
6l/FHRGuCmE1/LWZa6x+/BpWTDfEZCpSW34SeBwZWFQ0IfjENiTGwgbxEXloEtS+
YT5Q/M7DaufZnEsldwqD+ipKCGqXOooUZo+l2Drauin0GZge/LagFvU+86wrBAD2
iNzMiZnZg8RtPcUjWpr/cwWrexnqj8I1VFmmbuMZvAySTHwXpdWg3C4VTxh+q70E
YFUtZG1+iK3tYVS2VheLJ7j3CMBIxsFcgXnumYKSvWrr5JXgp0j7z67lxxKy/LAf
rSd7Lum2SuV7wZutA5vXLMg9RsblNqzXnzgtHSZhwKgTMNYtiryRNZGdblAuPq++
XTsxkdqWHhKizkAvcqklTkxLoSIGUs5YQ/G4UbFXvPI669hHJthiC2y/WumuGV/2
77P5Sce5aOx5E3qeXz4bv5xnJvR7qqQaWz/ESWS7w5tJFA/h0GE2rr9Y+un05s4h
bbmXXBUOGFr1suv3vvVBHzREK7z0+BMSklL7WA3cCYjPskId0OkbwJWYLAIsHiqR
iZGE2L6DfRgPGF9XZLGD6PmoNXXzuRbRIV3SCBXcsxA1wlgxNfqwhvCRbxOU0bY1
IYmxSQnp2qvuX4s0zUDteRTB1wovOAuCr96nvK2ZcRYO+0kyeF1gBBPLp+qG+XhY
YHBZx2msi71HL6swZAofaLMOqo74py+xbcQPucTt8Exxf0JT22SJc+LcZt4GjWDS
QsehsLT/TG4Gj617wLsujO9gSO1wki1aqmsESr7Xa587dhmHLAhDKYC+1rCSuWAN
Mtl5H4KVCDNkp2y2gIWythR2XRbzxiefQlQlhJsnWGv0dCT7D7vVoXNUn/gSrmzG
3CiDYVxdtn3eNCEP2NXqtCxLDHzfbk7FgW0qHZLLdesUMMnMpOjRQd+Uefd4Kl2U
CgSmafNKZ7al0Dr3N2vGsytqsZVbX4uzbo/iuYW/nXrRZQj8K/JkwReitfwiVvBO
rugRwuN1hx2EozlmPvuOy1PQIX2aRHu/MIPaVJ60IR4mqtElERhj/3Y7ofx7QLE6
oKcTdrsH4jrWsGK+W8jpkJH05hMdeOnXe6hz3vdYs2x2WnvXYoeTulbOffDAlGtL
fjf4hAsgzlzrpu3PPmgqeA8NRRE4T7UFJE+nYwSZ6LyD9xRfLRyLDDmmMCRu0J8w
y2bTjjX45U5eBocDZC87cFZHii5ce0uRU90S/WB+HCv5iOEPNALNLRFC9oVAnkVa
5puRhLN6GmclSzpE7tHgWoao0e1gnTigLxm2EcxpRDOTjFLJmL6Uybh93rkv8zBQ
rTuIjR4xXacAAnocVz5jlYBfBujYAKM+xEok22xXV5peoREZfRWKxa+yjLtCYg9Z
8cBKtXvmfKomjc9rVHuQw83igencSXo3m1Ua447779UqXZW6hvyIUITIstIxFGFF
R+nUefY6d2tOhKC9q7r01R40hkIY1uPQpXWYbS31Rhz8JwOaPFxJIgYpVIo8DXtP
UBNDlUDgZye43AaiBh9Dg7znzgwvMOLsxOg+AH8bjvCDwlCV1iyOB1TiowWBP57V
OiwrzyRutWPVgcyHk1yX+FqgC2tewrxO19GuqUWLrVLbElWLGQXvb7RuoZpUih2i
DSl6wbBrKRF4EVGuwIVzrU+iasl/fAa+KT8k1EVm/KMh6c9sFuQkyifhvC9C1d+r
aGJ8c6UzugFZJKmPwOB0HnbBBR8SUh3IUeszKkriyzXrS94SiZv7nGLuCkVW7LzV
CRG7MLtS2nZZWYfHahfI+s7zpW/UcNw5B36LEE+quPK7idNNAqwDi3uviO/yNYJp
xFM6CBf0c15AnZdJomOLrgQLJpaFmnj2vMfvbLL65frmrzmlkYWJiEVuTt5/peKi
ku8CFFJ7SJiM5b09+OqAhyhSQMl1ikglOurv6lCXmWHRK26o7O4sW8CDprn/PLeD
425twEM6HNFWI4CBqMLYUOu4IE5RLciG25qkawCnxjLJG9cmz0hdhe4rmTY6exsI
27FbbG3kYeC0LOi/0Nycjnltu2MKWhESxPFnH1pN2fODlcUvSjZhWxBMuwA3l5yz
PK7Q/TlKPAUMGPyXBtrkpzT9DPkqmoUqFhnAPZjML+HTqvFDutEtdtYU7wxGI02s
2ntvJqU3Ncyd3Q1rsX/ZfJD0h+4WbD4MPrXW1u/xvG+C8Gmej3gt5DPUxZLaiUqq
xCx4+Y9Zx/VAnyjrVLywOchGvLag2a4AdazqpLIwAQPm/YDBHJ1XlUkCUfdlPDcY
ijcfWk6rBIRg+3Pq1H5FBnep8dt/8Mfyt+8s8IXyqId8CH4m+xPi1mqJMa7rGgX1
gSJFM4OaF5rYxqH72AFT9E8Gv9xb2BI2kbY3ry0OsL1LZMOPUF5vdlJBXnVzsZhB
hP57OJThpD4M5jxJ89q6vujclNMa3eHEW2S0iL+0QpkmxSQ8IoHb45ZmZT6FcjUz
N2mBl6eo8UDTabZEXOop46IKnCr2mxQUNOCa/k0bP/SR+RyEd5/UHdwPgLlGXkIO
vwrD5vlzLVW0tDoC4+7kxE9u+8hhfY/gHCtlFya6wzS4MM6xvPRVpUm/fqIZaqAP
rRPs+SgSm3BaViNqBprA8sykCxL6zKnf8rKB0mm7+LEj6lsIGf/E8QqREsT3C999
25T2dCUVDPQn6gRcfOwrqwCQViYhpTC0Xlc+1wYmHPh2E0fWhdqbQgV3IxyWgB8l
k+PTcjntOU6u99hRHOqGR37FeGXiurbaZIactb217qcTQwSPjZ0qmXHWZMtzekYr
gtP0PRmcNP6gMs1Erc5OU2rmCzLtdHMfW4BzoBU5Lc5P6jAlJvtFRBXbfMZgfRfO
1TX7o5+gnEJUCFLVgT3UEe9L/g4srgcmZj/XE2h+b745veJMGAgKNDKFeBYK9t06
xf4OiwERSBtcT566mTA+b3I8OTxCrtmLnFoquhY42UsmooihD1f/xPHWPyDAXQAF
OAH7/rmI+4sceQUc5G0JtSFIQ6odc9duuRcR9CofpmB/sl7/6ZDnVv02MEaoG/V0
pqT6yU+/rwX5MviZodfkJfunRgeIrJm9J2Ayf8yPjwqM+UVq+TobXeonRbH8BQpP
fm4dg+yUtCpgsE8jbrwbQKtgGi5s/KTk+W8H0pTkqgm/u7nBLfJSQLYmyFeaApDZ
AHgmPCsT0zuEWA0wQai3AorjRddMkY86BNyJD2Dip76ectQ122EVK34MtFvhNRHZ
lwlwdgkDme4whKioyzrJsA8a3x2wUJbBV7UpqXAG1AXk7nzFINB095X184uhxe6F
qObygGhyPLBDU9/L0UpyzNomQTqh1gv8mg63s3PYLJbYiDYEJ7ZIxhVAZ988G/xJ
xmcx5EG2sVv/DafH2zrDZ8JPqQpxjNTc7STUsCDv+mhLWGNZE1SQUpAYFPIPYvPV
U5ynGzvg51OCCsrGNl0ma3x7R3L8lgru3K1EDa3g71PxcKwXTGZyfir5/yvaxI1t
kyuCD4+LLBuOHsohcXssEdoA2wWi3L3lPnkQu+hUPmbUr/c7xuC/CMkbyG4wQh82
U6jxxmvQjewEkTleP3ZEj6dxGzGyre88sxyqG+G8Hktwn4TFjt4fjgK2J9JZpopN
mJEydxyvxgvN9/oK29MPKrre9XcrSG8B2yDoRt2GAEiwvqZYn7ERpHuN9RgMOBqQ
l/FNikOM6VlDz4B+M645pD7LH6G1apLV9V6h2nm6fRO/NYfTUUrLduAB+biHDHI0
VhO+9ZJvn1x12NR7YLIR5yQ9zvkK4aSRNjFF7abgp7gNMevCuv0I2O5gP682Mnwa
iqHTvepQbBv3XzoJm01T6sgupWWFWyrx16BTHiF4LjnYd+IE6r/NA/WILtlnRiPD
64hRjJ0jYNBZ4k2hD9AOscIpAwqcpbwTa4sJ7w32TWtS0LlJ4OO3Vcp9Jw+EzDaq
4LDa/mkxDmO8d4UPBjDm6m4LtHpn/juaUtBxXv5i8L/lOvhx4bIN9Alg6it8XFKf
P1DNpgBXc3j9R3UFq+3BNWeYRr/CTlm1fbQ5f+R440Dp3RsuC0cPMQf5mynitU43
yEyOs/NTCs3b3lduHZi8oRhRab3e31Y75pUbYFaNV9ivbVDLrRKNX6THFHwAC8h5
tXIah5Mwxr5pSNGsZGMMvp4sXAN38W8PKSQfdMzWzF/G9ip22rmxKA+RBUwtgQ2t
toHZonXZypT5qdSnnfFnAfu+LKPbQ8Z+STatPV3SY5FlgPp/3rINbis0a9o5trcS
KHGliwoxYvNvWBhendMaHR+vPrwzwypcnQ5fCb9PMzTf4sOPM/yYfeo9nVfJA4zH
sPisaBopOBp7IGOrHGA5D+cS42UGaId4ARK1BQO0EjxeaO/TEhEA9MOYd0eb53Zx
IauIvZIh3f5HJ/KTt4ZrCgTOpzzVoUJU8oqcshN7QoYm8xTGwsJz5xmxJ8tU8omr
zJBf9ItNGf60MbsHBvagiD5BNJUS17dvTwSO/vuBM34Z08o/pFuPlTvsfWeYAPqZ
WgfLSzyxXXZJGmgkW/S5peKrMMfPTy6ybjL8rhhRttNGo4wqOZD7Zx/msWKZ0yg8
aP1t3qfYCsWpzFmXXjC5NI3xFraziCjqN4NqjZvs2XViy8M7iLo6Uz/qKpsSpRSl
kXGO4WJsLWseHo3PqUsytKCe8VoxtPhHZimdPgwkbpq1r+PjLzW86feJN2l6/at4
G1YqQxJjSTGUxHMawzjBmaejLwZ3xIPL/fY9mpR0/hhppCLTwjYzB8Gr+75+Nr0W
IKhS0kBBhPnWnAI3N7x91P5d0D5rIOuXx6ZQVscjsSqw/Gt5COhOdgkQjeWMqMZg
qOg+1SX03WxMj4gGJzFjnCflToztiLJZSwEWTL7UB13tXJ7UXf/vD13mBIHTvKEm
poIWgwQ0I2vKMzxKKb92trCSXywwhH3UpR7OgkXsKeLYOocQF1/9IXrfF9DKQ431
EatPxFLD8y8+Cjow3pxz7XNNfkMwmQDT8yhHdravfkhQ1Qfn2zSaQGCSH+Z7tpI1
/5iUj8bsj+trOha7dLUTjYjEsbwjZH6NizTSXu8osC1nhIEmKmaug97YQd7wmgiO
ZRtuq+6WJJcO7L2quyJUU1OEVOYYm6o2Wi/VprFG6aX1ZV8ipWjegyqHfDeDFuIx
Ukc1hPAoP9TWIzhp2FqE5/W8gItqtOXj05WSHtXwQKI3XmmTD7eDKAqUtgjx7JeA
LOLyLB+eSDmiuO/EQE1Sg6lxs46K6mdpcOB61YyzSVUQzJEqAnWfdUanyeZt+6Dx
JBspUbzPPPEt/c9u/3RaNVGKbG8xNiMvy8FIyxioJGhyJ0wiTu/hjmPo9nISm9kg
j1xKpKmFT/X4EEMpgzoXn9ZZVuWNkedcW9w9yuvWzTUD/H1myc8sKHw9szGRzRo4
x8OVjWPPaPFMndqYHHMM/jy5k7R/qNVsOdHpbtV652BeQ+Vs++7WB2BHyzsFIx8s
nrDqAdVP96rYAEUYejIhgORiCQqHR65m7JjBtIk9IlGc8WoFo4mIVV/gzr2CsHDO
QyZuUJK8sDevJxFXjCE3ZIzkxer4mmU2PL8RAetLKR682vV35LhyOkm2jYvZbXQH
LEeXdYwZRzlp4EIiiSLL9r4Cmgg5NWWrF1glMXDYfEoMavUcI+y7MNgUfnAOoq2+
yxSgNYV4frixDT6uc+LCeeKPFKH+Djg2syjOonBo4o94rPZEdTzJ/qelGrNz+4mx
9J+L/TBQ1ukvhl/xIwV/cnPadsx/N+Adi8higgQTcrgZzujPOYIXQbW/lbop/OGK
4eHy/NFsVj0LivHW8bQ2CMBb/RESGCeMH6yPgm9AB/LMRwVI1YA28sIOBLf6ilMx
Hu/UM3uDSS0Qq6dycKIQKWS3LHS2mRqYO/7/Fz3q8JgLMiRfgWCqBPKYsAy3UVhU
DLura/MmGaMehukoSh9vVTdvhhwUTr81OI/qvssw1o/uS4NseoNordf+moidVhba
vccTfmtCbxTI/L4bn0wTRII/m0VzFnd3Yckj48qqKLHPwub1roTIctCXEnRfGx4F
2ckEHQ0Ef05zvhXIdR95ayMZEfR26V72JcqNARfc/+CN6F3JfFagLifrUX//9j16
LeS/9M7wxZQ2IeOpJmWo10pqtEBrEQbrzYVv6TeH85H5KD4yqNEMJhRLlURGPeDG
hwugPzZEFkBptTVdqCwah+VmH3ygYyedJEzTo+Iesp3qDnU5Zh5wTaI3HLzlAfT8
7qn8Q8mQ4GvrOpnQf5xNsSZMaychFd8lWoC+Nv0VZx0O4eTaxQISuUpnaQ7Jft/c
CMDVmOlyn5K3KZBqs+AubYf6SPyA8lfXpHsiKRnmP3jzuO65qjLLTYE2iutiqZvB
o10905A+3ubFglifAOuQomF1G9kg48ycsvaMf5jGc8U3iBGCuaSxCTZmF2kw6Z3O
XakzFfM4esyjRvPw5HQLewiFaSqPF2XqKIvctJMGm8VQCo5tcSiH0sufpyOq5QUZ
2L6wy1GLqnfqNkhQm6grJ2uyeuK3evn/BF21VBDIiVXZnhCMobcQM3JxbEkQm6Zb
DcPFlHdzhBKCAP08HFU/fszFK70SbJ3Ijf6XNIw6p7N/wU8Nc/DLMCDD3+xDLvPj
z4B1FR2CixvJQtgroxu4TK7ngmg4d2r9JqtAq3NZs1gO3vbAggfbWeOMEz0CO4pQ
Ryb6zT+O5xA7zQJ1ybldSMTOnZevh3yLAp8IE6OkHeLEX2RBEa8fGJhcQGaH2xoV
9TsdUUybqwj+A829FvTE0sIopPQiPfvAa2eWhzq0OZbJ1vby0/rhNxkMByiIu51+
pHO0znmAW38neLaGuUr1/VD02ocnJF7EbKKopIAwFTLDRa8hRuxT7J5Z8abnN5xC
EJuqf6kGWjz/B2NV0+eczM7CWTm6jxRjfj2Sny3I8YOcZtqXwVIInKQUO+ZV/Y14
bU1w6IikgSEsrU16g0Hq2N5Jk2yzMC0Tty0yFkOCqNolp0PRg62iyzIOn2KKY2te
VFnlDO7Rhhsx/cezVwTYxapJMRC8fbWwliE0iqwkp981tG4/GE/lINYRlnbaWvlb
+2b8itP6WYBY0Wld6r9gDrBUsdKjZ3B0zb9TEgK5/jBFTiNTYciS8hTTqUXrYzFK
82+Tz3kEAuzZcbNTX6rwGljuYusAaG5cFfMYtDkYaQ5Ka/2FHwUY7cNz2wezUU05
5/HJ+tWfU/O/FwGofSNyby1J/Ruyv4Px1P4TxQjY4K+/cTaXVwGQP1b8StHJpNFG
hXHgKJipxD4ASmRqPNPPyMAfsV+EljG+/WnDXcOya9AxQRQrDgOx/7bPdaAFHlBO
H/d1rlGm6DFBIjclW97O0NweQ62CEYzZU2OyExb9aGf9+Lgz309ahaFayYk9HN/4
n3i4g7oHJg5OMVeTNOfN+6vEc2gBqKqHQEakW/9baybapVsPHEqbL1wldhQXvLb+
Rk0fUfAa0twjQUD28IKa+gZHz0+hRt1u62PMawcBa24u6ebJOnUx01k9PFJg/HgW
+jj5AARHgtFPlmFdg6WkDQOOKcWXgaBxYUd8cFERQqdkNyZ1k+3JozMI3K+43mDY
pFGd6iC2c/R4ux1x2kQ19ozaG9PoKpgUrb9u/g8v/pXn08zjMca9aEYaKmOWbSPI
7HKYPQZ5PFEhW4MLg7ENBoKFySc6e+Y6AWW7uvK4u1CJs8d02B6ynfl1JD4zB+An
bsDch1OxQmzHH3ceYWw3oS8fDVhyHPCjb5khTHXl357CWKiIpiGXAp8LUtTwDP9A
b8734gvcv/Uy7XqetS81bzbG9KqPZpo0tZCETYgw0ADZHfNqLCk40rGH3KgqXt5N
XYr6m++0x4SwN0txVqHElU71rlVQf96/48crg/YDRNGLF4wrg5OuCl/Yl7RSmDAR
gqtUHakF/8cH7A2Odivl1Ci5cZi6Ubunnk1OOMcC3JQf0GxTC+U7uyYg2JSqLDsS
aL9WoyVTNypjum+qO0SHHqPxomW5YjA4bs3Wfo3lCdyuF1XTIdtAD5bCdGIxiBQx
UPVUBvFp3ArhjNsBwTGLwaXzaHTw3h8VtS55NGNNARc+Mu5tJ53aov8KSHZHgahx
F3vA5zU+evc28de44kfGoKNdjdsM5/VHbtKwEOnYC/L/7jHcg2/2ccAeJWL0AePL
zk2AwG7de63/oNaMtN47PegBRI44p483jzQKZxorQagl5cjnORsXcQDGlD1THHlG
MRs7dXlxrplCBlk0Tz7PYkMoznkgwhudJP5NYAMIH7i4Bf1GnWvuzE8Hi0p5TOeF
yldxNPlxSXqAGNswzSUuDljM5/xGT3wRbS5VGS8RiMsCLcZ21NwsBZ/ohGMSyA1B
WOGjccc1sdd5ctV/1qQUes87Pih+JAKe/tYru7HdvXRiWX+Rps54fGKoM/wnON5j
JrJyesdntdRTJLIrGBv7JqJwh+isQV+97+R0nLwSnb1yZDpJagd3HgHbeYntnlAg
jP+eKd8/Pzg1cfMZTtj2OrE+nbbVgWf088pBCMFx8IFT5dyTwvJDTNwptpoO9fMr
Z7Q5sE1+FdAOo55hmqCi1FEk4pLhSf4wvLwKXmedPxDRrKVTc+qrT6kp1n1iQxri
P+/ZAhEKiBKYZfmuyrbnUyC1VV95vSGh180Wa83p0fExNo8wT8J/5ILcgiRQHX2y
pqkfSeLGZ4ZeJGPacJV0xC51RSKqIecANrCxszJIwwEquSO+by/Fdn5GMixnzQWx
ow4KZ9plBhB/9ld9fwxo7EVXVAsQXU63jp+xWwyeQ5PUH3GoFw0tXwbp3FeVYk64
JqX7vHtyLREJ8t5JpEYmtLByGfZkx97SDgRF/lkqxRWjlCB6is0xvBvawWFRP8+3
3o2DlznXxWVdyWwg/9lWK4r4LPvxev1VS9HAGVRIs4SyKuZ0uQFuuHGrkL5arl1b
SSxyifSWeyWuLBYWLxBu7SCNIOfZWVuUQkRhnAqTRdQLsdXOU8X4n/hvJzz1DS/a
xpMLTD0VxMNFrl0FdfUTGpmVVXHUyO6KlpBWKotEnhglzGcBOo3HFzVaFNFUAdEF
Al0wlV9NGKM9hxFZjh3cTTAzkGNUUIcFUKv30ddex2jKBq152axDmSRSrg1f51AA
CamCFJ1NNwxEmXbM6qvOwdzA1SLOS8nIKqYppddYmgEUg0/E+5GZaEdrxpWhx12Y
Z2ldugrEHOfc87w4aFym45/BVkkT8kfobXj8GHNVAChYvbDKwT1kiQAlJHOV8Oeg
RR7q/Fxtb9e4haOI+ot/6SMi+nfZpY7KFbI+2iy6w7i/W5Flh3p7phLgbi+QZS0x
dfUGCtyYHMA8/8wwymxdSBafZEi+Nqcf025g7t4qUk9wrzMGU4zpv2MOj3dzRQ+/
TW0sot7NiblyHmWhiXImSGD5jdBzeT+DYmXqfOFECyr1MBkIAyP/o8oBTWd6fS6Z
6hnFW/QKG00+366WTcGX3TsLV6Uubig4LZ2B5Dkj3Tu5OmHpk38vODD9OXOS3DRL
hItBvDP1nO3LgCOSdKodFO0wsm8p4patjSX6scS6vxCS5pq75T7x7gn1QdP+L0pn
lNzwoln+PGvHQvfDWjLELkzyYcE2876x/6+mo0pHqeq4DZXQNWqdaZdq2Noqmsp0
DiZZftayiOArFNtoZOM4fCzRD/QdTPFQfmli9Qd82HWD8hBzXQJIqjGmM1NH4JoZ
weEGqka0olDu5IzykjPGA07aYXYQEWjzWDJ8hZPVZfD0jn/9O1Rj+wfL7DHtpclG
Xd1sc0NzNJ+HafDnPGLY67FedyGwgYMkAgn7HA6Ev0ub42cwX1wdUICzrbU34Fna
JuY5w5Jlfz1US3lGRtyvpsDFMkspf7YqTIERv/2SmpCETTT6+p9mSUDjcZ+6ewg+
otrfzvhf5US9VdhFtv6zJ1plR/z1A8mybbE4MNitSDIupG5gWGZ9+Tg4+z2aBhRe
TJLAaIHl+Nnx9htHwJfTnYl156Yu+y7rpV6KFLI1VtSN7VpW9JyJFS/TIpnVB1kB
YBkTAD9bJ020l8zmgZvBquGQx/2kEytteOzoXZezm6C4tMcN1DPp0PM4R3xXQgic
D17bm/L2HIrVrQ6gmuWrxJsPzpYUDswlqRqS5cPaYXB0nuUYxNrbsHWtzjsFAFdy
x6DusYz9T7ZfEZdjinGNgcEbFgUCTM+sjPDj/pCsZXHLGj5yCRA4WWzgU/5TVy35
Of6JZyPaP1eJiwmFcwQr6g4WMXPkOf13fpyXBOXuHiALuGybQaseovieFYngEaux
wVQe8goNlkcorqvQ27hV/Ix4IdFGB3YxGKlNHrDocLrwZK5QtjlbWtcH5HPVtMMu
9XTtJlEox9KAcT1y21SmWuN4PFuPypKh7skHJfj4nhXgEa3fW9ZiqP96eC0/A3pe
K7Ee6v6zic2Oj4BOyHrouSsyok26X9EzjwlT5WnIsckOafHYGpPNQvGa2GzJUXU5
VYToEM4TgkqzvrrsRve4HieIIlY2ggu330z5CW8ehPIjo6JLSdQrpnZfxlQCjVtZ
oTLxn/2VZPkqd0dQYRB8v745/52LjPQLqjnPaLidQ2IDCu73BO6VHkWemClxKdGF
EwUdKpf7w3Wz5ldJjRGjVEawRLMODlEgdgrtQMntR+nK8LvqB+Zo0IAJJf/YhEtF
qFtilvyKWmXLDb4erjVIUMzlc46HYZctNd8ixEAQmwqLeWMFZDSiXR8K8i/jXw4i
iNaSDBsB9NJLO7D4vtv56veUg0O/qDeSBgYn7mgfwNeC7b6JNdpPD6mzz59Cm8u/
t0AoWW7inB8M0xl1gIlZ4+33e3mdmyub6FdILQRPehi35sBM5Gr4D6XHEHR+L0Yu
uaHQbhp3piL96g0vm2yCjvKwnmtbwEmSyjq9RANQGX0Pw8zcNpYU8UUDURErXP+D
wWicUGzjGX0ffvNpcpmSUqapbgeQzUt6TNK6H9EUh/Ab4Pa5o4AbH7sEytnxJS/v
NRiudUUzzAxWtu7sJulCDUSahLiPT5467VnK6j+JxZhUK/kVRWzJVmdwow1ijU2U
AHUIQ5ObOFhlIXESeIufrEqosaNUPsHtwDywLS/5e5vy1HBZohXNXOxLMLi8QJmv
tlg4ZHqT2PZHsWUsCHBHHSwd36ENCG/pbiUuL7ZWDqcXGPgmW3wfCrp5p+rbeKOx
7exa8IqLD9Cxip7f8oeLAYtTKeEO3m4AunuW92Si0CczBQxTABKv9ryTLoDFwyNg
k4gppyaiwK0Ea4g1peMJytKs3bWbuySKkWbUZbrCIjFg8J+aTcbwo2k3KH0wj6vl
NRkdmZ1bd15SM/xMlrzfZKTA/22106hIkVhGydALDRVnAYAMBj3hqOHY8OJYOBOM
WyWQ20fZDbl4j54mIdnHxXAsNsagu2k1UXFlh/rEfel1nIJVuVRruPprHKUqx1fs
Az6w/iPtm6m7eLMPL/2cLVZWKV9nopFKQhiSXQWiBuMg2C9oa7u5sqwU6dy4+Yei
EmVv9GDaAONInm9RhHDdHIYUDpLCaQgWar7Pz4FwCeeqrYAbk7FcVtOCMzT7hyEe
1As4AqBTu4ZNaTO+7Y3VMCmNoJoOorY+VcKHWM1Q8dM3AmgG10HKUgY/tfg6zJp7
TvevWjSvzyiAT9meg08XQ5+jUFApNAsII+bkKCPDIosRXn73/ONdvdT+tyU+L59i
nxTP9HP9cubdAn6aoP4iHcqeIpIqaBGfnEDbF33/ZZwF+GfdiLtxn3G935/sWBkT
VdiCSGM5A3VjtHW7ZQ4e2O1e22zA8wrMT1oYQU3+l5eP+jEwPt6XDUUh1PffPC3V
CZxFMUjDZRhAQbkx4jVvEZ/pjBoAv+8BDgt3QRZocXcYSrIfhWeo15A83s/12MwL
BEtigrMG3TyvOcFpDV3li46PmBAhxY3zw7wZR5fnbh2c1AQpydzc3joiPpOxSd36
rosDuIL74KgoFGytscBEIdCA0BtuexicpukMHPwUjUwI8YImRxjcHmhD4I6za7yZ
sxpd9WMbevr9xPDVrMvwwlkb8g+o+nTaZ5b6TNKjEeEgCXIfw/NY5ZFn/fQq8tik
yRdmMlY8rMq6cj22Y9GFNoJDFGA6OW82QGZH1H5TnTPU44VLBY5ZxmUuNGse9nVZ
SHzNz0FNqf8OtNdQjD0Cjhdr7V2Rcq2LqxLgjBMv8HM/yhSANTr2KKvKpa3Ksmpp
0N+VJrjTIMztHuGmnvBxt0WPOwh0xl1KZf086D8hEw/Iz8DUOxXq8dXvdwS29qr1
XzJgkc6UJEDJ4p77gD4b1SHxWmlWHsoEww0FsfQzXTCym1WZ4pR5lSG54LGCpuCG
EMUnxRE1cv5UaoWNBtlX981yf2HMZSa23NheF0jdGT21MqPB231yWVdBWohJxnk1
ZakCdccKufubroUNw/Fivhu05NDOhLuevxQv9sJGBiIWF4mKn5dj3bBfOVsqqUzf
/5ffS6tekG4Te3IeAYzT/EGVizw6NP/gnEGw3DxU7r6MuIyldlQnIVEZoibmMlw0
Ua8aX/aRhlrZdIANbTmogc6LBVeTSWhqsDsCVezydCVi+JjSLkQiS6Fu4pH4s3N+
eM717CqQGUNyD1grhZ2cbXmxj3H6HvRnqaYybfa6mZlu/kr+gXjJrb8+VAMIQLga
YmXDJ2SF7L8qgurDH6ddJ2W78LC2mX1vaWEyJnjQJP6dFPUZIP9GbolaBzD8Vr4G
17OmliaJ4LsEX54svXXcsef0SnXHj9+sZHn3Za+If9x5GesUcsZ4Ps5jRHM4lJ7R
FHuuRlTtpCGYwIdcoeA7Y6W94JuSyQF8yGWI8TIlttscJo9I9PJDVIYr/D+w/ePS
zL9GtOZsrOk/xP0hYywR7t8X1qX1O3kuvPkhpIakDgd/liLgWpHbRdNjLGKeQ8bV
3DvTsC8YUgNClx9is6/SVjI5TCNqR8Mwe/R0DrHvG9EngwWpLP3r1a6UE1/a/XcQ
p8CIEyditW5yzEvVjSiHsiPN2rsAqbDfV70l7Tg9D+D64APRPVXYTDv/IEUdvUTO
RSOPgdcl2R+mXnqxiiOoOyUel5SJqLuIrO580EU+PpgpSyHJFzyJKsW7kVtbXZT8
FJNK4uPugHX4WwpcIAF0Jqcox7Ce7irS8MH8K1qfdoFqltRbAhNdut61zz9mhcad
oZ3DrUJY7ScB7UcshU/5+FT5Hml1D8SvhJvp8CfYQonsDOG+BbNzt1f5/k0G8r02
1pX0fxK75CduACXUMmiC5ogoU40IYJnWPXfmglvMa2ky62qtXoiKL70KDNEFDdES
WxXMmvUHIzfyrHlg4OaXomCeKuOrO+qTVeh+NzubKs7qFrag3fcPDN/zAJo2bGX3
kktRbC7W5KbCzTOLkcdFGhKpfiQ9LNvCEV0llQZmZXwz8si+dvE8lUbzRkOKhu4L
hjaCCiFcpnZMtgh2GI5dgGnSBzIoAEcQtq3f6p56MIB+dJbh9Q1OZthyZYW9+ebl
o6u8QNRetcrZDr1sio04/Neiv5MOQ7SKOfl8bQwz/RIJ29dD98BQa1ch84uBqAGA
TfBxKMon0ECoUznjir+4STgRqablN4GLDDJe9PuZz8cZ8wuPb+TnNxng4bDB9xVQ
kp0C4bkiqtMunVEF1gnuIBSQLexBICmqWb+Gp9JfNZysZHxQ9raj0VEPmXrXWn//
pw5ZTwoPqNEMh9qGaN8iGNQGr0hb71+ZSCi2Ys3M5h7Tc99PYy9Wz4El2zOeCkLR
au0uaoGJKs70VNrAv8+zkxIY98flLqlbm4DuU68n5fpX22LKrqkdo4fLNellY2ea
yv+pgmF4Nf9xLI5MEYrGGdz3J/YRTesGG2gj6BOExxkjVPZdbXRzBu0yp5qEBR9m
xXJlJcXd/TdpWu7N2rVcYqXOR4GESsu39YsHSY2VuOR7A8fWdvJfMWwHACjJSF1d
TyDnH3GMdsl7kjfdxzvNaDaK3FhvCh/c7rHhUPqHpILMUq2oC4W5D8LOrMuDrOu4
yBJ1Im19UL3U+mF+nHNxSEVYqbsSZpSO30zC6g77QVlfcawj4LG3LLomcmV8tgvO
rm78neqiiEpzZELfsSKxkNViK3YeNxGUllWK0PE8AhFT3PuQaxtUOZB9FjBOpe72
IvKeCxDnNd8TJRHiqvy0mhsKpUkSZH5z+SHlAO+QwmdXXIXR3/oUVV35ELO9TGMx
iz/mSxXqu3c7NnvUaAX+WhJ4tWq973ZeeLHtf+ysDeAsJj1ONBGra1+yIxc1LXzL
g1imi1cPwB2rEfCxAsdTX1selJvQ7nGv+sktjswz8nAzrLpZB1JYqqv8as4gbNjJ
n8egNXy6Yq7gt5pOUgBbpMfnmoHWt585zA4fqjZIzAHebii0Mm6r+U68NhCrFiH4
Y+0qFwUxf30yglsu+wSxlR92X5TiqqmUsHUH4Ywfl8fmg344etni0Oa+rHTxQkcA
W+iCG3WTyl2JV7JvgMKZI41JHG9RJBw3nuRLiJP/0RuqL7NjqQVO1Jb9Izorv4qU
71bs6xMxAyRIU2bmxSzLuRImt8Q9wOSrePg/F70sBYvE/m0qYFnKDbp+PegkzkF9
PHSIM4p9WXBjgDG8IdDXp5wcsvKNnRIx0ooDnmakhY3y0mAEQEMmz5GXzg1dV2L8
/bz+HKs7aE64IA7yoiTjgppAZSHB1b4EnopZbVBwxXmM9zorbQBNf+k5GGadVvtK
QwUcvDwNKzrAClHRQTKfiEDGSBmSoexSmVbIhmgfqclHw6nqcwlwOn18mA5zB5CP
0dFtCrr5V6op76PnFqad7K28OwJamkiUV3kG2IhKSd1EC8ldBmZdkja1qOgQTAkU
mru6bhzV3+32GehGNu5rubEri7BEHE2rbaPleapfjM9R/JtLGDx7B9JIvFSp+/FR
EQPoIC3WoMXqOaFsWuBlpirDqMDejk1KubWS+n6RMJwygNwPsKISEhG1CNyR1Jy+
o9gGd5p1RK4jF1KB9UgSVAmLYYqByDVpke7jbooOab10XE1zbbYOg3AgW5HeShuK
g9w0Su5yysnrTYY/WilVSyX9dQj92Sg3KBTxkXVHs0lxWHGB//Tr1pJhxNa98co+
3o+QEk7wC8tDIamLhBFzO6BELCbD0n2T/WNW3Fbz40+YeUjj8lD2z3LCEKxM7eSR
bsBHQVfRv1CuMzc2wHqIkvfNzOGMcikAx/85v42YeKI+CkrTllqOgo40UFxHeJfG
aoH8fBLSlGqtr2A4VJFDjf1TG1E+upAFFv1v/T3tqyRr9nEiKYBciq6Wc62Wp3pY
nYJRk3O0UGVpAsjs0GGyWaa4kzCTw7rkxofT+tUS0wN+ugqblFRjRQeuNGwn/bFJ
PPUbKJGw41W/O7qTC2OR5Mj0BIUnYWXh8eaTz3/nzhLqbgB/5y87HexNf8eYfEoK
n07Tb2EGYhSkOyoI+/OGRoXDHrG/Ifj7AxHFP2pEH+RKF48COo9g8dgPg9KM0H21
N4azgw8e2y9Pxrb8uXkq8ru0bwnxmKMOk72z46KIhf3rmue38wEN/xrYQYjUcvmm
8FaA+EvudjKg+1RNZMRL/NcceGOY52JhzQm1/YG0VXuwoROGPnVfU8riDcDqAZPj
r4iP0PiUzu8yfC0Jib8YHyY+SyTgrCpgfiRQieN02m4gccgq7jWRZMAGqjD8SVUV
V6dl0A+0yRvYym5Iod/MOJilbZGSLLZajcJAi5qE6uFiU9CmbhHCE4d5hvR2HSka
bx7oLkDZ7ZbNck50fs4gujccMBHJrj4j08AyaUPFC8+GWNqQPcnbPod+5GX+lNRq
vo1QrShwJmxQzzQpASMEAEpvKxnMZ2HGkfQ+WbF1tgtCyqmYPKIirxqqWQfz2SoZ
/1I1EHnxOFtwYmvX+7f8FM1RSgQnqQzprhVNA9nlmDiSejBlb9Qv1h6iVJ5vzZwq
rDjHp/qyU5ru7PzCdWU6YnARqNP4sh70P6sDdRHM7yZ2Msa4+wABW657CEJ7qWyW
PeoPUPmLgeYtwhWJN8bg2jAwriDaYWjN+z4geDJHj+N+Hc+j1qbbwM+hiUwmaXQS
AK0AZ7532BXoaN9RODnhrwQXeGgXVG2bngwP4Hub4UqXLSp0aVC6Sjgo7GVjSFXI
J/3kdMUTQHVMGJ4qt9F+NmsTB9idCYoKssG06Pa8dV8WsVzONdxacyDlbI0QPI8y
a7ROkDlaRXQPr+mYf8uc7R6GKvcQmNck5+kAJ9+ycXUsw3SiiZ72BptJIY/4xljI
Z96cYKzeMurLPlRiCJx0ogPC50Jrg3m3UAsLNbUhMS2/gcAFYhT/NlXP2JN3E0gk
1iNCxUKdW7KTkBwgqYp764sPpuHP5FBBTr44kqFNBCjvn1K36l/qA9frEqtGgsO2
e8ihisvTsI0IXXXyn+6xwf0kwUIz+FjZQ+BAV8q0gjs2YWDJlvM4dkFT4BLfyi00
IPS4TUcLP+68HapDx9Z1YnE52ySOoTkYxGwXF9UfpHqc6hmbLHsoaq1ZHvG8RUVb
A4m0gFifq5UWe2PYjqEVCpQhRzXBt8XBKZWAyGJly9HqT2pgADKitip9sBL7SuJe
1mTNyNIsuEYcylYEzThdIMT6BR+ZMnEj7+yPq/e6URD/HicrWzBeEFW/QY9AbXQ8
FChR0IJQUXO2OtXkQt+Xev9Xm7LWtbEqsUu+/N/NXjXZzVvikEOmg7rb6SrRVEIM
jNOi5kIIqzvrP7+yCNVmZMcQnIij6OSbB9qETut573RZXSlmNppwf0aLULb2gbYP
Yi6eLQ3scJFiqTLNYjKTPegKg59kAdwKgaNIgpfF8D0rMX2vh5toc/HE8Y7dCDVp
ZiQtpX41r8mc912UbnAWaWGO1g1prOJ5PVGT2fuHZNS5ScCwo8uUp8mOByOjOBJC
Yh1+PJnnOwaksY1Y+KzGaIbR7oLqWkbBepgD5BFQbBEcYFVFwBpeg2UlJUg7WPzn
29UfvE7ft7FCT/OFaao3mO4BZ9nbx6A0BOtw42xA1bBI2aJ8MG5kW8jEM0SywAzj
z78s/oSkX1y4z4JRvfBqba57TwJzos5nMS0zcgqtjzt+UbmUoAv6eQv+fQJ7WF88
tSf/utJvcfKnseuHssIfFO9euwHJ0/J5ye/aNCxV+6BYwf9yMdNfz/fAPkWPzsQS
4GOxL9IQe6mQuWuzAea2M851f3NaidZjgzUyTStarHsklNMvauT6SypiwMBm+yId
yQuU4RidnWUDNc1sjvIge5YIOKpL/rXJjVa4s2S2gmuBxDInN80fWNgNsK/GmDKh
q5YmHMUIjp4JM3wsHGWpaEm2S6aVJ9Nz++qJielicFeT/ar+5SQghBz+wfQ7mJnp
xOvnmzny+SBA5wJqfGC82ubMW0vuc/iwgh5mc4NyuavxnUGFEbRgqtygpltOecQN
VNrF0N7KBXupQN8Wtcm+0sLFoWR+yu2Ng36ppaSoXLwdWRghNPVGOCFu/0uguAuM
/lsMjh7tODYxUN1DIS8hNIZj0snD3lR/BqzwNvMATKT7+geH0NiaNUXioHbxZxUR
W4UXu0QeG/2VbN4p1hMKaTdjgh8rfQwE8BWgJd49lhYL1NUAV0duaBB31qfzUDuI
6Q/eaa44rZUG87zatEe6AWNpS49nlAPT5oVNJ8Z2HuXIkXcRJiFvZAEF0OILi4cF
AInyo2snv6EOZDLZq+/39GoAkW1LwoV37o10bY6NYVIltXuSSITJ6pSTDgkwKl++
sv8liNJwosbWc+E+1FkpGaF3YtyLllG9NIMDi9LOWSAsftRS4xtRRuxJIq48bZu6
ilrWiRWX+7QnHf4sSjVrJ1pBoA2tbR6O7CJS+A3xvGMqDPUvrnKWf+oRemh9J/Wi
4q1EhFkq+Vj1k3ZcQSzyPs4/ZwsSdZW4KTbimQNduYNDeoXTl6r/xeOTMrkfLGKV
iPSZcl6gAkYmll0FIsE4nskrKKalcQmo41Mmw43/Q702455Z36ls/r2QlZXYv2DS
q32OuXROToyrJdt8KF/9d2LKGZDcaat6F+z82QlFVpucarLJWDNCIHr1gwGySElq
TQHexnNH3p4k4Dwl8S1D3R8dE0/dm61IvCiHwgM5Od0kfcpIeRMgiXm3EorzM6op
lVEdNOApWPX7gLVRYmPU+4afkQwHTn1oVJkBANhWjGOsHrsr+gQGVw5rwdLNJYb0
tIXbIpBHyAji/G8RGJnc97sHK9oYUtVr0IZ4bXK71GsqPM+EuUUh3J2f661d3pa5
+tIXCBdYdiDc+VI9FpXSWFqY16a1nF5vbcX36VX4lnaD4vpH/+6n7SpI0sswMjqt
8yGAi/4TrSYnMwk440BrX0XPfLS+909CQjtw5t0vNzwPpGJqBtIl/5jr8//AeKdm
t9HDLUZN938FOa7eNg6frXDKF7xrDodYWbu23zQ3O+uNd0lKyeLYN2xr6aoPFwg4
VznGwF7VkUvZDlMQ/3qY7xUFeWpV4VjoYWJJ+edncnAY5tMaJE2qSRfb3MZ8X4B5
myzBPssJueMGQ5afgR8+HLmbb3Z0Owfxo8QgCpi+4sKoFzbhdU1H8VxqxDs0B31f
3LdpUGaDA8eLe74l1brb6sNVujCg0h3cONdENOnEPPLvpVyP9FlPUwd+99Ifevw5
au3ezJdOTp/Vz3O+pKFqXJ1Sj9A3FFOD3YCWxjEKpY9J2YwCSkBmF0yxf5yNefWz
mIN/k9mCJ/Z+aS9gRDVl844Zr1tSONpAMPQ0HBoMIIDLZSDZFYDSLkCLMo2ie7Oe
AFFMUNV6AYokb7DhW8KwCiFQ/1cNntdS0uTtIny2BJFMvQaaQ2ClaOHIodgGY/3S
yyPGyos7KEFe87lIjDW1y8r9lmzzdUwYErwTlqG4ZK0rxrco3C8RIghtynvodyGs
f8Zy42EFOb6H3itOq080whk6zj91XsAd96B7z7Qh1i6lTDcYs1KTJbBFjF9dMvlM
fJs5EwOeH2/a4cSdCnocvw4kpqRCqKpZgKabRta7HEwK8swV6ymqrWlsmd/qE+/o
8qsv3st9Vj5y3ra3atujZ4Yq/04ITPdXbORhxzVuHis2RZNjhEpzgXISPeIa6lq6
YjaVYdO0SQZ5LTTv2naVWljQFTTvpTdysmxT1rN+YTVn+xLh1epsooeisfBESqvN
wOdGvsR/Dnyq7hIRp4hAw3amfaxCb6Jjq/jxocX50apbomSiOV/gUdtVPYti6XdZ
j14mogacKttaNVSJiDkOVPEJd98PF3D9ifkivgZwGp6zIJ57LnhqkIs+F6QUvYIM
4XhFfsnqF6hNHCjCxfh4MNYB41ObqLgSpQw8BfJLbKNNIwIauAc1VZnX1JtdlTxd
aVhTyd53TTy5PV4LUMNKfVYd0ShYmeBHsRehOV1ZRFByqFHaFAkFCvAmh5D2EMut
NvL93Mqbr8RpkaQU5GsEvcVxltcDSiTIqLzKXKqkTBEn6gm8fP1P7JM9C3JQedAk
s8xpQ7xrMUYRYcXeasETg8FnhiJuupMSY97qCO47Op2zYt6YV8/X1xoJkz3QVDeS
CES16y3X0Ls8fZCAZXdHqguBhaMytZmgpoY/XCwx1uej3ZI3Ej40lLFWafp4j9mw
qfo/mC8F2EfQOKQ5By+yvgGUMT9JE+kRrSDNMtqnM+TLPm+z4iWsTjDzPUwUTZr+
U8EB+MCgi3s4cdFgJBQ2ocC1AjciJpzcG+BZUyQJWKsVhl/lnF9+OkZ1s/XExlxX
tlKUT2f4W/5eBi2NQvjdlljm187x6s0xB1rFrGUMKfgomG8CL+gUo7QUrbX+6IJR
1vjSwuoibE/JWXT32QCfzheDdTiLgs8kQLQN8pZPuNyvpzmSqxB6+z185nI5qIkU
XsY08X9xIPF1G+g2CYN2LOJGhUxJyBwSUAlQe4CT/QIiximPtM8ms1vjxx5dxrvI
AwKsVGfsyCAll/L3rhkI7AuJqPMiL6YV/yYaEvF0C5b8B86fVbKanMggUragN4nk
2fSreEME3jEPJNOS6my6xDCWStlxAeEMxOl/c7Als0oAuvNCYMQApLc6YstHISuk
b3J6gepnjztRder3e5X+tLiGPi9N5tdQPYnGTdKW1CtbmXLYVM6QrVAwJWe7Yv5R
Hr4FI2ova9wMIzlaOOwz5XKsQcsTKne3Lq49+gG/Yi4/hoy8MK6fsBx1/HzRr0ns
38PufnronA6cCW1aj9LmfYFeB8z6BwhWx+gYmHVSx5WtDegGMhu3YEomswRSW0yt
Ub3b1Ue2HiB8Jed1XAXzHoAMR5/bxIyFRcx20/nYOrlbA3yHUY5JKrkK/bmHRrQK
j02yG7XIkvqfulK0BOSXt5G1HaCbOU/orTAXGuOZHJ0Fo8lFlDJQKes7zFugwaMe
u1huD4LS9m6/tpAy9IbI1hzDqB/PNJTJCYVEf3xpvWBVDBwPqOTVeKLE8ts+4dT2
XjStkgmBTPsqiRWIEQtFi7cW1lOAYQssZVDAVMZBEhX8GwYpE53m2U9vJ+eT+VI8
I0PM+UOJYM7az2TsMERtW4vz8Lzg985hmzoJD+iHFkbpdIUDkm23KMCfxsFVkU/d
/kwIRdvAVlT6PhFERcWt2/ewewmeHXFA+Wy/LeGqx6bLC+cRYa+MXUXM4osXeJfq
7OnZMLFs6AmhhkcH6bSiuimnc9emtGp9iDaKskaipuaQglsty+KsytV5yNHeLpIk
fkaTe8rYltOuyKxROwD443TagawZNWZO55s7Y43nNtzja+C3J8JmQNbs3ZVVUt9I
YFQpsGocBP2NPBSXDibztcadUzIPTiKQNqglOfnQguku3oXAxy0iTT+g5AcsdV4/
8Bvgwnion7HB5LezK3Zn/y80nn5LEwq6y73NHPqSi25mG8StUWBA17nTpUo/KKJ8
lj4p6Axg4DsLYnHedTB+kgqI/pW1YM3YNkbBKzF/vlvNObu7PXZV8UXEkFwVQqSM
esW9JLagsbKjAtblZZ3gZok1Z5vCXTHkLK9tA4KzOnW8zrn4kPVF7jyEO5a0AVIZ
sRbqOi7CAF0lAL0uZP15JX14hSsUmao8eC1kMPx8deHlNOzxTfLqji3GOU1sXo6P
24bXdLgz7DS5oXOR1iMjSpYnCqLCRD3x0FHhAWS5vaVeU/4QYaeYSbggJatqAG8L
gEuzDRzAwnm0TRPcaoXt8eSaqjCQia9nRQeQFgM4zf4fY8FzErPgZswWUkpnp8Yx
WOdyteTgKUWpKthdOgXPs6PNUp4vzFBVFkJGKe2wfITDqlnjrsvFyTQ65ffF0oit
BLgWP4uWlhGXw4Ty0UaLBU1R4cJ47J/JlSlI8dLHHEY+122pS/+26x+6s1LOP7mj
H6Qxa/U2IgKZd9lIcuV+tMK1yFbH4A6ebqE/MSbtbkHKOxOindM9wP7HAdw7znXN
UIi8ZPGxCX5JO3JHNnA6RaUz8U0192W4tS8TMdeRJtnLUgi8eXVtkIEkTA953P0p
6W6sTBMdExxgr0pV/KjZCDkIC2wUzUD/GEKECH3ZUkmyXKxR3rJWSzcWqYBTivut
F5i+1U9EZAF8NufpY/g0bQdyu/c98NLtFu3Zpr9NYDlxUSnjEpLW7Nf9wAs/XWbS
3xeDS6wS+WvIfeR0iS100MZwigdFHhVnk0Opt3waAPaUesKatNLDnKWBI+tFn/z3
VBFJZrGmSsT5HSsWHheOAS419Mjle44N6cGu6HP0dv/gHOcDbLUt5RTuTdIEPJjZ
xVzwsIHkDe7j/bVat4I3qvpjtMmOQYeok8i7GS6Ofrfbi1btaOZHBkYvV7rAQdrG
kAejDUpxn3az1lqS6xIdk3zKskNHYDv2Eg+7DwBq7tWJQHcQ6IIG1NHtxBhBqQiH
FcJ0gaKErjmOlB3okDBn0natjXi/mneilkj5K4jxE4un0bHYcCg6EtV/AVktXGcp
LfLMCYv26b7ArggwvVMweSYU8HVApVKLqXIlLBG5Vpk2cGmBFgog7krp020mM3+p
tSV38kAannjdwsDugZijppdOqizbtYRnTHcu52fQGyawHYS/4CmekMAzrv7b2IF6
Pe58ajIby6U+SlkoBv8SGD9Vkui70baLkuWK/bsK3BjMXdbI/Upr3YVjYYoFJUw6
ykAHYqlrbvR6GjI1yvxZyQYyhfme25gMtea1b/zIghjEeEoHAgEqKADgF9x3yewD
DCaKvYFwnup740qeOv8EmRxFyhxMplCEsaxmD+sIFEaAT07OUEZh6jiFZ/L0ddL7
vYT+sPg5OLjbefoXBJaaxm6tRAVkMI1ihENxp2j+M+P+cc0ubvDYYvu08G29O6at
ky1wFwsEoQtReEq4czaiU5JOYNlw+i85RhzoTHafOf7m3Pf3RKpYnsMK9kNVnLRI
ZUM+LxOeyQC2gYRaCqB1Sz0H00JkFKE2b+uQ5Ob1J1SzSfORhUQyswfLDExAB9pY
MZv2F5zqNy4ZY7M0H4w1jn5n24zW/HVGDwivkouO/SYQLsuNXAZHyxp9RnaimZUs
N4l54HcGuFsDGMtD86J9u49oUGBZ3KJ20EaYsIdidKUM7vrRBe7YHtEs6heaMI+v
O1Dl01EsjTNGNqqB6xzy+skDolr1de0VtsGjKuLJM+sut0aC3gV9J2dKcXkLWKKk
GTiD5rY74J8Q0MVS7s6CbYnHSU8AGikA3rna8x4P/It0U/34kz0q8WEbi46G0IBK
tnHMTaeQNGYhntD7Zo/zgRfHgBt3ocabzgPktdzMbOg1c3vTJ63c4SY0RA0IECay
nC3oNLZywPbZOGWkP7jcgGR4Awzr2UMUqI9MOjammqSp79TxCEWUS7a1s+wqQyZe
5XxQlxI8wm8a0jUCyUodBaS81fzPdId0VbcOCO4Z0to1F1cRRVcS8zkDSchJQMtz
y0lfliGSVkH++YanLL4wkFcsWmJPZCyKV/a5EBjKB6G71JUtJDupkl64+11KHhl1
PdP8kyODoI+yaV96tGRa5Dyid8QwU6RH8AfqEPmz4n1NGs3xJjRVk/tVUK/AFayU
2y3/taAkh1+77N3eLtMsqOXMH9CiaK5PsUg1Gp4un5VheSgB5QosxBUvLL9ibzr+
PPGFzbf8g37Z+9FoDl2lxqJqujnhtHclYar3qZPf3wXIUTyEB/ODn1Xxm35l8fXm
fpa6U9uLf6jGN+YX37aKCdw5SzAjfJotTmSKZOCiWEQ8VSJyeTojmc5qNtpjNA6C
ro4nsYVR56Dh7DzBqhknXOxmm6ZjhLcHQP+mLLBCklAsc54lpr33dwF90LAJO34G
adUfuEo5r13VcGlJnjnuiveStSsnIpGMc+RKTXKWANrQVt/BzxT2jdmRlGv1T41A
n0vh8IO5sO1H7gYYKYcKVP7HiWLvD+fiONkK64FB590pQZUxHDTfdB9VSC0jUpcj
uc16qkINNhbqu8M2T0SBTU1SVkgjBCgarMitwo9M5z203DNtXQDYIm/F30gSabhH
Zwri5DOjJB3+DezoEhqT/XEm5Oh8MAGvH9THX1dnhReFJQnpMTbFO+OPcbUra0+E
EYEaj7BgrNbFEqlDxXwE5oL37pPFOtFVkUNWxMLv4VMWFGX2VZKUJwPmZ/UJnCtf
DQQuZAavG/NEsRy1cwYOEccNGyAI9bW42dpf/GQAkbpQddtQxj41ufGSZq4FCnOn
I/IR27TtuE9MLrnCyYohZdW4ZN78ClTsjYlpY3oKmPCLsPjAuzdmAm9Bwv2oAP18
iyUCgV7bZ9siP3Sqx4PgZisZ+CnvyxoRNCR2XRAw61DKnc77jB816KX0QnTdCK3V
l1at+CNsYPHBQo7MyGqeWfuQhRIu5UtN6GeNGnpaqFCfAqyCWVyoaSiu1iTBT5y2
P289Z70DJtSmR/iWjZDDwfnudTK/NFgQcUqaaA8PDDmDYxU04wWSiOsl4AzsKARC
e9RynjNPUJmHnrHg8OPngD6CmbwbHPitUacl9gA61Rz2EtNRKtpRNTgr1Xvp6oDU
52Tc8he9AmOpJLDjYQ/Za5JLp8CHhr1CT6ZcfKAUQfzFkmL+IonRvufCHYmSDPID
DjvvMcA3FBahtwLNCAq+jRwbwJfLeyhvi0nPaIZ04n54fZzIWLoiGqo+wpGxhduF
SPHm9qwbjgcI+EAT9KYdPgShN2Jdwa165QDiK/u4Rnt9N6Nc5p0n8uI8gyF9/veh
J89YC//8Kwt2AEjOg/6MQ35h+q0huW/5NFgE5RcmI/9RshBpViUNyD/Ej15UegrQ
Ys9Af3fFW6WAVX1GQzOdW/PiPfW/o1UBE9HTomdQhqzgXvIoODSbkJxQK06/uk2O
H/2kkPHmg9C0BIh5U1//4RjFXP3I2TR2tAT8W6uYCCb5YOQ2PqZ6DjZYuRI6NjSf
XRKwatA1V4tdp3TA2odzQ3uQ6oVllBd/kfmc0hUlcL32NCnmI7qq8dUjr4R6xr0v
Zoov44CaRLUd6jhe3NHUSDMfQYxZIrja4Elq+5f+dn4TVYLOR5zPaWRZ/AcdR2Ha
6Ko9281ZeBtv51astTqb16Nk6oM6+Rn1HpFwYgy8ELbUP/kC67lm6VMPn03n1jtt
lMU9LHYYAW7ABhEEZOhthIHXIViehoQEMf+b0cmlvWDSHs3kfT+mfXb/18FlTmTB
IDbvyi0rs2u0wypZlNHHlfb1GNL+0XFMnJw6VQc5MRTmChkCPIyuMnaCGsqDX9jM
Try+Fcx6I1SFSGRCV5bFL/4Tsij283b1Ed8UR75C5CBo2H4E8+twfMIOU+buk4UD
bF71h/OZylCimDOpE03m/ZuPGYvVxfS2ejVEirXMpRgF3YOvM79qGkJnhrljZnwP
HkF+BzSfUCTFke5DXVjJ6m6xUnmLsUZoWJFBGBdsQGxck9/3JrZQaSobFzg5sQTr
pF7NXi/aAiivgIGni/qvvj6DkTsonNM0AQvG9uFo0qHLgbt5rIyyDpJTQ5P7VNRr
mrQj8HdeMML3aJfcBblQ9h+htWlHWRIOONTM+xkB2mK0NyfRyWmsmQjy/d6p8owf
TkBMCBF8b3ZfSvEsKFNGyaYZRF+z7S+fs8p6rSuta76kY3jchtDZGkxDqmEwrnLM
wTba8OSWgni9qj3v2WosqaYcTQZLYusff63PbmdfeqE67HDuz9XjwEYIJtQ5pKXN
5TQBTAb5uhVkLIhEjhiEbEurJBK+W0AA9alZcgx5fBRSdfW+l5Hn9IG2IR+Jqe09
FjX0f+a+SiN+04olle223Jaw0IFqBSDg73vcjS2hHqZeEUNasoOsvF2AY2VgSLIu
kfgPHEyXhglPFeXH57zR/n22Nt99padhAHma3mLz51Ypg4NTL2k+xJ+mJhr8T87/
Iw+6fAH3sgn//DcGi3wgi5Bxzln9emGo3hISc1aoP0N94r/JyBAfGkR6G2Fu82hq
gPRvMNcalnihUeHKkeuNjzBK50hhZcswXLDbrsJahUN3T7S35tTeZ8pqbSH0Sx2Z
ywC5hBCdsZ+G666Foeglr4tdFXymw6j4VAIpgDO3hzOS52rHqWJ/Yty/gOnoJV8H
yVfZolhGe14V5r+/xTs4DyawAZUFsO9CrVYBuHh34ai376jNBQxtu/UpN2b++np/
/ynN6Vmrmiagh9kJdNaKGML6mMbI91/XZBFBHIWcMDqPo1W5ZS/bixWjbyjogkPH
HLZOInp84QKQA5XWBQBt27Vgsl7RpPmyEoJ4u/xnA0YU+7gisrwQf22+C228MBK1
mal2sNvImc6HddldnSq26srPEt26nRQvPLuIckj8Keq5s6Fpag6PAInhTEQ+0kCa
ZPFkl8FLltX04dYzzqwHrbrSj6fbdXtV2BWCXjT5Vv9vZVeL4dAxDYomdkc0yhi2
GVTB/zuWrfQdRWz7RQNva7HaWO+4pWXbUf8ih9ykn5cVSwruWt6OZtLIK0YVO0C8
5yO+MXjDz0fV3RgnPwLpQeYPIBXo8iUkdVreXMzcydaGZ+9IPXXJ882PpI9zPxv+
hpxE9EtrSBFpPNsbOUhiQNWT76Sw3BDik+U84S6yw4pRIDpDZSdq36kjyvLVs3Ka
MRTkIvBTaAYEC2UsDH82vC4qxpbUkYnAtqkAkrFP57SRHoUGssiZT7fm6GHfmqE6
erG+jPSxcHOrJZQMFV3NZcxLkMXbYGpK0cr82Qt1h/pKGow/ZSF2ShR3SIEkEvvA
D6Q34tzVW/SxwlhnNDvHoWhZ3dSWsMEfRqV/dpqi0lCbTLz3Nla0ZFqNZd1ba9Ka
c66N6BwTyEyP8xpg4/Gno91SfbnepYQS5NQdc1m269RI4GKQF1wdls0VvzV/fHJ9
5yuvjQMi/yEGo8VSOmhF2IzUyTrzg5x/QVpRYCXuJpYNkiBxNk1k9rvivqJGxvGO
j1Nb1RdqlB8kJBMDHFSINRtYmIDd4iDawPeXoOPGuoRqlt3Fx7pSC8Uwh8e0SVtt
pbIpiZjEVHCN5kjK2Ykr3dyVA3YzDQemZ8tP3E7l8jlIjUoGotqZg2uo2EKFUC/Q
fz6ieKzlHMNV2f7Ki4nFaxpjx59ZwUk7OOOs6AD0p2Mt0Ihv2ZjysXoZQ5mMmIA0
m2YhaFQTqUBC6Tv2sFCd3GpplGfn9CmRbd4FGT/SfHLC9euTrOke7AlVX5R7hc6S
rCxoAXzjR8oaVcoc/V0GYOWu9/A1jbP6VgqhTgLlg0OBCOG6RD+yq7JkvmTbNBGO
pnMNhUyZrcfSgLu8iEGx2IoZ/CWovYm0IvCykr7RxWH+nLsYp2f+sF6wJgUyatmR
q6yimGtO8wJNb1NTYB2KJmwAas0uOB6iKSc2MD+Z4NuqWecl/wTlpzI2sMR986ng
hz7HKF1l34jBdfBBr1//GNKTfnehYJiTObdAOyYjTSxLpi2iMXABHRwQWZe9rVkp
u0UmdO9JZ4pb2evRZFACxXksBUBZt4zv26nGTUO4UcLtx57t8Mc0TxQRYjDISB13
86OHoejjNzhb5O/lFxEFlpBSOuoHTBP6R/RViHphy42T4ipSgS3G/FoDf+MMZxp9
Nm3ICswTfbDwSD7N6NgZOEX151XQ1Rz5jeVipQedh0L4VOeEBAsbSzJBOEchv8aD
yAfXZdAK7aJpop80pFSWT9ohJOzmsaXRRT6AsD1yTUTojV/HF3j2n/+E2bbIfCx4
0oIH9CRp3iEDYm93xKxLpAdQ1owAJbadfLwiKENCT8w7Zq80xjV2sA/AubWrsAP+
g5jPk3cKDNG+ANM4biqHPYseOHA3mppAHE6pxhu3oHCCpsZJ01twtO0VZXtQhrYa
i/evnp7yJIRUpDjML51QeiGAP7yht+c0bgDgEj+0+a3rk/qFW0uOKEfReddVB3pi
HIe3suUq8wrOdTUAC6jZ8E+aoE622XLa99z7M57ZA6jERJxzDBRIEufY48e4Xs1h
MmyONPi9n9++1WsGbf7dSvgGjRxofJY4JkWViV00BOVEjPT2hMATE3bk+lMWdts9
Ez4RF5Pr0fgWatS5XaiHorIGqfrXG8qildOTmyQCtb2cahP1FFqtYdzrc/87gGeG
RTiXs+qKmlcUiCnJlXHlzTcz6nwH1iec9Fo+Gc0kedn0dd3nFAGUtnHKH0TDh4Lm
YPa4XksrY3m2G91jSaSvHeK60vlDyH3nau1YqHnmtJKfqwRQzjWygn0r8+ER1zso
oat6EdG0/i5seMEwEvZqN2zCUF7wlD07lSNUSY8vJI7U9wkJr5zEsrRNutZTY97n
zLHVRdZ37a1fqp/Pf3+sJ4sZGjorsxCNdi04JZ311/f59akYBU5w8xUpmVmuRTfK
xEqWc4OKNbPOy854VDxNKOPxeuRWA9QTBUE6wLTFSCi55xazDeJC4OqtYp/qG/Zp
MewnYuC99H8pBsuMu98mJgXG5yOoD556Dvz5L/BXUkLjK0PWyRM5pdHMbv2TfkZb
tOWsf/6RHcv+Hoae+PvnRphT7xgoSgV9QyrlDHVQQBRMR+ecNOn8axMew8drxW1c
DHPdhZkMZIWsBoLsH2Tn2ByE/zADTw4/uBtPyVu8IsQojVqbjhrl03NrTczc3oNz
NFE6coqCubBBvtUktrSojGXKqWLetlhfoAHhOgpsfyFkF5sCC6CQ1DtYAbhQxLU4
8GQUHkLQ1SSS21npaV1rP4ONK4WFHbEd+pRlD+CI6joDC3CaSJM6fK70uAgdciGH
bzGIUGevhb0+MQm5PyD3R06fuA7wQne3mtM0hki4EgtOCZphklYbBx9efSdRYrQN
KLLqIqfEKSnqs0CcWALx1sdVaRG5rSKqrM2c+uSSBnCRd3E/x2LxxjiBGjC3AltW
JoDgK5YUiHvAUKHs1e5l1ZXK6gd2xyHErSxmdMESFthLqEn1L6sm5y/iEflc8kPr
+Cynk/82WeNGvuGlZEgPLw2j97Uz9hnH8RkroID0dDHSPBsRUlCuDwFCfW/AA5RT
pZ7IkPiyNw2j3S7FZbhwA7XHYXiwyDFEf+/tWUMfIgGnp56ctVsz61mHkuI96ONQ
K0YmSDFVFpL5l0eE2VtgMIRCxI/whnplWeB/cxjKsMwYb/yh672wIPsGCDhIXFIk
aFjSsnKswQVUXgZtBOz6xTG+FYSYJUVn3Yq9xySx9582jE69sranttbooKA9XO3s
W8EoGLtA3oCqzxvgsKvCiIfufjbupDzdc7Uym/T7myUwJLEJxvPojC/HaFEtYglq
Ro2F+chvABaVPrWL3o+WOYpfsKQqxo/B+AtXVE0/z1Nepbvp+DSFPVOBpQLL4ABg
zNIwZ6ty01ZouFlojSwf97PedUjYRCZYhR+9qjUNvOWkgn/gf450PJ0R8sxshPvh
9C5GKweYmPjFpCwFGxez/sdhecfckTl7v7uV4G4vzkv0o3ykyR+ZPQSzAciJfOBX
4BitssknnALLxADvObocsjfEP4y3Eh/3CSg8AO63HP02/CkyosNjWdFwNMD09UZp
6JYwH0bl0UFVXmGBabGOEJVzkHehQDMX6NnRS/0zzjOgTZy3BwZvqlj7kROxqXVl
GV0sGZ+ozrRDfeuQ+NgTy7kOZbO+PzR/nt7LELYREHEp4DLHcFdz5enLBj8bf9Tu
kLytmZcfFMQU+Z0Bbgb3q1xLJbLzr6ZkDeJ2nEqpAR6aEgW7Fh97yxcHdmbfksCA
yVyOtCI66ChpfELkQ8xbqekHO9OaohSvZaVh3kfWu9hK6bbCEruNmLPGVKHBfsXD
7OJ5plaIZh8du8XOYCoKrwCj8auLKAZLROic7MUFzqka5a3QlUIyTo9T1PvRy+KK
IRxM0pLm/YZz04+CtM3YGOcHTJNL/VaCagbX+AcNT0F2bJO6z+d4iBT5xZf/udh4
pet/OwIJLrrxeYfGxfL5CCFoYydBjP/09+LDnmKUYZvWcSxDPWjGiqo0CwRhvIeX
bnp7fMUL63tVP0RPJGL3JIFfDQGBYq7YKx8iAcmI6TvaobI57MlZ0juw+iyII0l5
5czy/o7Tvs45kaOYiMwel9suDAVhsWX6ltD6xGSwsN95v9I28zUbidyldKHONWRQ
0ClNuJJybqNJ1m0kyeeKpXIBGyEu9muvYHBY8kOvyRInUmAhqrD/5uvPBXac8WkB
yqsHKsY0odPhaBnSVKDMFTRIOktIbuaP5gAmODBPai5GBK77AbWvgCvmv69DR7Nj
Da6+kDFDFD2mSCjcTe/NrPweh2F4kYEOyUfxLGH2Hs7lLfd89RpYnrzCtdYD0biU
C/IDy3cLmMp5mhVg96X4tHpr97bNBU9LmkzynxUpAHyRN+McvpEOdUO4hblTxBH0
kUrUZaRXrcfhIKEPx/hNZ9YoKTFPrSWe/yUuIF49NzApO6nFrRsUnizYDHJZM+PT
V5o95XwyjdnSLy0jJuac3Bgg2+1Hw64aKfqDYJbfprXXPQknxZyQdUoLQz41R96U
qDOfUfsU/s0EVX12TlzyFHVGtmietjjiHUwZJ5PGAjEkyua7VyhUc5Si8jdTRcYl
snlaZn2+dm4p9MFxHLB0nC656Lb09s640btotZVn7Y/0AsoLxDo5W8a0YHiP22Kf
WTCeGwClYfsnek6j3E/MOGbLaQew8zK5um/ulzBarO+W5cin91E2i0IM+vimCL6V
qNc26iS33uvO5UTGSkebZcxC9bn2Px61+ZkqhUxHBjmu5/OXqTylYMRKFOcWocT5
isCOxn4xXoTA3RK3cMxy1qXgP+4IYHYy5f11MsT+dz8dNj6PJyMshyCIt+z4WBn0
vA3SBk62U+xL6N5KNoEnLwtrujjH4AsxaJK6CRnV+GnuMPgsOPwYjeJUQ11or0YI
soohsVkVL0nxTsQd9fc9LweIj4JFdMBQebf7kWdnetzIRX3hSWxS2DbtbpTZ+wYu
2s9xRzI6ZHX0JFKNMw98VZaVsJL7rfaiG3WOM9422iyUj2emQ9+axCvyjDX3ndT/
PWa5vKhXWHJLJuH8JivIwXgYEsp9Fq9YKqYNu2WaRakXkMxICjjOlzOnEsJcn1xz
8HfmcE1qR0g5JBhGRU2xmGT6huST77jLHZE5ic9r1D7Ut72Hv1VafOqZ/QXlMMLa
xh5P5CCa1IInmNUXh6B0BWChybes/o2Z/wzhggo2ny2/8gy53Gjz6b+Em9iRvRR9
g+tY6F3WN/JpOLUyjup4Y9/icAH3zZJw67MfgqFJmZqOccQYQVfXyNibcXeYyF8+
WJyRMIRBoBwS3hW3MNSrttc1xm64rKI0IKbHTpotu16R6sHXQpML8d9k5TJztGC4
aLXiw3QVxDKHXQpaDwAnrdnicGS00HZoxmkQwasEtuSa692TVJeqPwtPkFm4443T
WX8z0AMGY06lmfwTVJORtZ57AVusbwCuTjrRXDm+DH4+R/i9X5ZbZq/CfZ+H12Wt
Lkt0k7xvl+vjkVxUz0RoezTJJdV3t4hSlJszAUGJ2M6Wa11UuPM9wgY5QSbA7N4S
2k9NaFQSKwxfiE6ChuneYKumYuGUaiF9ZTrWOuJeH4UR/r5KrZjibM62LvPRnAT3
jH2egXjt9+yDp1BKjxOQm39PJ6dzZjlCjDgq5gzCXJ6RNelWzzxLQYLh3aYHmHLk
GrxBz5FRbIplcVKaFr3i2x05JjhUX5hMtfZvX+MFKA9zwXbLX/j1D/Kas1k1bjIi
oSyNOyHG/HSNZvuK0IeKLLBWOre/ChCpO6Dub4AmFwiCp9OsK6z/uBJEtxClvg9L
0OSAs312CwoxIzIe/FGsuim6dw6b2dVTGwtzng36Gn26u/0R3/Ku1aonuajPT9Ge
zs2/4U38GR7jRlwkCBaCFnbP03Ey7MxW6WIxvMOjyagWjEuWOIxF5s41JS02XDNg
ynn1+j37yfcM3c2KdMXi5mX8f12syjO2n2VLNEY3BFdiLekncRHA2MfCOlB+yZi4
8chCPKf5MWSVioG8SbMuvhamshnHV8uwbV9M3lWew05fmdAxnoDm52JRcASjrOeX
B1JfgVq7MgkQhsLOKOcoVaB67d3mn7Oh6GrNoOyoNpCqku1Jim1Em1OmPfp9KJe/
mTHT5Kj5UzSbm06R0mQexkBgIlINOGVvoj9vrqupZnDjQVjiYnDfrL1WcHUDC300
oVKSFlld0mNiArFAj7Vh/sdPgu9savlEXiX5EVxdP5P9jOpyHgZhpB1Nzp0Ldn5T
BSQIsTscR0MihZcie64L6r13e1HYFv462wLnXxbw0gnBVtA07UUE0dG4L4KkK7ri
dvkqSTm1u3oyeRIa67LyshiWqMmPmfMlWaKZKWa7N52qdeHeVfHMa6THs//7D0GP
2ZIStgvjVV2huQMF6sr7pPrnBjtmAtiT4ND5OLYcSmdmrL0vyccYCUOClo4isUgF
qKkcoukEdcNzEL8YnbKuCa0e+8TcUAMm/ahQLrhMno+3DUze4jgi1jXLBb4yDRGH
0mCXG3FJoYNiIHVfKBN1TpKq+oQA3R6ZnfYPi6jkguMnnuwCgwLLgggNw4NoU8w3
CbNWVGs/akb3dzoH249Nu8qj5RTKSHNkJsWI6sBgJXtAjes6aLo1qJVcEuBp0sgV
HgC29NcjSdoPrL0wgGLHlzOy38zeUm5drRfjszjfPmVFWAMsHG+1lPxxlyDbbkuD
AWBjM+diZR5/wYH7QY6MM5xXREhfSjwEuzaTrK8aPR1migcAIL7tbNVnDr7YZwGB
vXw9ii/5TT/JrjoYrv35cQa1ak4YJsynL0ubXHScHM3oakSq+vCyBJJpKYHoN4P/
YyUHLdhcPV6Pn3lRKTJCcJMkf0MZA/63cHaPW5pI8nIe4Jtfw03Q1ec6Sz9Q5q8B
+GDVTjI50wp/Q5jd23+wgvT1fykAcFEFubvvceXA4c9lrpIeispTimjDp8zQaOfr
klTM74thRtz35vQppy67ubyOEDW1Ck5feUn6hLVxv8Z3EtfGdBxM41oLMUFDybWT
lXrb/Y7EwkhSNa9H8IMN7eR1xik0SWaDiCLPjHb0h3Aq9+FDVhnNPQP29NBYLN58
NHBpLJHGbqEpNvO8uipTthUHWI8qyscnXxO8c7IHBPVJh60sTllNb/WIe7NBp3aB
iLOu9GpA7ipU82ZUsVer8cxbQyxcOwyfxfnIlxhyMuOSDc/e1r7xu1FlrjGhEaWB
O54eFVhotCIV+jIu+tR5n31xyit3C3li67asGDjX2w4woI/HptV49FtdM4TDXKH8
3HAgseGweX/nNAupMwePQ+oKxzSVVcDJ4Qmh1TITP/zkVhExV9jrDVNA7eUtHRPx
qzdeTYY1bjelOtS4Z9vB+jzrLjDozUwEHRFZooRgPqO7jrAE8g2OMXifOoKQlTQ0
krwVWQ9TBRBWCXZ/E6ZFPvSvz+pox1dzBHx1IeeqwENZg3m55meR5Xi8IfD6Jw1S
aJmtOikPFsD32zNqDAGAALb2WSWBQ4dRK2A5ImCJAwWbcYjo3C6dv5ELIdufR5jp
QBPpDIPU/XgsKvz/54y8+gx6HBhBb4yvgJeaecd+Cb5g4Xou+Z/S7TD2L2F/BYaH
BcueQQLm1ciAA+eyeIVpwB7AaMm/WAo8JqQA299ZgPR9tgzzLBrmKjkyOgGcVfOf
1ievEvfibK/L5kIWuBrCnQY4RkdmskTHxEM+uJXmm3pvK31cEd1GNbO7/luk90WY
0WjkIMeHUCNOEOOUcPHUjZ5wNmktqNidmO8fL3ZHj0EPJ2Znu2wUYbqBWp5qK+OF
1eVnu9OPScq5cukat3bKJAvnWoi4eVGKp00L9tgkELCDCGkcwbEJWLo9spEucL6R
53bsZLRSzaJpYt5sy8B8P5kPsgO8SRd4X1b6cHK4ZYMIb+2tGKStAJKecgCwx/8z
tCFab6M+4XDQMaKtflIp/36WTdN5v2KAIavIRy5DgYBzKKyK1UutzccVCI9OzhLJ
JvQV4WN2zBAugJEeThAL1KbX64yYds6NZjyrnhC2zIwPVnwLzyi1Y5gwaBiNVPjY
wa7mmY5z/bcgO3Vgfp8BIaEVeHXFoUJZ1/bkmVFpbnOiYKFJLPvyuhh/9CLrken1
cXchgatnh66ECQsuJpw2qILwTErxCfqnHGCQ6BxLw2YMsfpaVxOBiHUrhVy6pG8R
rjOEhywIxXWoIXY5F7Rd3fnm+5i4ZmG/OMuziuvDfe33h4pqkE+DHjWpE4blg6MT
2FSg2YoePIShSSnPSSOLhwGDypFTKmIn6GM8bPanfJiQSIgBDz7bQqBMp8ZLIqAZ
USX2f+mMLpgwrkYMZ2lZjUysGh9IBAcrgoYDjtXf3/R4seH7u6UA3yEJ+YIMU6AQ
NGWAVawf5dpCRzMaVXfcDw3IfDMMCv16HSitbZOtjl10piQ4UGzdPt1fpoG43BTZ
nIFkPXOhMfGDWip4jeOZWcVOI4ZmnvEszGbOOAGrVU5V0WfUNQ6BHUcgerL+CoE7
HvPBG2nPucAvaWd3lVcoEvFkAabQmYgewK9fgYGzsPaYRxECmkAckaZ5+tgcsLpR
m7pgYEhIjw+sC2XJmgFhP/xIX55trPyFj1SLsAYJfEgbH1IkinMlc4wiljdTviGQ
EhZpV9Kcqgbu8JZiKVUut1DsuCuH9ycwCN1OG+Xtw2rIBYNGHGjZm+8PVyn2aXUw
KepJZ+SDhhJYiCeeTi+MKbpi5WoenHX0wXvYqyJWO/1HTMyZWTDB9WrF88Sdumfz
HTAgf/vy30BwBfx6UAE2E386ZE01Zb6qaCr91MzBPThiHrvY3u/FsLyIPlKAKNx4
NNcDIHl885F1KjbC0fwL5DZEFvwSMvaVM0TU3uDe70C9U/lzDvSnq9NXpZWryYCX
02lIwRwEQDSt3Kc261G2cyXKxGNiI98HEmqdtAFybVLhEBsV5N1V53KCdJvHaCdI
bId6UP+stqWyspZpj/eDqcbfygzH8NqfzvJVSC9TOF0TuWbeCnZbAQLD0jDltQyJ
tK+QXknpwMYRbpB0RKNQpc6zRthxTMsBWeKlhIWq3G2k8HtCGGjkMrT5Bs7tr+0V
ePJgOFPwzM7OIgCWHlAI+7HWwxWHQNCADzION6hQJ2zuagj8jac5kV1v0CZs8E1s
jp89MhPDZ+fc8lvtpI1Du+Pnejgz+8MtpYu2DXKCJR0AYznNsr+QCHXgm6qCNa3R
Xb25+U7e7GfwA7bBtNbhZggUUppktKIoAx79OoyPCojGqqNJ51WwEY9rHKXjW6Ze
/vD6JPN+JFcEDrly2pYPutVLWkadfUkpMybWv9TLFQcbnVV3DbkytR8CcLDn1ssT
9VcK7TWy3T8Ew9m6kQae2Dx9N72VD/PyKeXbfTQpsI8f2tLGPF5avIukxsxY7xkq
AWGNSyYPlCPcgU7OxJrhygM26VocVJ/gTMgK9TyDAf46Lfr2u95SiJ8Fnsqnmf7T
vm0gNpzmLFXs0/yaUyj2MdB1Lb4K3CiaqgUz9XeIw3nXo9S4lcVLEF8cDOThaBGq
g+PQi6E02BRAcxsq7IOMS5FvL2g9A2D8G8pp19Stn2gVfJlacOPt0GnRkuFUOGav
xQ/CCbcn0HEOsY5GtXG9tj3TYH43j7slIqZY7TWo2NvDqF1oRHWIxHs4Oy2verEK
3bNOVqYDYu9BIVHDvgh1g5fzp1/PCLVRptCRuTEM7g4Ataee5cTFGnDQZIpUUPmB
sxydVbi3v7ma81FUpdt1tVQ4Q2GDPxf7fdZVoHqDoV17uAlnndjSTX3p0FGO4XWT
zn6u8md1ZGkGP7Q2KDFcDtMFt523ErD4kV70O9w6nLUInCkU/8whaGY8e962DY/l
sSsvfvednbTkzJbBSd3Nn0FD0WMn+vD3wmH5o6OWOmPyAfNzbZn2Krcsbgnr4P3e
SvTQ+TYYBvO9MADyEDgsNumKdGnlgSy9FBnAUZudzBz+a/mKtwDqcYDWz09IB4tg
uOV+ocXXxTombTRnl9KHup7he8y3fWcPqCecNabDOp7/erkJYdj4rkEdWJ2y320c
rGJv0Zss7wxl8PQtHkK95ApYaMfoSESMoWMSY5JpUWTBMIg9w2FXdaqCGjbHu6GA
sxk1ltzKSC3sZzeW7tMdLiI1tL8bvRwwklirmNFZtJXWPdWw7TfThptFGq2exxh+
CrcizOyUeL/PLOv14RgeBVxB7x8arG8n0L/I1HcQL3xERdpBGYY9tdRYjQxAi6Br
sSYjYagclIcWfYO7oCab5TyYc783IblJ5H16gNfw83PXce4USUonwvrIYDXaQ//A
Wc7xU1/jV9XvRR85JmnnsSJC103LAg5cEwf+50FCkp475joGArkF77VMhXbVyjRm
Kx8HMlWZm6KTv/APWXrCMtTKaVb0wWhDGU2Kt/QwQX85sYE3wiY5Jy5nrmJYIvdb
syEKRTChAGSwdscf2d2p2lGgGxY2QLh8ZRA67VpCNNUU9JlHtaOuDWpz31nVUXJW
159sxKcNtrlvEJfBE+6uPaV/w9ed7SkiXjvpqyZDQRbm1ipa7ZN6uNg+yyVM3R5Q
ejXbxntz+Kut4duYUmUcPyMtRg7oJCB7k++WGnl6KPbLRou1MfE3+Bn55xnWpisz
jm4eFN3d6JadhliizkoRs2uefPmJg2c5UlfKYnrkFrJ7rHRJiDcPRhfslrji5z3x
VeCuc7GhqAQi8vX6o1AmPX7bUp2qykvj5qSPBznO514/ni3AkdJeNbm6uOvEsVeA
/gnTLqcdoac1qp7HnxndmvBhZWCw/RShOsvLDsUsi3duCQQgHkCvklcNECM1U0+5
nFzxnWUSGP8vtEqNfvKKQZqYqaSe2S0O7RfQ8oUStcUFm20ec/P3zgowXMn/mEjq
WVFfxIQRoTEbzBSwVEUxeZdE8cy/hqdyZKoEOBtr+Fc9olzzlGj9J5I2T2bqcDlx
Ehj5zU24Hwx/bBDlElDVYyvWJiz1MevNGyvGNM0OxaL0xcsALqc+qo9LicJHMmiC
vPv0k+Arbp3L/KzJrBJiQfMYcjDaTaaDcFwj36BA1f7RwR3ONrGTf/Y4oZ74fUcx
6g7FQzw135VePxQC4FhwHBGSHTlTXGHppGm9yS5M82/z7HYPO1pLPy3aNTNe/Y7M
yIpEXp1mH3B1kBEEp1L2xmvF8XUyawScq19HbvaURnOQ4LPCFRMN0Q5J7ma8XTpx
wl3BVu+BWwPLHfYi6nJ6/YIP5OEEth8I1PwcptM1W6SOZXvUPmb1lmdU6pq5nC2D
24STyUxssGxbMQI9Uhm3YNieQK7456m83UJaMBUBWyf4JiSRaD5pvlXJi6Z91oMi
GHICoi5tXB6k5YTvWpZjIC4NPifdcH8qTGnzJfEnoWS/83ziybMaSOa6f95PBpyz
PHKre1s9h+3Bft+DQ5VxDnPgqPAWVefKNphYoNYsnzyBGXCFMCZyyj7cLo9yKJQv
MDnF5zAAvXiOwmPrNuUc7Sru++UZge2UPF1+5gfYFB3MxAbE3g4DomJlHzGYMEL0
OjzfmuwF+MIF2RXCiV3PNVDMPAZAIWywk8JMWN65z+B4d2gMmF1kzAsJLJ2olxIc
8sk5X7bVsm9drBNJAnKTgj/snw0cTBGqYSqRcVprAAd5ZC2nB34xfaL65Gtm6hnY
4AY/5fQ+SXHXxDq8X6ii1lowhFC4nPN03jLYsgY+GMR9rps4N5eB4oC9zcUU/wX1
gmWU/tuHF0ZJXRUCrc42D1DSKvqzEEQfkFM4o12LaVWiVixB/ahqfK7hPnRqyAAw
92AbkgeI+Y81/iWTEnzVXhiVAjLQGX+McaZbihdsYhjkGe0+i/pQkh9WAQeLb4AF
PTJFJtnDDowuk2bKdIa6/74untnWV/W+5Zw2oHJzVXOqGwSzqiQ3j1xrCSbiI/ip
3Zjs/qOk9GMi+hVCv+XzSXwxHvVMeO8G8VyqzhrtfDa8FoGItxWHSQFTY7I6JdYy
d3jc1GMwIkHSxNn/AZPH3ek3DFuF0fj8VfteabshMAyglIWcXX07JzKGa0hRUPDx
LhoNEDbTsFhWlqPMzgw24q5fM8aOQG7NG6NGOfq56Hm6pdDgw2rMj+g61Yi3kzgH
ALsBXkWG2F/5sgkr2IvKV352Xm1TbSycfMp43tg3bo+2EqhHo2japM4j3P19x5/P
68fhgODNoQxPgmZOg7tSlFMemOH35pX6g+i/Wji+r8BPvMiK/aCqKBPUT16QfQyU
s91g3vlOu/BlhCLZWcyqiWx349suG4RjVoW4cKrm8WyR3HMbzrFhDVxyVpynhp2m
pwgQ0Kev++3tFzjMeyHza43m1nsGKhjbeRqKPlLZCWsWEr+vkqt47gHJIYD+eNSQ
Oh8E6N9w9Xqq3H9Cduk7njpz1MDOabaUIdGXdT4mn0yDxYtUna+DrLTejJqw32tV
EEgc04S3SHKBX73T1OqMDR084Rt5wVmvMA52UC/5o74YtEsZp2YCgNktRtCu0eoN
80wdmYmCckRGXj/SUhojX+Ojd8ZeTaGpcJwplIaMTjpgtxf12kRR4nnsO90O75S2
xTU/9I2DGXAPXVS+Icwhop2vGciP2OP/IQUTHV71+zX7JcJNalC0U/n2DSRBFGzD
6ZXdkx3/H9O6vb1MDNbjnb4Vs75tu30pPMbVzTxDDDoFZ2cMYjUJ81Pbr6naWcdN
Xn7eruXxWeYLb8nJlC/fXoBLp+jq1VfqTq9had+y4lNMTdrHe5hTy5peapr1E8xy
ff5M2piaIDyGhObb1Z/fJ7Uuhv5ltHhoUXH+Y1mZ+v5CbChRWT/is4tUHzCfBoxe
jMoZ6h9SC6zV213lx/JbOCGNg3IJIsq1KeqBWjSDamfmd+m88O7RkgHWz1yrHhgn
0fjOiUK1zOR45oo0Q8Dz0XcuhA141XIUf/KtP+JK1GbE0uWBI0iZNCjAKIbX8OXj
SDkC+C/FfzcMOv4XTiDuqhUSmnrpHOJjeNhbuaiaLLtjmrqAB53Ojlqzwa8IPbfG
KCIo+0Us4BPvCFihLO8YlaadbumepnIGQ4XkhDow69eKvEqPmWPwQ8X/cSXbIOES
GVz6iE8mITZqIogRR+2VOHNdfEBIy697rYdLZyR1po6iHU75/3+mLb7lBPjie+Z9
4V4mZinz3p0Vr9TmHrqxzaX8aRLEIC8dcwLBBEh2SHlG/x5JNt/8Z7+EtMTIee5w
xRS4vDUV9dXAhP6YRZIPXTTo+T8J+BTVJqvoP6hNAsqg14JzhkCSy/kohzfwLhCJ
epohmdnAUp4n/l0EqogJwxSNX5+93ivHtg+QnjOs/dCfXff+VElzN864GSLGGbE7
WQLEVW7DuOb7N3IerAtYdbOkI6pKI4T+TjdKOPp7UHJgiozr3qgQn6K9Q7RoMPEy
H6IO/KWPUBIeX6stoQUwZR0EBVxxgOb5ag7OrH0CgzugQBaHR20LurCBa2XWhjBW
uBAY3FVNkBmoYAO1XzSEI3Nmv/LtNlK1zJb2U78A7WTq0ZlABwl0sPPmV7dQKFae
VAbupe9FECWtPrEvaSU1k4dtGVpB7QQxnecgY5lFXvgsIOtuxGTCCiTdw/wtGpvX
oBeLUIVuKg9JrdNBxfaLFbSYB452LhQCVcZ/VfHaNUD62QnyCcQn/+VajDavUFV6
AS/sjHEWY7J3FK0wjVhVKNOXpNzaD8QNRQWvbamiC766YYPU3Gt1jAVa4mo2smMH
2PIXkTU/LZovDTEH5OVz7M2Wrzpejq2KeE1LWaSKWxa0SWXGFVOXF4l6WDoghfzO
0mIewqk2mqt/1Am8uhwhGhepL5B74NqfvNbQGB6k5Mh1+LZzuHcDS3pkDTBbbwGw
xIPHGxZ/HaVJddVioZ5nO3fxeuqaZputdH7G6Vm0HXPPz2cp7l6UmttShwf8j5f4
0s/EZ4e32V3n6HfLBWylDEqK6uLu7M3qwGXtUP40saFCWx3Ri+GG5H4hBoo9VygP
+Ce150juKvjJOsLH05OngFmFg7SsQFlmIbQkeDmWXo4sGHH3iyOyq2txPWpNgRgZ
Y3fiLerKTR5+vGxYH7fmz1HWVHXtqu+jyjv5zHXpXEVllo1yMtA7FpiMPmj4zt+x
Ty92Qnd5i3fVAlhfpPztjI+fi1KRdGurEDQdVOT0ruthOUQbd+1Wiumd0vIz4Za7
zCDO8SLi5FZdDwAAaMLfEOOgflLqlrlVif21Js5BXD5C1f2BWrICXC0f/liQxCn5
g3LVYmOZn60dcCnNbYhFOxtzMxf+iZS5+OU0/i54vIhzi/l6xg97X1PET+2047Ya
dQNc1BK91B2ryYAjj2VpSnjGGtht0ddj0NWpDNg26nJPw/TAt1rl1TrQbTYo4zaf
rIKYJqNbvEOKNu6CVeSQhhejl/3WGSHKWGsh9FtVG3S33exRD3SuMTPqCXFb0VjB
JuesYGpeDB61vMAasyil3Hl4qgaEdwdRSFvw8DSJ1wLrUvOvIxZCDRUFGxFylUs8
9amf+7ojRsynsTODSUeMtn8RllhmMMdRpfOyjCHw01f26fsB9Ugza4a4K/DpwUsn
RaUG0aDWni42pGPmnz5IDPNzTREmLOBhz4Izzq/AADl799Iq0jPFmirvA4QIdtqf
hY0iG/eTxMSltC5VUwKhlJArDwzxeMkElKfEt4ZIFjtbauSDyzdDRlv6sBiyjSPG
L0AgwK8rI0zfuu1/xOTDxEXg9kbbKbxws0x39dTb34j5mjwM6GASDUnlsrru/rpO
4cKN96iNS/AIgLxFekFQfdts/xpRM2TtDmfkxpyF9QOMjirct+7Z08ePCieDBklH
dGfjY8ncp2+QfzLX+ijF1FZE5JiaeawC6jAYgE4Ic3b7rApAESu8Fz0WhKxFj084
YSup9j2z0dOoNOPMEAroE+Z50XDuHX311DSExTfcSZZoqFIBQs1v00QZREUfhtaZ
dlB+OzsPKZFSFLfZPkuiUJCnU/qwcPh5c+XRpnlCu6LJCpt6znRc1xQC3KE8nRpk
0nZpgUJNPS26WQem7PvbcOPQe9/va0KxcHgh4DrC+Y2syQxvQicA6695Co3V+nr3
VnSyXXZ1OyqXwH3RZugSKMWD8CEjfromCGxcmA89WItegMOjuRrGQEk8M1+YcZyj
42zV++UZTa782aQYIAs4EB/RxKBPeZDZ8TsqLMBljIWyOkzQD5UEEy++ls8rEM/s
BpAbPOmL+DCRfdMnvV7OB9Co6fdRZBY8Tnr6MYFz0ruDmPEBEerDDknFsbtryikl
f+T9nJd6d+Z3MfrjQbOHnbQyb6QQlxCmXnmQ5sAj4bxrPp19xPOkWhloz0QE0LUt
Zf9Y5Bg/OBjpD/jQ+/JhNlD1xRSZUAFPxnTlKHDehSoDzdaDlbEeM1/nxbK6KoTb
WLaKZOf6kjuqiXQPXTgmtVMwNZycrY3qcTCWur899/cfuDsULgRGg+oRGzSjDtye
r3fD+QQq22e5mBuKC4dUtioVHgLPhHitrrh6q0hY7mXHFNydxZlM6twQ0onAbMhO
DGesDTYKH01sEAENPUPCHwGqrRSkWQk9szzelfVBvZSse94JCFeOWXypYwcasn7p
koPrTc/UWT2/Pfym6sB+YxmojCU+SVx/IDFtj0TYSIE8sQUUrUvR55dq7kScziv3
lb5qIsn2n/gkbcis9iCk0kh0qmtQbPpwVZxfcTWwnp6edef5KZW77bB5hNpZOuXW
8o17M/IpsotB+S2uzExKmhCMbqVRzd2eCK+Bl0/S2ld38sgM5FyiNuZJKXNqKq0I
SOQGJYhtNMMR5G4hNjjhSf1WR0ARFvD5rQ4lJSQS2q3D1jcaRkqBM+vwrBCixmcp
XNmJ00Et9qvJ5kS942GAh6kUmuF4tS5Ow4JLkhyYmlCvnGXJAz+izlPK8AHJ0GJ8
60vW0krz7ye8CVmToaZG1Lwyw9JdxRR/qoaZ0/w3gPFYq4aoUP8zZkn6u1THnYLM
ZWzj0+J7P71ZAWAy2XUP9fNi9CRGVebHFqthX59olUGqmSl/w1bzmvgHYEIvz3GE
7hxyFPh6kkPriVyvxLM6uOUczxA22gIB4NzFCUHORd6rp8IkVsL1DsgnCFCo8vhn
kgzY7UsvUg+HbVFlfl0LCmo+W+KhO5VuBwtjxbbume6gTZeQUdTlZHaIVS0sGSOl
L8iTWexv/exCwjBlOb7A2hGyoK6tkFmvT7JRz9aCleqrPa4icmmFtEWdS7ulakBD
muB7M5qSVRC2xofjfaTnAoEBfCcIvLsAw7X6QLA24QPJnwB2AUO401gmDoRqbkiD
xg5pt2uMdtn+g+ZfQlL8wqd+P0uyG4YqsvGGdCr/ZjkD4HoMiVABsa2RfXPIInjZ
2WdreHYtx9Gq45d10x/C+wtM9QfuSktIv4IRZ5nM8bMGjsdccNkkTbqGV/TRBjft
3cX3j91XHP+MoedwB1g91oas2xJc9HslqxqLVKqWvbUqqa0Q2joUaWEa0LqMqWE6
UpzaMdysNSe/nVzEurCqFiMylQIU6laJ1HV0ttGeJ2wnBhgnjsE8SckBu0WX6k2R
BVf3whz6hotnxQAkAPbrm684MkjNKafpYjnoDxt/v6XNKv4jvOzMJv6/vg6+fHno
D0kz3C+6/6N7aKIeyCXHrNwhAh/fvfLdrp0oYXKhMREK20eTSiD7FPDJmCqd+i/b
XUJNsPqcMY/XcWMDlimVr1fB/wQ0NKeoMN6roh6/sfAI3kncSQDq6FhcI5HfkKmg
q4VO0Ha80Fr2TmIGdN9nCv/pAfYdX7Sdw8DaMRETJl7DHM+ojnBAGdMy0CfRxy46
c8jiKW7dNJZRDWxAKm28/xl8Ul3gFCqn2NX1yIajJrI=
`protect END_PROTECTED
