`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C5XDpzYbJbzL21U7mM8bLALLkFFY4EupAwvy9WsRB4Dnm0XmXnQLiVqQELQ660ft
wt6olTvgpViWePwTNcUi8oI3p6Aq3t0PpPrsF/Kbls/1rp9nrPNVXPdPSoW3qbNb
+wH58kEc7WlEkFwEPHt8VRqVaQfEb7TFoWHveuQTsSmxoCIBTfG2rDwE8rHSFr/L
CRlzaYtonZowqywMjSAeJCSjw1Lq867sO1m7BBYqee674uCG2YNDZXSkXvbkshl9
kV/m9IbiSsHJ5w9SxE7bj+INVMZ9rf/MBnsr2oECut/D954ykIrIzVEXcNwELoMe
aVkUQic+hc3LUmjqkzZRiQepG2DN9/bc9b+88QCPbNDEM+nIS2M62ekKWGJ3oreG
fvQC16E8gSDGUymz6tzXXQ==
`protect END_PROTECTED
