`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NH2mSUsqQm191svgSjjqgWh7B54V2GIRWwFTKzRhoUUu5lVnkBXRG8KnvRQCZB1Z
Qa40Kr72NoHe3pSrpiWJDtQiw4QIcELy4IRjX2vXBOzu08IuCa2dUWepHg3Llykr
nBIquWfU3gCTwgMlmTf35VlAw1N4EYdte4E4oDJvXuATYVSzage/yU4Y+C+5H4I1
MopcrBh54ISxNVwZZV1BkD3ZWqXS7wWx4uRr8u0xF5ZdIQJgMvdmStgFNtRkKlJy
g2jjKURwq2kWmhzZK6c+YSSz5uxeqcKAosSfrjZ07HZV4Hw8O1r6Z1JayI82DJ5p
xoAFG6woLw4e/mqeGzDvv6N2Js8YiqZoII4EUAl1Hz9MN4SsX9C3elVkiO10E2+u
uJBwi+Oyg2nI9IionSrvccCgGwCz9wgJTGAjfvs1NucOCZb3wGY1rIVyqSnvKQt0
QU66NAn7K6f7EnyUpMDKV/+bmnPzBzHzyPYBOBMjlRoXb47eKJWnWVDLzrt7ZYZf
F6u7B7JpFMtvTlmNnoB+gtd8t0h61J2vYxJjZLPQ9mNJXQAr2apLrY3kDf/liVLF
0B+Yaqgyq15YwNH1bd+HX4JBIvoxE9ploSKOYTA27i6aQiBYxqc2wfehJzx49Ckp
OsyJxaYAA1jj4rnCK2iowNvBOeFCgLi0OuQZu3fhhtFChmE6fbQaF/OIWqxk7vMZ
Vq6Betd6eL4i4UWLMMhIYiNfX0iNmZ0s9tgDHheRrvrNa5hLJKhF6uyiIm9K4SH8
HNljNwfT63a3TQ8cH0vwftsEUxwEDQiYNq/yShVL/UiIVvTEW3Ql1hifUkcXF2Pv
nmietDjKhqS7Y6SFtHCIZ9H4Jn5xL1k9oCC0KoOTYQspF5GOlX+Y3Kqk+YqQX7Wo
xA+gQjkHGNQ49CbtUSi8OHlXWlLox449x0gRjOkRTi3mqqLNlWchrff9SASClNFa
`protect END_PROTECTED
