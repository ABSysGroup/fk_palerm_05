`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zC2XSe1ozvRF79l7sDkKfOE7aAUFbq06c8J1aEQlwttW/vJSTwcNeVU7cWFEFShs
C6rSaZRj4btKLlmrSI69ZyeOcivbSYCVTdfezkpT3cCYD1e+kbkWyr9uleS3tH17
WmNnBrmvZ3P1VUDW4+U9FD74LRgCV1cUru1NEi2K+EeRjrfDrZpwP+UwkYDuZpNq
HLS5afGRUkt4JrDO/wPXE5v1X9iC3PbhMVl8ywVM/WJXP0W2ZDqh9CuxCv3uWH0E
BqVmIelDEp3E7vAaNE55ntJnT1ok5Y5Uqm7WxhRtRYeXOkbFuiaKevMs2yUE3B68
BgJ+gfnDHDkLKTBmRLqMmRe8yApwvkPKaD4v2ahhooTrhoAal2MFyaXtpmS11Ywc
Mh/ysKgWq+LuIKtzdlQRlbEpulDmRDmnNykU41SUScW4tXtuKlGFuTbxMS/Sv1b2
nykL/KhHr4Aip1cN6pm+m4fQGbO3z+fChzQMs1C9Bn3tRLffKxiWF9IgXJ4ajXcm
IAohx6JekmOHgzy6SGa63ilwPwL7Cwx0Z8S1eClUXJMBG4etbrcRpVmP6ptZdU07
VW08aA2Iu0757cwSt7Fckbib6ewwxOmDiaMg0AseMiA2GC7CzwKZVrSeAladK/kf
RZUzK7EtOirvXZMZSUV7P+79TlMUvYYEnF+n6dTjHE7I3tOSoz57PUgxsiP6cjzX
sIP8H7q10BW7UIE06ukTYcAmOY0wUk5EIAGu0qddaEj824mHe523NyM6R7ABjpxD
SIpiCy3vCenLvefcKfwR3bS5o0vKjWihMn0fD7lU2MvNhxhv5Rt0VbJt2fimrIsL
3Ipy+0UBjd3WWWh+t8yTZv/o27ThgdNVnbnxRG7q+mtEOJ7RtPUUHjQPGF8WGGxA
QjVxd52ncB9g1QuPLsIGkBR+n4+vigGKphGn2+YzbGEFy7xC2v5d1IacVXb1aoA+
AXPWoKJ/gdIlC/CBdgZ2FQKDVxDF6hzTJd6pYYBfLNNV65GyYjjfsuq/AYEF3IVl
9Dhla1QHtz6HiUk20ZYrCiEqQEUcLTfj2LCtEcXwxrY8nn6Q/EtBxQFc9Vu0UA+l
HhImkOCbSnKgf7L3ZGmYCcMg0Sye0k8srF5ry5NN4SybyVuW6i1D/ztIbaYB756W
FKMtSwqZhjgctkjPm8u2zs/09D4i1b8lrxw+h17wMNVGGQG3laMqTgbsmylSdlcp
cfGGL1d7Cp1UjpR8Gscq6+Lp1WXhQ0NQrvjJgaPMX8BWNX9rE1rUJ7PTXo4QGzCO
urf4u+6GjW1trKDV8lO2HBvSgmbGea07t1oxQhhnueEkm4lQT4tPwczx5SVwJgQ9
KlbQ7PkT9EbqMPxO8Gx5zL/5FQ7ouVt9fpy3aZ3jcFTOW2a4KVT1FXplKSAblAK4
gxtvkfWTgryDatFOuqjVq7jG3g4hnz2WmZjvaztRqWR6valxq3NRt6HHPcJmLFNp
yQPiCg1Oitm+IT2h49F2pqPS1AGaWMxr63QDGpKvza/6ReOg+XWNpDjeUpBwDdX+
`protect END_PROTECTED
