`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nGhf1FqOc+IpRRpHtXld7AolGJXlBhrpqF7irvJNT21yK2MhO+BX08RVxUGSge9Z
18mCQRTct+zUHyb8SyrUKCUHb4+UX6+6lVOzzPcS0IyLtoZwCLr3bKsiVJSPpb7o
bCQDNhX9FWwbRlY4P+Pf1OwXpwDuJgXZ7m4OqdEkUAaJLMUy8uM6iacqRtVgx2kG
n1HTXHcSnqbG+91xsxb+yJtEcx8XbLcFNd2LeOHGabd+EXJ9YAqDkZD/4lDRwV7u
2XDznjh4BlFsOXicmg3o4g==
`protect END_PROTECTED
