`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rJZrqDx8LuXTXC23VCLVve0YVxNlCtd2A3Kb/WRHobq0fkMLHdxwzBz+JgPEtfjj
CmjnmB6hZ4LBJBWTodRRqtyj80Ghd3qFJNSmXsOdlHOSl2loV2s0Yp2uHDTM3S6e
mPlvA8I4Fl9BDyqEYs0KE5EYdXqnb6YO3fdhw+mhuEc0m0BuH0AuyFZj7F9fNa7z
KsPhysem3O+dc2OYrKtTTW1VfgeyLzcM8KEuRAYSqWZFBuVBus4KieayIACCdYHy
dCzqk53P51pCmhHk9a5/z8Lomp62jpVukIK6U3UtZBeIpedB4nS5tWNUiEb5D/yq
GCg+SP5+TGfsdbw523+GcWlWGTFfFCzzdPOABIeJ7IttoYiamF/9g/bIBdWuAC+T
paYRbwCJvL+u01wCxRfCMf2KlEYuIVXkOd1M0T8Ry71UW3I0hixfwKogxBczvLVX
Vl8xRVMjQFF36pWXGffXF8bzYzE0jJtnQD6caEmdrhswAVv1oxBCW/tn27aEmmfN
BW50UsagF5zk4TQEuAteWMhBUYwakDpb35c5V+7X4nTfWEe6IzJYMnHwqmRmsSQn
HOYETeuKXX7aO8OlU9hHmTngbSzHXtFTM/BHE5KA8TN+R/e2/rJ4qb8aYm4+HJqQ
NchqeY7p+8/vkqWcoN/ZJPX5Z+D583gWzbfS1Wnzq587Zj7yOh9KSRso/q6OpVbn
Di5Kc94ceZaIZ8TrGg/c5FbXFZstxl40NX7qD43cRKg3obBaj7ShsrXgZAAofm/H
6VnbaBicjyxzgM1+Q6KGdXjheS3sjO5ZCwFleUe2qG/0h4yOgGN4d1UIDqAUa0EV
4sWrvJ2TdE7lMRZLASdnjBd6k9hxhxL7B0E75xcuPISi9Zs9xYt3bkswD1KnkeOM
NS9ki1TXMToUaFckeC982g0+rDm/EoxPNR2EIxNO6DI=
`protect END_PROTECTED
