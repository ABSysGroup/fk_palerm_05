`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aeEYg0gMRDggE27/xDOHCyQxsbc1SjLx8d/pYFQV8ObhfjNYs65uXE3iMohzSP2W
tXBRHvJ1pbBj0LhVkKK+kfzA/7C8P4SoJT6GmnvhAZ9z3xQO1iQgFRbev/1wQAB+
orwHadSZu+vknyDvlNPOHjfGjSEz2c5uxLRpW0eQjr4bl/5s0q2g6cE9fFQjtJyX
3VxajcnjMdSmV5EJda+8wLAVvn2XT3nmLJpuZQldk5N41V7EKo37rfK2SGiIpaZ9
EJZokoG7ZCj3T0jpHMLFHnqCLWRmot0k0NvCzIseZWE=
`protect END_PROTECTED
