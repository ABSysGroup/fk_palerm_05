`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NbsznqGKEwZymkR2DeDN6N0xDCI1naxqmJ8wLQTi1RKkBq15/WiFya8yC2+I5hsH
Zqc88hlCNJ2rvFF4eMITU6PgXiROcaB6ggevBMdXEdfkSVNb8JpUqQahP8eo8RWm
9Nx7CnOKh+/PsIcPn5ZrQ6p+qNZZwkU3TpaqVuKh0iUe9ZmA1Mu5aCNJprSYXjg7
wxaoexFuqJ/WKIsO89zXk7BrOy1IL4XrjwHyvejJsmSb6vMxm83lwFZ+lEFBVD68
ndY/TMQl4H0E/giPkZA/mVFiDCjVgf39fDeiqeyGNrzOfedkmY5Not+oB2MyRlV6
1vK4/r/MOIMUMzpm58Dh2zo9svZCcY0r4PJ950AgvktHS86qpoJ4QNtk4mWe6xyt
pBRxIOqdsOXUHg47gSIZIusE9wXL3gsL9vs1mOzb1o4KEwZrPLf/LUTdr8sd1F4V
TANX0kOE/fvb96bNjVLU85t5zwf/QAovNH1bDbLReODp5dUkPnnbpWXyBV2RTTIr
g6K6cLcxlGiSFFOLt1dWsXdWz7WMHVx0K7iAzI9UZBuv4YXOs642rmpxIZbsKU2q
JSRd7mvJ1aqwS3E1n2klSgs/MHgBSNPLJsq+IHuvKdkNFrucktnyrw/EOUThjj5q
PXqnRDu0hsPpaa/weK0yWy5e3J3RGFUvcwDDhKmIZOwrXP3IdmwO578IWtIJCJXt
9650IkNx3XJJ9ZTqH+J6+HZHgGdm+pza4u8p8QxUXcCbkg4/s4FnCqzvhnCfzy8O
Qs5aTBhXeJFIkdZMorde5CSv7XU2qbbJ5pF/HqFbRD4kB2eKNfE/r2BUc2rXRDlJ
ljvq9sVkWckH1zysWq4W/6kWBRzm0uKHKe3yLAb3gx3CAM8NBq4jYdlbQqeIG+pm
HuHIWIaEa6mUo4bK1XzQ/M2gQ+5qAuW5nE+DgzTFMcdUWxUDn7AwNJH5MBam5yCZ
`protect END_PROTECTED
