`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LITkeavHYX9yJAFGnA6rKBNmNcQ+i156utT6jflzzIWnowwnd8kq7mCGKJP8eZ3W
7wdyJ6MHmwIquK+3oLQmXmOxzPDK3+e+sElt6XHxmzyb4KW/JOW36VejcAWe3+Xr
CVhP5ePERVJuhYTBzDhR6o9PFEnMFXvShWsOxYxnm9gWhFB3gCnVDavxkXjTWGwC
4MhJ+k17YtC/F0WZHOTEWrJzZOtv7Jr8SyLf12eODZo47uhqmxX+R6lJ/oV5H+3u
eXpbtODdBi3TGrOf67mdTqCaIEvCOFrXYEynFvKaHCDf8iZGwE1+Et2Kl7K+fn0V
OaFMyIsGomTLzhgchXXcKk7Jm72NGtauIM8j2LnpGsuNNvBDJ38Vn+x9B0p3PH/p
JgRCEEgO3ghpMPc94u1uf3cSoRCbGXC45zatKS7r/52Q3dOeH087MNYYZfFxIMWP
ysoBaCSShmd13vDB8o5zC/aqTt11s4z2zHOhbvicZvnd32zLd3cN3iscyT36ABjf
8Dc2xDIXoPOipIhBw3rV7JawG9fqnxunXpNEuqhfa6nPzglNcPYUh+95vCbg/4ow
+/Oo+i6WafyofIiQ9Yh+hIxPh/FnCOMsahglX7qiN0yEh7T1/Y65eiXuam9PDAAv
pQ8sqa1HMzOT4DlSURtli9sNVd/TVKwOSa6y6oNqdcldegIL2Jp7InLW8B6S+miz
sBSv9DqqsWcPQ0QrXO+NmlG7Kfe5qxKF8nqJQ2yrjPQn6DI7K7VEuDWGyDn3hrBB
7R03O/dMey+14Ud+PYROzDE8kaFEVu60st0VIKXhWz9VPhmSphruyo5y1tpX628/
oaMJ9gSeSJu2ORspfi3/3ELWNxg1hK09oJT5ICzGyxUsMrtxHSjrtLTHY7Xuy7IE
BktPrp67OTC/0B8hHreXrcLDQTN/vpH+MT6cpSHkoNiHfZQEOQumoANHAaNN8+/g
KPE5ja0smmzXMvpKmvU6aCQ/sN0S5vibFePogNcWnwrG3eNCAXeirNdmKQUEUjw7
cHsCieQAoHvGDK/QRCWTqGk6aIOjuIc8gM7vRqoUtipjtah32mIxJJF5dUtmzzkO
LbV9aP4Sa48+S780/fzIc3PomWCTlr8ze3o0KIHw6Uo=
`protect END_PROTECTED
