`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9mskXR4tn76XFV46k1C37/BzpnCQ8wEfbxufMlr2G3tXJT58cIm7iiiU2gkGwJbg
oc9gpQ8wxGP20DDMvOMyiRbhSP/RToDjiR1HOc3am/TxjvW+gTOc8Lh8xN8DW8Nv
BVbk+bCzzcPFwLe0UZS2wdTFoAwyjDn9GEu+3+kkd72K8l52k1FydwYEtVgdaCD/
KCjuZOimKIiaTnAqDfi+gCNH/Jbo2xzy9gvsNJCckWtH8WGkzgv38lc6AHdw3Pwe
mQEU9+TcRl/UUGJGM4Ud3FSiTNKGns9EkT1z9/QbgdimvId+q5+Dg+a0vZJ3WpFi
MuIJzSZ0Im1a7VmrEBX3MISKjHdkHKtgs4+dicFmc7D6eTg5COvDPmE8MVCEaPiR
+QTuSbmOSDouQkiMHS7p5kuS48Clo5aRVISnIq0dytFEQRK0y9Vert0zptCHD4Q6
qNHNZ+SbY0o+3vSaRBYYAw==
`protect END_PROTECTED
