`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sex5zyt+P/dmVyx0/4fKdpOq3xB/JgyiwUB8F2lauKTJrXZlP951CecnLx8ghOQX
KQPKVhL+yJ0ifMA69ftZo4uiVWv2fn5TRlzDWbgplzxORREXMg+Es7mrO7yqlqYa
QnwVvj946/Ral/6vyQN9+K3otdEJ46suy3r55tIX9GnzH6ObC+1c+Id/6vuoBHLj
TS4uyXDSv+hQEhHvlHwjGn9vdO0BJ7BSJZmSzck9Tcpw2BJFRSTF2qC/TcubzpWq
dezw00J/BdTDwZ4tN3LFdeeUIZteWK4bcrggAjqy1ybQWwAWO2WlarGLrDkQVazi
usqSRLbFounGP2o7x2h0/MSteXRicE6jYawgsQ2hjB362+o0U2vg93OJbKGNwI1G
n/8KK8qk5lNasX8uYe32MkGfIYJg5NNDtYiMK0ONk41ZZP3XrVcQKI1iGpTSj3sh
`protect END_PROTECTED
