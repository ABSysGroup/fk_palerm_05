`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tWRPzQR5ZzVfIl0egsRAE2bzA5UKkHo6WN2GlmfUcTCAVPcnngIiCIc5xBkCajmm
vUDnaMcgsHy5/3QhY4ec6mC8w6FBsS2GQZeOGyl0tG7jOKu3ZXHR3qnfpQW2UY4M
FW52fiPMPbEX+zaYgkEz1qmiDiGTKR1fciT29uEUf+09X45ECI9eioAF9oQf/VlR
hgfVd7+AWMKch2V72+dcgzpTIk9q5tOqUyymoxSKYWB0Y/jWMs8SFEzWABU/kzGV
GbnIH03aDEXJIkdxt1g1aBJXDcwJaZlVnp4c8GmIfduz0AtMJ7yKZ3Qo/FmHJrPT
1YuCK3o0I+YdL1vZ2/TRUCa/BVVJlCTxpYwYZcjG/AS4gO5d01erqTpD4YGbMIRT
m5StF3K2RwLK7IX5udYhkGLRQDqhVaPLHmbUN4puC/GE7yE34ApYVi5B7s5qlcW8
z6CIfOg7XJ1TE5yslzJadyMhFeVIAvh68VtZShShfzKiuJbKfH9Cx/1WU6WNK3ny
3WPeTssrX2Nk0xwNwm9O4x92RcP4BYmYXh5oPM5qDE221qdpp7viccC/4TY1aJ1y
+NvyVfNLT1GDlNrcv8SYQok7WvQeTWl8vbUix0/LIRfvaqbTu9NjVIupijJqKD7d
vU8R3RS1RHJBklkXkOx9OA==
`protect END_PROTECTED
