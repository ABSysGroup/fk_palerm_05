`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tDp7h/f8yNzEhtOxyILUSPCMdu/1lT1WGcuHdMd6rjlwTzNPmKVc2OvEiPD5OV8O
U+i6NgEbk1r1qunhq2bvAqEBAQenjDi6zy6TI7TYn99o95YpM48+tNBzwwzVpUpY
a5JnBGfaQSeA6kUHsZBJPQSQlwv0YjC3hf7QXq/qZZvKRpQK4oAvaCabHG48cLoK
anOy9l2a8NXRjaGRIp7sRbEsjBaqyQDuiOdT3T21A3uGjnF9hAmNpJiMzT5FuNdW
kL2IzYv/pbRQvLHax9cb42iGDlGLyqEk9OxVKz/WpSNcXKfJW2eOoKAqdFBEIqIW
BG0YJneToCiT02n3pEmxooEangWlavtKdGE6jlssGEjndBwSFrn26r983sDlBzbK
pe4SuOjAx8dHsAVOnRMnyxLnrOWGU3nvjk6+DSPsePeopCQ2pTwTjSM9bmiTWMpa
`protect END_PROTECTED
