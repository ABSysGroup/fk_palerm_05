`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4wVZzX4sWdNYFTCDBRdVl1gqJhC73uB2R9Q77M0r53ssSg/TnqURTZfYgvJ7bbUG
6fXuh8PFqA6jJb7KqkX+tOGWRI0WKmEvhvH6PLl2Lu8W3Mnwjo+v8DqnzOtawD9i
CjhaGcuXpNKMPJP5kRKIbxDcwVZ1ESdGYea0Pi2/Gbh0lC1Ht3vUH98YmLnXjTKM
ooC+LJSht+b6tNeAQsW+Sgm3NIxabGNgLTn56xgVnQohCp4GhlSZ3wnkQtzDq3m1
0Jtv9oZgd9EX2eDKaEuNfdEpTwmiLxz5U3d2igqz10vyY4MYLWWN+rBQh8mNzYmC
Ei8HHDF18uuTYR9N/Fy0nWjJAlf7ONKBq4CMG0Dy5ywbRJ52rkD/FAI2+nwsrNzs
IcLAA117J7NOgIFVxxjojeEj4J5pEWYL+DD1nK8NHCI0TruLtKsgHRAxxy7DjxJn
yi9QJbmILVDgvEam+DEK4mlcZKfitmAs972L4Xqlbg8G00gPac1aVD6cCNW+NATd
Y8MPnt/FHSvr+AWGVz4Ve1LxmZTGJNnYsfFxekJIBPAuFXiCl0CS0AGovdPIWxyU
MNpoSrzsaYc6Jok+L5tkotzmh/kPCq3x7kl2EjbkIDN5iItnonK1yp9EUTH5R/q2
VBBX1ynamrzEIfEEVAGCQgLzjyT/N6wbjVKGlYLaZYifHXDXyS2ofjto1mkkHjcA
jHhy51MBRQGSoNcucX4SnQrCGWiDQSLRI+71IUZPkOZjo1FujXSrjxggPkGp23Ek
3IpXR+fYemRAAN8olBVhrL9eBSaO6vSHwwG6m9BbY/1O7/n0ca5LilACOCaOvRhH
82zczzQVm+KJD0OBgduzoW9oJHI8xHj4fQkM7ygvddgjYD/i9ibIRG62+JCNaoUD
6Ni3LthO6xcJ9ldnJ/RrPja1nj61YG1C7EHD3EDSDw39ajyPeJhQN5by1qAcvL/P
1XWs6L+R2W/kq6iQlX7ohw5/ZXXA9Hr2txKFLXw2Im0HyJJTN05cYiqHg47tjDFL
7L0y/FxIDoWKHWd80SDXLw4Cc/dDkLoBSqk1RhUFLBJIQJsRmnLekwqslo5fLF4X
WqnOsFJe37QW7eRvFqh2R/Gkj2xJnjgsR6Pd8BV2TNLWMVlkLFcA+HyayRx//swc
yDPuKHon35iAUEJNOT7bb1IysLc3flgD1CC/IECEMeJtejUBFgzaEk03ROjrxYn0
Fuz3Spb6BVHGOL7oEvi7WEYl7lgNV5KgSpC0pIswTsuJ8AwmyUC7Qc2pSQBI8E3q
az6tS65SeQgqZl0hcEyJ7GoJwMyInq4n28/s5I7jfXnClEDAfacoWg57L4wToWyC
JCveTaM9xH75/EbNJTTDYO/rJp9NZcE+3lyoKl7OUcIuVP9SazriQ6/VnvjDBVBN
P3kqL95G+tVXnGwA9/mi1Q==
`protect END_PROTECTED
