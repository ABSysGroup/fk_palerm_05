`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sDYdsIuZRxKZDfRocnjY67njVvM//FYQgpnirsL7FrcKKL6NdpYzynIMIopqlinS
pcRpwbsRJ+6vTxsjOBkwolvoGozdzVN+Xul/yMiN3aglth23AjFn6sRghPECIIjK
iCs1RVAKPOJwiAqdt2BiviLPofk1cZKdPLxcW6IKZCs125uiYlSq3jeRwrqRAhgr
n0HciTJamtPD02ZnR7+V1X6DNgIRc5Oe2kWUJvyTaj+WWpQg41I3smqHk5zzE4Kj
Thj+MFSivj8vvh+Og+iWiIEg5KsY31+uS0IXN9tDYn0n1Tfm6LnQLbj/ZkaNG3Hf
QxhLKgxRsebmfffQ0HTmjQ==
`protect END_PROTECTED
