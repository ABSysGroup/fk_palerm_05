`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
07CToq7CBa3G3TWfJccHdHleHzZt+rnMwrcuvclHdaLEuTD1iyY7rlyIcfFYbqim
lLRBGEB6rdyI+JuLRMyXLSz/ozom0xG/swxWd29UfB/ss8m2sA8gMJO8riM/rT9z
cZCtBlBNadfKTxXrB73TtgFq1q6ULuxE4WXWZmwDQsMi13qp2oYxaVK3Ls2RhaQd
+3Kj0JbNowIBvGiTjS7wO/RQGEPqQPpzuq1CDUdQjuf7tE/d0ur/1HxvyQc2mmKD
904Jg7sKktLUrEPsCfyjyAqIRoTH2tItDrdmBRCjZwGZcqekJUHo67LjZ0tG3pIr
Bunp6ngJanNhnV+hP+TUtbEus0/Sh/Vq1AxRWr5zzZ2W7BfMTPPmfFenZXOGo+Lp
8pqLx3OoRtijGs89Lu65sCsurEE42gL3VnpLHJaMGaYFCSQviWodymGA0kkWYx5s
86pKHBiz5vipzJ0YnSTBJQ==
`protect END_PROTECTED
