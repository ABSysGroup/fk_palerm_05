`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4DGVb90F4P/JideZqBm55+6fNEp7B1UnkFE7UwExSg+OyX2QMSCpQwS3rxFta5+q
qbFKdi1oq97gNTBjy4nFaj2jwJ8K+L9V+k/iWNs3JS5DwIfRK5E1s/VUXEgAqdSi
I2KDQoSrCFwnRftYDRspkWtij6O07VXOaHUPr+RXYT0VU8yhJJvvJm3QzJkRt3kk
bJ+HRzeyqfJHLXnY++1odZt8w8d8et8fzXYo6bqMEQzbpC5xseTQ/b6ijD7Zm1yK
Nb6CuFLMmFa+iM7OfEBxO9YSvf7jTxuag/tQ6Uz+AtzhejMwdhR5mRxkdCKreMvk
64s34dtCB+EkDlrzOdxisw==
`protect END_PROTECTED
