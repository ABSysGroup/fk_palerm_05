`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1aR+F2NFGI6AAFBjaU7dWW+oMhHIGQPtgC+KgTtDueQI2Nw5cd7i1qDzBrfXLKle
SLmJGXwVTaNK6FjMr3KetR2zi0a/AdmYwn1ZVUyeXeKhYrK+wiwcC7wV8sKTm7Qb
S3n0fQYOpFTQDT9HTVbquByWqCpW98gIXV7tsmMas1F15f332OivmoSMzb118iW0
jjAKQYyCgBE8QTCrcCoQlrlN7tAewL95+aRDGbwYohabw0cg3dPNygFL2XNu50fH
BjHEaPrww3uMwSuG0ImmEmwvEIX4iKK8ljVP9a0zqaryi0T6umI0xtqLTuGWKFYx
ssXmwUL6wp5c5z6F4RsJEy9SBMHughPSe4iJdM6dq+4eedVyYKqESFIAF5txnTQA
druqmFSR3V8teFeHCh4QFm6vMZbPbXMDGP0TP/5XSizTQmXCrztcitclhvzrFfAl
KnG/UwNcGDmWjktZVNYlOLkbO7bgOapc3HVoz4WnkI3DJSdvNT+Zof6TGosFt4OG
oQ2jvnnGmJft9AQ2ZTiMP8XBbS842iZhV3VfHnbpI10oiBGjuMOE+E/a9XP+QYux
pMZigzIS/lgC9mH9PEAwo8AZsZp/XL3S/JvNYc4OlOzYVZ1UvJdFhTaWaLqSp368
RNNl/iyaWORt9alW/NUCLFnKyCC8+S4+tFvSGA+e3qDgdstLEjSw1v2JjClLyLHQ
s4INYf9mZkfTs/Dts+YrHg==
`protect END_PROTECTED
