`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dKqpNN6ue6dFAUH0+jVAbY7UYMTcpmtmnecb4Uj7uZw6J6BzRw9+zRK/4zCuR/e4
xbh3nZlj9AAXBYhxuORY9WGNvdD2ixWEdMhGxRGSgEMAhH/Y/bISOF6btHjGW/4d
X9PExgnfajQ+MO4zwJyzqugIiE6poeaCXIs6HCUjs88VUWzrSOshgNibc5yudlsS
3GUdZCESx8X7PnKxfvvfZRjuCyBZ8XmgRLTSIzI7jSaQL/QYK/gMaj+ziEPpt0Hk
nBusXOoheJ0Ur7wDSruID3a+WM0HGpFKZljPK2MJSbrqa81e3entC5ik9dwqfHKB
XGE1Hd/mF1VeImj5K96UU5Zjq7fAtXrYBwvsZdGF1CSArdnNcrvyYiuzRg1UFTSm
WbB9F5U51pRPaVfqR6Of7HW/54Oi6leuRGzoB89AgNinwBn6BMcINy1mu/z3BEV4
zRsiJZ4Q3yEHAUYL5tr6BhurK2+JpjpEuyeO7/EE3QLBLq2wMQefKR+18NlDXPFS
18IqQlxaDQEGcgweXH2sh1KpNS/oZf2J6Bnrqaw5t74f7apUm/7rec2wvoZVQMHC
Flks8fLpVYTzhCvzIUtScRjGWDfHQK8AYPOKIKKjV7eiS2HI73Jt4LJQlxqa5lyK
XMEHes1hOnUimgqg/xEL9pHVToTGDy7LvYkXGyNVmpaABtnqXJi2p82KmY6BHyjB
x3OQXKtQNj8UritydqMinTZqYzS+BXnOJB9ezuheTq5y4WLTC564QJnERtPlLynZ
n9lFg9QvlcMJRLJfEteIloRGc4xj39PAEahovv4fY9zFqN8bUYcYJXCrvz+qXsA2
0V5qHY5JYbKSMbPOl3IqtXROcSeh0mfPDpre0tKiDWbc+amxFUxK5AsKHSftBfTF
YOQ3Z7TuyO/QWuodP+iJcvf0A+lluMQuMemX318lZjslXi/vDbyeFZO41y54Ir9B
mjXRqDq8vHdpyyM2vhH0sQR3Iv2e+glD4bHDKgI3nipqHTB4xRo2Vlk2Rcl+mnoz
0qJk+6pcoVFWJd9tpVR0w5CcF7RsPpdVlcZs1ESrjBQmWY4tpHsuFiEnESb9kZ58
XUeH5No7orZQC/WfcrQea/d6e9EPr3SK5dSLS8u/zRvyfAh3ww23nowEBggzbJ9L
CAwiItgqG+/9/YoDdVI1jRMZLzha7hlUKH7SWWn/HQh4q9X2tftkFBRldoSa2QVJ
QTnoU4EdyjHg+cmDTuvwX7MPq4NZ7UxpOgaKdDKIUCL6TwXl7Mr2JkUqz+M0uhgW
vhnj6pDuekuAd9uQfAHAqh3hRBMQw+vjZ7NjKmsnas+VxcgF5PGkwrv15n0SFszj
fA249n3nu1MC1juSt2nIcZFr8RPAPsLVOWULG/7Ajrw8I8sA/2GhO18jzFPZpRr4
SDjkEJxKSirm6kgRJWS1WyfGqVQ4R1sXSPxvGrlqQ+STCSMipciYQwDwlj3XA71B
oL0a2AB8wBXfTyp1zUpaLLBtwjYfvjctppk59ULtDMn8vH99KNZ+XyGWNZDsVMV2
CEd3IUqh8ASKCathU/xMJhHRMhRflEvbV3GvXOCW14cGXzT7GHcDHFtj/sVlwN7u
wiLnBIyqB5CPxtTuCKAfhW1spoS0a1OTWcE10VMlXIY4JqgBIDAaFqYDkP4cLnuH
1Ufzi6/GB1eNlRjzuzVA226CEXE3BOapv9+dZNvPWGSGGTZgbBm7dDWVSk5t72gS
wtxFDjfSYyXO7kDsPyrELjh3z7l1+OKQM+kjrjcQRgoW/C33nipAGgiuWga1ItbP
KYMa6PATJWkeAcdcPnihEWg0QnZoVpczD3NselaM0KJ0kHUNEUB3AsUgN/IaCEUy
wSjo5k9lt/gNVbExFkNVUJlvN7OQRn8M8El1OucJJr2WSFv5ZHz7kpm4Ix3GHYDo
CfbHN47B/1ehNFZV5+pFb9ErVDgmjtiZOsn+fyhPRd63My314Vn893PO193clnkp
xUvH22GqTdev1XRTe/XsIt1LjpT3iFVq7Bm0wr6pn8iOvXNGVoiLlpWHDmSmtkC3
oBCXpbvfsoln5QSmxqilbnS/N3okV5jEPIzJGuvakG9l9HLZEZboDPyId0xDSN0w
AZMczHC4Q1NrTREGB3kN8Bjs+Ekfg/yJkE1rvE/3/dCy6JTseCdfxvwdxBbeJvX+
aNhaT71HgkU/b1AclB2m7XMOP2t/Gyju2k1rGhEL6T437iabAmV8fcHNCPQaTdYH
1lA/I6Q9qPI+YG6uFsqb1Us4N2IM98hA8npd395l9VVPPTNx5fRmUdGjZmOGgpxx
u4YFI9VHz01DajKEoA34BVszrwCujJfxpKsLRsEW5ZX2SweLxQxT+08kSvVMeXLU
RmhNht2c3SySa7O0UY9mFBI7d2nMeqn7XVzs3lIROzvyKGszvEGUxeDHKiDlbdep
u74nrxlfD7m9qhbM4zVDpiJNHvxRtbg9oha8gZU11AlzgIrk2vSHjClehMe6fsFb
E4nMVmX8FUrmpTHVaxOYmBY0gp1aegufxS+/lflDV8YmnuFvdnhx99lq51gn1m4e
3RKTXUv8JzX3Nt/4DXfgwyxbZMAN31aXZ0nVZfxUB1K84QZjBzPIBZHzN6prQREP
y5mOT3FFasAWCDwFksOAY7xpxmJ6wTv+nRjS3+9J7RM0BhNtoPIYkjoV9kxIW15+
xBF40AepC5YJe1Ql6bse0XjM/dRdqonLwmsx2GgW/Ovz82NscDffKb96jhMxBkjL
+YzgyRkom42PlyAFCkWyiVD6hT7hkthaDYJUQeT0enSZ+WlXjOkdlW5kozancao5
unKHiL0Fsix+17SUDQokvLf77vFDHUP1xVpdU3V228NAOdBi+7P6bAwy2y+WuqBj
sVosc2RLev7hrictydgoam2yd/u1zM2NNOvHsUBpntq1V/+iqA3A6ET8dw58afve
LXG5ho+4lPq8bu3bHszbYHhpYFJZZunJytVxRSFIF8cw8ynDbtSIPwrkiPEkdKEf
6sdVHWRueLtiAexVz+RueLj7y8Ex6skUEll6DHwLEXEwLYstawcVUlFj7Yqe/lKT
1Ck8UPyytIw87kD8RHpfNuL8o56JX3/8u/rjAnkPenD3yS1foJ1ENdNJHjByj5LN
AuxWAWAWLPhfoOdobZS3DYvRgXbxkhPHcXd/dw9PpBXLV20rC4mUXWXOxQ2q+UjL
si6Ol6zm9MkSFigmwVgUMsy/U3eIEG+gAUFqZOW8HAN1Rx/25k4SQlC9U6hRyats
43z8HJNpWWFWBoF909cFHpRLAI0OdVjvLD+hh5XudDQMxMWHL8s0lR7kirQaJU2f
tZJ9m7bngfrEd2ZBfPccLNynDliTNkB0+OZiQcMdPQiIVsepqSlDJFzUD46Yy0TE
xxmsNC4OH0aUcprYiwpisXrSllqsZ8/iQFBgjv4LPJaExXs8HPwg1jGBVpzQuwrJ
1BrMae82JTX1beZ73sxQkwjZLplHfHLRTp69jzphtx652uXP2zvBSScr5DnHh2We
FNlE4CeVNUROV1jJK0hZFmnt+NDHiZ/KfJ/KLhUJ8o51gNUQbTLKS8CynRfH0ygM
mhtd+UIZyc7FTW4uq8YynZroZFInNd6JMxcI4eEacjLYa5rxdAtwSh7BXBjx0Oas
g5m89N40Hczr93E3yHo/FwB9mZ+6P07teWatKmAC6C8GHlcWsxxCk9Rh2GD22/bm
NebJi3+7a+EDKZ7FupIoeZrSPooyj8swtO9Aoosjw+VuWr+kXkgVNyvfyU8BXBwH
HsGF9SBMBOonGQ3JkP9rzL+ptoQ3PTkaZWb7lEthxZjIVPRNBvjoTAtLG335Aey6
VCUgO+c7PBcx1UNr8HpMlj8LdJRSzBXmkSMJwWklO3BdJyNxIrDiv+uld5hNFUVp
vGE6m4y1KB8PXRb96/7GRr1tc9V1oPD7EdmV/SZpGmbkMECQ88YUoITBiCPQtNtt
ocxnalH2TnrLf0ln3M0t/djscDiF2ZhgxeFDNbeVIMbGbVQbiDqeE4E46/m0g/HH
Dqiy0dqjpdZVa5Dvyo0X9S/njRSkhws2J7hHd1QsnBgOeTMirI0753PkLzwjZNUv
6tcys65C2MQhcjddMZ5uRxikA8yTHzbUkX5ZGTQFISrktrMF/kZ8Wk9LMpCZBLup
SPZEkMtvf7vdPmnGl6gaCl1eLZVj3pBTgcvNQopdwchG61CF3ClbxrGmT6wSrZ8d
TqOfKEwy21XaeQ8mZ5hNNYqa2vtSUWDBEd6/fj7yPW6PRrxgH7K78cdPD4IhyYg1
AAhL8XQbf88fWsN51vSxj5qui3AVw2p6aXkUHKq4cqSOqbTzL2lq1nmy3gblYhvw
PEByv6gKEnOJaYBjg43OqMZLL6hqldS0Mk4ZRUN8kEk=
`protect END_PROTECTED
