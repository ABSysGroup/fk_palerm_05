`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sp9yh+LiQQZet4nU64+IvwWZRHz1PCu1lKjvadTK8Af22W1g8mATSB4wJmvOkleK
9Vv82M/jK8YLdF4zXz2w/MxPE2me/5Ek76ro61MhfwYcY6yz+dVK0qkyUGJtWcRh
HW765qE8ojMVdN3aO0l6ypaZ2LDOCKekhQEnzMY/EHQU+FN2yzAPoI7LlkNNBLjZ
XKDbmw1fRpgxPa6FBRT1EgbW7CT40ISpGTGLE/QEoHkqaf3ezMY91RfUxAc5SAeu
tNbyznPi/vZHfxFz/OFnSiIPx3yLVRY4QURwOmJ7JSRCG6QVNgPaGeCB9BnLH5Ok
JPWgfA3warL/yDcmXWKDgc7D3egGi8rqcPqHy1Bh+NyjJNNxtglSX0mW6cbzM6kV
Rbvp6Amm7EfgwOdO+c6HqypHLsfnWYk05qZslB9/q4yIcrcdy4BxOfBoGch7ByxZ
dGc6ihWTYfzM1JycA4+T43eaWFUOX6+b1eeOe1Z8lY8UYQb+5lA8Niq5kf/v2Sif
UhHS0xe3oRc9p19Ou4RbkR8MBQfgtOptum9EWjLO7U7zqku+tAdKSmIZ7p0X23cV
0QOU1/TGRrPdglQqdN4p4oxRsQbgJuBRfcoo74vY4pD/wRA+h6y3wYuTFCLunzG8
YsBkZfTiBTkiCVQZtFlwornXv9WCWp1OLsG5dflBjVCoAfyf/Y41wCO6Sp9Bk/Fk
MMDxEL4a1wFlNpGkNmH4a04EV8nat9JTfwCHdKrdqi7Pp+6O/PZZEQE54JK4m/k0
WNzdrgQ7RcBjljSnGD3JuEgE78MyoBsRA9K1lt+8QZMDKEEZdUrb+A4xIbAYDqVb
0MnrhTpc67Qcdb1wH+LiI2kA5Ktj+wAvTC/gqWHxvW+RHdo60NQUhpqCILWz/HYJ
4TKDM5PChdxyqRZ3Vph3K69rUkmYLemOqTtWfmdhARSNJVAFAUwymAtoP5dol7E1
SGNqv0erlARpGT/S6c5uqtcpzngpncz3OeSHBVYvfYahSgq8P93CuYwLXWTdfZW1
Ni9Bn/Re37QWW0x6XAbZ4cf3t0ux/90+xZK7ptru4w/iSXvXwThElYEa7J+RqkjR
KFn/OnqMx6S706s6D2/u4SL+tPc1qW7cl8J+xRKkwrUqIxQad7s6DmQMQjNT8uQk
ZHwTFfZ+ydE8XiGHRMzXBqxDq2RTclc5mJkjOy8lkrRVutcZ4w2yAtgw3E8eDlBd
LGqDMTWHdQN3R/Na2TtqCo47mDtklRbeCDXHfP+R/x+0qZRWclXCJH7r77efng3B
cTrOnPlTE+po86T5dxDuKVAz9cqmKjv54m+WHtBq15T6BS2AJi4xL5z5pe8iRav+
eS52OBr8lmQ2l2UB24BnFO2ye880tAKeEQO48HroulY1J+5Ry5CLxeEm5JQTmSgp
mOtTcGGGEscnUrgJWUvXsIg7RXBHy4DEO1z/lD6LRiopLZL022PapvCkJ6YjpEYK
ZmvXEECKvCMVsO7l4l1V3fG/zeLdNL8HWOqVcn3aS2LiFPtr18tsG61AxsP1RlhN
XdGA8BlDY9hmn5kvXLpGzXbU/tHmkUFwaWoSfu1eQlSlimncpBcV19Qlv7Tmx2CC
r8xEOasM++Fq83hb1HlSvsO+gTlpy/cucXGBC5cCYl9OukdyEXDeyvgjIHxJUuJk
MKq/UL/bufZuNaJMoVKnqEXf2K7b9b0NE8rZ1cbxsEQxRcQ99hi4STdhefdLQjlX
rZRKZGF9iIC8NIHs/GtpzmK4qLhRm0IQaRoa0c76/BisCuhfYApMTWk5C7bwAR7w
C0icAaF+vBrS/ohF8oS6C72sbYl+6UP4EicZwz0GOIF4u6LL0oOjIRMHTf9QIkwf
Qn0pKen5eE3C00F0JiCvfoTp8CrQ6VJYZ4ZFV06wguPrzPZKGvWUzmyR1OFF/XGl
D/l/u5+tZ+nQ7FfviukQlWNNycszgTx7zzTVQEPiRhp1Rl2dLEXIDMi6DVY9KHXB
NaAkODlt/Ck9c/Whk1g8HN2/6DfNTiZuvepVqRyn2KpaocRbuF/0CvZ4hUe0LVf6
yLd0dI/+cog0/guERpJqGZBX5J99SSgjzXv/oeGOVRz+A/OfgZEwyuNGcEb8dd58
5YI0/FQpF+jCa9N53B3NIyUdAFWYL13Im0AyRh2OIGJBGVrqO5zeSdyv30J05qx2
Up0rOfp/m45IHwPqSLvJzKFJW4Y1dAtPS/b2N7ZMRc1MQQHHpjz0eEBR4DEK8SiS
9iqx/gGTJWCHJmbfpPwHclRLnrdDMaX0qHROTIGY6vfmta35invh/0uHRuo4idMk
IkS5+AizQBoauxJgnyKi9MZ9GVLSSqFyttwJ3bulGemfBGaKIN934MZ8yMtHyu76
m//2F6y9BWtp3X7if1UG5oLBSh2VjjnbdZra4QRSnzriqNbsf/OrfdRvd7PFL3ZO
zm79paeEaRYRCETjyFHGZkj8zhvCQ5pkz0FfcdyeBsXCJWaYjHnHJP6rRPFFbgur
Mlbcm/L0R2p6CwdeAu7H0t1W/ZkUQmp3QvZ8/oWJDwYbPnhYWgTSc8Bizf5kbGkk
EMTpT4uZiDri39bQvnbP3LBeyRwYwCFLKdbMXnBtQv1h1kNugP35Q4jHpE9omMst
s3ThMWj3xe/nRuPVHYK8CpP8XNLk7Yu1/K5fio4ISwmtFY+4meDpOFCLbJk67zPB
1aJNS2d74ysk2SiPtmfNw0YOguDChby+zHOV48bW1chk2idOAEM9baIDu3oILz43
6DnpgAxrfSxxa1hNPN4w6MTh+8fTPlysP0UV5VTVvd/oG87YGcVy1CaMfglZj2Cl
x4hqeqllfb4xQTQxzRmQmXemBehLI37eJjTIfch4FbDiHm8DdXyfcppYXV3yI34p
mH6hlrAv9Mg34mU6aCd1TGAuj9klpakaRw0FMbNfbqnhqptcyCKbEkQcLVbQlmoz
iziIX2GPWlgv6QFCAgPDi2zTtofBIz+MEuauIwCLEUAeTRozEdX8AY36JXP0pTmQ
y9xeycgPs9Txqu+JBY8MhCj/90BXfJyzZ1MGAHsQUKQ0x6pel00/llbNkS1qaeXS
v3d0s3tuo0bb3Oz+Krv10qzfeaMB8Az9qrYX4M86Ph5j6m7QyBPf8BhWlVWv6oP1
iWEGuDGTW7dVhqno8w/G3qlg3/HO7yomvLG5hPHNBcFe/Zi5EIAnia5EelRzlXkx
4drBc+MbP9P/fNtUZHmkt21N6vq7BMpYIjJRjiM5uvgpB0P4cUhcjYw10tMx/hjm
iGE1JCiayr47Aq5K7S9AFtfKyOj42erqevfGpit6IdmrGiP0zhgCku3zaBbjrgXq
ICybiOaCu9QJbgZoPjxlqYebHzvN6Q6O3VWZMhs4JQjyWw9VppI7ZUCd6hXE6CF4
Hx7cVpcU3Z/QzPX0iNvhqUqkQ9tgE1ooMQYGM2it4OVL1jMxKDcZ1j3rjfpZwb2u
Klw2lpWMLiT3tDloD4x34yMrWN6sULXsdoOPSFzm/Y5+dn4HRdks0u2qvjtRh+jL
dMUncrcIj9QK0w4IfACchkoA6vTbY5d5l6axNMpACbf/L6v7PFetKJRXPR0V3ykZ
LwEaLoZ5vwmRmFquN7n67uF5B/nDHj5KrJiFRaa2Czwti0SDvFZ//DisgZOS+qkc
BsjdoYU2Ut/p+WCSrX8rKYKVo/2dXoF8gIzQqbFOyNqbJlLxxgkGip4/CjNEbcnk
fwJgy9FgkyFP0ae+ezhYzXm+J4Jt3voERFSYJpgsZ6tvHxYeL7R9ww5lswaGwD4B
PtGrwO+EMiUBKUzsEEWmsLxFzewXoSFpQv5GHK5eb1Tx4qyWam8bIe/f5RGu1eX7
2Y133oGbSI5PTrM0Chw1I1qmb5TgSCy0xmdJTHK50W/GwoT/oiMW5swRgqJKdKfk
Z05B1O5wKb9G6JWDLdSQZe1XC9x2ajnr99hzhVKTp5YP96CFg54DsLkmn/4NLUUG
yiApzq+FwvNv2z1J9TlnRXDvOU0jt+IgRsHp1ReBZYVw42OlmY2jerF2g2gwKL71
e11V9ZHXwPS0Im0PdPc28dKMInAyT2pC9Bfct9KcDRBoHKBuQTLMcNjfxHD8I5uu
GAS0/KFLtRtJSVWXOFFhC7lWizQzRRlzEemFfTvwALMohZdEoUNx1hzgvViFRdMY
2ZHSiM0qE8ewY448akBBd0+XbTXpVlV9ujmxBvFAtfHQ+oh+qxr0Dg0AgD8HE9JO
717pocxFJjZcdMQNPosBSKNnBPiZd6VsFzQfBdfSXEAu+/o1tjncCccuWk74d6mN
UpDfMG9tqbWwT5AWM/pcD1w+0L4ZDyP3WBpaml54BMagpNM3q3gpDBXHlfXHEuKL
Yq/2GU82vo17k15aTf+EDqxd3x23nF3rIvr4muZJTDbKo/kL+V7EZtv8xFDUwMFu
01Q7F5H84i4Sbmh232k4RlvDNpg5n8L/5AaS4HiP9YaM84kadckiJKQSUYL6Y5Zb
xFDW0KmieI/f9PH/jtsfUL8/wXe6MSACYB+a4VVSzIahej+7dR/1s0PKeTSEk6MH
oQ3ArdQg3MG1iIrqydli09j0rq1aVX9jboJPYT4kCzlvxZpghXtK5mXuV3sIz2W1
ACttN/IGJYl9M870tAbQ8KypaXw20bEWX3MPpj+zxHg6YT9tY4xxjcWSeuUlpIKu
Dv2reIUfTi6oQLKdCOoHNyfosHIzqwGUxutJAC9aM3urJoLGqS1qOb/oKdsK3QXA
B9ocx0n/6I5QxAoht+qllT9HKJWIuTqp+tsSveRKZBarImuAXBCAgd3bVDU64qHX
NpQ2wZD4Q6fKxr6JdaGYZieBPGolMZ9K5GEI7Ydmyx60i4HomcFhXpwZ6HNyJYCY
qh5L+6gKhwCiBYRCx3t/57ak9y6S0ed5UuJqY7Q0cDNRrRLQjheBE1FPCAr59nD3
yxmr9KRArRlMQyAFMKCTrTVTtR4yiyZtWgUNCm+FnobOHErS3l24kwknafc5JYcW
law8Iv8vzqbIjYD7M1hyQhvCbI12mrkmrbSw1T3dwIHpU/UjDQdXIDPyFmoqXV5W
TEHVvU5Ti2wX01bI2OZpQR+icl0cAUhkXI6uSetMBzYuZ28MWomTPxM89uYwcYY5
DBHgwu2aH7oq84XUB/b0xF/0qV38F0XYm5xhb6c6FIubE5fghN0sU9hKRQusREo+
Uyq1KGnpl0N+INfc0ix5iCCHl0OI9d1zYkMVV5gAsiU3ULsfq71SFVffFhR86qgj
GVVpn1K39M1GVn5tMT8qPEYgZ/Mps0f9JpaKKgb9Gr9MSYGXXW8iDDU8Rcdhucd5
qE+qxUkijZJ3MwwrXYEWyHJ0M+Q6qynTN2+8s9xzAaF9D1NPTwFwJmA32+oh57EQ
8DCHRpIyKnT60gThQGSr34UI4Qj9HZUTH/y4AOPUHHfQMnvEmmrQpHqzOb90NWfV
iMW/PhNjfmrIxqey8KLNOXiE0LimaY4H8KfiKVOrODsVKfUamPoxtAPkagJBCh3W
R2PKFKtJP0hYZGSw+VaKnqGSdsrTIx7LEu/KyOvPjqbc6w3tAjYV2S7gngYyNI+d
e6snMvXcH6WXiLz2THB2TBFSZdXG4rH571361ON8gYTkl6mNUi75eI8cnMcyOPR2
J89SYzWGyzmPJjdbQkjhxvx5UzLVAn+6DHsxjm2yQudN6o7e6Q87DqWMffwfVZ62
ugIxsEu+jfxIOekAzc1WqvTmPiTp6/38n7LGsx65hRisvZ8HB1KzUEjkuoXBBDoO
uPJBiWq71C/KlXIMc+sOY9Bgq3DWNJ2xbT2THFy178j6yhrEaxwhKc7b0dfdlvH4
A2X3ejlg8wLmwNEZNFyvkpPhuUub9OpIRM26TW2DAuKYcgy697AbA59DK/hwKBTC
D+hdAzExI5cikpqTG4dvBJwOnyp5/WVX9EACzlyVZiAWLx5kYB/Zo2EmiYIOIXBm
sTyf978ACJ6YCh9Ez+qYExg1PdfWj3+NGvp3MGZApAFS2rNacTiNtNo/alfHi/jp
njeRcYTzK0KfBTbUCAhCydod0A77klYcZGg2g3QQTHFPKqUBtBBKCOkOkZAfonTM
Lj3amdruvFCix6tusA8mK/fW1yQ2ejMkTKYBvRZyi0sYbEorLV+HWBaiByNY5wgf
WFp74y52taaml6EnAwa9FpD/jrqKagj+7M3iSigMQkqLIAHejDcpHFmX75riH6Gc
aPPanLAfB0N1g8ywtKF/e/PW+vWFSpgTAuCk5WW+phb3IyzhPemyYGodCzDAmROn
fd8v9xKLkTbpIqtccdf1W7Talwa7w+6PsfQNj/29DjN5WLA6TlPaxqRcUtNk0VtF
QkDjTOLT2T6KOkY88Ogai5kMbEeXF9qw0MrmasHWCu7wAokk4OrBeRPKMYI0pXwz
NxNGNYLHwuSy8QLqnSRbTLUZR5/FesA2SgecSRlRFw4t3R47XSRPFa0+QfNnQjG0
NAFMqcc4NXDEFctPE2LCf/OnjqBypOJHDQ1MwSrVYasgb+DU2HC3M04xSbPOGL6O
mOv3A7xy65z+ncrVOnUAOqjH19uLisBRwXQ2Lw7uQHCZHtXtIpG5Qmc/j9etDAM6
FlceI90To4Ii5Iq5lcSLTgbcy9bKuEBeUXvbdBnuDOJvcU5UQsfSCPRRZgzTtTx5
qSTX6FJY3shYl730QvrK9rANfkv/WOV98VEw8Tlr1R8a92gmcOqXfmAQbo9JuyK4
Zf+ARwS9epAhjwR8sfRuyeuE991q2IsB8Pl+qVvZemF008M4iGJbejqkV3NtSkpo
UR5nCylVadRMsA3RJwD5H7jCT8e2jXSp0Y957Qpdor9ZZwlsOFbncD2Jfjrfh5Uu
155BQN+2+J+6FD/fwF3XklVIsM+J7+91DXV8JMV4bsV+E0Vnlj7KnNyK79iY5aqx
Rz5pV+It5fChpXp140HOrf3BALUqmuDOOnSDcjmH7t07BsDbrLYk5krF+JL68GWO
7p64EOttr3gGtNbD+w3b8XYX2ntGew+0VmLzPUDIQVD1U/2lkVcQh6QnasSDtzZd
y2/cbMubhuk8y+ueoek5U3zvV1c8KaPprSMACljagcUBRgLxpkb3Nwe+BsnWbFCy
kC3oNNvan1/lCqqsYLDHMc0I0I202eFMq8tk1C9GkrBhtct3xRfax/9X28s7GRZR
1hykbqEqWgA3jxQ2KY7rBIExTKGwK6NB2cl19/EJjxiL5EP3wiXyEzPmxT5Su+yI
5jTlfyeih2s76H3Ptq6ewCp/VA34WHmrHAXagCWDuhFCxAUDgccmrHC628wQXzO3
XePrCeFaZtzgZRuhPF8b8COXudq8wUMM3LimYRnqNCEv0oGByGa7ybR4AcOkMQ8u
SvLT0QC6PgG9YER3CEKbPj9E+mzaNmlDEQppO7gon76yObF/xceBJ1qf67AO6mJx
PGDI9DXqrLpASn2RHGqLlR9V4NXcRoCt91j2C5kYe7T5sYoDbMmYoiLJ03NQhqGy
lYAEuPJjsTZen0sxmRIxC6S1bhSptNmxAaZFTSLkyOSWjwOafIKTxCriyxg4VL0l
tURDOG3+B9F8feKnUWjKuaHKTJ7vvsfV6VGVwW2k3saFKWAfD2z1yOJ4SH5j9au9
5oRT+wexGi76JVlogzJ9fBsK/USUk+RnOO0T99D4yB7TyQdtHOUf6T8GFmg3PoaH
FzaCxWOTxFITJuTm1vWb8omTwKbZgJc/wxvyctYO7IsomnAhAIxAAMQDs0PzVLaS
8MWpN5/FTpSOKZ8jjhaFp5169PR6H3shiRWYARuGH0fo8Q/gE8vpfWUb8Fr4Ejo/
+gUHQzLF4oGtFTFkXHy4y0xyYeF66PcDUxVrZyntipCfpbSN3YPWPzeFsPP3cPLj
in8HRRqj36zkLMpomK/5WSUAfHcgfVWFoKzPqogJhwshtTMPjA6Sur5NcxWzCI7z
gxbweBIYZVzPb0JtMfyZmBQQvnRWTktGTu+mwKjkRpFQJBKDzulWy/oKyP8NBoAD
4MyBrgH0jUv5m+F/BToeC3K1YyIj/hvM83ghoajrIhOcb7YUqLyLdGzx5WCKagIS
rAuKbyvurLTx4AGAwjElGVDDnRy6BW5BGZRojHUM5MtyOybNUHg2kDess0OS7+Ej
kEYtqcqcW/zSKqascyeBiXVbg7y4YsNYMegW+VHRlBfV9guPLXscvUn8UmP2YTw7
i9RVxcORbc77+lrMbzKAnsyTG7L64jno0d72UUwjYLQYibfaRnBiYVNXg+H69EFV
lwpaXriOut/bFoBAKlarAbCWpdQp2H9dAISLf9Aeofh6VSYLQb/J9Vk3xqGQuxhc
CmYHfViAxc3BZFRNQ7pKEY/sddiIBO29KnhBlKC+rDwq8ZDnSPhNBgIn8mvyVkYA
OA2PWhwauFs0BKmQgXFYs5RxPnNxU3SufvKo3kvxWqnoqWtCIV+XzW+UhV50oF3Y
y84vA6v00cOk2lcK2GMkAsVSeQlXHI0NM0Da18rFZbJVouFZnu/cLARx5XRvGCUu
M186hZds39lQSdEEhvQ5BGgD/h1uD+Q2YZMc8oF9fjmvesjd4fyckS/2ElT6XTss
qvssNbRq7+EhL0+0buYi+xn9EliREZ2c1H3ZFeKRbD8AeTrKKCRuvqbCz0Js5UGW
iXVlPtwrDvyVD5x+tfTU1GejwW3/yqd5rtQJGdFWdPuCWr69NbT9mU/y2b3J53Y4
gU64jJBHRgKRg+e1FXygkdiZ791nKbajabDcOuEarqeUR0t0xTZPt6MGmIcDUuWp
14WOKHc/rJwWu6A96Agifh9llSROJ7MzBkpNpcCFTNwiAPUTletqeGQwx1wDZPq9
oRODLr2IJrqurQjkGwST40B2mXBYaRWXVHF8YoIktRsOBOQnPAxcrOEzXOJnIp0m
NgBs3gTM/BAVgcEq9vhB1rnNq+SOMJl3gPIyVVec51BLJwBX/J9b6xpVzMW10MyU
YnOkNo3Di9Jz4yFGQetYcxplcSoORLGhsTAKZzseHtqqKW0orRkeQcFY1NM0snD5
3Ff25jiW1PAsmAGPc7iopUYIbkVmlOF5HXaoX1XBpYqvWiox12bLNfQsu/wWF3XT
uec8pKA41lCeOZGmKvWcHKaLDGQpp+Pk8MW+WKAc7hVabYulnrYDe7V4C7qdLJKK
JiuavLwnnINUcTKr5t2bzV5uONlzqL+tm9He4A9gEB/p4V5Lt2LB7KJOTq8Z9iAb
D5XGUfvxSfJn2Q2v9vG59/iBNv9JSy0x1aXrfq5tROW19o5Ad/7pLqdEGIl6ByIT
VQrbt2oQkcJFW/0J5G2HUmZYpPeZQ6WeJAhyKn0FsMBs/V5bU6FBIOiJ6hJwP6GF
5PtcwlJpAXElerDyhBq6wtBZbevQ90tIct36KGIvDJQNSDVSteKzMHuvI2fOwTHg
MrFnWP4rKUR06RoKqTBHiplFpl9DveL8n9FcnUEUN5YrluEDssYJ7TSA8wUyImlt
2gOV/xoWLgduXjaieatZ8aMF90FE0oDKyyvIKDaBwUJ2njAehatgIcf86+w8RX/C
4J9kbeR/fbDClEbRx1TVQ1NsNF/Xf0HH4V8I9AOkmScvnhN8jnkKYEH2/yTKTyec
bL5yO9k/9CCitdCtqXxsOkfxxVE+VJFP4RVUzs03DULjXWi63TMkxMuIVZuL4zyF
uyv0zxGWNcDH93q1BlCpX9eBtaRvn6ZBJePBs8jiKRyFkn8eYN/G8idxnSlgc83U
3dJWuX0t+Nc+RTNpb0wdbhrVCBxEYzfJ+rnuWzFa42S65xwOKJkwTvnSk7fkoidM
YCLX1nvQMpJBe5zbBXavClKCB69tQLHRtOuMfG1opkX0jjj4jLfPwMTLBFWX4j5b
yIqLz0QixN9CwNaNprCIkOKXg2Orx6C3jg4TvOTuSNhNleN0sX9twDGNojRXCf5K
QsCl/OFco9ULtzTXPONAdx3pVQ66n8CGVttU3q71zxOKhTRX3Oir97OQRyaRHTSe
6/t5w834H1Jgv/mpu3wvuu7Y+vK3IHHbEF1aHkoO9l4eWhfqFIf9342hM43L7KRe
/j3wnhlDqqh3qNE7QeTcAYClC3FCMGxoAgra1VpRt4ESq7Jdvi6IQBlca6i7eDWL
mc55xapcOW39O0+FYW/pNawn+CprRCEW8RXr9siMA5r353QDetACWGhWypyEdwlZ
B1OIU+Fk3R/XsMLiernK4lxRUlxOFKpwoMR3A90BQQU3caBEmcKFBXs2ePTPouQV
e2jSAKKORezt3G1W35SHZtOyahxBGMyR/MqklBJGJU85tfgm53lRMYa8s+UVGgKM
eP+XYI+rsvooU0cqGxS9Nb43glnGI0mGVPvLjRheF78mPiYu20xIVo+jus1inXjc
dxp8uDz+p4f9Y/oxDKw0oMHN3zhYcO8ht7mtBG+/F3hdJsXD1WMPX2i7MmooNSr5
NkNxQaSmLszVZ04srExb3jACJc5cf1Lj93CTeCs/22wWWOHpo9HN4tkdwhufDh1h
uOIqFrlxZMqCX0wWj0/nwGZdXkvoctqyu2so1Th3LPhrqK8b40JT9bKyAQMB9FPo
Ml0qUXJOCvzOqjBPPZccEbtl/NeOsjtwauJ2UXLwi+BHfdx++wU+MEQxNUtcY4zk
6ajVBFbK4CZ6Lilt83zPhmQf4JxwqvGYAuwQuv+3ETCNrf6pjttboc7jGnuPoch+
jNPE0Fm55+quaX4bvbVHeR3VreEtW5xRmyc/lNjC43mDWZGyVvcPbeJEzLod/SKL
aSrJuAUX/MFClKysL0AOnMg4/Kp1BRBLsOUSlTgUBNkSHqS5dF+rSI5NtDjCvFtq
GAPdrtiWPCc6/OFTDvQzBwk4YOlwRofSBdNABC1fs2hJObS90U0GDGIaOGl6Rvjo
C+N1e5DV8hum7XSnE8csY8qk0AtUnNgil2LuKh+82M6Fs039ovvS5Q1WMH+FBbor
YQnUcRl8ssSRKelW6bxAXTq+90EcAprt7obFwEUttZ0IWA0bB8n+0XL3ouscQyVZ
PkSg+jwYwFM2mG87al+WqoAdhEu4/Ic+TlXvuiOSJvVd7BG46dRS/AtVVcviRzXk
4/K6+s7KKr1pX6Lb9MosgzU6PKZ3m+HITGhX6GVlrziH4FYSi+WfO0i8xk3Q7H29
yEFjo7m9caHth/IKTBkHdY/EWSn/XXySLXZE5rSwQP3qSBRxlIkFQRwk5u2uQbZk
O05WRpdor8Ec19bfboa9/2/dSc0uXbaFPWV/eN4QLkXgKyA8UkIjLuHHXGqrVE6U
GBgVwMnrWFP8UcP9Bqe9U2aZTI43/FNVxINGakTQ2W4kel3q3iUlIwRYkjqPoybC
K0bhvvrlOeCqRNc9P39tG58hES11TcAuCMTz4KRyiu4axWdIlk9aR0mH3yFihgbb
7zDinnT1Ti3ifDuyU15IGTImJSTTYuHSUHJypjW6QWyE33rMxRcPopRSzlozEeXj
N0kwBtkCb47hbLIHYxf8b2xA9BObQxG1MjToH8yEeMUpq/Mm7I5z0KqKj3gxcV6L
/9f6Oho6F8Du+3TVfF8zrQvYr7DYGDGIYoLdJU6VTXS/PZ/YXQqJ0rh5LM/2VqnC
BwXJKi0qAaaLfc3NKGXUjHHONCvZ4m7MNjSLnwqr8JAfyqqrwmw+zJQuBQh4s2IY
tSOlYm3Z8ISzn+5OdeQIDlXNkXlnQ9qGofod8IY2WElenHH4JmNZeINhPi3iz5Np
PllHDRhyosQ2YyYTis/zeCRaPWYpxBmh8jYV6gCctJSVRncrjOfsJLUG0VyLeuZh
gjK9HcDTL00C3rB3uzpmZMo7a50j1fDFKZIMyjucDPFrNGk466P8BKvxx8u8UC0I
Bq2IrVFC+o86cYgFwfL9KWalXtd9XofItWohYSyX81YKLWQrGbgyXO3Ct2loWPYH
rldb9tdIzYe8WxosTYibvmkbVIK/Ur2K8TYWuXAtJEf43BTQSYIY+WzQDs2dvZ++
Ij6rFdlxz5sUpIAyEXlNm/uDKkPsZmj/wcbLHXlZyVVXkPm75YcgPSLTW7tT9x1l
n5Jg060qfKBGXA0V5lCI2/qh1pc5b4edbgCexgDtZQsHsI/uaq21R87RvpySRDBD
9F9VOcj0JmS8LmjzEjRsSOu6MkNVCp1S51pdHApTEY/LN1ZirxUlAce8cMicT+Ib
9CCXXGSY8ACWE4fX4xpm5gyFzLO01Jzbg5rMVPkDHRCSWILWLdwCeBDLFfUwWr8O
/uJU+uHJWplh6zZHA0b4tvTqiSMrR6V+JzAWQ56dEYI+Og2Y5jFkA0C3LlahQ+6f
/t4UedkgdXB5Q/BHPR0Om+4eOpGFo/X4ROXhOXz8z0/v2GERI/8CPvwU0+e0Ix4d
GahJ7/bl90FyfXOxyON7usSeYYooiGKbLXOxl0eAXd2oBqepDI10K6xRXRDaOOcH
oZqS0QW2Ds8Jwo8aCfOdKEuK0W3dOIiz/dVvWkEd5fK7t7QO53+BzJ4PjQ1AnpsB
5f9J8jWoudlrHftZWy6Y52jiQeal/d+hmFfoOI5rpGj97hf2PIXAcbU6IdTqFNPc
RH9yEKZ6VTn5yLfLOplhBcwp8xhxS4vKsghtILiTHGfVQDWwXAD6KGOZMa3EH06n
vsGrHophR7TxcQG7XGrrMgTnjECkQl87xfpzqI/CSC7enVR53vvgXHlKRQhCvhIp
zhUF+paVZKfSG3LpaqcEBn0eap9hCCV6fRqRRFqPTs/Yg+6cqMmSh2bHYx0gd3Sq
fYlLiUmj/FuIwHicquYCpLByNEhYia2/coBawS2TRgY/cvP7TAhL9J6jYmZ8Iy+r
lRSODMpn4xqIAuYsX6Z58CgbdvapX6gJ5OvlSUVdaWYgT3jSkhMnHXJ24bH5J14H
+skWVxf9d2+asm1cfpRm7IMVmPH0D4Suxc+yuVnt1fBprOfBknObTes90R1EvRtw
xR8TfGWzgYWIijhHaV+R3D2ozacKq33Yta8PxY3X2jY804Y6ur6Tn/b0PAyYRNPB
Hj3yXEeCu35Mp1lSHuj5yes2Lf1II+t0IeDgqnTM+nIe99ZluuHHZpAPWbsjMmKb
0F5HboVtQI3EdJwWNFmnISeMQRevXlRKQRDQbxrsp+DxXJsEGXSxFYvSiNMmek9T
8of5GcsTISHfl+x6qZFbgDFM2kYnSDR5s2ow9pEuio+FCl3EjydcnZhs2ZV2Xsmw
iE0NjYs9qw58JUIOryBLDJiJuSAYaap5Vq/tzHjkUwVfdY9+ZJ/+B5ey1t6y4eJU
QzRndI0DX+yw1i6MmZ2jOXguEeNV+NUTlV+f0HIzUPqTVTUFKo0zF4MMOQMC8yxG
bGCGJ9EMZrjxwdNjQT7uoLeyLJnFsL/eHIG0tM5Vprlda8P0f4EbG0P/kN+Mxp75
fwkBRpJ3tePQaNn14ERpYh5vD/Bhye9rzu+dLRSQGlSAjUsU6pJd0ec+d+xIUt1I
wPxV8iKdqJg2CUurAckOr7qM5nIqxdH23XuPkEiab5uMZ1mXLb0qNmAGDn2tPmwW
ucQ7DAn23TMdo9TS6RocySfU8lmFpyfe0Szljfeb/wu/GoRcxJO6Thyw1maffUTk
tbskVFOAWQpO45RtICCQcEIjlYRl2drNR5f+3Y0A8+K4DBXbaG8t05Bvl2TF9f7I
DXmoege+kdnbzkV/q6mtFd1tRKQYFbkj8KUKmyjkXQ3LqiF/61Ru0Tya86CAfH01
VapTEFB6MFCP/aVQ9DLL9g0qoDNun8d1MLoSGbxAgYxNO2DLJ0C1HfgvKx9foVXa
4OvwME3m0AFzbf95b6ykbYjM4d3wR6Jz+cVScELHUkzNho8pAA4skqocG0yWI2GB
2lwTVOqwJcf2mNf8mPjuCH+S5zOL252eIqLFveITOmC9JZMR2aAKtDfAysniyKFV
lJ9gZB22pxtauMJbxhTWoQvGtVr9GmYcqN5hnHYjFQl598hJqD24CjuyA52TeNiv
E8XVUc4aia0YqxfUKDJaZhQKtgf0W6ilLDUeB7d2KMPJ7YJiRTVStanAJWHPPCi3
uG3wKb5oJNcuZjUJ5vZLf+pu6IPuz1CpHZs9QNJt511onNrrd7xqOFt0TQ6c0o9e
ze4BLqZwjy1h7t1w7ciynIUAp6qAP3tZJHolpiY7YHTyl50OiFxXPK/mmGvkmIts
HuJZp5fcK0K3sx7hkMu3BpdW4j+IJZURTrqBFa69DdbyVH3FgatcF7je7pN7dz9P
LcrStMUgUmxLBoiZsH6xWDGaP8e0PzwgZ1CmUQA4F8NfnyvJ0yYbKKddkKGV0i/4
p5UWvDKhgobzzmsOAtT6ySKmexLFWAAmNHTEcHijFnRagujCudrjo2TThQ1ltWx7
w88g1UP1SdoBbhnfoka78Bdj8nlFE0QxHUJwvvrH6Drdp9M0roZ/clf0vtQm3Wyv
phA/Wbtfedc/FdITBwjQO6IiW2Js2UkHEJASKSfb587FBlxeS+FXPQwrpzbtuFxk
r1paUQUCEgqZsG7zSr49oKXQ/vEqedYvjcbZIxKMEkqtb+NznIVeqLjZ3Gg9Gjn4
kc/pu4FV2f3KbDVA8LeioFbFb6UbV/rUEksKqLqzCrYKSyuS/nlq0Gy34E1W+/Yb
NRaASoNJA3Nelt+V9FtqGiRXCF7olUL1NB0vYzadQptcyNacKvXbbiGQPzAYs/7+
W/Gevylza9pUArmLj7/xBnuKqY8nphp00a7kxSbVsd2vbP6i0mL9VKqVLFLetYQ4
/Gx/0wGzZRreHJP1yKkWOvhN1C9+aaR1iBNIE9BFqPq6mkbyf5A2Vd+j8QHnvbQE
fOge6qs9GQpnvHjK85c+utrJnqGf7q3efib4GU4mZt2EwaoFgEZPoKsAsUC0JH/P
rpKrqDbH0phzA94pgBJ5bYhxv+O0eJI0Iu+Thy0Cr15+wMewdlbtx08ABU4kYE6k
5fihbbb6Wj9GNpR29ial++VLA98NCN1ARKHZSZJOVksRtcaW6oIJIW21mIxmPWet
HHs/5p63WB+DhQYkcLalRaBGun5rZgZlFH6TwqwO2tnjsrucbJwQOLj1Sm/WbXl0
DxDeTKhS3qJgnByVy6x3bgnrIpkEnR1+pWhnWKkE5K/NpJoKYcTFnPogzwUD/abO
MHYQfZnVgONfEHSGUUTFZaws/pTn8qiiVmjmSGggBpmDCaZvfQfZy1RNBhi7ah8B
RB/raIPVVA+og97ujzlUHb25hlJIsYxV64IZxxjWi4lm6W0VQ/i8ULhwRFktgQAa
H2of2IA9K9ReyY/IkCzA/9DWqCR3h01Foz0AL3+LuIquU5E0uNW6GuShVJqjO2SL
NIEm+HETSPEWDu5sWHo6p16SbSMIHvWyinZCtkT7DVmvXLPY0XwhdVltpX7pBbZE
K2cC+yPSHjFlJMlPDFdrwzKLaK54CPdGxB7fK/IoL9jUSPw2xL8S3d018qJo3Fa7
/qN1ry6ZWG35PpswzUMsTN2oOoDkYOM7GLlDb0W9BmWtMD7/kEEaDP8KbktUiG08
I7ydHzHBTKOxTKEkoFQUwuT5Ty3wQKujd9uNjeU5NV/sbC2jv3lrxieQwfFAfsyz
d6MpQtfoX3SSdULaVL9xsca5iZ7ij1SOF8FtDj5Bm9A8Q9Y4d3fT5KmeHDrvWwhF
DydVQGFQkm/r/7JEFH/HMLX+CsJzgE4f/No3f0ofyb/LfSGUGLgxmcvEaE0LsXaq
FSYUVLSpruXFDHwIbhY9VuVUVA2Wp78es2tpdHLhFfN5eqaEnVqlAdQfDUPwqIJP
+qski4cmJdgv3VxS4b121RIs4iq4pzbShmcG2MO/OdLh3+fkNPb62O6azBf6il27
ASe7EaJ8Nh982bTLPd98h0SLz9Yw4LY876FSQZfAO1+g39LvkvIJx0QAXh3c0wXP
5Sik9jqapm0Q0Fht6yih3DYNJOptbdXIkmTnLyx7cZSbRvTzIVbWMAvZGpns/uj6
l7VPZyrG1JhifgMPf6J9yRanCxwBzAxekmNkAfOxj2d/ZsSqjvoYRVtA1kStI/T7
mHGVkgwlpNqWagp0KFT4hONp5aoa3WOhtr0upzjiqAvlyMLsFQXA5SWAr9fHLInH
Nkj44XywLzn+5Qb5J3PKpcqEiqgxI75PQP4vEVkc/50/Dj15wIbWVZ0f44yyavEb
Br04UMbeHqAy+Fa459TedZmTO8q2IRTIUEQG1SRAWY1m+E+F5d9b2S0Tzz/JV51E
2XD7k0tmmczu8uFsBSyTSVZWnsMi1fc7etsZfyDfqOPdZjJkzcruqQhd9GpQxZ6Z
v1uRRMJ68zrof3/lfsUHnJ9gOxF6q2K/Hkh345C0Wx+xVuSFqQ60EVGdfyO9P8Th
Jxa5RXhrjKu6T2J1wAWCV5Zr2L40sNqk7Y6VqkkS7SQJce2IXr0ybChE8FXDb5VI
wSmTxziD0pluLUIJUYYV148i7nPvK9Aeqkfvys9P6XioTBGBdl1XzFmx5bKX/jLX
2IEYRmzX7lRRvgelvymOFUM5OPdTGkSfsmmcyNWVBu6x/h7bDyloZ8zMU/AXg4Ey
SeBTZdkLjkWTsB12sNOgVCryfvEU3ZLsrZavuZJ1cgquhyu4v3qJGk/PqHt+JDGL
jL/MyPo1K1rIfwpStOq9A1bMKKqP1ESTyfs+0KtiERNdK+HSrCBLdCxeN1aAVPlQ
hIGXr4rUr72fGFS5lrqUWakLhIVWYjKEMpia39T28NSQnkeQLrRfjDKS66a3GJEA
Q0tm5SUk98F77reP6Eq5jshjwg3I/0KWftgepAe4YvaN/QweKqzH3TfTqSyqCi9J
23U8sdHMLjRNvc58/kMYJw5XP84m644kI/baNZLlNa0CIezCQnvk5GDoS4oKqip5
gk/gpzZheIPzkNQxckuU2e6TkfbhTBStmOMocX3c53RxJ6LWpwDnrGJYcCqZY+/B
sMdWXrr3B7xO9SsclvGyeKIMctBrsGnAyLvorMbP6ZCmo93/3Sz0UTEa9PNVVb8o
aTGYr33Ej6VHwxKN4khVXdHNCpf/gTit+PNSAYsNvzo9GuJMPbWxUnWq7oS5JF5u
bmkiC/1HhzZkko8EaJGLgaSpbwR6evaJHgXyqZ7gToUhvl1hLVWliepFbEBi4mKZ
AK4JoTp2TX8O6VrIBKYWVp9wiN6aEKFRH73yzuZQLCz3WgciDC4/DHIefQft8TX6
ULI4M2Bgo/OlPo8sVQLVe0kuYF7c1HX+/VHNBzZnRl0YHI/H8q8HCcqslxD9t4hf
fp2X91RKb9SQyzA8JUFMFnFOMMrMz1WC4Rxc/NWAharC7R9+RwAzYjoG+ZAoaF9Q
NTy9+XPT1f4mtYt9yvbmz390VO8C8azxoUlmWgW4PTEYLo3Z5jH40grRuJZqi9/C
vJJPcOSYqytULu8nwWf4Uh5grBx+7atGEYIcSGRJhO5pWMtgXoGo5r06ouXOFriu
o3/3OuW99crmKMyqv1fOLkV7nD+scA0mm+Trvsu0ArKAd1RwQw/nJWO+JgKEDAQI
qin0om+GAuXlE8KwRJD5qLLqWI7wvWv9a1yYK/+va5c8E+ZqGw1SekaNOXooNbQ9
ByswDRBvoD1vJ7f9tGBZ7YFGkuIYi1IBE2M5+Mikhs3nZILT4LYcXdRoz59DLiwg
3XA1Bq6Ae2ti/fOoGPI8rVnQJ4Oq5MkD3Xqx0yqYckuGhfGW6uMCj6y4f6C4NVYn
idCDsGgFhn/E/of58tOTrjvWl9zOSi+sXvNhi2YwucNQ3dd250rbplYIa4FtPlG7
TbNXzosFMFbKD6Z5qeNdvBpGQiSLeDOATWbGBmjA2Sb6+DUVmfQ+iifE0DMEucXG
V72VY0letTGo1duFuLNp7agKtxY1kvGqKVMJzXXq96T13nRcOEKQbw1M6IRax5V+
LA4cfjh8K4DO6MuML9liuqQJhZkr4bJL85mHsxYjY3p040zaDuK0kB4N7RUqhlyc
9YeLRCtP0fAK+ZNrsFzJAf32Tvv8HO4CNBJWH7lQfOSARY9naGUJopFhGODi6G7G
KT4Aezyr5ZRwCHjmYz8ardl9fjTQFo7AzThpBpuoczUQf2vOiQfq+ne4qEQVfVEI
BnS05TANrYY3qNUaLcQyp/sDCs+nRkNvzqV5K2qINL3kcKdPGiIdmzvckOYYjLrL
Leb2AM9ss4Xo8RkfjVQoSk2dLDu95/EjsraIXgE0cTiwh63BH+enMzSyacQkPrsS
j9Gtz255JmTVvYDVaj5JhZeOzP2jO6qOfkFSDHl9Hr7pfLQk9bQnbg3XRaceZX8I
PB4xayXhHVIhFkcRU5uyIl5XWbxQoggLmoI0eDtyIUMz9iPOfqNu1vZ1cQDmwf6Q
Pq8aiITDjILKtC6flL2N6celGqLAlO7m+3llBVjXsm2WatjxCWD86JCqVN3ww6MR
DqzQKOcschyw/h7AAMZxNZk757kZKYOxbjFZ0kcufjx0RqsuBz7/iACE8A1b6MpV
5CaW53R1EwX9HK0f2Oh3eTaXZr02h/FT7+oaWuTk7kEV8vEVylEc4wxiSxJv3NnY
u7wUroJHvPOiEAIX0AOJ1i3UGShRW+4oNCStiVDKwD9tgaEwDDFGqNZdR7aeOWU1
tMdGigfazK13alg92OahOpvcGJLhwttzuAN40TdUCKIBIURHfP0v9o1ofNh+iDSE
J64jJqUCl2JH2kx4dQ4yVIf7gpwza25hvrNZNBnOBdFaTLbLeYsNiB1cM78BflhW
Pv0sIz8uHHjweGQIMJBJyhWlYiHahAvA2vboATbM3VQJPzzGLRY5wVN5CNLq8HiZ
zCAMU7VeMdsGJKUdQFERQ7oIWpIs/SI4yW2jegESrezlT+IumjUFuCp5MLdod6FT
xW7Hd6VHOp4bn0rHc9wsxDrUHkUnR2c1m8EmPAG+6AEkJtliDhSepwilia8guHnV
Wcu9v1XRGbEOA+D/M5CINCKiFmMw3dYBy1ClRc/XOGJwArgj5STqynMYZKMAQSOT
Aqgge0Dxf64l5Q3J0Or1MoHjO9/qmg8Y+kXP47ElLCLvCDhsfSWWG5WEVUG9qYpm
InJBHOWy4sbBitNsSVXl/N6mVGvwZsCi1lyHXwh/87Kp1xFinQBt+xAzuoOvXY6R
/CSZdYmxj1HXxp4ntQ//GtA8qsiWl1spwrSsZQE331NQAtVD0tMcgDbL/Si5lcK6
NIPocOTqOMlNLkROz7DjwBmVm31Sw4nAFOLaVOga8mk1nmBPO2cwV/kAepnR2cxK
/H46+3QyBOEmZYMT47uK/A/VLrUD/zpeToizzYdu0cH4qjOdgy/xIkX+D8QZzaEE
MD7uCD6FaOEfg2Ga6J5fXpIudlKZLzdjXUrm1qSVGNm/5nivLwLmYUeBASX1ek7r
oQGxikejtSGSFyvjxvVIin3vLTuhuWcBsmRWErfRABbBz2ZGwejCV2L773xTwqPM
UQw12We6rQp20XD+uNvLRMTkNriI23dHJIbMe829FWqBpu7MYfD/9cJ27pTbazBl
FMaewiqH7Qw9BrOVIdZpH4utlejGeA8t+y5Q3qvqQVvrnPJsUfcrJbaMneGcbZ3W
JsYjPWIvqiO8LjUpysoxCJt7sbqc9T3+yJIPm14ybCgHsZ8/sHscPRtBL2Qjz1K2
M8BV7h+T09yNpxCnaIgjsLn/dwgieMnd/iu2KXE3+7oPJqKulL0kIPYzl+reyAdo
1COpoopyEl+hWvl7txPcqWAe0peJ7Z5CTnWSek/KTNks5tUj+U9Q+pSHWrtOZZ9I
LAt9mSAuEfABYgJFfLODGgfzOt2n1CmmsQHkJ0HnZTAu+mew9i6R4Vat7/Y3OlYy
akLGEvMbhaEdRjUh4+exOJk+iWa3Q0xPUx8RAGA4rD0quxuvwXCf/i3b/KGBeQok
Exu2BVsivMH2j5aEvb6dNWQtNGWi81/OMTI1TjDn+ryDKAFCpJbb33B0eEeT7+ZE
INlTb/61vlRWOAHMk/VTCNb80I0rP3/s8/MWnp9Ad5NsLVFBPgM9irtOMJWONiur
PLsFwGukuWr+WI3U8mnUSh+SlNsOsOfuW4IUmi1ftKvkyQIQsIr3lK4M5VBdz54d
NOI+uN6w7hHeMjixTF+0aVGKM/aKPC2sWLspc/HkCyhDzugGiGaAeeY6Oq3QGFF+
afKUgeJbVOYgZ1lyanUDNPWBQfUol6fD4pkyPeQKL0/hwmH29vI/Z1OgtcF+a4+Q
pndWfEbsAaO2eZG8swge4UnipzX3kejJs4awb/hXuFgjgBeHXknRvRSdylBfZS0U
Q9xmKG7m+HpGv6ZSlx+5/RJcjTVILjT2ILbgrybnoBEIsPOm5l76knCc4Rh+HHwQ
YKHvxYgiCFsPwfaLqct3HfTXHWTBrX4EW0DM0OdxrccW4n3IbzzkCe8P1Gt/75Cs
feYf4a0bGvgycwET4hiSCDBKzrtpWiNgq6PFSsug4D1sizQCSX07zk4j98uAQrwc
PpOduOm+8vgisot59ScCzYcGfnQoP5ElgSkaQzI6aULQBasS3mBZjjcPhelvvpsd
bttG2YPVD46VR9nvxbsR9xVsfSRxYldiO3a8DNWMRK7H3YaVUIRYKjVFTSejjf9+
DgrpKZH4pv63e81jv/ahkt6NJN5zaFwGa2VraB+CphlTIAwLFWyxlB3tmBriFaFu
sE1xFC4rxL4LXNQMYFCYAb3Wx+hpuKUcpp3QAwozRRbr2gn0GNLVBuCPNGJ3DYca
sZkMrZXgf74RiwudupyTooAiPVsQK7iQL/CaAlnZUExhQDyIBGNo/Wj3h1PChh6Z
oZT1j0yn+2jMRfmuty/SESF2Uw7CtxEU+H/pgCbZuW52fbfzvxQ3diT1OaT95BZx
y0aNMucYDsgKpXAHBrSs3K89820TGsQpjUJuHUNS9KyBsM0rxoOBsSTeSTaPDWDE
hhm+nEPKSGkG1nHkQaS2rFZ/5GDRF0ZNswHIkSR2bK9jvuuKDgTkqZGTcdqnt/GF
2rCyD92PBm33mkluc+fRFPOcPYxbCFpjsusG8nvahFG0mvm7NrxtGd03OQRrzvUv
bfrfvOtlz11dLl4ha75EEeIK2g+0ynEIxUcCQwbGue/tsEtiAa2iH2RpbLcY2qvk
YQipYqxczOhW6p8SFOGKUs5r4BPIkcimIxlbVrWN+gQ=
`protect END_PROTECTED
