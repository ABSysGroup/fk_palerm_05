`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T4HjcxjmLtMP0ZyxCDy3MWWcAAqsLYF00l0PZAbFEZtM3SjOAIesFZUVvBOrDat3
gwywPCES5iZ16hN8XkvBnY3ZMp9U6QUqf6Yocbeicr+OknR3Y2cAutUzOGTvDlaa
F7mcK83G23d2PuldcRsPMuTg9o2lQ4Tz14bQDwKz1TniKNJ4BuYb+RLmjOQF4AUo
FLvHiXScF9hJEYAwXsL86eFmdnH48ww4ADnRB7SXhivck5Ka0n8DsDEFnmuyXgoA
DxdApchyU3oFkLZlWx3LpwOZ5NOtZme7tt6P59vEfhRN5BKxtLojiRzUEYJnpicv
UHAK5La7xEgx4o4wzlrOyURLZzJm/Mivz0pvw/DQpLaEf9tY6Qa0uIMb7c8a9jUJ
dOvxPQE9Jb5bkfoVSGq4ZV+51OD5EFbpDnFcYut8uy8MFPSR+vO6GvUEVWTG0bT/
`protect END_PROTECTED
