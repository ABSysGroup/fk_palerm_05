`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T9htB/89daxJ0AToin5objwTHWmFNB5/P1OtKI7+sRizjJ6ymHzEHmvAr+AlN8CA
YOgQ/5DQqFA+H9v58MiMJBSAqOvjugina9LDnLXx5r5YFHdKW0nsc4GE5OO3iwgN
PUtjDW52F4oMGHFCN7x0I8da4LG1uC1GOzS8ShjbnhCfI2jlYfpUcqMfhrCLrbRE
vbW860VENgWgn3j8W1oQ42MTp954Ki7RbFBPneli7ti83mdYzGwmYYIgnCmnBKVO
hE11S0HkwgPMii4SSVlffW/r5Tagv06lsT7gvOawN0Yv7lyVJOnLi5i6PqYPwTuJ
DfN9kMoZe+Kcw2708pzyWwNFY5sdBIQHwP5Vkdyv5RiuKVC50v6KlluuqkKPCXwN
nbofPb+ir5JsmGJNjPQpcsjwfBdVfnEngyzCzTfjoXBhWq3N+wONX+Gj/gLX4/mz
xDOSI8Pvqc/EjJ1dXBOfD41umRtzYWT0hg4nAyLNtiDTAToynDT8lfEUk+Vl2OKc
u2pgpK3mCtk1XN0AZ/ZbJorCXOsD6fbWOXLGA/gEpSirSgqsArjSnD/T8fCAY8Dw
iSd1EhcKEofKlDmGE18g8A8wfaIj7dd3+hOf8J4LQPQiCTMcknNlINTk32Sm4a++
VFFuxM6McwVeMS0fKY+tzw==
`protect END_PROTECTED
