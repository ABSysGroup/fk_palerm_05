`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fDOBZEj85wQ9ysgPh2tiHfVGnkRzK5i+3v98sCKPhK09Zh6Ejt2yeCR0d0nyUSei
Wgr8dQSbweMSVitqsq/E+eOqgqwKQr95PfDNxHY9Y5QeuR19oSjxGUfvtj4czNkb
ctZgeNUXoannapyO9JxODln2NT87ILYVLn8Y8tSk33o+a3XQzK1Zrpr+1wzatDE2
pDFpiyHaLqDs0ydcjTCvSNIjmypcBF720Rd6ugZLptWuUNDa9wzxkLqLTOqzWKI1
KSuARONzdpfeTHhHUTURyJ6zRpDxEwvWINtUlitodogOWkpCbEi61ruIwZdwPnWQ
DHMJXKtxuv8tQJHsEoaFfbnB7AwfySo8W1fEt8FjfGmm8uQOgzGwZUSAbA1Yq5iG
Fo5qqE0WA+3zAliUcnRKM53rpyKY0RJ207XloeYHLNAIZZ6mxmBEXY/uu40qvy+y
881rZch6CLqK7fHzUyN9VNUzaJKf4KjYJwAocjkuQ3K02hyeCXbn0e1UY/Mm2/v9
uMU66vkYMCZc8MUGIAZ+Qv/fX3DZ7diz8ri9ZQxkCFhUAUK0ZAl3PEq0c73l4h1b
`protect END_PROTECTED
