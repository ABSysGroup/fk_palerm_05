`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S+dtbuPefOgx1iRtCo9wIv92wwrZcWjVcd0GVnjB3hRG1gTsnNgK3RXIFvit7GwY
rmW6zgL7NnHD5uiA98aMoUgsU15ABXGuqqR2dHWbrTa1wisbsPzqyUBpLHiHJIXT
sa9OD4SLa9n/26RTlM6eB+5tzxVJ6LTufE2vW1oEUUOhgWr60dlc4nV4M5ttJxtf
HLEpVvi6lBxFmhr48VH3zx7xYFssZ2bL+bt8uoNqbtmoY6RoTD9jBifcZ8RT5Nr5
fqdPktu7yI1ZtVAbH+I7dI1dXUhGJDT5svwGP2NbXWYOy6KrzUIbPtw1onDIjaS2
jGJoYDWY4hs+FVgco/murmLUzaczRCuMy3cM9lgBDsppkh95GBv7XI2VRwHXhODn
qvXoyhjOnhB3aItpMnRIzfpaGt2ei5nVfW5f45g/VPWxnZpg3zCJ22Bn+Iu7xpyO
xg8xg5VPkSFFuHrutv7eFwbxp4Fvw+6WdWIZ8/c7xEXp+bPPOwt/tzwrL0VeOMgp
U5913GdPhSHuFzSQMWYrTYQmOG03dyKHlS/qYoELrE95sgiHtcoZY0lpxe3MHWMv
Qf5XO2PhyZIBCtnCziMhSKZNKF5Gs2aIX5GCE3WhtN7xaAmHc+rf0xOl4W1uF9Jh
hVkALa+W/AzV5XqIOgwAW20K3eiQVxO5MhGLSl6Uh+pbf5FpKS+WD9eL80HS+HNf
CvKzhASQ4rIZYeIbasrfccu1riWQljQbIAsIiKCE12Y=
`protect END_PROTECTED
