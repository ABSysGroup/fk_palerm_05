`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MGJg9dvJ5JPVWpKXzoQZpm9wRXO9VBAh7YA7PAXpDIjOsgqtxGYGvRU7zSiJnzAS
DY/8simP3X+ic0K1ciS0Ya1dH8YZ6ECUf1KCZK71diIRfeL4ESa5Y+g8BCg7DF9O
lsNXybhr1M4bhomEl5pVljC17Z44kzXwUJc8VF7KYeZKyFGOQvV5hR4AHFCVA/dh
TvD1lqAIWn5iDSWZ2lnzmRCtCSAD/UlAumvZ0wYJBwuYljMhG27QHn2EeezEyFVy
U3HAllUmunTL1Aoik9mduEWLA4owfJ+QDqHsfjz7yFptXTb5UWJu4d79RVPJHcn2
cSvMH4bXXiiTK+fRLKVWzx2gwTvwCvvMZZlMNkSyMUhyH2olKlkuyx4hzNdIyggz
S/vk+NgDuUpdRzCSrTGs4NyozuCIKGqfg/x4ytQffPL67MZOXv5sr3IAmj0bv5o5
UqKKVfxj/TjxQTepdjRbjysIuM75JhfCce1KS6cA0VectpBtsZbO+r9nrSOvwZPI
clWMv/fbXXEIH7Ro9Un+7qH7PZrw0lDg9D2M9LI6WqTJSFsUibqG5a8GwRAib+Tt
hIm0sYfnA6RcG1GOVCxsBVDPIHP9087Y7mMR4mOV+ldYs8ypIWZfYGOPZFFkkWf6
QPQtAxBsfzCWMqHXp5+8dxUZGFBDvLIEqEU8sFIsYQza1gASAPRtd4gqLAbDU7KS
0b3EllAjOGNMZgQd1F1ReT90WRTFRtmpisfXKBDbxhnwdgFIMGookY/EowGyPL0R
yaxmhDBBsxCiJrix8lzaiG1/ncu2ty2GeQ5vjD9braxoFaIH0jIHW8DywGhfN/th
gU1guPzaDGFRiv3noq7/dFJrg4SZUeEPhdximGhPlEERhKeobgg/CX+2qzbHxr0l
RzIbUuEI/sSPFDYLJUzJEAnuexxuDq6NlBX0RO/WKrNxQ91Y8KNItuhLCp8jcIOc
GnL22vev9zQego6ybJhZUoRsml4cF1VC0+3rMcsRoJsDlppo6Qd+xjKVhiaOw63x
`protect END_PROTECTED
