`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o2ah9+60bBH0Ggr6+JLoGSMKjWOVbzwHMQSub3gyAljx/jrDBBv2HoDtqtx0PPha
RxbOqm6PC+opLsOTXAZqEophZxi+0bVTTWZn60eOWWR88pT+gVHaqYHGDxP8Sd14
WmOKMd2oG0/2pNHocZv5ktZKqcFu5NBAuI9iy8xhn3ijhV9RCr1IRSmDFXGMobxP
hor76q+LZv3m772/5XfUm0XBZhdBlY1LcQNF7HdttWMbxElD7xdvGxLPsg4pkYdi
9vdr3lN7wdTfszzdF9Hlhg==
`protect END_PROTECTED
