`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yhfxQQmlTOStygd/l21BHorPV9mSO6ZK24+RduHVUqxmFjV7iqyWAlwR1PtZf2tB
R81mmy+JvzE8u7MtwrsF4PU62fNOWdfceh8v04JPvIyMRnUmdlaciKAH/ak6NCax
XBWaf8yyvjZS0HCvy3Kw5z+KYjG30cMAeXjWBLEejziD1RBOkXSS0ZaoeaRrC3mj
4S3E3/At3KxlpaYq6xGlGlVlC43lOFrB4fWfYcVsium9U6k0MEfQHygI3mgvr0XO
JQtOM9jfoAu5RNCeGpS7QTvva/Mli1Ff12yUgfNAnzJ7lijrWBjKVbk6/0z9mDP2
jjiY1OO1Y6SXUCDdQdUhtd/fryrZyQfnaBn6FkxlSZqgOxQXBokFcuhTNum9qAeO
gcQWkoHtsDhqvceDu/urcPuEnJwhTDiXgKTBY/HsZdvDlYHqa0d7c075n8IIWxRW
fsSVkOiru2WLn3//Uzy0RG85llBgXz8e9Ya4+RFrXZ48KoU8Tg2A1GBpQtJLhJ2R
akycENQyVhL3bNL3W6bY+PYfWpzQDk5VoJuyrwKk/iT/FoIqiUdxdC1RYYpHxDxI
wScholmuC0nR0S43TZva61N6fxCZeTlRsIMxtWTXkcpZ+KhXdDCNfrmkE0/VM8ZR
+X80PSn7uAag6Fafro1EuLfYVXvRCHc1mA2gnMXWCM+uSJeuXurreKjiz2kbT3Vy
+EtwN+CupbTZbci1geSig/mWMOp99I8yLJUYEg3Sjevh8KITUuioYIJJudwa/8CN
hnDVFlatpPWQnU++1XeyNsg60Y3X3IKEzpmhr+B1Vot3lEeEJ9CGfJgFPKVPIQVf
mVNbTu6dThVupzKr7Sk04hPDtrbwgId4vC1naCPhYHIFYzG/Euwuz6IYYxBSztGC
5KazXPjMru8Q7pizrC7y3mfPL/Wvpk5Y61tBWcmzP9mRf/JRRN5+7iMmJAPSihvi
zjDLgVK3wTdTr29wPJLnLwvU7jKS77zKel2HHcz2Na8JfK7RU7rt66bVZfIo6QWh
H8FrI3PzpQKhGXISlI/n2JE7EJivGaOkRSSZktfttTxWlmEYSkCKRByw95hZ4D2I
4bFr7t6klg6nc+L4cS87HH1DzSMKdPvIv53tEq+vrI1iDmCX1OqvaVdMfND4FNgl
Tn9MuysDaN7baAgln4uXsz7OmhfsnMH/ZKe+WsBEgTM8Sd5ynC5PZovYjneoNijY
bobeE6y86hH0JRzSH2qB/ytHwdiHQ0k4dYKLOpFdCupEHwXhTexwXwlNQ2rm+R0n
ljRivHsLPGlFdjOhK/8o6g==
`protect END_PROTECTED
