`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j3qHkDXFIXf2yk5ltSi4hb3a46L+N24+HgYBeKoquHsXj1IDBOXbva/njTrsOxC2
u4cA/hRKMzT+Vw+LLfoLjwpxksIotN+eAQ/aTp0lXSu9khBfceSf/xX0U0d1Wd2Q
okI5x2EwH0pC2yplcCYQeNBMXm916O1fojWvid9GYb03/ZIQawiWLk1DOAMWByQU
O7OcTqj32PNpNVcjI5+hCWOW4RWalHDPJp9nNbzqzj//kLEy8dbInUkok5vA2C/C
zf5/eRXRu61bmOFppOOoCbEPvnG6YN+GgnjH1tvGeXt9OsnldObzEXD6FGbR3cgg
pJqt0Y6zbFU+D4xOloHz4WKYydi+jwvFXIku8y/J3cpUs//mUjnzdKsU8G1kRFT7
OMDHZE/gkqlqGR6OO5NVp/N1kN0GI/nVRXrhfryXQlWcIU32j8h6im6/0eqJrMpu
OKTS9HEhZP5Njc/m+Ojhccal9JcY85uqqOOM3rj3V4ovJ7CR3rd2w63SyEx9Vhet
U9feNPu5U51OMhqj7yLMpeQl2/SNIzZ7wxuNlj6ZLBKpLGOqZNWOpzJGYURfpBFS
NEWYVJVXGANB1YH8v/q3NDWyVxh1fvDgX3k/Kq7qm/EQg8qGlJpuaHwFvgaRd/Os
P+scXr+2Fwguaeq4RqQeZNtHiEr84i/hvarVxiLYGkT0x4QEsfVdbf4BZPghZ5ma
/AuvqQViSmmkfRTdxn8wLgz0yYu38eHyh+mzuRMvQP0kd/OFZkptuB0rRcH36s1H
BNKij5LFRPa5GlkZrEexYw==
`protect END_PROTECTED
