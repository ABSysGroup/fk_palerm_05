`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jmjejROIjZIuSJ+07O48tEJpa869FdjLctDkXbttYSHWN6qoOF74TeEiZhBt4bRh
bQNl3XQokg3ZrflDLWjsIyAYJySfirI2lYik6EbuM4fVJQY8eFYh+k02WUW7x0o6
JnxUUD2Gqqg3t2PeV2D8awHMW5Sh04O6Z/nkdYUtQ6PLWeGQpwqUzO0au3Rn+Uy9
GV/+Ic8HS+uUGx/P1VDZ6yIY3AQSaDehL+ADV2CP8f/3JdtgVOh0Xz0S/eety3f9
RFryRLmY8Z+FikR9e+ABeaaL0J5Ab9ivMx5m2iExMlwGvXImuYnk5dbPXtqUDZoh
x9x16z2kkiE5xc2iy1oUZP+EIT2VgyKDOXHbFcyosu05wh2YkYX56d6Lp+4ctX12
9W2S0Ld3Lq5nC1RwQbGn/oCkJmfEa6uxvF8xeRhzx22W/RdtZJRDvMchR7KDQ7sz
rYutcej4b7OBqVoELuJFn7KV90SB9NJdJnKOmgBM+WqhsLaV2ZTXTNtaflFrdP7O
J2eWvfD7J3G1dNX7B7bQK5fk9AS79ASGrvfl7n7j0DBBnMReFGkcS93r4oTb6FJF
wJBAbmLR6tOnQJ0P1Jl1i8yZ+jU3QNKTAqgqgKdsbhcY44f4uUv7XHXxgQFIeaAB
l1MbcDPNsFjjG7axaE9UYHK423N5rGTgk8KQzuniWECgeTa12Yl+ZoCC9ZYL8m0Q
11W0gVQ80j+QxptB1xdyq750h+kIh4x3vegFAvbinMooP3/8GgR4fxf1HG7+WZB5
iMacfhSVdRrOnRVbQBp1O4QbzK9kK9PX8noUm4dnhYufwk255G4CGZlwWmTESwYU
oD46yIsU/VMDEuCbMXswjghRHoPUaOO+OSKt44T+sszj6NMc/n+3czm+mwh/DZWV
eP61BP4UbOfhQGFL4tdL5ujTMoxPQTQRXgu1evdIPJPpECngzCf7EE3jcM+J4B44
5gGpBzmrfxkBzxcRpDaDv4GhufgkCIuR2/KlGt9KIyTfLtmW+9faFzDiYdzA7lal
cfwVrBe7jUGJLzkxVOh+ctg89+SfxbNoZk+L5X4czTUdfBW4gmrcBSOjHhn/2IZE
s1Sz0fnpPLpd/7j/evGennwXsrl1q9vGRlRMYBygKdytpDVtPsVIVCmr9kkkEEij
q1wHNPvbG7gyisH26awYVsoYYWnv//TipWuwpe2ZTWqv04ac/8cjZe/mV40JSAyf
WsG17tCf+o5SnBMpWZk29ie+c76SVjs8abDEEVD6tqJZRG+qEvmBnZFNHL96wY4y
PuQp0oI8hIhS208VO1jJHRjSeDmDBOGxk5S+IpJGOd6R6W82kgqQveZ3DOHDx6wf
3q8u17R1nQWe2yiel5e6JcWCVqBz53C21dSLi6mQGJcg4nYPXb3qYN5EZB2j8NMd
lI0FIr1hX6p+4SS6+GF4S2BhCZcsrwum7/R891bSepgxpK8ycUJ5Upyxf3Cy1TAh
J1sq0miGxWvUPqORPOXw7CVOIpIVphcc0K6x1N3DNvjFhbKF63TTSIwAfA+wiVcK
hR60Cet8X+9GVZFVC1UMhVxi3rHoJgS3cBdr/cTmfRMlnSbzTwtnJP+NBJwfmVO1
hf8E/AMiNmo+uPF9kvRW5rw1NiJcd/XBpShDaTcK/u3HJsRCni51IZMV5YKBovyF
6hKJQZdnHF81DRMXWQU2H/KVzNwCrNeI0Txhh0r5IS60IgcFTBEhzHpoGJXAUXzK
GDnK6eTkIxuRf5EyENcXpSunbr1dVDSdIDDe/0AqQHbZ3vVNizXi0ypP6hCduMO6
Y2bCenBMpDNoyYgn2AVLiPPAECqWenUiO56hEI3c3xladUV6qFgOzNYv5WIkOxEp
FwdVVO2GZzhc1N9J0qOBv9Nn3b3FMIlKtyAGoPTWnw7Wv02Mm1aNQzL0Gn/2yuMH
2uBsuxW8+ModbjGY6Ziao3rF3piV1wesphgOaUfHg0jAk6cgpUDruHIisylxKTJV
XT9m2pu2o7u/MsKEhfziWw8GxVylJHpwaSFM9/cjcDt02hRbMPZRo5SylsF+zIxt
a77xpb0XwExtDv8j9Ql1T1rd3kaylwXQj/RGNhrWJ2NdF2CNKdITnJlSQ+33j07J
nkk+LgBxTtDn9ozf0Y31xrOIfO1u82o48SRIoUyGiz4FIxoX7txWoIaJa5aySzZw
ho+f5KB9U3/c2SKcqzcBCn3fOgd0ZTSTz5UinCQgUK2/i1QeQ/IjNKzdqrZ8ZeTc
a5CGz9Q2gJO5/fNkB6p8Y6fVlyzzCfp3KzuLpWjTJ0b3MV9my2hZ0u1OoEMF8xiO
neBMRJe3XFOOgBCpedXDYwN2Xlb8UdrhEHfml7CPYqSB66pjxC5KlfxagWqkQ5Py
tvJPhQbb/PINJ8rgpThqM7eAKuuG4l/MMlZt50qkHLJ/e4cfkcyQv5veagO9fm9l
ex6aGgzUy7A/0gx/gQ9Tjhqwo3DBXtARJIhBOZtrDOR4EctMEXdX3a7890AB83b1
uFWeiTbVHC88rKQG0a+nhYdHpiLM0z+qpkrSQqjn5u9N1lqQA2813rBU5Kp7UVIl
cvbJFVeeqlrZhgjq/RXrAIRnTpnH/nFFyBaKRPS5kUAY+O3JictIWolPPP0Lw/pE
t/6WBQ1CucZL/dLmziFLctAK5YtL3n4zdYhqSRczsMYFQZegrwj0ZzU5iQkbVKvg
U86ZZng2beaDfhXZ6ixpZXxcJMJowoPoEKrrbbo/jtInX61dS+Lv7oK7qIeq4QO2
5PBIeUeFtifK0CzK/ydYXwZ2kLwRIkWVvfTEdPRe/sUT9fX7P8SOWLXjIv5WE3hb
99NDdAYxhqRDPxUMcANTvq9qZ0FgjJt5m/8ycihGUn6DD/liNKCQ5TbvOZuxt3sU
J9B8pIsBujDsVJ5UfHKBPU4XBCUV7vSWa+NpoS+CY3pvc8KrpLM+i37Pe5SByrnT
MsIKnzKv86IL8gx96mZzU3YSWKvLwFenFdA8AZu3sE7/7EBZXM5dHNbb3SZdIqd3
yOIA5wGbTAGFcZZH9yWs+BqJSoW/XP2AvMU6V8aLZyhyBdsQGD54t8KKXjTxyKr7
YDq3RK4CBzIuYKpW6moDVMTaCnvJQmL6kyEqXHwKOo/oq5PKJIj4xSBOZIfwOcto
DhnzEbD2rhXEq2ATgtKYoQjgOhaa9JlEHMzBBsb6TK+gs+M+xtXJKaGWmvdAP3LF
xQMl5W8T3FjjzwtI1i0KF0LVcxHxx3PtRELnopBt2iZtMPDEUSizCZVgjxXPLjzD
nIhhQIOxKoho2HB1+bnsGmhEiS8RriDMT5zSojUhXTFigtekKYhRFxXZ5lItEdqo
e/NVtiXX5f2tePOLXUhE91uKIu4dZFKRjK98pCFhNcrNg5XfS1j350TLIesIHmxz
XLybctw+EwRu5i5gxxN4qGBS6/Y6bjhX+NFM60b/lG2OcC998C50J2Kt+EL63klM
lf1n7GLdgXi3Gw8VQDtL9Sivwzv8cEfb01BhKVbuX7oA5z3eKjq6TddD/twUIhBD
jCU1CY4aNfAJA3pVyN4Lt2RIg+NUTPjEW2gz1H19N6UWaOFtCjoxHHlaLz8idpfc
GKUCyeDBR/KgU6u6TNCkSiSnhcn/qjPm8VuOkihUtmT0/ZUIMb26YL6e2qHjCRP9
JwyLIZL3d0QiHiOQ4i059i617H+4R12CfSsTvT2uycynJBQ3tWCDPbmToZX0Re5L
N5Pk/xj+Z9jJIH2sOXwfMpNDrusMqdwzQL4yMHF5+68FmdjwweV4Q7129npW4Ufz
eSA0AELuhf6gV6pqogtUB0OabnTG022FG7Y9vVdQNSWwXVCVzVy7H3wqUWMkcTeR
La2hf4Q/AjVqzONuEBkAuHjlW08NxC2yc8imCHwfw/LxGPY9UJZqpWUWRPGKc60m
ujGRPvjtsW0dWjq8gWXjKr6A1FC+LSa6Gjhc5ytWYQRU3yZtNgv6JcT7qLFJWm9G
8syFngrNTvzAwuZwnLbvYXSj4j4A8P2HFgy1ZcBiHGXv4uA9J9P/ZGd440Bl+Egd
Z52Xo0LZ7pp3wFfsbqA+sljet+aJ+UhxShB0qitumZZsIcqswNMal/PA1XpfS4Ei
pAV5meh4VQQLLb3jX+O8m7BSb5EA1ItojwPKLgcZ1K2zrDI6Z0nhTvo9ydg+tDHI
fqZomVNaplHfrpk40OurycqqciPln7TWKC+SFoTf2GQ=
`protect END_PROTECTED
