`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
biRjLejnSUNK2QCEQcuh7z3ZX8o/5N0tALEyBqnqYydCVcje0ulMhxqCBeh6WKZq
abcOS7UXdqyyJjKbJi2lzmztqAR6+ADYaY1Eqy8P5MUDDmDGLb2CLGs/abis0Dq4
0XZTLNY84+kH2FAuuXLJdMXQyakIH1EVipIr46VyafYBoVvzv7mF+CxSHGc60gHc
EoZvoruAHpmpWpY3IrR3Cn2MfJ1p36+augLwsYSEExhM03TAe8SWjJUZlZ5IMH5/
yylUQ/WWUIljr2vtdbj4E0BHaLcE0QkRlRcxpM3OcT7Gz74x+PEvvblNu7MkZWaI
T7+d0Z8x3Yt/8Kicqu2BSrqe+aF+LYDDWb+49RLH8Py/Y5GQc5SYl3mHrvBGFcDV
pulWBYWL+aampnFqa2mApDQpAqdB8jCA3gYzCb6wpwzG10MwVmhxkQVqOZBjYa8/
Dqb5q8GQpjQZUdeH39g+SuKnjNp5TzqZY8MQfcnwQr6vx2rtqMOXo46dg+nx0BB8
w/mdtfUx7YaiRdYVqZbiHn+7bRaVVM4IB/eVAmJtrlqoTyexzfQ6bQkg8fYvbV88
42/jbGYewU7cIGcgz9a24BpDZDdWG5e5jWnKEZ3XTzANE3XB567LZkNCA+VdRnIG
/G66daqgIWulkGwglv2OgLaGR+1NX1HfxTgy1JqpmTojY5ValSri3/JJcLPWHlba
6frHXWt9y1mqg42nCLLtePcjK3dSG0TRvY1mjmSv082wJ9IZz0jYQp2Rednw7PfQ
e3Afxe/8M2l0ASVDuht6raBHRBoDJPrmtxpceiEkeem3e+0EYtOYU2bANTQ6XL86
/xBqeimL6/p6BgwtnkrgNPqEqErlAa6i0ZVzmIsiERsnmkWFqBJn4JvZA5NgG/Lw
f2ohZP7QvthX4i3kX0RdiQ==
`protect END_PROTECTED
