`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SwUBGJFcrlsuxEDJynmU0qnlR0d8H6ZCAiNZ2Aj7p2EG4GxoUDMvfTL2lultvtuy
ND3KhLHB+ziH0AyDMhwjLCm7H9GFIZiSnIgEoDifIxm1PqmpLkzmJLDcvJh0ADLE
H42sgCHso3K3kVm2vLD7BYS2rIdzWu4OXAhaEHnUU8OKAIHsZ3V4ktVxqrAztS8S
qZ/hg3LhaQnhTZXRxjmdg9GJZYjhxadvZUdKN1+dNYDG9A5TA1oarCJ8xHDwtQQ4
yc9ESJHLzi2tDp6N1t126g==
`protect END_PROTECTED
