`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ySfxTtEvLsne7tFkuT+qFIpmJduHHBgmMrZSpJKsT5WOdLU1EaF89iuVqmVpaTJa
2d8gRH9izcM04WCT5vN4nZj7CC9J59Ma2o1B4W4+TcGjdb9ZQxfgZXaoxGezkyRi
bDWjRnqpLU2L8gnBUzHmNpqYrIfa279wgda9PrWXQvARO7yJW98vsW9n5m2uQh1T
FzoqYi0bng/9BvR9FHTZ+M96sizn++w5OSAKsFyLgx1ztKBXbscDTFqh4qyKM9DX
5ZGfUVdEaOWrYlmGF2L/8fdngObtjc7yCvaCgrsscw1DvFpWmP011lEEh8zaIcFC
LBoS6wFXgJBODPXXVZGxSpDZMFIb9CX+pJF3khJbpRz0gXB4ja2QwXB3xirVjzgm
S2nX8Fufwi9Ii2DKpZxWKKHb8JIhgsPxyxdBY9lNJqfgiR70VEjR7AlAgPpwnHfH
Obq/V7FBxjvBTfsJhwECRI6OfIM/50RSKATDTptA6KM2tZ253CwPzCPNmFqufSpv
27EFYIG+Fc4gtdjrzh3qVargWDcO/uKqhdjw2rVLBjhBas/krfGd20zvCUi7aQCq
dCEXsprolRgbk1nyL4+HUxefVGYn0Ts33HlN6IrJEcovfVQeVcqA2DJIxscoQwBD
AjU0JloS55Mhwr076iMfAyW8XKrAw6cBu9OzKLodnvuGHNG+3mcxIBLT8XvkUJfi
DGoibJQJ++5/SykdyOOCCv/5CLolac2qhGBQlUub72rmQVarjYP0M9qRCQ6aGYGl
9qECPR+4oeLrrRUNYLXZ3ueXCnesSi3DeeciQTP9j6w9QIpLIendar225HwZbJ6y
T36ZbRGxzMtmyDK38uL1IpBQVkTn/r58qcTfQAJ5gAw60TcmBsm0djdEy0NmqIax
xKWaNW3mUeRe5rvlJE1BFDduqrYK3JfWyaAMKE4jYrg=
`protect END_PROTECTED
