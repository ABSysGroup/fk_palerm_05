`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yntDnA/CIn4RjdDly8u2e87i0ge6MPfoBVORP4rhyn7d9W6rbI+e0h0X2YMKbcwY
3aik3+/sqMHYWtTOIcyEg/cPLAPxPM/fmBtB5WpBPn6MszXT52BkD0BddJPnVK16
ddNPMGFNftDl3HaAKAsLqDENBVwbdrJWeBqYkFWDTewxAARhx78Xn4Dp+jlmD4+w
4q4IRSmivprLKgVIQ7/a9QocmZz7mcAykb/sPyleWdhFuRrtMYVrXTIgl+GxWcHg
t2mXVI8R/NY12SixyPUW+yCi9vRj1+jjMPOcG1qBl9h9c+4OMWpVFMxaOfrBxani
OTz16QmAxTbNuiYo0nMHSDx+DtshdB6kLUwBR/uKoYCkeziviWQlO3iYP4LcnYI8
BBMKI8HIcNtq60MDMKVNVkjtTYZCMUctF3q7clBBbfSy2dODPCIVW76cOdjJRSnh
GmiMMBqNzcrJ08iJVvZO5xxVS79MMSVqwd2/I80oywJ2rMd4EnI18hwQatQZhpmN
XolzOLsICgsSW+Z4MdCD6IZ5xE3r9yJKxB3D7DFtMc/exHWBTta+F837GEiYBDDC
IufZtBshwaVAAW8P1uW+S6c3ZdV2h0aqaaydu8ZMNTvW8NBTxVkJBf0FU6+xDTne
MHO7NCOg2igS/LBjHvT0oPkn9fsrQRLhSk9hHYqLO2FCliVk7aKfa1O7lUfyUtIP
Rg++L7g4zyVJGvJcyodldIQAbJJhmW4qzL88py1MoL1S+jregBVZvFHD4gG0lOu4
DVgR/uLHGhUC7Qp+Nl99QFiKegXuRfalR/VSQ7uhKhh9maKVMWgyh4RKFnW0FFTm
Jw3Ehun1201qraCo2JMlexJLgrkg/wXy7i1iqBsTGWRD3aQZi0hft47csjmwsDiL
DSphMyJA3aQ18JLVp+eSXAP4tU1zzcRkLDzboQUaGFWXUxwsTltttmOze+r5q1Km
tKYGEIpTWtspFMVOU67bR7rcJw0OhavbGSdnZYZWrj0EpfBrk4D+f6yxes9xo1ep
i7LWKPicFErg62NHZuIFA+yLKWQCL6UrD+p9XsQCL91X3lrM0kRMy4MZUIDXJcoY
dRjI1uCAcqK+B6ZXOuTU+EGfdyomPan7KpljLO6Id5NnDJqZsLC6xTqQA5cnbeKa
8TmviPhnRtr3/vFEYU2BnAyuKCKQ2+CEX4BmGPgzDxrQBCt3yDYvAtwLuokFQbAj
jmbtRX5/AEAQs45r0M0DG7buRt5NRgHyYku/0bCX1oOgNp0v0BCot6bdPee7MQG+
aC3L2LZgGkzqNP2OMjC1nFwkHTK9yx6gXEOPLjNKyqtHV7SpJk8RBO41G9bzK7hv
p7+J6BdZR/VE449c53fPxNPSFL7CXSt13oGxcWgAqrV5zxDpLndpcE2ktkiObn28
HGYbhZv4dMVhJRys9ucnkIiklMeCnShWv5qzhO4krrKvwmpo38tRi6f8lFvl2kc0
lXHVyzvroQhmPfdRegEVU7h038wRoDouDfrCh39s68cw2NV/Fq3m6t14iqsEcud3
Z+iz9Jj+gvFZ73Lz985Xs8NetmbzW71Mm0JsKZ5s129nuOrR1l1ezBFW7Uk7KmNE
EbZku/nAiDNE6n9xQ/qvc/AL7acBAsjAZvRJgqKWHEqr2H5F9aOyUT0iD7CayyYD
S1/hSwYpy/Ux7NZTphxBwtt3i7/fnZDFOZ5+w1gMH4tXy4fAoSgMYsTce3F8H8Z4
tTjDSIJNL7PiyoDFBAjWxQzwF8A0dl1lkB16D3D0YRg/IEDQnFpzL8Zl/39/m0HS
Xt8PGBhqIE4vHLy8ufOgHbu8OtmBH/STJHvtTtPJTh+C8dhu8PnFj2UGyfsyIUn2
zFqtuXXt4nB2RRv2pfiBDfrQu5w5l8cy/YEP0vdVOZrWLIrHwSl6aHZkmw42g2b+
miUJLxFyGVMWZTbuTrW1RW+JkA1ATNfO4xaQ0kYHtu68rg5zqnhgKonMe+Y2N5+A
8kClcLK+qcfqtBFGQ2rgIYxV6iXYJJq1MJiEbzoOwXTUehJMQLlLdU3ml4rboohh
DhS9ewmJ8b9nusAMJ7+OtJ6xnYHwPc+NxV+kkG+UHyYVE6xmra+4bi5KYmFsj20d
WOAPOhTQUjov7OBglEBS8SoYeAGiGITkL0DnNIfkn8EYkDvKeRrCYByl8f3/2x5k
F8gUsM9/XkDh/tov3doXCnU+2rY3uJIfeHCtA6t1lLKu09u7+aCs1Skd5maqIRWQ
58+5NjYERB91qjOd503ZBfY4LnySg4VfNefOPNZvNVd0noADmSU4XhL51G8m62zG
05hNH5UOp5MOHcVWVIjnH9Pz19dWwPgPT3SnFYwMQQervGCA5AdcZ6s6ayiQPqcd
Js7Tl2Zs5Pnq9FQSXhUavzCqJPGPspzzqVpzOluKVoWOopJUan2v0nHX8A0lhu4f
uH/99ZgxfDTH/3ghL2W4+/BdWlmoip12uK4GCbo6NjA/vG9W25wdJF1OYi/1aAaS
13c40b1g9iuTP1dbrSq2BBVr22hiQ+xyKWLXwXXrrbiOnELroHeva8ukhWJQ9wBa
qjJJ0hm7TgdixSKdea8ZSCetZU9TbSgtbJjRqrhr9bwItIuOD0H+3LtNAC1y0er6
nmV1K7i7KIevlUYe2in0QIzoN39H/W+iuguXDkDVJFKGrmzNsZCe49y3i2Aiy162
cyPsRTF0qFou3b4DjgoIxTa+OgGyDkWYt0NFNaOW+jAMM5iCCX6gFh0wKnGbkCmN
hPEVvWk79p5sjkZZ8DkgJREnldpoXj7V9GbMjVf106PBmSx+5jgLfviHEmv6TA7c
mbCBs+R98MmCxtVt9UUrmg6kuMdaVkDb77d8+gNKI4rvUrbFn5sYM9l8DMbniuNL
1FbXtl4ZbddF6n7fovecE+y9LEW37yjqN8l93NKC31LZFrsWIkL8hHoJReFWfIVq
I9zerDWkPUbQ8pSTDe44rdYwofCXyUjVq225o6+4H1ORBSOPQe3OWxHC945rsbWY
nGHxAEOkAE69bnZ2TwM88IRPI0FxdboE1naB1FaGflZaIyz66NE0Th72j0kt467P
RW5H2THlyvxMkwkv+sg77GOkR45Mqb120AetGFfrHHjzhbPPWlVMSxROIneGBzyb
Z+iGHsQjiaZzkcjOrWEebL8l8ShUloSyXYItuHpKZlFJ+535FFRLfVOCbTJeGV+F
rx2o371D/0/+4/QmSYJpd+8dVGkLmNpEeImG09pFtLfgPxdHf2AB4/MQL5rWIUed
2GCFL7ra0juHeo8f3XLdHryZeErv0oNWJHa6ZS1k4/5RB/jdCRB3Nx4rUsKlf1XK
HzRtW7JLkZSdUNC0+W06yYL22PMJulpxXPfyU2RAn0372bCCpC+jfw6vtqYdmDE0
dol8INGR9KXZO+c2zbQuL6lkP5xGF0SgT2jcOQ43Kz+vVFPvbF1l9Ha3/BxA//I8
CEWRRjQKN+yZRVvbC3u3PY1QGOQYRLvjLPde7CtdWtOKAMdbb/lLsk4RGZVscAJF
B7EpxNuYio08bAnUN5anIjtoNvBBLK0CgeB8mQw1Hi2rmGD+i8CcsJSBeJUr131n
ixPd+UFRSqMXazcEmkaXA3ipGXW0OakKO8WWX8MiOAdgH2fY4nu98hAaIvvxSNQT
GGz7WQHdVth3Wa0bn8223RNJB/CVEoXpvTTE7NbdC8qYVz9eRpz2EGfSdHWivNLb
Kw36r6KjKROewOoZwSRTQHDErMa7ir/ZWAfTkcAEEeNpJYGKRIANechGJNn5fUml
OMBPN+ZmVhawzh6ztsvYz6uO1BO3KW09hYUK6BEQbfeL+Ci4gMHUVuWvF0nf8++m
rViWmYpzrb4EZJWhNMRAETak30MNMuNIct6kqaY/r+kqh1jpNzWzC/O5VnPqKyNI
F/3gb+pDUY/+mWrqwJ/QR5BS4/fkjaxk3mY8au9GqoED8ywssFzksZJ95sjQKT9m
MQ08ozMiZB42uf3C/n49oyRqq9mIc0KKHaF5w1PZYTRoDqjoDD14tHqA2K8ZCwJF
kXHojWeFrHEge1xAWQwXMhzj07dC+N8eVsPMHC6LEtd2WVCo/MUaGiW0yqX08RoU
cltvcZalp3HRpejsdbE5/LEZE5ldCpY0BqFE/pfBIn3WI4GGs4G3B+36287BysCC
jpIksW2QV1e0iS2BeNJyAu2hMhu3rtG7ZJ3uroKhNOOlgc/JpPdMu7lhq5miSWpU
nAxdTqxLWJjzMFBYXI7WJ6/PYeCkV85dEXbz+rdtB08ztbJoNWiKXjk5SXshlFjc
DyW+zMZLm/SjoAimb0R1nQeVUt5L2Itf717gVtZh06Qu5cdPxhJIZgu3/k9FLHtg
EC+8pkS2TOWAQIEadP2xhPuxrAYc/dBPYDI+OrBf6TrG5FqJpJfaCF1JcOX/ihjV
EPUOSTWP6p0hCa071r1VyhECrxMVQ2IO057w7cOH7YXv10l32IZMJdTBzBNsg2OM
8i8kWkMnGHnHVE7dF1D9czqp4p/IyjD04q7XFCdd1CVpIIGIKEmuOt/lRlbOXQAq
WfahnWZHh4vmbPZOz0DTk+SbzZfE7ZSCNFTdVxGWYM9BasMYwf8WJ5bSOiAM1bOI
ARUwmSWd9WBeHE4xU8AkchfATdq013fzC9z6W4/vIAN6HDnt50NOaoYBiTVKkK73
zSgOsTk6C9D+9DZnqANmFLZ2e9SPdNkxMob6G4GIQ0HMvRlyoiRFFwwja1dEEWkU
MW3nWZ447bjJFVnCNGUVgA6ociGDTMTIwHIWADkvY6/8pLt2sJz7Si3sTQSKD+5G
naCRFJ/LiKE2O/Rf1wOdGRqodcmHgL1a15hnl+pY/v1aSqvUoOP8QnfeqrPg3gku
+ie5vyljEeFuM/WNxjRB3zHKMZSNgGdGaZpPVP9GNlCsolyHvBwCsns7cXSO/aMQ
35TMB3f4OuGY/T8LDnnlG+3L7us88bWT8g5LfIJXuCJvc4qsZYZ4ISC2AknCCbhy
01HM7hANzPLd0ytZgLAa+pP4o2RCtl2ZCS80lCsabX5gSB/BdrDsx4xn6Pc+/Hck
obuWMOO0TiEN/ht7FTU6sSQBJmGM4ZgwxF8I/5AOSD6McQ494755JwBjFaRN/KrS
GxB+tswJjLP+1IzDtXQa0E7zYR7NdsRxxi/fTLoVhLoklpQuWesefSWWFpk6AAZU
S2fcVpg8/+oD2KCdDxWeH8SMEQYAuQLMvRNOeNgeg0mO6LEoLo4QTXmIJcJVjeSZ
+PRyu51/mNx/sB5hAhyEHQWHvYcJl+LVdJTZpLgv5EOUQ/IzHUQZLoLix/Y7vqIo
WMMdQds3an4Cpl3A58EOq5dlYp490TOHRMwevq62CCz+gdl1KZ/2csKMYrWucLKj
uRBXuyhSZJssG3JVdeT1fYlXUh3AoeG8XqMKN5Kt+yW6Xm+P2OrJjqc0UE77QUBd
yGfyOFeDhwgHHNHlQmhM4IyuVdy/JnvbBdtMu7CYY4PvVNKuhqz4l+Mz2/gMxOMW
hoVb2V8/L9FAbw+PcD1duJgqQ9Kl3iNe8tfdcDsdnzf6XRTw5qO/E43NYPyJbyxC
vUB8sqaXv2JDaj7sWisq1vh/wf4SJ5EUztQDoIK8Dfi+stQTtHOhA8T1INS0NL7k
62EyyKvn5DLWNh7scz+K31Ja1REf7FM62qeaiRwI26/Id9IxFZ5UtNGV+7mJGP9I
Bj3V9Dn2I5kcLDT5OswkkouIoWmktz0dumjuaAOAzcL1s8p99MgbDfdNyrfMfdrn
M5TxOOTSyhjMZgYgds9iF1mX09pObyjk0ONaxj756i/w3VHF0zI4CqFfgyOjKfKi
4qdl30NpJNgY1HwY7veREVo5G2XwGH/6PxS/bcuO3ZKJC4ZFVEnOp39OexX+vQ6g
hmAcSRZh86Z0mX0VE2upl2t9fzSi9aBImo47keLyuAEFTCei1jHNGO3OITyk3RNT
AvaYI9xg38jOOE7qcAYeirWGpYdXB1EDCGrLeGh4CSPAdrMzEnqLYj66Liq0N4ds
bFOjBrrOAHq0zA0NGZ4XhFzZdJM1RSbezFtmrRnR+Hivc05AX2UjB0CeaRgWBuvE
7F6fua7qeg/dmzlTZJ54EekJR/bG4X1d23rv+vXivuOrD67hJOXiIUz8ODLLQ9gA
labLHVW6TEB0tqSuaAfkeLAH9fXoF1thLjnrmy5UDNil9EnUp2TuvLkp8q4uwk0R
RiRJQIkXi0oxEiMLgz2KP3pkD5UiyZ2+4FCBI6ybm3flyiHr8biB3LyXkbaHYZEo
fKQMwzv/97qA9ASnvpwMMhJm3ZS+cZzkBnqIFwhNrq+mEtGoRYcLzI7c0t/BeNeE
9VQ9xMmWD3mEXrdF1LAtC0U1joK0xm0kYzI8QhPj3R7PCr3MclYxFXZ0/DYEVC5v
zKHdoykFuc7D7bHut9U+l98vEsGDKgJfo+vuQF7+0fW64wjAQq3Ds5H3JB5Nn+KU
vFRSTZunJhfAbWnnF4xLkescYzXO3/n6GWpV0am+5euw3WzDB5m+4OPDwR9CfoeI
5VdCvZdW3SV2di8+5N3G+usH1qcYi8N4B+e67JhOwBN5s/iD6nFCoyTzOkUqVvxp
3buWb5SpPW+/xDhN/VlpHrwbj+JJ5vGxna2ETSMRNBzRuvGOjhqmMiHLe3aQANpv
SOCFEhnEyOqD9R+s82L1PYs+BpW+ZfOrNYuD0DvsqsWQ4P9aGPmqBek3nQYlxp+R
nu5zoDeg9vuA4MPaNLPsiANoEytEdVA5GnSmOaHLyjezkBqoOA3buJWL+rKl1cac
ZPMHWGTiHfzr/RpoeUV0Nflc8yhOHrq+d8t3v2adKzcbjMHcp57pTvt9lDuNtaA1
5i1qCGJUpLz+mdujG+gQKxKKBGKYxQgVx4Ypv5Fcxgbdnca08WmDjyHGVoz9xD3T
V73yJKaDG28euXjrywPJQdzN5DhtrxQi6DRgHID2w6WVutTv+miJBuxwVWvGk9XA
lFzEeX0It6s2TDWMSnIwe3q8vbYvNYTeqP8hMTBz2Hjs4TJnLj0a3Zd9BxgeC9Pj
B7XKl3JDOab3JyinMv07DjEsJprNNF9rZGbBAe18jQFhQV6jP7X059zAV4jGjEpL
xDuZ9BMMQKeGiMIG3kUPB/nRVmMXWTHRpvmmNTSYpNI7Fdo3UfM3LCAPnwBwmohm
AjlaIW72MW4RI9WfBfav2shOXpUFmBQep1K3E2Zmp+Zwhmd8uWceGYKTzcYYG11q
ePy+BwGJxee3glIclIX/ry+8T3xHNh/a6WW9U9x5a54dXF6eRALLK1Gc1fLUmWul
Bqts7k5BR+1yu2uqwmXu9u+Dc9T+g8zAc0fpXVdym57pzMkxjqcjaJVN92rO75Ep
2x1jyf2gJCLqr0xOhyQonhAUTD3dLxWs0FzTarOKns/SbW0EliS04izK3iKZhKd/
E2PV3qnMIWlrB8r734nMSnhSAyILkTdzG50rxQw1R8LHgq3hF4AmSk8tH+30m02e
lAT0UU49dBNQZjEYFWdMo6RyBmZDoeAj1wv2g2jlQICQjpZ9jfYa8ylJ9rvI48fT
K85+Guq2/8ippZOzNQS6BsWGoH/fpnEtlFLUvwr+/XUGGGXB94rT+o2warER8H/t
61GHIFLejT4EvP1YTMtHNKKkpwh4GlChdyXLTXNztZHPBMtFSi9FBlT3UdtBAS9/
br7OP2/uFpwu/Glud75rqlqSYJa72BZSK1KxUbk153pEn3qZR9GF4hRBKaGz+AMK
vomKGFMD3puAw6z+PyjRLrsTH0cG3jPc2JEMgFfn4GCvyLWGIxHGNQNtmMO4Bpmz
E/1nSmlK9Rkmze85r64q5hS4dOSH9n/l9MbEKdOTz53b4e3EgiyJL5jOWyJcViEw
/urcx9EFqoICCU58UNQFl6y9sdLajvwKbYSxK8CUzNEldqx7RlrAsaKAT1TLVGjl
eVG9O7XyLoBdywsZ3rWASvhnpKdZFmvDHNS5q/XgOG41ADYRH3QVwrzz6cDB+xDC
ne1a2l2mlxzm6+YN+DuzFvVEOtThLguOwWlvF5oXmtRA+1rb0ZBieFWM1rjvnrlV
8aNsqPna62l0zk8utrr4BusblEHHLIpDQnfoV/MAx5r2DitzKhEOnuet8SooBnLz
LwqcRPfjUtWwpkfC6cW97UEDSGYX1JY/i8hHzHbTlj0pQpr8ShHmqcrshH3sMJle
oyypB8DRTQhqwx3fYQHTK+o7gtqWGtVMw3ot/TD/7xm/BkfVvVr1qkowkKvd3QTH
cKkQjeYMURXtb2mgA05Qmx0auMUEF9OrCtVBGPHRiasfyhDHuVpi8znE09z31/Of
+WDg17NYTYOyNvZnE16wWBBtf0HnE+Tm2hvkZiUvl2I540ea8/1vzLWfL/+P292j
K27via/Bnu5B50GSl5b6x00OgzsHmGLtRL6Qh91Ygh1Uua/j7s88/SiL0stfONIL
xCdlYudiIu+IKZQvsuxIslhGRiASuUyS7EhRxsTCWllV4Rxu2T+piMInqP1A4afD
btoLUODZ1SO8PekusSFznJy/mng8ys8/Z7/CyuK+ZT8aI3pLf4dR0WKx4cchmkrc
HAJB5C9Kzi2Bn5wKMvhejJcrosE3vLkzFc4JzYxziilVR48KeDPZJ40toHYfgT+f
D92M4EbpgCgyBaezlqs2PvC2M5GBdxwiTpbbZbW/pDg202O4pTT0/2ilaE3FLeTY
nSlKIvaePM9xwFouwTn8LD0pYIw9E6Kz9miMuPazijXOg5vnM3bw5DrzzMN0ocio
k9BEV9hG0iIs0wN3DNHZVppjn8o8kH/A/PuohBVAB2tzqeY6bZU/dMa9j7Cwm82j
hnfbcMwEavASTqhJ2EazzTwuMev+bdUWVh/8M2QwADHB8Bn1UckgDc7Fh2++IwSO
442cCjRNYf7FBovPsb2h+tG/efzIXms/nZ0pisgQ0KlmOR5LJzT5Il8JteLUZVEz
6a9Fnb1WyjHXyRHbMMbXSlh1o5/Eivs5gER+MhrKDDLuJ/OodS3J0MOjGfl7A3Ad
oUwSXvmWpVRxGDhkHDt5UhvQiItxHxC/Z/Qqc4j07uv2qvnq1u8S40wgqapILeCQ
d76eQdg3j4qZMza9NkNHqw6574boO8qLfmO7E9+HTab3ELLsOSStSbUBKSiLwNdO
5ZLo7DN+aU2DfQIM4mkYhKHU5fi47J7qS4/pIKfZBPIlL3UyxSZXCE9We53gxj6y
5yt6uCCwV/6STdK9DBr713oZqeiNDBbBfoMQugapLqJ+mrYUCt0J4scnMgOA0V9X
p0lz6PbwcYfem4XQ+tdrPUaMAnA3KCTnOkAXGaU4MrEouGb3eIkcp9kDe9A7wABF
TsDM6Nd+t2LuuWSdiEbL8qEXJvUt+rSCR6E8W23S4406mLKDurtYxckcX8AnUV6v
92JKrtNQX/dBWgLKeDppcaI3fOefHTfxcQ2QJeLnuJgQdsKxLkJT64Zrqpe465Cn
X6d4oe5Iyla5nkY+OYnLi8Siyv3k6VINME9C+4ZW0VqpR8LkkmOw4zo7Lc7UKhfx
st9jMIWPDDl2iktZRAZV29vmqAG0ODzeGD3G5M6h0k1PWwwAhz+Z9sFdIudydWng
rkLhKame2/Bq1vbzitvPVHEEwGVoG6stYUmoTOTJEetmMtR0Vu+DPeLMeXrL+1dB
tQ/ytQlGHZvWb1f7A+0xZCi09V8P982NYhUmOFF6t30zMyO4cTaH5jqPI/FLcU7E
5ddLzKrU4GQvovls8c7KrfhMVR4tGts/OwCDvCKoolS9jNzJDRwZklOHugqGx3hm
cpd3MaUfO13W80wqhk0psbA457k+oMLPVNw5BhDOAtHK7SG61to3VA8pnkW9ZrmH
y1+vIbRnL69TopUj5do9arZBe6h2ghpFgUxBU3A7NyMmoykn2brmAJvE3kZu94fo
grX89bp5GssJwJx4yCaq6QzfyVeTCnmv9346r+czLMdAghnjTulgk43T2i0ecop3
jfvd+jOwAX1wpULVTVO5Z7HT3xnxTkRyMCqjLMLW/qk+t3AZT0rqo7NrrzWAeaJR
gUQyWNEivNoK/lDP6ZCXWu62mQFRNJzzq0WJnN0jhy7OpxrBbyTn5ETMUeknbV7r
r2GXn6Bd7ft/eXKr1zFzUcY1y/yteObRP7RdbiYyHxDqSN9maA/Dq4DL/b/lTZ8s
6xCg+DrBkJd4bLuZvNEJ0F1U1ascgB7wjPdMbx+V/pCjQVFJfmXmCGPJ1jMs1WoX
N+Ar+l443GG20/8KlDSXVVhZg2nYSAuxh15M+WGE0td7IU+hsrxLaReZZXMpBaH3
hEKwxgthPuIMDJsc6b2IjUmcprJr24LzYpbHDtITs8Q08x5IHabD43OuHc+q6p1M
iBbnnGKvyAB12X5TAjPf2fG+IJU3Z7t01CG531jaAHrd40iUvQKteubkzblQYwnV
A1TaJnlT6pg8mY96V4Xwc2Z6In97cviprMRQPBPtgPtmHI3GyfkxIjpU0R6BFMgC
TmcrdHCfvVyoZhB7EeDx1+QXSt0mmA4t3+E8PvLcLyV7a22fLtdhcCZCUcTxpL9G
RzJm1CJLk+N7JEdtcG0tHij5QNjKSErDn7oalCCu0eGWCJIC88KjQ/LErTmHRnY/
6Boyt9aY9Jp8AWJxhVmwcXuO24YBXfANn7DpgsE8TU1XUlZ44trrgl0YNGFhnAV8
+pB2oEpHtyaV/k9Ucn2C6A+NsDdsYRlV6MTT6S4lBEQNRRj4ldgRWXAMtN7ONw00
fcdNgQrbcsIbKw9vgrrz24VAlVffeSLZqhOMRKuyj36KzDMX0j+S8hfuAZC4vyOf
nZizl1ofuGxWOwE7XMCthKUAyinY6K7v56Vw4/on8qYIPFWRpHF4jqYCI4YUDkyY
1VTWFZCPBSfJDvfKGGDuGQY8aSiljEyhitN7nMgi6iBD4b9JTe1ghVPsVQ7OTJDn
V3kD0oso9teM4ZlLm71xEzaoyFTTaZFFpBCDJ58CYPd9gmqwzuuGr5re6kReTK7u
bef/503hgICMI4o4i1mAW8qF9fZfphCm4qgE6SAc7n5vEhW1ZVgTCnR6SI21F7s1
IZ5QIhfhCmRRd3UbDg4WLwBmIYyNTQkUFwSAhDaHupQSMZINaKzyw/r4Ub3grMQ4
QtOMJHt+IEUi2WMh/HBkqO5jkQg/zis7aPka6q+W9td9ysXQT0FgB4BpwECaUcUj
0ZEuRrdPb315ciZVPv06OvmH1FpHWc25hor88XFv3LjxYWwTGyHRFLIqe5NAO2TV
FLZMoMwejxM2clFmXyzuVr7kJV9aG21EgFcseOK8+LOuMn6nh6S3BdaemnANjYbA
osu8+NKuivbZO0lZZreosiecqQCBEIzW72Qr7tiTBz+AcDAYSW+sWm1yH2WKUTP9
79YBg65uMN3gMvrP+C7WjKV0TXiSHrTzuhMQcRrjGjUitKmNUSdP39FFvUejipKB
3cff24kH/DlZlPTK4HHIzv0tQooSBywXGtgpbfSzEsHzdnblCxJVMpwZvGvRlH4J
OAFTgUIvxlUTHffgDNHGQjz70PtE3ityVWLbpHuaN3YQex5sRZ13ON4M4Rn0LnZA
dq0SVxC9QldTZqKK3SvBaLmV88BOfF/6UBGRa//HwJ2j1XXz9khDCYZBYTxIXWax
rBJBOQFU+yq3dEj+Ot7SzGUBqVP9qbCC8l+0eVSIzue6YPr3ZTgGCNMYw+J7aN7t
KHPfE1mj+Xv5r4AAR6NBwBOn7OT6jqJ2V8nMJv2RlMaMlkxD18g1CKU+1WasoRP3
YFGusj4rtXbNqhQYM8IQh3XedqDUlSeiUY4wwjQZn2P4wmPFOvdGxSmyCIG62sJZ
rVjjpEirENeO7GZDL3ytfEFDSLc5fmFLk/WSLZbAnOVfuX9fEFQKMtICG0yqg4md
hED2mez8sxTb4zhMx/wsPSXAbppLZLeGAz4WT16mUyq2c6ok3V1vFAL+GxJuCUe3
dzZJCerf5az4Ai248tbIx3PL9YfS3XyagTF3DedcraXTpIctysOSLX4Alnfyjf8/
mvcUaxWwQo77ZWDnfSRVWwdaOnNu5DBVx7U4MINHHlI5LT6fjcAJ0zdOalrnJinJ
OWX3uijbzezRSvMIrI64UUhDDUYWjd8VUkJFpNGEsQrJd7Q6UwEfJnaXiJvw30a3
sqsezyDTh1/q5whIqRGxMEbnEXp1E5/g6Z6hyaqVSq2rES5IdV7Zr+1PH0hlqXAP
UK92qHUmzAvseBuIcbbhLvlJEGEvK992YqpdN9EMX5dll0QrSvI+2R2v6Qg2bwns
HfQ9A7Xt62dIOBkkcy3fTfSNRrfjya5Gy7O4qA8dAyRWRBTAgS3GHGn6fw04Ily3
Cq6RMYf3GAwbH1mYmhMAWzlI1qnuCCcJLqCoD6xmgtpHyMEUccqtWcxmk3cAtHsm
Eu4JiRWwDJ4SrLXq9QMfjolBK38lfruHN5ozrEy61/WM1WHdAJ10mDUz/4N0DB1d
z6QHeSY6X4nl+B7y5IaZy2QANsQnn9SdzVKVfammwKR7l3rE2Eexq7TyAYzbJKTr
bHE/JzF1EQFB+1LG+N0n+LgJXBetFsXpGwuRlpZOgzinUR9fds0bY2IEw85P6xEv
e1FMoS8D4J4V/dgKnz3C+CJvbk4wBfbnUiMAyB6pDqOdF124+gPJUMar2KvfjsZd
qYrAHE4/14xZ3nMW+8DhlyyY6wdfC1egdCZDeapvmD455C1BP1I5Vyxav9b6zbDf
OGmasCgzvJbIXhZwJ546r33g/cpiMclHcf/+T2ajA+sJxoaXpgxbLQnDtoLKuwIR
HK+yOI3Jn2GM5UDQmxVM9rHkCpcPDZZ0CirO3Ah7fxlbjqojvx1qE0j1BMnoq9vw
GWxolf8kgGNMv/37MRNjfsgAP4ikL4Tw8hIMmPt9ZLg2ibPXqZxUm5eQR4Bt8uAa
dpZCMgrC6Y7NCH572DZ7S2XnmhJWqCCLcfhjc+zRMS4ySWNYge3vwhaOXKtMAmol
Qh7jtzPhygO2xCBVzUFJHxxbmcAdTzrKLLeCHbuct14IaCaaO7WWh8EcFXKyAPJ9
gLljqMlAuaiOxTqdFvk+Ol1QktkyiEEo81s/jNWoykp7rT3L334Rs0IzJgPOOv+W
Bhpz0xulRKJmRcJ0iVbQzwYMm/qOEMpOi3OVD/mMu7WTV1J5xbXPOfM7kyYDoE4g
jOYRvCXhhWf1lLikW/0oyDpCScuHI0EKeI4P1Eco/A5Sg6MHhGU2v8/q6GOdJMOe
eqmR3Rx33NkM/fTUGXSfUdRg4emnUrqV7KFr5VC2zKrpFLS3ZU1sUQo6aMZaH7yT
ZlQyAC+y254pL76KLAhYbcYKDdTN6JKp0fiZyEySg+B0xWNJNI7TL+hCBXuOB4lR
tNK+SiTQOWpxKCLXg0uI0tMmWF0B5QafjZEwR0ILgiwM6k9WpfZwX4IJuLsFprIu
mOWCzS8I/5YeWu+cKb4HbUMYGdfTg5q6ePMtiI1T+sGfAcEcTO3LM/ERr64U0B/i
QMfVtrLeBXKD5+TloGdixSQuBl0zJMq+rsnSuRNUWoplLMzD2JDq6n2XRJWyuzCK
keEmKp8LBJE3Ts8AXJhjergSV++1wXXiSgj15rUKTaSoUWZ9BuNmdoi6hPQkZw5+
zKRceNSCDqLIOXRjgnp66/U0LJ6PcWlLKwt7+b5OgoOx3yumeAKBhwavaSk9ocfS
9Bs6Jcfdje5dF7/XOhgEiz11cGGecmB99JbbwE2LQKWr9ALgfUKFplrqWOFvkBk9
YnXdwlVwnTmp6HRklA4KpCWEcwXsbqmwBQSKNJpZyG7Xqx6o/LhNSl+CRFo7dU2k
D9+FFc7o/qwRvtnuI6LCKMn+UuijdRSGG3Q/3MlTSdZsc+WHQpxAjbglM4J6Qg7J
NXfOSkzOBcceoj0cVf4DgC6KgLY5JfPPBpg+9A18nDbfqZCOsHWGiDS+mHkrGggT
EKWWyn8vSP9JHBYIi44HYTBy4LUd9MVr/L8jRJFgulHHqjA8+6WKQZxbfrQvveEI
llMYVY64V/mtfKNSqvRcHtvDUywfRRYqbY7ADbUqtyCheddkakxUgXHQN2yqFf8q
Uw+Suzs7eDUrDvCBJpKU3436IKr1XjyNTqSl9ImgnfcZ4RikSRtAa6dRq1iQJkrp
CZbJEFo63okck78wqPBsBFXCTE7QCOoOs1X0i1JVzKo=
`protect END_PROTECTED
