`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u+iIcLgDLbPglc/PjD4bpdeUtZC6ffvMMalFpGbkZhUha4WKQ2qjEp5rZFDGDP1r
ad5ml3nfmRFd9XB2ceAgigCXDk3YgmBAAxOnFoZ6k6mU4e5h1Bn/8gFoNGEzHnvT
lemvSCUfLt7/0RQU3AYuuzwtFbmo7ucGoNw0N9mgO9wATle0Nfv189WamVJMrgZp
x6H30tpwHhpLoI4lStsK5rucZiW8cs80TZdv9dZZCP+z+2XstFpMg7RW0hiBLcZA
zgtQRnOyQeNkZpJRLjYvTKNMETm9rMWoBHTucRpUeT2sZ1BD2Ma2jZATJKpXn6AF
gTaQLPsISfimHsdy0VC1QAk42sfDy4V8H2Nt/81dLCsblKuNNKDO+2SfBRMhoDaV
cg6mCtpx55RQk/CIEzanuBtEQDURLtRRYXcFUoXc/So1eDTdJnqKliBkxxVfKMwY
6XawDMVf6HI6mie8LqGw+aRN6Z8fzVsBR+RId270aevVkQ/+fT91Bq/JWdJy54Vh
Fk0QIzb5ExXT1WPkIcGbXjFP0VVOICnkgt5MbkguxzC3ewTJiwX3EuYJ0lwieiQ7
B1G1+BcOjE/qqhPuQCd0rooVcGWJASZ5RUp6k24aoqMcUlnflvjpyuNqHECfbM2M
xSSUbNN6iFj4TeOFerdmwBQzeidFqYflLAX2r0AniO2gx+cGkU26e1o+vCTgXC5L
vxHIWvQQ1l2YuGbEdURQsJ4RX0vFkW8WR4rOXteC5vvuZAWMWDtoguzn5GYA66aj
tPN/gln5aOMvrWqbWZqko+2j3mnpER/pELJqEYxrbCqUcYMju7arMC8E0x3PaHyv
0mh1b9ZRlIKaE1P+JMQ4SakWt2uM4/nQ92/n0PwTK8t+eP74cjjnvRMD+kke7HuR
ZRQneApN/n9/2Fgx2COJshk+WDC6EuhNWdWOsm+wlvKV+T3762vfy6xtB6hiITk8
CLfo9Hn9e7a0NYxaSajuExZY3PSDLCqMFfHYxHTTniXC50jqVPwW1Ombi6qQM4re
VWrR6CeIoufKeXl8jq4V6v2lmh1cNaCrrSQpBYwHQyOD1M3HAxVRf+mjDg840W1R
GS57yS17QnjZPRolhZREgJVmU4xKhCjbCtgyYHiyNftqpfhQcYYq4C8i9+j6BNPS
JmmAqqVFuIXa2mrg/E/ugJAqulQuUKaZCvf+cqfjdc5SZr+VJtWypg7CYD10Uf+h
V3ODMh5hrWYl8pgz954Y5TJCP5ASV5B+YnQiZJ4bLlBqx7oybZ+3KU1kw4281f1S
u9agZsKmC5GoHoX216susRsxeA46LFXHoTkZw9Q4ZoZP88XSSKfR6BGcySrGVhVY
RgdYr0XjUFkHIz8qfVhJyYXp+KWJhNrDwPHNSPaUsjkMkJa0NdgXccY9rJp9yHgF
yqgO84f5loMnZOoLRfs9rA==
`protect END_PROTECTED
