`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uod3oldGDwwYjOqKCb4MphCBeLOGKTGmsECGhAlgjpXeBPxUzOs24DG7KE4cVZJu
XWVqF10BXBoSI2kz+3pDOEgVd32WEQRmF1k3EVYncmGIhh8l6tkikxOsehZ5b3fU
CF+vsJCM832kjA80JgzD7psxsVGVQ/ufPrxXtI6FPMc7sQm0j8EiKu5uAjvMN2O9
8vA+8P2b8IYIhd0FMAy54leNLVo1GTZrPypvyAMJRkgfPi7TB+oKL9EBWDTkJupp
X9SK4bIiUOun3NTID3cI8vX5uP5WieJCVKz3fUx28fp1QvKNCGfodNOpC4fqazF8
zVKhCIC+jVZtWy5/PpBEN3GmBGMRQ0UDKaHXLNX+T5MtVNtLCJykcawLUnXvhmZU
LMbbxe5IxKojEE5jddfUqXKomH4F03n73TUtnNElzgZqaIoYWohv9fDInCCVhWKE
oP6WUls/aLmql2mSxhbDz4EaUPobjjSIRjgA8nzgxABX0aGyw13re2Ned8A9ojO5
rBKZVQ4atv5Rk/J+BmADy+9cKj1Qivfz6zH7QEWf2NIx/H1XjiH5sCmj4MGMkURd
XEFwBqT8pBEDea4514I2cwXvydxK7NNaW/OFsF4gH0nyspwpmDUeVqZgadhBXO9r
EaW3lJo8CmQzJN86GC50g7FyeE/eCND3zl83Uf76uMI=
`protect END_PROTECTED
