`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tZAVMl2mxp0xBXsYYHE1d23cyM016JNF0r61YxwSaLqjHZ9XHnYQjCoOtUlpYlJ4
Ies/C3BtbPEDXBaZTaJCD0Ah1lYWkpK7GIaPFgzTLiI6eayyRB2Z3O/wQiXhtitl
T8Yf+q1SKySBWtE5cUsqjqp1+tumSyp+QsBwZaz3xw44vDGAbshSN9WHUOvAQLE8
ZMGQSAaF1BDuyniZzB5PwFWJQ3de2CWiE2gR5vScaVONJSjRVbZOd3Wo/zK1ljAX
DW0gFn7tfv5CcwvBeNylwiCBMocwaDMUrEzmQPAKg6G11hWHu5wqbvbwPiU0cSId
kutChLZ1+w5NGCqu1iRW/wNxSCuzSn8FYE508uNbwbjUxW1I9eW1Qu8Oq0fTSENl
6t1ZzsA6zkvp19UFSQBXUEGIorW/662X1UcM62CVSaPiZaJnkpbSWE3mEiO6zKRf
`protect END_PROTECTED
