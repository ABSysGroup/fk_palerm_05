`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ub5YBs15c/tb4W34BvBxVo6ynF5We9cCLlVbZBJJP80vjKPuqb04iQl9aajTwd2X
5bWF8BsCNx46dmMid9ye/t5L2yLVLs8pyQL324fu0iC7poZakSYIG8ApzrRuLqtG
9A9Sh38V5qjC9wi7VDabNyA0IV2OzA+66iXyV61HcjGOciDBJiVrkzgfISCBfx1X
OyGysWLyUJKZgAXD+GWlq3NgzPFN95r8PE2OqiLXHePmQuXPONM5MdHD9NRoJZex
v3Ta3D97FsDtDZK4+EDDHXxuOfnCNM8VGqOec8/XNT80hwFS4Y9+XbPdcY1EBImJ
f/iPq03A3jeAGZZLhkVUC31AK6OnSmMEEAjmnCHLjwlZ6rS2wp/hC0WlowoblIYW
uuzhhJCe/CuzSHRxIozQeRNp3b3mtO/lpnIHuCwwJJNtP0FaJ7q3MjrIORg5Laj5
`protect END_PROTECTED
