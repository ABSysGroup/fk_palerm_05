`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zVb7r7e8IJEtOu+D7dKDqDqhNcUIvSWNPJWUTGq3WcBXFaNUdJHiiQ0D7y9hJzY/
Ud/L2+NS+ExCavU/b4TNSpy5SPPCXz2JLVieqvfN1dnI4BX8RAwq9ik6lzoRJdRX
PLqbdg/Xs7jSNVVA3LAvWyRE76xsCzxBeDMJfc79VM4fLUmIba/IWe3DA+Q+x1XG
gYFPGDqXV+4JntAWSyrJvxkFOV9V88/OBKqqXl8amB53U5XJMu2DyV1neTtZksim
bYW0XpiMVev3rT52npDecckyzsaRFtXNUK+6h2/KpNYpYmr7U5/7cicflVg0dIr+
+IQ9rrYBNDuoTYx+SKqZhJ+nhEhzXCW3qag4GeUWb8kRlHfa4z67vqmDOgw7Mx3p
bKqdl7nIbXHJ4neRezXJNGCBF520EJ8rcL4G0yAgklCeKvNc8eAPbzejivJJAMXq
OiBvcFVtUXKF4omrfWBuubhoCc5CTb72FjgaPh4djlSmHErrndh+Y/3VN4v3t3A4
MW2oK2wYv6LLvA5hab8dNVVGMFlT5k2FGG0V3DVJZ/x3eycyS+et66LL8vOOypAh
teMA0srNCCYYkQI/+/BwHpX+HeVH0Lxgub75my6Y3bIABFOW20qvDn0Wk/VSo/F/
vJUo3pof2IZeeO+LtI6HYjs9H4xvpRLXdCLTb7ofuSPYg3PDWWyVA/iOTBsqzR6j
9GTkYVXerUDDZLblIxoSB3hZFD5Oy0OpGheyqhMNBYkbneInjSyRnOaoeoue7Avc
xsxER+E9ACSqRAj1AIaXSiaJDgvjkS5NiPve4yX+83/XT/MdRDEyvFNKxNbuZViO
tf7z1Sl6IGvmowxHbDp71qsm+GJ2ovSFFRMAY2ihZf4fsewUCqCjbXfQ2KhMxAnV
HuXrA+DPsLzIeQt6cuKZo4FNAoraXoUsZ8KSwyfk95WkmB+iAzTwJNSU5BqmERn2
EmcwWLCwtMeL0Aarq+OUexuZRkyNhoLWD8Iyhy1qmYVEIonf9CuYfObGHkicFto+
S+vYPcO4XnbyU37U43mCeGaGVIWMTdRTc9iHbdWqrCn2hIBjbzH/skczNV0OU/Fa
R4iMwne5MdpG7p8xtWetwc2sj4zyeOn+VdzhCyJX0LQJ+5PJn/RnJkZQ0whEXY8i
OdA/BV1xcTcidIAtM8RjC3F7XvXEIlIW8IUa2FMW9zF3Gabpd6xHbDViTtAHhwAN
+dcyH/w+BfgDpN3A1vOAihD6d3KQODnZhjhxz7OuwSZpXRJBzxRpZtrevLAwLBpe
/f+blU5Dtt3hZcJ5tMF5txJVbQAovN1fyihn5Kz6sJ8lXhbrnUzNEWQb8vBC77r/
pZyywga6C0k2JN0sgefGfyXn5nQNB6z3j6xZqvVIFcnQqoei7QmIIJD1D31bzmQg
+iRwQnIbZpOHIUwR+UjdsYuXWwu9I2Ow11tdG8y8c52Bw4+nxvSwDihApz8Z35K9
SE8r1rjX0RHzBOGa59nnvWqIn08lOaZMONgvWPntOPoRhVIn6xD/uhecMdrQNAVQ
YnEhAT0K6d/iRVwBF4QqE+6pXOwga3PD/WVvdq/83f+gNvlhH9v7pmoVlmcIvMfT
MLUqLkbGDhV3BXlphYWEqPxm8wBzkQeAS9Amxw/Of/xT7eqkGM6vobzjK6hrIc5Z
O4uPNanIRljQPtQMvPsCXrs+34gJPGnhhgWPoTh7RY8GnyhTSZOUKg4R1ZhvpMdu
aYWcSNMrBzJcCh0toZCibim+844lPjBSZf4qK49dYf13HmaRlATW7qtqmEDuDuVO
gm9EI9yKAUvDQsnCFrsWNOKR+9LaHO6lCYX6Sw/ZECBtnZ+eP2W6CbrXygNcVIlw
6X2d9VeqoJC+qWK+nHPlgMrD0uT6NHUlllDhPw422WbICLGh+ItarCP4WS6oEQqO
ciMT2tCgrWJzPHZMUcYM3lMuX2zrCQz6SfswbtN+NitEH/fr+ICzJZt8RP28VH7c
0lCKaG6pac5kJ+1MMLkzk2XSjN6x0ecp8GJvZVHkHFeERVZI7iEQmjnmg8px2AcK
GdCYuEVYeIz0rEDkusu20nsiTYItg0D5JRhc8GIsEVZlYAIpM8GhMCoz6qZ38BQ8
+CCISLpTrelXkQddndbFTXMyQi06Vv4uWZLNhCHZLoX9O5+PsLbp4OEDL2zYtsF8
pVo0EM5hi7779D2R86cMcGvgheGtqZvulRmuh46O44Bv5YnPMnRvKm6XBe4tLdiL
OkUNVUI/Rmi7jrcG3OIugqyide7pTnerXoSKPTvitu9hrsLI+gnVAYQ6Qv5xA7MF
wN65/jwjv/h9eilM3dKcVdcWD2FSWgFBVUVpfXrlkIRpYD1Cx8lbCOVMsnEYCLH9
dxXwIZEIsuHhE0gy0UneBpgFAteAnzdPMuao9KjIII/9We/c9PzutYwi0u+vRVov
c1m0YtuzU94ILtpNrz18W4dF2oz8xxerm8wRHxASMbJA+yUKw2SMJD/02d72gg/h
TZ1bafQbC7V+muBXnWQhchE4MbmpjRrvHEA62ZbKTDVc6p3BPkyNRLpTVW2aIO/G
S0lnjYZHP1bBwIYMYzUwTwO0Z6F9HnbYssDq3G709I9LLsZudvzAyVDvFpMwkB5/
IW4UTeiz674pfNjHtzvq+Km/BvKwN6oC2x+91+3wteMbAnCXHCXXpQbREUNSBlyw
u4w+hTTfsguiDJM3tW6hulQHWo4Mlz+8O40xg8XZe2h2g413xzzzLTzFuY03Z/r0
/xNh9uHRQQ6EREQj+w+6n233MiOX2RsKwe58OEWMHayL3WExPM+FupQnt6uNhu63
JYBZeUeEJrnS/MH3YIb4gB6cT0/k3aThBcbqePdhVyBVpw4e8gojE+ShZjSD4cDK
rBTExlOdFBLCsBCQo6ai2uJ3OZ/mq0pugYq2YRGVsNTZf+4esfA7zVBAFZF23wkT
UUptSEyIOp7KfyIvEbcu6/h+fNB8/SxnzEVYnKhMV7cF5wKE4X9Tl82o8nqBTNo5
aFWKgl2wpvO358EPEyOSk1LUbsN0LbkcXRvABaGQmwpH7s2GdvPOq9s8fsh2a7ie
FDQ2khkqFX1SkIFADG1oWcNUZs2PVQoO7nwhZ85JS2JA9OI2j2ivsFHPKzS+r8Pr
/KObtoPTgdz8hOyMvUV+SeK1mJdGF44yNytQoJRkrThD9D/YYH4EnI5m92yktn1t
GgLJAtAKuMrD+6IqWDAzGxP4bZL2Ivg/hmEEv5atI9LG1lgEWWHgwaBRr876Saad
fjcep7XrQ3q3HggF4XsxiB0/3rXl+4fqasRQFntea67HEVakp9MFgkMkqDcnz8lp
hfPXw2ABf3T6HxYQqRQTxRevBOsqdrljto9YnGuS2Ezgon1Al8Pf8eGN4uE6+Def
X8ZbdWyZPMZJ3x0ryk3nOadOBsLc9aiw0A14GeVjizATBTT1mcKB3qMnLut4fRbh
mfPPWmp1aNLbqzHeNgIE/HyopN0AN4T9HeonSCpSA5jt6QUN/ZrIp5s1YOKwyR2V
oojNZ7UDGHoYPY2bJeSdJ7fHiOISwk1oEjyBwB9a9c80yDFshVf7aQC+Rtanq9sS
FuWyQrhpj6bbFlMMckWTR4ZVL8JzbrmBSixfRHJU0yFZQCSmYI7q0gvqax6MstDG
BjqyoDdoUpXEtv3whrYLI7EF3gHMNV2Ry6nfeJKRhfKEI/KDaGekL9aKzurt1ke9
HgA6rZxLW7nBQlCBEIt16Nit0bwg54xZc6uHgVuln1UmoZsofzzrYyRw6YjMWJVj
muLXQomdghRqJoeaicgLih0cJG6M8gpUP86TlnAl6WhyCLzmXeb6Mq8hR6w5iw59
V3GCNH4FufEJlwZiT0gKtmR/dl7xt0hMAXl4IbbXx4LM4yjj8TKKgdgFvzOBFVlw
fDLoynLGrLAC6X5CI1ae6cRBlaNr5LJLTz46K+J6ng1pK5tnpVOnrwsgZWqAl9zj
+uqeRMyXBKaHiUS2yMCjaNlVs3g6ifE8vtEpXXgvOppHsiJ0OxThB2uYQObUCf7b
VgNA+DWFYX+wKXO9GVyn9mF0r2OIkJEDb2GZOWy8hRxqrexy0B2BcRXEGyAzWmk3
5+lfSAFYJrJ2Ya67ynNcuF2jWnMbRSKYbgiszGKdzTSYLf2fCpT2D5NXG/+pcZKj
W4KLdbigLNc/m11lug7mqMiqrhGZ9612SVeckyCfZxIKcN6ENoj814msRta0izcl
/T9kUMZl3uva/BzdP8UlbKLMcDnJrdlbUgd00RgBXMZOE+Jy0BE1tiTSCqxI1oQe
JLMqktCfH+D65D67ED2vXRi06q2PQtXY+E3phWBQAn80TFNYe4nx/ffck2MmLeot
8znmjIHoPXrm/2bZkESVpdQbUmTkmdKucJRCQZ6d3jR/LEtfatJI+D4yP2v4wTYc
IqPqEHJxPlRYZIhYqzKzBY264BgKrPN2QEEJXtHhY/ftbWQjmMALK/epiqineYjn
Apl3dCdh4RdhxH7UpFCQa7ljZFx2t4+wnvj67SJ4VrW/Uw/wpHbAJIOM/OXtpHds
NWOLww3Pzmy3Uk87RDNJ05zRGl0kVEBZoxg8AY5y8w3MvcQDj3+A39RBGQNzJlzo
UwoWBvWKcDW/NnyEkYt284pCacw6ELxnd7MZvbEx6D/MRccc83hR4tVWi/kKuhpY
XxvZBTIftpIn1PcMv69zXc40eml8GNPhpy2WDHRQN707oup7HMmUUtS4VD41jjE5
ChVb5Vrz7b42oj4OESz/agSrnAkhaQfHx6jZyefQkj2gX7YxRlZYx99ULPJJ6Spv
EqK+hyDMUEs59/58QACaW3xHdU7eEVIuxiOQe4kRrfvqRzCRXscVZJTdhsVZFW+9
N8cgLa/TbVSrZWgNKxiTqhbZxETBeU20OyqZbX4sVV0KhNM4ejnlJrMfg8IEdHxc
rZhzw8s9SAHduqFYhFAoGCa87rkaNES7Zjz4LkVISRFU1X6baNVoWtdFfkbGKpgZ
PQgBPsKNWw3/1YLFqNDrljsMXnR04m1bTRK6eEKjDBNOUW4jV6TCh7g/F9I1Z4CK
xU5HBmdE3kUD8M6566h/tbBYuyMBia5dMdbkE3Lzxp1s0uqmf0psQ3DwJKvPN8Wk
qQfAcGepfUITflmFhTMKxyaXMPvgTevwqVulixVSi2Z5obdu5hsBLINxYGuI8RN8
HYMut0m+qT9Spt1NL4n0khM+X0ZQyYzZ8maOy5RtQJgTPSdbSFQ7oG0TdI/cvbUS
sHgCeVBPjsp3z83mdBS/28FS/pNo7/lbIIaQjwzWOdlmlA9ItmB2qhpDPc1jP7MH
BULgDvGB4V/pi0Xc/Gj0IJkzBPkk8Gw3c0NKrB05FRi+TwH2l+KZtbrAkIwPIB3R
xDpj1/NM3psBUTqr4yfylekPuNnPJTKxyGqebLBZGzVLSE+DegZEeMlLBHMXML0c
/rx1wH1OCvqNYGZJy4j8NWLbNEAwmvjOkT5F+fkj8f8fXbiy9fUcqDUUorJG4/6Y
qPWFTAQZ+oA+1OaJAwPY/gKp17WoHUZKuSV6y6UyzpgH4hhAnYsgywpdsF3BFTqM
HDZ7bKt6qSaoCpGpX47HQKHBDaI4Gs5KHo2an/cGcezPZT2+DSj9oG9Uf8RT88li
TpX3W4hEL+3UsETU0Lu4hNNK9tn8KTXny+4ss428WFl/iN5g7IFpali4jFcP8Nbi
OTDu9in1gNkeqzKxKQnZ2ZkioiW0L4QzG9Dg3Z032PaeAq1PsX5qd2O6eP7fBufu
22yO5AkT4IT8DJ+RrosBMYBqJJm4UTzVHULDPR+N25c3cRYHqodTIv0XHtFRrrCq
u566kemtpq1vamKSipMzHXs59TC8NMhTzBckN5POdPJ/+TMKjA9dqyIQPhiJZeiz
a8qTVc1eCFufkqVmY/hlAFN1TCDZVCVDgpzB+A7GvJCeeNegfZ3PR/0N6SYI8/AM
iUVjlV75vYw8yCTJfVsd0JeOtQNdY1b4TRp560dDTS7gaGkygcS5+kC17pgdK/3o
OepVe1kuOl7jxAokeUvNEm1RTyST4o5/NMKrIVVo9b/vHjM/bDP4s4wOXpKJOXTf
N457wFRg3Y8y8rlBzhTD32XP2WCw6sO3ZWLPSZn99fnyIOcRJ0bRshoat10xIhUO
zLiUu/AyM8MerxH3EQ7gqovl/MPmR52uWNka0+6ghwEn4/JIO270dGfOZ8nf3BsO
Uhz3xLWwE5F0WRAcIuHvpdDI4jO5Vbe9rn2ivFytlnvxoCin8TkQQF0T4omPNQS8
/Q6ctyUuLeiA/Mcr2+uLkhQZiOb2GdslKCfCbSAGnYW7OM4roX4LMV8tLQ+Cm/Rb
+ftUUWBfXypA2y9gWW6c9dKu+TRf9Rvj8n4SVPupRgTKtSwB9RkB04M1uehDOqBg
NkvgRyQPF4oY4E+b/rQrx94BYBSfIalpMLyFFQI7mCpAYW+4Xa3Yb7kqpnz3TQsS
eqViJtvh7quTplR1+22WnzKUyn1uocIyvJBxJOoPI+HofW7KRzL7apYswMesjaaY
pm0efsK8gkoagR1GZR9x/EaMgQ0wvo4jBoBOm2YJjf3q85GyOsyGdd0cZyWNHAe9
WuAYoNEr0MegIdKyDmnE2SEKsUeeIVg/QAldIii5hMuG698WakKL4CHGye6VcFMl
rKVt6Oy5iVgVZWXyEvfILPim2P7CRYcF67qoqG8yDQX0U0l4sTQqJLWnmjoGlhya
uuT5WCa5nojBKC40S7s0TuY8d2KI2IlzQ3ff8UDDETnIiJwssxB1V6bk1JGuH/Cb
qVOnTP3itowMDml/iJNX5HkBAsGK3lmEMTCDHXYKse6NZsp5FJ8zTNYPgJyRd7tP
MfbBHekgQi1StGl8qwr1rgYIfXdbKwYtlMYaaPEjm7I0PUkFyXklZ2FJ983fpSSj
KFxd3g4re+OW2/EGSQ3XHqvlQDkpe9gG41vUvambqfsqdNg/iM4+RX/HguXI6ok5
tUP0Jzrqqs80sKvihSQWQ1Ht/MBeV/zj9utFKpqY0NKJOJ4PuW6O2FHHCiIAipmK
24P1YDoPJqokpRZQwEpr5Dki2iv36xxxbGV0mL2d8l1waW4TRF/B+d5hQvgZSdWK
B1a6XYjZyT2ajzXdQaBjc2xIPl/EZePBFMgq0BFbtUXiPIlb4bSdT+eAcIj/KdT/
NdVNt836veu7zLx6wx0GovWGMVuKcrAh2qlcMPIqdUPupGNo+KSIJq249Fn3KqQz
edBRSpeE6IR3A2StlPNx9S1lllbYcuiZfAx2o/a6VTsxD0w0ePVaiQLLJF7vbUfC
AhNxqSGVvrQTshuagBC0JjY/T0Vsf5Q9RR0BhY7WKAe73Vkd9cwC5enh5k2YHyeX
fGOZlH2AbBoIS/GJvRYptHYvP50Cs+8MHkPad/YNoymPK0omSDnnOjY4oycXehSg
knMpotQHiionPnt3Oj9UXj80NVr/uu1oOC1tl1SVQGiiOQKw1QiR2y6rdn3X7o2w
HJtaB5PrLiuQjtJFv9ErQzxpcxvLyybyWj6acWAgfSb44yWuRAD/Eqw96KnEqkdf
NfO2v2ORwcRj8PT2dwQ+PcFp5eC4Tc09QjaHkbHXPah2/VLdAVhT7lRs8KlV/9Ki
H+2g0N8avOVRnzAIv9jw0jOEBpcYxE2jdMcaNeDrX5yTuzt49XWgCWBcJF5pxxp1
xqDtam20S8TeKOnxftoPm41i8p8GrJBSssI8aA5p4WqEpmPkKy7tTmyskv1l7lM/
Gt+QRoxIR40mdaIFUf/5aurbgFKK8cPZhHGU7jZsKwgGyWErfEiDax456bfbsSJ/
ZW22eVLXBCxy3FPHiba7zLOdJ6dsvIrYwlo4efwUjVTUqTF3+s4Amog0keiIdpSq
+wSdlp4Ly+5DNePTfv6D9trCG6Q8EGrwBSCu0S8wMC7QkDvKSaYFivAExsRnARC8
EmbJvVQzia+q61QpsSrGD5G+pfrD5JDtCtU4TXkNftae3yBvCGdbsTjekmIkVvuK
f3WAhIefI7qxnGPKn5IHoNpMT0Un0gxei+XEsR2e3NfKrO+wOKoHQ0ZacC6rTiG1
5XiPWpj0nV4nDDY0nkSAoRMqIKlxyG6d+i0JyOePbE7m2RH3LcLK9Y5sspJpQyCH
UD/4L+BF5ewrhCYkrlIFm8lb1GTj7UloscJ1N1IHczRBvI4BpuLJIfM3/zXN5ccP
scOo1Pa09npyW4omLxHQHlgKVHObzSmMt+yni7KYg1ZDA/WMBRJkP962LfbFsiO3
Rp+Uh17lcWe5G6BSaZVvJs/fA2RUsv5CAW5/PLbJkeFqB6/G0M1Gfc3Ml+C3RDx/
EtBHFx4eavWdB2IvqO6LrOyvSPfnITywzQGIWavu/6VFisY8PsHoN/iJnIO1mQny
H7Kvn9OMVn2yOxjtAFulFzK/cD3uU8Rcv/tDPYmhA/im9/NEUloY+iiZAIvY+uEV
aNBPxZGErjl9sRZgB/Pii3SlySDD8wWNFThswXYj/jSg2h7/CpO0PuLShJ7Y2Irq
rXnLsgGqW4CbmPPcWb6nTkFM5FQwokONNhF/ZCvuX/pmXYhB6K+3cmKQ43Wuw6c4
7lxjCwtpwbgWqlktyrMdRiZuBpksqkJC2iDx0B3lp1qXxihB31/fLZVkER2YmN8/
evWQC/ew4J9HJWvRrTS7Vtc7xCBOMC/kpENUU2L+gZdggnyXg7S4dFeLQ0jJ8a8n
ePu8bEsT3/qhmb7HNIx9Qj11pkF1fNx52IyC36Kxj8nce0s4vg/2H61NV8q7/Ffr
9yXMimAJ2BpmdcHIzx43P/PRT0R8GQ9bW8Vrd1ZnHjZOzaDNSMRsC4BwIL+7NTpQ
kPEX2KcbFteoYDLoKYlDH0DaXBhMOqXNMHUq32uFt8LrPTsOrrlSErs8cwpfXG/r
bamQOezWU8+a24g0Gs8njGiv63Sc9CNg4WcnWllMgcwblbADtAK5Oqj1HauUYEQl
iAajvp+IReZhq2dUNTAXNagAzr+TwrnAYj1D6pJzIKniwHYQzAglrq5uKHksDx+6
2kfutjaKIX0lbsddi0d/3jpPped3FGceMbO0sbMnECHrZwjbF6/NX1nGiDEXeloT
bWaOLJ70DMGJDQluehSdSLFzp3t0zVf9WARfPjHg6KO3ArOtO0UXq4RzbsRi0cD4
87RSFH4nBtPp5U2xLOMHrI5YaYVsj6/Gm1OCt01mohITT2yct/741+CXgJIwJrVR
F8ZQaCl3X26OTC1kNNblJLDH60zjfCu1Q1j5yyC+i4uQ6BFYo730Oy59gsY0mitS
gn81Pu9jaEupUDUelkpr6hYcaQ8h2OAjMUc9jca2dLWh5Jwq2ZxKaX85NSTmEBaU
9OLFRleCBCAnYnSg3LNbBF9ONGzPf17qOffU/n//1V7cpPGPCCMJWICuRyJXN7qa
TcLmADnrZgiJzWTuVCbPsDTNDPgg8uLBUf/e299/7q/gkAk+sAP5An1Kua6hGsbW
NvpyXibsFL0KynZOF60Ej/lOXKVXMa99hXPF9daI4+lXJtb2dXmw4dyy3jJasjfN
FZ771gCuECKmSkBrNuBlSQzmE+6R/IXNTS5WAbXXNxEAA3YcGpHWgnIWFtOOadkC
cW/P26TsHfZLz+WHNUC+t1nZ+njjMcO4D6yTIba+6KPlhb5pFvZf3gfP/lpoI9vN
CuyuBEAnIHkxUHiX0SwE4uAnPXkyqv9bf39aNKOmDaMzPelTy9isgtuIfSSoV9xi
pvtbbBBERicuhvBUjzCXHfn7Or04dOApR4l0kAX2Ewc/wUp/tKl2TlfQqPJB0DXx
qg2zfR+BhOnZlHqZyWUZR7qz2rz/yzpWTttbWS2pcX+KG5GEZBzkieFlKCMB968u
EiWHcli1Deh46/qxt6vzfS4QraKF/CpsRg8vBRMIfKNsPD49MvYbwUlCieqrSLZB
+85EeiFlrvD1yORb9A/l69/ccGvBDNedpCSDZ26OdncQuzFkiBJqy8pEYz2dyE9s
D0qrsStlU8wg+pr7eegOPpzm6tqw41bCWeQVHTWc3ycAMn01zBgBkHnzMMgNvhG8
lBm7SYiNNrKj+w7xA2ekEV9el9ZDAffdYkTVTEZg4Z/gNODpfPjbqc1neOL0f/SB
7/fiAHAkJKEIycoQfeEqLzxvfYHNVdCieLpuRhORZIZFjqwm5P146EmRDFqXEdRj
1yuDW979h5fdYX/w+Ss6WP/cR3qXqW+/Vx8j/7Zuzoqdsi56c/XRRvZb0aWb/sZc
rScD4go1IlfpgzaI0aK3A8f5Be6wSxUVzYSjxAE9Uk/m16yDxnDbtSOYVQJw9diA
5O9+TdeZJBASqBw4fV69yeLT5W8TKBgGEzdg+Zq0nLcmcS7GWmOBTvIUPblaVA86
19B+iol+fT7ESsKN4wfXyIXX0sZ702jaaDThxVvS0TNAJhfDVrjH/Z+o7vVWjv1h
fbbSqTZWM9BfUHm2rp5xBH7upi+6jWTz2R/U9A0WR24RGZTETKTMAQZcNN0BVQr5
TXTv2p8IZplx9G6avZ8QXhtMFWeRN9THELasR7aNqTV7M7b0jnuzddvwH7Cd+mgX
k/hLNXfLeEh6yY0DAABlTEn1ysd/mzfo/GUx5BvQWg0PApWzoGtWSAqfGcjwqvOA
UOlbWwRpKdxHCKWHieIR70I2Z8grpuatNJGq3pBFWyttBYVNVDy7RHqpDihaKS5C
oA7PTY65JFCrCUfMLFSE5jk8jNLlnmA/aiSHpcxepNBMyxD1u9QdkHVruFuYY9s8
h4AGGPHz6jy8wdfYEyXusNHjnntoDw8oTUCTZkQqozG+PEdbNx30bFTP7CUIFZ/b
h8ANuQ02dFYFDFOwWTjO6Wu89/H7pCxKalSiEjqO5s2s89A0Cy52PAiN9DdNtYnB
FFib8LXL+NrNd39SkQjmxm+8rE3tSS/SvNIPerTUlRPtGUUABkp5g8chDx/ARwN6
iCpdiqcgFpYezeSdbuwhlVe1QrQaAqpqgPnuCnKwIDdmSX3jZGmbBcviMGZcP3Ek
GebgImJmGsWoP7Sxk70uLUMZbStm5sT6DnYg3PpmpWkZBrTSzBTgqwmY2nNwIOmO
Q4ZKPd03F04ccRyCwxfcs/swYU5BANkiRnzc8dJ6z6TimjcVp6ExzVHyHFchED0R
a6ea7DM3w3cmcM8vJleSjoSZJ6QP0LBMqeWTRbWCPpUSrUNiwZWPs7PA3ZQD5wDe
IA7BLHMV3JCCLNmrOSyqBFakhe0g8mWYWJZQWe4dzzZl+eZONlahQu0mv31Q7vRD
ji6GrM1Q/ybdqELowsKmFck0sNo1j2OnVf1oIyC/v84GH1dxO72waaq7IjC0Bj7T
zXcbec1LpQQTjMBBp/R72kpkuNby/YmVMKxkLXkiSHE/eXz+KlMAZqCcocX7BRyX
YFqYziOXbC+ZqwqcHWtuS+LYd4GSsJYZk3cZlnjH95grOHGVccnYVKpH6bAQJEZz
1oXkO/b951RwN8s9avRr5NngbJH9jTl+3A63O+6OnAm/JOjZ2FJ+i/Qt7e26OHHj
BKiefh7ZMiOmJzSyrO5CLZp2C3RbzIOrb+luTnFMdJCJL9oi2sl+2YxoDz7ISdfe
UezvCvjh2LVZvzNZ5jXQBdWa252zoLm+umZxYGPz/EyLQxXi8A0fkHggJ0ydfa4K
LVv2skpAepAZBu8EZaYGr4v69fQ/ad/3Gj60wXrAt9ONU+M6kLFGT9+nifBw8PKG
RnRvGftlzySZGNqw/5Gqzfu90EY9fIPqcB0Nofjnn7XGt9rbDP5I/htPI3Z+8mgX
/CuJn2w2Ecghb99wx0O4GEdNACoFixhC6abzG8WsOWP9gWPh2xc5UEBxLxjPoluI
jf8/ObeLHDfn+HAZWSsntWPcAGioK6jo62cZ0AX3m4mIs7u3Y9WFZm/yQwzpJEU4
uDj24rN6Kuwd2AOaCE2sMPmdoJBUPilql5O8pUzLFc8XH6ScNDt0UvWVTzqlrnmS
HITNIWsnaweCp1YziQTwaKmt1uuJ+9gF86G6O62dyQQ8YPDasqMwtfv0oGH1xSHs
MCdA8V5ZijRTkvC7ZOleNYSa9j2JNEBkMEDhVRMuFoiP7OkSOgEQmlF1DMmlT8Jy
se3YcnZTJ9zrR62XzDzfIVbbojVcuZFx20dY99vHrKJpZgLKdQfCLJai0nbh1JuY
Ba4nuXi9wPZuPnhxgpvsW4GlbBxTEvUMX7grKbO98uzMXmO+dY866tuWIYpWoEzS
u1ipI1CulUOOc/z3mV1+8BFw4LbtxEGX+Lb/1QZdGdnHMV1x2ZrH0bvy0r6E9B/l
vhaS/ypxh/gHESBVR1n4OurRG0xNB4mvzzEHSBZYxKnJ2Xf+6Dbi2Ka1XjTG89Ig
EMfT+OQNfZOHKGK7g6wx7nkWL/mR2FtRBR8ChPnmDriZ52Efk/orvyB2u7JiwMsV
Y+8Zu6XsrNh6tuSBUSEsjJot2yNgOskTMBni5BkOPAluf+XZwPLK1iZcPNv3zGfw
aS9lsMoHq0rlMV2nJbf3uKnWw5jEV14eG1IIezrl+cYCLfinf/JsoRf8agJkR91n
12QcS4AGHMu5dMg8+Bf1fuedyWULijGI7KIxmauoA6XHFiXXg0++mzPysAlRWjOh
cVEKhc7X2/ZCBUxmUTn7hOY9PMtkNI6zDoEX6EALoXHqGseaRbY84wnuip0E8cJ5
N6yL2d2GBoNmkARlS8929mo58axkQGYmfbBNzNc75LkRryfcjdkctAfWsvEYPabl
ZVsp2mayEWFC0LB6YB3Ubg/d8nWIHnYI65z6O7WD74L0Mc18XHs3pXZLFBXHsBtC
MpUbyYF7dVZiA3GEiu7EKjJCd9ht7jy1dYUoizu1ZRPhOWk1m5DTLvyzwSi7dcOt
mwmCuTWE/T7Kmejz9WWSv7miMGInPbz+MXS8pQ0TERQhFUMO90sAL5D/lzsPhZoV
VxNJ+mvziHtzdy3dSLw2BDde3hUSsV4+o53Y6fnyECfWmZ+uDOZi114llVpbhcMR
zzQaWKj/yF1022BpNwjGr4cxRbQhkDycALhOKOa4hpWQ7rIdkxRjs4dZLYJM9CVR
6gXQBFNyVtkaYHTr8Ztg4x/IkHF0h4VNPmkLtkccecYh5hG9ayeRdJZavBSlOMdn
bk26e9yGtfXFs8dKi46NPkGd1jFwdZ+YITunKn7zoz+vz6dG1uBB6JNO+tHAWGuU
BuvUQ75tEw8khoRxqEQ7Q4pLOG+gR/NzkGrrxaKaoaVUvgFTURJWZXQfKX/POgRx
n7xvVCKnAiwyHVweWVyrf0FjbQl3o3fzcA4WmiPuqt7RCjsMtYOb4jpuAjt+xnEh
W2CTW0OjQPbQutRu2424nAHRKxNMwOrPhYzj3jvWB2oxW6lHV003+/PwOscuEmk2
jvWnzdsQTY//YegledqGRYbk+Ovl2dI5EityAKkLOp/sZ/Hrtnz446FmYReS71+f
q2/efOCiADZ+IA1i3JymiQvw5b4OBz+pCHdhTHEpRK6+YnMTbWKl/3lxep+JGlV4
rozNoLAebCixFinWbeupBTjsv4QtlXWuBzJ1ctz4U7MBEVlsalW1tUG7f8Xg+zjT
jpOv8o7I2BcDOZtwWvHIykwkI629SDvD3CBhBfPBYuRgYg3XpeUHzoNsRj+JcvTb
TS0SDrQB0kARDIaTiFQeX2M17xEOF3J4UVFuQGEUFtClV412vA32TWOO3LiOveoX
zIiHR/25vWCjNGZTJsxrXBI1wPLSK0QwUBbgFGndDb/dAao0C3+am2DnCtufvU5f
Xkf3s9xz6lP6CiP5GQZJo3jTarKh8XDL1kxrRAFRz4zSPgSm0IxVFBsdlRgC/U7r
cNpJewcaXwKdv7eeHpC/iE4N26ZccxXNXAz2iBG5Du7USGh6DrF7t2CTCGZBurlz
dCfoP3HYQNJsoPEmemFHUWt83VyMJ2z0gffh5mE8tL+Ye2hE8oGxvKuuJz8djTx2
iG03p3254q3CyIJHBmpfY/LHEa6GFC9QzSN+nKFRfu3IcytN7VdhihkVB7egRoXl
55qysh7cS2tO6pBHQW9j1Ce4TbRVcPQ475uazEFW8wacGXn0R0LE2G7paj9An3Vp
cEhb8WHj9H1vKSlMeAXFmasEV/77CFGpZRt9yU2QDeymOO/1yCjTxvWrhOsEaNqZ
jwhQqIx7lV2hy9gpLk0juPeSAmJ3K3kY7ilA3f2hfMJyzmNHnhlq2mPqBUPoyu3F
PYAaFdsdKMkqmWzE9yhFGIjvYq5j4XmLoADLsiw5J8BCCHqbLeqYNtU5OMkOd+i1
4sfhy6Kdcg+XFwjxIgEJsgZ3Z/Yrws2FzAZcKo/dmKHx4ptvUEixWD49AZOEhWRA
3JCreq86I8FoGPbk6d9M0q+u9WRpge8MdyFD7DxrH6UenGtjwUs1ISh4YnkXdiVT
roUSOK+ovVE0HMCXSiXQn8Rt/dnsG2cMTcJ02A9W4SZrmU4U1pujbdBnvn51vJFC
ynxjppcM2rKuOBU2JAUG3K5BOs+shJSnWFGA1S4Ggl9T9hQcCfi1CTUzAECdTpho
zoIqG1LmsB7uT8PGKZpwGmbcw2bNpxhT73xchOMD3ph43S0agnQ3udkT9gAXI2u+
cyCkXxQP0yWYSTnYEEXqcW1K+lQePEB8tY6ovYiTA4Bw3OXVlutf+IZrMBy0S6C7
tIhpbnwPpRtYd1P1TSQDIi3k9fFN4uPHF3TAwanIePLh4B8/n1jN0c+Mls2C28gE
qTC8cw67wA/99zAL6FGxWtxecILCoTvtKEvEkbjXz80VzKnshO1KigyF5CIiCxuT
VlB5VIYal1Kb2SuRibK/P+I5l7ZSk6B7SpfvUfHNPP1ZnwBcf8VqzQEIOScpAt5G
L2ZshVDROo0qBRIpeKKPlF3LgE9LYSBNFitR8Bl8kyCKIFCOwmUxH5l80AQhXAkC
lyPrAL3uGJaIqnXTXb7x3HdB9UC/fVash0Eur6ry7763faCy/kae4WL9w+n7ZIAk
lP9K0Ay5ycpm3JPBL73iTmwl672dEbfzFpQsFs92yXbzw8R6UGb9TFvDn+emWKaP
LN35/IPmufq8e7wieTbh3a4gz5ehqRbZ70BOCSJR1Mg5fMNRVYu9V/5k5Kcw3gW5
JxVDao+5/gJ8gV8UCypoqypBsWsCwnvjUBuwZZir0ryRY6WrjiJYuzC3b2f241H4
`protect END_PROTECTED
