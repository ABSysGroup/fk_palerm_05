`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Oz8A5Hgm37kYjlfhnrO5g5g+2L2hGGp5bfTcFpojiGNVUuNSZZxUqOUWXTw4RwO
vhmI+r1LFhQyuT340hEDbADu9OimiNpPPvoYrcyUdglTKnD6nIZW7TwhiiRCT0cs
9hT5dLcdGs0h/vF78LC9SCMoquJZ3gh2PWa8ERCZ2e5/egmwIQh1DcKpPLDHwRg6
phPd5k0YK2L0gYYvm60JBsaVM7I+17/oQH4nbGtz4VOwSH/jxr0oH4utaJWYn7z+
LYuYiBYgAHTL43jqcYEsf92nALoDgs7yyFgcoHOiCnxmT6AZN+cdz4BEHDLdC7e5
4fNvqz0L5b7vKOPT29IBo+95cYn2DcnBXFsBiEYScH3I+Uv+pH1K91CBSAob1+l7
mecBu7YS7nrccAbAxsQ9RaNIVyEIUvwFY8peiBKES+xGvVdOb1/UcKdTzQwLSyxB
8CkI7M3nT5uSaFia4W6pRunEJVc2OKj8McxAQWgtVleCLrddTTIlPLiEcdN8qyKE
rnJZrZHci0JZ4Ba/cOPhUVV1TO/I2blXu9vQJiYOmCMpIKpIblr7tcYAgNvcGmbq
kQg20LWNw2xZCgqUPGlBveforHRpCfIFwren/BPFw/fN+kLEWF1PWO1BL5QnZjN4
3bgeYRBTkQnhKxWwspFns+3SI7z4amVi7Nw+Hp3ahahGJNxIsIKLMeIAIr3/Jcoq
DFQXBUBd0QIS2Pfv9e0P3hVnUGHexv75zVb4MUA4oLR6BhPRcNrdcAeIxDDJ4ctz
NavqKR+26jABZb5gtKV8Q6lUARQCjAWN5A57dGEWRM4tb/104S3Cpk8/0CvBFOH3
cT1VdS9bvgLI0y2jGbb1GI0dzE4hW3T+rGhqFmnHT3r4UJeNdhUt9aM0QaHiqY8S
nfcHQkUE4xldd6i+UMOZxqrt6YSCDIjneeTb6vJz/6l2Y6W8JTMnYjvFkrEIzymH
6t7GRU5Xr+mS4j1HzjuOQwcqDB4sNrac1ZgKvi27gG+qelnvjcItk+wFAteRGL9d
l9qzzCPAQ3iSVzOxqz4mCJG1lJh/IRZkJD9qpyLDuFIzWN6T4vMnIl23JdhlGSGp
jLIqywGjvp9utXqeLF6+ZwP5RRmdGiA1D5BRWkkkxP5tAvQjFX7GiFkxyFnBLzj7
9iFleg2xuh7ntQsZDoZHFWwBdt+MBakEX67E54yZ/iFdZ1JoVDYEGhFCRoj0QUMB
7Gnrj19kPn0zw91IVLrU4uDNB0vQ60qKF2r6S3uvwGtprR4CfbZdVveFSweoVl+D
YIsmhN9fhH+PALahDRQDeY0rW+Mnx4iyjgqa65eyEMHH8rWjbPxq/fYbSLNdUM8c
UQRchdL+VfF4IJo9GGg0zjDIFXlaagF+tFISXSZBLlJZUsXGUXtLYh3AHn/cpfAd
HolpptzzAzexl3ruqLQ+6dAtEN22g0OFOAKbL1xkjIBc7osbKG6BT1I/BMvyzvdG
Mn37WlgVjd2zR7j/1PRTG5g4UWtFHPGpSxFIEx9LjutR7FsHPR/RKR/rD5uqOOcB
J6nEAZwcNi9Y4hpQ/6s2APDHKMXHG+XnGJrxHqZ4Awfv30T4bZmpnvHryn8RZFQ1
KFyHTK5g+90H0FmXSIkTWmJWPlz1XIytro82SRvLjNa6GQ0ba53Wvuf5nN66bMse
Ol1Bh9BE6zXMzKZ3w9egSY5Oz7IinR6W40VJjhg51zSP2BZ5RhZbOY28uTVaj9J/
7N34Z9v+NbBJFqJb3tRdsfh3AcrWDCz4tLVKTGgQ5LMStP/d8ne4AogzI57l8VN4
d0OtCyg2tVSzvaHIeBT/EMrjDFUQq05hef3HuCFgBmfQBvFiIwz94LD9a/DgWSDe
cfYIDx4lOZSoRyZjlsOl1X7mEoh6dny9IjoVN91c0bpb7sRTitfF9qxC1GtNLO4k
Dt6xPRBUawVELtqML2W35bjirmgHTdDOsT59Sqb98fMCIRAjV2yZn438hxjfSqrZ
c2HECoiJVj/yOopwmOGDT38dcjvkqLxjehMz3JjJdDRfR1VRqB8519ZAS1E5br1w
CFUFiomrfUeldPEK1YwXZU9yp75o+SMlArCLDhpAutyf1wwtqRto/WvspprJ+7gc
Z+WR/X5qqNfI8jomux7im3RHQvpDi+JbkaKpdnRMZbkJ276WIrsOJr1a6UN7DQQg
jNwYsO1VMQJaaRiByASNictNElWyxLY8tvYrLWBRRqWGdgfquQ4Qh2tFekTU3Q/l
7DfIJq9gkWHUEA+jkuORKH2I0lyOyj7D2sIgYnJiZI5+vTCULm1D6QdlcUCRHXho
LCsLnpF6Af7RMA0ZYTk6QxdqRrNcVd0b20Bc4W82wotxdK86DaNi2/NFj9zhMTn3
ZYgZ+0Y2zyBUdMH//Nezde0Fk+Q28H0CQ7JgZKraUgXOcWcJdZdTz6Ym1QbUu/XY
CCuqfHeuLPtWzSXpviCRnSlTS11bJ8KRH6hbxwnqwgtlxGDuSWF+gWDY7Glc9FDd
Kjc53HcATvz2Jl1LO51TxO6KNndfrqQ1f0SyDLEmbC4AyIiDvM41/nH6CNedvv24
7TpayCuJhd6BtwAWiRCh63D/aBwRmk8c4X0AR2ECUzpTJYrRbBXPy6xw1O1D97qc
PAr2RDhu6lh1s2UmBF2DeNikrQBoCY7m2LLbD60PAAE4IQ41sdavV0sU41GHR761
vZN5248drGoNDQIRA7g7P1xWc/TGOsOtFa9ePdMi2ZrKQFpIbqcPuiqF/I41Q3Jf
ZNywcxuPS8da2GvJSvWqqn83uPErYW83RVhjbkLHuxwlQRmgNFvtmFxymtzTnfAV
7XNsC5eBYETsQns+Q1jlc36+Vbk8QvyTcmf2g/yvWcDrdgelvAQuwP0oN8jQ49ye
/88D20nohEAjsotnEg+XOA==
`protect END_PROTECTED
