`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
phrifmGdepSIVzJ68gl8Yebyh6luXAqqI+Qz9HxqLEiyqB3NRZOjUy7IZ9lNPnx+
FG+NqOy4pe1Emth8SEbTfE+gws+djYOpVnyfpYfHtdu96qSqoD+x+NyWXdQm9Jmw
lCB1fzlaUWyjgob92pVmiNlGzkjGuo6upOp4/XIcptXLuHhHSwLQqVqEGVnuuzK9
6+mrmCh/42nzDdpd7gXX+AJ+OAS1Xz2qaMU8RXpnbZmP3coGdiRzNT7cTh9r8EUO
p2GVwdouL/ouEFU6FLh0Lw==
`protect END_PROTECTED
