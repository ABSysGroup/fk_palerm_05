`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OjLk5uOZk7ZLl3uJ9m31JqS4UXntF9UE/bt7ZaXxDaKEuuxAiGkeyaNEQKWBP0rE
ferAiOTcBxjCbf4FyTjcGKK0VPWUHpmAqyXdnKxy1JHZbijmU54VRY3UnastswDm
qKai5D2kRijZ4yfs63t2a0n+tHBdyslkN55qv+FVtu7W9l/DnPxDaR7uktVzvyGl
gR/iUNry7eF5o6laDtfVXjSCrkbSFQsgC0RHjIjJi+IxM/i4bX9dH03HVttJO/RU
T2yzcXeI8nSEVmwuvV8E4A==
`protect END_PROTECTED
