`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0IiZLZwOq0AKmJhD03Kw2t90fBiB4QlCXFkHilaLNiJbgc6DVl+ZxH0AGevxcveS
Wf1XuKocM/8LwlNXJ3E6h/TLCFn23axrrWAf9/uLZ944seUv3J2FkW+DjgXIa4US
ZwTDl0RTXB9uY712o2jDTyHy9R8ol+uH/2O2kPR/BF1keet/ts3uyNesckmrGePX
SgmMgzBAZ1T0HdJMQSYTIhYo9gqfL0DGciSA90M1RwubJsj8qyn/bR/UHpcj1RK9
nzurqqP/pfFxYOYtqwHjsMNlzqTjlw4ZMIDLxHIlJU63O/SUWo23SHCUAEmtYfop
DsnzqJcFrckrrv/FBBJrSM57Ee13AwS+fiWAb0r3jDCFcB+DAPsDTh14lzZ7OwKN
ebkTLe2a0CcZ2XXFPDSXf3u4GgeFnBFhUYbnK3bHE3HvCrMCyUYu7ndtQTYSqWXV
1NHyVgQIbc8Re90sceALo2aoJ1Kl7ePhegKFkyJ/E7f1StJZ8YKMvvb+Oae6jz34
tAfs5Cbq8jecbRpp+SNlba32gO9HWw463XLXyhbviNGeD8qDD/4QCTQ6JEE4I9NC
uRjgQxZU1ERoVkxb7eeF/zEBX8SjBDK+9kbaCgl8walfD1LrgA9rrPk0Msta+T8j
k1cvAVTQ35A60bHCLF0CQxw39T48licaXicC5qzIdopo5ax6x1+dUOxtn3YJf4Qa
neb5PycGzDHrjgDx8ZIuxQe6HD2ty6+S+VIKJrmODf7b1/IQJqXZvdeD2pAIgeaz
ZR5OayHp1CgUfd+OI9k9bUVFbcQYn5vArWGi/AJIsOJEZZWJ4qFpfL4xDKQ9yZ6U
72SpS76dVgOwWKfvkkRQgEspO5j2MS4wX5N8NzuHF2u6vsE2p5qGNtf9ERYtbTT1
ETHpQVZBc2S+8vZwwiSVCkM88lSNRpysHGDMWV4VSg1+SA1Fv+jZT9yeg8UZHyzF
emCYiJ1NgLghPJewpgTr2VQIYly3WoQnHdVfB9z1qGFEU6IW3zNgK6ZE2ERoQYSB
2igeEcEbF9gnavcEHOLG3AwGFFwm8q7U3fd1CBxy7t6dmUnbwpTKysvQtO0ntgw4
C7014e7+ea+DeFRmx+Lo/f1+hcvAh3YR64RM644O8BVYXYiPw0uvKqqZQRInZGsf
ZhXZCAGN35lmVSshcTcijQTCAqbl938DBbJFlua2Ffi2QGmt9p5K9+jxtPdfPW/Y
zPMb5Pz1p/EutUjTkrQVCt33Yge7OfTSIP8MqtHYgNChpnco/X9dpveLKYsQMCEL
uBokpTFyFujgjNjHUG9GfMU+fyICLU0W6ApfOIhvaejkG5e89mc6mINSZE73a1+/
DOemqsZoJgulgK3CkUFKhC9zXhKiV/KgZMQleOD61ONbif9FzRTMcC6xAk8ZLAVt
aAs48tr/18sBpVTxRWpaG9lLC83x1XAT2p0eI7Nnozt8E3MWSdMecsoJz7+bYCAk
CtqlNE9TWdSwKPaXeVSFZ3I4K60fojoyFoGmbeh1SAk0m4UyDkgdn1MO5lFsva2g
+nsfZ8tYUvFuZc2RdkSAGQx5d95HkLlW2toohppU7OY8K88z0i8my8XuDN/mRbnC
0DQ7YJ4Y//FssBiNDGKQr5wrKr/q4iVSkUtPs79tQ8bn3GXteNhw3oU5oiZfjoFo
6UGNh+0gprGVFttZG+T/1yroAaVUwB0Qbie1k6vYL08UfaBMYm7sJLPT86hxTBTp
jIgdlf2ePQaW/ZAEPzRAcTvxiVeezCy8snf07MryXEKYa/KJnRDbUNRRGJuSYwsl
ioauT7OvEFvg7oYTZJo8Fg+lCZxHL0mC3WJmFcju4cTyy4g2Ra/gOsaYem/VRbDL
axY7c7KnAxuvGPiOBHUNRDWHaTN7Z15BJsXvbqUYAnhnYPw3kQ3YsRv2peX/sQgG
xJ15I52TM/xuhYB9nF4iQMyY12Fp/DyqHgjYny9ZoMl3wAKMukYJd+WgqEYGWVFN
ca+1E6CXleRZr0bHVk5siwlpujnLInG+lr6F53m9D1cpwJfvcwp5CfXN2mBuKNI0
DyaHYnAmTga7keaxgbRy/3Y2ub/eDXNZ6HSTXXWjLznXKPekf110XOavYcXadLRl
PhsKAcTxnTDUyJ0NCp87mdBUt9Lnu9YV/rjSR3dlLowzHyL/WQ8KnCKkYoKAcYxx
bWXNL6asr8ymCsmSQJhyHDi3cpPFbUkr6v09vK5ZseCp3xRXUrFCHRc4FIFKKfLI
xxL13TYRN+ntprKaBydXms1P1vzL6P0QWuikOdhEnz/rRUw4HWLTNWkC3vD+WvN6
Uhtpv7C9+y59Tt3gKNHCWHWOZ8d3nOO/2bVyrMKovC98I6TMS/WKvD1opc2Nnp6l
WfT987FRRobzxJeQO9W0O+ii6+9O8F+ou4sBR6mlc5OkLbduZ/ety3MVdEShmqce
yD1ZPeBo6t1cqnFbRpZ95JfcCvxy6Kf/sCey1MidPx7bI38E5mKUeFNEB07R6SaF
lHzH7gGvk683BOh25bw/b4R2h5BgpgvaikzAnoshPklgWeEaVg1xghZSTz+KWRuA
khucenZiHXuzTW0uAao+ffYKv1BVX67MacN0goXUJED/GwBPQlcCpccUuejI7ak9
pAYhknTw46EhWASthnM4+AKt38wLqeXPMo+xJSJVD0/b970AiAEMCD5L1MTthNcG
pAt51R5DTraJq/i9YfCoOwWLSBMMTkGPJobodRR+td2DbZ2HaG/4szvw45erDfLO
METdi88x0Pj/2pJSP8z5/2YLRY/rbY+RwFVnsrK3Y4QYKMDn5ULM3FkUZmMMhV9s
i0qBiskQCbemX1lHEO521lDHi+T+mCBkWgQxt0ueCEjnSQaHQ/2MWS7+Wzgb3ywK
qrgeXCZDCT6Cfz06IQ7g38eJmEHH6SSRnSr3mlYeMewsP2STJoyK9Tuf0tHBS0QD
IT9Fww8lZ1RTec+82ZbmIg1S1i0KGlejt9o43HH9IgQQB1/Y5ySXUttwNairuaBH
GaLvp6SIFpjMLGRT0LEfGJ04GCgEC8IWp6wC2hD+ho6UFC4Q/qczeM6i1pNyo883
v4yKSETO5M7ydwSSnwbbmgJDnqd2TE2R3erRQtCfg4tNz50btDS0xIdJK+4zQC6u
UU0po9Ns1UbvKnTylEzK9xIO1RYDJE+VDuzhJSscB5ol++srpE2YcwaogbzhD4+f
QAviywifMZL7JtSaghqCmMJHJE/H5QInmrQo7Rfp5Z4nTyJ2+xz6lRW2keqXzh25
V/q9jIX4R0LlfC0ADE3Cj9J2PfYYad/wBN1+yVN4eb3n1H5+CmbKmCWMY31YTum/
wgL7dMa/q96P3KA6SziWmjVZ3iccK/iv+b+kONnVL5gAvnfC0wyAQoSXdEa87/xw
RsczcsCfXAlqVnrf9cpX6gmHjG1iPPcWGiNG8CsIm9cAv3Q28skhZqIW0IQGoM9C
G74KyrxtZ+Lj1AhaCNUJv+gRc8AOPWkuKoKhzW8CjCDGCZaL7CVjksXUPoyyRO1X
4i5vpAOXA9EBZ3cyFAe5hx35QSY5JXtyOSucpsLoGKVRFfldiCVq0q97QDGI3ZBA
om+iVKdw4qiAlxCagi10scLMDGKAkzSKQDVSICmas7L8UC23G6xAWXYGV8FSI2rK
goKaFJWKrdNR/s9+oum1ow9uyUQMMuKEEmQ7tjc6yTd4ljcOt8W+3HOA5KklNw+e
wb+i0SdGKpkPv+VZWQJQeXBG9e2mkhr6xCItaucvR5XE0H4dV1W3GOuVwdrS0OsY
P926FsKEg2/jXzYtGh5LA5mDdE38BfZvZVkNh+IgtlOhDHLhsrg133IHooUM9IB8
+TOmS/2IjpHCSyD97LmZdGqIvCU2WPW5WW0DaZ7ET+RkR/Qu5S5FhgHpME9htuNI
e1I1v0KtHe8uMYMm8Ixqd7tMx4ANpzej2pjA/LrehT0XtBusSNYB6bDF/Lg+Mjqp
qc/L7mD+lYCk7taZ7IsGc+JW8EfeEBNKbdRYa/6M7QNXNd4/3qSPP4UhPdX/BArM
plkdZD2iMapUfwC9CJ4ASF6sNJL9vnjrtNgNlWWecj7tyvpQmmOT1OOTLgy/AfH/
mOF36v/Z5BH2p3OZ1G54faOVUDZh/Wex1pv6IfELgeso81z82Hhou0GBmLEqLL2r
3RHzog7S5jZVK4I7iUunpiPkybBOjGQ337eP9Pz3FPOHTbmEP5uG9I5vNIhvID3Z
MPm4erJ3UFMEepIKMdY+9aHoX/785w9W0YflKUuSdxdBRNkHn7og8/zO5xQDzrS2
F8V65GKKZMpYF/CrNhrTCJ0yXl1Fte8LWQH+8EyDFdOKmjUH8qC6bT+Q2IyhQqve
VaZWkrxV/I4cYRzQUK1jaTDkN1WWQu9yCoDMzNkRG/WFxVDAmE8Ka5DFx36ADbTR
qmnWciKG+5HDHoF3TMH1bLX35JStZQl/lzKpiGoYbu4cqoCJ8Zt7lUIJQpgcH1Du
77xFufq9lb/YRUUugWfLS6O3pgcVcXn9hn8GzYXmaQQwAo+zd1RPTdV9bhHcb7/P
gMwNxSx/q6EJ7uB0DJiSQn85Nr036AnEA92nlvoWhEuVoRxpY+LiCzHTwgn2ByuY
7GBGcxNfsA7p/ISaQxsW8K3n9ijRsqIXk19b+MVnh3G7q5Xp7zAQ/5o0ps13kfI8
dvzX/0UpVP002++WuPSXxG8SujYGtySk6xctWxdYFWk+CjbbjH8yT/4fOIwV4rDR
2rNphnpcQ4LUXerjrNr4SZ/f7xe+9YxqO2RPwoeT46dZJcJc48h+CZWSANlkL0Gc
kA7mcwRw9SXvbGzoOW5aDAARDmQjOnEjcXltOQ7i5chl8zzNULqjlDlQrNI5BZUz
aX5L0g9Sb/p78m5EGbU9JBLUY68BlFebieVy+Q7eX+x8gznNjmpFxD5vhpHC6m2C
frkhKztJfSI8RJAcdSPrjRAJPE+9kZzPzdPyKaMBliw1JAm/LcpOcv59uwbRzXN2
hPKk9NU4K9kHVRh9atHh9+ayjwU+4/wM5aq/lppLjFstpND/Va93AmDd3Wy77W3M
euex3/FCV1M2rfqeLskMLEca8dTRlfl5ALFWtMEk5uhcx3z83ijcrzPpg+UynaHR
dqL7PdEpz4EahE/74Z04Ray7JOHDGxMChk/UpY3CgB4XbXURuyPzhxU4LswZLnT2
BEk24ICT8BaT5hCtnk8wqI/OEn/1bWFq+MmlpflQMMJ3dugg+hF6+qmpzTrfs+C2
LkdVJPZxK0bZDXXR9PuhnuYxmAupN/YRQCzUTVY/Hgfigqs1lZI/oXldxtqozK+G
yfdp9jGoaXPp5CMOQtG9dzVbXjXkKDrTAxpdQamyRpHaIrVo7EooiXdNoaVkWLZz
nLnArt2yC8c29kJvfo5rUvv8fnaThku89MoDjssjoUamX53KYcp+E6fQ0UAeCbFF
/Vrq8qlhTYuP8m0TNU25moY4zLzFvzRTDQfroPDq/OR8UK3aBQUdHJ+SW4koF6w0
aBwkKicqJS1UO0SqOldpmVatjJVnT+NZL2HiaAFQBTIg/H8gGkB0fOCSNnh418an
tcWUNrwhE0GdubAvtEwuGLdjZvur+t4chjnZ1P4CXcRZmsPVy94KtraJTgsZfd3K
PZTsaVILPmDRn/LMMp0Hv3jjwxQehtDCYZN/TtMB6ggY0zXf6nBt6N2O0wfoy7BV
3C9SqFLRZQ5npqQPoiTc9vEa2ENiLY0xrs0mlOACVfkvIRuhE91oH6mSVmk3Wv91
HIodt3+LDAHSTR9mV0r6eVfud2Qet+GI9NqNExd3aisqmYjq686ROLnqRZ2pMCRh
L6hXBx4n842/IpVtohz0nC+GBCs2djcfzJBR9jqW5OdwbSBjX/R9gEopE5xjfE3p
7ZplziB9x5zRp27Z38oMlO+K4luWzFYD5ZwfqeOgjAJoNdzWpVkNsTLIjLhrTR+e
BMMIHZolhZjLXEjB6zu8KlTqt1Apemy/PePS30jibCZd9mlligSvxCvXHxCfIDVM
HBPVDk7+MR45ZTKjLD+p6PVxZastjrzvhq1X/MZgyETRU+lsDcUPt7UUdvF7Qit/
E3HqmYt7vvdIH+wWpUty1jyk2apFV3l3jcT81Nt6XKmbM3MfNGCGGFBc5GFs+BBV
iCJ5OzJa5Olzlx/RwIe/1urEeyN7CPL0ROZevhsew1WbZlTOKV+mHgnPNXDdysTv
3wuWT0thzS3AnKE0Ukc4EElVS3NBMdVgBoifIqXcnm4Z06MbVZefMKerL+8Rj+sF
4xB/GzLWj/aZc0MFZMPZXMBdRy2KsDguUwk3CiypyalvdPe0ORkFLp0OWiP3MbG6
kyfUutQY/1IumZdOFvzINls5dBB2xfLNFkwdqdw3DGLWkd3BQnM3cdFQAHlSNvHj
B8kIaoy47o6t/HFHJPG93cuRsK0xaHWUaFRsDehJti2/RxbTo0uIwyTloC7DRjOu
0NHGsaRZTx01NAZNv4fR3G8x2i/nSDApUc56uiSJQKut9jee/OTy1N333y7bTp4X
2yT5pv4EV4eHk4rjfmS8XVZ6TwyQ+YgsPcAMzG6nsIM=
`protect END_PROTECTED
