`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tmWXnx4UbK408IfMWfKsLxCF1Pd62NKCxtJHXAH4gk9aa6Jw2QT4RKlRzqAri8m6
8Ecwz1lN9XOBXJjTml1Eqro7oPAwT6OkIYJZyQi4TTRyMTCK/pKdAIdRlGMA6ntg
BJceo24F1NcGWw7Ycomvw0Y/1aKXPTtOK+GWBIHJVrGkEKpB+dvPr0gXPWLw7iT/
hvSKg6zdoEoBwqPFI96q52ueKn5r/GNSYeKuvBW2MrCo4K67dCBQ40MbXle8+USU
IZcbVFnlG4KA1PApd0U783h/MAtRtVyTV15KtupyJeL8QtgJD7yaDtkxFfXljAU4
6K8oDXoHg+JqtfdUzRtpOkB/dj75y5cIcuPSaxVKs20=
`protect END_PROTECTED
