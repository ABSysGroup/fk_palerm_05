`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cXntYT8f4wGX7/49JRovI7g8m1zv6hj8kEjEf8NvCUZ/UP8F8RlVsvioOvLHqYgj
xiJVuMqeQhLsr6iNg8uqbsy82lYLMynwAx8lZGUuo7ppv5FK7zAKEqFkpnDSqQix
/FLx8tJKk1hU34hjHA6p2DUwtD5qs/Wt9p2U5uxFkLuE53a5ouLmFCua51ZToVRU
2LlxfUFodesWHPTFhquaIrwIgLgF/52PW4GV9QD0Pg3bBM/+CVKGoDwpgbXBcMxi
`protect END_PROTECTED
