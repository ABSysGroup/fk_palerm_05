`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
boqf5/mHlIEQNqC1f4Cu/vh326Qj/Wycn+6yG2lwS1IuNGNjsz7IrZ18LW1mNVLC
vHrUbS41ppP9t0/AEt4NTkUtUcuB9SkYGxiyIeRa5gN7Q4dJrTwP5AnGHW6LRBOX
3jGQ1bLCHuXZR2vT7FuLsmsClVfli28gThU6KW6zVRcYg+44aPBpZK5F0OjyjcO1
2RZvi8pjJXZpHANhn3E/InB54bZWwy7vsb9rCdGswIH4BHhOiIS9QjW9HCdGbt9P
77qv+6A2BuoVQDkr+3osARTD4u0BsAePUgnxoqLfcRBKQLv27V7ltiWOrW7IRqse
1xtVR43qg/DRlliN2qXIq5zcFWkp7ECTDZEznOKoyjHWtiqwKkzkGj1IVN5up8Kf
`protect END_PROTECTED
