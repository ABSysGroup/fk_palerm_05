`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9o2aKURIueutrAq7ST5o8AfEsAvtdKA1UeTCyumwrSyEQ5ZFZJF0F/n8DSMkP6EQ
2U3z/xviVd5jfXqbaXiN796+jVAYHLJkqsTRnqJe+P5ZX8J7naJLvq9mdsl4ZK6D
Bsg1V52gKcoA0DQiuv8wC/l+k8XWzyt6JvsVMUFpyf1kdfK+zI4yWg6snVNsqimI
wRCU0vYB62WEV3uQ8FV1ekpLybmyk0YiuMslsbMRXZWLtrRgqsL/slKDIvOnk81s
aY8PB9XIAST35bJkWlqk6sxMBEC7o9XYHantBJn3qKnbukN8XAeTWcqvvd/7L1t9
rAICK3caYnCk/enJm0imlgEEWMH865cvuZt7x6uTyAKLPz79NvkYT3G3zp1SyCpl
QIWgYLxL/OgDw6kTTM9a/nH7KDVGB4GrBxcJw7LfTjUOMDypfxAGCPLgpcMQk3lY
L0MLyGHEyMTJ6a1i8wQT/2YVG4OibHA8WwE9pjJSkzq5j6uFgyVR+9vqNyv8j+vr
loTvXd8p9ukT70ae0dxc+lLIqt46rx8EvfpxTob5MaZwSbWgHDvMqVJDf01geCcg
1szhHaeCH7KU2xuRYMh+mvbe9PFbK/MQNcWqpobUQaFrwxzbAC+EgcY55ER5jHEx
g31BAb6RbFkRxmJBvIqJjEvqz3IURUvGa0fnuwanNjFeGgFhOA6Kv96B5lt0r7k2
poCLfA2w82HlnqrRMnTC5fo8D7VRYBZ4r1Yjm5fW12KvoQubCGTz8yZ/8yX2LnXR
jE9Ukn2LdjnTZncmqwOJYrRMH+Jw/FQo5D3xEv9egoJTCBQfK5fj/GjKHN+83Uhz
oTQ23gBCdQMXKee2tZi138RwR7ygcSwYzKNxow1Q+6XavgYDOm+kg1it8aFtPgFr
zFYjxrHoQgEmdj+Iz/YyT+G3nSeKYpSWyzOyb4+wYX+OT6WPPFXQ2dywdInAK2ep
XZdwE83puKpggUQFzV/gWG9i2vdtF2HiKHEwEdnLEE7P1HSSgBKAKxxz2uGOzDju
FgWMzbc0lnFPLzF45edGPoVL2nxcQRdhfAHddwlajrXYdIgzQS4uz4158Md8y/FB
D3qOxk2oIBdH/2RaY4Ilf8vzY3wselBLGFvewB5Y2qKRlOW0cXMQO/9GnnBBJIDA
5JDKcxCGJdCeYkfukOzTE1XKek8K4tBVu2rIitU2jMDxa7PlyG97dvBCwoF0w3wv
EahawgQGbOQo6pw4aQfohRZP7P6UMvTq2uBpfgDXONGWi25rhpfkmKTLxuhaMPrM
eFv8k4MRMFiN8t2SdstkVsyoXeyCU7q6s8jd7Hz1gY1JXfugI++UM5RM5XK38Utu
NAExUQbECn4VykZEHG+YD/RclJbtS1c6BddyrMti7orG0nvF4dK/oHHJVBKUFRWi
DM8b1zo3xa/9iTgVSvQvuqiXVAe1TU2AAIfVA/PyL5KpRIn7+CKwIamb0gvgYKh0
e8iTJTfMa9cRCpGLWD5sTW2qXxBRFHgiGshNrq9WRXESYe6SBxDUONXeJQyt8tI3
OgV+ada8zCPy63aOZGUHXF2RLPZToyiZduS/ey779Z3lNCA0JA5R9UbU0ENkmFq7
5+bA9WWu3ZVg87totgG/NiEtatvaqLJUqbjSInmLZbAVmga3HO/leaBBBrVjjmuv
zXAeJhYFG+xGAdOHNVKhiPpu8tZj3PyJFL5e5Lgm43Nm6JBNV3M6kXLGCOdGnsuY
T3D1da/GcSRhbHcU9Idgpn2zH5TrRzzg6piQh/h+KfLkMgUjjVoDhGleleTfp8De
CjvUB+mWPQRRhPkG4uwxoabvNfgVGLRWurm1w4vlr3qW5+AosD/mGrus6TChsof+
8hEwRUYMlES4X8UO8TlUIkP5tdAjS3RDHLtkLyQGTaNwyaM5xqWl6JoAqGCFbmth
yt70dI7onHF1XpFLFj5b+1gwKRt/XL3ZOcDvK+lnBS8umA+q3nTgBzDbS72qDwrC
DaIL+Q0kx9NVw4zlsD6QKCRU/Hk4LHpeJe8wa6CYFHGV0TCc6F428/BXUqHK+iLY
itmu3rsXfpzPfPix7M5a56E7Cfy9W+3fP342iho4Fe5smz/OZlIxRG9zF5mKyrCn
D1oVq8bjNdcjHmTHGiaLSKDzmQ1Wh2HnCvG1Y5AWLzgJmfdCotQIF5Rz/eVlSbrl
ntihZfeymcHcMEd5nnEaNvLgzfPGdpenoDLkQBCVUbRNtke72lAbPT2CDfLL1rqa
QirZpQlhleg54VGnqzE5PqctUzMVHRfnvuQ+aF5BPnrdYPvOKA+sHfzmJH683Uk0
JT24GghI9bFC38WWGPRycA==
`protect END_PROTECTED
