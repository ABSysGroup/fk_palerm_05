`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y3byqxcw7gBS3oX9CfbIK4Izn6Ix/fzigI2BKJ0tMgoRD48ROOjnYoNJX/zMMIo3
qgxethb4z5KjQdArGGur3JeZ2Vk4etHWGJ6AcwmzLgjK0ThN/ypqKporgmHA6sYo
GO1nQexI257OVdn9iFLbVkHgg6/IufUtDgCIwXzSZNCGMdY5GYwYCP+5SfdIev5Y
2hXc0RRz63WIVfBFFBInWMTSJL81RZfYe8g+VHrTr6POWz3s5W6JmCTej4jN3BYr
QWT/Ue7lbcyCA0lzpZeglBa3IkMa+xYX45hIeLmI2950WMrNF+Y6nl+wDESp2VwH
ZgpG9+uAy4OK5FM6FPVrrQl4anhzFH0R5qZ3BU+SyDoFv60+PQq4eerE/0lMDRcK
y38NlS7pPjizUTCw5kFikwdDboFIxd6TUz5zVYLHbUZ2x6Kqcw7j76XAH+v7Aaad
cOQRmuMf1WKtgYDou2PMkIovpVdhV4R9yhAGdJKLblliEGIXkDswR+K/NktWmYpN
btcy+X/QdIkTYT9LqtP+gW2jczIGUw0fWcfj0Xz2hjvjC6etdawuT+bVeq29nmg8
wY7DJc0BL+btHu/Fn3DpPVhp7bJjvx3JCUNLpjVgeVz4VLZuZqjqEorMkXSE1iUj
/mZ20bX6sIArIwLyAAyrdmGNMcZ7UpP45KMGLV81mguTaD0kdF00IcpWnNx3yh88
GNKwzWODMz78oxidK5qsD5xIrc1zN/u1rpegjIpdh0BU8rFPONyVuNjvhrG5I9tT
ND0jsybDf+CsvMtOaVX0nVvisDwnnxADJi6WLHu9zTGYJ9qs/xfCEm8TZlHFeham
JD62bGsoj5f/6/jfNLGV+qQXJs5MOTcc8nrSShXWzi4=
`protect END_PROTECTED
