`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B/+RqUApHHxYPU5w18sCH+rwUWHOmtDjEsozViDmmrNwZXlfFXi30CvqxgIHKX6S
mnARpPX3Fb0oKA4hebYTNe7CQ5p0celKaTCbKdl+zwVzAERu9v3yvYNU2n8JiLHo
lYGrriq7k8iNB/n8nruFXh6rpB1jlnhhS3/W5n1iRKLvUOT4ny/H97716ynRNtPd
kRsAMrnKWRlOnXb+rVBtXZjIJZp39Ys+75gOzIz5SN4unbDQfwk9Yg7sH4En42U3
NqNvNJkQOsIr4eL5BytWhTWrADNORIZ2l0xxW8fZyQLlDwU/IHe26WDFz+PnIEAD
JyR3DGMXiVtEowv4wcGSZCDwxcOHihq/Ys09tCp4elRZn4/3IAvwoidl+ThZiVaG
i1EmbZFOpk93A5MMxMaVPhjoBTQ6JZwVE91RtC3vbMw4MXqKBBAqsvVh0pflfEm4
NyoaFpyci5Zy4WH8X/+3BKOACAKn8iPQ2RsVPUfwGwtqRWT9Q9ZSHqPB2M3GAzLv
Ech7ET0qxDSGNYqiN0c/ObriUaOe1KgbOYdtSa90jv4dZ7Uqt3/l9rY6U1Wyr5CP
atfHHgSJgCf2bvSanzau/sDjB9eFfWsYKoeuF0gRkBFmmSlfX2NQ4BO4vNLgxeIG
sSkeO1kvnvx07KWWYIVVl9k6/pwyFVDkLjsMz5eMta13kRFtbMHrpVPomD4cLjK+
asg0THqT6hXXQK/4Ourimyr7f1020cVqG5Ncznyl+QRQpx8SOnE6TKqQE3GJmSL/
EJnrzzY99Dzhzd3RiYreD8sMyRB5N/SWkLoPWdFsjvu/yB6bNT9zC2KXqVNcIdy5
Nzavw+43czlwn8qqYWvZ88owBJ+inufqP+GPfuZlT3NQgY1FoH7O+wqNzwWT5h6O
t+XM+EfthCbxQCD5idG9rDXZ22XDO90d9wD2JzBB6yTWxMveN53Tpdp0haac6kiN
unE27GHF5WMstCn0dpHsefSY/Ias44Q7UXBFxmM5zDctl1s4Z/kraU7AUwg8dA9P
HgGi/OBfT+V3dFQoi8DUOesKdM+kKsAvS8w4iwqQqJ76MxWC7sne/YuZWH71UZQ4
El1GiX+YzogpBKwD4n9B8dwReiiJ9J08W8lcyYH3WK+sMMgTEiilvaZ4zStslYf/
l4u/wnvg6/a99l8AHSJNnB96ZbYyzjxzLf4ai6r2C0eYqzsYCnzyJ6V+aLaqB9+I
9k/vX5IfvtnVY3p6iF2d80OZZ8Hj39lMCRRmNh71q/FiQyR0cnLBGjoKfAyLWa1F
NoBDuywakdOt6p8RiYi/4UkfMZC1L70ReG4fwUIwCQRznrem3F+Mx2Fdw1Tem7oM
+mdHFqRwUh9jOyFiJhD1iCwHdW0yvWVSYwjPxbE4UT75ny4sILXbyDX53IFdtDTl
nVJU/rWC7vqXHOXQlp1kYjnf0X5mN0SIv5f/+RR6yhYJUjMlxsMQPPZhBjD7N3Xw
bC5AYN/i//Z83kVWC8tlHmAW5vcgIEE0J+V2n2J2UaR6csO7UFegd14tnnp4RahT
6dr5G0X1koXmgjob1575k3zpBsZtR3tsW2N/C936FykR+WEVSnNc+8acglSL1mXk
8Cy2z70LCJlzIhp9VdySz+OqIonT4zdMVZJKhWck6ku4UVdU9iK0TSEKbuFKZCuV
luYICUZPqTz3cIm/bt4dzXaUy7bwQZQeizuQUJTEV68iwvdDQjZG9YlpQFOaM8hU
dEniW8TyYLuMB0a0sFyBACCCJD6eGrpJwpOuBoBi04iSz8FuTq86Y16AXRQHpaH3
HvqYz+XxXajvsTjfijRjjE4pSFDS6FYRGcu9U4e6DTxT6c9ukfNAMXcG8GSNmaV1
6T+ZbBY8BqCRIDGi0LTa4msE4+ez2oqQUrxl7FqWS/l+dpdkhHoyW+Fm3+L8ruFe
I/YBpOHsfH34acp+b3IPUVFAUBTVNCmzZ8DqnPfBaPS5HvVeLyVW7VwlkIKowEah
8iJdI3rLzYp56St6Qp+0R23pnvLmXBYBgPeAKnIaakoD5EWX+KsNtYZogtg+82h4
FzYHQjK59nLBBhwp+aKhhg+SG3PIMoEaKcYTjEzWmWJsHZoaJWSGa17/OVk/dIka
cxsvRaPkYUBilD+tusZ9NYK5mJ/t7wjcC6ZJ1dQyGhN6utM1jpgvA5dLE4kQe21R
3F8oEXLPB6HH8DeCVmjsNeI3Fq/BrLOIxpoMqKqioKBp05oKRBYSyFU1jfIrCQG/
md3X6RowYHZS/N8MmFg4dCP8Nstubxe2FVr+KP5WGoYntq8V3JWg5bkUCgR6I9Hu
2gSbM3Z0h+xYY6UsA/tsYLgs+achP+YqidAEWlIJkOkgvSPAvxb16DXbQfHFhg7Z
AbpFmJ4x20eZ/HSjjOJlyPDDglKnPcQFfR8KJPrw+OVzUWr/eOS1eq8Yc+boUG+K
YdeKuPTqklue/fuV2rPgjht8GyG7iF8fc4Hc++ajQhatoaRt4ZylVN+z4Noy1Dz4
PjO/CS4KsZmAQIu7EUli86FdXX1l7r9fwURDGWyQO1I+h09Ct+E2UW2ckZY98CZ8
NZBd5EYZTd0+MbP0+faRXAejdTIF3+lUC8O1B4xNpxgDzTXsFbfmORhXYLnD5EF4
JpgHDoO/VA2cTXM/OMkLcAsXxieH/+bRGAcZjL5vC3hhFDUm65vzpTiTAhcbf72l
SSSzwAJKrBT9Yth8UdOjXRDybWTgYx96fWYn3amehh/skHtl821hfLTp2osAw6/o
//gfwnL6UMgDYHNVHCUIKRlctYQzP15ZMfd00ectPOKTIZDFzjiRqfrAceiwbNQy
cHmrQLzN7obrpnxjRD75br4rNulahfwp4qpwr8Z4mMylypykhx06LoxL+3eg2G1G
da3k6zAsNtmNMvIyJ73q+ZYI3FzdgOebDeASsn77QkBS5fXyf4Y7hbHzBfAFimIW
IMszyaR6x1mVlwzNccHzwCoGQ+ZKBhz2X1QLGFhY0QxzaT4Beic2JJ+c/rl2Vv0x
gDYS+FfAsRdXjOgba6139s5RzqDIpP2NVOhthfmQPvafh+avOV3bjALvn44Bg3EO
rWM5yIosY06cY7+qKdsEExlXABy/QoghMyH69mOgNy35YZ4p8lN1t6jdFx/Ly4gz
d3s55SRBfHp8jUCpwf27QUC4FUEnYw8/p55c77Ym0yfK1ojfX/CSjJHuPoaNX5cA
hXWRHQXHlhrwIVXd74+U3mtql8IuxaYwEi5Y61s8vAn1AtO08g3ma07JBVe2v3rV
/lxxStf0deZ85M3ZX+pl/jinmrdbCO5pC4kRGKWUD+DdPPJZ38WTUdhdSC14CGUG
X8gdsKQv0arMPlfCnBKzVATfXGdRsppiV6XcCTAywFtuUJ0yHKMahkKziYRoeAC0
an3/wxS9Qd07JjSbd3kf5e23z5jBNRYOPl9Ag0WY7ooNRZCQ6hYxkc1ZvyvNyIHU
YmCwzSq5SqwPEEQ0zZmGJ6Hl5EIEpSUyPYfn3DW6gBI1xqcaMtuC/VtMxoGzESPO
nWBhggQajF82vFvVu9RBagii6mOo10PENaVf6yq7au/Ugn+mqISrcYW3X3m312VS
qGXH5H4tpDSTazgqIZcY6yDHPUO15bUcY8dHdkojDjyjDyQz3fCjGyj6tnuj34jY
LSyPsQ+hFlAvKB6gZr9l459kmcINeib0w/pVhOeNqyMAbHh/bKcbBtBaI0ZmpLsf
veErcqVOO3ZnlyN6G59bxRaU+jdWn/0wRyLPjtZaNXOR5IWmV3XBxB2K6Sddw883
OYiSWnYpnWabW5qbM3RURFmw5YhnM58x+fCh9RzLVwxTauDYWfiwE7oXUwNcK/JM
DEr2LFQCui0QPSzqV7RgIsa5zcWfWjUuQLufYS53YRJZI4NnycCb0TRgGcdOKrnB
hB+B+yD+m52GAcRKASn2rXKlhl5pUI2X9mzwvORqqjoPtTVRWwLJWPMCiapu+AM9
DNx334t3R9qJP+a8OIToY7vqiNbq6TaKp95YOjTzfUBBZNBQOQYRKalBlEOUjMzb
gbdaTdl6u/wS8fmVbD8GloAk3AMNKiVNnnsl+1GLgTLFBgJLbMI3kYNyUm8QC+DE
7nslGhodWHzRdhKwtRe+n/TXEbWH8gpDnr/PcEM5CjYuM2Pzv7Mu62J1XFRi1DCE
lBLS8ie7fwprVMUYFTsg7CfTjvC245BZR/rOQWDAaHTEkz2ucCcM1AELaj52FbRF
x/0XbI4VQO0x4hOvliRctgA8Y8lpWiKoKpFdL0RGIGGacwTsR08cpUGQqVeVO/JQ
nMRf+UQ5JRnxn3ND/2YSPqlsHaVl+Ljw3rSma0CSnBnZdSk3hlNtl5xc+Ireyd/I
7+OwSHW3Rk7Sz8IBd0uXctaCDNGbE2c+hYjYdoiCHIvSGwLRqadI0n9vyokIvLyH
/rs3Ix/bYXfrrZUtp3Cjpg1N2v7hU+EaiThvwHSqkM+TXnqK+2HCB051Shv6q9Z/
FvH9jcYBBvMdHCnFcRP3tiR+lipxnCpzfxzx+hNqXCbXR8n3W/kxLgRvTczwGopu
6SG/hJk89edWeNZxoJsdgDwzqFqHdZ9prR8xf1vyFdh0iMl4mokzoiABPlB7u4On
mRg8s/kYg5lO/kFAhieboOeoynVFFTYTi/K5kjqsoBBOSVB95IXX3Qvdss2vBJRE
oSJf1Qt/az+33mkzmO5RgD7f9IhwHoVQw4L+9mNfIKxTX8WWrhX1OxFQbKeMxPEH
X3m25Yjcl0ee+MdD6sweF7SIKcnDltBKs2YQEGPuNy6zs5XLgyBX9rvJ3PJPI/34
6a1iCJuqZNMSFF5MavCXs3pIPJsuxQqtP/62qn679THeEtZThOgyvZx0UiuHDkfv
i5dmF43K8n0O8crOOD07WRri/LP9xJ9MTmvuVoxCtPJ3pW8kejaleR7R2Flh6Kkd
o2rvl7CB3RZKlwKnydkK5zXZ21XCN0EiAYvso57vofG56Nfnz4oq980/KYgKAB8d
l4Ijdd/xMHMkESbdXtFwfN2r7LZ7pl1Eypi8F3gu3sk880luH9hGl1Slf4J1fdhH
nlZ9nRzdCleDEepOKN0FZPIyMcCVX8pA1i0InSrI3m0nNuqnNWWexkU0NR+zblJB
VYVs8e9R/vISQLfBVlHg0Lmw9LNLsozOEqupDdDAoS7HBR2lyVikvgh90TntOqsb
k4GC8V8V5p/0FtdksN+8gy2NIo+7C8JUqSbGQKqwzxOUQafJFq46bLpdjqLT1Eae
bj4rLCVJlrcHmi1P5632krs5DCx686+0xoO6DCXNMVOSXxXfk7hVgzXLjmW/DpyM
nDMxKWaOy456HdK2T7zikmdItR3m2dDqIYlbFQxxI4Xku2wH/9DlL9Dbqu3JC7ab
fG3Rk8SWTTB1x5ZVQhlO4yK2m7vTsE4XJZj+CvCdimE6WH95AY+L8HuWxG5+SSR7
viDNB4w5PDn2fSpzFlhriGFc5wdTLXw07UuD1ewLvlsMNNzEIiH8bR9hsPRsepuz
KY8/oJBxZPY5ycHP13b4sjAJWZFh+Gx3aGNCyvTV+IpZyEZ9PHCn6t6JGGPvpCjY
OR7JVE3gIPt3ChZKhI2sOYkRx0ffTMCgvLRmdXfW2kBdPxLowa4hprHHA6IMGzlX
mvYeEc0HTTh2tG0AygFv/0P+Uni0PaD6HxWH1yH0r3nsMAsfBS4vXcvnBp8Mw8+2
UZx2H9xiObcjtKd1QKQaue2TXkrjDJxSVsBupV2E4ymrRI3FvuDstPSOGNT7AGcK
eNg+u9nCURleEEdprJmLEwXChXSMQ7YNBjAwc1So1ZIje3gwFZ1Eg+EJKOhA9PHJ
uROl/49t4xlFvYc1eILyDpdr+J5aIn7gGOMTm4BxK8lPwvGncvVNqEOLih+DrA7E
QKQ51NOF3mwjWXPOrkjnceIwqcOynPSi0DdC0jTx8NSXviYtm4IdyeoWhcSUjqrA
TPtBpXLN1wZsnpFmOCgGimbkDv2tq4RtHfLg4mVGcAoVGQhIY1a2xyWgabUArNku
IxDz/jIPLoxCNITRJV2qHzFTwI2Z7SQBzaSkDOOLx7Wee2oTHZt+LyL04sjWKKn6
F/rK/9iFyhZFidImrpv8/wDWUk1vxOEIjk9A2OfexwSFAZgxKJfgvnSf8nyDtHLP
a91u0A8YPeJNU3LgPlmsVKj6RisghtMPizVKdkVnkTYTimb93uzuLj7VCoSfTC8o
4iXYRJeF4ZU/EiricPz4XSzzC5YL03FCgkTY35DTXk91/pT9h0jSu/f9sdKW2sjw
JRsT2pc2PJTdT+4hL9HIuJPPtgNEqTlDfAUTEnbD2d5koNEoR/gqGOtKzI5vURYw
il2n6viqHoIXaWAgorn9+7Nc2+pJUMnuHPXOY2R22eBAAk/ZAo1XQVF/54s4xRnN
mfO3QdLEP4LxNh7CkWEoNcUHMoI010M64EPZ//Z30R79NkNIYIWR9SZKpHg6qxjk
imDh8cJALmiAvu9GYlzdXR3I8lOYW9rgfY6nT49bN0u2A2BRcY2Ggc8vrpCjEnTg
x9lAt90QaApqdypzA1oAqNepXJwaqimqwQfbRvVGYbhV0KkY7MaMOnreaGb4AGet
mLNDi9BWW45GWr93gnETlrFAarchYKrWnE4C+0oARdAPgA8/kez3074bwYDipOwB
pPFrJiU0EJr7ExzH+ha25+lgbDnPbkCMgJbOSTxh5BAPEEeshhfV8tZD2bH3msfu
e0Wdd1DOXRcqS0g9Sup3fmsL+/D8nuk5IPpSzKBblcQYG0xDMt2qjtljPrgjRa1U
21FJUv78TKT1xhQoin8lwLK3QdyNiJQ4epSahy0kQF7iKuY0V9TQIaJwOBC533J4
OzemgJA6/70Exqqe9E3hlwhStZCWbMxu71UkiKleti0NOKoSpE8DhucMZRFzW8OR
N1QQn0w4QGmOdBDDrooxIsoZlNV6Z/xHRzJ2r1N4qWbXOlcTeVMwejpUv7eQQuK+
eQoO37RF5nQMPC54WaCIY5ZqkBNckrXj7NcE/s8xmKnKPFrPw3LKH8jNmP/W7OLW
UqaAU00uq6VySPvcSKhCXeRYzQwrIQ8yDFwCEJO6L4aYyvQfgCpNNY2T4lpfsTdU
9rHPWufRNx87h6mqWscrOg1TDYeHAKGbCsXEq3efoLuvXSmBQjeKSeCVPmmk/QlJ
1kraw2uCTLG6I3wX1xj3yLNwl1tkdj8LLXDqgEs+vOKSvNf7s8dsIRSHMnihZ4Zr
/BE9IGTf+YgMOXUnEkdVYiPqVAKeqlwv0KytPD4h39bNQK8Iszsf0F5hTbdJiFuq
V7MYe/wRKtJebZlRHcDyt0RC5j3jYvj2lPT4S2uUDwZkH5gYm95BZUtRAxWA40m+
C3/dKPHKSuwJs37E8OdH6E0NTMOsWONIpnqEcpbv8ZOXP5UKKXfypPPKAYxcFl0g
Ro9Kv5G57o2AFSe+2jf4HtSo3nQnF1hQNZ90Dmnf7V8B8uHAjpN/T8lnO5Ofh7tI
9WH2riYU8Wp9ij7bT2Pu8pDX/WeOOwuMPJLLwLyeusKKdW9xiKZ6IuyG9RNe8H6d
4YkG2E73yw6vVj40+CBAhMC6sIS2JQYo0zA708oOOFDUtbKOB7mynGTD/pyzYbrC
Xerr7foYD5eNhZLkPlJS8TsojU/QwmYnVpRGEIHhTQLsRbhYHtaBFYSPp4syQlMk
8hOC6xG+zxEpmKjKVT0NdaM5+vCTC+7vFfaThyZfaeIOeY/ZkvyfCIrgXKVgiTPX
W1U4wxedi8SOExM7kLlkKwapjNjspsb/H5Cex2kR2b0pwrE2NKQDikxniiz+d+BM
UGh5WQowfw63QCz/0iEi0JzDzYpwOOKQ10JpD7I47jZtLXp9X10gnhQSAqPTgg5P
O9RKGXOvnWYQtzMItRTIvenW7wN3+FVCUvjAqiyE6ZcSHXKyI/zM9bnGe3lsZgAp
lLPPpdbfAFeuJT3FSutgl5MM6iF73GnPIlWA5RGPzRSoHozmRTzC7kOi9aj616CY
kMc7R+6gaPUcE6VNbyedl/XgLD1PiQDGLQjmtdMjudbEdRlJ/Ke4Wjzb+MLLOv+h
ZcX7OOmzQWuGcAfzSTrnkML7b4WO+4m3fSm+RRzqgvZfclq8D+Lw1fpjJY06v/U5
aaWl/apegSpErH2hOv+zXCl+RKwvx3WF2DKoAP/vSelNXQnY7Ea8RdfVZKtK9KHK
wFJNNTwBI7odGx08MlREy229DQnq96qkEpthWc9xa2jyzyizrz3NRurUb4MN9YIZ
XaanVamESjL9xcvivdIazkfgJmapRdaNmoROWgxdcyRGDDl5SINrcUe2A3oKfaOy
QEdINvWKMZt/oXRwipS2OAwSbfgdFJ2G4adt/Ojje98O5C7Gw4xWkoVTKPL0UfYd
NnJ30+bssVJUo8qBU/P8IQN0tSMJkyWvXt0ibR7xxXgRr91zbkSn2u9OFSHBrBaC
C7bhb+8oo5re19qPO0iucROG4jmDLLK4kY7lMvjVdaT4NMal2Xz8bNwjhXTcRJjG
3+UOmcc9m48wIxjC5BzIgeaYjgZq4C7Og4MWMfxjdHSbXLaplKmsh+Jjou8rKSeh
ivUSUnhf2YYzROle5RpohN9BqNH18Xq0ZvBip3InEzodmmLdQApweTFyHXbh94gP
H01US8oPAuWwDcbtRY7ez8ZOncH2Y3sVX4ftxXijZBXJQveYoA+4bAbQV7yMO87j
F7v406D9KFT2S/ul3Jxj/0In22rgPIZtEdIlKmRZznOsznqKDrcDOyEkkMzJmdaA
2v6xYZKV2yPJdALTb/VBQgyHNzNq1++tNeDXsRNMtKTl/D+17Uev4ZrW1MZK0k1L
KlO1XD/IkzaUaGbrtBpmfwz8fQ9ArypMgCfOPGXzDumcR4S9t3nFQ1/ypUPl8gsW
iSwRJdTlhsELYkc4sm8lqTpCumv18CulLyMvS6zZxVzIjR6Ul6DAkzbNTSzwDBt7
1DKxlhE6Zp9Ob49affkX77caqpGlBGEV1kU9J4Vqy/IpV3OrPazyeAcFZFClP0Ur
CzZ7YYZGbdiMbVtZSS1PFmk8QCxyKUPR900OTQifnIhvymvDmYBV5kKMjERS2hPB
/kdzxnubpn0Zun54mNnbbjDvtJAlkiB46w+JvpvrsVoAZt6aeJDqvzqXqaWCt76v
1izJ/TxO9aYw+iw8OhN7Fmo7PlcKE5ZFPPWccG/sMnh74WN75sROVbVZBWt148h5
4rNsFAdtWoHQl72EgXps9V0w1htfXuaDrM0chh6MRC8rcf6B+kh7DJdHXTGxpYB6
A2Grkne+WeggeY1ZSXB618EPnzuoQGqvtwzvECWzxPtwx6JLuRQXlKQSsj/HBV/s
GbqqRoc5iviGgjdG6BvBKzGrxJlW3PAeQMDluqlZLgJz/DHDDPdJtHzYb028+q/j
FEvrvznQ+AoGtFfH9p9OgLLFjxwGSHRBeOcwySNT8KUnKfMc3gh2MiFISELVtREz
BBxII1GJo19JYTQiYdXu5Qehsro+J366UlwtoUWDyJZKbBQfeDWo4NUN/74NrQhx
1X5U3EzoWzEH5+Oz1Gc5YAVOiT++uEhIo8c6bw3C3o5jupW+Drpk4cxdJQrGS1aY
OoDRILwuE2fOhfazIN3JS01Oy1PNVMjAJmjQUIw8fAzunUFTl/HGcdht45nQeRcZ
a1q4E8uyq9WM1cjMiqqIwZGW+Hb0N76aPtLfGaKFhK8pKETwZljhJFQ7l58zAuek
dnCApJMe+PMq2oTxxHJnsPUJu7mcnLrKj+6hwOAOKyNeAR4ozg3g6y8r0b0rectu
7pagzYc727H3Q+K9Rptp1g1M7kwA2cf8+/EIBLLA2ORcCWD2x/cCdlYj1Cp7Z17u
UDRFQBzQFldu6Wa1xaBXRsw3S99JGYp2RQhboIxP14toJtfAc+C0n9Qri2aqFpzH
cx2QFXb3n7qCrv/edBxG+AmcMip9699o41vjMB2nnQqKBTnCoBWl9KGkgzgoPbXd
HEjOGoQYetSpFsCO+NVMWrU9xradKbLlgdYtAr8ztAjRJ2E1iChXWRJork9DwIyI
hX9Zohu2XNyp+zLXSX5fFnIPeLw+5bAsWt2UXW1EM1xSNgpOJSE1YqyQl1gL1Nau
ujtOqRhzYwe4M8gi1fRvppgQsQryHPdbDJYzhhhwxqbVMq4Y5FBWvH2Cht5W47EZ
1t+5qOcy8r7VxoTpeDySiEQvuksCKbbqOagGGMZw18orhhEHOxszw1x5okwLCsoi
MmwweOqOhef+iebyBeAauqgfY2+fTTb4cawLwgmeGo/0F918Ye6YCzQqnfyK65+H
f7Gx/illk6WW2zWXYkhy7DVAMOSc36MFc8PFBrxRQ6BDJQFJeRzikZdSUMdEmuwi
82GpryECjhaiqe/B0r34pVXk0EtP28VzRXcNrjIMGuLPOfjDEfTal7j1e34HXPPs
m4Do3saLneIkxLReIHrUEdEXmIe+m6ftdBCoX72UbhOxbITcRVjbPD7Ta20to5Im
oU/cpWLpzwTQ8Etfzmnl0aiuidzdL2lYb+DapSXPlHWjkmSW/ao+miulI1AYw/CO
wo+xboLfY1HTvnRnF1HVX9eYe8IsiJo0z8qfxnCqqrV9dblgZmJs+mYshSe0ENXJ
c/0jEgYQLFdk87vF/FjfGkiaJjmPZElnx/gunVCdRq42ZJJbUlV0OQLQhFLG6SZt
pwwJp1fCzuWYceRDorP2Rtn2aEYCsXpwufeOH0Xh2UaE/m5yWjUskxFzHiOtJz3d
ERMAxdtQAo5No1G7UeBcYXrJa2ztFu5RsC4Yl1XcIR71+NV47JugDgzRRBw/ym/v
PIbjK/+y45qysfh85z4FLw+xjIYMCBwSOLLplzBrxVbDTfgaqwqkeGVa8Irz2VWw
4TYQB46HW96GaOCCnupdnm+S4MO9kVQTbb7/7oVXKvo47tf4IEGTHJPt9SdI9aW/
i0g2U9swx0F+75Y1dGG89uYlOciGAgjgooBzBeGOhj1/4p7IDjQc6v+svKb4HQPv
cQ+650yn8MNRqCpCCKGidpy/oTczb4ZsKITRxLWik52MxNhGGJ0sRRmsZMldT46z
Tec+AJEIOqqSxgM2HynC8kfAS1tiuzav8cd0O6UgX+ivKr555MAaVEuTe+guYqEH
679gxEwuAdwbHGovISmF8lZ6daeS4KSeEa+rwWQSdf3mfiMtUTucaxbxQ3vKXuSA
U7e5JVYs4z8IaMhWVrnJwOLb5JdN23ucTZ5GtxK6/1STK2oCIY9YpHYiILe+q6jb
G0mhl+0h2OXIstzVejUfET9Pa3BksaamfYyKieHgraqFUrfo2891hE6XUBOtGdMN
Vl8s7vKKV0Kcy1N6Q1yZNewT1T0p02TdIihWmyKnk2PculCBFI2w9o660iHBI1qz
jM+IyqJlf5Agf3xNYbwzBzOmUEZYYXozJNDh+A0M/krKhmtx3crl1f+vaKwuOqKm
7g7TJ082cpt5SGeQ7Q6whMYuwnddQza3AXmg+BKUtwOPTofMbK/OlVAJq+j07sHF
DNl/hh6kZgxXZ7TuIuUCNw8BpDg0UCoKLYfMx9OVxZQk3gGEOQlF5vlF7lK9pT2x
HodpKNukQ6lN1o3ZtSl0X249uShA/MwprvTykFLRpOM0HVnyReSFBrG8YaQd75dT
JB41uJceE4K0TsQoAZINU3JAkxGMi5f6Aw4XrbodBRcdl7WSzuvxG9zBIEA0jRXa
8RtjRJTHVS3B6MT/n4PzbzJ8fg+8xseaqACtv7BFdGeIZAsUjkUKH3zKOGM8QLsZ
5Jmh5h5jjN+8oCay4kJOjfZAHqvkQjTG+vl5JfSxd8irJYvsAWPez9ieBn9yHoBk
NXRHUtvQY+Lgr+zuKOvbTV3XVlFNff6Zw89gqpx2tGWRuw/5ys5WbC2WnOLHf49P
86S5Gh/iW1s4tfbkq/F1XNh4SmODw+PXpEY33b5p3lSJs4eIsg6CWak4dLsRG2JP
iVp+OZlia/dFmNJ9GinAwjcRBmaKiW0OOX9cBhbZfQcjfG+fCLHq7fs7Y2n4bRp0
K9FJB5QamrG7QufukZOiLIAkygCBSjaSJqAa256aKVxxNeWyU45j0jU+EvzUdcNs
Nq5a6xILaVTVopUxK7WAT6UX1IYOZFs+hvXs6Pha75R3pVIymLQAh59WM32TCLYA
QXOSsZ8viM49egja8F0PrXJqpd/FYhxuXgVCMk+xbRuY47c2JiccMLut4mUCHcSa
wl0716kR+TPEaM0LL3y2NXtOv9AZ5Z0x05sFu2AR4Col4MbD+o4nmmmBGq5GCLhv
o5lLy7Zs2uf5a5KWkrBMYmBihTia6xNXtsMRuHxVxO+46X77N52KLCep/DOkR8Vs
2sg1gzkg7nyyk8mAS9S0ZN2oQ+XWJssj6kFo78+pEeU0JFbeqrFnPD4QCMQahvui
IRjuuCGFojHX4sLOY5LYlEiCZAgmmM8lBANGUWQ380UxjUno1cFBKyECS4xC/Oep
IUVeMe9wIVv0rODfp9HgSGVKWT2TGxso3PcrhHO2Zs/bwS9NT75qSpUiRjVVxgly
T9WKipjZBJeUwxx5M/BCC6THMETAtZHOBkMSLOZQcGaSmySnlvddmmM52kSFM6hW
lJOLPEeVsU8bRlAioJ9KTAIrktWRZXTImRSxxcWV1wDdtyGsfxkHcW/7uprkxtMP
+KONiGM52k0gCnbizVlwFCKQ1W+PvIllY830gkIKGAIgALFzM2DjQ/chs11Zn4Rz
MrRl8phm+laR8BEnGhU0CP0dMW7ZfigRhlqspCx+SKubQihHAINtYmEG9xCdF5pz
onrp2S1A6YJ1cazzWTykHHrrzE2zYmHRDcgYjAK22Kc2AoAh0tg6Zs7BydFL52TU
eaj9hluq0wXgd5oQh40+UZEEctSAKzoeYpyRdkLpzwsqbvV91c7RAnuFeedN7dHU
Lg4i038CEcutti3qMfLZnu7+yvjks4STkoOaa7J/A3wykXbRiYbbV7G7Gjz4Lr4X
ryWW8LfroUfAE4AchgEqmcOzWA4X9iNR9pUbGTD0vv7NnarbGAyxmvo9nRwXpOH1
YPTzMhIZc6ExZfx3yoEJ1KMCi3FT83cnWtXSbh8EGYou7g/Hznqkw/yyfUHfKrv3
olioYib9MMJxDF5rx3wVO16csGwD4bKME9XHJwBn69ED+Kz5NLJiG09635/TUBjL
RQRd76MB6QRv+x5b6CiMb7WTefS/dzeiJUDANbLS5sRWyzRm1UmHQYYHs+kzzjLA
MS8fg0yuvHmMVhEGLocYkYdvaopPAKb8bXFP63cdGrefqaHn0UPrzcW1qYuj30x5
XmxmNVzIZ+FTE4ic8eRqIF5BvJGUUoIwYUATxfyCY1OHhDXk1cEiqfyN1kF4PYS+
VV3s6NpPZ+nEnpcABxfoXBYDqP2ETV0Ws2iyQEcbJUVOvCE5PW+TRSue1arK9t/M
Xr0PHUR1WZk4K6ZoiovpKr2LtOAFxgb+3anIAmM+ew5YN/f4ZyJQeYx+Zod5lAUW
VywYQDZeOZo78JqMfG41nmUO3x83Uqmopd+R8Itw0ewMDccLDKhKd/+fHZ081Sct
5Ox3h9DMYyGS9EoksZZIcJlaOsNSVfBIaEbSSS9CE+ZABvjFZwq+R8Ha8PJbrJ/Z
T16Z4nyKnLl5Ljycs4I9MDvxeoBh4YHJ9qjy5Wbk2ZJtP5x6ijUa0PI3or6chEIO
rZuGy2uQyu91q9bvRf4VI5/rQ3mOQkV6I/S/Nm/IwF8CIK1CQntZrWE1Xl5nf2KT
sd7mexVOuqs1amN/PU+1+wHGMzlFn3TCR7QEkwhCVVl7PclyIrL5DUOcfpm6vYId
RNfcSz9DUn+tYdSMRj4taPRDbhTWTJxnUagMQ+0Qgqm/B9iCYFTDDt6L/C82c3Gr
FUQpzJgXZ+Vti4qXvmV1xWz4E6q7lPmL4n2iT2VaHcIyptIKaouTU/N4XLjxxPRY
QQnzgp1USPk/ONjzZLws7Sg/kOPloZ5efEw7eL5gh4M6NSV585tRqJsMumuiW+zX
aRVjKukuJBX2grILRmIDUx4RBdH0iL20DwMBHvgmME2WpQ/JHNgQUIuVcljYKmdo
JUAh9oOf9dEHF/6CKpv5UN7Ujm++QBEhGvwHXjcZQZK0Jjb9w3VO0cs7wz2fTqXu
59DhT58VpOtYprw5XL7autw3a9Q6IP3mYk7SkpC2qTRjfXk7F2hX/OgW6w73Q87h
dcYtX70TgINE2KqfyWV1mw==
`protect END_PROTECTED
