`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gtiyaJEFUE3vMWlL2mu2gVD4redcHmvpDtySzOHxLQN5NUmF1zTeYF9GytNt81jZ
QBjLmHH2nB6kqbxOzqLLe+ggBpJX78I5gdIxU+622B9fOhNOZ0PNw5hwUIvGSbjY
tgk1eSmYpG5D6pM9aNKEZJKqPD1nFSpPuAO6kt3i41u87oXHvi0SGS/yPVH8OV5c
vOu5KyycYzM++sK5SoxDeWlhsSdwvL2oKtCbw7KQz4wD+mbGG2lneu6lILb08Iqo
FjJAhrB9lOiPcBaTpfkkBno9lQFaccrr0EE7UcEROMzl0Hm4jhJcgulcQoUjjhNP
256Z4hZxQhXN+s11/7zIkQYuIc+e+WdKICvdWXgSu60RYz7XmYSSt9ijTAHlKPbe
xDDYKnzMuF1mxbKnuE9aPk4mOqHY648Vduf7KJDJf96CmWxWlSkxc4o8trLtp7q0
`protect END_PROTECTED
