`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Opcfd7j4Ea0AroscckvesqYZi243F+nHIwsennfgUSKWjnj3jrhfPHYQt6yAkaRT
YrNezEiucIBI7cYOokWkv1Qfa3CTaTq/z/j2/p8gF6nJJQcPC2uOzmuUAx0+H+0s
pqncPMpS+LXErH4j2Gb8wrxNkSZwK5+w/ism0Fqk74ovvBfJH3+lWoc/VgQh9UWY
Uws40F20wEf1NKue7VM8kFcybR1+q1DNYyHNLxzl+5j4ZD2KFKbefLvrW7RwcF8+
Ku6jMT25B4MwpknzNyZXM5dAP4b7uNPN8DQo+gM+Bfzzq88lY0lJDWPNDrD6JD9K
KxKJ8a89hm+lYG7vnubrth2DF9QMx0wX3mYas0OaTCih9hzJDHY4wn6Zi1Fz5COY
PhlScUyuOpARuftpWecx1q6ezX0/7BoplvCHLCM1MGiQaaHJIXebXDTj5AdFFkt6
YI/xSeWf4I3R21PWB8KFXSW2ICL9W3mDIbtxWXD2Xvitu1lkf6bdmltNsHGL6cVO
5Dihdjz0YMXmfNNqzLDKrHEElFotMxx5DQ5T2jVTblc2xN+pAtHxllzON/1iEf+T
NvWJHjjGaNoNLqWKvChLM6hJIGlI3rg9seOULkU9V66rXWUScBjR5XjAGLzTkb3A
48aEXtcVOMOlDO4p6wusCQ==
`protect END_PROTECTED
