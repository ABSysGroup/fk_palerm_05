`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OShuy5YtoyyxeUYPKYec2jNx/9ZxWwNobEtoIVYYWI2o8P2OjoJhClMtfbiHVOIN
ZV+/WSKrbeimj6HvmDmGCRNIBlxITYDCt0mNu4qS7HGiEAtrU8SI4Q3oZZGHn3dW
UYIbpGv3hedcZ6mn24WZYoegZ/e+CzeGTGeacc1Xyg6fZWZMagEPMWInmy00xr6c
t0WN7wxqbFql2Vmm5SjSuo9DIbC+/mJCiIyxRUThAXJgFqMTShOdv6HlPJst7RWT
931Df284xCnDgI/1NfwaEUZ3vkUpf1xWEOv4QtBfaz5wojBPwmFVBoc8H1kHX0hW
X0HaNxlKNPB2ITyroKCCJ3YmjvHp8iagZjjZ8N/yziL6TybzDDlC/QW2u9uNMCDt
qe41wkNMWRMX1L8aDknQQQSSlIEXUmP/XGiwllvAUjfSiPwfkX4cZ6kPOun9h/p7
VYkyTKoKXH7JvI7TT7BEG7JsQhSBBoUWq/tEQip1Jip+yMHYjRfByIGIPjDpCiQA
UwRJ0X2Pt4jqCT83kk5iyBlfMv5/lrE6/azpSQOZvBID988IP480uicphgIWqgUk
jPPcDVCwCLEYADIN1tf3HvfqzIFKYHfECq4BzCSToQXOpZatcX9OWJ8ZIwCwMbeu
Q1+Oan9Ff2iPNBx5rzeAbsCufts6ds2cOFYNKqwwJMVX66IOCo1QIV7xvXR4VoSU
5ZEIAdoanPyZjZ87a95nA4cBrgPi7VMvBiJjnd46O8ZlZk53d88uwiCXe3sT8Y3f
WTxqTiWsbG58VcEi7tga3kD6P1U1nIu0O+npoS7wnvU=
`protect END_PROTECTED
