`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hq3YP3/3t9nnrWnM1KDYn3liPpcjtqVtkiHlW7sCcFfasDgQlSC6DzLUoTLOY/8P
1RVamBfkdm3UsR8FcHPG7+hW+2vYcnKmD5Q/+t4alsHI+8oCIHNo4nGrTm5Ck0N8
vSRW/q0czLCO7pzDgpVzePTBlK8eyRjP28vj+5ZqMwujQVmcc3cldiWVzf1MFACW
28+YUJE22pF7T4nsrvODnYOPNR4MlvdU4LaACChznQwFv8reUCeT/QI/n0phqsoq
RLlcmqtvyo+7WZ78kZER3J9gyokCpwO+jAfzpHyz0JjsxIADGvpWlpNDk/Hn3R7O
Iy8W9LWiBs0gJwmwHefPxaQ7ZvsabWZ3M16UXh6w0TkViX7YABOiIn8nlQOxXXcM
Qfqj6w/+kCWfoBrjeE8fZ04cuZNN0VLouHbCrNvHvmkCqnIzgGIMqyMrzdW3K0SN
ORvMPXeUN3GUMtqTbUfEGE42PHt8PoEp1ubWdGILHjV/tMfxAtlgtVpsLj5cYCSb
vvB48j4m6kKrEqPSql8nSHadZ0cak7WJAyHSMGlah4fDdj93Q1+ofrLyOKK17Ec1
6IlxMPdCyodIzHi30cWSjwG1F2CyE6HnJokgNEIWJrwvaqbRJWgwt200OMvvvIvi
7VFDokzubI8rLTkBNWBa0A==
`protect END_PROTECTED
