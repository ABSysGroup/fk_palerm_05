`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
umC3Gm8GJ4HPueL854KNKaNBsE4C9pxRqmLrQzAP2gut2c+UiQ3UByNDD2oaxS5T
O8lOIc1heB5ynD+fUGDh8FBGFcONcaORgynQHMj2dz8P2GGT9F2Ft03o2lqUqx4S
5Z3XsPxoQucMN1BQtLwrFjSsMu3me0Wa0OKqe3a7Aid/ruPWDPkfciZw2iX+utej
/O0GODN4E5C8sDS2zQP0YWuoEo+VXEYXSqlzojHWfi/xog3zMxINef5Hweq6bV5S
qa7AEShIHqpeiYqEaLTpJM536Q1VaXxI2pEVSpuYmfvC0Kpxn/idv5tU6dmjUhTJ
MCeX6Hk2DrCa8FUGhGXyYEbbHwuqg3NrOH0h/UPuKwka5d+8wzCe4G9x10z8jqjI
nGV34iExWhMbMYE7ky2GlnEQvkq0twGHgcRd3z5CAH8Hz0O0/04jTgiYezQ0sKO/
6P9Ak37VAiv31IWyDBuURMfbDPvcR3znfv9lGAOXq6Qlh0rkdfiMtKvqPzRXhlgP
XwAOl1zoKUE84f42vbHGGmhATKr7Hx+QX8eZ/UwCV36RDiuPNbHbx9+IHW76ry6g
ED3swByzDB1rth8YgvL3lukR8Gw/Btu1wFRKm0UvkjlCvEHKsAonnhexPQWXW3Rm
Kxyf1zO2BNg8y/YnysN4fVE20m4jc+KWtE+jAtjzEVZg2Ad0jlKQX3oF935B20P+
wxlgfTuoQ8CvVysrhggL4rHxr8YGALPQ8Bkr3HpLqhoWmpwlteUWHABOkdAphvfI
izCJtVDtdSi+Pw8nlg1Idg==
`protect END_PROTECTED
