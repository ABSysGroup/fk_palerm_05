`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
drMYTPdUSa9wXVCqK4z6z/MnqBwTU1iwJjlJZKsF/jGjwjvWF9y29eFJxfkCA+Ko
I6BRlsfaH6zCJDmm3TCHnU4Lw8kIV8LZkFxTd/byB1RTsbXd+zY/y2ufy1Ix6NA/
7s25wXyfnhYQBKV6FBS3lKo2LRzzoFHrURzoZEaEZnbDe73en/pLbch4hfxDkPdW
88F9kcGtq0W20a1joPYdL6VnBaS3JfYiVIjmmS0UdOfMAoyiB70GxAm8qlat7qyI
8Fhg63hCYyLw5laOND5iAjBGxbr2EIFmGiiFx/nRq/1uNOqWhqfpa+nHx+ZIF4QD
fQRUywdcI7ZEsDbEL3EUGTi4tMxC94CVE+FtQtr2E3RDrd4A/IkmLHgPqR12uwE0
LinvsNxpy5+Vo/CmzTJwpeJtnSDHeoPLSUDskQVneQ+Yhz5MrXeS0+Ouu0TVDru1
H1LhkA1FRDfV87NpEQ9KHDDkeS1I861NmOci9n3g2nfbUNIHLzdvkTKHZmvbGgep
7do7i/0q7Ekg7jq+0msy41ZA970lHoIYdIK5XAN4IC82DbHwE/mnnPuhr/IqmbJ1
wS9p2QAL1JZL+lu2EUMShq4pMXGGuukomIE6OQjdFN4g99TXWHeJcfrbz2kfcwya
5XbzxVqq+6Ed8Mzp4wo0WNPL0LZQnZo+ZaGlFgyecYfnyQxQwoCU8Orz5UtsT/Xo
i6oieX9WtDCZZGVQERNgmLYqUiI4jortKb8jcX7enjfZZfi10CyqNsqiEFENnUOs
UBpngyWT2ZUDDwI0cdGs1T1kOhKNYPF/NzpY48sPPeHbD3mvyDDgVz+AVQJHm9DA
`protect END_PROTECTED
