`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r/3bw2V1ShFJI/nMgN9wA8X/aSO0StUKlnXWgWO+EwQ3dqtbxv8TpohCeuHYj8p5
e3sseQFJPJiVxB3T1fqN7/fr+s5yKFR0jwA2qWVx/0dGeyFYpAl3I6ViGD4+FLqv
izRwIFOw6xtrTX96qBM4774Y5rTFlsaxpeSq0lMaHRh8lvhHHSSnIIdeVww6nc/C
KTk9rikyqgEbuwbzsDqYH3T/JiQbftgv0IR1bkYxbkGzC5o2KA/EhAbZdIZC0H6c
Awy8fg8IRK7phsbpNUDjoc+xRrg+8JxqM9XLf5V+ekdX7no/zyIHYz9DYfk+F+dK
7ioltmmyVNoMnOPTaS1GYQ==
`protect END_PROTECTED
