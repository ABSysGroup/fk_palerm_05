`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LQYOTT97r+fGyUxHT3IVs24DioTwRAvRNnJS5Hk0HlGZLnWqFIMonjNOuXfLmFWw
1C86V3NyAAvaIlKY7I03AeOyg96CllgQ6kSvHqIPd3nHFKkl49sAEtsVzqy8tei6
VofbppCugjlP4CsOF7AxS/+zC7ULz2JKe7Q1tDrK9AxyFwVDkqC67LQFpHaYlhfM
Pjm0F+FwIkeosw8VWVQ9xt0Py0eRd1xzzgWENoJAPpmIA+NJjA/QeTNKZd7CDs2U
tDW9xpgyyeU2wvpCKZzRggwK4pCO80eajrdvNpXDi3XGWDU+tneJ0PavhhTbLNnw
s7ar5ApUaatuS+AzP5E8YqW+foD1Vy4R73TdX9mdenfeqpDXRiK1SWGWPzdwGBti
6Go1F+RyxYCvVx9o5IhpZoYAUsP3yJJLMPjrY4ndDgaanZpypMmtSUsE+sYx/1YJ
JSiH3RmaDrn+h9teUaUUR5cyxrS1IuHbckCJY2ibYjhGTQOFLbhkiA61uNau+gDN
iMAqsBAWTpfiWVaPuwjDnciWRG/AogujQ07ugovNT7W/J79UCt3vLPm1Mw8TrIk5
yMsB1axmFbiht7/W6jcik20aUefR/zR2thl6nXHx3nneaoJzqRqXQorflKpFf3U+
Cl2YUKyxxPnUykvGTmjXZJygUaf2EQajFF9bwJsvBwVrp+ySJK9I4gR3J9NqDUlK
ys5fTqW1WUzZiNIkqP20soscVxM/jXcPzR/pHWB+QsMZD0SWk+2z9Vx3zSh8fax1
knH/mRZQ1dRJmo5yt0ngIw==
`protect END_PROTECTED
