`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sbE8pn/B0sZ/q5pJ2DsBTkDMkANZUq55KzVNz7KdmrkaK2crmOeL/PsPPPVTovNR
0yyy0Fz84h+stzrKjEqa94AZYgDac64FFHvPNR6xbpCcXFUeEqQlH1HxXlElwT70
0IN6bDdlz6t9HuU3yh0Yp71I9ZjKgijDnpPC6S3mxG1GE1O9aylrRhugMU/f9SY6
kNKnL+Pik8VUsHJtk/554wc2gH97RgOxgad1/BFtOQ3TRPHhwJ2S8S2cW5BHJAjl
YX/ynwqgSCqUmUQCxD/G6tDGWafYQp/cJvY7nMdcAiHni6zaeKMZgFCsT+ttjvjn
HqAVx6o/fsgYJPXwGfBlm0/Ba1uR5Vx50jNxjonCRLbGn4WayfF84mrbYk+gPvvB
jxElhGwgJZkFmyt027Joa6h+W1AmtbrMfy5Gk9oZtKWJivwuhfm8kgj7ugPiZsxA
wGMjJDyPLqEh21UPUnKANiDElA4+zQ0YRZOy2F+YxC9UCJFs/qmUCryT/TA7GA+w
3LUzvhMozN4gMnVCDq4nqHhATfeeM24RTC3qZVhTaSDkwzTvlfinsltrzyJ02Q+J
rOaRFKIpDgxPM4r2CkFfGuzh6Pr7DMybwMxeqfqC5PfOWsuCGjXjFhz9z6kqoCUc
yA4WZ3e7JjZ/zZ7ZU4ZD3uGXZ/jmssG61BtxOPSph7nlzFUHNTll5RI3Nx1FYx4N
Ho3y6bbbQVxjgm0lli4BcqP463xOj1gp05pfMJ/Xvvhn+9ahSMLGaIjQSLcVnVLa
7SpdAgqshK5GdRBCHlZiNj4vYyu160+SXPSvw2cjeOXwmhjHAmIRWoMunxWOwpPn
oEUAW89zI8lN2XjDN3B7QnjvHV7XAhyx6zPFclC6rgxhEjAdFSxtDDRiZ5lXx07Z
dOTqh6Diwz9FQ4PK6AP79ozvOsgJ3+2HayTJseh+cOTrKGT8HT3ZFwZP8oxXpIla
tE1MSrMcT9iImOeCedrcf5NmqDinmWc+WrOe69MV/tCmGijY6iX3m0+RC5cDl0o2
RRN0mHi5zwXaXGgmSfeFbHRR0Y+e4lTgIa/61FQWK+vSvgqKqvU5Vi9GJLIJB9Zo
KP46zyNyN59PVmic9tvoUF5hL0C42yNE2zzl0BEfYBQBfm2dWqtq1Vub7hFSppE/
7pW743V/sHFXGupqYA6zPp+R3aChBHJ7wnH1OqnX7PnGHtTw6FQNUm5Xn9e+dKbK
gfLt25bX7dTk9rwqu3UTzr+S4tFU9rI92b08D/QznhpWaZSAvzvKms2mhODxUD01
nyM4UKvZR2liOeEU5t4IH/ZT0WMt/LDFIWHr/yWci3WLfDVjW4oulcpFMCXkc47O
OXZSH8Lm99w+iCK9ydkcTp2BylYJqTaNscqup+mnja8XgdEVaookNjsisznBDa6M
gOtoY0+wmu5KVanLZ5zTwqK1qRj4HuOiNclzq0p3Yb89hjZiwbB25Q5gXm3G3X0q
JiSxAm1y/1XJ4/JNptWtWioSXYV2evhfoxOwT30HErrv9r+N6rQlFL2S2nJyJ1V8
lqDeBFCZaO+UvhmtHPN17F3h+6AiHjMpzjxoRzFASUF3q2csJ8/cdLLUL4QasAyJ
wZRnPPL0RfvK2T48QHBisGTwDdrr+JoXJbsslxQJcotFAxQjYB63PjKmgknsa12M
D0wNJj7fWowIyCyn2LuqLVf/59ZQCkOX/pmHjnY3Ndzs5gdnm0HiHocJA3cBgSdl
b9Z71wnVgYJHxtlak+Edi9/AYm68RI33dIsKL12zPpBzUMMh6+IyM7S613JNldRD
cUrF33iPgzwNu+yln+NPFJCFGMRMpci44nJsB+n8w5HiYT0pgCOGyeiF3KaOa8wx
3LfzWWraPODzlzMioPvtjnS0O7nMW36KkIddUQAnstmH9jgJcph9dXIdzo1TMg5H
OCyej9319OJcHexunw0/8IJrkgkorRmz7hEM+S2DWBarfjnNGqwQp7Pq1s+T3TXq
/AyIKoBOhvdROiMkNCIGauXttjA4xfRZ8n4X0BTtlnm/k5dlpCjigEiIa2EhK5J7
BSt0eXGHFDhF8Y+SG1Vmk1igu4OGQOnf22zeIFc5mSvNnQUUBxD29jXH0VAa1B47
hANXiNsKZMtlwYYOei2YDhb7KNqcVlZV44lNFJiVrsSqWxIFXohiS63Xiu8d4bqs
w5UvCgn4VC2GMWna4YbgLg+UnbgmOMuiEk5gXakDr5ZvKJNnCegW/JJ5ha1YceVe
XbL7zyULthaDakT4xoaTI/jzKsVb5xV6NgcR2pcHUreU9lwiQML68NBXU8opsUz2
RkmGMKPHs/bA1LXkIdYdPxH2s32+3YVnHZWVcg7IOiwIykP6KG+2pEAlVxdKDgvn
Kf7yngySWWVWUm6UlOlNW6tdVUPIdf5TLyFGLrzPVIJQOmyyYFnVJ0y+XL4R50gJ
4z++zIi555cgfjm7Ae8PYpeO9Uc0aPrZNWMXuRPpJcbjvj1kyz8Fd/FeydrVrSyG
fTczSwtD4eihRMzMaikF+QLV4MA8wqxKs0/km2zPUI7kYgTMxFwbcrXqEfnVw3wn
gyvbEBtreC4lFBpyN7sPHVWVzy7KZL+nX/KvNbU6EFKpQ6NhlUawR7GdCyGlETUP
fffnFo3F5eJ6QzZtjnjuP7wTheofOCOk9sUnPFSVp6LTH39UfRlwkvVPHbgK+4Qt
oDBrm/lXcYrSJ++rAPUSakGEc5CEaq3CQpQGmutVfRI0hBOvSrMtNAtckiHKrkHH
XXKapdQxvBvpgbuNhPwgJrDB+tRzOCNIl826Vr8hsSbWlkw4wrFXPCm8zGAl8ZVW
ZP2iVCKalMk2JqCK+DcJDlPgiyTHvauSss7O6Uezhj49xFmdbBG0dvYAH3wMOn17
LpBby7WkN+rgP0RJv54iCB1dFX7KbS2wYVKRPDF3ik/N7GMWDMT1IcVD+9Ujt3W4
LRW0jj98cf1v47IlVvx9OkvkdyqmCNg9hpZecxqsRrYUgO4bklB6GU1Chd9o9Dm8
J+Pm7AFRjDg2IXgB9B0BkvVE37bbq2pmV+RwtkAkpsE+JfwTBLMutUyggFVBvaNr
XiFwVcwpE2tsnrHvkms0hnuCJVmIWSP8orKbT3pXvn4IL4PzlWfXGjnNOwi24OLc
8nFpaCIZegVx0lLgKyieaaBYpHLIvQ3gTqYvDD6e7OxmoxIGdnFUOUprhrOSwbtT
2kkJmixNnqW7dK6vNBzJAC+L//6jbTBzoVvccTIcpfSMvN8C/N6WE/K64AJkeKny
G4VkTT9sMlpk+JjRvZfgOu+6rqpH5zVJPMziLv2vA+yoeADBHLsNGJjplE7SCdBV
9mQ87RNTD3gPC8H3wsv6YpSlfX+872ELVrEvAFU6x8PpljradLW84ALmiq+A2KOI
icVl0vGSy5wAs+KP4Ncrz8Lb48pzXPiPl8re9dH0BUrR0CyEXRfbPkier82ERRH3
p9APm84/SI0arMnpRwY6lj/ltPnNzRHAYUqJ3ivvH7Y6uawoCOaO90F/egU/syIT
8iBjvKRYKLG9nz+VF/FGeWr4UCG+hzeuOQ1jcQe6dceg6TYfSqzvOTnD3lG52Fcz
rowb31yfMsuY3zCDmnNHUVEheaOgfNBlxdHHube1vpwaV87TS2C/XnSMGltBI1Jh
IkdYkanMsapIKHF9RcYD/GWHbmvPFE9TLpp8/me1Zu5zEZ8PP3C22tkESkBZ57dJ
5FBumEL95GO7O6EC48ef2hjIgFmwd2Uf03FQh0BhWVOftmPS/d6x/0gFCJTElilj
+blSNGNGtiqIZYJM0x7Grmo03a9ZBiYeQFxfwbziZ2QjlFBiJat1n+pDRfPcF/tX
qa8/1da7nmK97OdSQWVBbe4TxRgUPNavQeMVJg4nmwYWnGq6OxPQV9Ckt6Rme5Qa
DIGdKKCPEFlbS79YztFWHVuQCn/MQIUJqDql3AzDityE13wVb5IQUuzPYkPcXAWR
p5Jj67aqFeYC6dJKcvQrCgX7o802U0Kddk+aquGpglj18eCDS4TJEr3h1U2rCe/j
fn1UyuduehUlGPIHEJq9B4dJRLnuwK2ciKt4vGCb0ykNkXKhevZBDR9tk+39bRpi
pm2rCDxPjLgJ0Zto7g3rWLiLFIdinOQdQZzUiH2hq4bkh1OqAqvzJyOfWZjfJ4W5
6XO1iD/cRSMYxBGpRjw2hDPemAFGGCMp5AlHKjsZimjsWL+NStfKrcI0BRkQQBJH
WxkRKkm0Zj44vbvQXaYZen61B8XM4X6vE6mXCXT5T0qFcV95+c+OfNx1UJOznPb8
pvSy/+EqH2zL5gveTk/4r9R8NDuQSaGOdG7n7lPt5uxqhcUKJ33/SkiqRNBlXsF3
xEuWRoeJTsHIaeJuhBmB7wC6eq/JziLH80/e6xz4py89qaLBzXvgBQ9kihVJ6J7e
fzTAN5Zv5dCcYBBvztitL1Lh7MKDUD8GEs0XaOEZXHENh6rcT+cx0EPoTD0kWuad
k5gRSGTJ86qQ7+xFldj0MscB6tes9GQik+RiGMH+ZUt+HaDbv151wXjlCTIDxObM
amULJs00iSwRL8dZjPT2Hlx4xHWgk3syW+bD+oG0zUs2LzU5awPE3kX9jCv8xWzY
uiseRubHAfnBE59WgB/O60+w/Uo2I57M/32yA6tqXRam8Rx6wmLtez1gykMwCJHh
cYcJoSW4L7/7ZqXkpz2Y2xBdIEJo/MD9C99W3CKaTTpg9lLD7Gh+1GvomdH5v7C3
sJHorHkrSY38Tld7hELbWp4NEF3zzUbKaZLtZC8lEuHz9jpeubVdBhFVlF7tfxfu
aWP//gk85Nj/wzzXDBE9zpi/v9DtuaD/Ff2Bu4TtQvr5SKJslBmoI4RN/mn67uon
/oAaShXye9WvL4dNrg669ywjUGZ1zt6dIKjTKGbOvXqtKPPaesNFLEc0FIjDZXu/
OQWfSu2NebL+cs9hyqcluZoDB8KZg2Tby8cKcTgq4okPMDJ9aR34ITHoXVvqg93V
jmX4O3o/e8dUBOFPzABcuGpV04u/MCu2WKLt7nC1VPdHLa/GUbW2l3lAsXpdfSn3
1rfSF+YUpfPSOJG+mUCTncnzkbrO3XhDtwTP7iAwsJopiDrgqUgbuT45CNsZTKuM
1BIjliki31i/6mAUKaYGZ5izdocCMt+1byCZ1CXxc8QzRzjbmeZefMYeCSuYs2yo
o5gsdFsznoV7owyratEkmEnxA6PdFLECsNm6nXpcIfwVSLSBZfIPch7+/H0QUdQY
Y1BxSU6m1yVMxenanZs9qsNGVtsJTr5Y8zlqwpQX4yamsiD5xZbu8tgmI0VMXc/R
Glu81wQnEQy3eHW88QOI0jY6fecPeYy5idZBCL+uXfeS7XfCCkS6Yw93AsgXtjsM
ZvbbGeK+LlMy7OrsDDU+rfbwS20QmZlV2VxPatBhbZblzMFgZiOeG8XoW50goWMb
tzGpoCjaKOtkpQdekB1Pcfw5Clgu2Vo4rdCn5z+bBrHOl9wilHZoDZeGFIPib/vK
FDZlibMV9q6dMPYbNVp1thz2q9NqwQhWK/mQ9b/z92+C2ddGmteJWwsr0Amh5GHo
P3i18ZOwo55DerG+OoRiugs5oAFLbF8NAkB2o/I+3RC2Df7mF+d+MO8WSFaNPVx2
bavNmJLHOSXXWgGryjAvRQ4Zn9PWVuBTkTXW9rjtKBtK9N4FykqgNpMX13zINUU7
wLFpEAgcsAm5R4We7V+sLBgAN+BBqc3I31O1ooM6OMo8whvvA/v9ZV84yb9OzQca
jnFlWxw8SFPAUGtT1kqDJqjmtmkmDaEphT3SFXEzyaXpLeyOjRHzdfAptdcgX3s4
YhajJg53VGslGzoE0UUQbx8a6MBppWc0lSyN/im/FXD8dkHPrddk1mje+lhvgX4G
bcio1QzT79Uzjbdfn27M9jSU1TYJ0YE1SbmF3jXssXNw3AxVbaqLKkM7WU+73c8L
5fR9YJApq0bQP9/vQg8WCHFMhQqn5aMqcPs0GZ/+R/03b0/1YcTHW50IBaWQxxWQ
3Qw+ALpo1nVYdm0XgPDQgwIIuFLDmwDFiM4BQQFz/ZCtavoF7YG9NM3x2V8VaNEF
Cvzrv2rIg+HXWIzu5gjxSOBwkm4s2J7RNahH92mCLTA+QTU4Wcu8BL9CQzfiQWJM
2mv0MQuW8PEAYlW0sepKfWx/7/6/ry6hUIEY3MTzwvSQcFUSB49QYINsBCNXeHxC
QAvw782j14C8msiA41u0ADfBf4yMkyTq8EXHlvcpfouqDAI0e2tbVz5V6isEYzIG
uMnCETXewxpf2J1ZV/sbU2uV3siaZRMnT2F8QhERkfsWcmgXEhZasaTERvsINu3O
QTLrPLLwRmULo9VjziykPfHcCouII84oXd7/+WG+Te3lM6/a5dgqGzD5NkSEb0rD
+BNLIG9k85TAgIw2UMn83seTs5XKvJf9r2Oj5550KZs6F4Y7/5xH+570HZlRJbHW
OSzmd2nP6LZSQxS9JXI0HDsp5MChG9dMsnn8vXVaK0aggN6XBdDOUWKJdlv0EH1Z
xtZ0Cf/YoNvGh2BIoqemeUZ5Q2ySAuCjBhAWAYwZAUy6AkDXh8ybqY2GKeebtUo0
ks7kzS2ob/+LCrAUkGcLQSXUJWc7flcKiIScWGOYa0dDjbzKq8r3XlpOhdGj6RDJ
bH4IypHx6Rnvw70eZmh5YVzB+UwGC3qMy4qs5L2wbWJEdQZVQDjyMsTaWCB/2Zct
MhbnV+4/DqhBhZS1LVKicgxuMcrXRt5wacPHci9FBKNQ0ScqToMvMrmZs9N1a/xc
8f/KI/pgzDv3JyZMX0EKp5EauGyalv5wFEXiDMByPPalKpV+XiDk1e41YIGWykzp
N5tmr/xzp4rsz4caluKSQ4jhtv9T/sOylkvJYAhCTz36dJalkvNbShVSK0hkjsjy
b+JTYzC2wpgfmyTzcVtnDAtYSuuLUKT3iRLN3/LydiqhclBa5Wb53FxzBEdzqxHw
48YjvZGrXyf27gto6i5Fintl4f/zbYTWZTT6qD2YzALXzbt4EXWyunGjtjlr+YH6
C0WNcjcbMfZdyokz/CCmOzvIG0p4Yq1eUWOCVWq8Si8f69kcEwr2sMjrVSWANd8C
r6RYXHC4BwwSkLXJ11ea9nEWbPwD0QmejFqc9/m18orkA/ZQc9Rn5+hBiBFyMuVM
1/FXrcLjtPis0yrN8i3IV+zS9EtUobpZsND1kutVYOeUEYfxxGbLf/MGutwMnU9P
3SCiXgUxxmj8uxBiBEfl9hmhDIU3CbZsMz8HPHhtx8yb+YbDWMI3q+DS98wefqUV
qXoD5yloyucWGe5J249s1UiLHP68qoO7lRB3oYJ6Cc/bs4QBa8HFDxS49oIrYb8g
R69ssdfi+xAiYKSNZRxwpfqVUxHgOIQ8tCHwq2JnezIKu+9/3hJa3Zb31EyEDaJQ
zVh7Fj11P+e6NIkGa4szLQoxh4+iS5T8Huz7d5uUcoeuaLy3DGogPb7H1DiWVQYk
+hu5Feiauc5TTURHFOubWbWDxHgyY2POaT+DAer3Mzcl65AyNbMsr/VyueVoHvNB
koCzAF7rAlCqmhDiRswHXythnHY6v2SeIy/0+ouICpbj1Fd1FW/DzYoTJHoqFO9j
0D7I1iWuuyJM3NxyD/8wUMBffFeNLfpxCQLCPfjs1FVowfVNo7j/EuHLMwZqN0Sx
IoZ7v1+KJfYrrObCWOPo2v0/xLcnrOw6Rw3v2t0JXyz2CcjDP6AifYoBkPEIOMZM
VLfrRJf7yAzwtX+E2kfcOcU5qIaNCh6MQ5WBYO1E6AlA7MioTbqBqLqbQzTrz1kK
WJv9LE/RP+IY+qme+ucIdaw5AQvoCo8tVWLjg6JV9mkCUf12mZq5C8yV1Sgfpw7e
pcIAzSs7v3lL+tCPcHgK0f/SHVbKY7/aQE10cLab1+RARQxs9brl5vscGocMgP9Z
DLU7AjeKVSuXGpQ2KMTU99e3nKQTfbp8KQTtC27EvES6/5xOdmw98CaXduv1qfxi
SzUkml5ljyWAYLbCKaBHDAtqtJBuGNU5Y0zzdv9aPjSKvEnjvUX83LWZGZxr4kRM
NAoNLCG6Gpv+ZQ8DU+TEU8Pq02ari7MGnfFfvDOyJYHZVGvgs4PZ5foeUFmpT7pP
dyhDV69zIlaKIn2a2mVVMtKwZFFthFcwERd4RhVSUM3TCLi97QXPSq+Mbz8IWsf3
25d0jzb4Tk1FKcsLyFI9OqcsZUC/Xl+sYC+d5olezKClsnLpHIPYGkisfJfkB0w2
Pavp8GOJfzDVmQe8G7fR9upUTR19rezt8rHnQo6vwdYxEJx7XbkFgL1ZRKnaTRvI
EIs8HTZJLTlBmAGTKhyMD+aQn2i0Zmq2EUZ5q+7095Yg4FIIdn6TpiFG/IWqUxTA
EALcFBzccIHpspRvXV4xr1w1n3yQKNmGJooMB50kh2d5ccp6VNR2jorcgowXGYao
hkun+32Q2Pg94FeWfDUZ1PnrypHLKl8QFYOO7Ej92Z8Id/QEWPMAZ4ejqZ4u7nrF
jZiOE0N4BM0jHEMf0EysetJUUn/RkG4bcu1U5hLjhiw9893Pbp8juQ1tpn7xr8Vc
qJrYvOT+kzB301o8YnJEal/Ty2gFnkjTs0lN7xzth05GorKdwJZ4XkATH3wbuqJv
873cbc+S5JcbmTy2cJ1tnXoDCFFK3CWR1H5tzL5/mLQLXptA4toK+zrWk32AP+RK
nYRlP1CXumHRS7gNtJ3wtY+ndLiNc7mjc3IndKMpxEt7e94uwDSCDcDpqU9cFbcv
Wr8F+xfXSNlDcwHi8Uqo6Kgvy42e6zLCTJN0Zou/psPBIdN3zYAhhrkMNhAIgApw
J32dqxOBdpyy2Jj4RriHX2TyVZHxQmm7PLhRQ0mYdbh/U2Y29KXIPwYMK5rb8ubW
V5q0H5Ksbh/HS7CZEPR/CN2PeaUrSFX7XWctymujPNaICKAnfYByIt+dYYgqazvS
mhRkTsxHjbdLtlsTxyvvaSTjhvTbqyj4SmHJbchaj/Y4hesmjiNSA+y7nNj0FQPl
0GuOtIpSBVH/jyjNtbpX+AyYgWxe1JNQQy51w1qmPK5XhnzsJXISNG3u0jkW88uH
SsRmTzGMICbY9fWJxQaDtN9hpxrE1sxEH0Tt4Wom0udAmQp6NccXMagCn2FwGRWt
sg49XqWFsGU0NA8kNbTjogGLWNFgFMZAZNbqxm9H02ppMvJSkS2d5vBlctxof13W
8FDkl/coibvbBbX5Ekw+JLXiK2ZoJFx1onF1ZgmGEq8sP1Rg7l7hm3U0H2AxY5TL
fziSwEGVVMkpgmOEblC6GkO9ZpgATi0f/NWIqEFh4P1DqK0zUigZBrMz8V6+mIwx
Ol3mEqSebx+LwSKimJguNRtYI0yUDsnNQIXztwtA60T/1szhvVyS3e/hzsFGvsQ+
ZD+2J4yXcH36bijJWyB81bTyhYhb48ze007IHBSqeJ5CPrCZ3dwTbk/RWA1MPmCP
nc1ju9JZm70jVLuffzXhyag8i9T73Rwta12rFzqorMNU2cJ1V3gPGYenWHDCTRo0
2P7htIYMxOA8yX7qwa4sYrd8jr6BmJ6px4vYqjTSui+0tdiveHWN3ZrvK4DfQinr
x//hcmjMB0cNNNiLvwtbVemprNk3dTynaK+EiKWws2xRKmp0lyQV8VvP+0NstrfD
j6IeJneClXZ3hJHzQXx9MQ3HzPvQtVhttC6gii3eWa4wo8hOXtwERTvNHpEqA2X1
FZr+KImWsV5ZVyEBcqvN6uq6RwgKMjGMTCsGuHzN54OI7qyExzLRAB4mfETBYwIO
NRUUCrY42UdXewqe6y2/8tCjn6x3ACSUCXUP6Vs2ss8WNc0oqo3TmPMD7W0EOcaG
43sCB7dArm2Mb9uIosswSQRmCvqBS34CRMgK/ONoASGSYvBQVTmioC2V8zmxXf4E
pUJ6N1bAE46hB7yQtNaDUYvf9QNVtKeVbPFzdw6/ZJXbOD+EpQ0j3KLGdVqSaFhx
VBxF99U7uzzAPjuK07D6nKILCDfKVmTHawMYroKbxn3PcRuhUez8Ic7WzYTLnGYY
z8rkqzg8+HUd1h+L0jYfm9lWNqpF63hlrKcpCrhGtqDGeWY2utCQCu2w6dTmC8M3
2iguoQkwZzsqc17u92n+EIGz+FM/V3GvFrcOkqHS7sOBkp0x6kExGHqNUfUX21kJ
uSkCKVr9QrGy/0qvd1XABdCWuizPmBuVUD5EhR8JYmJLEEMduOY6vt2pMSGeuIoM
AqEqDoTeqNgvad4h0vjpuJtb6kVY9oICk5kP0OAfgS1FyNqaMr66gmLZEFMVKSWO
XPA0/9pDUwo2ZH+x899oiQH6WPZRYK7CmH/OyCsNWDUElZmJN3+a/0awwXJXEZH/
mM2Zqa2ITAkVCNF+HW6+QVVAlgxdmZhwUP18IKG+Lx9JIaSFVnjDffW2SEbexee7
aH76p0O7mE6qPBkV3StCg6hypWrQse7KGYUROIJ3CZhlKihk7ECfhxT28h4oEYo7
qlZ4XZ0F8r/9nz4+saNa5HNIzO6A42o3zL8agXNQxlZZUJQVcCiigE8FcaZiJz3d
ioCOXHT8zCjo9pMoz0oTeVGOb2el7Kb92D81TN8Kgk0oVbpadqk07scWfX1d1hJ7
wOq8g9BxjS8FI/95YFopLLzU6KTgu4E/PDR02V08Ci3Bop6lzPcHRo00uGMIu/sr
IPowPeBDFat8A8wPabB886SmBUgntBMi0Q5w2DPm+stbO5GXqDr/lmFsr+olgc2w
oaLZ/9X/srIKcS/ts7GYuiOrUAx9C3dH+k1PEB+mq4Q+G0TOpMb/En7wBXsK/t0s
I5y60Rub3nkyQLTnNrwMuB9gMBLnbTjVsT6ssN/3mKPOM/VIGrhQ+R4cxs2krEDE
TmdIdUMP64QacY+2ohnuKxFNxpDSxwOlNCusxpOemmedeQOCJnDiWcs4ZpXeRrrb
pBpbLwoGiihE3m2GMGVwhM3O4RIG0HcdBRM7pxPJeDa5PcXHZFoYbm7DQhsJoQXx
yTxWk5SqlcR3cngzJTBR1yPhbeE6TpKL2xenFb2DBN3t/Be0OBNjkoxe44dfeKb+
H7dbsOhKDeZMCnSCLxiWuIH2U5g1uUaDRc1OonOMOiw4RaKVL+/bxu3L7XYPg09D
Iw/I3brV6TJ+D4QEMBFQe1uj3ON6WQbHc2ppF5hLVHEdeF/4jNKOgn15r0upRdAT
v+tyayf1Rq1DmFhubmw/zFamT7F45xRRJ/Fnz6LDFP5p4CVVt7NdDpnAAAiX0n8Y
Al/7AXx5ESJQ4m18NFX7YFiJ3YOw7utP58uDCAmFjSIYSdsJKBHbDTEJMXDxGrgo
hx7gAWWJccxcB87FFxIlv1ufYC2WL5VnmySUNqcqa5PEouRZQfSPqzTwBIs61WOW
Y+Uw5LHxana57WAzdKcNYgzhIhUmqM+VJRHo9O2+J0Ex0CZ2Vva8Xno9K5ljfyx8
c3KpVDEb9onSmsJbhcBoWEZ5Ffh+niMH04oTxXrRRzGBiaHGb06/AllZQgJm9WaT
Q5glZRofz2d31deejJKAasRG1XDuj/XsmV9HYqReXQzAxJikNjbGpeRWSEpP8dvQ
hkKhITcIX496bFp6t1Ulmm32uUG1DTr6ptn9cfoJwpS3ixm15FfJ0FllQ+O0PBpG
x45h8TUW+GYjGCqK+qxDdjuIIEot0odkRe0dWv/f/475o2YRzfbkAxGpLDq0H6o5
r3Nsjb8c2PPGC01vfDnNUFzx9a17U9qR9koNw0imdnQGzX8S6IioRcGGGBuiQ0Sp
EefBtEWDGsA2YbMeBqaSAJNyMsNUVPTzExEZVf07BqrDFhX7Uhn+n9DNUYxPhkCB
FIR0ZaJ7oLd7u+1CzfrZMAeRxvaKsePN/uhTvlN0ONWGs0W2qCsxU9h4Sx+zMu1X
K+1XnMu6GnIEJOKeg/nUGaFJgcUpu9sqf9cvg1/Y5lauoELDErrOmLYYi2sTYsCt
bixLIktQej9UlWvWR8zf1YjDx0s7mPTWMQ8/Biqmuat/BQRPyBQVROV03mDZ+CVE
APd9OnMuL39StBq8NZwIU2nuiv9DErzbTxqpLCh7Zyp+k3EXuE2Kz/AbO7ePXcsR
cJnKmnzgNMEkeMj/s2OmMyQsj1jw2WfHXuHL25Co6Org5re7u+J+Ivbyf2jh4ifZ
PfJosFZaRgCQcXRINc+stKNuLpcRWKJlxm3VubMkhfVFSbTeOj9U+OBXzj9KX3zT
o5CEjWXz1BQrhGBFt21BNQZkMjfusn0g1jRaycNMEZmH3LByPAEwiDFo46GDYeL9
OeSqXPbsVaqPOlwTrckQezVKAP9sqE6bWbQNfYhVY0WsyjwWdX79+mKolmpqLJ4m
E0jKddQquSptWputpGOawbDx92U41ygnEYaTv+LsuTS6JW1NluEdUWQcmOdeNey1
2XUXFQG6Xs8i4jITgkrLzocdDgvQ1hb31+k9DeLHwntFaLetE/rWa3GpRIogpNu4
vZZB8CG8rmNG5cLwql1vcHyZqVMLA7nFOT1Re9gOqXgUajW6cXEAxlige/lx6I7N
2oHti4oQoyYFYcGz9Ec6yMCEXUTsSZ+Chw3lqYNHuUTUQhw/Cd9I7KGFTC7eQZ/W
4+yVUfTP9RpInHN2gNZ2N+dnbB1SQp0Yw1dB1OPaL0ugLkbrEx7s08LnL09VRwdb
THCy2/D0SoUtFdlSxwGndYRkHS2cyqoVP9opfVdUig1jICFNoUynGhmofKNRby2m
qr2v6tdBN33G+2KDNUf172AHR4twdCLtNR3BZGcC0X1w7mU7hsS2Dc4B9eHx1qpU
uJxqrL70KT3tCL7vy/J3aAYXIYPCpwqVB5vJDuP8OxExOKCssaU0JnVBqhWqNpek
9H5ZR8+sf9qmGjo/YV/J9+aDW06KpxnT1syYOJFaBZdZy7axO57ZhjdRnkaNFlvB
0bWgQSwtvziPwkW2cLg9PtLBw3B/Tgr1iC6dncAvPPP01vMBm+v+IcnJ85dxChl0
Pq/Xw9MndqLIsnL2ae9I96SPCfTOWItgBxg+D1BYcDNq02Bivb/pJb+UTugdOgjU
EhWEZaVxnfzrqLDBRLZXSVnQkxcFeqhvNmfiwqFg1Pp7LHd8ZZBRz/RQt41RdSMv
dV0Pnf1xcH5i0v7QlU0zYwdmajET6MyM/3hIkjo5zpcv10X4WX8uCNXBthTnSJ4S
5+lpCECCrzhdZKUsCnZJIpwweqLM+naiBZ5qJ5oYM1Nve1w5xmh35iH7FMYiW5Ly
cuT5SOeuMn4heNhOWTpr7++4SiUGA1Xjn1PXh+iqYzAkWxn4fSKXWSVJIK7cs0ly
vOTjtskcN++107kGbaU6oy2N8Yvm4wPq9r7QT/nvMtcw/Ru+V72xUR0H7fwqAofk
uLjBY7WUfAru/j3IopHL0/GAaA7BVKD5JDW5iS8rUzGLEHfXA0qCTSAgIYLWYCKL
iOGSoE30j0l3rYhX1noOkRUdRkByqwb+9bWCurZdWGVZaR1TPC0qruoWOQxWEDbi
p/8f7VLH8f1Rf3gb30jD+m3wmWAE2RrCMhKBN5m7tVoSPaskPIKL/vJS0CE6WzNt
gqAzlXP+B26PduJG2adqFPRR3a3bdIYdAeoAycx1NVWQ0tvi+qcmuBo4p5JADj/x
DVGZvYCUeevP2XoKyWnHXE2sbbMnykiKPC7g8Rr5jPon28HQQI34sMA1FpNEZqDY
Y35llTmZhZrSC8dO6e2RHIKinQJXl4hyD1tlR/hDibzVjEYXwDU1QRx6CvAEGr1W
QvaO+yaoWfYj5SLW0LuennY3NWOu2ijEfqiOCQGQQOlyg2XXXl6SjpURpmr8FxZj
o7ELbWricWYrKeyndUThp3iliIzi7Xq4z7aF9G/4c7xO8RfkXV0FASFcqilYPpUD
2jNJcWr3VOmvd6LlE0LUuZW8SwGg9FvNX1DsQYImEco70VOxwDauSWXGG6U6swlu
mn5ZTymoE+hBq73MYrZuCB4dWu17b3cAX6i29/NJ7KDxv7/WVmTm8AkHaoFjlPvF
eRAJsVvmdwBV2nPHuUGskOg/VRvwOBXsMEgW8lYkijzTsCurE0jVX3PHidJtPFxn
MorSb2zi2CdpQfseO/bBdnDDGCbHXBEI9zg6BD8lMwTQrmKb2wbIxKgDUJeExx4s
0NGlO2YyRoifmuONF3HjHypQbd4cDvXctUt9861is+qUieZOrtjn52Fcl8yIolKh
BxPGpdGeLffg1L+B/EFu3xIF6xV49CyEUV32mr9UAHOdZ8SnAIuE9VChCf3mmY/1
0LOmVb+qyh93vWP4AL+4iFwnvPWEMhh7bneGJFLx3S+rY6I9AEcAEtxXdjyCbLop
HlVmhmW78WwKqb2YQv7i123y3yFLmSZ8PjgFMo4SQRqrOUgUG1x0dc9Eqop+pMTa
50wNz3kt5xYkjki+tLXucwcuRDNDb7KZFSl044qjkwwJLQOoDFsWa3QQgV+dzgCt
QNrsYOzuWnqfjvb+Y61ZnjFhBr1KYLVsjCzd3loW7gyeeaiDDRbCrKpyC+Ox8+Oy
4rYlEi5olqUdsrmGjb3h4oiTqdEMl4pv52ZS8hCjuITD77mTuG3tBAg+I3IChw7i
H7I87Zyq0YNjUY1y0kRSQOWRYvGDVSROJTjyh6iUHVYzer6iOucgAZdutgIVXgWo
USi9VduOpkBfLauq2fY7O558wgRWI9RNcvRTRdXMuO+Kfkrrs0UZBrl/nsgDtc50
sBaR9Y27oFUa0crRlx6QaDFi5MUD9DZpZa23bnDUE5Qi/lvep3XqR7sF1nLfTlnt
6Jw9zp1xxPrxXYwFYmV/gtSqi4yseK2M1xhNz1cl7DCzZIqpp3Ixe4KLQsVBPeem
c2CZKq7VPg8+/4qsztnzupDOTw44SOxMPpIxkFOC7bDevzFj1vGZsoLlZWpnmDrl
WVtT9ZHIZ+2VB5iRtv+czbJF4qrxRkiCgBHmcpnKQ12Rvj13PRtzn+h8us1NsXIs
Vspmcef5fXT9TayEoTrwBY/2w3F7ayJq+nBKUGg4Ot84sWZjN+RuSGqigGSU1OP1
PZrvJFC/DgLas2ZBVCrPSarnaeaZhGzAz4ATI8cGQG4GOK6Zg9lSRfWThSC+aEu6
ThcvGq2df5a70BhbS0JWkGCriFY6sg5Xz49pY6Ns2JymdnklbJhsP6thV6W+zgFz
vjsgxLwcRHzsEGnW8vVj5dATnHFo7Zt01MKRbuRwER5n2NyoMo5lCARc2mer/Yqq
z2ntFXOjIlrl+acCEjCqp4rpYPBnN5LAaJJtJOSyneSC3uoc2O1XMLbqP6NglA79
qQnC/E0FP3cD4CfgmEQrk7Om4Or62VPeWxUOtfQmZA8HnXjUhGBONrcDetfgmTmg
QtO+kOFK3z6FoLw7zZj1kpVU/WlP4vvVoQS2Xjz9FWc3l2IV4dUimKTzFjVh0UJT
IwJcIYhm3XKT2R/BVpwRTQ3NnH87Wc4I59mViYgmTeFXyWZkg3ft7EdL0zBnf/q/
HQu0pg+sHrS/5YQpOGrk/JrRU/dxivJeA9CMVXlJ4kIYG96Pdvb84rKOXLFFd0cH
kSL2sSgX/FWdqGrl9+b53sXmwzTB6+BbIuGjIiT3cqvyo2Jl4QCScTiT2UoB24aP
CdVkA4n839nf+c/2fm9lmzMQQJJozXU/jkNcy1L9ShW4dYPua+VinUmhZFnAwmcG
tioQpdrr5ZoV1AuEqOvckLtBeXmeumSxiX/9xyCfRuLfT/zokhItmDcMI9ZERtCW
DGEBrU0yDwf3C7yOHiM4hG/bE13L7VTkdpJvSjomwvuVAE6BYivqQTvWjz4E3hdM
IdgZrcd2ttRmKIapAzAQPqt35qM5XglvGYLOnfdsA7BbqcqQqAY2s3ohMNJUjGVj
kOsQiBz9aLJOLsoff0HqKLQ2h+htW+jBqSoJjmU+EFc5o5eWIJ3ax1oWbyez3fKW
ZKKPE9U5fGce0DKG6K3Lce35UGSA8m2U0otsGtbTJVWPBMz3mA2iGPO6pzpTOJ93
Kyddbg31LS31CzXukBrrY6wJa5e8eb1la6XuW8PpMlpkRWdECUCgAW2f0ByjbZP6
hcSOzrWDfnR9ujefDDEI2OzQ4PoS4qT+8OE7K09qyxxTVT2WwwfvXpE5Gp4tGx9g
1dJLBuNO0mr0J4B1HgsBiK8Plol3D+GMGD3UdWXR2y9ssMJp6A86lHgNRtp6nV3I
pa0f/1GBZWPSpBPja6mNbn5VeBlA5mCvpSO1/QKzYJLo/aGMWwCFNS86QPAoTgHi
pChMyuLVbsWFdHuGEoFlJwbB6oXy/L8F9B7zTvS8YvhjRVbnsTYdS1H0olY3HQLG
oi2vo51HWw1PG9LCviYMhgUQf4BJ4ginFJJwqEUjrf+8LOX0O9D7Q1ZLRaVO+EVr
7y6iykUUth2nF11NbpIdV4KrUk0sVkc8eLRnZ7TM/sevtRxsmSrAUHvMroNN0bRD
y2tBN4yWWMvQcpQ61X6Fifl358NFAt5h0iylO+7Xjj4JdHVLpBxlPWPIqKmZUx9g
Vf442XYQNak8i0jHsORH0YL3ixNHqSTO2cBFLrGD1YepUh0sf+nQX9Fn2lh5ig32
Rax7yIsUL/q3cxwzV2vc/BUuy9WxWSHQlQdnZcHDOQIY+hWMmVYWkrQtOEWN5H7q
YyAvxQ30sKOc0cnR7r+SHCNhSP/TQ+nrwzB27Q415eXgw0ubcyID6eomBAn4P3uS
aXBigCQCMlFoxI27qCaOzflCmf4N4tfrlicbFA38eY233Vr8Npkcq+AsIhuNcuda
rslsDrVIE0mf0kK2ugQ8X74wSYzmsqEvYkftfjiHP3azmPHlluwLKVMh9b13I9dL
fV6IGNcNWnt0R7Smu+ARpCIoV9I+0xPRuSeOYIkcYsF+EhdspNhu1LKYiSCNLcQe
emwiZF1/LPdgwrZgLhqm4jDGbHGsfyUrnk2vPKFz+dw5apSWSS4CBG8dVVSleH79
f+K926sBNXWYx9axqcke9GEiJzZZr4/GcWRIdss69Lr1zxNFu0vC5bDKou+5RzI3
B2hRvwekTGhKpNL0ViEtVK+R5d2YiJuOm6mSXNIXtaT7p0uEDlGICeAdL3QWvNf0
EDlEW3xRmL3fPz54KwBIiUSfyEIfWt81wAh4GX7ba3lL2M0v+h3wqOVaETxPbzRt
SGpfajQRzPG9ty9YwlcbnAORa0Zix6tYvJC+V0BTy3lLl3M8ruZ0UiI31XfsuNs4
MsmYE2trBwbzBI0DP3prDgwLpwxYK86XCum69iePYny+UZQgTpf8BupEgTeg8hBV
YpW+utwVSq/htawVwG6N5VXtqUixRJqv4YAd/IRcTGiFCPqc2dct4tSigQDL7jUN
SJu1b8lkDS/1TQOHzrHr0zx0UpM4N0vvt5KTpgF6/6CbExSxJltzw0e0BfHWHz4F
on/f3GYW4pc6U29mkECLxbgstmBmA/xU/Oij47X8+nNVtzgU688Na8C+kGG84cQl
B5ExUhe0FKeMkIM/hk6oCy8YXILrk0IyyCxHR/dQJ8wnBRA4vxtkhBbdegtRhOe3
12MVXyiGbnTwp18TrYvjdBD5pDnI2vOuQaPXECpDycwc4STeZUahpO95GC7zxAnF
5J1fuZIHe6Cf/pdSmQxnfr89e1R/9N7mm3phCVxs4005AcVYSnDDkW+OCH/9y2fz
iIgFY7J5jFOV/02CV0ej5fC73ZszAy4QxkPQx9MA1c5OKVYfEow1rqrG0hk+dftV
XyfYDTLhHA7CM5NdGgXDXgnDqxinjovLjzisl//9ioSOYOwnj+gnIkGl6SpLbx8w
M/gaTB131T+ayP7D2FY7cz7WfotNnneQsmXNII03SCOiX4UvDegvlQw6E25QA4Cd
eGaDsQ9PHBGBV2CXeFkZAbtS2VnpoUmSM8wh1AZEyjmMn5as7OralcnBDexANeT5
tQsDREeGBr19AUxxkL4w8c3G7F/aIVsv084aDucgimC8bSkN0Jci1vYBySAcgtuK
x3Ta41nCyEq6Dod8S0rAxfc5AjYCfCVDS2DaGg42pzvyJB0cL5BLscVZcSICBtDO
qsfN8yoURk+F7ThdEgAlONqH/ogl8LN7PEQnl8cqdbX7tKd2HZ4/sm2zGrX3FOTQ
od/3pFa2y1AY6I6kaoJA1O8OOqf+gI3LGHNyVfpq/0vxr3WE339toFWiE9hSBcAD
tBxV0jdYL72LbjIXzV6Mb9bE/ZyvxT7eg91bntpipYPIDBve8nWzvJKTrRqgIWod
v2eJBCsTxHzl0ox39JfjW9MGTiaFEOwD8/03npfnQwdEPKDYjitN6ENaEHkDde0E
XpOhLL7DoMdA+Vediu4lNgBjV3TcWeFMZoGekE3abndHaGpeoJw5TjvsNMeTKE8z
5NbVsnF3SMO9s4mS+ljXqprBUicPpBTSyST0P53RmwnUCWIZbH3flAeMSlVXS4ls
MwYZcJGEHNjYRHUY4B57OjfafA+CsTh1z0WcRYvG49+qzL9shnomU+Z29O4eH/Qw
dgd0flteaflEn8Qtrx5P7obY6JsQvG+oY8a/hzKK8HU90LwUEtW6Gy3Xo/V6UCxe
+ogLAfm/YuUoNfq6LTzOy+hjljTA3J15C5ra4GXxN/8Hxphz/3QIL1AaBgN/koLX
9/bJzJ4eOrtDXf62En4fEUhbRjiJp5n0XJLap0cvqPEy37zWJCdaIVdOYvvS+GNQ
s//03LnVWh0DU+uYTO3yA2r6Lg5chlqBpqB1eudYgfEzwNXeNm/H858W6VHoDd9A
F/NNST3n8njV4Rrn+/suhJ59PdWfLOhtYzX5rMefWiOzbx36R/SzVnvxWzV5XHYN
d9sARYwp08H+2hb0lThD+d4pstBAme1WuFptDN/Ka7Ebtz5CtFavdTwLWFlJqGxx
eIVq8F/rae42YU4RwpHGkxskV/06IM100BmRFQojQ1G/zqfKV4v9VOr9rhHpFZ5t
Ps5oPBSfWySfOhXnL0zA3FPpfwUBP7BZ/K91eMIX0NWfRFm1kpgUv1YpHNMma6JZ
7EmwzJqzGFirH3BfNzFd/6Ths9o5Q7uQKoyjAgdzLRy56tx8BCNIjsFWoNyTF2EO
Uk/orcOQJMAsxvYZRFQgU3I1psZiY2NBNCHANaWxsZylE0o3Da+yms88ck8icQQK
2lVZx/Zi3r5XYGh7FquR4H7fKp1RVslrSVfKfpF2VvQ7z4fFq5VrZcjAX0ETbMej
avquni6turw/Tlexv0uhgUioeDQK/rfzuuZCQry8mbeAJHapN/UfIbHtDgLoPQYw
H6n/a5aaCxGSka8SQ/DcQmFBIY8uQWf5bKKJzwea3ZTYYii1E6OOaGy+mKr8TTzL
D7f01RjTX6yD/a3LYfqDP+rKkOO1s4KJynM7pt03zre/T8W7lvHqu8H7ATNKfAER
BX28wuw8hDz8KC1l9PeO2+hQFpJyvYivBq3XglvqaZoHWXTUddJLWgiQLCipOZN2
EcZP153QRuyktkWvVmSJOD3r+xG9F1aRqG+DmTtBX2eQ8FaCGgJCmh4fqXUiuZ6K
/JDaPObCQxIWDqZ/hwWudMyYC9gr/sOdkCgOpeIo97S0Q6M9WsZ5/HcRhIIPXKg0
9YP34FoHLrBq78o0tpX6/dvDpks6HNBz0z8Ej/2xaaB1tSQUk1u1WlLE0CT9k/vQ
7pz8zHLw8vFeF22UG+C1EwtqjjoRHewU2Gh+BhX1mVHs6gPVfMYL5a2CwsLqVlK4
B/UtTHpq7gjcq40VbNsTsxG2zh3FpDQ4RHO/fucf1gOJZk3406ZYaf5ChT8ucWk7
bWGl4DdbiGTTfHP66iQmDwF9v1tpsuhdT4xm11xUMGL2/oD2boJD58rIo0DaNZVX
cMnhMcoMSZDJe+ocOI7NlqOWlAvk83HuuJM/5TTB2KQfxuRmqWoEPdplbLKG/YNg
WHa0MLYRjjqYO4MrUetv0AlMrQYzSFKBRNm3NBbAsx1En4R17L1f+724SVAsQuHK
GFpPhYQUiA0/26ipUr4gAoKo/+bgxwm9IJYKDoAb/ILHIRk9DE6+3fbzU49cyO8a
AehLPjXTeLmEnD+PdbcM3wzkK5D7p3WxxlGRAJS+9SvpYw7gvh2lind36MWn7qkX
RQGVhxuLCGtAzMdgtFa2Z9r07oG5M7vl3ypC+j6nEJYZLL9P1P6/xMJNs9cC84v+
QN/87jhrf1jVB4J44dHYpb/xuB4zN9NzHsq6UTVHoYF8CtzKsQj1duj9xOeppx0Z
OUPyZlH8oMqNZNajkmyAZ8A4zheyk9KiWwY1uKOQ3LtodJuU8eBn612UFqxBsZrl
FeArp1D41APQUub2hiRmONBaUsrZcM5Vcgw9iRuI54mXgceYLtSUIYUR+2hiQ7+x
81PXfWhjdL1ex+C7T/Zo1rlL0Xqir7QXamd5oNVJA4egWYtpdnoOzH7Tcje5vDi4
PdyQ/r+/wbUHAgtE5EyIhipClkaiXYGcDmj/3M2Jpz5OpsZDvfbxat8TgS0UKUQ4
wXXoJ1dJk0qjOzIRiGLBxo82EJIKNAGJAGVN5xWQSqjCWoAvY1o7VCw+U8nsOLkG
vT6peWgDRQPF+MZVaepL2WlFJAnfiw6rKPolrxZ3ZZQlVU77gUeSErYjGefsiXx0
0TcAd0zi/jpXmtltZl8rI4lXoYcOzN5qFeJOiZMnficBMowvLNPF7SMh4nJIawHJ
kJw8vXXDOnOK59+QEM22AH95ftsudrVrm6932XdD+6b9JUxxZwNAiM3Qh/pSAmik
vxnCCIA8org7g8d8ysn+K3azXhovCz59d+vJkc5wHIa6CjB1revITN/90pYeh5Vh
3s8oIvu04LrilY1uki2MjQiS7LvjcOvif2IxNjoN4rw4iZyovivoIQNsy6/YKGwu
KMwC6p5fK1EWxFMChJW45vxgbWWoHKFmtmfLyaTmsOur13tgCHOE3oE/6CRxutfk
qgZMFiqL03KUlKA7NJv/7fRj/lxtxnII7JOl+wGRcF6pF7hmYAhw9yUQiQt/jOZe
9RFfHLLk1zCyn8gwdFk7EG4R0TZasNo89HqvojZMHualv8cvN65GbQOoe6dVN/l5
C/Lt9bhrE2Y42w/A9+FKYQZLYXsy9DgMfrkjDdg+l9Q0RsXEnq5L12+GI+kIPVOa
zwciqg4BQgLsLqFnbU+OhX07+X7IE9ezPlmr5+l5MxFopBmlNw6EPL+NTDHQpfPx
Lwek3dy8iJKYNZ1H5+kXjkHfrJ0Cmm2+op4SIbwEND0w2RwD/5D5voAZnxriqoci
JzyGs2jlsJpguzQccqQbDrDygiH3rlLX1lh8ZSThrP0iPngaK+tATxdn4ob//4fP
QEnGGGHHKaahVP9bnIxkpglGqcWkySsOT2rLlWvHoBrpmnuHcaii1PieMjK+XeV9
ocmzZG/oXo+AUPZykGbtC95Ypz3AgkKwfxaLx/8AwkaPrd6Hsv1P0JnSFbjsNTXL
zKN/2nBT93RlqK4SyyECo0VbrmEcFvRZqnNuOCLvcBYO1Ih/Ju247aBH+pO1ybJZ
a7YXIymXu79lagmFDytgG+IHLC0pEm0LzT3SvvIG0KSpX2u/APbqASEhXvKt7YVO
pbSFDTvAv2r6ZF8vanBZih8GhFcUu/Vw4EXHtok1bLUlvxkA7M8SS7O2noNxc9Uu
H9In7uZHEUJ8O8lEWjY7t1Y50d5mZigvHpR/9I27/VkjyRx3osNqBDuXAbNoBZm9
gWrAKf9dDUmCIjdc5235nWKhBwAJleTSD3uiWgsqrFpmiPwoy4RctE1Nj05eXctb
ClGJCMSyEkHSE+61jrVcGyB9bSbRbjR9t895aCczrLGJAiYgbeorTG+Y+4ZNWc8f
LJ5SoYM7boBIUP6ajsRiSSTdWT/NhQIMfdXLQIEtGKtJLpUsx9uJ9g4qlgyDfLQE
fu/u2ScObflToFjhCXVE2fIUzNgogNVHBLhjWxp9Orrh/pg6EK/+NK7maz5/XFMI
TUGCstCOnXIge/YzIVux70liswGnKqnnIdbBgHmqIB5ehO/4lPldyq+74BQOnatZ
gYPUmxNioIBk5k28tuptXbDheLlN65bmfgb4E/+FN5u83YYeplQfCGtB+usfVTPT
Lcijxo31TFVDc1O31/kmfO2pjXURDy3GQmkVDWt7O4TD++BIaCUq2r9ZCLaWoIrn
2QkoQNwnQVmilYUVIvrRDbDSJEGYKiiE0m4uCIAjx6V0xlA9QuXjV/v2lViXoGuk
HTLDEMgXxi2csJ3ezYgQAOgU7PXw3EYIHAcXLML9vKq26+a5A/etQEaMLQx+nxLi
tKwvsNTADhKc8dxNCwuvEPgZNrT+kVKSo1E49JWRtvqJEjzUc5n202HowJFNe2+3
Z0nEVYwjLxpnfMuZhG7GxrKWCFnRkp0odq7DBxI04E+MRtkNfF7WCCccGem6THGt
+FfSchtC3DhLs0tOEemAlC+ETgRvMLm3G1PH0qgWXaX/kUSYLGY6Uo6szmakxXsc
oDpCgj+PYvgrhwoK8MM9+A3dFrIc8FXOK+lV6nTv6gW49bh0r3+oeh4ON60UAlvg
Gawm7Jz1dFjm3bzwudxouaB2m8Ab7sRg/tOh4cv9o6fmt/2s+XB6yntHcMiBSB8E
SwwkXQttrD7TS2Ig/g7jxNUTNUADZJRsqy3R23SXYl5GJUBpvCCm6gHCoQhRewfI
fA6X92h/kxlD/KeASehp+svBQis0QzxYwEnIrhc01/aNx1V2sAD2WOa93XhfEfAD
4PEnDsTvfTZHk4EZ9VdVGRyN+QByUzh8Bla0JSci8o7TbLPCcdD6na7TMbGvLnug
j13SA+CYOqj6TfJVIWp0dp/LY/RidgL02AAo0MWFeZRv2G1nJXhoG/juIVnNscUZ
j4pResGbVRlIeVmSjzxnrO9fnVK8IuxbcIKxSw79ysMoHrodneYo7q+SFL9ivuio
WIU4DN8Q2D3dmsVT0nJfTaeWuvl2J4EAZGVmS8vHkH4kfQn2onnVplJ41OzaT0nk
FIoEW5cJAv6goni8P9dXNvrTAezKxtO1K7orrhh6DUrb8mCLXZVBDKYg/lyLHb1y
tn477diuqHKtPvWtzmh+k1lX7HSDFxiF/3xidsrMJIKE4YDTjbloyj6Qbo9Gi3bW
skfHr81fP7OAhQ8vnWhOcRLqu7t9hf32ALqyiYsUe7kRfjt+nrWK8Pg2WqqeBjMk
IgEYVpeGky6+fsuu1THww8H5MSWj1X/XICDnVNmIvQXYro66tyc7QLVYEGzUVYxo
9X9aqmKQuNwAfbXz8FBX0suXgviLvXCuiOWOUzvZdgikZahCJlfA0OcjYz/O+7V5
9JWeySjl7NDkRiTz3/vrkBUoG9Dx9gCzLmT0OYJYF/O5A6u4I6QpcGssTgz/qz9h
bM0Mj9pBg5lDtW+m2R3FbmnldhkKsqWCSEi4QwHvwhvplsCKUxOJd7WvIXXfhZlW
kS56Kv7D815yt+YdBYJtzDpIXIcPITRbyR1BoHVAHfO2nRxRvsndWdrjFB77PpIH
9SZEGnEmDDFlj8lcKB9yTJpOLK2CfSKpYwVaxmuzHYfIY1kAoqKwn0PyoZHOrWzc
oXe5qrwmbTUP8F09WRooQY3995ZUaIYcLt9a+DOM2X7Gf2ZdsfG99xqaEJZbEIx7
4uFgd4FOp8wpJCSnux16LWGrlsG0ryTvH8CpiCSsh+IpVQvSied9DgNlLXuq84L9
hBXzYzQMQAAjmePpkHASSrrYSttAy1bPW5X5i82fDa5mmJU3ou9/JYBMS89pVAgs
iD6GB5QBiASSe75bmvPILDOhRs1FZCuuQZlXsID29QZGP7Nli9JaJAGCWjxL7IoO
q5XPqs+2X3tYgQq7AuZuRSW87ipmHkWdd3ukt0SSI2dniICvlx8XOKLcI7Uyao4G
LxCkhnHTXqjJlMNN3GBmYWOvfH470qr/vh7CvUuw+vHEdxNR9Pw3YNpJFjnH29Aw
0FYETh3OqSRJBvmp38xr5BTOT/1u4fAJsCfgSbmrNltnmMSxywmiBsCV5iVCgouu
Z4Q/snoUbujFnCmsYgr70i7VWC53tJ6xz6oqiGKQ6bJ8wpiEf3Ye+D/InSzLdhHQ
X6z8V5LDqBLPvk88p9KLc/bSGcpWxbAO912pzPaLRMXLNk3PD0iCNyj2p9w60swg
LKdigNDSN7yX3A0L3OP9wImL4YTo2MGGSimYsEIaSp+2BTmJr8OCNSbD3eC9MQbK
yri1qdhhcGMAzVUMzHs0aeo3ukVU8wX8Q1nMkTJhjxrRGAHDcompJIiVC4CC1hTE
MXQ5n7CTVLrZpzXUWTblL+LIELXlWyJ0j30isxmqdKv3qOevhPKelII4zcGYvFgR
pDlpJZcW19i7rWL4DXgZ6yQHq4eISVtl3anQmG25hOXIUyHEJ06UBTcyHZ5b2j+x
RaATvuniUhTu90mcU1s0f3TyqtcAQLUMIIKLBQgWDLG/kC6Jo5JXYMSX4JE1nCG1
loohurPDygmKrq5H0q5GdxWqnIal0cIPWg1WUdmE3mVZXOkSmwH7pRuwfuYXZTOG
CegMgYd2OmgtRdJuitQCQrxBa2hMVYmstqtSLaJeap/oWsMQnAJ4PTZHax+DAo4+
OnkMroowa9LX74X2C3ZySzphJVB0DoYL0Tu8W5f9FtWXPG9C0iCLatauj2S835DY
QWaz8jeJxLZDJC9aZnvSoGpAMsBnl4eP2Nega5rhOVNnaqVfyG1PdJqimgob4r4R
MN+HkDK7hvC11SQ4HAJ5roG6xw3xKhVdHanUgwtZCm+r/7G+GHse0kaHWlFUx3S9
GggwvsW8zFHWjB9f3ifGo4QeGQO3pyQ48eo1f8Vmm4jPIXC2fb4p7pnQHQQ8x9I9
KTVd239/zPFN+78ubBmu2bJznmWcCsZp8Ih3YDb3gv5l75JEaPAdnWl+6BUYnj0T
/7QOKVzBW0syrw+RW8fgadbuRo2zFjHfefR6Odz0iCGl+IY0ZSQzya0ZKitwQHpj
ALe58GW5020M9zKGF/EdTQgXnMl6xKNlP9w5R7eZ0hyPi8Etp/QyhugeKo14DcVW
HWze4I1+CXLV4xN6/YtOIuGT4XjT+W83Rv1buOZmRAohBVq68OT/sCNS/Ym2SLVi
yD/gFlScIpXfBxuoU3Lkx890nG2+19ZACtn4Yrzv427U4Gol2kbDJoCJQM0k86Sw
2wquRfYCVjjQWzwOPrnPx/DLEZCm8evjxoPIgtEkJaTk+uedUh2y8BQuQNb6tTFL
4+tLozbczZ1UBYQjgqabgkoBrjl6d60H9cJOgNTCQdNvUwY+aF0Rs/IhnTAqMImI
pKLfw1h2KGKEpdyw8ew3SIDpiDjdFPrWKx/UI981T3AMJ1jDJoPVWyE6Z8lZ/PLU
I2hevmV3J9nJ+7vl7KRPw21/HXBgDdGzQmJqPHEh1304FkikffMtNjFZ8fmIMRS9
7NmvlUfgjix02ARp404QCW/M1bWHK7030uIn02N9MENICj16z1xtjntTmsuWUkiw
uYsAOAkEbL666cdJ+9msMqhbfacKrkH15pCYqQFUEXoPGDpiNneJNTNh0jxHeXWu
021esXg9LJclq0WB1mot0P+r5cRQV9c6DmxclActAeUEfaiIRzmaEnXNAdEPsJcP
QUTDmNQzOGxVBByfQrmB3HOgvzSLUyWQ9UeKb6oTbT0DFX2Db014zXWm64QvFXW8
5cMEYb4/8mnYxQusYL31FSwlkxKlR6xL9Q6K09U14+40hjPCQh+8wT0cvWEoG6YK
DvrHGxW4RIdFJsyWX+Kt6pcljRzSQf+50lakZpjMcZiPuFgQVoqWVDjijD49utl7
E8YhUs82RZuRNa/I4QiJqa9KXQr+lC8Eu5GmIt/kyotlaQcMkxyjnMWx/6GbHUNB
aOcmYEq9oJKHMEj3+qMIiCn0LFAnTiqhKwYnTL7fmlcZ2PPX519juZ70+jGZUFVP
dUsn+k3D5/kWRIXWmbRrWZOUlcCQEYPSIEvP2AoVDlQfBL212i0glWRSahqogzr3
Ltzr5neb6Y5s2zxpXXADmf5ia/0DKDYfJEtniE/xRqInkyVPQPz/zHPzGKLcV0Qu
hKaHX5XVCOT2D9Ng7zfYTgtHOYHVXHwES3glnuqfg7GZFky/7ISC2qscLmNHyTPn
YhySt4VX7+qSZnH0uTBtjehzlvTWJqwSmg9Wf5335QcmErNeLCaRam7xUl5gqeRu
NVcJq8olvmIbK9U7mD6xc2twEp5fIphtGoEsSLBt9oQy4rFtnclOq48QTm6eOODe
7g6yCdAry9/mYSELAbEX3ocSWWShWDdqyFy7lAp0X4djynEtMd15rtqUF69O/Sur
GmK33yExuS2QoHk5fj8O/lZgx6hb1hjkkNIn/hEek+F+Eg2GNOQWZdNEt0NNg86m
b4QtBNfzVrOCFMF/9qwprUzs5Mgv9Z7aBOQ0yyOKElOykgoKyB89p2r/nNz4m5hI
dsillrIpOQI4McvG6VMXwuppGhkrGNFtiAdCDWrVl3OcPtTyMKl/WUOuBlo+5PbT
itG4tdosV1sG4xGOvk3s46TjmMVqcC0BZqowgtS27QT3ihWxIitY0iufpJqxOYhh
BPprf7WJGV1am181kb263IITbISg71jBMxJld2N1V6lNpxhRQsHHM+1LbZTSj6l0
SLvKjMGYrUlKgX4TOY6QiPFiIa7tylvkveW0q+FOY90wGPJPenvqgtc4uAWAHfw4
2r0wChQf2OvAK7ozS9Kv2C6pLvRkIvdWvtZ05tP+wp/Fo/HY1bH0+xRT4IMk93++
3pBCOmfL5hGejQM158gKeOIsHcsHWK1Wuf+sFqmIxrkdxxXzTrbQU2kWvTVXRlBN
hHS8iIazcKs5NHPGtSpC2p6Y1LDRFXIsZvSoiIl8zUYVjXReMVOb1toujBEiIP/9
MIz6PJZwy5xRb9PeVAgAcgVlCmSQQvTDAXX4ZI7AOcXCWhB3OfUNiM2knBUzA8Vj
941Y0jHnXLGdk39JvqHriYVJCu0DDyJELRvA0QzjtAwXW842B2lpRJTj/PQyMfjl
D1uGoSNtgzBMAuou5sPGnZnfamFYHc3xbSGuk/rpHoC3DlbqY0hhdPtJuOzhzd3r
N6VCuaby6pjI7/ANFHHyBaLEkGfevADNhv+pRrY/6J9D0Cy8oJUAC+5jLjtB+WPe
JS9xIZVVm9FaTNDZ3tSEEEK5Upt2g1okcQ8IiqfssW34OsQv/GPbDp5Dn+dIgMnL
EMV2Cfw54Xzo5qfDPZRkKRDaf7XIg0CMm1ntn5aoO5gWP9Sz4e3NrdWHmG15XmDP
1F/RLMOx4ODgzpamWgLMRWgtnb1ZzCdr9AEsanseD537j4l6jUPF2vn3fAu7s8sV
YQIy9lI0e5l9IOcr2TKtY9YoV1o0a69rWh4JU5HcCAMOP3rvz7pAfL2HpB0tWwdI
VvcuXC1hABzzCQm1zTCYF77dsCh0rp0H2LwCXy4eOYe+2eZ+WgZ51gX+cBsbw2WO
BKPNfS2P5mWYNMPhzchL05Z8klOL5ds7e4RzGr3i8PSS4tZUdWUWyKXXjn5RfE3+
tDFxW1OyvTTrH3AxrN6UD+D3vYBriryFFjA/qqP0n+o0ikd6Vw1M14uv2nG54Xg3
LWlYfi8CNsbUbno/vCR6QmhNLG2jzU30sXmlHQq02Aa6Q3GqK2FEi8JZx/5wCFuN
uDDB8OyWMHsOb6ucUIWNtRQitY4u1EJs/SnGKo7k5ZPvD1/YwsoAm3zspoLDX/y/
d4KeN6lsdvwWD+YlhQsq7INXyvOS4XJU/+Fki2DlhGBsP+fr2923MdUP/rwuf8hS
6CrzMq0EDz6UE96DMhosE7OpEps7+p9NjNNlcG6pR4glU1b+33XIHQGFIfc++hSf
aEIBf0hn6L1tZXoFPOqMmNVDHNn5oPX6/3ZBF7y9pguHmiSg71pbdAuzgMreGg2Y
CVZFIhJ8phBan63yk2cNsD5/3eH/xm7jgaii6Kk2XYleBLlBLFipPGkGgfakWNgx
jYxsEnVfZs0jHjtoMyyoH3ZZJZrNqlZXduA1vtbebiws8b0JiDSrz0xwrYNi2Uie
tkbH3B6fvy7QV0ZcN/F+DrNFOxAOxsgzaT6XtN+USUn1fBrBmYjh8dfRguyLCw+5
2CvZGsJ1ZapZBsAFoEIvNCA7RcSaWdAdtelZvwhUJY9CwrrlIjljGrINn4oyu4Z7
TBe6Mc6UBkTOPhdGhRh/44I6ORilMskxzCTMMiuZxou8LOuLJY9EIVVb9ExT6mOv
rUEO+ZKhQep/wJyrRf8VTdxqvxJFFKzfJVK4hKW5QsKAhYr9DdSfqRN/8sk62e/K
m/maYYRn+tOY0/+T6YQTI/k540DY7yZRa98N2mgjifWCVtWIGtAjZXgUunOG2cH+
44tOeD1bELCAW4qWW27dDib/YxOHIO0LpHmWBlfUDt5K63pAkIv6PN0AJOYTWXiw
LOjzwSaOUnpPD0JwUlKUbDSsEdZRasgM26YsTyBGTiDB532p/xrpmrhEH8ZKwPuE
pZ8ygSv6uiDTPIKIlupgLj3TK3l6yuhZ5V2cHxL1AoPsP0ASc3LKLch3LRSwJ4X0
Lfp0hmoT+KFPPBklrFh+6SCSetOcskBduWuqKbEtFpSrwaaRdUIA5+7dxPs8hHpX
cUGD2PxLFPhJToLf/ux3NjRkH6VMXs8sGi4eunqctF1ypFun/O971JtkZIgFhun3
XQRUqmqtyim5ogLjlK+4nio8Ddk9wJSheiLM8vvbDdb7iTqjo4XL7t2TxL2X/T8K
/qSd7r3gdOS2ruCva4G56tAJmCvI6b6ny8tX68psGWODn1sf3akuVbAhw+T+Ip5Y
KCf9oC9ymlOy8XdrYufMJ014sSwDWYZEpHXSDCYDIU5Ayv6+rnLjaRipdltWPifV
dR2dD8Ev0yOlRCuUD+Uf0Ab3UCIFGzIzINLU3GJ0Tx6Z8vprxQKQd+3bIVF7yc/P
cqu6DdJVZtlW/E3GjV+quMnWKqVDO5TzmOL+XHzAZm8rmLNFYf4I+1EXgrvCU1m6
nSyRbZGNOc0imkgmd0DpEoPtqMSV2uaQpRNqzr+SYlSY4VjwOXMTL4XArUEuhk03
tTxMzunifiHYJZAGmxGgA7GRNMtOagaQQRfa0rQDEEKjEFCxTfIT2NaSLAgVr8rq
RtqNLPiXhESFEDwkMDHL2YROAQNScSRkJODFB0GvFBBJA2EdfxTc5TqhrDrv1QU8
APvRHHxYCO6euO4W0KR/6UGEU+MvJuU+GMLopWE+P8jf6p7C56C3njX2pI2VGKn8
ILG8V5/WIb/H+vPdINmXJwjxLSj2trsTOwcZpJCF9KmLz6/2gbzX0fasejdTqNji
GePjoGk2/gVf7gC0UMd3XSDrqIQhQMYd3+w/Nkf0fZ2Kgcm/ojHvsUn+IuUZCnBb
8bzfdt/Y6PgW5pEEe6a2xw==
`protect END_PROTECTED
