`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n06rBZP/B7c0C+P/aI0QWWZyzbliO2iKDle7u5tmBizjOJRVI7cXFey+LIKEyZGf
sqBQ2LAmbM4hwgbGT2+xWCu0qnmsKojA5iEwVX7eAtcnGxeVSCHOz10VzuinIDYL
ZQaS9w+X+2ZLT49OXsgKXq74cH7xXL6apYNtSmWo44TEp5GACjdigKouMNKvTaCF
hoLoFD31t+lbgnU4v4+A6ctN5wQl4HNiO2uLWsF83+FiIgC3CwLbKWdB6hg6CUxF
utKyXOaIZLU6+aZvBQKtRfB783mcbJ5EnH+fUGP1CUM5YbqURIPEF8lXUAEds79m
WPYW5EQNM1EZg0zBXeXSp5u49LJTh2Ah3Zosl8Su2qYjlcNGs6c0d+UlCd8ZyC+t
5qwDja1euDoYH+OMrk6BfafRSMTblutfl5zUr4JZj6uaPfNkQwoVd84jgT6IRRl7
oeJQEWNdb97250my5hTep7SjrrwTL58Yb3AlZV9Kr/afIsizLPz3N0zIWPC2uSBx
UYlWgdoHijS35nWd1KVVPoYrebKZKepzcTeCm4HFG/b4LKUtU5JXwebibiOyERpL
btvbjewjN4wylS1FlgBGwCRYJAnrbBJbh43KChf+HKrIeXVMfxump1r2OXGYVx6X
11IyzAf39a/8Fa/NwruB9wJVWIU0kFdHM0cW/C0y95437oQqc20kSVaZsVEQl9MO
y2at4/FTRXpMx8YzZuOwOQ93Rv4ZDLFQDIiAzu04SaVjGxLQPSIQ6aeqgVoBhOGX
50418jfoOfo8VSbnvYUnnTGmMOtSUZs87Za4Y9f+5KEl356o+Xe2iY0QLDGoCSvM
LfCm4ILGg8zYiId68PVtLQwQ2KMJ9eau5oTwxYVmDktxd0/Zm1c0Ex/6tPsnlIqh
cs4w5gwUjQHtnQ4gNO9zparUwAxxNRS+VYW9H8qMfDSz492APVExRNlAsJx1yHTx
kYMfcHVvTP5m/sIvb5AWjVFpGDN5VjyS90Zgg3zElXxXkbWR615xsSAekNDmIynR
N10tPGW6+r6zZbDQ0abwfGVTJnXll9efOGZDGOca3Lp5iPhFlLPQ5UW/6bqQSyPS
oobm19sWwQrD8y+vR7HZqs/JowL0FD9j4mr3YDkPGAcW/2a+a88ZvPCUX8A1SXtS
Pm2Ru6/HKzSb9dkYMuQi3l3S2GoU4kZCXITuQFdZZO2dGtBMIBnnM/MbwF/q/qWD
UDHwMbjFFfLGIfdHdKz592fXryuwoAMIy51Q8hPVh5sn1CDqpCl50WFWdU+sqy0Z
eq84CqyoAHc50FqGhS+BqYqD+h4mCB1yNNOt/WODkbkLMG2qrbUt+ra+uiYf1OgJ
9icwbXgicr5zDUY4wZoBIj36oFJ5y4BuUlqRTW+sQYw9ObJsTRO96Jmc85dqlpnL
9AYZQKfaoC8UrTDTB6F98+H6jFcz+HFm/JJhzWEZXesAYnTA26u5wIB/61iVfVOK
z61qyJSYXoTwse1l84NowDL2lWu0YfS6yZ+nAjyFsxFbF7euvjycP92paJHm6/OM
h0IaBJLphm0JloLJMcDEpOP5UZNKpCzJi2Ey3ruU199VJFC/PVL7hwnWjN6mEMlZ
3etvyrQlnMs5Zi0t4NgAEGZDYI/HJmOk7N05wH6ZL4b7gjyJhXAyULriMJHzHlwh
DypUDRbRN26f1TdQGWbnc82xfaZEOvFZOjlrSILkQDfysWzZlPj06OIIIeirBzou
HlSLxUzSleEoAQdrsKaXmhhjqaZMpuTX1TO8rI5SMhYNQqT2VgABFkPkfzeiwbxM
63/B+OIRTpfiPYYED9mqy1uT+2h6Ro1+wQd1e93xrdCnwWaIllOvEPqJyf/tQpnt
SN/e8rgYEhwYtfBsFSdBPkTuKnRF7GZU8syApapaXD1NrCfQOq2aAzejtBNw3p1l
KImzoT0wBsWOxpFyn2BQ/8wGqk4q+oTbsWsFJV8pTiQ5udjopaAdDEP6XGesTp0L
a6oSxdiMF52p/XoSSD/ucM2nlqzzyJZ5TqcUm4IDyA9CH6GvTWAmShkSID79HGbs
RwUqHXJxgVNEgC7geaPWDT6nNHKpNZfvpzi528HlCtrzg1+ArFKU/y2BZ6azZ1PP
DYfft+CYbPsn5w6LGLRVPCJs4FBfP+p6sVsPfzUG2g/DDb+awnaxmZ3HyoVXHm86
Le6r7aEFC5B68obueGmqUnDkJBqamDRCeM5JIHWYhjIQQFo4iY7F/OQ+BHvZLQTb
r8hDx8hB1DbPL/5t8JVnQknQ2pEx+ACsheTn2BF/9DPsBr6/+eCyHGdabNTm/4Kw
hwNIRVwgWjETCtzib79mjGZ0VyQbotOdCXhQXqzScP5G1lw3UiF9cIZjd1Yewxnc
bsY/+RxqTRek4E4CnuIUx7Y1oWEJO34Y91xK8WBqaEjywaYJSq9kj8FHYbtSxrZl
4mq1zpvxC5gy+lFuVsSPXynm7IiZ0jtgDC1WHvG+ScyNeR6jrM7m714Yvd9B2bmf
DWpzLcPLy+KMuZ4/LANK2b6oj//fF7+4B4oLDDJ+SsZE2/oqbq587PscYCrUrMg7
qPym/eb0J7MBiS181U04Rh+DhJFQLXRPhkImfqNRGtuZGiRHhjZpG58rBZYUTb6J
qjwR0psNXPEmyEANZy5+LcnOUhks/DAMKV6RKXimpQ0CKJOklTw/siBLTqXNmwaw
mj9jBgU4lOrXnkYFA8BId1rFZ5Dr+zKWfIFDdpz+MnK2Nrf6KB8cwzSq3pyJQ1u9
tbfr9IEb8+MjhrEk00qd8gkX6OKY1JvZBQTTf9P34vXaQP1gYkMMxFVa4Vg3qhVD
myqdgeln1xjS9dkcGmGufa6oqVyIe1yGBNk4dT/YOIzTGKdI+Hr+rF/9ulkh7N64
o2o1XTzdYqW5O37l2WOSyD42itlxeGyb+2PaAtexmuT7i7sKYNGOiZqnBqBMVVlA
CyjOADXWrti34fdez8FmQxfZ9rkJq3+blsGXUynR3Lh+9nnVEs+h2JjuRhxRp4db
qKBju0Me1LCep7zK+J375KEmmG7or6bSK0w+q+ZqM1otk2jlOG6335eHi891QHb3
/4JH6IIy0wxmguPQGkZCu+0JPkWD9uLOZ4gWPhI6Dw/q59du0O9d05RVFUbbNMmW
t/+mA8dZC+dnan3PdoeaZPq816s913/hR3nG83pglT6xwE8yColxLy6O6kb6Dt3o
VTj8x+a1P88ljXx380MlDR8RP17bWNFg7z5Q+LgPF2m4UEQvheX7Nk6CHoLOWBuR
4s5i5MHrg2h4WFgvFWvPg0Gxk5vysg5iVOdD7y1v+7snyucXyJPGfx96wKUalwLA
Is+Ee5tyDfOED9JFSZe0ezVqWVb7qhpk8SsUBLl80ryg+k1uMNKrDkWVtEdootSm
qi30FI1qN98v7W/R9yZuMX5Up0jaexshFZKJOYhmoPgWRDbCPsoc7vwy9Xo5WtJ4
Qb8bqxfFwREql9jr0h6zjCr2vK/igj3nP9AcnsvPnRW0/aCyF4XKDxnNALRT4CcZ
GJWNxWikKLL0XQJgaGml6JzD+v/SfRvKpwrVL3iDmJy6UBx9nV6rPe/C4nkgi5MA
i5r6LCxNLpUAXkFTJ9Kdk0E5bcCZ9sXQjc88WD2p+wkY7qff/69X3/lf8szbI0Go
DaUKmIUFPhut8BaNbkkOvgR8ZYlkOfoawTz+iNDBIWROSGDfPsUmRpLqjmdyWULf
FnKfsY91lrDZ4ulfFywpGiIraDSAZ8og6hhxeFVYWU8VYaneUg5XhyybrLudieaJ
FHBTOFCBpFonzBPC6F1EXKMsE0WNa8fhq92Ofg1dQ5DYIiYKysjTnUpmqwXpRfZU
BZSxtbEtuVMMGddeJ8CZtIx6aeTJMAv8wCXYgAgkGX0cL5WMLH+XlyQVmdq01hOV
ir5gc7KIVtasCToSYmib9nO7VFmJi+SLksd5ZURbLdmSpKDHrNrrabxBl3J0rvwQ
vwdMOhX1et9whJGc1/KzY0GuwmSPmJWqbwgAQSZRUztmmz8wdZZTkUZFnSfRlYah
rB6Zn5hBZhDDbgCDub2kQbHwI7DNTtIEJHz03SZrzLXjWluwNwY5Zng/OdoS94eU
rHywvgbYoPi6rdT2NPt03WXGRUZqhN+C89D6oE0Ec+WwAsnEj0RvHWGNOK7ePOAX
vsYOGvjfvrIwlmVfXAttyOBRUABKvg+fKZ6qVlbsLAMXEBH14QyZ1+A9VT6elav9
bRFNH9TxcWrWKHy4N18gNGJBl+zHgx1RAnDy5ymdBWXxlFhoogSZafjkck/C6PiT
mAN9LjsRYxQyZy48UF2YCSE/siaR9mJaElJD4hxWm4LZgmzgh2X1KWrnqOrOsNv4
NX5df8sA9Emj/ALzEiMV7gSSIdvPDh6GEM6kqJQ9BfvibPfNPt93cc/hAZ5Dup2Q
ch9BT6nCvQp287/bLGjV1PEwaICg3pblbekhXTzMgpEw2OYqh9FEb/wLlvyjmihP
Hb0GELS8yov8y2w0bUWbOVzdDhW/tJJKGwSgIgM+SUzjB1pbOeGictYpJkE+aYa3
ju6blls5J5EYcSKEJONQW9AmrRXjlgN/e7zhaLEy/+nxfmavpbUI3wzRzfsHUSWX
Y0NRjJ+6/L6pa81yaCvuKwn7y17N0dy4XaL1IFfxt8Uyon6s6Rh6ktppaOWWfJBT
Ux0RKL+UWw09xW6UD6J2akYGMsZyGi7Yn1w4QbXwffP3vZVEHfzFiKP/CX/Z/3Tr
txx00gsBCwAC1QL0nlXJdPqLliMVfzAIczqwW99kVMMs8j2xHPwmeIXb+K+geEHX
ltN+rhlg8HaGQEOOmpzSNpJhblhL6nGxw1qNLzkft9nTiRBYAlqNGiNXI22y8NnJ
41Rb9K69PtME5AMWXF4teBx1N0HhvUoesGMdGhaQwg/XWKa6JyeZ9nbPD4JDvBbg
pYBfsX3mSi2N8K09MGtZ6bEjBTrMKxAfJGDZE4DFFltsUpPADnSwdsyYLEwt+kvg
3B54aZr293nvo3rZdYE5WPlSj6YQcsQPtIFkATXScYHpf777Vp2Vv8DLVRnC8coK
QH3BLNhGODNv/nOUYB+pQuZkOwG0J0HHq0yV2P84ugj62RmACpU8v8jVeUmkrNOz
wWruxV9ux/4QZ1fuU4AA5d3Zas8yICnqN5oC2aftoYQsznTk+7bu/unc0CZIwqWV
4Mo07JSGXP2lI+9OuxDCgzNmxfQ7QbIM47tPLdfW2ket1Y4JtWUPF3yKvimM6L8t
ScLpeG9gEhNQ374gqiipl/rANzbfWWXxpHg019aSp9DSPhWhab/w1OriPWqb6tkF
j1S1pq3kL3zJL+063Asn2/hGotKdNSKkxQh1GuVlbaNFR/0oBwiiN3GWLFOnzdWb
o8LFurp1+ds3UVeua6fVzMKm0Oy8prMoWSEv3JdphkKCI43pgHTS0yX12ZL1K/sd
ikNjd5/6Y5ERDNh9+ZTNlUBUHi/HC1Cyvm0YVfP3X+NBqdrcTgSUx+ZBA2LgAzZT
JjhXDDS/jvTkqZ0iGxFWrRa4r4JeAXYC/fsiDLJRAB5K2wqP+Yp6oq7eOb/GmGyi
QhTEM0usLLahh9KTVIlVov4fZ9Y7XnLJzh5P/C2v4xPJFogaTWk5WuXSFd/IONcu
jYG80wDuRcELf+ybUgfHhrgzrVduEGfSL1rRqF6PdrW4bjIO44YKtoY1DEeWBZ35
5SPkZdxN+77QTN0QJ/6U8gxFc5xy+0fF/OKRTKi6E5tvjVM5NWah6UsD9cyFEODh
jzsJJhjsuAQJGtQo+cITgibAzdI17PCGiBx/BshLGMIhVi8YK07qseaUxhatlfTI
DqelShi6L2rlOBRjwlmNayDfbaisl9Utum5Ox4gQOJDOtczlYqUz8m9nydl7LYX6
Q9ilCdv9F6PbDmKFJRr934bPPJzzAjXkLXH7E5HzuahFu21LPkLSyZ66J7t0L7Vb
Mu5b4Ng/xc+KhK1uA4qx3JTUSiNNNH54561MpIk5MXQL3sDDyx+JGFDXbAOyZyys
M4CiKt8OeI/SjQjQ1CFRDVpgYBp6X069ePt10hxQAQd0NECYpxlB6utkqhiwij2S
6lu4OW/7EEkkmW2A10+VMpzAy3Kfkhnb/6ugpJG25Hp/DqC+US70VpcqqQD9QpNY
Mc/oKjbkp3/uMUCAxE8WFyYZ+U6KMNi4iFp53ICXg4Vb+Tu4nrPJZcx7VD0hMReY
Oc4qicKENgbcNPsMRmmd5/CdzNaKI0F8EKlxwfBCHEdt0XUWfatI4P2Pfaal4Akf
RTExsetQk84JirNnnOdLBgo58LMHuYOtgIRpqd/zWMJjVPKV8/I78lQBTVY//aDi
mv+4JImPL6tFqk9Z7PY2am/qjVYk6fpiZ7wBTLQRrx92uTSKlo5UP+lIM2b0BA4C
CxtyO3zgT77wLL7k6XelIZC3b6JgZdOFJ7BDPd+MI+193wL2mOki6tJI4LT2YrdF
mWDyEKFt3Ky9vOVuJPjI8BeeRBr/0mcZve3rtl9gzejokLF6kjZdlld/7LCW0CYT
Y/0XK6eWmhwFRgEFTlC3PMqexQWDfzrAhJOWIdsmDIC0C4q+/Dp8R7E+z038NGyH
tdvP5gV+J8PRInYKvQQQDoeRAFd8WH+YFpOu+ZLuIkU=
`protect END_PROTECTED
