`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YrDoJxCYXsMSwJbmp78CJJFC4gyW6NJkrZagLJ8GWrFT9TKzR/Q8YOay7fNddwCs
KcQl890+R9OodWb0oryWFcVqU8Y/49xZcnFMCQlkh+6qfjbiiAgu6NAEYN/ciMVG
JyYpHgTnCbieI7hUGBZdZ1XEOjntCgzhsY6tNW8Rz5oThqCqpytzhPNF7AVftHhm
jgB6/ZEwNZvB2Cw9qXZ5JZJRXRc/dQS1PhPU5NDAUIMhf7omK/4Dxr4+lnLDfux/
0sltc8jopnu9bjuaH+LUZ7hmP+roG6+ziusIeSbL3abTvMQL6zsA+ZYPW6Hrvo4Q
aBlFt25XSpVHMfo/EIok9SEY/7wn7OW1uOocjAYbdUZc6otw6TBvbZ4LgqxaCQNw
VAXMx8uykvWS/WTMSCpPzehZvMIvYSNN1IH7vADIlHOwhDU9JBMUO/CpeUJkQClI
JdUeTkWniUH9G1MSIFr8AQDOq6YQxnIbXPlPhBXKhKscq4OeoQ6Scu6EfJ8v9P6v
lAU0HQ+HK5ezfRRYuaxrhqshOdWAb7zFsDaXhJqEDzz8iFZaVz/wkWTixGMHAdNs
Ats/OSFf75gX99AtAMsbO/2vL4bVlzw3zt0jWiejr2QEQbzxSEfvRAG4tqf4x46h
4drUDMyGjmArEhryH5Rnu6FmpeUMfuPiwI8zsGSp+hhsmycauO/5ND4g0353YXq3
kT9oL5YluAuV3xE9eETS8hEXyZ1EPGEmzNJ17jCq/rMdUW8u9hknyu+dltDzBWLb
P8vLoMCPqjPjGLy8NtlDg+F8RfufLRnYH2/y+TLJ3FxX9rn2KwFTUZgYgQFv4MWF
+OMkKu9vndrK9FBTjGxOHNLyeo3ky3ozaIL7WL3ym83uDM+/I5Hudl2HCihd0eg9
/zORh3l3O32gcQtvHbzc7dGcvzifefhRc7VTPyShINKwlWq/pRV+HF293dg4Oq3x
C1AM/ENNaMUq8/xXkIDO9D2depgf+TJu3FdetmZdBlvEkBqpbz5yEQlNhEDffKP5
e+9EmK7YV0zQB+TM4HtIYdxFGDTRSVF44o0gZH4VbTD9od69D2U4giEN38FypDJC
PfbM9vjfe4y7yzOYj468UVrIzDQRg5H1LpbkYHCKlJ+aSc80Ms1IEX5TKbKdW08X
dffzPsUbS7BstdCCF0uJleep46Sqdnolsy+CBOtnhEY=
`protect END_PROTECTED
