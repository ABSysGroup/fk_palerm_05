`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4hE9zjqaPLNDQO45SI1394mm9JoChVsL88+FzjZplegV92LY01XJqNn4fUPx79d4
M8QGPLEGAPmSJcOopxu+JFWfbe5vU0hPfkbUH4seJJvKRvpw8oGX15J1ynm1cUfe
WpXMwWLP1a/MgE92HU2rjgBYc++YhfIUZ6dHiH6pAEiGdbbB8u2GW+fPP2w0Dthv
ZQfFnv1Sk9DVwh8uYIJ6eRrO1BBnA3w8mB6F7YSkeyPxmce7vk/CRTs9dLetYL06
+ajOxyHGkJhTJvFspdbD0rxwU8nTxv0p3XqeQjgDiE/FfZ0j6ZjQxtu/qbfnvXlR
4kdK47JJTUpT6h75yz/WVlG+ZEDAWH7vnLVhSegX1Q+XzPQtvNd+9sSqKY0/IJn0
As6Nhqc/WXEeJGSSycDJpbWWUl+4UZ2P+grATBAyYrAbwy5w4AdIijvKx6soHaY1
e6jwWJZYItKrDtir5gwZpUzncGt7K8EAjBmCLu9PqPoohyEOMMhKRuBP6pKcs48p
G2qr7na5S2NZbROrgvsD4Xx1t1eObwOf1QbikR2HmeTUmO9vuGfA2++ggxgmw/Te
+9mYV9ej+TEh7f2z2yiJHWWdXCcwU94rSPUnBrwninqE2I3MFL118rBLBv18qPkP
IjsI8j+vP95TG6P3HcQEIWcch1YG6SHwJX4GR4IACxEarH7s1MLMd2Ng+fZECK0N
PgINYyO3MrQBehUM1WDhs/QxmtrZY+AFwtVaLugrmcAajcsTAtIS13NPTMPT60WC
s9rJ9kxOWR3LNOgARhYy8CrGwzWB7YbtLAwW49zpy/WeByuV8pOwZ3buduWc8db5
cje68nYtDZrpnZ4gl2cvd3beQ4NntmJ5AgSrV247PBjqnwwIhcX1De221JZAmQut
jO/93OsVS2y/+5NdMzA5G5QPp1C/N+L2ZMuTuLd9/NKF55Npc/tK9vODDfzifbGn
ocgz8GdjkZPxGT6Sg1leNDmreHyOT+Jhp8QTDZCWZH4DJH6WpHPFjRogshjrbD/g
W2hKpaDUQOkJnzsXRI9hNGjXqPV374mRtdOp38G3C3nDbNWB5pHhtjS8sdSN5xa1
SSj9+8kwaIgGKXghPSvX7lAV1SC6PZ1jMPbrNlR8ijKHzdbIi+LRrqp9AXmsfwwJ
rA1xMMwW7c7bsnv9Rs4UUSI1+mB4zxkTDa2J78TW/nh8p1/udyaUJS9z9dLsKLcn
9XV+a03dMFlFqotE6w7R4StS7ruI9+kWGdGHGwFYenuUD69VvKq999UEWBqO/UmY
k5gfcMeIR0/zuMw3l2DgvJkYdD47Ue/RPaU5Idu/LxMj3pEd2Ks2wP6yfLsfq6eQ
rNfKiDS8DHZ8yHnEhwmahSCDIqyrjXgdVO1Tn+/DN72JFSCAxEL8C3ViSgtGpL5q
5xDUZxhIkpfJPn2sq6EfBbUiWUXQXi8bwGMM8Eeyr1RFkAwjKiUXn+UNAScnj7qp
ks8NuD16oYkx28TQEQ+oXuKjWV7Xt865rU1I11QBLxzk7JLho3+OMm5Xrfpanc4B
RxeodATJIyyx1EgOAc2WoDMDyBnIPBdoMpR4pgpaXYktbdSjfQHkgzhPgsHKMPrr
JaTWhMW8Oq/yaxt9nd64bcZ1bnX5NBJjSfs5JEKPfWDxtceFxiyIdDBQ4gJZAU3y
7Exeq3njiyaIxFhUzyjYluN0CHJ+Z0ItVOtOk+z/lsXWF5wHEHZxC/O/THT+2gOM
EUybcvrwTNNKjyadT1P3jWynMgLEAsHagTDdhToKW3IgnczxWisZ7x09kb0NFTFG
Zik/hBkNFWmYtyZFz54vNOABZfteXXuTsYWLw3esIXia7LqVLwjPQS6ehSLVUheU
Qd45/Ax9geklLbwE8hp+JFBDTp1JrKq/NNTN4OzUeGAcyqcp8st0qZ3axnA6CowS
WaJiJLhetwWu77KJAXq8sT8wq7wYvMz0ibFqSEsibXQb9l3OURRrRAw6qn8Yq4Se
o/tzBZoQ+X1d8dKicmRC1KnaiR9QkMKfYD2DRHKrAUMKXOMF8TtZihwYGOXgwg67
xFaQ30oHcR5WzqKSRdAMjJ4NIrr8TyrkbObXQrPHY+dAi1Jr0Wcc9z2uePkPRJlm
CPKRo84QQPzzNCHdKGxvuS8anMA8B7QaU2swnc9eOHL+czP6HtxqQl6k5vnHarey
7O70m3wOhdEbl89ddEbjQK9i6yjSMT4JuKpVczG1v7lkJQb/Whdl9A60SdHsiV3F
S80ugIg1B1AWGgqrYQQBD9zBhqYaLxxmIZLtCOMkDC2XL8OTogLyv/8zQopyphtF
aJIGuC97k+BzFYjxVKYJtamlgqo4CyOQ59s5Zd+N+F7oe7u7vgJtstrDDDP3N2we
1f3LBoE6alT8MCDr7fWl8onsCOceeQX4CJx5urGfbHM8Eh+aH2eeMVfhmIgbj2f+
UoeFCucxj0f1oCcbmetNi1QkfK5FJz0WIR8s2TB3EjIUxu3IRoreeEkR84Q7Kp/K
TZ2HRwnGwtZBzz4G2nUuenrhxEVR1tC5EYzLHf4bmlSd85TxjzTyppqBlbmBicgh
IA86bSNCRpQq4o50zM424qJJ1uj3PKLO9dNc7qzrR+4XmKBvd+5L4ra39ZhhcEcW
5JB5dI9R4y2dxCxgxorsG9Pg2KWHyAwwKHEhgVf6ZlwpG6dMjmCfeshLH8bDYl/n
bCxmjTdYNBppMJCNUV5Fb8REFDVJ6TaAVPoTvP1VygIxIQGxAgiXzbnq6UaBviiG
GM1U8gH+vSrtheSZOc14j2jrFPb10T90BjAh44LB+jhxKi0mSH+aX/LwyK3BgwNq
c37frOETooa0LXpmyaHmdBCO8qI69+VKS4FC+rX6CM36h5YT/2u9d6lfweG3Vacl
WaGKcwdacO1THeqGKctWQRY/Jb5QEobKW3g7Kx5T76Pphc9JLxjFRu2cdFkSyl72
xA9LQE7Odkw5CXxOuosVCzIS20FQA08knON9ywBuUMfjXUFqRpRSAHABhCElV5ua
kDfoCQyPlC2lChN+B2GPfFRmbj0lQx/1RCRXKPYIzxFTHgRs4ys9r7BIpl/v4E4Z
4fQlDB4S8d+aMrUXsRDIbVDPeXpchJ75QJWOkMTQeb3zy/0X3wbbHyMgxrBWdddM
E5XN45ohfnHz85s5D4dceKNhGh9iXphPk1FC9o52md7zJSD4vIryyhS1njU5EFBB
qpGVcsOHMlB1gUjUBus5SK5BsToUdSE5W0TlGo4rAK+PH5z3xM2Y4OAs4iRpoTJU
wVx0zdx3Ih0FVQmGPGDo3UW6qjEE3swzbmT5Cal4HG6jGEz27e+vi3PropCe9onc
PDDpgn0n9DYpNl+J37oDTvZtwLV6hIqKR+T4GNWhWblWpLwIwwZCujFLWvBmo3oI
tyikT4zqP4iNPSmEIgAIa44H3LTHfKOmh3Fu5edbPk4xOeDh362VzGqsB/wU1Zhc
BE2QuWqv7OavUOcrP9aQgC8T4ycMoMkhI4/CGn+OTueFokAcmK+rWRF7BTOTfkvt
yPVBgKxZhV/SRHzS4NBJEb+FucpSjVyfmFAsD6KD8b4WjryWpDDE3EVCPYJqpkEM
JetD+M6dUsy3546GczbEym84bsdDiNJ9w5/ZuH/90yIkMSjnHA6E+nqqh8as6x42
giJaOd+1SengxNbcnjN994Mgwu7JdpOI+2OwtRIl6wxIUJMBU8AKQPHoj6YRnW9c
UJu0Efp0iy7eVifr+6/5WQMfhXgQ9yn4YiPcWJEvf2vtzi6YOq1rBOdvnC85dFYQ
50zufVdV5BwUBA0BMS6432ulhLW0ivp72SvsJA0ClYymSQyvvlEtjMc5vmbtvz25
48sPScDndOCfvfN0Sc0Oa2p750KRoYy9IG6ldUHrzzRUZOSlDGHfMkluoPC/Nkix
rt2WpcudN1fwdX/m4Qe0LRHFbLimVT0Dk0j8oybgOkpAcIJ9yJfODxxwGNwyfkt4
uQ+NXJx2wORfRF59NcsQAX33+qDTUHkIAgQOoZPICes7jTlA5QeCXx6dZguj0OJk
C+2gCaBMH4LqMpL7CNs8377y6d0v5rxA5ErI/6XYfG9/WVfzbhJLfnP1IeJ1pPMH
tqZ1dREOvOMHDWnGnZXam+0Stq4gHACVTquiWdeTMJJmVM/6Igie5nloNgb4KxUl
`protect END_PROTECTED
