`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F3aNP6rqs1WLXhNfULG4i1LuK1L5iX06LKSM546NxzoQ28djRL+/3BTtYHgIrpA4
y4zJHjg+eIYLwK005cCwgibNbIfUw0+ZdVR4eNGRxNCqLawobTQgyd6IFyxisDpK
H9R11jrXobZBlsrjpW4GHpLh3MN3GhR+6BJwVm72FArFpVbk6fb8bYKkxpmZCXfc
45z4QYxZo4RSxaT8Q39XbndvAb3wzhYrXQ+3ODA+XsuJPtJGN8OmsaujcdCuYepP
Jvv9boCXmjRCiXILqSoUAg9gMQ10zIoObuLs7ForSRRz6ifWMcvCSqs8+8RIw0uI
cP4FPHY1q8JQhoHnJmxGwB4qq2eUZV5gNpkcraPpvkeMwqAFySvuctfw00zQKxfQ
e+eSoG1aiRYcaM50+BM9TYgJv+Ec5u7L1efvPi7IBlSIrp7B7fOi71z99aUIib/q
OqfeS751879tZ9ZkGTbVIYAHbe7LwzoPNkV6o37Eic2kGd2YSIoZd/HvjgL5nvX/
qt+tUIWsuoLtAPJ2waFv3VE9ai5qdTUq0upm4TSw1F2f2o0yqcvqY6EXjE2oOU5C
c0If3oF9tkWIeVxK97uyROh99y12Zsr/T212BNg8Nv8QmbNpm8/x71HHAw6HZG8x
JXbp+18JXfgwcOPxDv6VIJF4om6DKUJNKg7CrO1IZcviKD7wsi7rkehtt9TgVX2B
mKcZrjhEEFafb79ifCvb/l9w91+kqa0mya20Lhks6M63ykVis+rRij0lYejF1nuK
TlUf84d4s0bGvDZNOEO0JyKnRRUMydF0Nde/AIdBzAYOrcK/wyx89cIdsyvKX0Jc
z5cpONIub1dva2YKdMSMVnY+J00SXaMIuKsMsAhSZ3eSq2qF/MlVIovYNpzX6CQ4
RwtbuR3b+IkEWgVA9cmbolCuM4WaSaRaxtPK29hlxgyF3fQVGq+sg538ZQwnxypr
ArK8t87DOQv6McTAzFJ8TDyPks94Ku+Wb9xJ/bdCXq/Hz6Xma2bzj4VOto5cJVLn
LZTZyzzMLgT6KBDrzRmdeyFb0utMws8SxF1zm4DwjWgjEJge+q3mbTBs6QwB8rTy
KVQzHvID3NqRDLun1NeHV719JtGEo1V73KkYxHxIIWx1JubP3ylRvN0vNt7PQFGF
QAVtWzV/IhZxVb42UeFu0uT3bVwb/mJJ+Yrqiqv/76+eu2EqFpPMDKIUy5dx+fI8
xzNUhDUEsUO5SCiHgw0l7gFXqiuI64I1wrVyqvebUQoPUioFjiLcL1kuWbKFD6Rp
GIlusP49TxZ3vTpDrb7Rn0QSdcn+s66ysce7cuJFxMoxTTKNIGdbsQ1ZX4GBgzvv
TYzsfeR1RzVhpZWuCecTTVvpj1dXEINsUjUQfFxyFtE8VWmnDm3gUDLgGDosBuJm
3fA+RSQsTmdOYzdwUFRD9BNX1ujK9Gb08PwRtUgnnASB2YfaX0RGyB+IRu4ZlUiW
bu2QjfSHfIPjJRbpgn6Y91jrVrwDY2ibv4Zrg1SBkgmXTXK4029LAtnST5ym+ahu
H7eO87IsCpmqONrLFGTHFhdf3/EjpI4EuHsOudRXqH2Epo1HNpo53nEYmzQeHOrm
J0aU3YYZ2ilNo2Wz528YfojjiQdE2sr1VhCD0ojufhY/mugl5YkJG+3uzbdAABt0
oFntM05SkaHUduAyey4jPqBBvNpSHGepq9zuvZrKhZX+Pd/VBYKZArkyLiwBeFqE
t8ouH1H3hAo39m1KLCYwFkFo8iXbmRpT6IEuZBGTmT46G09mySrJkwVBEZsIOVd1
lKAydaODjO3ua5QWIZ8DEK6TI7LgArALg4xvuQYvwTPEtucXnYNEnx3yewABLVnL
Jz0gbthdzhiTIpcBVy42cMwSdrTFzUn+W9PfISf6a1SDjQDLayJRErXg9Bge932W
Ee6tyqQSDFA2/DgIzLEMw+u/oX47LtU8ATWxiXOTAqijMooC/g+9cXEKdo9NSrDA
WvX4WLwZPfFy+V9LRP3l9weeKRe+36QEig06K0epENhuFdlLx3LOzr0Y8qTY66GP
L7Q9ObN2PmJpTuYxilEaXcuYsKHNzEO7PkEvjxwTjrmL4uLoT7OXRQOXajvbZKhQ
N1sv93K50j7IoPMQyptgHRGCuqRH/1RIwsheq6qr4cnFIXoSrAgZ79jg7Z7autH+
oQ/qCFpWbdsUAAjdxFK9nhLiMdm5Y2EIcsfqLgzuWHNbbBd1Bl+armXzMZXsKI6y
R2EJuFUgtkFnqOxdp6FDw1lZA1EWwrLSmryAGFnEPXfaEsubMzlDOg2zY+HOgYye
IVj5Ru0A/k2zTXxaqbYHYNFdog9Il9cUMFKWDl+vuaUoZTEpZKnMHrTt/IbU3lYW
lR83zO/Qxcy1BolKSdWwz64Dg80e+0RjM2n6XTJOFaiVPn8E7J00gy9rTZpO4lJR
Mu3b7Y1t/SayaWsecy0ZeEuInMWdNZ0oE2NBbIEuuXb12j6K1Gbn+yoZ18lMxPLc
utROoKGgoxV3EUWZ4aLfgmqkfr6PVqJ5+gEI+spz2iJXaeV6CO4DRqEcF//nd1os
PTHUoAvHFTBtn1B5KpExMIzUl7htv6XsACrwsJXtIyPqqWqaGqaU/J7FiZk3whxd
lX94Blz0dz+EWWUVZVaIKy+jUC7bGleegEj61BP4y4wOjDBPQ5n/es4FA2Ovdwmt
2GTmkzntVZZBtv425Ly7kSSzMSyNEnicMpFulSbuwQ7BGcWi7KUu6mjh9Kjgnvuc
ZHBzeJgyf6z51lIVVcGd3m/NMabzSmR46OvcFFh0UW4DijgMwLtAMxTr72PCNPqU
JIahBqIosgaV3akBlMg+dlPO1ZntFcJuspaZvoun1+J8nJg6XmREVQP5ymOCHyFJ
yh2UMwYmTqfBBnXXW6RDkabCqMRIdkC0Y9oSgKPoRnj0nMBnqcnE4wv3UccfCOXx
Onl8C8+Oaea8XnRxBrf49J6knsWTx6i4ndJvam34VvR2TQP6LeHelJHfFKVn3ll4
A3i0s1n+fA4jVqJ6Hu20d1ZZZEYSskYX/LpYOMYdN+2eaJ+28qgFFiQxwIf0MFiF
SJ/kkY05pUkzVMWvQspbD/3gAhiNWFgx9UxkbQzcpetPH9D/s0gLVPkr5eK2Kvtd
czUG2oi+WK/z5unPu3WNyH9/p85MnZelugKKhtZ+Cu7NO/hL0i9XcVGzNM70spE9
sQzdg7w10wIGS6acA28No8sL/iddHCrKePfTVeQkSKW9mVqNWvNbT2KZ9EQ4fyUR
7t0JAfzPsX1WNwkMsA84h5n6so8Jq96ZtADxzC3ke39FhTi7uUkTSWKhF6aFty8P
Omf7qUkpJgYgeJd5lZbTPF7dCm64G5W7AQ/8J5uR1nd7IKZ0Pc+rpTmNANlGZSgk
mlL+hs7Uz0NabPqBGoO4nDvLjwTkQ1DFKuCqBSzfGf7t7jDZphVaCIterx9cCd/e
Tm21daIE3VWoHnLzYRYJ4NLeMP7271fjZQdaxL8anFeGfPiWa6+MayV98MqbT/hI
RZZP4svTxdpdtPqVMIPzHpr/YPE4GwtjObpxmD1eC1/8eSS9gVw56xuTAJ0I2vML
SL10oo0RXCI2+gIccZqrBVizsI76DfEnrSlFEq/HA5hfWbn0sbWRYEdgXBo2bynE
h+jWFonYPJT44LIb5Ce2FaQ4Fwib4aSDdP3gjQ+gvBIaP/wKdyh8DHmLB9AEQllN
97zyklPmC43YKNfSLVAZ8ctJlHK9uRkjvwmVUnIXkjwDVjd4B52UKaNBnVIS+N0f
2ffjY8VP1VGiCxRNfZyKcL2ihnIjbLDmSJhTT9Ok71lNuRr9mECIKE705L1ZRnq6
fck2ALAer2TnwtgtWvleH7GQOS8rZK9m4Sz2gO85pxJ1O+O6HT5pQQ//eiOPxJOY
RYHwu1quyou/zTmgbFwhvIHt/0woyNS5E/LENni8b/vPcU2cAlqxbDR0iInON2CN
6KvL85iKm5U2PAhHQryzajJqjTbAiKb4ZTQ862BgE5GF2nhduiHJlH3kljkoHTil
Nboud96zq6nEKSct+UpJb7rjeoAV6ZRuiFctCRyYWwmmIdqwNytU5S8Ho2lzmiZf
y5E3LkieAbrI07YBocLFhoIigCDQOu7Q6q0uh7zmq6QvNIiY7x5tmH8fA8pMur41
ZeGV9vLLN42DY9UTFjRcy8RP71PERXM8O/I5TMIRFFj3q1WxZJ2ymMLTJ6/upjGE
V2oPSv0za7sQAA6+v9zN6KmcuUWK83IxGraI+yXFqvx1W8HS93oLnUGFeP/kkGC8
lXJ0n6hJnexfscBj37tDUfIm2A2l901gvrmzvyju2cpcNE1AosEuZfIWv0Vaa0xM
IIpoBpsUkc7coyGNc+KT9pKGGGIL200gf/176ejL+GKRZjK8P6ic7KCST6Bcu4ph
BcitNemcW7gmBs3ktdO5lfYbReUHcpUGgV0LctbmJFBPXZYJiB9I3f0O1WKU9b5h
ybv4VebsiKJY1NnLLi4WDcidZBn4T7U7gnEs5mddwyTr1FReFnVGXjMx25Hee8th
p6Ge5zoufQ6ZXh5YiA7FTtdRXUGBNGSM4k99/hZXh17ckvfr6FHhCNI/Cqpdp0zq
MJczQzCehZHfhscyfCbiB92gfkyu6a2vLr1TYBAf6qXrdUiIKh/DGC5qAZHijdQm
PuBd9bUsc4Fly3YQZ55huyYgC1zIU/s4V5q4jGPgRkQM0GVYFsVUP2UQ4bdxdHJ+
47h6q2XyamZbcv05r2wIARt56dBpvAlUX2V1auuUEs2WhPbsg1S5iCbZ6qst/MLV
1OR44J9eT+JOG3l3yZh2wxKoE8jBDrGVAepvKG03AgtctzywhU85pW4vuCOhJ4KZ
yt3w57Es7HfAMxonh6SJa+5rBGybEBAFN1lXKvo61EigEBWZSEDi3lp/Jx9rNmpH
1w2MqoMY9E+KWz0qvBH7Zc7Vwl+PqRn+oYLq6/JRk+S2YCR2WFs2f5z/WEYMISYw
mNP5COydNUrbgj5dzJ0WEvYgNlcpIWKd7gs6brBt2DmiQS0QfzsRZu9KN1G1l7SW
MPZBJUEzpszVmnLOpkyQA3NpOy0SB/TRrxLMENWiZBGw3pQdK0Av5AAO9aFHD1tt
JNJ5awsB+Zxj0E5KZZLoLg9iy5V6tLr2oQOVngrNNzL/ZS4MNLSl0leW1eiHra9/
FulaabJK/ua0DKwYUWkY2nUTnk+lzBJ5fqUMrdyXF01nm9ozzMzNuQFK1as10zI8
w5H544cAzSVyMCyx3Hbqkv8wiyAqHUad4dlSuEObkuWhODzZW1YYXUjn3mOnqkPF
PJWcCCvXfZb0x1MWY0/M/55+GjzaT9z9lM1zXFzy1UW5xT68D+ahTMDdFOa5XYKL
HDazLs7R0NwWqyNZPrtVq4Lxd7VMSzKsXHM81MxcpM+RqXZJqrayRXU9CTyexhcI
4m67KyaBGUEn2HSygd7UwEUJg5QGiCoKjt85xi/gx3GRomzDxUmHBi7tx0/NMLbB
scKxsTi2X8IAba+XSeOBZoAP/cIHFepLi0h49NdoP/XA07sS4uK3+b/q7mdjlaTH
OKtayGEe4NuErckbywQjjoKI0U0bNyNMZfLWu6txVhOzO4kU0mZDjI/XOZtmEx14
gFTj50vvBQa5g39O8jlgFLq6zO9Cjrt2UqGM6QX6rkAww6RS9GN+uiupvnC8fAvK
ehxNOLO6H60Yw8MZBYt0MW2V7u2Zkty2ZApNdfOROTkXJS83gvGWAgijSZrKThnG
WBml3vJNvKvUgrLo6+/bFA80Vz9PDibJyHGxQoSxC93VklF/J9/Yu4Z3KHR/hDOl
Ryg3vOnX7IdXqvI1tTmi+ZHVzhsjoGrseJyAF7gfm/21ATqMvCDwhEMp2nFYASbQ
8CfenFaaKGbXP4GYIh4moZ8IY7cBlsjhkNFA26sQYDLSazEvvWIzMR9SUFTgbNkZ
/9nFVW9Q0t0ZgDxsrd6aO6K/SUC1ON+w/betiecwijnetMXR3p64Fv2B5WYva7gS
PmALKNuM02rR2d9Ken4uT9fMos68MedJkP2XnQF5h4h6OCuWL4uffytW+z5pdZAB
s2EhcOnHQVA14+4aGpD3KuCTtS9Ok6Ob5yFsDt3c/tY2wxaOUkVpE14x5rGnXHPY
vaulyaWdNYVslutXasmzQlEhuB4ORI/APOcbLl1k/sBp1ktRQX60AhHP2dFvH5ty
Y77jmmY9cElnZFQg3La55perqagbR/iMUqcUeo2Mofe6bDezk12jfDkv8mEu7z8T
+EsdrWxAKsrmZnFVA/mwL2g9O/mxDtWb0M4JL9h+X0ZqJGnNhQQubhrLz9vtvKZb
zGN6xjDOLdpJ9geMfnCTtJt4mvVAC5iAUmKfk9cV6NP1T3pEt8pu0lYuOfks9Up5
IV2YXFnJzeqgud2bu/cQlJyDtC0tbqBljzSZU3RUjPiHi/jOfpgi8hWn5hWugFrI
TeFKplJj2COo+L6swL3IVqpDfr+/Ms4924DmOM6sgHEXXLXqXcxQLGWQ0LqdTa1C
r79u5oxxY9BK3PTSfJHUdJe6m2Cmn4zq6KWZOxcUk6MpnxuyLdMNRwPsb/g94wUq
RNpVWivYFyeHXhO4dxkpt/4kLyFDPw71ZpcmKQYOGqPWHJH0GmkyY12+cM/iSN95
OqI6vxwrxCFrvycnHj8I1Wl3UbRlLi8INW8QeYzzRETkf9fmDPv/jJ4tk8f3yI+T
7TreFIlZ3ZBVVNKCGnv4RD7fB7vDbyPC/UFoYbMjy8rZcsD6PM8hPibDn8tmCD+4
YyO/CsnAZcOa+XQK0E8jpiTCuH3cm22oaLFGQNRyyn7NG+Y3rdvZaykMW1LivYwJ
gKn9UaPM0YK/eair7gZHeGqODfgAZgQpor5xWqxWE7ek2agzjfMvXbTOP5Ze4RIZ
1IfEQCvIh1FCSud7VG+8Lhrq04xLYvhdbwsL6zXSuKVS1/N5LIn7jD3QKcOOD0aY
t+PgGDEoQ1bvo8T2zgBl/L/VS1I/PK0hgaTKIf2Xyqij3vB8beMUsH4oq4cG+cyv
KhaNhS5ED0lMJDRNcyzV0tevSj3SWALp9kWz9jejNudF/SUNXIVTX8n3ryu59JbB
tsG0QSpTdofetPnW8FPNQRZSBr4NmbLMME/dp/jXZxEvew6hu2mPOwjQuOKJvUCW
aFCT3gpiQcCjqiPLzSsSqBTn4WPP8Z7AKe3Cc5MSzM9fL77n9SvSWVcekV8hFzfY
GYbrmhva82F+8Sah8bAeCx9NTUrOt5XoUm6gdjSAQud3Xw2abZ/j3tQmPFerboLG
2TZNwVwgonbv4qQHUpycqcu9FzVH/r9l3vbrIipZK2x9SrcrvNrp3vq7OsFi8nwn
z+x3vRNSAjxuPEMCtvVA8MHAZM8NOveAMrgP84dSB+eMD+6fyLymCJVpeGL6XSnO
jMNsrHNN9sGtR5+Pd37R5xTBA5ISo+QvNCNcCAQruHHeFkb9B+CulqyYgnrRlPqC
9Zvu/Yyyp0pNJuZftJg2i07KMCHRjX5rYBQEhQBBjth6hRd5TkJBwPSv4s/YBftX
MjXG8PiLDoW6DOCirViz7DXDjGgADJg4CMlbKha37dyyCkIqaOq+tXVMKoulkk9M
eQ5k0wI5ETbrlm28rG8TXah0gBnnBzRsDKeVeFKWSqN8OSxN1poBb5MZfx17T7xf
qIB6xxMxbsWrRnwfIvdfl8oiZT9PVUkCEoHoBzjXxoCWHdmdTnB+sVj9Z4utb9mQ
MnbdjM/Wnh+aBruNKNvnoNloZu3u50Lz1IywZydwmy+IBR3thxO0W7oNHGfjb5N1
/boLiZ4SSiR5fwtczo90vGuFFGsllVESejb1k/aTAtTwe+9qgBkr7otG0frucCds
YHn3Q+8ozwbLn8pYudKRsYWGlto+Po3b/m2sCx+PqC27Ya2bzp7h3fiF63tl74Pq
isB8FCKrbXt3Ed5NApwaF+qsvb3gybLX1qw3qcDHL5tj5FoyUaRA5bf7/bR7FTSK
dHT9nmtHd+XjU3pSzNIWbpQ63K0oWUd8OgfUI2rjZ1MRDLUaq7UpefWzheG7gRMR
0LC5FO9pimS0pr/UBWkyZTikdTweLoPN5z5/6QOMNsVSw7gGK+zE4OaYp+qSuOO7
agRQrQDBFzcwEhjmBcU+FKUgENfe0U5/ibAvzigRag+9nOxyDR7dwwiAK63JiFwn
/ihSiN9syYz0F09SEUEbrlItF6fqicDmy7tAnFdpPKiknT5kxsapiRRDPxGa4c4w
fcwy4hR7na+ge6ilsKEtJ4RO9pPGWg7W0vt+0MO9adnRx8MEG7C6U8mRO8F5N31/
P8NfTjlKD6+sEhMivixDm3CFdG3Ykm/nd1u0bgtxTwAT/geNze7fqX/7DQyUW7YR
7pGKTk6M9LD/UuX2Xlq/r4mXLHaLEFO9tCnTyF1gIgYVT2w3EbfHR+oWhaUsKnfl
T36allmmZ8a56jJ4gpFf1l3qzXKw+Wqpu/UI/HQ9NtdmyPLb9ektd1ma7RlVQEKi
5j+A2mZD+vx9HbwxesiyT9iuIm5KCbUL1AwFOCrJUvdU8UBBMdrbOlOnzXLVft6n
zvQGQykovEdGI/JVEC4ceUJMxV4A5QyhvJka2ArlhPeSK31H/OBaOkFQ2w84ZLfm
MbnidOLEGx6A/BGwMRnZ4Z0UiMAeq/GxmOkDA35LIAdSwF8TjBFoSe06IqA8/fB+
ni8MwLBLvrPKYSANd1MQT3mIhfLPc70o6kncGHSbmmCcjtpS4yOh7sZf7QOX5Feu
iD9DI3CS0W414L3UcaqL99oOMRUTiR8VfTpAj9/gXDD2soTC0kPdfDjUfNk2CS+Y
nziga6697PGMD1BUixAHo2pEZKTG/jhqaEMoYpzGizqdKxtnQ/ZkWF3loOU1hV5i
oftMAP5GVINMBnkDtK/eVe7os5pL5e8Sy3cY9h7H4htE6Vw27z9Qm2/oCJLerEY/
DyTrWLkalfdS4PqBB9ZF/JXOeA+p3sSC6r98V6+ifYpse2lVz38Cv4hEUQv8f8bE
F++0LZK1otQoxryMqPdq6pbj2juDocvXJM378fWBFFT+0qtie/4pbfaggjR8NLBc
xMuSY/srU1XNUNySvzN/BbBj+ow89OgLK5mj1lnl3x941vWmnupJ09QMvQUlRHSN
4UnifQFHsfjunyZmcUA3jR3wNIZtTJL3bjIrED+cIB9oLmxXqd0w4LGabinj1kF2
WNhtFa6Tm1IO+dIEGr7cRQnvVRpQtBPMzZRtuklI1+PUV+yQ4BXS/jf9Zs0i3hZI
a9C/vVuPxxMJ5TpV1SmNsGNk69HQuNJCjlzyD10GUo8eLY/vwwQ+GUsA1uDX3l9w
gefhpJceK/7miYwnOIA0e1YYI0E7OFxukrytj6uR1+iyDttCGO3XhZwY7c/spkIG
1p0Rv4UM0lHgHfiw9u0+C2RcXfqxq3OJZAwKLxHw9+O+t+ftg5I2o0XYOwD40s2e
IV1Y4V/Ie5ekF6RkoqHOsg2Mi9Ou6kqZPpO2Ym1CRk179kDxTPx+5tzQSodof6Ot
nvTej2YeiMky7Bl3TyXL3WfDPv1mbINxT4JauJSI30ZdIs8j8CZ2XlGx0IXUMOyz
9yjmNT7/ffyMF25Gej2RkpUPeGqMzVN02pC6qPfmjIP6YE2bnlo2yTAb6qspgdMn
l/VlKnIoX6ObFrPcviBzBn1yMLlp49l/Juus9CRUgsfQkrUShxWwfEAuh94ytt0i
qKFUxRwKUa+my+CC3nG9mO3Sbac/nZl1+IACnheK83MAP7TbhdvKYZofjnwhlQ2A
qxexoadndLe/Z0NQnyLkPxaGZ5zi3F2aRXdJs1KlqiAlTzckC0ucgT8b9KeTCf9Z
P3zxaweebUW/L+qU4F01t12D7Fo0rvbJqRyuFWTXRbs8OGzYSUnt5c94ERNLxF0L
mf8Pxcld2PpYAqkRcAK/4WqJ/aeEn0CM1Gu3WACjodUxbORxOFdBxZBJEOLBQfpI
iZXnA1nSEjoqAfUCbcW+njho1WwtjO0LMIC3MEerOuAMLmC2LN5tJ6D59yvNkrwN
gf1jDiDsZ5SwNvKwjkUE2j0VP9yIgJQiEpiuaGrpJYCb7RQpIGlWDCu/O/BTkrqQ
ru6IBemdvaab6Smceqhp7L39e/WzDctMekNMYXUXwE42EO7ymLT8i6cqR2J01PZv
p3n1E5ee2bMHgTuxo9C2i7oEqpv45jWrJCNIBf/3drl3QDvYZY031WUCOt7ukLZ+
M4tcVJk1GEmnwuvA3BYl9T8X57gY5+ihjTAv/iehN0SlUEFG9w9PelmIJMTATLjD
Yw/DB1fMAOjL5gtQIRTSMxLTrtSahLTn1msq7EWrKpeVgCtMNtL2dAwQdFNtz4mN
b2d7DCw2pFXBFVQZOKnXHmSTHrcAMq75K+CZxP+Kt+X/zohZCc0WEDiO+5AMo4+K
riNRsRSC9Z29yoIvS+28VY9McSXlLhO2V+1h8pLmJOIMH7UjFbYfRRr8WJjGZw+R
r5PQmDkgIrb13y9qz7RjyEJEtHSNWFr5CH/2FPXAhdOyMsU1DT9IQk2maIKtZFkn
QgZ8Efdfhd+XWHn1yTwWzmj4lLlE/wh5ycIFAc5IhFkS+7EB6ioRn6jPnBPftOwH
EXwj6pEVVZMJCJQxRS1z8Z/XaMlr+OIlFNJpC5WFt5CLo4YJjFF/pxduk8hGpMIN
uWdKlIfHeqDRapP7WHeHLgIFPcfZ7Oo2pMmyakYC8DffV1tldK2nD0S0XUVJ8vO5
9vv9sk5+QbsLcuQf2vuc5BWZBpBtMycxvlo1gIQBPX5NMLl26mOUOjZ1/0a+Wzvp
3bz0bX0A6q09Q+JPh6V9NcMAFlXljRGHbjLi989MTvzrun+tNEqr1jiX7zl5a3ei
O/mFVWkNT0A2S5J5y5TftHdkCY3j8aSGZTP7Q8CtNxTz4CME0iwGcKYhEOoK291c
FNRqUf9DydGhQpL89yWgQWQTymVl7btLH/S6g1fby3KFaaQHSYcaYRxK5dU28PAx
7N3JVNTh5AK8tPfkN6pHO4JXdHjFZ7n+ZkkyjZvXIQsJInvseFJ4eF6N2S0VRm8A
0BMvsEfeM+sSuX5POnOzjGu7JOYaF1vDU+IpO2sFE756ZFYTDTEXs4fvWO+X6Upq
oR1zwq/5KeGtJkTGfT+KO//xT7sCOv+HqA0pO9cSLyloQq6pxbxhT8DQa5nbJw6w
2BC6vvAJjSKPpeRxa4yNeQfwRhbbKGL3Uid8C+v6gJt2xJsPvy6aDuxmWEZQ4uww
RCHMoDDGo5HsVUGIJXYsXqoBDhOuSttjubMGdvxNhPktI49tEVO4brg3JTMEhRu3
ZQc8mupvwHmLrnYqeqfCcwnPuDkJESbvKc6IX5hUqLkTYY/wLPpn+l4FIVAxCtQa
k5dWBmWMWxrM5W23IehOskJqXEtnfPxNcmdU40dlSE6g+kvAK/DxXVFcNHptJtiC
DZKW0drMezHRz199ccKpsx7mubIAXeBd5kKpvpDnNfkUvUbhmUOzCkx5DKKmlvON
70/2kXIsN4L8MJWBg3ziBWtyT5YZ6/AeM+FrSwaTa9pE3IDfiBEiAx6+43t/guL8
QytEdJff8a9+hx+bcWg+HhHRmmix0g2lfD/wa2g/4FeBEmcLVYkAil8CGCjhK2nb
oDdTcxL0ESHuxE0NJDXEk7HAkpMJEVUitPnqlZJTM79RXHlWzHgjgK+Qk0/qXDrS
hG8wyVcJ2jQYpyHhZoLeO2i6QG5D8NEmylCUSJRFPw3mNQevi0pf6lmw8LFzvD7l
bACw52tJZcRUT1UUrIvCm7SrHABAaz29z0MRtLjNBZwywvfOtJl6KoIkfn+dpvaY
M9iy/8q0EzUaRLlpJQOOPHGB9GN9ArkfqjrTp9f3o3VKO7JYrpvCWTTfqn4nGaaj
6R+K7PvSw7w21IVVi52qryi5BpMw9/5lmx9PBZJVp2Jo9oCsSJHV8tv6DlueicY/
1r6I1LD0j0xx19khdK6+DRHPVjNbs80X4yzDWKRrbis82sLrELrwEzMUaofeg+pf
c3WBpB9ixX8QU2fCOb7hZbVVfohmK3ppytKL55361k+e/mzMZm69fMzhnIfe4zOl
tOGIApf9hBHpduUERvyuIeUjmVLxaTiS0zL5JQ+vCCfs9SQ/LMroJs8YXDHpn0vD
5sgOrUsRkfnOtRoc1NAenrHgTMwAC8Cr1yaILvGMyLZsrXAn1eqDmVJ0q95CV2fj
U+0+9fBzWiU76Bwf1A2+rFjQKPzHb6U+b3cpZsUbiaIKM7lLyDCH0DrKiMFFkz6z
vmjDdwKzQMTvkkZjpmU+dAnGWf214IOPAc9OkSLYRxcDFxFJfTpHOEPRZDhqIgFM
JY/jZuWSNrVdy7r3g7qPwoPQHruev4qIBBaWwikHJK3s5ny85tVG+Hc5gmQrdtK3
3v1uY2uvB/+xFZccUuQfwa6xQ3KIlVlhGrc5CWOXK+UvTpK4NYdi6wDIs1ElVoUr
5KAIEdlPE8iVmjUmV3T0s9me+spVkMIB84kNswkJ6ymvHYLE3ddXyHVE046Z4QQI
KpqY1CZyB4SuxS2SRE1KJ6Jyb65uEs5B/ql9hynVxH2BncyEGu69Uo2QKEs4M26H
Ui4L6RDJ6FjqGXwGXGzphEFUR8SHype286pq3vAHeicezPQX6iHsGA3pI9BBzKsy
dE4XC+e8A0/hctg8zRBQwXwPhzaUS6Rk9wCMTk6iVZ0topqgr2Wxop8bktOwpa/Y
NnvhyhND0eVU7+MNKU9MaaWafi77OyPVz+8FhuN63jcKLP6/MiyicMmn2T18KVJ+
3R009cuFy7v/KcdnpJzFuO4MSYRM6mCdsFfoRbdXNwkY5wBQuHg8YcLeYZboBmhU
7Sf4ARmkgFWzcw45wN8i3WKTI7jBhwOITBUQ0ARbh51YKrGJgHeohrKE+x6Iv+QF
YvXD7JuPZA7czOr1DJoOvUENeby3wSB1f3foMg0o/zU/EDgW1PN/Y9g0rhDRKL7R
vjyBsTDhjFn2nrMvWHrgzKJxB6iJJ7C2pSx5UFcn7bnlFtJKd8IfVMGS3SZ2BC33
GleN/9Tpu0zPwRarL9gqM8nHcNrCmvPVk0MOVhXGGG7UH0R3LAC4fcJ+js1g3eBd
vWKUn52588cNfyr/wXmUj7Ran5pEpI+JxrxLji2EqDMgZ8Y+qLvIWHx8lvIEcLEZ
wnFoaJJKikZ9b+9rZTHADKVYBVs61tQGZLTQ6hkfRkYLTEM/vHySmiUIluLlfE2V
4Iu6tov8F7p6tnKnKgmQaouebF6CjX+24AmllfarbHWMYsBo4LP7XAEJfIGdoZ+c
OZvqKze8nM76hO0d14Bxaq7j+ljFcOktMtp8wWecrqF//MrEPcwhGrE8tUyMjaGW
Gek6KbHNMCHfr6hgUrNt8ndZ6NQpcE/bglQyWDeuWX1yxMnn5GKaoAveAd80shqv
7O593rQABXnw9OJWWDStgkCk+dmZF63csJK6rqfZnKcv/L0PPy/J+CoIz7Q2MfFO
PSJqR3AoWjxzZC9u+RyqUoMD0cTtVnSX3p6nO+7nH97e4ViPGvJXD2MbzorDl3Gn
ygP9eeBEN8jFOuX0UPKclIN7mpwaMqXbIG0g5iHY5Uw1YZqt/0GNO8/7r2H3uxEQ
L9EeJrYm9FAhw+TCm8XO5aPwNUQG9yYFGeYt6jB0JWYHtNCfYWA0MnU8gHS/8Grw
Tw1SZsd5vQy102S6nNedOdPhIRR74Gl469Q7bhWCFS+J4K2O6c59Arpcs1LWH5fj
MbU1r0euzARmVgM+V0Py40oFP/Jl71yTiFbXau74uZ5l2IpBO41pa89H8rtl83Gh
LbR7S48MQ1L8PVcMl+j7f8V9j4jQJaFL6GuYHOITwFlKK/mDkcxGsSo6l3+rPTXI
JG79hEO+Mr31eeFN5GRJB3VFR8tneLO+pHwgUsurQcsuP81OE2S0QAMupwkrNrWl
HZB08uYidMjBW8dltuoEXbUkeK3ei/0twPlPRjjKAlXngYB3de0pRwCdHgRTecym
sWw6bNcPtCZPzWr91NonsuEoy4EmrtmxaTu9fWyQWQZJP4rjhinTcFvVdNmRNxhS
C3tz5QzZJGy/CQPJXec279xzq+OGfXQwXCjdyA2ij0Gw/0W/d8Tlbev2FWUsGvJ5
lE6Ej9yIbYq1kofCcn1TtK8YTJVrG+VgczL9oWls4o8u0CE94hfqwCEvRjCMRNVb
vgXc+ayaNkVo96GS4caqG9OH8OwFwObbkAcPb1aS5qoduk6DByW2EYIpAKoauS+k
5hMqyYVcc0HDEDvXakgphirFwvDNNE88WJSVb4G40TmfCPIxVeQ1cAhRKXHxgth0
7u4hRKzy06PnEtmFOvWlGe5HIs3yYRaP66df7RHlUvxn/asUk9u86Ixt9Wr48AjW
0bXWQYB29Pkng+FchRzj5G5VNaiR1zz947S30mIi/YHJegDT5V28Ypx/dH34A+xb
umNnOA8c1+5DzuiDS6fhzU8TcdGvaUHnOB3+k0ijWliOqAEWSQpyd6gznmaaHyss
BDK0Yiv1Dkhg7p0KqoNwRxBnzq22/gCzFoMJhU76jn6JMqeewk2yHHAgB0ezsW5l
7IHuadOaJRNMToC2zk+AbyjwjFDnVqbtltel8kAIc1Hll0lEhLCmRZKb2KNmOwGc
E2PYaAr+Zog7D/6spuFCxnNWZ5LsFCpRSDgVCbX4t43Z1SJ8pCT4LvpYqUtLLuti
q2aHdEJ+uwOHuyuCaaEx031I459C0Hdg5Klhnp1cgK45kb7JjLRySkYNUzXjgXWV
WCkgXKG60IAbK51bxpuB49h2TyvAwtx3pPPRp2KOhBj8YyQgeGHjPv2icOJ075sU
dhRJITUoo1irfsZJfNL2dGFI3zSZhBvMNRo/taI7GABjMogpZ1AObmoDEc+VnXa5
BYOBSKORwaJ0p/Ise17JIit2CdVGGMP50NeNJ7csZqTT1dmcGbs4E+VbC9OqcyaB
lZOO6/A9Dz9rl4UuuP0zdGj4CNSSAk5zDDmf0ih8qvEtauEZYr7jtaPUhw22OQT+
EA5OU8UPvvjIqUa0qUcBqFPbagiI7SU1Tnpkb5VXWyXykqNo9tbl5LwTG+hrhSPw
ZuUT03XcA2agHfCAalkAaKXyIwzJyI4nDeNiZEsJYmX51Sd/UHv5pbW1FPy7t4Kc
urR278reyXCQBjLCR/JSGIeDa7/eZSnOT2VDGyvMgDLrkNxf8alz24dHL1/zTAMe
/IrOqvz49y5YPmbYlkn425Ic1ZPzIKTBPtN8uDz7T2tzzXof1y6144WrAfhMrxHw
hbW4jlZrmkwb3qVJIXZp1Fk4SK5Z53wkoEeJrxScLqIzUAhb9Xq0X+isd0IRmiFt
/rt/fx0OTeZ72FUkDgoCl2WTP0dQavJPMsisifDdthMQMa86M8EZV3Ccmx+HPGFq
etAeQ+kVYIAGB0fQxo+cRd1nPFGa7Evl77Ff7wl8Nqm/sQQyThxjvCh96VdoEW8K
XCYNQ7I9PR5l7RJXsIZ48+fLU7tvgmcwQXOhWxBcDWRJhYFH92JrJcK0MVjenEcL
NF3mg6y0geoHyrzl5vXKH1h8zEj0hXQrPYC4U4W2pirXP2j0aepI6npGFAOpPuYp
ImcPYq87xLTxugmk7M0R5NfeLjvWfXi6Zc4M6cEEJ4IJYQT88dKMQ/B0FJw7mAxH
KxUEKyv1oY9z34Ws2LKCS84wPlm7c5pQGEpb0e4qYQFf5oBJ96DDAeYUbgkAXF/p
qHrIbEcOxtCtb2IqbazfhMccG74HNzIlFkFTLTwjGZFgrcEgvl/A/uEjeUuC1rO1
vOjHUIocXinxEqNUQ443FOiSZgeu9kaVONcUMGjXp4pE16iEfME3i6HcMtCZkSFA
kck1M6j9LKGw1o2/jVbDK8uYPltC0omviK2goOxILg6oe/IQDu7rKv5PeRIrtkpy
7ssg5dMizo6FafQcOuWATDGPcZUecFfqLD8LQsq4lVpOM3QQQ/f2vKRXvXe72xvT
02BRxrox3Uubiec0Xzt8Gc/a4Vd3ZPMe1QgRkhOSPwVWJjvqnJlHS3Mn2NSe6Zye
UNoykeGlrhDTnOu1wx8g1pzDhqz7fSe4UYQI/yuALZ5DZDuMi3Ih5V94tjvygHvZ
z63aSwefEDzVVAuXCBkySIxsMVxf25PTSThQMTqs41HjiFBiUasgBrEyFz3UJtF1
mG21BemIPMyoONKFndurE5zleeEYZtK5OCH1Z4YSR0XieblgcyQg2Rf/5nBmULRg
1ULR6xClnejQ8uYuYShFfcg0zWaLZ7y9E6bH9M2MAVxp/nvF8JkY914dcBZ/b434
QNjcF/bekCKEMj9JcwbVM1EJUPI29DLA2/5TUIDqq7nfpiy5dyj0VuVcAEEesCZp
tMH9TY0ziz5AmkWTcdamMoFywZrrs3Rht1RSlQjvlrFOv9ZZd71xxfdqcV3YqfFG
xIVcxE389BspvT6dnpWmJSVXLM27Ng9vrm5jfOMp6LiGrMHfd5qILIxfx2Bh/dqr
YM96Gnsrgufxlq5D9spkEUjry2S6SGnOQyQo75/dFmU4PKfxeuCixpvIvRJS4vVO
PUiKJyXXGwGjqds9miCIXL7ItwtfsUqhTRU8CRIvTbz5r1QSjjthmAX9rLlc2LWS
1r2SUAj5rKJGUhRjsLz/uRW0YlfQXm5WK3wgWbLALie/9sJgaOHUsJslTxqKMNoL
ZNAbSNF0reCIyLlv4iCCXFfhj3R8nTecLLY8/yliJya1Ci9vuPupc1hN6iCZqt5u
2KsxbWf0zm5ZeN1XcyotE9l20lGPmqqtCoWiGj6+3wGYy8b8urWFHDrWKi/U/z9Y
2/QgNZ18jcSLUgBuqvdE8b4Yks/dUOBToHZluBsqfLdZ7T1XEaILaxwSy8fzzefJ
fBNQcLn7SD9w6ed95IJBL49zhzcaGjNn+eZXgISUnOhXLs5epyokHJfFqRKV0YBk
aNHbISLND+IkIjqUV3m9Np3/cW5jmdWS2e89Rv5XPESlBGif6c5xy6R16X4p+cgc
Ji290RFPHOCLTkzYTIAALjhUq7832ddkq8DbajWcsEh9oVP8s2IwUWAcsa/RrFrb
v+qdFK3RzQb5X4ucYCIWFlvGrFmOwHLhICNIMtva3vmsu71thYf4qFMKy58DB+3+
nPKZmk30mlL5dCQu3H0xf0t5eFfPJb1+wdYZ/vrqgBenqWPWdvHIN+qj5vvgaWre
fLmU1zDA9PJ0rPLg17FRspkPz6QoR5NhlcOMZVB6CmRXuLnQHKeUJFAGmGtya34W
JtzUl2k9vBZcqATWX4uB1vkHfK2zMNK6IniOdIdw413W7j7pho04R+zNiWHTfmSh
Gp025N7QEByUACdQcffMkuW04kqChWWbu+rXQIRmd5YCjh+NUgzxFtnWps6/Tq9c
CHoRMCnSkN0wYGiBz+//2WtjqPDHDQ98FGI5JbbQEzlF96jP1ERtCvWwol0CjURN
O/R3t/Cpwq4OX5Fw/0+Avy8Z8c17BOu7+h5O4wu4NucKBkao624lOEiZLqst6f6z
bEij6RAp5OXUZ/Oo6O7rvxxUMC2FwRN9I/W0LnQqnRMavqejcHos5aB/fNQItVl6
ldy7sct79TYtD2RkyNAfHUdAPLTS7DDqyQqKU+TES2DS4wMgG7kSbcgYtBLi5ejd
agSiX7qqZ3PS/gtD0yiSi4onUz5IUeYgqiUqK+N1E8x2gmr/pPgMNlUHKZ9c7BSO
SRS0gpwWzb+U6AUehoV6EiNWBHxMWEsbblnHZMXW88XMWEhqUth28qbaG0vx51X/
ZAS3ig0cmpGpgmR1zBB1QI/uYSaTwpaBM2C0wHF2OUdzLtNOFGGZRqG/HwHF8d9u
46+5RGji+hENrDCN/0gfOFrH1lrEeokHp9XIEv82kjjUy0c3it2k6sI7Auxs8kye
CmfgTWx46/7hsSi6A3wRuQ==
`protect END_PROTECTED
