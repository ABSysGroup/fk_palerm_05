`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8kd2TxmG6AylXxli7CQ/0WrZNuzf6NFrNFrORVDsW0/9pwU7BRSHP1Yq1Xi9/976
xaay3EEJEsC2Wyj0pO+lRfV89Xa1nzNDsAx9O2de1P9+GhyW9N4MVmbA+r6cFXYB
Mz0Xl2EITan9JKsCvQKUvYf4bl7VYnz1afzMF0TitTDbCvh333zo8FAY4P5BkY2+
xJteRFT7aUyce7xPKC+/Yjui/lnRgQKeyTlHjG9cJUy79+r9Ux4MvWU1Qtb7x/Lw
99UVMZ2MfCtrjt59WN57ZmC3UGUaD+My3MTrju4fQIuR/tQFwn13pgdcoHhKgXrQ
aV6ZzFgD/khr4Jx61UTcM3Z7fU7DbaNzahHzzXl92TQmZ9ebFFfLNiBp61+zjE6R
e67fpAEBAzOOvfkJ8qtpz2AA6GwMaBRAKK6njKjcB1WSccLoKnmtAdzAASKewLup
f8gRUu6hw4f3m+sFQLQ1GP9TkB4zfDW+VWsxd3/1ErVQIthqketaZ+tbuzOjK5H+
RBShqIsXu2YmlBhrtEVVXtwr2iI+EBIVCMV/KPCa/s3/zu6rIjdrWOCRNDNDVfzT
uMYB5LPDZFFELRy9mJ8dapooqnx+fsbouvA/bCJY9eagnPjCvbXp/Gteg0NQziRf
hFuOdBLqeDiTltYgIAXYav0LkCuzVnJUiik8GKnEJdM=
`protect END_PROTECTED
