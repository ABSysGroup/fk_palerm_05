`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/IrFXQzszFbTxPPjQBmTwYxfgH9qbICfpwpDTFcdROQCzaUusCQTSunw19isahSs
FYG4+LDOquvHQQ3WVJKPfmdo1PcS2Q+FrZZZB+pawfxABeuNa6XZgpqkf9Ly+sZ7
ssUuQdTeWsGjF0hl/96yDflwZ3ArU8fyWRiVImVFDiSuKM+NlOi4XKytgHUtbefS
sHUSkAQTMHJp9RftwocO1ehBP/1lP86VCB0zMTc31q4Ui1vqYCJwXmKZBWudku6R
YFGzf6lpfETsGEcpfcWpAugL3BK3gL9Lz1bhGfLL9stFgvk79Ix/ZEZ7DUga91L2
E7/evzqjMDcP5jQ2YgKk2g==
`protect END_PROTECTED
