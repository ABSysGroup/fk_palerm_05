`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dmvxMRJa4kpu/wGVNp/OsqDsk2lsH5XgGpnWIAF5tYNMeWGd3oMrDg9O6ezAnOG4
sXyY8ZMtwgoufoTX5A9dzEyGM5o2NVA8wdZ3sxOT5Zkm919fY5O5/nNTLPWiqQt7
Aec1lHM8SACcY/ZdBixV/J/C6Yip3tx/4pBrYGPSVuosL+UdaFZfbxriDL5GNaN4
5dsEEWHcLsS2xfa4FV0vEfYHhQoBns8MTWVFgh46bhgz8O1++VSQ4/BrzAnb/rdF
lisZf5dGhZSB4NC3Mj/ESKpCOH4MRPVsjnbQWfiqBGtas35HT6roVCo+HdPpcEla
OQ0KeVxLgMfEP/VZGdTVRg3DdrphY53KLwhNa0XENqKl83vmljkStbjCR7gn6rRV
CXKSf7d357UWs48hef1DPDCUPWXWQ1jqwHl9sQTpImkW6j7yUPhceMKsk1f7b8RF
siUn36/aGsAhngcWn7TZt2GhdVFEMy+qPcRd9/yL/zGkcdEhIZ71XrZxwwsxnzfb
gqePasMR6GaAoUsz856hvyT8cT3G61sfBomn4bh+8N99O3kui7Xg5A9ljXF4BEsm
UX5pLbG5byrURI54SwbSRN/AEj6X/EmGmKXcGiQ8dGLeK9zHI/gmQ2bKjAE0iBv7
euQPXM9rb94FklcD4o2rHmuO7iG2pWCbvZu/gY6nOZFRzrHSvgcSED+oPUZYJgwS
VkFK1qpPi6A0R8i+zoXH/LuiIcUiBRdyIVYDg2pgv5RlZAzmbZlYs9PsKvuWHLP3
u0AE2t3QvhXbB1zkcc/jjz6xgNZJc3KF9I6JfoalQfG1tZwv2sZNKdaODl4U2OKw
r8Q4KE4uPSg9miFav5D4Qs1cO8IQGTbB1UAh8tst6OjVECW52960ZxoEIRnuxWVM
o+jKJHT6065O10MOOKNPeh2RzUwWHAaZpQ1C9RKXuceFHYFbFOh8eq4C/eXvCP9R
a56ARwQ9gT/Ee5HcRBG4l1xqjZ/tE0K+D7zucFQnxnuMycsWbcw+PcpKaBhspAz0
dgWeCaCLJNzgmnTsrWg0giWLXhhOKpDfO5P89F3w0hErR8Mqbk3KFgJFLzt7G4qG
47JJT/9M+BkW2tethtX+6JKUCb6I/tSiQAdpWz4aHJIG/HsFJDw5/YFjJCAvkyuT
iPesmV4HhG+cJ0m4oISUVR+DxbTE4edivt0cGV5tR8wTwu+akmvKzFcK8LUNekPH
4KK+hRBEgX3uCHRi8iqmUy5VBUeut50etvEL9qjzwJGwMs2fnvqxouwW5pf6qpwW
fTOTHwrKq5nY6xJPhmHn1m4LQpVPjwl2vSR73I9YRO48B7dn/nvADL1kZHMqsAfR
6UO/4BJ6N/BL3/BAO3oEoLeKRNgRXgg+H1akgBRX0T0AbnnPGWSQKBijchLFQxc2
ucSIpfZmQNCbBEZWzu2TSyHrHM+bAIwFID4TKdXgZIPZSTD/V4XvE1emh9ZpIJBx
cEWhNWsz6UQ4LOeJvrvLorJdGyLz7Co9VCsKtC7OwAHKGbgXjvvIhnTiVWxmsjMO
51TXnkcIR5HtnsoUSjmJYvjv3PXSlAuO0sbrDsOfo+k5QncBsYD81C4VfUGoFuJl
MVQlWfycLzD2IMtESPAsYS38jMc++pdHzuFhhrte0GClNpND9m7FQYD7uN7aHKoo
gwAUQpJSPLTMmagI0UrQ4iS9RJRs+L9NnIHiixe5FbZQD3I0FrtU36Hcb9V2QGHY
C1mZYARzt1CXkJfkcnyFThbvrD+Pjkoa6BldEBnSwW8hHrE4+r0Lc89QTDMiacFW
4AvwolCBCnDwV7bLe2Z5Jfd6YwFI6pXWIcyX0JWpyPT3nkLN4x9R4wEJ37dpxqyf
IfOPOQqb9AqGNFgBCiZM/DRyX+JKZH00qyaOSR4aS4W6Rm4iSB4HG0YqypfiqM8O
sV8UddNaZG4rwnlch6TLGfEkVWmaF8cn/rGIz2hnuuvYTFy6oEZk5RqSSSekrMn6
/8DhWbgN1y7g83YBay702q3fljgRw3jsGtqh2aeT0R+q2m+roJDOFVRPtQPi4zkv
wsA+orTF2fk+CCnCOpQq7x4+yvVjp5eW75/ZPDu2+xnLOG1gR9fu2yxxPuWVftKF
LmuExJOwUgMBPwsMAyy2Md9VnJ7SaTvObOHEUC7jMjSeS5oPApOjcqD/BToPHtYA
Fqi5ln1FTqnaOz9GtGrJ5gWbsYkA+JWhJGNgVeihRc9Ttx/ImdNEgG/c65HXVXr/
bAFc2VnwGuBbrzNB26py5xfUnUl+5egJYoV1H9tfgcwarBSc1rmbIkc8sH59NqFA
CewRWPYCFVVpyPIOgGCXZo2IYcrhbIqQZMZWWBaP2Bkdm0v+5jJNP7mG8myhP1oM
qRvBpPOooM9NirnzzTW32HCLFRFNZ3PeG69Y+OAcb5oOk4G0XtiPHg1Z32Wp79ly
ybSn0wPSIRu1jHCGP2WZh8ESwcL8iJBht4m7O5xMx0nVMm667XZeRjy3NtjD+yBt
Mwd+U+RqYMbfGLhlyYuhalBvUI8CWzDx1l9sdgklue78RxsQKA9Gbdfk9il5Y1oV
mLq8G7x3Nme1oSCFP1libvo+Ykg42z+faJ2e4Bj2a0nvG2zzfk95DsqKOdo1JjLA
6pH1CgZoT/zXiBWt8boTUutEt+oA7nWr7Ti/8Lafc39OwdgKHzvRRkilrc7sYXpw
yPBxpE8NWWU8f+eKp2SksdG8wJsKq2BI2/2zYNQv2uriC666aU4RBKRNIUP2cYeU
iQCqvkHhLlAnQ3FsCdp/g2+SK2JIQNUk5uTbC0BTnud3+EbT8kM9QgE7Gc3/5wAt
Y03T7zFhh4XfFT/3Btfkjmy4QEfSTAvC/CTHgNWq3z22HwIAaktK8WQFwphby7yu
Oo1+MAKqUU7ZxTDEuUci/jFzWAD2A3pBVflLicDtcDJrhMuf3S4yawy+hVIDfw05
Qq4vWNgftgrUY/MtHhe9xcF+mfUUnFV+N0zFj/5jvdojDarhGbic57lzKQpKauGR
SEWtV0VsZ8ZKSW+aesQhL93n+R/akaajG0MnA7NlHfbibyURJ2Z+q89dvBBYKMF8
6CE79znE/tHrWEGic+eQ9RGD58cM/1NyyVfEDsDjwSsXgVnuTPhvpiyPOA7BnJvG
d+7zCQ689P3gSNKtKuqHrCyu6nsYZUi4WLlriWTgSvUsYFVuWwxuePgRLR/kysnc
wWLOmhW1upRVYuET7TYsk7TNbkjF5BLcqwGEFS3J/6Jf9OgarYfjI3tELwhiI7fg
Vlc+rVAbZw/mFPnm1mz5qKYwhp70LqWOjC4XpxKv/F6scaAZlNtL2TcFr9+uXEUt
B3CMVfZORi7cDohbEiw7RzOqKr7QOai40F4Eux9wK7rg3MR5DRwTpcQ12hDnIxcy
vAPemUwJeo21JQoH9QjUb3yUahL6dE56KgQsHeGO/lWdkb9VmX+x1f4XjuYM+yOY
H3/6wATIy3jyLls3BUThRcxJJ1CknGvf9LxS5TZo9mRclfd8Gn9Zm946uvuptZbg
FqX1T8jxQFWSBVbA0wABW6f8jgyfg3fnWdlsY6zCPXt5xPS13RmyNA3pBkFwrkeV
rqYubvXBp8WiQ4z6iAPR40dExU11OWB026SF/xISgqw2DYZaohzVbJe83c5z3a+n
EBFDzYyRKxY9qUmNY1xIoddKcFyJtT5/iq6Rdb4cGk6naOIaOFc3rHxAfqbKAhzV
gjKGYfqVxdRl8KoGSAJqLsdHZPeKzp5IyK/jssKg2z9/Dqbd2W5q31PfLeYX2Z8s
EiyNpfCfrVvAw7zuH860zna7JWccUBHuYkLMIrsyMcG7HK3nUlR/rZD7Dsm56gR6
ZFrReSMNjxKF9Pru2dJvjvS3FbGz/7Mx4lsr8559msxZtkW+kJQWPGY7sPQYku11
P+9HTF25Tl25U5FG1TCT5YOK5AjLNYtO+nmWi5f3TBxLyiyE5IQxMxo94cAk53fy
F94MIH3/sAkVJ7Tn3mMga50TVbxXKYW4eqtRaQRqWjtFz1PVRQd2xEMwgp0j+JRV
WpXOmWqoHvY65bMQWCF3+geO9GQgDz+OWUHE0Y0am3uGQPETCScwP7WRwxvbCtXp
AB9iqds/1OxTyD3+WK6lu/KQ9XUAP5OEyC1cXRvHdobnKYx2Vj7FyMPi3xoNC7YD
wYdbi0uOP/Nt1hQULrMlowa7conU9JO/cKyFyauz8jGWEkG8uAJh45VqHOxXgCNM
g2j6vfp0KaAyKnAMKUQmKC4bHQjfnPDqLePpSniflZVub56PtksHnpTMKVD2tAOp
BpuQn7t6q0M9RFUSX8HMBZ5SWckC6y78SqCzLktDgf5xlZlBAkt93Rdlbc4IqLnt
grptI7zOMISWolB+3RlEgGeLu9daaJRNaz44+nCXKInUp206qkL/2eJ3VZRT8TU7
BqqgnDHqaRbO3GgfeRE3My/f3HoqrV1LaQwH/kMUXMGicoMyNzlfkNgmQs9+sWkJ
mqNkvdrrkuFYrzXv1asFlvMUdTl76g36e1bMFZr9TESe2EKs+YdVnYOkX2mtSv+y
+O/xUvnuj95NHlCzdRrnbnup73gTtoOTMnXlLnhMDbHrnhrrD7UgC1FedKec+kMI
ImnbN2CEtuIF8T+cXIeXQj8YitOW+2fxiKoGB8RGJixl53AURttAaskKD9Hsvshg
p+MtROD+09GUYIG6MoFuMgB1pbefcKG1fDdkhE70LK/+r5uZNUJxyh/kjySYJKTM
NLTDEDeqAHUZR8kLIXp+ZN7ScpsjKsJ4/D5PXEPcLti0SjFzYLdAcE3FIBWBm0Cp
egg3z3ORj1osqZeoLhdF89djimUyl5KX4s9rAMGtqO1eAqsYMmNWGI9TlrhdRgiE
vIAjfEZAzBk7oTkgk/A/lh5d4kuDuNmDyFcD5jgzR8spz58V+Ms8cSE4Ab/y5mc6
SHdvppjkExNCFa0M5lSByT4lGyxpgjsvQGfSk9Z1vKVPuOWnRUxiHZ+yxkWvjhEA
5BctDbtU4A8EyLzir7ijs2m/D0kqyxlqAUpF5m5W3VuTH81KIkgFvZDWqWKf0oRa
2I9o2yyTDMFwcuzVJeweZAQyeWqvjl7Jvc85oSSuV5TAJZV6ZOIxy6WUOhz8Eakp
XzdFIVFH1J1BGFlUPFK1tHmegybrXO6WA0F7nxJbjBzjfC8LZTFyh40OWKAhOeQe
yhwpnk8w03+c1LLDst8nnuIuzrM8mE9bHIxlOasndovAJt6zmNvH/Q6Sci9TOwFW
ecPPRO8s9oNFx2/crkMeA4G0qgE/2HGqLuhmwY5PXr4PIMzGrICCMBuI/5vaIloj
+CEb/AdUmmYjvx7TkgaFxbOkGXRZPLYJEmv+yVAIxEbdF8Q+UwbztdcsaX0DSRJk
SBSJTtcao9IzPeHcIiPKQNByWX2d57nPfN2nlq50reiyFn/rbVsbkAQICRCt1MDQ
qS1+gLtbZ6/n0iyqxJX3tBnmwHPP6EyxUD+R0usbR2cg6+LQ1fQIU927KC/UElcX
d7q3ziwJJXBZQBGlA9OlPY2a8KIuJXDyUqbZVrf7AX9aUcCFoEWLgGKnYlM+i8Oy
fQ2RJ0MVc8SuA0TJn0wvBcsLpy6FeG2UMOSEVB9Hi7I53OBOO4MAt3rduEqyRtv4
zT32qzsMn+wjYpHpMAb3duBcEZBHfkWNKOHDwExwpjGuyEPLv1sZNqE86x1o4/RJ
RCaqstl2b0cLkFmqxx3wxhoruxRc4jlBqgolujTpW9qGjMzTDEFhwfix/vGobTjf
b9TNcnhYu/O+uc8pKLoC4G+OlXBZPAgW28pqX/EaX/qSoaw1sKSUUUJpgqH4Ej98
2qTxoQM0Tb9OwTUwc7deW9mbhBmnh4g7ZQJAhe0ii/JUn1pfDonkl0WXYxKMz7G9
e7wTo/8G1NoQi+TCi4WsHRUc4K2XG+HpA51D2ZEBsFHhfcWr84rOww+LzL1QafYE
1jYW9SP3bcDrLVZhhGRb00nMxyBSg1dHEdvjBac0Z1SbyA3t8ZINLXHu4Biub0s4
d2XQZ/CwGi2dWv4Au93cJhY+0sdIXZEhN1MZbejvYYXNTuMv3+9iFjYfPp0mYBZm
I9MralCWGPXgwwfWQE5a1y+wvQMbe0BNCYkFI4sbxwdWkA0x76rhLFA7mUE9Cy5d
mtkITwyGALaRmydtSwBPVdF7IUjZQMpzHDcsqy2RjVdvmTIEPDCeCb7/hH3vJ21L
shAbKh88comprUCiGg0SQ0629M1kiUo+HU6o/qFHbn2c9GGuSCVlhq2XqFCaSgVm
6k2wWv/sRWa46T+2QfQBFLw5EX+pCY5FjEZhQGxraLM8Pv2j6+x5QXfRDv5rp0SN
t7PIch5zjFSr2u7aKDVXfMDTGRn/WC5vMaVsYk22QS8ItFFyPwbEpF7gQsUPt71w
z04gAnAU8+/mvwgFZoMUelzvBCpTU6XQsjv6AhQXitZ2Gxre4cQP6ILK5tbgBaUy
n4ASgaBGHw9IisNYterkMwppT0EO6bA8JoLNPX5NKaDeTgWEIdnuUyTyXROYyea5
i/kPxd3JAOGzckJ+vxMkN594LIYSm7F2Kvs7L7vpKBUzX/gqlEhHLBLok6K8L5x8
8jvR24i0eMLj1e5GDk98lgtiqI3T2oXNW2Su3r8oDFQdvyka2M0CoaiY50eohviX
dIwy+l7UwNIFxdbdbk43N3+wWfN/rAD+NY9zhXJVOgeiloK7/1rRqMrzekIyD7Zk
NVo3BBqLc6kwGKZAo0IyQV14ZNbW9aS7yi78pAVLliydR86+ur7KL+xlutIpCRUw
Cdr1dFaPMX//LLzPUeJHxwpWd+qGO05fWw3r/ScwVRjyrTxpU9tsMlOP8sMqewID
gxBBwLZ0Of/oAdXs5LwW+aGfB9sGFPjugxXl66QVhHxbZk2o1Uio7K8AqirVTinD
xz8UoCv1e6Yt1nLx4FKAYpLBTvuUC/32cg6d3DwaXogZNrfHEMu7eC+f3JKFuwDM
l2Xj5uyh9Bh2qDtKJwcfJA7hRj0887ThSnbaW3RyGcTj2ruPuQAZTkibNCrEbJYG
xzQXArBjlaTcUjSJAMA6aUTIshLf/Eh62CwL0xVsGG53NV36MxDxj5+wolLSUdFh
9JLGtc2pfNXBnWlnY4+qTgbWkluHJ+2UALbxAa3Z6Pwj402yFVBDEC4nUUIQAN6h
VRVA68R4xjm2VCtqL7pxTG7he6qme3TK/9qGBcG3CWzZD4Z4L2bROCdRbWF5mbEG
5n366MArFjbAMH16oXaJnqu9J8ePYP/1EpejXWnN4fQGWRdRp0P6I7FTtBX1P5rN
NDbmwk6kP8BNFC5djlSqVS89zi4oU+qEyLu3G8QHVgXDty4rCh7r97OgRCDQrzMx
73m4cq2e2b9nB2wCkZauPlGxpOkL80tDXJWNcmdymm0AXuWg2HVfjxVTIyBVjm61
9HKWnW6nbrAY4jFYcCeZDdO+XxvWYGsI4cIGABqC7fFNVXYs9XEZSZEJP3zfI/EO
xFeloBCzh9DMHPTOKXueIh7oKyDbKEAWMgZCVfJmQQlLvpPtK4J0FvQfGxUDITql
W4oTtVWJm9KGyy8ExxyblC4+q3hdAFuFfviE/Dw3IsCbDq/hF6nP5YgeZY2duEnt
/uBVWXDk4a7PZcXXQ4R3/IMad6itpsEgkuD0crHmnbjRYF9STwWz2LBcwnlSMa1R
qqvPbYa7ZrOqxR8qMjaQphaC9vtiWWCgguxSG1BVEr3A5i0EFpX/upSkWk+9NWD0
YpoInovfwRU51W+1FVWIFBUfCfOeGpCYS9O0jultsMrFIBFl2cPSk2vAdpDcSTME
/kLAJ2T81u1KBR0I7A8wGPyryIxmLVVHPoCCzA586Jd6U07dyB2+Ih/1sWJY4+GY
q7OopfjPLq4Je6krJNyciWRZiW49qImEyvHHNeQVdKt17CsXV7s81OoYecM1nNRS
PTQ00b41xQX57HaBdeiXWfPD02GaPjosNY6IED6Cxj4mWKY8yhBd5IOCwoiGp5ZX
IfTg1Bmyk6RY4GAHccVwK88pKoWkOQTkmVoUjpeDHDUGW/Yp0fo89v7Z7d+t16Ug
/l30Xp0e+AVEaErNMj70vzSGzyGMPL7SmSxujDbYAONptd1cqNkRDFK3bytYpU8I
qR0MXMP56PnGZL5WonGeitakM/dHc6vWasNHjEbapNllF3ffuZnVT7uO1xynpU2A
Em1mFPpmkFLLV4WdgP3vjDu5i1Z8jMueDMIXC+JjXSso0lMnTpDwT2QuHPmVBLms
aiLaWtj4mSTh3/HK5uSyW4XZVREASiUbieaE8eUVgFZ5Pbibjdd3YfCe5b9ICJMv
0OupNqXpZsI3PwwsDDrswcajss12L4iCfw8zSXgWyS4t9/DjT8dlxC2FoJlGk+8y
4TWO1p6Z3uQf7QQEY1zejeoxsOAl4lfzbDJDYVM9/ehHu2c+85S6SH+Rfwsg4ocL
cDfsS8d3gRAX/O0dmb7WmO7fTiHo+59J0f2idcO/c2x3eobRnWxD0//6/gtluH/K
ewaZqzXeA/Jrq0Re2NrZzue1+xLW72plh3dW+0ayR3xMJ2p92s9v5dhYkslaSQyH
lAeDdyKuEOnlrpTSXIsPytofgWIMjpHF7NRV7kZGsyf1z2FFDcDXkuifZXghMxo+
aPV9ewGxnJvjVV/bXVaqt5YFXv4CXzb+fSem+BHzvGcEim0thUSX33L1KG8XJ2xX
WREqwTAgzi4AU64RErivYtX+G3klKb15A3fHbTvKxqxYvq5RLKuQLrC+9Q1SxGqF
U7q+LoLq3oM0Or/dD9rjl2NFSyWBPrwJsGdyA4J/NnUrIpNtam3Gi8fJItBz40h/
lIKHQE7RFoDPQLuCs8bF0uKDnew39/FPJq/yamNzYWhGgIKuDmjawKzIPuyCLeDg
ehDdtO1HQ0bMqpEQQHsGwz80qk0M0kwHJ4C/N8dTP3Ji2+Ijhol5P38+oQGeMDRA
/48GhKbzV7xsRRpb/RbgYH6+fY9JPr7L33mQoJPvyvv4folcqhTPPbuqDfeiqRK5
8Sgmta38PqbXhXactKf3NRnnxJ0N34iy4/4qmLHdM2Boz8dwEnFnIcvXXPLS8LUm
xmJCpYPQHsPIInqulzyrgIYX+SJpH6zy2RxbXbiBvXsYaasAiA7OrCC9YsH03z/m
d8O3bWGMhxlSitoT3JJDEpI0L4+ZuvoOF/Jw4Qh8xFAL3tyrZKHS2UffIO1eLR0M
/Epg0YY89B9G0rsCWMu7sUAJSSkhdZ/c0quiLZkqybIEbpdLZkOaMPGepECuDKy9
FRPateqmRhO4x5lqUu4uEAZ/zBWHX9ccwq5l+VegHkG5L2ZAhn36GHusGhtrChE0
5vHtooQpPNR+b1UswLOmkzSvlomz+6KlX1Kl0qeWYfxK4tuAtCMLPFII2q6HN8hX
2LQa82IDDw/Mk3G34ULOsjnbUqSGDpRES6LD/IGeLBVITDFMvfF9oJCKbCRtYUB8
DN/2+UafmlG/Zkzc5Py5uTufucMHZvHkj6Nnj1IVW7cz2Nvq1EjSYuPvFGwQHL9z
Uwj0beHIOnejuj5QKglLHLDVeX4Gl+LlQcmGxAWPbmty2nm3DRyHbJj0SJHyyvCf
Rgq+lujAHd514wHFdH8Tr5Z47UQ5gfq4e3N6MbkY9ugwDQe/3WneRaHzqR4YIb42
8j/uCISZ7pVjzX8TxYrAubeJqKIlkWcF196TSVG41NYg49PelO5jxnXQxFLh20ge
iY4PWJpLx+k/Ppm+74cbJVA6W2NZakgrRTQ72BYoDt3DI/StLDeWubZDkrn28Jun
+erHhmMZylMQ2mCZ8J7QWu3JVlU9uLljO0rLdNHUZknpHQ32r20NE+xf+w1QwNn+
YICaBH+JWn4YaBZSph4MMfkgdysbyHix/j7sX23tOHnOrwGusXEUVeY6HZSbJTac
MFbLSwBJ/E+5VolEzIo2/UD+WlKzfXJ/zQVuPaAeZAN6alepgXI5beZLJ0Z6LF5h
6+NkQTwqmjg9Hf/bNb4/5GM7ikBw2F7BNxIBc9fQ/6atpjGg8bujRCIn6ARsC0UU
C2z4OkkdpDJg5DptWF565DWvqgnJ57t26/S+IndkHT7gqrWiLva9YGN39/qR18ai
2/iIqVI2YGZCteUS1zoFN7zmvbYQ9qpsezL0Y9AGe279baILTA3+N8W4pWPh6sOV
Uv5ZM8oYNJBZi5J6YIPlD3hMp8rzyzgI61d8xtNddMJr+zcX6FOPXucwHMyK/EBL
H8umUDtW1U3JpL4PRCOzxtCoMEaapvMboCcR5S7PLQ6rLdQgSw/taed+AboB3Mh3
Uiqh7SbNJpQ4UkVx/I6pb2OiNqWoovHdSVu/1XHbUSOXsOMcgEtbpvfnxfGS+jGg
xU1QpZgoj5fY8NeT5+bqGgFOMrlaI4QgdXQrpO7I2xuCqhJJWZMZAfskLdAzChVM
BkeK6HoyAfoh8jaoXSIz8dSbxFEVfFeF+QMcLicLLjoHfyJ+ae4R6DkDQOxFLBRj
gwCVWM2LKJz3ZxwPdbdu/tHUqAIVR0rS+ZhiW0rJIyngpOYsV9Oj36NHDjdwyFfs
kWbydS2LaX6HYReAPQSVrlrqG8QuemGPneDRUibxEZeHnrZu/riiCWuTduL/kSA4
QBYcJGy+ta5wCsaQyAxqQbSyLIgW1cV4v2l4erlXdTcswlsm3/MK/o9QvvvBV2Y4
cohFHNCyIFH7uqzZl9i3pFIgQ6RHRTWxd3OGZ0CL1OER/P9HtzJVg8av+xPixTdS
A+T+vwY1GwRFp1Wo4b7cQqvz/d6dOxwGzgDkPsUuO0nzRxQooHxMJqSH9m6eApn6
JC/wbuuYhnqvfKkZJb1g1dugerzCSf6Fj0LeuiUdBskvaLvUJZA5LM5H7E5dgnbJ
HD9nbhKD/MGBRZwyjE89yxUgmSzMDUJI8422PBenCq8LSUjZDOsGuuFEMaKtCJl2
N2GB29kkPkvJYUG0KUqVSoF74+AQ73iBaQ6+J2rQRoCy+nE5qPzjjEagdgayTx+E
aDFYMtWFUdyXLjLSlamrJpC9R4tfGzcMcL8IDiJBVEyH2w8lvuNJsZiJkwcD297L
viH6QqiqoTL3WlKR9WO7RaF4mlHMQyQ0CyWV3JavfDqCyoaCYH/nA73bmYtz1guY
lrYqB0jCr1P4tOXB8MkewXNKtoStueNvXF/z2YKzAuJsFiTztvre3L3hnYv5rbn+
fSXOWw9XJ+knCddkiRvyk6+7COLtLm/J0IG52F/lBFFxVwQfFt4dz1gRZD96rMGa
JWiI21F8Eny6baoOD9owW4OIDgQTXxgc+YL7eC9M/wQTFJI0xt1wcsVkxs++plkf
P+PtljDO+yiLRBUgI505eFsQZ+rpinK9dtpdOeDh23rc1awwbxNzMU354Iy8aYma
H0dCv1hSfhlnDsMUjoQ3RuOMkpG+EquJYKO1rS17ClOjJe8AX2yGMjYcC8cPLgHp
V6iKpbyUeSL6+DXIHgkaJ2ehlgcHOW2p/OBpUuAzD9A0hn60drbRbnH6taubnJTN
dljGa2EYQcyjm9qN0e3+liCqt4Okl5uij49upMBmdiM1kQEHiXugcvFML7GVL5oE
jYtR+7/a6t/TEwwsJFTlUL/8ps6Q8aL668ZyU1PT9DznvfivJXtmXx+G+yOXIkrI
R416dIQ2lAYshEGICbtO/tm3cTSRitYs91sUm2HbgmAl1ToHt5Gbc4fL92sIjVqr
+jmn95C2j2kSlf1iLP2vZbKeiRju6BJHiJ8bxVHhDQXfOFi/XFIJAuRUhgCIkA51
27MYRalgrdMDuunWcP7hEqgwz05C1S3NFk+5YY2+xLNSzdeC8SKoFoQldl9+JCcs
MxKAN+f9JbRvNLct/H9LIH1vaQ20DCbTcFFVwaho7Q89PruKVTuUUwM/lMOhFOZZ
Nwg/h1EHFA2UkZJ+Eo7KXf/pyZnktsdOg2odd6IoFA94stOawx4LT2oLKBhZzL6j
WL55bePIDAHh/FxU5uRwF8w9pJGDsa0PTb4zcadFyJH8QsfpfDSrHn+Sh5BSPxL6
o4XHuufOYAgsQUtUlnOYGPqRBje9wwFK2pxvuYJoNWw1/T3CMj9K+mwegWJqXfkw
XtaBZe0XcAq3O04oDmG3SCua9sqRxWfC64FGdI2ouf4YfKgUzE5JX8Zf4LU/H8OC
ytvldxno0yEvyMK8H6nwrR/qQkrKR3X9AIVpbv20qNJugrx9+/uzbU59dvQQA0X4
NNeJ4aL9iJlQQLfhqvl+tGwl6qdNz9lzr1BlURMlxFkFmRf2UXxhWKZuCGkfy20J
mXZFJvJWfG/WbKVCUnumzaLyb3RY3PoJlb+Z3l5f+c1SVv4hckPVa3qrs1Q0m4Tk
pzkpYh33ImNMNaSLASaied0+TbbC0Nz+XBmZGANsXh2B4k38wu2BY/clGW2Deg8f
NEu3qhOcFxojPgchKGKB2VQRGgvf09jaZSBzOtHymlAaAeRf3QnyjawAXwnZTm5C
leNQ4Xks4xXq4CB03JbkhRXDqvDz9xILKYFu6vzqVgrdKGYnUKp2Cr4ot8Yvz4Ms
0L8uJIxNTP49z8zdyHQKpP40SHLrRhwhPaiiswlC7cO7tcQ1sxv7gMi5Z5WMPb/n
kJdgI8W6I0wSzMWlbpYN8zb2TSsFeHNTaJWeM0mxTLTzOYK2UTnoBi3LvrEs9YZ9
91pVhBe/wazbPAy7oDcPoovi2UA5Rmq+L9hqPLmy1fgrmm46g4cvhah6BtW75uNp
CjUe+zrpdu04RDIsTwEBSPVM92/wVwu9CXSqZg8CJ/9mj2ki3gV1VUrMEWmdOeuy
99I121PhZjkU+i33cLK/6l5Ba+Dhf9TjPwkuFmhhUq9r/YbxbkrFX2hWXtc/YrEj
TaL9id7uejaBSOhmlkyMKiwRtLbxvCwp88CVWmqaf+FXmZ1EKxCqu3gNLCoGMR2k
b2VRedtbQzAsMJOV5iD8pZSVyV186Ttu2NhWCfw9c50qKgeiz2OiTkYzUNpqlxvP
AwJNjb/hqL562nAz0bKOe63O3EHtthaeQDtga3eWd4JJ6+kdpMc1z9nHGSEDrlo7
qxEtdUMOGGXUGH+ptn2DcYpUseVCnd7NGLMBrG9Pt86YqjAN1MTnUo2XtB+yP1Pw
SUwVQrpbhSG0OqXLznfmtIgtYRkHeBlGw2QTTayMwLo6kXzGO4isaC8nNtNfLj9X
4UdZygg+gvF/rQUOtZBIkQrjh4O076aw1QmyWavG2gxZsU6kuGGgSs/fz/geCna5
D+1y7Th2RbtszgKVGfmXxP+P+n7eJ0a+vgWM/Ef4gfgKPv81fFzqDhG7JKZ3r0wh
d7tUx7Ji+n7113cjTzOJM1L7B+UqPG7WQ+W+npqtVu1l9y8akpoHfC+7U8MJ3jx5
FAK3aATo31VU1WvCCon5O/7czD0Z32CZqj1bvfB1XrF8Y/WpDoHrNX9iMohO/F1a
Z6kpHw7cTTgyVoCDDASqYAVGBQTUT33lJs9o786zRzqvz0mhnueRGSTIPw3Di+hk
5msAEuwEbPmmvX+4HPBo1YZm+q0UAjaPD3DGUSJtZcA1FDC0ag5Xny5lvO1eoU4P
oB6Fs6fBOIoTHNyQfvo7KFfyCr+Yn2jFY54SXZ1kvbwWGjKkhd+QvwGQLJXH2K/Y
XABM5p6nPmnQ/SNhOVUhccjXk3IxEXr8vInU9elUnUlXb7xzPlEbLShVWz2qYLnz
ONDVgJZ7chL7UtD6QchVNMwbqfhAGeFRJqCcgxIahmydt5AoCN5CN1hii29ASlC4
KiMONePxVWPUYkTQJHFMtaIbLultBIFNAP/yh8bJC731U1sFOCEOd52WEG/+xwHd
DHDDxjRZfFQlmrlOql3EtxnybXPYyvAztCvIYNWNKYEb+R4qvdr0Tv/nvkh8cwLe
0TX6X7ymHMp6ZHZs+KYG7MDqaW+e5YXFVOgJdydWbyKRMjn3/nUpcv/BB6bsG6EZ
fxxIhq21Cm6tU2gxe9/A9tr5daYTw0lhJwTcOCCVfacQzHS8YIKcaHNODOWnlJOd
jBvjYzL+1h7ALECfUfUUJ+ROvAKLiVwIFNGgCxj5z7nCYY81lCYSt+fyZjfxEHBp
n8gFJaZVgHuUjvqCOr1TzLeW6MWqGJfkzijICLN0uqmwDW7qgGHpreVq5qWn80IS
Q/AXXyq+cDQNoqC8ALsJKORFqc4SZWriFMmFAt5pvJfrdhvG1NT+oJ6xtAfycXu2
WX1eAP4YghkBwMtGGWZnzp1u5jmMklp0RXpOO/7pwmOIUj28loyO8qh/joSpwPGD
Fo2gx/IJkbpjpxyEfrrrlsFlRL73ujgz78kHmD1jUcgmG/sz4p8g956LRXotODks
4bnGUIC2mV3RkFnjsvPxD8iJ++5gtOdevKlTzqwYUuUKq9nK3bpNUi0bMWnNz3lu
ktEnwv2YyXZCBnPAk+WAF9oxvwSf3MVYzt6+ixbeEUzhDAeWM8jekj0x7MDHvD+Y
sUqJsT8QqgJPsAFCNvwGvvj0+ApCCrPNk0s8abI/qK6x0A9qI9Z0db2jC64NI2UN
XObMMJOXuyc0K0GQwS/6XonsqO5mAeVCailmPHq5q37kt1MZO+AS5eNC88ODdJ0+
QByX1sqWcp7+qg2hUo9b235k7oAbh/LyDShBBKgs/DDa/9WeKjR+Ly3Y8dAs4HJd
a0XXLLEc8aEeoSuYMv2SG0t3nTT2XSwg7eItmasWWpfjfhf8QX9Yn7Id6F4j0sbh
GX0yeuEz4cRx+RVqn6c2HhHzAoOx8S02GEsrh0p5C+aL50VtvedfndwhE1sWvDl+
tjYzCFzykZqdFG4E6oS/9zku7Ec18+gXzVsqTpsHM+EzpkG24O2aAztnxd0TrphM
7KM/W2b7IcpH4HMAuX7WXh4Rd2tlGg/eOQkEpNZx8kO31I6wuZ9CkLiIsUhz1W1n
facToMlfrxPxdLRQQg9gVDtfjTuBa38A7fZxSnLz5P6LxW8OPHOjznRFvFexqNgy
bmQpAznh+loNXmJ4wmC1z5zpNmeljSz1b59XrEbUF+PkUGxNtvjeppu4d7yMZV7a
EnzsBPgO15cMWvc4Z75QOI4YNkChSXBRP9YvJ6hKa6aRlOzyqingRVWkT+wjes2C
rWLccMprflM1vW0KYZUQwsj3uOB1UzONV7+jvV2KCIYeVw/dbB9f+L1jA5VdonLL
R+UByzxbKvfPhrrlN2lXKmXlgH+b5Nxk3Y9eb5I2Y6imf+rChQFoNjCYPMR/8UCo
PCYL7HsOYG5T2/TtpN7pNH+yDLynyApTaaE17wZ6gQxLo/h6S5GADqDjQCajgTRH
9srbKp/aM00lozKtxXBhvmMvZciYL9C70xi5eT4PBRpYKBTO+RFGerHMiRlAuSUa
9acVLTwzDZwQuy91h74ZOmRJwKZ6E8PyVFvVjmtHmRlhcTSsnOUtyjkNwwpD2cu4
0N9eY4DQnUjHvhBEx/qD/44CL7lg35JeKjlPi5eBkBrLoWmHB5gXMoQt4j/uhNna
kvD61jcMz6Kjbaq8wt7VtKsOmJcrYpIrgFJ3imZ6POl9jg7U7rCgrgM59slC3gJQ
TaEau3BTlphrnbEmDZrjOgmVb3yHgDgD1+qvdwyiaB+wqGlkHo8VCtwUW3EvN+ZZ
Q2rUjxttNnglgKQp6WosYJ/EWQ/YDyr+jJTv62XbUAJiNA3DOnNZiVXpo3ixNWns
jjxBWhpHYQRxBomj1DbqXm4oEqOykBO0zntHM19LJJfVG0VuCxVzqNHbKnppfNp6
8fzfGpr/wMmQIJyQHyYRmEz+zRYcLGBzZ/2Nuvakl+UObAGQ9iGTyNXl5fC2poR3
MsjHmHg7+uhkzB4JnwYOL0tfnYc51rWdDSYUfxqtNzjchFHw+XoadGWSZymt4YTr
yhaqmbPKjsBJOD4UpR0SfpamulEJXMuiYQgxIl5xW6yfewRhJIm4iNHfSmBuLVVt
d3E9ZaujpxPZ1eUCwYewlXd9D0OngzEeshc9/bD4ElZf+mdGFYGeIlpqoajQHrFW
RV/llqm6DtVCrXX7uC6aKGdKm8SjigTaTVZuwU7s2oVEIcjGUPRBOr9SrwgVhj21
vhRIfFh5uDBk/NHx5lfbOjGD+ps36dM1yewYVNHAxzwHuS3Cc25BV0MYQw7eq9vH
kG5aM4rc6GbMQlaxzVjvTNnPfHiE6roPUAzZGXi2Jt/6HnkCf1OMTpDuWlvrnSGs
8rABdJHBVxodxivhenmC2udd1XmUFk46+l90/XqbQ/ZGqnV/yj5wg2AoaElpM8JX
OpdweQHoQb4xKvHeaH7kav260hq7c9rTW5KHAhT9XNXEkWuT73iVIZjzHBvYekn9
Gjt0plqxWo/wNzSZGW9PJpe82EcO13TQR/7XdsnQvSitVK8Z21KFKDzgSWEuLs5G
I6xYrJFFoGuiBUT0m5cTq8qk9drQdVZABA46/JTYJhbey99Of9yGP0osNz0G9WGB
rkdEmJsu+Q0Fx1Mps22dna56kj8RX2GPmtqmM/Xq7t1uzGa/uyDSmDeIhgE9e9dU
IycEev43dsHtK9Bx7j8P6QDlVGmy+AnRlX/4K/Zs4D4GkRj9cjxQbYOlpNKhl4yP
W/V5Vmm8h1SfjQnnIptJoa3JzygmKSZo8mdm/yB3pK0YcAxVkEXVh5P7TiN6e0P/
KiFSuP+Rzoy3RiGkYejGYcZYTEFWZ5zRBwOssjeTxdOMZ09qYrfb3Uv/yRnwm2cW
JHKtmKP6ovSZH/aMVD+Wd3pKFSzzsLMsCu3sgepKe8Tfce4k/6QqstRpXqg/N9i/
zlhn6MJk6aZpI8cHRYyXnjYo9VzpNXUNQfunmF+GZ13i1ndwTSx6YwWo2K8k/2xW
c+xOayT+5pV7ZDfR1uY9ojBU9NaUSufW0XYDvVpdLrDFeRiJIna1EkODI8k8EMPg
HgASIk/dy7KagUobfTEMXDZLqyXTuvAdKhpaJkdPJM75Nujk7TJaN47xfapkbem1
EVQ6DuAYuP7UTVTqmvL4wHcQQ3WXeILyQiNPNxEI9N/i42cPim5CliHkg54p+2KE
k6kFJEwgQ5QT1ZTrKLCCy5EbwnmU/jGiJBkgCBqrxKqwMq/wPzOhWgIpGyULalCp
Syqu0jpg3Q4VizTQTdQ/yVNSCW4yjCanj8lWNEgF6hon7+kA3zG7HqIng4ZiAUAL
tiun2ofQvGwgw6XLUzg27m4Vux4BCqy/wZXiRRc5gKmmjzRGR8C5oPTHwrnuGxpH
GNgmGeAqfoKYxNKUDaVlHK7G0shp4iWssxf89ON35nZRyM1IDlQ8gE7BW+XPlJsc
Q6GAT6WaRhs1OwjmQNIkn/jJoJn4ah1AfBXxTR5OZKCdA7jJWbbrx88Vn5dnY6dd
xpzydD/kuZsJiBa2+DqmdpzjY3y7lkXYVfBnb2sANGQvIFcTFcSNGYTbXmenHj7D
Vf4svRbbf6A2ys9Jc97YoTQm7OIhEja7lIA64DGfgSxFOIRtU7ISd/Q+NqiKLjLH
G0MCfizcHtPMbZF5vkjlut+9oEibK3RkWVRKX/8RI43MHjDX5Qn+m3AiHUFFPpFl
z37+ZPLWos1YFk7DwU5h5WaCXaHjOtXjKMYc1dT4E0Ri7e/UcGe8pcH/Sxj6w1SU
1pXJTrlPZUM92lqWxzy0xT7HYQBzjeSF32nU7OIOn+g5rxa0V5b3nLUteKQVScSE
kqv25rgPzFAsVuw1RIUAdja3mOWyv2JXNIEKyoB4caXPmYprIxpy1DzuYrpeYZc+
roI656x+4iJza7jM1kxiH7WQWj5c35a3YHRZw2HCWB4qHdx1p6uivJG4rifnDfOr
MB6F4SqvR7PxDKb6tW2k7nEMmaawFzqBqBOzXW2MHmw++lb+6qxsFFpW3i84UN5S
cXCP61JQYsZhZLphQG14+g/dZr7H+pMTiqYq7JG/j2GBMk2efr3bnAqu8Uo+WgWy
gjMZGnqdVOwimCaiwBGcspm6tnbilTx1fmj6zFkGwH0uLD98d9Tl0DKFi5Xp2zl7
ZZD88Jecc9I6g1EV01xiVIklRJsSeWWgVifro9o0mvGCfrxzNXtcTnU4lqvWAYUP
0WK2gaLN0pgsxc4JeEU3b6sz8Xv0kR1YnSFwVHHdjCc9uRLmLYFEDK1lO11LrwKL
GY4cg87wmbwANIlNKSmYUeeoPyUjSrCuKAUi6B1slb1DIPLaltME+jiN+GAW0ZeK
adhFwhHykmce6XqnwTI7u2HyMDniFx5gK+waEoLaE2x/3HwNs9ysfy/usUO28bPS
Jh+KfOUXf1BDG3puIVzyxsrqrauzEMRRZ9TcKokIxWL7SMNfDlr3RiXXhwn1VbYG
02n/iQ2DyMt9sL+RDKL6+RG7QjSeoEr1bqF5GXvp46SBd+X5biLB5AncQJ0DPgwi
nKiqIlnPKdJ5cAo02w2w6R+Uakkzd8IOtO6o5HIsu6upffVLnYPL1ATrOob0FK59
0jedjib5BIZfuhR0joLukZYYlO3eMUxfA/Di1lWZcjMbyLU5OqgZ0fMm1VHInSua
2B76ReaDbvur2OE8hT5ma1JgDDtdoYnRdBAAqFjMqEB1tofSmIexAw/TYEceLxRf
PsD0/nCeAlcit8ngPKeM1ZOd2MVRoZXqrHfaAe70RyQiSpqDa+0eVQ3XA5Joao37
/JqwkLV2Gybr5FjNa5/I7CiFfmQ4QVN92g0fXs+2i+uF6H/zWBbTUK9Bk2xexodD
FXphHjoLEp6nI8GbHTKbsF4qc9Th+hoYnElwgeQzCNU9i/ENr3nMtZXluR5Dm7/F
rCYc6exfmtGAUnrTHBO3Q0TXUycjv3RhtnmQWC2DgJujZhDsc/cUsS/OmOsdQGQT
cKSUOJ9Mo+lsCwL/OqOT8PlDCCvPB32NW0RbJHkJ/JELtysSzH9ORSVxdCsL0qkg
TzZjQi4weJMd9JnU6/bt6G54F7Xo9tb0EWCxcGemQoelvwZc+JmfYGsOb+JhzJSW
AjqprYbm+HuuO1tFVExb7rWTwSplAlLHiFHuBOwXp1E9piCccNfs1lh6xD1vbMLs
SNsqOclJGFOHsz0iuJUROuIQZL7cVXZs7VdPpX5DSvPppcHRGcjezfRTRdc6TN8J
9A5vriss8qhRRASCDbnvjkMZEAgf+6/z0n5RBgVXSEx1yYzGUYlj2c7u2ODOJo1t
6AQPNrEAX0fs4fic2jpdJBuuWpyBCk2Ap23g2GpPbPMbXPZqwW4selbyEYcdken7
l8MyJDNaSMVlmk8pBVf2Hje2GuXuQq3HJgFCthJKy0LBv9sRaSljQNrMLNOHIlHN
n0WI+Y2hm2pqrtYH/P/EYLROh8vfIvTjiPxhQn4ud+liaoCHy09tbuZKq3pwqJM5
0NjHcQmJj8n9D8FtjLxDh6btr7Rx/4yStWcHceRy1bSR8hUhA9dT6rgycDFB/CJr
J6udWCeT+nplXQjR5WctRKkUtJ3m3Dm1O1MC7Seo8c0wlrItPeOjlAyq1rYY+/kt
fHLqcztUMxgQ4d8wSW80hPVnkl96F3n9M7KHiIR2Fp04SJ95lLQLeuG6DGxxsaR5
ltnEWAKiFn1TikEgfTfh4UEE89hHu/2usyeaS9uy+tYf6LTzN4X/uhyr0PFCg5h6
h34YwXiydL9hJ5pbsi3SMyeP5O/ivfHubIvcgz8qJMS5qgNUIPUqtfTgFtxweoUl
e5Y333dlhmjPnRfGuaYCG2oKd582jXm5sfkeaS2ETKXQarX4gVYgmWEQ01ilOhO+
mY7rRr70ruOKARu+TrwgS74fM0SI7oLaMsXuRu+cAcbeM/suE0YyTTzEka9QOl6g
3sS7J8m41DU6Ket2VHdzgpbg71IWYV2vkBApEn/eYu9YEYVLq21LnAVvVqEt341a
zEnEbMS3wgvYbgob3FWfaqEKczbPcNNw6sFcHTY+5K9afRh+OrlkMpM+6ucs8N2a
7j0z/GumtPyTl8DA2Jx/Szon4oMSX0ncuj6MkrURzisOvO0trde9KnpnTowDO2YQ
IMiFQK80AxK4Jf2Uf3rQCP1RHh08vvDIKA1yuvV2H+Ckn0AhhiZEJHaf2dbpmDYC
98I5cRoudtFazkPSvOY7J9gOsvlyNUsuH/sWm1ixhyMjnTq8CLOcCN6q8eGqCF3K
TOk002OwS9THjRZnuqpXF5TJODNMxO+gki9ZpLWyc1oWYVssH5P1EE/Th2tLxrEX
nQxOwzGZqMYf/3JpiCaeISnRjargAxiQwsooX98tEsQBWeqpAX8a5I7Ri2zaOogI
doUsYfsPXpPYzcX24NNb+3Lc8RuWHVZNMvzJVsVVrhlQ7kJ/eCdxPckUMir8+5w1
W9XlViLhDeoHvxr80jTjFLaf5ietdmH14kRhEXdVgl4JPtC+fHopcXJhfqhuVu0i
0rGBB094mZlKG8XmdNUoTwm46CURog94iY6VBq2ZsCHccG7s/ZAnsDEGMIG1+3xn
+30awSfxok/ftWKg+5tvZJwmG0JtQISNPeKxRscbkvRTbZBj6p8s/CZIVKW5j+ob
Rqg4l6DTaAPoGFQOhEF+RAyzNjk8ZLJlFF2LLXcCTzgSbjIwxZl/AEFC/6luvmrO
0/C0WS4LoLeRUszoGVbZyy0rpsccnFHFL9+3C/78zLfqxwx6okNlWOWJsWCsRf7L
mqs9Bo1FVXi1rGyweOgy6lSkGM6i0gxuZVwuxKooDNUywIyceDVhXuilheO51AM0
oHPW0U/p5Vi5dlAT1hO6WzmignZ1sO3rJaO93C2Mn4H3s/n2lM3xKTis9Sgk/iMZ
f4/aKbU6VBYQpW/JcpnKMpMYH656NC1HVJPAzN/AjHl93nzFS6tpBtKZm2ufiuwW
FhCLgeixKGZGiMoAuKOemEM+NksaiGpbblSm2uxgEICbU8IiLshZUTOF+F33l2MV
tDsTPSAPyn9h+UsoDL002QsLw1KNcHH1tyj+v9jLpzlpo9hA5dZ2qdjp8mtUg6zL
Hv/XA8ffNVijSfdUNa9Z0s5kS0o7SevIDDxijSanujgFnYzjhenJvMZDv30i1XYx
uBHOazQv/CDwLXIlpHmnIecajbnXUmN2AAab6/uKVzwjeS2060IX6jpHmdNRCVlg
gbTq8UvzRtHhIzEVTBXOzCB7qIBR3yocPKKqpaFzYJEAXJVO9XoXNuEeMxZmBZ2r
WYkZJAzOkdGc6kIL3g1bb2HQpA6gKWbgttNQLPqK90dEcg3oQNJ9c16xGWzI7t0c
yLgr845+N5N77UtOTX522ivy6veGuj8f7tjxRCAaPAfldgT5nLnrUVX/x6hukXRA
8frtNRcm6e2tKNCQlP+geUCclBuob2biIMslbUyQeii6LDUBdgoK7eE99DSR4SgE
p/5sAparLE/sZZARl8X5+r37ZLwGVSMIB35hvsKK5j8PVMXKskIA1nD9EOfoioa0
ClJXYGjK5hiSUBoAWFOxLklcVt2j4b7AWZxKgjZxhQH2KxdzFrIS2gAFVw+ncWko
fJNB3oXycvSb5IumAv0Cgs3Dzh7+Z90by/Q9x6Ofysf0gHK3tQWKpRhhITpZW7p0
RNS10ER0JmA1/90FDXJm/APXPCES3MB6Q5H/PQzuWjbzeOdVSN9PhxkEN0FykCNW
+Vm4kPJH4k8yMN5OCmt4RlwlkO97xU/1qnt2e4/srdKiAQMQXufuWNxaB8Z54pTe
dKCUb4XwUWOauaCC+Go4Xm0HD+c8TBAVzxezC3zI53W2TnO2uMvUciDiUFBkHkfn
A+wr/9s1hsmu+VGAnc+JPG4ykOEurAX2Kl1jLIymWFxWUZKIA35p66SV0lZVssux
+/67vUaPLB1s0OIWclRoYldCC2QIoBTmc2gBBMV2Xd7ysXlkSFd/fxvBYyb9jbJj
Y8jps6E01l47vpFP6wo47EHTCW79w5w7ZzQyTYrZSCgyZ6magpAg051sml8ZGvzA
RhNx8uzDps7bwzNRZ7a1yNSYxrIm5PKnIDEgGUxji3hMTNUuuehNTfRdoPp92Nvf
dUbWHKJz/7U4gnSjzf4yGbBE25CP2e7MeDLnEQrUETEo3MUjJH/deFOdllo6GoIL
myYW6pba4a6kk1Co7cVBmfOUqBD23gumhQXUUKIq6xSM8v5FlO0QynAAXLuNHWCh
P2hizITuizoOiI3j6DjtX7mtA8O+OZ9x20GfUj/vz2sxJCJX9ADW+IpIRe+iVyYN
fE4+icPN2pfVPHOle4d71DZFW296DZx4BmLwrZE9SWe6rKWxFZvPedOXjoCzaXZg
dSv/sumKm/Ve20+PQvJRjFCrMOUR+KW/YIV9NEArAyw1h57XiSf5f30TB/ZEPzg+
Q6CeWYcQiXzCcZdIzqcTgTTK/W4eZ5O9qOFOYGbnuDDbiDxMGs3m7nPAFOO4Rwcf
0oLEiQW/z9XMRDa7eZKhhKPbbI8FtPKD8n6wzmw9UKFrbTwtPtvuI2tyPt9y6fMG
T/pe+sH6KDMUIl1/vhXl4GfspFgwIZQ32UvTs5RiWVbgCvwAqc9ez9GPSsAsoTyu
uiCWemZ8NMe3M38pSbVC6GZ0gg1gNd7qEJLHaX5v6Kir7iApB44VFTbmV3L74wIT
hEfTcFF5tzBd4OUejK7M4/FWBmGHeL8GHDiIdTfjjc3Z+FM/pH5lP6vKmHeyqXV5
JDW4tergWxXrBh3/y1IIviTrMmyoz7LQVQDzviKxK1ii8qc4+aN1y24a894g6eZy
vapH3wp5qsxMyGt5f816Z+kjBmZUBFshQ3bbiRmLO6ZXmDorfTVFq7MBqqyG3R39
xhUfQ4RKFEaiMmP+XokazI7FVuWzQjUgoiXrSlIf0klGbkWdoofr517CFs8bID0U
hfUvMYezqMKwOiisHBLC/yAx4Iz2Xq34G8vYmrEJeIjTOBtyokV2RjMYXGMELtj8
8oHDD5mPdUbrwhYXHBjfwTEhAzeYT8jdKujhLmqlDSzTj97D5rKNmw0OzkAHcAUg
fNtDtnpacQswfZ4zen/8eHXidqYVMBkfqTZVLs9Y3LrggqClQnAW7n3r/BSboxIV
xi8eDSPMdwbOHSerwmWfboKY09vpGw6OhU766AycUA8A8Db83UClp5GINNt5Ykx1
W97ikqemwARisIz4nuIHN80kGNB8R369oQubcWjFvXc0pAau2V99RpV2G6BZ9Jn9
AK65rf8qYj67g1AFZmHjOjezK85k2/trEeBg3kh5L74J2ESH03QbIz777HDH5uRB
7yMo25Jfk8F5hj/05DgGdagoGqDNf6t4Wuao7/B9dykVXTzBVdMcp4hixT6/tkvj
CBE+tmzIChAuCU2BnofZFQcOS5jzNO1bBjbAxJXTOvvmWRjrX9peYh/Q5V3TCVsc
UOKGp3tf7UVLsg/STmgLwwmNO7corWtBhswB69APfwkMe4IoTGGj/HTLXsgmeCA7
tkns8tVmPE9s11b7mOIscGMIQOZBBmBBZ6M43dZKs3lBcDzIF3YBjEXXBqmfmzs0
lMyPZmSs/LE4ygzeCo9NtRkFb4XByyvCNiaEaVc0XAXAY2OQAUIRsX90B1Pnnr41
r118BD83jYjE8CKB+iuw8IV2cBwvf66ldz0UcunSOJMrPCwt/x9vsbqyCdKWPPem
G3VsCOJ6i/TwaWfhZLCnKcPpk+EBZcDlggUMHfcbxdXHun0cPXQGgEk7MlByoiBd
J09zQDKhUCy2zkdvU3CvodznBxuIEetEQg0sGe8Yx7aCcmiVf1lMeYxgM+b790sR
HgcQCE2lPhl+8IOPevVEsBrtnXzMXvZ2OgfQ8rEIDJE09S1oVQR/Kb1nmkbTIjSt
Oaw6rrA+g88X9Ds1F1anbVPdIM/7GF8vhTt/owwCRNMyXlmmHdo0+DgXE2oTSnYr
JfJYGQGc+HqFXiGBNVxm4lxdUV91XkFP8Xfx5DGigJtkTRCKnM43ZeuzlKLauO2b
vMCB+FIKsBjkWgbbSy+AB9c3H3ntqFXRAuHLiRheXq3cjhx8VdwyjkAx5D/gSLNZ
YQ8wgBGspfIduCVTQwJh/OLj+2MKa0C9f7kd+GcjTH99mxXz6Dd2PL8IJd9vzmMv
A+rVYrOnbE+NLJtHdxsuToJF2UsjIBZwQiUuIn1D/Cat0QagNnCXfTeE94u3KLRW
i87glJ1++oMfe8u4rUtzs6SsyL/pzMfObCvOG7ExJAqcr/DDjnG2rS+Mr3leIOOC
qu327vOARpO14OMKLJOi0b6EY4Qw6e5GLGO9mGnNzcJsJHHMvc30pDyLYMLVAJi/
CUsHFKJl0Wp8pICPldDsc3IW4U2R4PN0NGWAf1OM1hrCPXTo/VCK1X2q8vWM3ZTw
yQpP6hn1DtOLkTE5jekJbjleE/8uIu0qjDjsVJTrK3amn0WBiB1fthlDiEbkGcih
QQoW0HQhOtBnrRtznF2RaBQmvOVVR34/k9L2/QQ6vdwBHBFrCwfHtVcHyReu9a9H
WRc8jMolGgBzLep5u2lUY7P7mNE2XIBZ2ZE+3f4jR7EgOuWb0bE6sA65FPRklZhP
KJl0IEffJmBpOkxyvu+L0pPeHuixpJHBel0BYk7P6MmGGuGBM5zKbZiGe5CoXmuN
PfSDa2ekkADk3GZfwyLmH6QfzfLgspyk8F42ZXHYkaWK+wpmYahuATGxrUVJKSpA
6WRGD7908pIqQY5pCg3hh+oiueFWRNna34PMjZ+J9ZXgTgsn6ZaFPaLtT5AjVotv
vJ0NddWs0IlJWFsKfXbGXQlHWR6NeXjRZ7GQ/g2gO/o9X27pdunAsVQ2aFVPtb8e
6/lqp30aGaEiVsbsW98L8oK7xuLEbCIbgxqnxPbBcNT/1dy7Jz3HsdnYXHdocD2B
rTQ3PVjMpPelRk1xAlenAdCAINl9OdVpwgZyzj8LDM0+d76VI6lo1v4wi9XeBgey
dImkk0uQPaVTM6M1+zZcOxluWd8f759HXKOTd/Y7IomoxZMnEWIhhFkJOhMG/Fvn
3RCVpEMkCCY6ROxhvYAXWt73pE/x/geM5VGzNth/ru5y3aXW5k58jBOSFXdbyDjw
bCzkOVQjefbm71A5Dn62STFojoVnMbVFs7E0UdWClVzSqnNzcSxm2dKsRyf0pzd3
zuLU6jBXndgshESuI2vYechv/TscXarbJWa3VbaE9sxOFXjuVNBYHxw2jyYWqoib
SvcthTzl5Qwa3UWd3tMApaGk2xgFaU/JyHgI9IsAhs/1LH8g6QoJ+j+MCEtD9ljl
dWjL3dyEL+WNWgratFXXT+GcmER6gFFoOEOVpjmDXReIgOh9nTLhtu9zyA2OGwQ9
VOhFsI97SUq30QhqLZChRgIbgp7YHA59kdL9Gw131fG8uicIhcNEbg2tFY4Agdw9
GUjMYi346OTqJnvofUOnHRrAGB12Vlcza/6KlomnfSxfRkpEZVTtmN0v1TDJCYfk
G3tyAUpdwJl6+WG8zdd3yDOAHwF0USu3HEEpjiC13EFkuwOCq16VHpfdppOioIxB
YQKq6nlJv8A8xSnBc6iBd9mqmj2sWWnDmADT3Wn2YzeNsxT/E1gNoN2yCY8ry/pP
m6BoWMKqKxlydHqQv5bt2kbtKl7EY68Y4LxpmInDk6JL/+pKJz8RnomuX67fZGlJ
6oAjfgKk78zUY9O4AiE7fWbCZAPjYccqgIFGRi1AiWmltWSYtmGmw1yf2IR6w1zX
U+S/MsB2cC+Zu+Dd6lRuJ8BN8QsU1pKPM2AvbqW35Np/WWJdz/ybBQLaFeCyduEM
KiSYCkPMQTbEX/JcVuT6SaZvRf3wCsfYJLfuMk6d4QFDcEDJX+oXernpZ+O2Xz1Z
ZV+MD6CnIUO32k6seD36ITAN1T2RddwLJoT/dECSJDxtnRQqC6pdHHn8Tlj6SaJy
6M3B4lGdU8t1sgNLsTktAEdFJLRtA7Svtad38ayUvT36EFAh4GFhwItdEXvML04e
34kXTu5YUFxbs38ugziHlu0C2T0Ya2VRZZiT1Jg1y/PpgYFf12NBQ4XLGFeKEEz6
PbwEO3yt1lZl45cYM2sSwfZALZczzOosBm9VttZNSOeu+MIv65gV3NZSJ1UOpcXz
CXINnBooj1e+DkI8LwFKNPNhejF1HJXcwQlXPzt1y3JBwlvL/wTQj2ybck0Hg234
M46aP9Xq4QPkKaePXEIa3/TgeBm5WSz/+L4wu18rWVDR19DaXLMwXedCdpzoiKTh
uTiO5psTJtLqE4JctH1jhPih0s9uAkFS6/WPXvO20JYehW/+zoAjUxPgCOkONqIR
TJJ396qxx/JktgY/vRn/8NrDbMqfnYDNF59BmTTZbI8XU28hzfJqw8KOUZPrrebl
4s6ol+IKXMIFEsDVeWpTQl6KF2QNlpqe1L5xxuWTKZLKKflWyZdrDBMMeSP1bO1v
gFP++f1IUfylJVoof0kWB/YTuTVVndZVEjBrwBbvbP+Y+BjxDbsgOyPqowv2e85w
IhypAQUFYtFcAckVd7YrdJQxxkTWFg17JmJry8DFywMyAy4VRn8AjsPGsT4kDW3R
GpzHXhlLK7O3TuQwqA5TYjBKh4/Yzn0YgSWQNUpVDoWHBzU50ZzhGBXn/xUiLcIu
wALNlkpwptXJzUfyPaBqKw8lscH6hac+OZ6l2PLCHCkYiLrhMwVFwlKTYThz9cCH
JeZKnd8L750/dMxJHYN2rwRFmTuEbYJaFoZ2KS9ty5pauB3CLLTE/VdRF39cQdnq
48nYT+xUQr+cACAVHTFDFTDAQ0KhZcH66JRJ6CTCwZnYWenQAu3QVyHiZosCCuem
gsfyWgmPABnh1uMLsttpHHyQgF+aUcPy73+UCeIEE43LTcuyaLTWeOADyZbvrKwC
KUiQAZMGLqgHPbgUJJqeS8VMTWEijSxp0rHmD72saA53Ns425tt4rs1NPy0ENJ7T
WkKYIUS6gQwiv4vhkwYHTtLqlIGkm4PmhYJvBC9/PSAUUgwMYgEsP8iKcj4E8cuO
iT2jkk3w3d+zV6sIIjm4iV18C8Ta46H8AFg9RxJdpTI3VGnPIWjnqKM2phK9E9kD
km6xZA6T2Orut2rubf6vpdHWf7ltHd8v8RM6MT8aVLdMxqHef//b0ROv71UOWTpF
Kmq07scSfopsYnoCcWTHTL47Arvgu5a+6HovV0T6HwYTvCUZpvputhYOMjy7BU1q
YbQX7KCDfxVVfF8+vIPWfWKsw3urCWyqUJMpuzG/6ncHM+Nx/BRsFKIReDlNog3R
8fGD6oD9UeuA6K9UBDNLRP9jw/VhBU+5q+o88W91XjxrinpsZrg+of3rSDoaPzPZ
oyxqO7CsT9hhRIkxrlP26tCblXiZMKmUXKBt2FEiiI24ltRs6JwKBIilP2IXRf5p
ukVLALsA0ETA0EK6JcMfses+L9/hxQNI6aSfDuhfWZW4hj+i/pdCk4/ecG10bNKJ
9xs8eHDnYPdjIoON+22c+HZWKcgr2Zn88Z1FL/du3WDwv3YrwpzGQ/g5So8W9XY5
LAcospzp8eF6Sz96LKMZ4PtUToWE/unuPWzeIPbMt2ukzC3BBegnYUoQ1pOdLJJX
RlVWTaSrgMCu3o0jC4H8kXepHKZNyxdSrQImZunNAEdKxMLwmhFMEbwHYjPiYiiw
vZcSzY6lCwIuvSOS/9Ai3/Ih4bEKvvBJL85gcZxTtGGHaUt9NfgEUZ/FU3leAacg
pekiCrsjX/ZUUkJzeVHexzKoHt4GeAsytH4ndQBa9oN8Ucdzqlyibq4TydHiLkpI
ryAr6yoYjBg+wExFuPPt1szlYPu+CmTKzrpLHlzL5qveiJuiOPryaZZKKUVihHnr
6UxFvLbzNMRj5dVzly5hfBvnXQBtP/ofYtw2IMOHYiGWcwWn4a9lmfLWc5TCo1Bi
cPyJdKSDofGWR5E0yz+D3sGgV4vksNOcd/Jh1LXGoiFNA2vbD50tbccjLvGVlFaC
Xb5ogUiKrBGenLqmTNudjMDPwe2dR/HAeSyzBn1aNLX52ch8Pv3Q4scA/fkVbOse
n8SXwdwwI8vCPTX2oTz+meczZ/X+tiKGK6AR0kQvdj2ZiF21r6Vy8UoabwlB1Vrc
8uui98HAKT2WtFdofYiAt/0LcrFpHSSMg2zr+goaDMelLqFVPBakHdLuhlgtKEb9
mzWpi1ardu4L/Xt0xevB/fi4w9D0A8yY1rtxskpjb3dsKn43l9lP6bkdmgNtrr1x
0FvnQxFQKawhcIO/wz6D4hIksJ5rXyQignawZ+SktlNIlh+0i/38Db0Xff9JmiqG
sDB+zuDrJ6WPteaQuKXt9dnY7F5uEMvR9DXfMEFQeFGX7iQoTqFivTA6K2SVsHQH
5EtQFjVjN0vgDROv7fSlAy/0eVt1gJtFaWOcigZXtXr2qNjjO9MbFpQANPp5IXas
XRo3qHDBQaJvnXVhbIwya6tq8Ogm98ksIRAaDuYcPrk2fuDzlWgd4M7cdIjvFNzu
EuK38N/Jo/iRLPyCWxH7u1XO5QeYIs57kR1k8C0n5wUkAbizMOp7UYiIQY4Jh/zy
cSwq6+3I8HbiPrtGa5Bt0cUfsWXiKx6DZtkk/CCYLMuGatkMqmxpc+vOMc3tg47c
ht9YXRJ46TAP3PJHPF9+nEb0ZFdbEHVba9itGCp7GNlMWNxe77KK+wlecI+1wPZO
jElK/stEPkcr91hDXc8ncqJl7rziVLH6z40sF2LH7etITmCpQ5UC2TIcUzcAJnY5
QK1gMyPl2jGfBOqcNqUtZUX/qjlkOWA5LzbchLZUGLMGFEaT95MX0JKOj5f+qAeG
H8eEV8R3Ey0izhKvLtnslBdf7aukcX0KOIrLr9Le5e+67JI/Li46XLpQxltEZyTL
rsk2DlW8A8bVj98pEQZ/LRmsPEc8d6txL5lQbWyjhmFQgb2Fo9o4Qgp5YdVf0UII
h1OHr9A20W1UGAD0GwQdbzoOEvdJ/KNEFcEofsXOeGql+nE2/gHGeYEyfGOf+dKb
iEzGpkCpUvTPGiQz85Ij17VV2hyqOuDdDnzEmxBELInIR53JidEFv6aD2WU2eWKv
6dNCdu1h2wt6t7sVntu9+ePMlexJuigO7pGy4Gyl378HaGH4mEfBmrbbpZxZWUIa
p5BzcxaHzfATf+IQXrrXRL3JkPRtDGPRxAh8VDpX+wpEADckrOze5zaAi+xWMq8f
Fd3szeylEeONI24sHza7OQyaUzrr2bXobfKncJgoxYPqS9bDPo398LJwWjbzbk+6
elMXY0uhTosylyHIEU0XUmZf3HC6epD7LXrHAovmZsbV3eX6SmQLY95wrSA69t3L
Q5Drkxlpgp3Ti7HJkx3udmy2SfrKDcF/4UuHZXs4ZgHpeDU6rbtr6R5PFqGci5UY
zNzn5tZZt6+hxNiYQ06p5D2X8sdgiisy3qn8iTbbrQLKobbBrIZvFR46GdsQMZ/X
QKvUu3kh+0qMJ+z7w1sQaAXoXYF9OmO0sMUgzwIKvcBdO4W2VwzVGp1VLn42fP7D
bUDLXosZ/dASlzIxRA0BdvIIbJaqK1MzjKO7POY0bc9aDr/jWb6ZIeYRsSnfHx4P
fjBXym0eGg4huZKH3qE0GgFB6FeT/TP4uQfg0pbJXMDfTrrUEK9gakljDMQcj3VK
B/xqVgBUH0F5GuPceRTe9fqprZHlfKm/BjcZIBjjTiA+B8ZwXszL/ml7wicWWlHg
L/coVUAHaz3mUO7TwPwTHCFP14mWla6PyGuauEB2u9CgZCRmKXOO2dm27p/MNyiZ
rYfUnZXn2i0XzxOYvfcnWqzE4UJmj6YlgyWN3T3OWMkHAfdKLVf/9gvJPdtHCze5
2aKQjoNyxOdEGWaUbSFg+JwYC8tb2mTILQNUSy7Gtilhtsd7T7qEWYwKll6Vn5VG
7fEmHcE/3gqQ1bL/gV0FIUY76oQimb2U23j7MUloMJmeO/AjTOib/UutGJkzmnZd
jwpIxMJeat493AkPBPBfRo4gvUQpRUnpWFm69b2du14KKDky6Ro9XrrtdNvq+Fqe
hYGma/4r4B6ID4d0vKO7aeQX19u0RrjUpFR7HtSJZm7ScniOL5YVJndaefGhLvw6
tx25h0/VKxRWc/3xcGu9nIOXcUxOa3YXKkmRUBW7mdh5pOkNJcCem1oVpnaQBndB
ljsjW6u09B9yA7+SDSfaDUqHn0nNbKvBUShLNuFz6E00sqKsNPnRQBfuRu9WfFFP
aJ/h5GmHY1pWMrt36w2hZRzUeRaPZMZq0oQ/VwWimWN7Sc4eN7hgLva7TYbJoWqf
Z1SbvbcE8BYW54HumR30pHGVwvRfdNgo5KhZuTtEhsqSIq4hzu196ejVFkZDnorz
T/2o4SeI1p0+XiCAX2gHUnrPbqt+Xd1Ht4yS1oI/dg/MyGu+NI3iP3Ld4pf/59h8
belHZbYovVYN2wr4PhL3xzBPhryreSSn8cptvIpOB3TAHm+FFNauTrTuiiTJy4EL
vwYLmJHhnmMSxbf8WhwJkUTVMDWTRg3zl0xSPnnFXpHUUR0+iBpckuF0/V/XtgCK
VW8yzIQH0hl9ioGJgz1h0L6fzQNHD5W3Vxpb97ABy5LqhuOYL5oGi9NJ9lbxgz/V
9UNzCoiR2UQqD9u7+mtD53g5+BtwMjIupW8t3N3lAoi8ZhyD225xhMIsnczaVzyu
jYvawtnrV/xheAaffIKu8YqrT+Lr4EhIfkukkYuKFoOUcovHmeI4Rk/T36tzlyFD
HVP61rs6cH4Q6ZA0JgUsNJ3+nn29IcECc7wXnmAXmqAaNjXCl8bvB6noO3NZjSi/
S5T34IhFdTZwhd1NwhTiL+ECFkyckoHU9EUeydmp10D3CWkcVPkidatdswJ3oVwP
iYywPMjPqHqHUhCy/kVdGEzf98V54Y6yd9oJnVBhSqyiLC5Q0pUamQS4DaxX6HP3
0Yh3KCVcR0mYsumwAaVmiJXq+NL19mCFcD5f3XE7WEIFS0Kzk+qu3cGeQ5Z8hCeB
R/fML83930anzC4iz4sqTX9l1G4lPfTzFnqxivgeW7SRbM1/PnbukXXq96DGGZ/A
e/l0roT/d9MJsZg8HWwdPCczGwBSyo//Yoph+rRa1Dhb2q8lC8J+kAzYy5QsVT1B
sIOCvyu4QNxpWH2oZX6NeRRihoxzJeMpoGzeaOEd35ExqF2ZKjrX4iI2pb7VupzL
HsKw+/BqO2w15oclpMnuFVFn/kQQt0d329o4kJ90ifqSJ36APjoP6kKcnu5zIvRU
JPFlUTNpBGpJW/RgAkein9I85u9FEoFY1nWRq/76HEAB150b0UZpXIXKWKoS/HTf
aFgtCXnG6sWUwKKOoNerKbVYrSOk6ZCaYqQQKOxd7dLYAPNmGa1JYCfI7S/krmdZ
ipcD3+GoFO5KUxbb8hRSOm5yj7N5ylxmGysGDfaYaFuSnWHlz3W4J9ht1eKGVSO1
GBRSOsZHOeZDV9ffvDbfBHxvTp2yrbTZY5o5iVADIVXf7c4eCFQyBbcRgF3dDLkN
nkwGXPy6IPwXAlzaMVApAI325YOnqQMX/t6Xl3mjXvPUl8OLDJop8T+OPjG25eOl
MUSuMHx8lXtLzCTfiRUnMYYl+MDdaakTGacffiVrE8+SJJs4+keGOWEnJIsLXKEm
c5CVpvhO9KUfOZQuvTmXCPp0K0MJr+aUjeO/C1v47nKaZ7IdLXoDwNlIO5PCqF/Q
MgpYDNa1c+RR3sBk/KOWsqRLYsjSVHTxfzDZCSZ2Zye/lmZ/SK3VKIbzZy0DvoQY
TKQuk6O0BO4dq6WAYXH/A2lm7kx7grU02+7JUphCwGxMnpGy8f9oTc+bqbMQsAZc
IpXGhxIJs/mWBl/LWJ9Y+Q/VgvJ7uSJa9tiPHgrB4RHIJyCrMLHWWr3u8hsqqDsO
l0YKjfbIoByMMG1+s8BqpDnzk31cWVX6cMGQ79+PhNK/yqlB2Pi4pIeJuH8VmHGP
uvhbVhEGbmVBLm8Cs+KZ9eMDEur+Mhm3GGcvbqRAx395PklYKqoDnvOfHkb6PlrI
JfC8xCvVo0fhPyr0pi2HRUU8HkmiZGTMcfOZq6G30oLvtz1JKoLZvc4q2DATOFi6
TD7a0sPFoZz8v+01AVjLC9E1aYr2xTN0M0KRxPvGQUehs3AuPjYLcOaqbgVGSdBO
dlj7kT/OI+/lrdwCO18DZZqNTKYxMHoeSt8MpjlNNbQPxs5lqZL7+1UDcKmPUuzG
4f8KNRJklzpwFtylodTM2eLc8vVMJBaoz66cZz0RakgUsK1ndtDqHWH8V7+iaKfW
GsAxfBOxHK6ZXxOj9EYoCS43WN8UsiPmYM+wT8E4YQ1AS7x3Of+t+QauYswS64fP
JQlm+GEwboDUT+3rSAj+97YlFgRJOqWBg/SWYSFmUQIvOyJ5GtXDY4VrObuTSvTO
NW3p/kuGzA9HBf+3CUH/hcSo2UyCrv3eUAUMasVbnevXgdzDE2OzywRbacAHwpau
j15JlkLFILZJ8sBwb/91jNAnwXThUBYe4QKEjpILT+2rMJHagKH9CuVVDknHKl4q
FKVOldRCm5SkAoUmRVAAnkyOpTAq+TOno6zWxbXRXYcFQQnfQs8l/hLh0LXhzSSs
QtYEJv2Z1tefUeNjmsymgfhbY+5acZ6xl2Ru6DK7YTiEZbwllwQoOMIKC9Kx7CZY
LlJr7wuUXEYzm4EvGxSpinNa+X6b9arL8p27Ufn0fz2viJGotGwF4JhazirUIUZn
UFmqHG083mO/JcDcYkraAV2Euw0rGUO/S1vUCOWRunVtY8YcLL7QHIwbEV1/YggF
UcZWOB9xbDT2uQu1ow31hrY6I7nBTfjtc8Lt6tDqWyMnaMVGfQ16/sFgF7/DBye/
YdGkcrNHZQLsyoKk+C3s9Z+EmLnqmhzs/ftR3NeCpzMPx2GsTB0ObowQVJrLgMJ1
rwj66NJERa5Bqexot0bPFmh1w7XA4v6H2lCPIJY0vq4ggep6xXpWQ3xPw72qE/uh
0IHf47y+UumTKurhPARrPfqzT1MZAzpkYBpHC/6HMM/aDW2bdvXjKF9sV3fjE6du
bS1DiR6r+j2S3ygaari69Gkq+RVp5QEvSjRsUBby7t5roqSsYqTlaBQP2pwre9fE
HO05K+TiJ1Mavqd7hEHUYIL0d2k2vcgo022TumeTYiArXLcFpak+jaxY0xDQK8in
dnBsv4RoKxlfeFzUML6b8H0YK1QDXJ5b0Ykl3ww3CeH7X1SJ7akPAGi0/cF9gpO3
6PU8B9n7a1FWGM8uOyDYfWkKvdsLNr9/v8ev8PBfu41lJi0jfaEaSbc0HAOK33k7
BXPGLZOpGQbCJRWl6/yVtuziHwJ2tGbpGZfanG300kEwkpOeWOYs5QPNf+JimOrs
jFixdL6OZCZ7ED0xKJIqpbhbza0ztLn0CDVueyCQKdSLXfZAuQuJMZ9yAd0dFU9H
ZcUuoS77g+/vhXiekKaDqhjZodkQEvkHwOElVMfWf/cE21L9tbmOmQL1zl/bxfRR
M8Oi+frsGr+zlfvpEgRULEcpc9Q8l/AuVt8yhp1A1Q7z5jGQ7YsimH7jydESvxp8
yGj8klo6rjC7BBCuw+Q+VFzwANHk7eImg1oM1L+0KnpY0kyldrZGQvICZMtXwIEQ
/pWOvam6/rYvEbZptPnIM7ArwqQ/ykIkY/OJOM1ZCnAPSA2rYwx/x54soICfuSfy
r4FtoC6d1bPo4WpPu16Ni33aqUOrCIO1JcLPvo/jxjrqkd4OBE+KB4INSJRbGJVB
c45Ycn2njCEkATHpNz+KS5hgxB7VIrB2EdB2OkEdH56hYZSJks+jL3Ug630fLlmT
8paysr3/DXiCT6oWG6goN5HT1MIEbeEz3sPlhC/WYsZomvd4A0zvPBwpuPUCHV1a
2YH2FVtVlDrhLz7ra5X9iiW5AigOzBe6eKfNpel36FHUe0CzJyNISa+f2vrkDz6H
Yklm3TKawokcSskS0Hw/oQfJF7QRGj8aDLLNEQw0Guy39Qp5MyYixa4xN+F1HkCh
7kajOiMsBImu+1hDW8e2vNELL7gkc78sZn6k7wrm+MEENSkuVioqtogTgNet0XtH
J/vB6VtipZYqrtI28c+CN/QVDkUy1KYNa98lr2zsQz/xNfNF6SyDLyXPc2j18eDk
o9JmwKAM22L3cVp4vjR5cSh5UcIBRwKbqaIiVw8IjkK6DXMp3D78JPIfw1nog2LJ
iLTjRP2g1+scXXKL5o8X51J91rS6BOI/wCaF55Fm+t/2FgeXlrHCV09FjDOsBPWZ
3+ov49nDgLDERgS5PIASpDB5JK0thJx0xCBok1gSQVjhlor6Z7nHqiKz9a9K8VqE
aMCt2GFQTnUkxJMgGTzZNFmZvqGEIbBVNxNW5iIPiQXag/+J0RFPra2MoQimifjd
IKMWSV+oeVjqW/hihS4IUPNu16s3bpW4yoKzOWQr+lgoAwN0unW7TXsgARzJuhUk
Sqmlv18OMyzFXq3HrWxvCTw1vpDiiXIjv+jUgIZWyoCU/HeOuj7a9YVwjqERkKdM
bf+elVaTKBKKFRa8p6+BGLTlKS07h9N+v9G3pkzVeTh9z1gkWQcGTQ9x0+cNI4qS
tANgwS4b+K82hkRoZFDrmjcB9NrsUefzWSbT71msk7jcamSzhCadFfWd+Yco5xQ/
DUDvTv44CeCn2CEMH0HZIr1DOFqqU3M8vFKhxOcQj0JRSXKuAQlXvpmIGwRVT9uJ
KqxznLjVzdQORedyx9+bMc9l/bwRjOISdv6o2AqB+brvz5iydHuLgWET8rfk++Kz
tK4w18C4VT03R5BiWBhnhoSDeKjJTXS43/grjGdA/8v9Aih2U3aos6zzDmgEx1QI
pReOwHJX8nyJcJR/cvo+VhkK4bFyVsFxggIcRRsfPBas9MMjpHldw+NmOdgIrih+
BwpjDnfm7O/iwrvSukp0U0WznX1m2PRVcAEOjuW5nEDnngnn7Nb65zuu9VtfmM1B
bcdUa19KXaClTDQwvcPbrfJCTBQl54dOmiBEG2jrOXvnwqd/S3grwTnoCH2qPYYF
SBxyyTJ9xnScfX7xfhudkrjygIspk2fPztLfgjPh9d7IQ2NJHxglTIIqoEC9eLoM
udxatMOeqzSRjFpkLxjUY+yb9ixOZ6kr1BCUmQtJQKULS0dckRkavZ9dnjzjDTSW
zukJnc8yvqgaEzNHC15ZU41xuvQTGCO7bS1GXlWn7VAgyPrKkbe0vqhn3acjwg5y
So9/WAc9/xPfJsRm5UYnYXmkWH6Kqsyb4vdAZjRZVO8Z+rIhW8DmFSe68Lj+IA5w
bX0X/OIqCQU8fy6bnyXHCpVO5ag58SaqvgTEVUbYhIPzYX6YAKoqxsidLWcshfVD
ghVYj9MhQT+XaZV73L1ytOnsDgisERso3haGD+qB896equoCSHUoAft/F1HFjnei
tGxOFaChWbsXuKGGOPUaaaM4evyq/IiGfLfyEKQS+BdKj55VHSEBGKISY/qm8QKI
okfGp8YpMLc3AABG8CeGMZPGJHDDfEA3Q4P48ey7Nq2Vwx7lR2MsPD8XmE4+VpQI
0w1lAGKt2VWQ/Phh4jmRAx/3RqnuGMXL46rIohxsriISuEGWsSv/EyMr9iLZizms
V6nN0cj5tr8ZImxPbsZozbt+wM9ximoOZZ/FjLcjwouOj4WTTXlDHzYoGYAxUQ/4
bKsZR6ZcDSR6o2MbuRs8HNwtAHMrsu0B7GlGez9w9w/KkIvHJUW5s7g1VjyGWmFN
zYHDiwUnAnFeeOzXojfu2b7UtAIqdc2nSLisS3YQ7xVamkhIvueGEDtZWw3ez7hR
ZXll6SK4mafRVnYV6AhYpWtQcDxBips1TQeCBnq/TgTgE0Q2S0HuQS1ZKTLjX3XU
7eQRyFW4savU0V4fPn7Qfu0OiB/eE8JyKG98z+wmMSK3bRyXn/JxkPiwnQvwlhKg
8vq15phspJscyofTQMCYa5gXuISa59K7hQaTPBJygyCdrnEb4A66e/Ivbz4pdIlm
5eYZR2CcWNg8yTX3ZOxwhr/4NmdAHVNSAXvSuzo2ku1P7F53EV2HEU2PlNhbLK13
OjnnTgXv24/yVI2sEkBsuA2Phz3OdcEj/1dVpRFsxYrIjRmt9iq09ZhQWyVCtZYa
soSYZSvm+K8N72UZ0Sda5784sbBnygP7R+ao16qNkolaKnm7Gsf34rjjWwZdQYIy
o15yNpmR2FXf0sysoezX2mhI4hHbxEsXsEGMnRSN00BziLbQS+QRVY/pFJoPiJep
6+wFOKny4N3GvEL+NbEqN8qKGMg+YSp6RPpL5xA47xOom7gZFS55R7EktGP7x4z5
sTmzY26+8+JOvbo3hTkWUrkpC+T4Lxec0bq4MIy/qPzm14la8buZny8SQhXrRRQG
Hp+l2JWBSQ2AtqqNUWZU1Al6SFti+bAjHBjE53ttoIC3tvbCMfCTCetl4m9pRty4
ym4fsmT4ntTjp2IkdHp/hQObSrpUAZ4yz0TLcYezOgh897i/voUl3HAU2cFiBewo
JwG41Mpag2sSTLuoaXUwSxQM90MZYq9xo0rCzXiqd1UNuzQFvXcBopNVbLbVAT2J
W2vA3ZOYGIbBadLmcfdK0tF8Liz+yFOZ8B1bC5ExupE4oIZWLBf2KyRaFnTQKBj5
fZ5oolboOB06KLQ73vrRuf3n+LCX2WTkaugi5ccCvt0dh52aM94m+g7YdJ6btqH2
3sdykU190n5/nXL9tMvD2hD3CuCPnJDSHXDVqD7PNsUsWetJJBJ7GNxCAIo76iQF
+8ymQG+fRGQ8/cEjgNC5xOHLnORuVkBH7ltoPx2exnX9+6csA2jHUfowxClMbWFQ
4HEUkuYDOISxbZfTEDwM6ev2qZEEg9HKQBMbYnNY3QASmWTN4idNiVkd36EpfeBh
VQ71fkScHMwI3tBAaZtW6v/M0vDkizpw/Ov25NcoG/QtGc+AOZHC8JM5pMJp92Yq
xG0t+2fG5OjH9aEXN88TLTH/mu2KKDezK+Pmqr4g011PLdW80M9HAb9xqgtFOs4Q
Fl8ZqmbuPZtmjVxwwCmhlGlv4WTIEOnaR+dUN+Ejqo3wPstUVc1bPMXx1pl370n4
xCbyWTU1nEnhNVnCL38C0pxVGVeWhAP3qj89LsigvwaNBhPveWm5NemYBw+pKxqk
s6HBkcY2LpJMjmVxjfqQtu6GQsmfc61Cssdq10yZDgpkDK5DiWZDlxFoByMYwuqG
L/9FWEVa7FRwb0buWp7G694HbR0yVp+Fj/radhcvRvP8yt0cxYOoJu03xN6/jkDx
T9hHognfVtM+qEwNd8CLkmxr6K6BLPh37QDVO0bGK9PRFUT1Gw9pw4bCtSH8gpYO
EaO6fARuITvnYLEaVPJEF/ffOUmG4cldsIrIIfT6HRbmBoNIbznud+qoBmAQLyHw
hWgVu0dzE5d+OPYG+aCN6AD5nBBKGKdHocyeBpSh60Pt56yn0RZWjGJyqmuxz11u
9Ret2Asx0PgkPjzJCPOqYAoGkN960/tDTvcw7ZZGVZ/o0m0hNXMUWbFvDOOMZ2JJ
rFvBcSecPCcF/766Vntl9Q3TGh6Q2lozmippoHOl9N5uSZXc63CpPnJqJ7wLUF9m
AUBNj6LdcECg2/ONADFoC1yEdHxd/EGJnV9MN+/s/CSjuU1cm8tAtjeLeGdrBstr
pmc8QAIr4tBxeRjqaPQplXBdQwnCFN3/NMz42mIggeM83kIByh4830clZawnLaFW
hgzny7IfWsV7L55o82Ninj8D2gQsPQRQHWFL4p0B16y4HpPIngWY8V8QBrYlihp9
kw9I4xnxz4jU28ZTpij2Tsj6t/8jYt/jNiDchWLLioCqrs3QvH66tijbdkdd6qI5
24od+43/JpxNIXSiP3NAZl3MnT3CTfzOUaqS2nYXi/lml0Z04+6mjx3ss6hm5leo
Gpo8VhWmjA/1s4iy50QQdjGlmyTNU3ry5JqwXCyrwyEurkngDxFhrMsTw+w0wBhM
KzOOeHCRXMdjk+0jLNkhQsEclpNUWHR+dIFuFvMFzDPVZFV4EIeJDgEOCKtcLAzY
FGz6FayyZjGzVQ875KULMCihQ35/8z/4iVeOSVegGeYwxIlPPelvSuuZyGAojQey
B5gnaPI3ZKcKOPkvmeXHBDelRtb8kqmSQqq1ZhDWV0NySAwb10p8YbLpIjmPHYyR
DEs9+Um08v3XZs15+k1/WR6zzjon4O3EvkZAkEjcXts37ygxgLCFPJSVpta2oIjl
k67EeH54p8HZ2+8w1ihFPivxiSo0nWOfNW++Ia2QB5Sz2PQqQpYdRU3SipvIj7Lv
CGg0GwKTfYZbOZK7bQUe1FRn5bhXmzVr37RJHXnYRl/731XzpEV9UEJ6nCsG+caC
plewH59lfHdr3jc8VHLpzDkZyegJgL+e0mHKzbyIZEZzytVR/BZz0j5X7gMutkk4
Fw2lglKxOChVFxSin76aViqfPy2nswvlvWytNs+RkutyFZFJSdvaVVmsschDPbrF
PIr3PtOsKr9PGKXAqjNt5j4BKXDOt2iIfiGbnCqGk3tTQwBidXsPZmrHLTAk0v0Y
tyEWSWvnVVOm852yVz/PHFHFoNX4fBli+aDgMzknKwVW4+UDesKLPa7gr2diIeKa
7pzgfRh1slGsplD08ic00XTCksBuAfEPfJvvaQmhgV9CM7XHCGHYfdX4fK/690lO
y3MACnKwZpR9js52F/Bpy2/nFKlOZpYTXAnAvrDCdcjT2BAeYKr0lX3rxAHMzFBS
mX0Wetvf1cNoXIdj+dfAcR4fGfNs4OLF3UgFDvoQamu9CSniRQdMcsvUBOPK5+Ks
Rc9T1vNkVqPNKd/bW4wo63Y89sp1ZvJM9TgHXVq+KzJYxzqVbbPG940tNmQKokdt
UaQDimr29VsWdFgDoBo08pkDJeebip71db2AyIkK/LunT16eMoA0X2OnxL83Rhia
kyYr/EYAhgX6ntZGWnipBKRZqlOMn1uVCwsnOXVZnQ66ruPanQfjn3PU0CqVT6TO
B7LIVyF+m8HOv5RlIslN5dBdBgco2i4e1p3DVnKRZxP9iBfIrVB0Qk4yHiRx4VTm
poLTvCGFuQCqvOakT6i009pB+NWUpaNUU5B+ZLQiBcStLa6HJyvzRqdDgEIh3jq/
cJEBeiHpqCRbQj8O1ND+ZgWQVqzeaHtJsW/yb8dK3rywMaOa6IJapmQdvzRaMyxB
zqHuxQHM5JdN/XDqc8wzaAUZYVx5uMaQyby82j/3m195mbUAhT9b4+nd0P3TMvSW
7Il6vcK74jnPz8yIow9J+xK4UUcK37CxZyRR5djugrqERkdNWsrgaoIP+d8DiIST
784M7XLjdJbRI2ydrB1Jy5y+IBHmUrv4+0+lIujEYCTIYplTEBeCm/QXcICIKhZV
xleZsQAT7LOHSgXHlJ+NhBRfq5mDVqlK1D8OA4lpKDpvNZnURXZJjg4TtfP7goU4
cQf172lw+fYY4kbiFAeRDMjQSmJ15gRD3Qnc/dwUHdvOj4uwzzsZerchuimp1nHo
iACyxqBXCXsHhJmif+xm5LNmzYJrp9yFJ0WnRvF1qjrvnkPyS9O2DfnZnTr7bHiQ
TBSknS5cBnkkWpBOrWw3mlzSG164aH9TM33VrUrQLS9fmHFhk9wbM5evc8s1btn5
I1CG/B7zjVEzws3mMk7oMh+tIp9zgb9JHWxp3BFNqBn+ySlCp7PiR9h20rpZ8T7J
SrUIldZHDwEQfgjptw73aKKaifyOuy0ST8pSWcy777m9Andtk694fiIqo8Id7wCV
w2KPJXp7HtJMM774bqsyPPWgsULs9gkL0H90egBdKHGcY+wqQRLl1gvWxhj6QbEk
eqjc7ToeOn7XpGgP6pIgyRoBGKeQ7dLhkmgDEhdtlhUQPKlOHVuwLmW9It8Mf2vi
+0CrkIMHZEvfgzmUrL8Voo7B/YLOQ7reNzmC5XxRxNkUp86YuLz9WkeS2OpPequ0
i11UXiNf+twL4xXi0AHs0elxVQEXTJbvrVb7jiMFcwNj96y0YzamCzCSBUahtbc/
U9DVAuvfkbUb8WECaqRUnSwc/MvM7fFJ3VP8Kr7MzhESJXNZHosDadMlCqwPQGMh
xO6uRkfmgm3aChDE8JqTGxsDNG25U2vb1miD1POCncT3ZoxetgfNsd+MSW5ewGvC
APZLisFqV2VyVW/oXv7nlqvfLk8y3e6E0KCVof3kN0S9GtjTzExN7gHBJ4pU+bVT
MZcZc0xe7YYHMXB36wxvFkG7PbK6R9aj9Sk6dkHFdtDauHkPuXWxBbW5ok7BCFjT
n1OM5KuESI1jIAQaDNXAXp9KlV/2Yt882SoRDZFp9kNw12hjN+/pFx2qoQ6gWb0x
NujZJ6FaK+SrmsKf63H1ineK13mq2drsaTPsbRDGIN13+6nzW0+rTRzCweivy/8/
7gP1lrO9c1JHiyWaO3HuaFGZpBa9btOVsjT+4baHvNGVcUmY5HkBU0KXiQ2CLO4g
WkiVXs1H58VkT9x/m6yBmrbKSH9O1rpLhcJTKkxBDhijjJdZlD6XK4OvGKai8qe+
sE5v0sC10k8ZkQZdBf2lQ+iHL2uktcW25vJcD5XEgyLjCSaR6bhGUuLXfyAodiCA
QWHhJw6XMyc1Gnuj7/YzjbOcAl9G8/9XkjDIjeARDyzFkQ6E1G4zuLSk8Aef9Cgc
K4YRhlN7Ng7XPFgm/knmZY+yB3dom6nWgQB5G1i0xMHsc4w4ZtOIX6YLm9Ibl0Rp
uDHC4KYhh8RrjxuzAsAhBn924vt4ilDRcO0O+5ZpE23buNeGqttT6a+wCuycjRfj
ghLfBK3hPWPClKZ2qHM50hvfoA+nvGwFK5bURnYnJf14+amjTg4ermGYle243alO
oiqs2xtVmMc97kiPayFxd10CYJ2e6w5sLzZoIFQGDzZItc6lpmzsUvp1HfLzf2XN
VQ6T+qvitZ47Xe3/4jLLbE1ILzEU19cbBiFbyE2sWU8CIe5AgJbeJjDfA3Q2T63E
QVgQEvNb21tF6MZAmWu98HEL3epLzz1jwbseGzJmjM5zsTZz/RbStyXSXH37JD+g
X9XNovB3iIZJQRDAAncYR/uJvB0G15GOAumF36rZrvgPLuIc9vGXBETshqXHsRTf
BeE5cyRGK7ft5Ba3Sv5BAn9d0+9++18L9urlldjD4e5zsNqMW4IfigyM1h73hdsJ
P3e31lVKJIFp/CNVOUmYpjWP0sHIY/eXqbL9/aNW2uIJ1QxHB+87iIa16M0mGLsD
MO7vjtqB4BA5Ijbrw9JBNOBE0gjrxUG5B2yjHQD55koHvSxNJ4JyfL1g14LiJwzV
/tYXTAbekCcPkLsAomXfbFPnns4sDYOWmzBGuAw6HCZ47Bw7ERwg9iPekhZfasod
hj64snTsbzyPejrWDqc+DuYv67WWhIGeJaLlPkP8pQxRCTX5Yg3hp+rBQEPoU1Dj
FxIg6mZPhVtH8N0ufXP80k3q0+8Mtz87HClHJIBOwcYLJ1V6BeUKMA24CEEUhONY
5jzCoKs/XOiZyX/IZRdrsDHpi8SuPqSnXvQIeUoY9VEg6HIzCD+QBTVRq2cOjx+y
RF0IOlvU70uJOAiWp/1+2kjBfjVZSgZVnmzNJUOqYXX1R+GBmzXzcZSSloYPodFd
A5/kH/6spXXrsxH5bWboneUIyFHTPkNtjJoXAHEDfhhYa06RQrU9nIzBxOo9mQhd
qcXjs6GtZTU76eA1RdQPVSmH6xEwOlti2wV/4UbYVoGCDE/Ti5tCC1d6B26o3IH1
mtnYRiC77aGUGveIjTwHXOObD733f9uQFSqIGUOsA/49LL+7idJXE0vXWMQr4Y+i
f+HIO2h3ZdWAWViIcmlLOMGGeM7TkIndpymiV3e1WLT/3DmUWzHv8g7FeVPTIU94
BUeigZK8I3qe/GSwsV9Y6WLJIsyeCT6nbAD4yvzHNfpudSKdJOSteM8qG9hNxA4/
X0zPNnTjCf9MxnKq0cq0UdzssC/g73KercuAoOr6iN//k1E4AzXH9lb46u7jF+QW
bTsekqH7wuVoczbYo06tpa3A/Z8YUZpSIYoPNx4+Bvk/ydoFi6JxkNjS4SApPSLO
Hox8rTKcjp4Yuu6FgDkAIHRPXHyvjzyjKirD3qpG6x05zn4G9tLl285Wqjbp12Hl
6I6KZSyoYPJgLLbtOaxqTKA98yzqaFWtINQNnYEXiXQLEz3bShA8XPxUBJHEnBoR
G+tARxDu2WInFT/Boeb+pYzXzfVUq1dkjpGVNXKKfaErFjA+F5yOsu5ybIllssFL
MxkNiW1OwEmCQhzImbnOeiHAXf25QiB7NhUJAenHCqlxMeckwgbuEVGBtnXD+bOD
BdYSbdUc89+qOFSplngWAmu33WZId5F1Ay+eLexvGEiLp4BeUJuXjqH4RQ3DCWfc
HnkTepTfCWclFWu1m+o2lxF0eHbSCadM7JJcJiWm16ou2w4mZM4VipntsocGSUnI
pee99KcPpyLV6cS70eJ0HBMI8cigUzEfdi2QuSZc4Pip+Ug8AEYLx/Kfzn3e4lxl
XxSeAuWtp313L3OhXS2iPxhWeSN54lZOoTEwHUiQCihohoAs0CJZ5h3mxYee6thF
kCjuxixNH/wRIFqrRhIN4+Z++2efthoov+lZ/AM9oC6kAqVWbx9E15wZn0BVYQ0Q
KXlzGDSWvqN8UHSBBgjeZ8e+N0Px+U6UnHRF1Dufe+iy4MBqSqe+URGSr3qkg6p9
WPHwpcNnvzgbubTjmTmFQNTF6XU2maO4wTWarXVlZZB0MhF8zWzpugwO5htrpenR
dP89ghB4M9YfagM9YqqMWfhKfd8GpxFdLeRrpa7aPWEX9OH3BLEru+W0Tr8lNoYq
lEL2TnK6FsB0IFKVXsiNpLpxte27dqNQcBFaZ7j1Ft5Tfc5LuJ6cYZWLuj3ReL6l
TCw+l6iBotn8MS4DGX8zDU6fM+sTVFpebFHv+aDskmgAr4qTyXaaEXlHStHbCD4v
B79x5eDmH48wCGv84Rz861qgpT52vliJ8nwYlELBelWJ4hMI+QlwI2VDdWz5hQBB
tdJjmSNbLj5nYV4yegxu6w1nrJeir9Kt60aJtBQfONHv8BFZEXK0mYk8EDMxLfHe
6B3agCknIbsLJb1YRKN3uYHAEwj8WWTPLVVsILkiLGVJyrR6RRg7XnkCxdVGKfSo
+VBitdcJ1NCENh4VKKfVlJ6Ns4PUnplFx7ZI6g0sn+Cd2ZB5ZZpvmyKpMES4ixn1
B5uvtbVLyLKgK04CkovWzmD8EUtbIpGC9zFGHDYKkRDjQY2NooXZoNfe6KczhRBH
cv68AN471YQQFR+deAuVAs/b0AO9Ph21+DwIgIkfofKVbgnzrmcRkAa++9BPxzVp
54HVq5Ex5g3UL0CYjZlmr0PCMbSkD4n8l8b7PGv735c5FZ8FjWDorbGOB69Stlt5
zOmWTn+U9qHW4v0XslU6mEKrRDZnF/qMtD2Mlfl6KXWLguwEzpj5tfct38/FpqGD
XY5yfILTkkq2BlGzZ+sUUyp8zXcLN+6myYx9qWkRUUAT51IPhEsKZJ5FT9INnUwy
f8IL11pjc7Nq5S3bbXn/tGYjgVw4o04nstT90JDSwyAfmq4z8NrBeNEhHgsmghAD
6w75U0qh+zvLiu0EyIXBqYmNunhxu0sYTMVlAK9CaguY9jCZBVb9aTK7c0Go8mf9
Mh6nOl6ZymVgT06cEHOKTSOFXqtg3Pxzzn8+5db958QUAGbD5+Ui7MGJNwuA+uqm
s5LHuDM98wfcpuAz0CIz+D0wpcyeACsOUg0vCZmnBnVqb9FfXnRyD6iraj7HsD5n
TCTKkZ3EAeq602SY6op49jiz/8jgMsY/zb/zh2Q3CTleUS5k7/mCHcM+KeYji+Pg
HUfeKSs2Ooh/iPsf1CnApS/IGRYKBCRjQRTZJ9mR0mjAdvYlcRY3biM3XC4w3aKJ
eEobSqLknQRqP4HfDVgk6VedoUGwPLiV6EB8jxXlHr0TZzSNcvaYUjuok9UDM1uz
ixuSoln2+UcpHmQ2X+tfkaCN97yA7J/koNKkSjynacuzU9HTQcvaZ5Bz+sK0q2fe
K339EOg15mYpcY5AYLDcPbyCCwUkedk3std1xwlVWfoqiu+9FrS2Cbn6AXN5fDNP
xSzHkbGy/1l3Ma1nNwfQv6/qipZ4M7k6lzJNnrGgoaDMXO69d1m9FrwKKxw8kBa7
owEiRFKN0Lgs7d71t2L/GUq3EWEnLaX5iqVUBOdkBBHsJ5Y5wSi23aYtFS5ui9JZ
C42b7YVRGowSBLOeNBMBk3waP4FvDXNLaVWuWDbATcWNliJ4/UW3rrQWjLyVm3gV
L4uyLSnIkZ/7UN5C5sPtj9IK9b5DGD0yE82Z69C9JfECO6QD3Fu056E1wRAHGyLl
SquOmWnwaGK3tSkjwRIgm4YiFi+hvH7YWx/Emb5g+yP5TrY7SnwItWOUCgOz0BYc
gVEo9gRkPSAEJTlPvAwwJzi1lWQc/VSdumBPo6Gt5qVBZYoGwpbdlGdvWnCKidsI
xVdM6uyPnzZMPkO5FSvw/uBBooEc6F6G7t/nZjEPS4/0A8WZt2n32KnXVS5ccRP4
jmEOrFWXgu09p6VUCQdFzPxIripxnm8X1oXvacM3OAv/n5nM1T+WFoYq7/Gs7rft
CmMAzmw0xKBk7YSBQMSD2Tnj5TYDRUqOdvVH42G0KnPt33gHtAXQ1jkIiapCfSMK
udkY9Doa/mwBkmPTHSShvFWqGPNZ1qfu2thnjpbdLrkmof7168WK1aUy+QfE+F9h
dEOg7F32LJZ5eZr64fyRGXATrwiUnM5R6Pmlx0tPNwgRkliAy5FtQrv46kPcUdh/
T1Nlbhh7x8isn07pSdumHOAd2d/R58NXkDGcOBT0HIRvU7B4woX5uUN1LE0v/4hw
NR0tcY2pGQ468i7rbuZfPFXoETqdXhEj83exQI4GLmA9dDmQ2ha7ucvz9UA06F8K
EApoLiXTf2IayGCDgi/3Dc7GRHu19OKBYMPvLX4blS2GwkxBkXcsrSjVsr6RLXXp
Y7NIfrx9aLNnRsrbSFqB99Zr3FeR1HKQkJBqFBzWLbQLCC/q86sgxzSkspCvFUBQ
rnD5KDWocq6PQkeT9+ZBke6WyuuC3lkzZUoV3RCj3i8PsqbNevzBjLtxZDXByYxH
AMB8W5x9e4gb/xfjgX1tIlvSFomhyxhdCtdN0tLyr/QYa+Fv/iZl/rBwFbWIvmRv
GzfD/5sFD578bfOi4Slq3hllRgqLMu0xYDg4kPqHuOB8uT/D3xdMoe8+SAHxTT2q
J6qhu+y0peaGzDesoq9yxT2c3ScF2xzRXsIYiEa2PmPN2b9ggRth9zIOZPKEzjT+
3aqWmjHLj1OhQPMYT5bFMhqlS7Z6RtqhSRNe6HnoFsF5uRqy9qhpboE7wMRu2szX
qd3TPBsXxpBiZdAa1QFF7EKAMb2BMWZU1HprdM43dvi8sE1bRpqadM9jI0CbiHiI
m7Wz2EO1UVPDT+IwPyCgwCJfu/Dlzc3kKMSBZTiYmlaxa/YkNeIpGoWGe4T+WEAx
vlotIDYJebURtVmFftG5TT0gxWR9PsVKCs8gX/vsDXKbBnyN2emYHqm2iB7bPBrG
rbmqewURWBt0Ua385+cJK+gm9oV4S9JJAnk03Ww6TVR+6UH8BgfQINHi1Smq3R9+
uApkR9MOdK3D1yR3fkDJVOEo4cHIDydEeTsCsqWlpCk/j9GOqm/fRiaVbKAAUXlF
DQJTYyhvQBZhvVLLa/8pT9cflUC3qnG6qxZIEIJYQHcHIpv5Tq7ulBtIYDHipA0Y
1h2tdAg8twiqKsAzkLAl9NBuNF3aPo03TeWVOoRiDr8eYNZvIqt5yIkJ6bZC4+JF
vf6+XXsKXb+QaqZj1KGzj/3gItA5phhge99hYGPcwdXoI2C/FoBXZlnXK6PPNZwx
lHTeWkZad/G1hxkrHn9J/hteX8EeGIP42gBkxssrAVl4HC2fD3OPegrkRih0T+SU
wm2b0qzkEw/93nT8fevDiwhBSCufhkINw5MDG3Fz5W48XTqiSIazJE/oArHNThky
FE7AKyT/rdJeQ7lmKa28ptdFj/1JBi1bz/GUdSNjE6oEIyq7y+fqCNnQ5y866iVm
d1mAwrm5KzGIbwcQw5C7K7L6LL/zk/cvuzi37QCI8YrlAu0RZUdT6bSkd5IZLXX6
bTO9DgNz6Qk2hqc2Kn4QTDqYf1FV3xk07FTJGnRBhSrN9/r+Is6iHFiEE87AR6wC
6DvHeCCAn0qaifVq/gg6ZIBIITv6qwdiA8JDVQurkq/r9Far/EyYZJto2XvpG6+x
BD6kVOuFG+Z4L1kGwMJ4CDuihAmZVRUz56HAKzHORCX9ydZ9DhBw8YaZThWEf7BE
S3dZyfvI7m1xXSWaXQRvz/jfSVbRJURxTC9CbxzcoK3BeOfI7ReRGsJl5JLfMqEz
CI0ugQzgd3qtQJrsdnyK8hyfJObKi7zKfNn5NoosvLl4bkrct88yFUEzUZR1ArSf
nZWnHX/tvKpbRV5jG5NmW6zufsN4+dKq3NKCcFqfAmgKiEXN2vYMS1b8Ia5KUirX
l1XUOXFZQe8GZ/cDS4CXah/5ajj+Tprk1UUomZNcACPPAfr16P1PKb7mujZN2dpz
zx3R9q3fGdQ6vY0bWc7iwMq83VLNtITBPXfZMFBhvtT7GDLRs2U2te8eInXcMU9R
PIB09QqGWNiTI4fAMw1eNNAqckzAgmmRzrIBDptC79/L+MAH3zy4hmxvIMgLr8DJ
4cLBHmxlW+Uybj5f/lu6PjflUFn2ZgGscXm3odFe3xnxg80GpFI0X2afHEIXCOJM
HyKN+6nDTeDYfZVWpy/5nVtVkI9SSoTHu0RTei8snz89hMULNgQG66cAubNq9c7H
CBHhl+RctPsnTwtiS/tKv5lMsvdjWPPTH4km5y+FEo7u+tvnD1fUhU6NH4JaeiTe
B01joovn5oWcWCGFdVZZNzWLzYYpo5YQiHjKKP4G3av3rhuN3ymuVksctA0+fIM8
GCpMs0TzW/qETQ9sLncKsB9ZN2ukPUR5tQXC7wE2rzrXx3fndbldT/31T1JcG+MO
VfMmLFSHFCX3OdoPzkNRcI1gHINTWu9wN4iE1+/YAJflwxuZcgqOWTTDbEdUO6Jh
HO6mHImn/1znnrWuXephLpHUV2bxAXo87W+2/AmXCe17FZi74ksz/+nTuqvdHZsg
oiGw8jI6/Lm4iq438miqqHT410gJ1sp8d/hrOIqcwg064m7EKjyqb/yao8KYH/uP
LWCevK0wrMLOvcwWSVhTgK0b4faFsyt50fbC3K3m3cPIGUQWnjARNekC4i/z1JIN
NA/Xoll3NpfpbOIe5/Kc2R2NU/fejWqlnQJmHkQvQ5zS2nGOc68+1eecbdlMyQCO
veABN22OjEK638RZgxpirG0dceaQa+a5xKU4rDqA0PVObVZqZZ0ozNWvOFh9yhlu
RzW+d5/Ym9C7YPeZrgOEVc/S9Ak9FDBDyQNdrnJtnKIK1CtYsjQtGTnA6OCxnE8r
6jHSTYoxIJTouTedMx4ESz43LUJEBFKJN1TU1eI4/SlADol1l1o4u1hsFIrqvfNn
VBvuowtAB7gX5F0feca664ZqJ3bZ7+mHIn2of0zP1EDslTm4rrB+auZgFo5DHq5n
oSbDV1/BgWMLECfgyw49p1MxdPq/wwV8QS1XTwA0sToueVPTPl0oZwqiKKsR8sRz
TEGt+rsef43LlmY4T0g/8WvfZYJcNcjTOd+Mj8TrfM/QFsuW0Y/Es3v2Ywj7s4sz
NkMeN6nfcVBfY0wtjpmiuBtW3gJjj+6tkv3TsE6IOXyAx+lm38LfXT0s3AkSXkK1
umex7D1KzeH01gOPFno/GYZgJgYuGYNdXQViFXLaJQe/CoiaV4O69+8EvnXkMXq6
XPRwszmiegRlMKwKHd61fXsVZStgQkE9Z2oyE4nttiUGAS+x5KS+H7SB4jnM4o0q
BNk3hCUTNrtUCyvdbpQKuDuixcOATiLiERzqDL4pkqW8SqvSEUEhs1Zfawioe+mJ
hKzL7kBCT45DP+bB1ptrkKTG4NDFEFbKZ4DLjbDQ+j4UAHVIGhwC0Z6sw5tDLhJH
zuGbxvypeYelffUg5J4diNoGgXbtT+hSnGuyKN1W5pk2BnrZbiaxfRDjjNbVKI0g
DXLNkhQT5lh4GrPvB1oEoE0ddSs59js9UL/1ZGAgPjNZhjV/H/XZqS1Er6HLycP5
bBzFNxTDqHrwk/eIz+HmEblWwuuXPBsPpXapHnMRuOOSlK0v6tMOcfOhHZCPwwb9
ejHG4VgLHdzdNA2wFDE+nhhFLr9arNcOxEkF6CZ6yU2vmm8H4ypuTxr65jq4Ipy2
/Slz6jDGn3XZsmucvkN11Ju6ylPDNt/qxIPO5rqDZb1rQVFarFU+ofg6bj9uuot0
aot8Mq7oXayAVoXd5tK1XjNp+YZoDRO7HGo1zKZNLCKU56FviBgKvtx94DpaPcQ+
NDdpVR3s2wpo3oewmpEsTrGdMoaANq9WqiKuUAZPnxf0ganbG7wd6LhYpPgTEUbh
Y12d6jocswT5vV6gpkKAd9CXeffcxnTEzYRv5NP4Pg/wf8aJVjr3gIcD4tEvjw3h
bSunBjC03n8Ast+VkPMTBBUC2p31wVdGg90OWcbuIEeSGIsdXNEem38PjACmlLxp
LQTZxCubWBpu05ZAkf//Hviq6p6l/SrmHVOzIudg8jQbUDyYojhNi7CgW5LWYK7J
RdPbD15fWtABd1gedL8Hqrq/dTeJVDkl47Q5hXlfVGUU/L+Je+GG34A74fovMVjS
lDG5z3mGupk1+eky3Ximo6RY/bde09F962Nj8SvkYVrH0gAf7P72tybLn3bNLoYX
oLPNAYyL8I2DMt4wEahcEZHEUlOM7kea9BUb61IzEndlifcjuTCXSXlQhikT0YG7
Pub5DnqoDUKkkeRDcPObMkrKjIZSHn2bp/I+LD9csgzuFHHt0DnxCrZOvogxfxvH
pX1LaZF+8kiiUY4WRlaq0Q7oIq4B82/nV6ooQDy/Ueygc9PsnzAZlKQDyU+bQgjY
dOCKPJD7fTsnkbmWPSSeP0BYrV7aMQCJs+jYpnwiuIuJYXyU8kz8p5VJ5+gbodLa
dPgdD/o83hQn54SOYRFmd98+ybt2ffDRwp3N1p3KzyS838QK3F//oowdkF7aNNt5
Ltk+cAL2i/SMoSRfyVbOHUroBg5Qf6wzA4cBt9kbsyvUDqrh0YczWINS3+fnWVxq
IF8C6tZoJO4KeZRjB7VixRmux4svkBtCF+tR+LuDlQrzu0ZgNDP/ogFJTrAMGjrN
q+NkcM/dx4bT5Mb5w+gZ9ccL0ejgqWf2tyLXiw3QyMO3GNljdwIPQWYjfvWno9FO
vQa2ek3kNcAWIC/xqLt7jRbKAZpEBVU+qVwxeeHDrRV0ffY+JB9X9ib+KrJ6HcwA
83FDv04qAzZ1X+/NWsrvpFqMjJPi1O0ppROTK6gGETuNPlRF8VgjtEddbpkoNbAW
hOhzZq+mlQY6sNcMq/W44ml9TjeWTTDO1LfnObT4JC5B8qJsukwG7L9R7P0TSr5V
dNyH2Hbxe7M1LWIiHvWa98KiEPFXVThZ+nBRkn+RLOf4fEfQpqNuso6oDFnC7w8l
GAzLCRhn4CBPzG8i/YHejLHk5tsQ0LN7490izk2B6mFPQReyt2Zepq9iiD7btZSy
t6XfXb9iusRRNlkesI/fd/9tXWBRAihfpJkJ7b8uATf21JExw9jrZqSvN8QlLalI
eC3B6RhZ+Ccnk37JRIuZ/zyEJjoSMqv0Xm5M79C6MJWMvKJ/mEXWEZnfyCa8IpWp
tXxWcXPVT2L1ESm+TkBQXTfMsZ687qvHS4zdWvLaWOS3iuWnf9U+Jn0EJMfdRpj2
U07OMdUgSFh/dstFjBraXAOvPy/xSfWZdW/UcRsQVyP2uhJ34BnE3BLmOAN6W8hb
tEKykFZV6Ah9UFCHYPMjfo7h6KGiDQk1U6Y3hy+IUa60ivkpkFdjP3AFgkY6fWWc
WLFBwpZdmrY2aEkjmWvNWGCnSedsT/Ywq6QY7bGs6zkvI1MVkyy3B2RkfwfNaUca
wXGgYUWxIVNQL9bfg8aMg+8sg3HUBlJQU1v38UR7nVJYH3rgSWV9Lx+mppOl7T8p
AaOHAk05kAhgoa4IcLmGO4y5wihKsplDhI9CUL0XZ8nJrFOtHA6UFMNWTopeckpx
UMeXK8kJBJVKgvTw3KcbBK1woIowj8vkYbK0X5OrQ2oKWV4C+BsGsOvjEyG2qnio
7E1aWsZObYO7loLV6THf4V7wb55k8/kmn2N69Q+eCSdvDwCWxiTh3KGveTychGp3
RFTtc5J7Zd8xS3a7X/ctnWXKbXG6ZtJeaHkMujOllvpTUe3rAXkOftmYpW2UUkMV
p2cRDb8g+AkgKaDtZCwLikxoDrkBQQ7AZ8O/VG9fiH7OBDsgvb4ke+QfavorZINA
IWYW3w0Vedkn4orIX4OHHgMkoH9Jeq4aV36C69CPcAVnkbwpsX6XXpFboYC9f6JN
lmbYYT+azG8TIPO/u4mxi/NPaDmd7F9riLV2K55Pqrkp+Xv3lqt8P9Ut4DkmQtKx
JVMjiwxOabyFs6eVMG6+ngO1T5kwoPwXq4BIRyQMYy7HjK2tIAK8SbnuBOtMc6TQ
ZEFt8fP/lmIN8+NIVqALhTJS8Op88EkFr8wklgkqJaa+MlB07l1r2EmQybvJvB5p
HQdyBPo/0P50X/pV2hAny5RKSVLkxxaxILg4k1vddaDZT8RGIacLbEsI5HFGInBL
66jFT0Vx2u80rWBqikvHhFD+w4l1MHYbVTLTgdUekDAYbiuPx5PN4AtwCxmcET5F
y/Q98PbfdqqG7rZ0y6m/n0fJqoNomR4vwYtlGeGVexpgKACWzL+sXrHeOT4TiNPX
Ylzln14Ehl4xi9JZLB0YoTpvfNdJq0K9MRnJcE+2yEhXniQHaf67hW8y++w8m7Qa
0ln2HVeeGI9XwgS/jWnQd/T0IN5MNDSkzETdhPr0PmWBGjYl+M6HLroDsD/9E385
+qun036OW0L3fTbH5kK8qws0TQmEfmZgCGw2QL9cc/rmjlbsFMJcmcuPxvn6PqRR
UWbFyunV2RW6UB2EjcU4+lEvzE1ewrVXs6GjixwAoaeQxOfPBS2ovUwsad5g38/O
ZbvUYvGgLDNQdCmGLXY/5Xkn5GCCNBtp8GInzkiYlPWjb7fW9uHZbMNh0IL7JKBP
ctZHCspu2nmwCEIbBpkQl+NszWyjimTlBgQL9XYv75Nk6BDiZBUScYbNcMlq4l0W
jHbTccs339Uu5SEgGrcZUutDF79fE77+ESAkcP/k3Jote5CoY6ccXer+7fLUxXbD
0EL7dLTbHsVWhltPUHWrwUuCj4ZAAF3AaNY6qXEaaGDnmvZIPSW+InFlRZOY7pSM
SN2cwdE4gCDuoCE1SD3HMUR7iOqbbGldmz0KeC5Nd50v8Gr6Kx7To6T/GCHimu0C
fL9J3BbydDMBIkub+ff92LDa+JZmau1G3B5sXgKV4We+twhtxrIpHd7iEPeUdaQl
x44c6Au43laY91bDF2SeFvAD0bs4261aa3+20A+mRqWnTmR8YusaLziWmhj8wKB3
EL2LIXUFG5t+O59vH/yXyDMgdy3ub7e2MMgbPXEBqG9zZiW3e6KNEPIr9sMgtAX2
wql++WrEcaRAaw2AMShfbyX/qgE/ahGEqB8eiUrTlb7ZnV2sfxmbzyygbDgEjjJz
5FigrYujdIdfWasxU1uQN4/RKg3Wrenz7Gz12f0KnozREinUVUGSoKFTwAWG4kAu
zOgoth6BRh4Xy7HxRmIpDIMP5rNc4s/a2OTs2sEVo1qXyTswnGqDd8+8GFAaQNZj
r/8sNyh0wxMHk60o+dVstSqqcAVGm11G5STgPncLZh8V1sn2Xw6AeBjzUgcnPhuN
cyjW6iDj9w0h175et63lQ79ldVX2yAik1qD0drVNS4cH6ieE6HBRqeBc3d8QovXO
Tkwg8KVslcvkFIKaHpZB5zWzNrDPnlMr3HZzO1hnqcOM+WIEP+Nse4Mc/houH+/I
JqjY8PWkrXj/7i4Bm2ak/l2nf2mjcCmdhtdfLleXUyGiL0VUAHVw2L/rhBNjZvh0
TwoIopaytkL8ZwOpEd0gEmajaoESrKFjKB2qHxakMjG30QIZ4nvdS0DV/thhXr2T
fLqcWjHBASwpzxmdsQkFy/3MGYI0LK1eeF8tizh/zO6txSsaejYbuku325y/usaV
WwznPhKqzEBVET396Ujagfgj5o+vUFTx0hODdadtEyD7ptk/Br6mHutPPxMImp2p
Pui3CWTAHZVfv25ZNP+t/RgOrtLTRPb2zj1Ql8kQPv6uosa8opKtllCWz5j2jERV
0535oM//5pT1Kz+1KKEzjzmVc4b7mqkCsM8gfFrOR94Ku1YNJoMJfXPvIJ476FAN
Dgv4wMY6YuIAVRZyWRRjJOHiQCV1+/ysVmrwxCYATag87TMEfJwkYVNRS2OcVSdA
aDcgvnvl6WQtbKGzpP8thcAxkrvDvILPG2FtpoHmHs1xhpk+qAdStoJa+/eorEp7
RcPHn2NPi80n7SfNjjQDcywJNi9RZe+NSjoSziPZz2G1Wf8XxecNdq36OTOK1UrQ
I7cHbxqyEUyNeB6slRlCsDCuPf1zttv67hd3XxHz9kY/D1fX/7mYQa4Ha5DzdnDT
M6utlFYnJXVT5LAjF05w8M0Zkix2/bneRUJrO30aofclxOcKR/eCAUftnOzQJ1+R
enSWqy7fHDZs0IQO1hJf1K6QwljEWpNK/J5OVPpALYoA60hE2Kh/sbMwIwhLo0sl
o00BB7pytaqIgKXRLvkJhH4lWzICncHG4LilISaboSTH0aIeUp4lAc0ujOj/2/Gk
DQdETbSN2A8TNXWKypb3WrntaupL0YPQShAz0hi4SK/YX/jioI6KxbO6jl2Vb0mG
ADWQXBuI7d6stOATAqf3euJMr+OrBFod9vhzOOgfnnKHAa6DpPwqttvmg/nefMUr
htv9miUSR8ez9IjbqSb8TDTUn+Tokpp65CfoSrRFFWq+jiN6bEtyO52MX6OIJ6P1
GuiMXlonK+Lb1IHyQdz57159cUDmvFqRuq+jilKSp5iRFagfDZuW8uTMj2x902lV
4syvSQMmzH3cXCCXuIM6ilSzbVrZPfZuKuRi9P3iocWoyPWFDS99hietHXhS93nt
X+EdusiXEp7VXT8G1Mr8tNfGcNvmi/qNyfYi97YwdidRubs3lcmAD6h3VIbm7I1+
J/3GrNhnLDbCw0aq1i3f/e2gUJrw3ef31Spng8PjKqF4gju9aAJLGfW/qWXowPBR
b5mbCvyqERVHTJ92eCc97HHM+BGruc2e9MlMY56MYCbpkfdpbjGU2ByrxJPbHGq4
rfkwPlfidSpiQZQb6SWhRC14+kAKwEh9RysEHZ18EOr8NhhBuLy1WI7pIzMrD6Px
hy+PdAfP9u8QvH+gGIKT0/n8fvpE+1JncagRogDNjMj6mot78uJojlUbdsUxqlo2
SXTQ0RjPI+F4aGnS+1yIHWm4Dj2Vr63IPWmwQA8mb4KXBSH5QnfUGFIFKoRdLTyL
ZUP0hP7hJ73tHmpkn6NkEC4kcqSD9tuQSRlYvCFN8WxCx8jwuj2Y2QUdeG1sZeHj
P3QHf0r0soz+o/1bPvzIdNQ7eCPe6WMcuVIkJV0zbxps684TXdViGpSlUjAYjZ9a
wEH7SmCJWwVhnTt+p03lNQm6YDryqxhcqYfO5rAB7VZK7FPrKQi2v9mjhfk5Q4DQ
GPoUP0/tmeBiQ3rXTqh6JclbTwmCl8wMchwwmvWVe4M2fJTtowx43xSiJwvVGaxi
V5A6ZQYS2mXs+t4mN3NFPspHyArHHp6rVnkN/D4WforuSWLq8Kof48e94JPKpcpy
g6G3hVwOQnL3gdNSFlKlYx9IDb/80A1dSdK6nm95LwqGJcjzZV3Z+8Jgh76urvaI
w/KHeVvDzwfqJrUU0xnCWiNaiQPlcAvxr7oyL5/m+oOSmJUDNK4CS1gsiF+lvr9M
GMyIQOQ2CwUzHkY4Spar2HNIO35Yn1U+HTvRcB9PVOwChqMgIwRKUjoI+dVCW6oy
7JvlaAfdNJrUV75kxM0sXtloBK3JbdQIXGHDmZhEMUI9Q3WrouVEvOcIu79nAlb3
o2bw3lTKYzLi8ILzRDUNOaKPO7pHcmU0xtrVxZU55kSrIUFVuQs4F1iUiXX4HTng
LgfwMzpPBlqeCqehXydzNhGV0L2ZHBh5jidsMxEt9YemJURKLpruAbUNOL5ORKiO
j9Oo+9DyfWyA324acWc7danNL5uQiV1RpW6bykWZZ/5l0nMxsOhHXDOS9RfPWerR
G/mzSplHN2n4KU9FoJUnrhbJo10r7qsjBltLC+I7Gki6WyCrmGgdrNyyyTysggz0
MIFdrzyBMbrhn3llzdjL+3SBEw2OCIdN+jUe3xYtd3keA7RIQkGfnuRa0YHSxcen
o7QjmLiMbVmwpuqXFElUCGXA2C+7VdMDwk50V3MnHzJnqlfXJvCMKBO1mntyB0ar
NG6kD3w/LmcJcGe/blE3yaRYoWHKoE/i9cLQaJwJo43ylnQF3vCRuDCC2OvxcZcp
njNGTk9u98F/dKWYclONLWnXcSSwi39Jr0m+FAp/qw7v+tNr69H26J1LxCMv/fHe
9DPVzbaASQwUX5NBZ9noc3JefIlygd3cFcpchLR3HcDivIoDY1jaMFfiuV4Ifh57
l+NIn/66H/NIbLkzzG7+In+VjetaFgxqQWvOEBQ8Dqxv8hV/v6Bl2ZQZuixeRrFr
Ra2G+BiJtez84HAsvVTRHCtks6T6iK346AmSxeNvXDR547yoA4ZtZ7cYo8VLrc9J
fC0PuRGfX6mB7wWCxAk32ru5Xqy0lYEVMIC7y2jhtaWaHipAToYuHZWQbzOy0rnt
eFs851pvedeHpjqa8Fqm95u10Rv+G9hN35EydbBlu5tI0RBCz1T4SY8N4gygwg57
ZbC+KRnXd5ckxHqWUIqJgOv1jrZuTqnTjDS0lrIEr0WH8hBVhjkQzgJaym4vikY8
/qwsBmvRgC2Ounx0biAFnYqHrgnLCCT6du7Z7rSnAEZmfmOPqIMLyo87f3Paqq0Q
bzI01ON50VtO5rOPDzN680Y29Jar1+9AMRXgt+wJXoErXpX8ojtzcyU1gbEwLpg+
QsgPAsQmaTU1GIqwGEUo0OQa+a2kbrX8rIwjYEVHTqg8IigbV7qDedZEeG7xuaEP
BCPDfP7UDxPvYiFbguvl2hsjXF92GinCb0B9HnRbL4ll1OGnjKWxYAF87iGDsQmX
/imAGC9TpHnMYabsJk1SIjm+BMvB5aCEQWBFB894g9LYR0uIs2ZN0oOUU93H/Css
VeX1q0PRuwdSHt5A06uLQSv37T1R1oKooHSIykrdIX2Gk9LUsInSZKmmvr8JbYZK
MWFwi/JMlol9JQ+h1qZZvUBpZ3YbeZqqpomDAnVca3mbpEJeUXXhE30GAQD5v2/u
IfZeef7s+vyiQFG3wcyajEKGqXBCtrxLNyABiaCOQKhv76JkOqwfs1EAL8YHN5C7
6NWdf7Ekme0fjKRBT8Z6pooMlVn4zsfBcd8LXIrH4erSm8hBdEQdTT2G8K0ZSkTf
FiaezKvzvDML3vRQMmXf65jAwkXw0rqCcfwC4BbXShrb/FwnQJo6LYtKw5+9S3/c
Sr8TChBUSkthJMdhBXIInheDOhYZjYHFoEnqbuIjmrjvqXXQpOkM4aRPaHZ4SHxR
UZWUhH8kxIOYfT5WrhXfQw9hj1EIjcCJIe/3zgFr2xexyvD6k6nPfi/FZpWNm/+H
DJfmj7JzemtynN/EkYZRGcfJn+jmOCOw3cMxSI/uJCdaJ4+irAsvJ8QE+cuZjX4E
8gXmMqoPpM5iBI621v9ZR4/ScLgDJxMitv+b8q1EDJ0u1be0YdRqo/hc3ToFt2pm
Lqq5Jkve/QRlOVkh8kCbXJrAuA3+/GJxDMThaD4hGrGaF/Hu4tgMQV8jU16teCWn
Y+yQSt7JsNKcAYxdiAkohMdejB7Lh38w2r99sheToYgfK8UYDDTPrUY4cR1V7TqM
dcL8csilLsSK3E0DhbpUfuuOjP8we+8Nnub1JEFvFvPZUJM8gWmte+at0CgRZDy7
nKAVQ2pRrj+8AEDrmH/UDw==
`protect END_PROTECTED
