`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nzkKtV8K1ilaw1GK4r4+x3uPJhMePg/XYU3K4fyg1wb3lIjwdYwcEk6g0A0RStFT
IRl+iBvWJqerYLZKSOOfmFdXFxy8GHdUYt0vGSLzjKFWy8Cf8hJsLofiS2uC9Z0R
KtHy0EObO93sbcpevz1Nr/qy1Jys8vPkYwvzwSbvw4sKrwmSaTQFamULTD9jaLNq
CphFCuQCGq+yIFsvk8dfJe4IrraIqImVywjPhddBas7GX1vOpdLCWAyQGzxwf8lT
`protect END_PROTECTED
