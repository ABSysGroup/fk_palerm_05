`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/NRViwd6B/BVmt6H6BA5CrXf5T5cCa6OGejAZK7PhbfRy5b5GKu5fVbJVjyqqofG
ccoVcI2Ifc8eN6llAyPTYD78ST6DdR2mTMdp6tJMwhMTqrMXPSx4ZKWAatPCjdLV
eqI9JfglO+7xBYfTEmRhNELWNEkkAEKBHO8rgZooMpsbFTtY8gGlYYIwDnIxfRUa
JB8zqZjsj3YYwZ+6pCFNj8Uarf3t1F8RXuk/LQaXW87kURzzKLUeWbUuXbY/oVCW
lTdax/ruzK2btK2/r0Hk4KLyC+afEw6Ja6MR+0hT0g6wCBB7ZaDKEn3L/xHdHGGH
MHyv3NEuDP1d9KNnGvqgQq1WlYwbKeDKZH7bADGVXudh6aTO1PWPezUDbHLcwx+d
Ko3KKnTh67NJIay5K7Lu3zkizgW1HiNvCv4+OfmIbMUcbm6m9G4QGcUjWTc2Lgo2
5YRjCdRANxnNdf3hPndJ+0Si1pC5zhuFZJWZz0dnHD3hsh2lkRvV05GXnLE8Dp+7
6QMBv5GvKQ7K8AbfoF/4gesAwtJB2n7p+sY2F0d0TJi854haRjwGuuSTGe6sPoBA
q7nEShKexO1+KCe/JU2uRXEuZp6DLFgXrfFx9s55a62s6i50uT1Jk2pHztgJrIri
/ovt5cmdwWHSZPhSaljKEH5z/WZcp8zpkipGk5vMbESfTS83urz6xtUowGWB6IBK
M5vRYSA8i5aFXwsQfAiuziKDKrA67PsNV4t8iHr1HA8IZV7Fn3WmBWFerdHyWu+s
iFWv5uONAimGZL1R5qmYXQ==
`protect END_PROTECTED
