`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GHoZawuh8FrLk4qcfgztMNI7a8GWJBe9oEC1wzsEbZhqDqYtjIAG6tF8wZpR3pse
ydjRbybViddEric1cCF2vBLPfS8iTf6PB2OU0mAQvmKP2dLKtwlljJ248nM31ZXY
7pbNnu/BVNlRaGDKaSJBmt3rFSSAl5+Hphp1ozhSSMtMYZn4wrBPYffNlO0uNX1S
8L3Pw/crOdseSBlYd9OSa60tvlyguNa1jR1kJIvvXiP84NCIkRYjYbMke2WRiFYW
wpJALTO8jfzXYs2Wyo8N0KYlb6Zv8wUQxJa1pfrLKMKh7T2c00xVqGZy2RhuKYvC
nT0VBzsV6zqJMbqnNWGLyGtqIPzVAd9hjkvZGH+BMzoMKMLqksWk8s33mtmNJpUw
jmRVcKKxzoBCXk+LKPblGVgm+lf3WmQYk9mW6TvtYtdep7v3/AozWDBL1d5dfxpG
XwcorOTWE3KKlwsL+v17nXvL0/PtamRZCHGDayRtcyU=
`protect END_PROTECTED
