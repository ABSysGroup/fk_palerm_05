`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hCPPjAcBi2jRgHUlGxBhhCyD+wmlbLyFgOu8lSRFGHmnhfAYPw/TDiulKtE8Wgwz
g+pSRpIqzK8giNKxZOMS5I6HrqRc78RmA+8CFLkD1sTTLuTTMltjPtsCwSpUAZeG
2CJaTGOjk4SKoWMlGSaN4JXnme6WBFbAFIomOdaAA9QCQ6eH10Rvm1dpeIZ1PD/0
l0vTrc8xyT/BXlfLEUcpM5QQ328pIL/O+CyU477DwVToWYCaL8QxJb8bV6Wum5cD
5JbO+9HepO/WCmtYMS5Lrgcf3yBeIbSVwKQ1R8NmKUDOakiBTp9YUlobm0dbzQra
wiSVBrjhM6I4zuN/drTZkQMZTtbG3DsZVDYIwGeM6TZeKKIMYrGO723k/yACY41c
3FjTI6HfWtUk5aOhSnw6ODkhyKwp3cCKXdKmPsK+lURD/qfnJIEUm5JVOWmU+4FY
PkDlGWeyFX3FOqW+BFrFww==
`protect END_PROTECTED
