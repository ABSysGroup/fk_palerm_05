`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vfEGtzgwTNKEinvoxL2NH5UTFTVs8Lx8hJRHctIemRJEslxjMJC57qcnra4EyE+u
pn9V06dAWG5gg9CUVWjLBFGgpZVEKXdTlSGXpq73r5njypw/6kvouD7JkqOMZk4Z
p93k/CGqA5p0P3WWhndsCu1TqtC06P9kPv+85VdaLkewg2rS8KZRGiNfMtP5Q2c2
TBwMOOtsJgeVCvVo5apPrwp9sjhuT4nvpUPqOyv9IUwFcBmhRBqEEkQXmgOObfqO
Ak6cpriNphPOTmxKlBVpijK+ZfuDU2aBzr3tYoBCo490f2opazrJ6i72X+pBHghk
FQtSUEdFFuDiqTEz5OIe72ZIjUBbn0FnqA3tPyMaYfaDvL/L8Lemqk/V8YKVBRoz
60N6IM/XX6vm+q/NWuZxBWNZhNuCuBQB819yancHQukQEXH9xtGzneVD6leZ9CKQ
`protect END_PROTECTED
