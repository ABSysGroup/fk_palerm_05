`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2S4ZbytIc7mlhqDNqw9QmVAU2uLNPrblPHyXYxnRCPVeH4VfWj+qkIipPXq/JAeR
9G6ug3mm8LBDmkXH9QY5KuM0/+LEjR7HU71W33GYTQQhHv48bVAZZ5fuWN9Jw37a
oHa8UDoxIa25fAa6oCkDJDjaThD7meEig+KYAhWJxVw5n9LaNLXU35F+xnTLRKs3
IjQP/tMmwnMVQ6QNlyiPIkPzY6SjFdUG92tLVxhJOQgYeUo/+WAWqSwkhzfAZXMJ
RwyI46h8bjDGjqhOyCHKCA==
`protect END_PROTECTED
