`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hLhEH1h+F0KtjtGxGs6sLVpZpziDNzavOwElIp/WaY5sAatKl91ss5pydwop66XG
0RPYBpbwR8LEbnwUMmED81BK/S8wZkO+QKcXE+xBurHcvJyfQewbP1S+TjLG0s5V
dy5cn+yy/wJuRB/xhnSvAqCGyUrY5yk5VpURPuPNLPh1CEY1kIq5R/LVlLwztDSz
FJEKkoH36pFVOl0zRdH36vCoi4qjUc08oGgpHvKh+DY60Lz6Ko2xdMhvSURhBC1H
z58r/1d69JqZxnwB1s4qtdMATcgH8HTF4TPHJ1VWe3hccr0180N/Ln6hlsD5RZzz
zT2S04dZZyU/f7rCbTHN5bvba+phVU8E/NmzwfRwZ8O6eKsjCclgAXM3QwPdBndV
mTZAgAUrwcfI5+aU6z/2UvZzepV9yguq1/ijmlEOWbEivgZz7XChkfuc+Ev2gBOO
`protect END_PROTECTED
