`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ccjqwlJDp4KpbWhzuyoBzU/rJ27Abcr9VZGt3IgKQYOriIG+vhbYJjv2hI8Fce8K
AUL6SFmgFf/ImOoiug18OBKtlfMCskAyg/k4o20y2ll0aysRGQvbZykyJtVBcGrN
q76wqMlbaH4uR83MaoR+W/PaEzK5MayvxOIH71QOlO5vwKWG3KIm/VOzBa4U0oKM
O7eNtVj7sYNr+DJUY0AocAskfwKdyKBHuQL+tXsdh+4iljZkeolWDce0Mh3MsLUI
MFBc2wlKTN2j2lBF+jD49q2WU3Fgf0oZ+8677s4Cae5apmzBrZFoP2baa0XVZTsz
ex/N2i6g7GcEI/KeRDCxHZJQhqI5NC2+YQABh1CQ2UujOHNc+vVFSWLXSYTJcbHn
NNDAqQDFoMf72CfCMhrrZ3sTFOFgSWF5+DS90qNvJy9T9zUIvVZLxwGViUtDZxO6
4/JrwDotHL3Pyw47h40jQbP+LQ33V9aleUnMAwvL4dDRhoOS4UMFulPbiFXJeyyj
Fh0Lbz3aKsI0tNssTiWmgIm7nplWTIbt6pdMhz90sJXOb3vp2FhGVAZSI48BLuJk
ToBnUQmxdPxqoDbUYJYpPYL8T0DyJVRdhy8Pfa2XxXUha4aaMYUoOx9x2WUJFLp6
SLw+nueJjLcJSNs1qvzsBKsG3Stjcv+9/RMSOsl4sk/D/Ckw3o12iySvGIVGvsAa
gwIrzzI+vfNNWw4MfCVebSRowvbHeCgqVJkt6i5pddyHtf+PFpRvkO+weSvE7v12
6+gUL7hhvQUuLSSd/nvpRw==
`protect END_PROTECTED
