`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GS1yXjpYOZYeO6GvbhQMXPcoGVmSA5ch8mFmM9Crw/bFIlYJ3bm6h8hk48ul7TBq
+JiKPhDDSZrikxQgdN7KGgF2pq974krlsKF4X6ELBmxuAvGoRKmm/7U0p53SMLjo
NGUzHZF4nHuqCrOSn1YSmKGEeKG5RvwqzcU0rqIFDM5H2I8vqDSUaHL/THo+esYk
lsHDYiirpX788Vp9r5uumLDvtLpDTY5CDxWIqFyrvjeGe3oeAAT4sGgm/DOg8F/K
`protect END_PROTECTED
