`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MyW0XDv33QVtvUIFzVjbRL0NWGddrMcGIWEIcU2rHNpjXwPsKOHZuro87BLkIbR7
UhBs/K4jaQ/B4Ko5onbTsgvXlokEl7QWh8pKKDH1vl6NjI6NaZUbshoUgHSRnv5h
v4Hf1zurUp4qJusp4+lLlCbqE1rjIQT1752LmHTke6O1sjqxBvHyXVkECkI1oong
xqKIrJvxVISey++PU3Oo5Ys8L/iHN+1+nEOHfMys+Px4kaMkOS0hNzCEwWFWHqJf
MPDpdyxun1ZllNosYEd3HmLw0n/dv9F2MqyMAYNVb7CcbZ5aJ8TUHnKRB1+fA/ce
jB8J/pj775/OqgNpwo+Jebkec6lrf/GoqDEAyhsCgQTHac8me7aRCA3HFs5v2PJ/
tvabBofJnp6qwq5cW83Aux6cRZDcNEYTVGAozBrUM5+0OqQY6DPZdHH57IcgXGqb
iz/k43Nqg5lsBt7yvMsgifitBF+lPdrXNSmp23QarzVlri01457VaPtLeuuG4VA1
Iz/8td/FsOoykMPbBFL+HBezeHNLPRQDX0AH9Wavso4nvTObVaYOnlwzKpBYjQzA
JEExwxtO0GL0p6luTnSPoiszcukrWspoz/7zO/tvLSy+PpnVArgMRTnPV5vA2AAZ
tBVmSgD4/AhxkBmsGAe4rsQverplvDRn877blhOnsAMlA0ahF3KC6ryd8tEflsEm
VCpxcok+7FuQ3JIUsVAnoAjZjAO+TKvNivtwK/oPgw4=
`protect END_PROTECTED
