`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CmeOdwIp1rF1rK3/9V2XD3QgCzEY1H7zTFjtQ/CivQ7HXpvRiBe7eu1qWrh0y9G2
8Yd/oga2Cbpijg9Ez9MjxO2l3vqD9Md9WiXGFR1aVDb8uaJ82VwHBwP5zsuWbKV9
tbUWH243nQCnvpf1UlWMS64YVWQWZPlkQ2IONB01czvkY8ID+GL2dS04ChZ6xQiF
o1TyJk5R+FdJ/5YR91Y6mBY+8u/EM1LprrNEDAngGdeWRHjre9bpienxaYiu6TqR
dsRGk/wYVVz35IW7gezpA3EzI65/BN1/YA849zyoctPIB2YX+OBE6Schhsn+LkCV
6CCYlhjkJ/s7DdiRu7DvsSOOAqC8yaqSpcdJlUhqmT+fFex0hjo+DHb0p8E6iiXx
xyxuRh6MYkGxTiMzFijsaiw+wW6kDBqSdig8TIrnj7dfru4Dm+4rFQqcPhVEFBz+
lOLuozzFLnnkUmgP1TRIC9nLL+2Nmd13JG8/fmcs13Tw0jD5iyBZvzm5cmJGEZTS
P9RkvnZF4BcbsSroMmm0SegOGSLvIE5z7AMMq1FBjvs=
`protect END_PROTECTED
