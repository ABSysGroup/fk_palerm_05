`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PD40bbbnuJe8tl9JJWmZhglPoyFleAKt1UHvVs6mea0F6vIaFTXZmb6hkkHy+eam
pt3ZISFOLX/4H69DNr3sTZel5lQFZT7L1miu8xfCQCChm/y+UGeYxeTBPwSv/bfV
AGQQEZ5+MRI9s3Ps7hDYfcD7aKjfQU6O78NDdI6/mhr4BeUjjnNmywMcIoqE8FEj
FoLlR2aGCHbGII/Q0AONffgdxEzBttJUhQJMUxDVoeXlyyfZpws9IM+hdIpmRcat
5SN7deC1fWZnGtbnfb3PGUgEaq45w6QBBVn744R3atxeigPQd6vkkS4///N+zenn
fqY86vlhG3KM4uZs0pfHjHvskq3qLlt6eMyBqkxq/i19SolTsPrwIEJqZfgYBC7S
pUbxh/4yqxa6o2Kb5ozVFVmg/R4dy6zxjEB9ZWCLs82I9zWAp5FRHF57D8+OO9kF
C1Jw9AGc0eGK2O56Ti1LNAsGz5Ehn+s0ierJavOhlWBy8JQt5Ih0Yy+oQisnR5B6
DzhZJl+ipMbXwMtLAqf32GGW9xSEwOUFAKq2JnQ+fHo=
`protect END_PROTECTED
