`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lay3QkKsKbJVmSai2HHwU9JE8dq3Hri0noCI4id3XsIgw+bu/AHFf5uN4CnG1Ea0
OuILCnhXMj0qrImJpIwQxpKSIBbhKFntyLeHQmijqbLct0goDpc6myXEDo2PHp0S
mZdM6lseLPm5AnPYNxPgIyR3dvOJp/KMK3dTHzBiOdj0xzI0pNg2lsoxTznSOiXE
/ctIl5xkA/CMrf1LVxTlkvNoCWy4URt8AwmCvfrtdwfbqEani6Dv2piS97EDDr00
5D0HxV1auNszfMsxosAQn2dp7HgytfgDGvTHbKgm3oW422TOokmocRLNRo41gHkw
O/EU29xNG7NK3u2joOIAmwjjIf5qNM1tx+l9xhQ6TqX9PEv09Rln29xvd0dsFq9p
c8/L1zjR2w3Sk6nIjDyNPN85mNyZGNK4QfyT1Rx8XtGGBnKymy1rjYUIgn7DNQNp
7XhEV1hJ4Ux2g+Qxo5Z4LxI+Jnk+9VoK8OP9ltncfAsq4PsqLypjsAduqeUv9etC
bqX4I+qQ4d/kxtgCyLggU3VKgiCCKWLD4Sg7kDHgdn+jI2/sv3T3d2/MWgeU6M1j
RMDCLFkMHVduj4xHKOLsKPyozYF2cOQAt5JpMo2AJujbguXpYMf/IErrZUuPPzom
e4cvPhEOtW6/a7WrbXZmt61nLSn0qT4qSg04Qh8fxh10Co6p+WE3phFXIsvNzQzq
EIq0mOneJs/9kR3ezW4OtGmIuBM3oIVnL2yXkO4tWKBpUMOyD7iGXd6uxmtatKc+
hLC3A+JGH4S9fC9G0Y8tAFoPA9R0CrzejWipmZBYPK9sCKxu9meRV3XFlXjQddUx
hQ/VeSa4S51Ffkaz+CnNaaasBEvm+olqnA4xCTjvcFNexQxuFM2wYw8AH5gkKdgQ
HYuFz9VWLKNfHsUnrP7ivrsl8UakYPfTQUXHi4YmwC1sH+gfEjnu61v7jZhybe2y
RcsFIe8lc59zonMl83U7zZbps8LckmHdR19oFdsudSzr6My0mtluAWIRgCaCcVSF
VIGTqm2NG4fSPCV6gc10R6UALD3FlBuvE6v08Ikj1WWzipZUUlYo9ABPpqiIHCMY
oxw1y+DuFBCRcM3lzem/6KJevOKowrkwKceAPZyIeD4AKz3YjfPr1m0SMsigMyvA
mFuNQE6dH99euS6PuEHHOK7SzD6n/3ZKHBUXXhlGOghj7Xyt8DrlDYaRhlnKNNh9
Z6Meo7OApVoR/+Xz2IXbX+Bm2olnq4h6mHT8hDgqzwwPZagEexv79lImd5LCUV8b
FoBa33gya5wnn/oEys7uGdSpfhqRKP+ZRc4Q3dSOGudYb04FdDFs6gELRC65DZPe
t1+ldlaP2YB+6ydzF+ddrBLoOBcg8eUMeXbKB6U19OOOqTm52X9dzdJq0GI9zblc
lurh+mXM2d//Lm7q5Odroam3XJk8UHm085rOJDlEfYuavQ/VeTOopfebw19j4jG3
gxQe5ykthofZPj0mnDd1v36EjcWt8q+yFCPRtj/f8y4+1KEKrFQBkZMYD26hWJFJ
vhS5UOcHrXN4FafE586biLDUauMS/vM4KwWC+b4A9A34r97AeH/I+ROEv6d8jdme
5Q3nz3GWZOFWzsDO1Zr9JoTl4sPSY3eEZ4sOmH3xd7sYP4qKu+BaY2HklLOdMSAH
QHPbZCgOz3XAqumO/sAORujlaEemHque2B1mBIwl+lkubjy4lV2NmnH/oDx2l/DN
YATcx4s+smbUtJs5i0wxYX0Uw3JK3yksGXfqE/cS2391U2rTRehOhmUHFO7JnJZB
Wiox9eed92/sd5nGzYbduiqDzijnfDeaKa8ObbA5zeABklM/tFH3Rr4N+6O9LZii
N8qk1ManzEypKAmWqs+VBNHgDG3pG5Io1oBR9t3Wabwat8FmWpRkti5LX0Bk4MWs
PljoQ26L8VkCDfdJ9L5CeeOR4yG4WCgwoy1YwAJwJTIeXFeSV4tptXKG12WVn9hb
KFXBr1lpclnupVRlhLpCnTde0QprMnBmhifkR3G+Zivli2myTkWYkbyZtTPLiT4V
6bv7l6HsoHrxUh8sRWZWr0Otls7i3NvcZtdzBL8FLdQg+fE1PRVjulRT4MrE2QCl
6cOSBZ1Gc7Xa/CttGIfVYkgt3rLGPXboJJgwbQ9YaQtiLp+LKRS4hRwSpQ4elKm5
Uh1p38nHVGmIYXyz1t9iuTlTLMjY9C3d8Rh/wFCDASz61CdGVNJWnOb4MXq/uktv
ObLFxaNm0K4Cp23Xrg/ki2JCDImfsCuu0hr+eZI7lnRyZf6NTZz7qdXGlLSHOHsq
wKHdktEpC3i0nRuj8A01JYZ0IFSjSNaki1ig/DtnC6otIryOzGN39ijFDtZtFinU
2GsL87mksNpDSbYkijisBFH5671xcTf8UhjdkzRI4BURaS1FZ8eKScKoLgcMTfr9
LdHNHHyXynRmPgOcngfs8RxEeUmET5vPmGoy3Nkwx9q4gc2RGNjs6sLt53VTYrHm
7p6TH3hoYhul1/GKR8gzYzeZpiRuSj15S+r5YjKF0ufqWm2GL61O8v7hssmT7gCX
7DOXbA7OPb7HXxKh1S97JDmU0FiwSOdSypthRZpKYmnkzk8c6hpM0oJ/T4Irm8hS
+fF4P/A2dcDQ58wfac/Y42iJX9G0c08Ay2aBRWBzSr+/Tt53nxGXqNZHi41RiB6z
tMkgZa5byW+7Lfb5v5na/8QDRG/Cnga+YkvRsNWzgVrjKTd0OdQdLBJ/dO0xVMr8
bSn2PT7n54b6lAOKgMZwE6wg1GgIXqKX03y5Pm7QqMY5USv4KVVtX5CKX4uxP6d4
GhC+cT2MWUJxV2eIRf905eq1rgkGtG8asRxJXxxipp7BL1ySlCm5d5ZnWUItVz/a
udKGNLP1M4nmyfBL8XSMtjAHn2tvGXMR621CErIopvgWcFPciZz+lntzGiJDr0ax
9OgTfRL7mqPT921Sh3uBnPlStONW+UJGUzXi195iLOV4QhtJSfC2WDIP4ModXK4l
t2HnIHUSe2JUssFih/NezEQVGNyRg5wVxw1WzbXbM907Bx6lRmaqjrEul9EmrAZ7
gEma5OGhAXULQJRdNSk1o970sTefThM7Rbh6x+wWfKRKOrCJRrTrr8AYEVXbFCj0
TNFG11/Xi1lvvP6N+t3VlZG/BNUhYH8+rAeyixgEAVhYCr+PvkpYYtD3OJWW3XUl
r5W/IlHtSzrf43eOwGWgeJ7gc4FsIQZSG0Do6sjfG7wofVQfu7tOQ5RSDagaT4J2
dpERt6jZ27EyAWL6l0wWI9/Dv0Pm85cAWNClRxzO9L6nXjF0zLCO0cjAnJuTe6yM
x21FP8csKtoKk4QC0JEd/qBJPW0HeXqDJxhktO8iYHMBHpjyYGuV7VvI0cRSrR6W
Rvtekqduhxhv/hnT2RSLTgdHLbi8fJlMCA9r1LJEPPzh37CmneQRMJ8xss0Kqdcw
J52E/PCmHSOafwkbS4tIT6bHj3ARsxIS4pfSL8bhwtqEGjtFUeY0gpLPeZV1U2bK
8erFRLFyVj9mxYvMzEDjoFlgficop/zS3DhrfDTHvxhKWkeCViRZFhyjJV8mLIer
M3CZugiE/hhQdqpavw6JEIrrg0sfjwac1hfWBi58hXYtMhpwde/OGIFQmYHZWN1/
OC1zGN3/FPls1WOqhaZe1Japo1V80ZsiNKzfV8z8Hfh0+DymETYMT3YY+kYGBWY7
3k3vimLWJlNi5CanCZSOUpVOJm7EYOfZE6lMYy+AkYnviwM8pcRhmkl+e3keCpjj
heGV1bu4BYJQ9X3cfDiylSppapUmb6Od01o01ThdeQ/swMg8AREFdGs88Mf79r9x
mZKiEhhbptOcfy4bQkRna8X9ELUbHblZII1dLuOMupXua7Y4OTKTUmXSz/05idJp
FZgqZWRyPaNDCOFlTNVsso9hEFmd9h2ansKYokhQU90rp+ZwTkOlIepQOmS01JZy
z4BWkAgEVKJKRsxRaUKhoXBRpGaKg1ZP5Z9tfIZxRlPNX0z+uI6C88YSwI2/5+Vp
TQDBwAaCJRezOOH5Dsl81IKFQW6RWh/C3g9qUV+ea2sZk0/ZU8AuvlhHAjxF3dG7
mN9bolPLB/LGPuOkrG4Ho3grz9bdysc80+eW/N0evThDqG3+D6UouSr7OcR0cEQh
U3aitVyAuGrbyVFrCcS7d2WIShHRY88uFnWT9UdO31EViI+DCtxiGEKwX36HJ1Xx
nx/JXd6l967UH39X+ClOj7KleLlSxD0PhGjapQqT3DsfNM6JtH8cfzW4Cd/XEZmB
34VijZR3Bc8y/Mfy95ywnaB/bMufCVrTkqLSmyecVdep9meGb0msV3lCCyZAWFLA
Z1h7Y3L3lLm+WndZV1ymnLtgqt2Pnlm3QdOsBfftu++kgnxH7/785Uxh1lqmOp7Q
LDI4BMr3yIzJEoXFbOS5TOJQqohf+KdLzjk2vJgVxggg24X/CVIWEYrAusjqRob0
/Szp6BspM22Kx0maB0dulOw0XJES3bNdpE4Qu65HYtxkHcjjXkskwqB4VktPP6nP
ICyrLEzlmYgKh2Ar/78QSLdje6no7rv9MDyN1cubnLxE2JQS+lR6ALeZ6X5dJYbu
3sE86QCru9cjRoXCgJqZiUOfr9HeDFDWYiAmdK4oRoKHPPjj8gj4MmrGnd2JVoam
i7WhOluG10F+wKpwY2GNgRVajIWxfn2CG5oj7S52E238o6VTtpSO0fu44g6iVZ8k
q8EpztkXkjnRpFU2sF5Iq31HWuyskUHpcBe0GIEpEndk2Y4ATrJmK5w0TGaAA3oU
8md98jgQ8Di+JbE1HaBFR6L9gafx6ISDRmnQhzfdZcNY3bWHCAUmDCe00n+EsPEB
RmUTTu3GHUmWZf+IwnfxiqXSNFuP+g6gR5QsY6k5Dsh2kg1unFXQhdNvFG4wdnw5
dUYotoGpNfQESqmCuMWEBjSiIqbjc1BEcn1oZbYuOet21YPkMhLStvEf40y5Xm75
AbRW7DGK/tPEZbCFNTU7kvbKSgu/Np2oHJI2bNJBcq9jeUSgVLYWXDUE0bVvj3pp
ydesA7uTqOWzwXRiLjTMKaWcPTE+MRs9ni5N5SPKnvUTOkjbss14nrkRb94M6Ubb
QB63WOfYyEpb0RFZSEO91mKFDQpjOGQ6Ke5Suf9H7x6/VbyKvX4yt3j2af3yvPFn
2RknX4zeVy7nPkt+61G2z7txS2arSmBWrGFGgAuyF91yzpjXYYIVWRo7l/nNlt3P
o1deSJQV3pkAd/iKcvQ4aqJWJj0Htfiu0omMrUEJGn2g7NjNZEsh0HuXRcbJFVHE
qkt+FX0WZpa9/di+dWlxjGIDt1k4EM1pxLRjyMKIQnOod/2OSbUeYLZuMzO5dum4
YFeEnECSffQMPCM2gjQgyiAUw9t4GFjwKsbi2Uov3BynbMgkiJHFgwexXD9uhS+I
0ozICiA3g4/2gsOLswRqFpRSrCtJZQ+dejWsLYQpJnZJBW4RQYTRFNC6anXIcOfk
YANnx+CUSLaOSZIhOLjmVgg5TBuTwwDtNjeXarIfW9qB4mikgHJyXGrHl92Y22g7
P0Yoc5ZRAiQBBTBx1zObjjS1rLs++9JrA0R7oKrLCdwp7fl3kR4p89btPxufje6W
VZL8c4cZhw7wbxphvJmxAlvdWdb/kzSwLGUrkVnoO2D62fyMAROaCvTIWCnhLz4s
ut/OY8Aysk2sNBXI+o+2BO67AqPTa/62tgia/9T3iWozFaKMo2UHCkyntc9y/xuF
SBsRlSqPlQ6SGHJ5XiJd+hr3S3JwYowsuUkHTc7+wyXAMNs18GUsOIfiL7Hmv0Z3
GrF2fvf9vWInCta+hNCfplRCsASB+/F82joY7/KkEbD37wSVhqdIa/RZ+ZLBAL3r
Eo9clacMjvQSwnAwKXg5+8mP3kWmwLcLlg5Uczsv5ENqtusc8q+nzQFaYKjpr82V
aBlB5fJFFzeCo3z63suEp4+TDE4IzMf5RnBFx5MZxoYs3uD8sthpbaQGXZ7IZWch
Tbnq3vuyomB5uekT5iU4UULdLmA+TqqU7V2dZPVrQflAIF6QaWSosZXgjPz6oHD9
aud7VcOkB9W/pnvKkgnlJCMU/Y0l168JgT7CjQmpgDEO4e7Sb41jr5djtcP7q7vW
C7sdCbcuCHNy3ObArJZek1aHM2mPxQ9IVUIg506+6yb9v8NCPGwXkU4stdFB1Ozr
DS3llmFXravF5amttrWdxwcGD7UZVVQxsv7wlrrRKTlTQXYvRBnVUpClP4HUzDPu
IPlUBhY4tl8yr6WZ2xDHVgv3gmrWPvRRcXxVikZi109gZsbf0msiV9qj/gyC3Fuk
cg2IieELys0ZcAXfueqLYsz5JVVn/034mdF4t0v5k5Bzdq5/MnHuADPCe6BzUJSd
ZHL58YO/DWWGHLF9QRqoWd0dPF4ZpCBQxDwbE/RnaExkxlsQ8eClk0DWx+9x7cYQ
5Pls0CUIi/5XUFe3nlbGYbGo2QymR/LxtAg6MdPxn3ehufwqMlMlrjgJsRYBa0tq
okf5MuTzKnH/USp7Bx5otrn0wgvEWvfvf6UG7EaTiU/DykyOFj3ZQpLIEBt7C2rw
1cEbvjpPegM3NA6sjFoMRbKz2KSK7jmSUIaFkK4bPz6QtmWSl8+BDnOKvxlsxVYu
MJ/i5clmrvvJqXewuEOTfgZ+od9fkLHlB2wsmyJjU1SiFpFk1iHanfLoYSgMfjUW
hcAh1tbwss5VhtP2RZrupmbAGotxyBuDJTeeBlLu0gyaTJTyzI51JjiauUgL9Ix9
7MIl1P931MX+oJI66+SZ3XlpL/g96YFu3thSfnVgaHE72V1ZIYtWGWCIreQIWN/p
L0PK+1cDlucs9jv80eSh7HU0jRQzHWbAdcXbTabZTDBFPOzQAvbe4ICTjOpmZalo
4MwfC0ZTn0UKwkhLAsBEe//LVJLvoNIQ3RADp4bn3y7iCIKbI64V+eRsJMaoAEnd
gFYQMgoR5XTKN6IiSAcxCR5ubbQ1Uc9EDZesOWexBZ2AlXKwssdVGbjR1LO13sCj
AqyX5IHntad1p4lozn46777r1cjFHI1NIhR51hiZbK0FuEm82nwzsfI8QXSiAotx
KmIiP2GOb7f97jCpZfDZJuo3ZEy7CTjX691XereeCtTfGIUR+J+MtvOec4AwhgNN
OY3cbNckohQ0CPAnspl85fzrBg6QVSCdEnpamXE8wUFxE7g6WKr76q/GxJup4GmB
LLLiTCwh5Uc8X4HRzueyCC7Xb2gGgEUobgUJxqNTQgZFJqWb0DTavR2rzft6kCeQ
AtEgOz5yeX59js/5mr/djIqPPBSmzNYNx70A2Ky//By1Yb8uLiSyW8BplCIyOp4h
vo7BGbcgzahYql2Rge2DhC5AjxKgfnZZcJglzjDDz5BfyI7T3aBWUwlyMgokLJpy
wjIXPx2NJzTJ6hn06WdJD69Ltxmk+Qv2sA7kcruxorlSKkiYf1wibl5vdenecLk+
eGOV7vtR+K5wic33n/eYaAQK6bIVWAujWklyDLrm/R4Q8PqQ1JozLmYH2OcziPHJ
9cCG1O0ArRXOvfQzbULPLkLlSHQmzn8lUnlM7Z1WOTmSV22w2j2HmB029YxdX1Xk
6fQ4qgKzcvWIidavkY4xJjGGv5O7l4Aafz7CwyoM7dfjeLnVl9T5oUwG1WmMQJP2
+haBSstdXkhUhUFdmt4X8Fjr10BQmTpbR/DqwIMt+gpJngGbLDejff89joZeXVlP
PbMIjgi4nOoNNPVMoCzih+WtrP9joaO+vTSd6o4z8yACwSDSnt+Ke8mThvlZMWLT
Zd9qAHjfnYDtowHaUu1QDlghP5Gj3/C4x0Vcuix3aZWoQbJ/fq7Iki8VvcR26Pwi
9REZzS1Sckc7ZYC4YQm+DKk+PfLSJTOSgWuSk8RkR2oz1N7D+chhg2nRf/forPqY
oC2rSkp3IoNAx172aBOKIaAVJQsmjWOpVG3uqnhAfEsosOvDdg7eacIKdARg5FRc
m+6PhdRKjFFQG8NCbXPO5JZxqJ3A4HDtgReHZhRqpstKQs2cRMNGNynWWprv3A6+
5q/RPE9XExw3lM8Q8kDElBxMNcoRnk0zJ35WwQ8zKkwOcYVM2svMmBWut2wOt4gC
PbnXRw4OumavWiMSBo/nJLZqCM/REbQfwGzWTKFPA+Bs7k3hNP5DcAh1LltkeO/o
+Auv0vFaAD4W6rScAHeoliRWPLdmH/ZoX5Y1RTn5YiC6DeRId/20BuxPdVDBYxS9
h6/uPH1wqWC8c1HLbCV8jvlIg2ADAsYb/A9Vxjm8jA2hkaVMo2Xp6VOXFlIIvZc3
SpSVRrwwyoELBuZ9eJA+Zj2cd/V/ivyaNI88DWpiKbHwyI96ZeJjm/HTE3CIL3LG
BXFzVtaW+L0PXp+P5ZFaH92iU4KXq/KR369mLJa0c7WvDcrKRyrYkVdAxQUR20Pn
/imStgQF1zz9fM0t8Wiy7crFrqAdj0cD3PhnLx2r7IUOfJ4d7O/DmNDUk00UUryL
GQI6O3KziUIlcx4b3yj4ncAD6+Ft3jYyvjIqdO3BIpbtHYO5vxo7C4tcWVmGt6yu
ERwqPzzOAwWiquSdcAYmuQZ8WPK1LLGudtCfc4TpPXYE68PF36Nljk5t1EanuFiL
T7JRgSB1hM9ykeELEa5sXEmM7eHuZP/0BsqlrSPd385pILHN3nwsd5XLVhA7JNle
NfbtvwhIxT91zPD76a2J/0dyKrPmrBT+9QjsN46iobbP8jg1FkZ7OnRsSS26C/7H
55dc8Lo9bzPOOObqX/pjm4vF9nxzGkiPm1TPBkv4AmcK67f4ioKAGkKgolrUeq4I
Kz/PUo1w/gOqSgQtq3F8Dh2e/7DawHCWFZgrH+Ws/Vrf3ELGgs7PXGMs3qsa8eb3
gUorSsAFinJ9r0mHFNOocyJ/U0K/YQ253Pg+U3bx0XOUeP+EbLoSYnsRVpWzqXNj
MlrAzsC50t0eT4u6mf2q3VgkfPHvPdiPd6Zzu94li0Ov3+B/ZH6iZ7kTI4guISTJ
ZykGTHP11k4k/yNr34v2JiAi9HGIFz8Ah8Dbg8zgaCpSl5c9D2KEkPsx4qPEmRmB
4/gHbxlxB70d3zh3tYER6ukUvt7CGspUFD39JRNY2yy9KGSwWQK70rF3IgpMlWKp
szF4paXcDo8C870AqlyDgp3Wc+BK+6jFxVpMivTHR8Vq3aEYnz9y5XZa8PRdGfFH
4iaNamliyQ8wMJdOzHf6qNBBvwXmw4mlrBrTyo5JqC7EoKktUCDGTQ1LtxgV/R3G
perh9Dj8vKZqMesZdxkAi+Z0Ay4gPIyV4Ka5sgIuAMauur56M5xt/6Vy3XFxYBfF
xRfgA/EcG6FrGYoUTaBpy0tHs/fSOxj4Bi4OSPFgyBX2HeupQ3xGCssM4AhvhiZ+
UwezV7vgSp9kWD7gxFk9LbUlOX2sP/MD17F6IGQ7B8h4T9AbCAMa/4NkOhuv7e9A
FmFIsxvwXNArI4tBURGm0pPLoB1ryTiHHkcNHVp9UaJiPvO3m2C3NynxB4LBDnbz
zCLTePgLKzxpPboaGAFP+CaCPsoCybABLRD0hwEEj1Xw/DPEg2FMCt9/vK4K7BcB
noyTn3S3kCit758YmClAWv5+5UULVtMsQjJKDQ8fieQ3ZW0Zvb7VwM2Clko9jx34
eCJe+AcpXezSGevVZLpL4CR0JE+Ibcz3b6D9S7+SqHQh+qv6i27wE3APn4jxiz/U
hHrlNmKlwTWkx9jTHnoU+9w/cyhreVGx6yQT3xC5Nr4NcedMTtTBb3w9N0k0GwOg
MCt05y57/ru1eyNKMUSUPDMIhoQ8VPa4rOWcO9cOS8QpoNuRaPG1YiX89t1dkBPI
MKrdFOGqRADpFYMiL/uV2TOI7CHHNOB8vOxWwieHQDye9IdxUcVYNvRbBIMTHPh9
rgkqb8ejHM9+zxIR44YmeErfMsJXvJ2oJx75unlf6rW8g7XDTme1MgFXGpiGK0Bn
Q2uGOTR1HrOpT5vlcQq5FDD6iDXbh9DM7Wyq7w541vDe80T/nLUtHVI+6KzgsBAL
beR9TJQUTwoKs2c/w3TW6LpEprLhncA7e8B1oGANzSeLcjwCKp3y/Odm77601dao
/uRYw7w7nVhZgHDFyzFCrw==
`protect END_PROTECTED
