`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eSx6qAmS6uyG7qv7mTSLl1Mn73UT8JfA+UKM4Yo3TKYvAwxv6jfY0i50J5Lv9erQ
EFBGHMyNdUXGK9c5O28ZHaH8W0mNDMdQk/PF6yk5d+EEXXeku6kwg+EPcQf0APJx
RolVxaTWwDiFipQz3er2qroPleGlmaCpBLvdWflkQlU4ch2Ijj9KdVZSNmJ9ZhwS
wtsjepQO+dkuCB8JHqyA04MGb+FnPSszdy0UfQR6SanVXlkMsEJwCrtz20lfuyPD
RHry2eS8lXIYptxXFTmmmukaRiTsSiaD7GuPlsd+N+pFGS2jT1hrNComQsNVd/Pd
Jm94bv1K+RXjK9Qn+6wgBNVRPyL4fQceDqhIT6CjBDz67XpYg2plSpgf4fteBWDC
mn1VQ+AK4FuCcJfrwZ0T5tgQ6QhQOBc8ZMZzRNDc8rDLA9vGhtsjjsl7OZjAx9qa
2XxrnDhGAx2r1PZZcwB75sxKMCsY2eIWkVLc3Zixnz4wJ4bvrueIk138Sn4SZayQ
NMZtI5sBWByP0g+wILoN4s8b3ZWxpDfGIbPLEYEvAfO+Xk4MREdJAqJ90rG1w6zM
3MncBl2jiopNfBzu2B62dyzNlB91/GxK9A8u3xrnl1c/6kYiP+NU3/Tdwh3ucMyC
WC8o3jF2AOsgHqNMVRziXGQJl2sXSCb9iSArErZqPDbXeKFoCzeRSokAfsC5/3KZ
5AmuybkKZI0AEpUpVgrkJdROTcJ0TR6DCX8MR2RK8VZHPPxAV7FNEzEOUSxw4TKH
wAaUNkR7+JZkZ8BkwnCWQP5aKp2NcmzBwpfuYYaD+OGjC8Q2MmzSl6K6pFWGWyrJ
D8tihbKMn3AjVnZ3v1xvKs/rrOfQF8c92dKPhkq7vc1mNaLyPWNnT0VPm4E0EJgw
`protect END_PROTECTED
