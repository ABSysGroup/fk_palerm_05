`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I+VE0MMbxJpKTdeO2rswINPGrmRa50fCjzZxwamvpOtYPA+/Wea9gDyTyqNtK40o
SZUsUNpnaNoljk9Z5AHYx9lelU82ppNsM37YWZOhcq1du1A8UjKTFBPvCT+O3GUQ
IcIdfaXI/PJEz7mOrh1xxh/6ZauPQnfym4yJ8RjsyHGPN5ifqghWNTNvPyAbQDXV
NnNLLBFxoSaolm/V8agWgouebCOFSHkph8QUfYTe3HVaboXA6ZUquWsMFPql4DMH
2u+zFP7C1HMZly8VEUo+jzWGOAVLO18AiccLKLHqCSm3XSNnMtRyAmFtGTUpLZc8
Y2R5MoVKQVj9oTWZ2Sr3hFlR6H31xBSL0X1hI7/fc2SMiHrSWURVeassOYJ0ALX8
jR7c5eOEHkzmMUvbmcwlQWJdJLltBE581r3KkdeQ8/o34JeNFi0U8uRzRvmYeM0V
2eiQz++W9GklK8XfTjhfH2wqeEfwr1lW13A5wJEPk+73lC46ke5EH6OzLAFoqxry
XSv1AdmZvI9onUofm216/011nBekQhmYsCLHS7dR8dn9dIfylph4DxUoi4Eacru4
aPgsHlqVEex2bj4EaSQQEJRrmYFMpaRcBbrPf7WZi7OvxWos1kVapM4cB/U4Qd+x
X34yg1jCKm+lQ5uri4ard6whcQRV5tmC9pSpPWQiZkk9epbfGKX/bLBRDoBzZTpa
F7B8PfODATrfhDBaTy+VNtwrAEb/n9kXax7jG8uYdVeiHQN/sQnEX6sv7EJAb2pz
dzqBPD4QfFL2KzPntIOpFA==
`protect END_PROTECTED
