`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Y42OFM+/p//ZTTTOG/f8BRtmGDbUajA82M/b4V4aktz2oA/F+DfjxQ5N/sqkhTe
t6Lw2d7Syfx/6SuIaLG5o3/jTbZ+X8qr7bo/C6xmqnLhZOdMT/MuFqU4MO16YNg7
YS2WNOIVgaB2gYatc+eI3z5D4RL7Tm8xi+0pIT+Jlk3DylWIgtrschE1UAVtXySY
hA5SnjMv1v6SsrDQ52gPB4ha/EktY+lkhQ9KuYmXtD2abYZwnwF4TbBzRg/AGBL+
MLoXRHZa5MUHA1d8iFAoUa8eWo+8oIvwzXmXlIMRR50oZaZtXMSp7P5sb8Mk13vZ
HsC86ViJ+ISkJSqXJ1Nc7nBnzDLYWykgEoNFewFiCnaf1YZ8h7FpkskafpUCol7i
WLeUkFqeHkm/k4/9M4Dp84NDN7iC/BmGdIZw2FbTSJwBLTY3+Uc9zZbr/TEHlCrp
MVICozhlVMIno1ZOMFCkqFGszxYY7i2tDm2woPZKB2YlCujMn7L+Q7B26VBBxD0J
hEbiJsq4hCKwtR6UTo9bcYl9AK33oIKavgLXHWUC3nhKLwYcaJvc19wiz5UinBAz
H1hBsQF+leGqxmmEHYmpAJiX1/H618BMwuoUrVi1CeR4Pbk5R8wMEuXuMv6xZUBC
fMZGlVXQDMpWrKgNl4VO3FAIPp3UpbQYcSXCLUCDfjE=
`protect END_PROTECTED
