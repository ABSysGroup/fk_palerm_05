`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Of6U4VApCgW0Nwi59dBiJM0D5oCktiliy65J4qprMX4bGbxlM/cHgh0Vl4aVsrt
mRSH5OFTUI1EhNudBl7QtXcPHIUjjjUx+x8oZ4ooI8kTLE6/LCXmv0lPV9kVn1/t
rWanETM4nNVgzByUHiUesn6EkLjk4lV3LvkwO0WEDFYenWIOEr+/UOqmFxyE+92p
xIt7HwyPkCe/0pkt4iQ3eE1rFwWsYA25T/5X1oGxGyccP1GMYiL0kFj6IzZJoCUX
EpdENWnJz5KQdRkVSj6Eb2sIsrZI8STmsH7ij6TwBgQ=
`protect END_PROTECTED
