`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qG9+qe6GuFuH0BjKKl89b3W4DUbVrGc5ZAGbNsPLew1d8cRkNHjoIL2EAMrUlPaP
BpYrIu4mF3lMyR8xH55WTs1ANFRjqCFMaKzUdXjc5GukTP7TvN0ouqY+h2wkQoG7
/hmbVm7jo9NeU7o9fHhJdQHPmGFUY005Z/CBzxmGrcmuvRRkQnnsnaqXb82xGctn
g4xlYGUnr33s8NG3UEgMzge+bYO96bzqi4OuWC+GgK6+LKh8hDHC36QGvT/rOW7S
oWNroJQBT58NiurQMKQk3MNZy9bwWw9/1EodbYq3wjMfdk3ysgpdPX9z6370Des/
4QAwntEJs8R420SW0y4w62OBeV1+Cc5J7eAN3tSl2bluruZmpecXvytLKAnyrq7d
WumEafLWXwlUXHGSA9ksS/jr/Sj5WvhUQhBfYq0bU576epmhkvu4wnb96SCh0ub0
XgiipS+ymSjCOOwga3c2JIsb9rTO3jgiVm32Q5SMbkQtb2QL90O+p3hSIe4lYu38
xXJ+cRbFqXqRBK61r4RufM058U2TmL21o/dOCjjNTmo=
`protect END_PROTECTED
