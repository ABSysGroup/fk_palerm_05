`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XxfY+NPdPlgJlrW5z9lDqMQDNCzVW+mLPkKS/diFc7VWmd3ZuPLCavzos4eAVqtT
zu5/yiHngdKp3cdjKOFYavGyPqVBO+j8TyhFh2nM6cAU8Vd49RUN1efnFuA/Pc1s
Lz61XT7o8vQQ7wq6hR43NCGYXT2sr4BJZfWtFMwtJTm/JNtYEJJLVYba3vUKU3bv
7yPNEbZQ0IrXjNNYace8BvShKOKQnQFJx2Bse1PpXxZeIj7GqiZTCzR47enrjSJn
bnxpq7ZlVT3LEhszWbLulbywiIerjyvh3VjwqCVZLb4cIGUh+ND8SrJprv+nkau0
0P6vuVxI+DA+BBHxLPOwYIaUzbCpZUeYQ10JHWmXpqfiJXY89bbqruoMaG1UunN9
6+XmFxAgsk8+o78XE4ArQoarGb0S+d6TQ4U6/YqhV6LxcuZ/eFzhsRwTfAVS8hJo
5ucsgPUvMTZeJxmrKe1RWYAqvqe1oYy+cVA0j/Cd6btH54NvCyxssvdnUupeYHA8
cDKQQkla2KpzahB/3sagL3T/dVIOsqWO149yk7s9ijzEybJ68c/ufZgwVO+Bdxnh
/n0pkVNVnbk9n+uoset9wV1jN5k9556b364WVICVhJpSO9WdhlmwzstW6nVCHCJ4
MbymCQ6xDTaakZsBG0iFSdqPddtVFW7hDrzfFsDw92Zo+3aQdoBwreTy3qrK3yHV
1Mgl4q0nXiLHqH8l+rLtH2yNriu+9FQVTC2mFxBm5rxEFqkK73IqNnAQFmerSD+V
xQmLgbErEr/61l13W4rtZ00hjVg3dRQbu/qM4q/qbqHQ2BvGye/2ocZCPzh7Vdg6
YL+xZjk8w75igHl2N9gYpVSRHkhhGJkO3TDR3hwcV/OMLrWaHCUhPW1pVD8CTIb2
ffO4rjv9A4aoQG30wN3kw1BQpxOVLhmnIW0tn9iocK/9uXgxlBGfScN9U3+LPvI9
CWdIfENuh/XeKacSBXnPWrnsTUsvoa6Qadi+WNVR1f1YuQYuL76Q9xkLPkqdxQ/H
yg65OnHux3Hzo1bDOMD5Z/vesHgry+N17zoBfyXgtCCw34muDXA2BDukSP7T43Fw
LBIZ5r9bczNTMObJE1ePPpiKMyxEhjZpE1oeLgjtlMA2lph/d81DDPSRZUr2EdPq
N/5Q1AW3/3WhaSnEYcMPrIn8XoDw/ge+VgKcaQR1mJ+0sDMoaHNMciF1aX71saAD
YYwCZh7ftQW5oDB4UhwrmEsLCYKFthEkIZ0aNWdEFbf02SOE2/J1RvCJZykTYaqD
NfToD9IK+zSN2w8e6bLiI75UfWwy0h+Ymdmz0svZfho=
`protect END_PROTECTED
