`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fmja/JuOWwchmawv6xA1hZ3GDU5L5i2qsWDZpCYcTLJ65+vYr9X3JoymmXLlnzNg
ll73x+fPd35V+PbG2d08ZV8IDFTONpwZkqw1VyKoeo71/pJSqUDK6QcMISgWH+at
moWKJWee9LDGOIMGnkP1vst8zGMf+suefO/u+BAuyJaEKOeTvSZDPVR6CJc2uuSu
YuBI3+cgP6GeKvMD9rZe8SUOSLhg8PBBMKW9VTLzFv0hofvWgAhwBODNU/cZeR2P
+1KvbFEKS6ayBoaxZdVFLNXVbRUNRXJl4tdFyjY+y37K8zvQzbyQbJUm3TFeZMHs
OgWDJGRuaX9Et1v52jUL8cXAG7feOV9luabpM45byn2DMFuAHhF/5ijCuahtESaB
htddj+E4C3cWNT1jcwL6C2Lu27gpXAaHQx5nUykg543uekXg2UbSiUt6jyLWi5pp
E5G1aeet+j3sqw4CLiWoV4667p9vPYT+Dw+cxUdIHPdM4hUzsCgLdf7o3msthdld
jN6Nr2RmowVROHlnOguquzaHQFRU4zsc9PzqP7JIHOK89ukvrXwSOsXOvhHvNVsB
WeS3Py/zH/8B5VdMuiqekQ==
`protect END_PROTECTED
