`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nu+UN/PsgaREHvXI5X772+x4xUk7dVgvF4YEbakgl16RfMr+yVqx0EoD6EkiV4Te
ZGVQUmpbsfzPY+ttZrqw5/qnvAMkE7urtJBIf3fENfG7JpFzge4lGFLaDnKYuVSR
6PSoVjXWHY+SHaHxfFeJ0viIyQNzQbT7qT+XQWn2aRRbHhzzB/ly2k430E436tax
1MbKbLd+NeJzOTq4XP8UpYU+RO22kYzEosVAK5VUojD2snhpYYHa44r5KeQYQTqG
b0P5srHmdwh+cTlddF/dyL5Yxl5J63R+wY27K8LnF2Dt0Z5lnOELOgTqxeVz5Cjr
ejLwDFUMWwJD8MN+DD7OZSLl3gUFfg0j6/7eCotN3/HAZpr8NxYUxeMfZ0VvYLg7
jMiA8z2H0PYAcb98s8o/B8J5dV4BzpYCW4pD9ISxHovDCDk4r/XlG38mWaWeB9IK
ja4s8zvOoVbS6sZk35/3knn7WdXg1S3TfGbjYM63x2DBNvxZPfkqWFmUDb9T+NIc
rrcOIWtNDI4YB0vJo1tl10ykXrWEPzoZVMrvrfkXbsBr2WJOHTWtKMl2zvuZfNim
SL/s4GcNacI61/X+B1G/BdD8qtpRMDpXuP3Rrt15gLu5iFgqRiQH3vuSg0hk2A0f
McsHrC8RAg4c+7QH7u9e2g==
`protect END_PROTECTED
