`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8g9GAIhEugdJS5selr+hhy/4j6L3RgedgmeVg7W7VoqxjG+Uw4QDPyviE2GycDgI
Ouu8A0JK3GNlXM69hRT9geAYBkT8fiKvZQx0dNz7E00jd2HLYzsr0aQdzxuCHN5v
FW1LbZW/zNMlt+NbFgJZt36ieSUc1Nfo7rkkrs3sEyLeAQf5zcrzO1BiuDZL05MY
U0cJLrgq0kSiaxjNLWJTwMQupQzgQkrPg/Es/SbZNwZ2Bf1IJ4CUNfUzcDRn4/Zo
`protect END_PROTECTED
