`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DGcQPqQammTuJz/29Pt7j8JitcfNYQ/98yUilUWGh0r19lilSHuEKqg5AsUra7ut
eZ/zKiAGw/g6o5X6O7fuo4IRLS27KRUyENZFwd/Ga1/LFGcOuJpgXK7oGdQ9XGTj
UiBgUPuhIZLzdRSx879LeQc9CSj1emoamSd6TIFRiXyqEGG9NOzvQbFIgqqlgIOH
wGhsrBQRumaYwPQUZJAaAu05rSVP0pPzNRGCUQbNQ7+AJUjAok3G/RvwEv8kfK/0
e79Im2X3MWaM0JxnbxDi1E9eLdzbxHNiZMPs7P2BJYI=
`protect END_PROTECTED
