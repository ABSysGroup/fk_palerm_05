`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h1nL8CFEsVgbU8e6zc91bgsZlTk97+av8UgOTJMoh5S7P+YeAvlUB3Rg1mVQPOeB
lF7gHW42/l8KWQh3Ef/cIzhcHBsW8VfRiAc8MlHL0ElkjDC5KP2UWu+Jj0ENDW9L
d1xjsO0dMK7jPHeT+lqQ0Wz4NPMQ14nu73HcI2iZJHfeUaLyDNRWy7/hUylsQFSx
pS/iGUyAJamdPiIi9NDA5Vd7H33hk1CoYfrSPxlyuEo1GvZi7b9DkvW7Jp5V65mY
J/ek2dgSU6U2330a7zYs8F/jHTPwkzRwmcS905a1yF9MbRekLGqt6TIu6XWfVM+U
N1VUFJpa0B35DrEAeivKWLOpylhc2D4ady2x2JUCRHT6bRdJr9WgVip7HByYsPPp
cGVt+Bi72Okgk9MIzEqtMfhLX03xxAwjLjeLXqf15YFFWX9i/1f1raZasbFemeNc
3fWka12GmMGZW8zPH8OwF8lHZwXGPHAL6N1PKeNOF/UELI/kGMpY5828k1GLNc0g
iHuV4yY/ed9pkbUBFA0gUerxk5GGFQbxsjCegE+YnItIOieIorcFIy3RKlCZs0Gc
s5HUvfvPydw/5L+ep1d374Q0TtLaduQHTGjXraBSYOeXKMZsu53Pu8aM13dcbnHn
7bsLVoapBIUD9hjNz91jGytPGU6Uv8Q3HSj0k2CNAEJuxhY75WpqSx3BUItHqGDC
56MCmx869YqOdCSA/IR3Hzb55+QoUXB3sdu+JpIQrxn8Xxtn/lFqEHkAFTlviflV
x952po839JUZEZr0zNGsF/bcDyI9hsv8Yhq7kpS2D3g=
`protect END_PROTECTED
