`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RnchtwR2xlTuBVzF1Gd0J2B5X+siu/8nNqT/KWq61dvWqvJyKxiFIkzoVco4qgGS
ksXyvfOqzh6WqWIuMxnH9gy5eCcsESuOMtkW/b7s0aKXl/CKPPPGKknJut8lPKHT
c6u0HCul298ReljE5LODh3CY9trSuF53pPH8wxkZYnPUYm2rz6jbSnHbHWs7L+Yt
1Kj5W/7nfiGO8LWAjB380TpvLuiIV2Ilb1e12rhRiQC4mGjfBFYRwOU4CUFEOHI8
x7HwxwWYVsDy2mEQGZEhIsAnv3suyAfFt04biBiL8HF/hHYSypRk6WYRsc/casfw
WtIsTEiowYmTiKwb0Doj8pVmdFaUdUgYAN4WarjKLny7PbW6ezPKTZfB22D2xlrZ
Dsk8JGgzJAWeFm8hEeZyMRgPEiZ2rmig+qANJaG9oLviWQSo2WrKbg0DQ74V0cxF
9qfV3WhJtQb9RGCxKGMw9bDv8tZMYYzbfeZJdkNEVYFG72npjGn2UCUFZDllZQ8p
CXVsj8KGj6lZwkpP8rvuh0Acd5IuGMn5ydxNlvCTgNAWCAoNFxpVLjpUp9iac0Kw
CrBi2joYQijXWcFCvI1v1SbQuWAye3B8NGtiaSGXHm5MP+s+v3k6/YSWyiJrckxO
vT1sb+2+Vu9uvObuxocDG6fPP0gNwmQoP7vdnq6K/dl/1pbvBawG/ZS95eG/nqmA
S6bqu/DKj+O8pL08VWYwLQ==
`protect END_PROTECTED
