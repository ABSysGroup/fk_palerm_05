`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nqzn4lXg66hseXGu8iR+37pXXOFVKmL2++QmdemjnWy9Wz/H0B/OGEUQI0X+IhPX
SrpX12Sl9H6vQQAzbj6/yZaUOpC5XkPER4k+fF5YYguJbUwdcMxf6ySxRdwmfXXj
dPCDBWR6zgbanwqKkCgJn0X9224mDERIDs5RkQ0rbHR17pW1YlQccWjc6P5WWEVI
MIKKJa9jhz34FJI7O0hRu5GsFe2qB0tDdWBeqknb42YvHQYPHVI710sCnLOb3v05
Q5/AdT+CPo7vqFeDWSYp6sdRsY+9l3+A9oaHpFWoigvTdyKEri/ouFU9/TPsXCm7
pCF4c556RmyA3JyiGpbdjs3ZnlZG4KUJsyhqK3/sNC4r6dXEg/VY4kvfG/taJY1j
xQhYIXTCzKQCCdM5/nMxsBeL82Yd93A/pcu5TPKHpNegFeU0fojwZmu4xilEt8U0
eKd0nfxwMocNa1pO4O8JJ4GLIxhXStBLhv45FGXh4y5AbR0psP0YdWFPiFWmgoH/
gkDsIso9kmuLL7lVrXr9bS7+InV0nd5G/grYKRZffBYOy11+cZ+6OuI4h99edX+A
Bxbgc1dOKjMvMYQZUM+7XG9LJFoo3VDmiRDU0f6XvPM3Q/e+F4YspCjlHl5jY+d2
7qtED9WSWQN0ZUDZjEStGLez0IYQNuvHw47uJHvGOiJ8kTcCFK+7DiOyzDGbA6ww
2pdNzUoX/QuGmWgPn7f8Tv5+UhJ6BkQ/vaFOI1q6RVDzsEDfR3C6r4nX3FF5A17i
ug2PkmolOKb7tgzs671K7gDQlCXxFr09GiAQxL4pewcprkP5P6rTfA3dWnjOmKIC
`protect END_PROTECTED
