`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RNgG6vlYPSeF1sfB5Jgfd7d0urEYx+gdyXnB8/emiWCadPQYBg8p6Bjdc2Zvzkn2
VpmwHGd38hO2NCISWOBOQyIuOAMhgktksRtZ2bH/LiI3J1TujCQBvvfv2YtJ1om4
qNNE3qpIrAI6Zi3Sl8Cc6QkNPH6FTKRd0v3h2ZhJ0yA9DFgG8MV1A2xwtSyqrAH7
Cj3NC8upgQDSKx3PeMw0sA+DBIbp/dFoxRFdmvvNpl6yAoLX0/rCKPxjJ+zFOaEG
NZ5j5TUl5UHkDN0Q/vu2OHbIW8YahJSm8lCoyEgFbrFQWyJ/GMIQ8d1cA9VJOHC4
PcQOaGVm0swgxZJsTajkJg==
`protect END_PROTECTED
