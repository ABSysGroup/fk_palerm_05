`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kd1MjaftR/W8A9kLhYzOWWBam8MVYlqXf7i6BgH9J4a6G0OC4AA9C6o9TWHouA79
uY5K6BQhPGoFF6+f+J0OLyeaU+tE9SQpLcb8/DBfS0q+CWaDWg7d7h2Z3ezeEPgF
4j7K6ZkY4tHatkTV+3kpiq3Ry2aN1GOC1l72AuZKqaCHFZDInMbDUxBDCGfs4sdv
+lY2q2cIloXI/6IyzTE1Jsy9TYyJH77ZRf63elwhxlUu9zGG70SDLEv7rWPPqIja
kQBjTHwWCT9hqVd2EPpP0KSdlWwdp84L81EZ6f2RvhhMD+fNHh3xUP3paaXGm8iO
uMYW6GxsSVpHtA/1AK+MmuYGHyhvIflmISCJVmX6VJvtezt3/U4v+7juTGKlS7MP
UC8PA3W63opBHudPQFXw68rZN5dk7NfdlY4PScOHQfMn9NO35322SoikBrSkpAOx
`protect END_PROTECTED
