`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9h1w1VOWddVoEdU26XKe3mJUD+dKtCvdbL1AdFcSXuGediORocw3rqVOouG634fR
BtcN3hRXYuaJnn5xlCjqyGrOP324KlP9W2MGaYmMJiZ4RCSFp2dekPLsvC9S8hpG
DAdLrgNBTJ9u+Cdvof4CmoKyjhsPAchq+FktnfaRzkqnaCFx/gjazi24hNaCTvcs
7eL487RteZO10wpuW6aDkkA0JlF9XBrltSh/UM6bwyqrBNaY3Xk6gR1z8G3T/P5R
Kunmi/aiUMZmoOc0qdU7Ru+bRQGyLW2cCQ0ofmACPkh87VSMCys4QoE1q5ghHREt
qWgwyLNr3GqNkLTqpa5ZZw==
`protect END_PROTECTED
