`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u0ck3Z8K13mJzrLWJA8josmRmduNwgdEQNCn8MQYKEEPTGVLqzTks3SHxF9UEfrD
6WrMVGbcPC/HcgDvZeB0eqz58q+fOX2XTjWfzglnUo/s8DPfmxfAIqxDun9NOphC
UPtLFkhl0t8Kkm8JFKb6DlRP0gz5D4iqlcSpHSHPoimwBtv3zlIirk7xv7iLPZt+
d54q9U/iQF+BQ2WsemEx0VktLfKJmwi2ksBE/I+/WxcYUEFFDUnHbJtS5fCzPqio
tGuoVgakZ/+vfjRQk7GIxNYQRmAtf5D+SMNryQYgs4ZLuxmZpH8dC1TQ3KyQ0/lo
Xi6CmqjkNa3+nF3Ia6BqrWTM74xT3YCivTiIAwHPihVx5nfUxdTNKmJgADfgI0zP
IFvbl/rY8VM5FmTP5tPXE/dY7Q/zobx6X0QxOHfjr+SBU8B6TdNNKcPGd0H1gGal
AzdKT+tsc3358J+NxXHF4vVbAio5u6C2wW5grQxqD7tTKHkyPJWGh4peozEg7/Kq
/PYo71eOh3OcrzD3UOHWz89PaZon8NcGFGfsSS8LrIKh2WTIllAY/6TZ6dhPMS67
OSnHf60Jj7sDj4xYsCKf08tkcZbzZoLsU1a+lz5VOfwlxByX3opBbVfXyQXDsUdN
eynEAsLK67yF6Jf2MHFREXOhLf6OwC3Ejx9A5Prj1Y+Wtbim4yI3zY8i1JVVc+N9
xmTM5gWH1Z4ZMRhx0MWUReGK8n7loa9voG5SmOPCzDrwfYxXAesn/o0R5eJIJra1
8osz4WcG3w7Tu3fTrxi/iz8GoezcBPEGMNM0qG4meQ9Bv/XBd34p99miWTO3MnZ0
0yJ5K9eIrzWmzbNopnCL+sjHamnxX3k8JmL4eED1W4G2ZPcx6D4XE5syMMESlDaX
/mcIcCr9dsXnFEVGyoo99tEFwL/prWjUx19Js/Bb+fXIU4eS285nVCVJ8QEat5u5
aMpJNrTSIgMM7Ycw7uSndEAQHVFYQlVjqOY/RjLQFM5gBC3R3xBWJlPf+nxE+ULp
hO6A+fHaDV4CNjiVruOV6oEMn67jHdiL8ugyTERwN1YiDLYE/ly+IJlNFil9Rtzk
/kWZnS4F2crrzgc6yERDUD+CmLDcWvg4WJYx1DCpTiCqRzptDNdv+DjcJ/0bAZsy
OoqGIRKpFGttctPwQTNMjfoTj/eSm926OeJn2cwJYJDqOjIbQ7vM/QeGQ9tsPgvN
mgOJmcCNhMozSKHu9k5/vAJ9qdG6h+aBEu3RCU/PykI2FmqkRvFSeFvEIaKfdU8h
GBRqchEcUKjZ9YCKyORpkmz7hjKfUOCmivikYOI8B0no+W0BIWbkxy/zHHmyMywU
tg5qmR3nBxWuMdW7iRiK8rLt5zUKt4QNHdyK3We56hJb5A6xGiDA8l1fRuD05kIz
jpiM6nPeZ/O6slQGRtBeJa5oOe9rgdDJizqjPOJkNIet/5NlhMBNX5PLze+jWcDv
QlnFcJFNRaGKloWkObVO1gI9aj//rjf2qxm4Wdv4wKXZeFqQhD+FyAvLPbcc59kH
JudHO2rY89rc0GRM123oxxPZWzLfymQiOM0TCTk7mMCF2OOdBwHEeY8sx5wfqj9T
2JJ8sGjlzji5j4jJiAiigG07suwatQvdQ7DPhAADQSoh9kBFjchfpc77fpruG7QO
S7aI2jAuJgVTZnpEj+2iCQqDYtMq5gmWpSvNbfa4Exo6bU8Kz9gNav26QdMcrFCs
nZ68dy2cdWYSBDFsEnDg0QalmeFHsao8xfpNJc5Bacd1GluTzXp+c6umVLctnFvL
0pgoWKTtYtpj7JiSD9MD1QijTgt0FMm6ITzHZPRup0AacKTdQsWf66xkdz7FdTwW
yfah8f6aeE+CogUhuzCEX9lyxco7oMKhyPWpUEB2rX1UrQaZcvsT4vCfnnVI6b/Z
TEFBP5Dk1smH40c1oNiAFuCiCKFHsChQE2ODj62pPE0o1Ksn87qqRa8Qkij1oYKV
nZXeoiUGZY7A3x3B9BkpymrRsad1BivqXmp/FbsOQD0iKVIBceDx17cS4bO/kDex
AodRNlSkodlAVVU741chFzj+WQY6Z5N31RP/gYW7T4kb7A6RjpWOHnRfh4CXTE6h
SBPtFbxbaiPb864PdEY4BA==
`protect END_PROTECTED
