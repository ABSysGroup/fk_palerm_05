`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OqWPZX/PmOEDuTGaykJ5voLtS+bjkTCUFwFYy6pFYVnHA6L7pMN4HeoYNI+5rL2B
QDsasNKMMb2olCB/qXYb/V5mPYm5bX19MP4+z1+PmVrtemtsvHLBC316jX+qZnt8
Sqv0tMuXn6kWVykkbnZOm4oVHBzuERG63QEsX6AIzZPQNMcjddSUaqVJNYxoMD7z
6EcgAjT5bIR8lRXqb/dXl6dffspaGiFNxqCs5t0zR+smPqojYXw6hPh2khRlXMNF
o4XjsvgMDsuCQTSdfkIp5m2kn5CX8iFc/eR1ypZGzXAKCZV0Ake5oN/PfJkqryIq
SoXFlYf2w4GPmkGJ80N1vP6sbEGbVMa8P9wmfTUT0ft5hDQ4FF5QXAm5JWtnMJYm
sCbiTQjdVL8oh7bhg5mkQ6qoFjH12l2cyzlMIsKE4Hz6d9oCbZsPHaFyrGFuJIqK
xdu52/9O76WZxjyiRMva/BrnKoyxsBjRWG5vm5Rni1s=
`protect END_PROTECTED
