`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZPUUWXr0syY1iyWGeGfbqU2cHGA+GKVLK7pXx1AxN53+DP3xfzrIHdvzDKggEdSb
YdGku6J09z4zYrJx9VGnOu8uu+FeGy3H6Ci4pDE4U17N2hxJ/LT/JoKcNS4WNeLC
lZVnKH9Kwuq98xeDyh2jCfWUK4MFd+b2MhhhbVpXcqJc/dgq/qBpefFLkbLaRUmr
4V0cNjfUPgguqXqmW0Z1G5O9yT/2aU2JHG7tptho/o1fNGBDyVwvTB9EQI1+LxnR
uKSuhjaKJ3lFNlmWWJunSyP3tqPOWkcmOOp/O8cclqX3ENJ3u86I4iMecWB7NU8y
L94LfGlBTlSI6rp/glRGhOWRzCbh8jLF/o1i58wRfCnASoAUhKBKhYT7MUfkSBAb
O+AmX7RaPb+uuXfUH0icJnWoIs8p9OaT3hUUcKxBtk/UX969hSGHTRXrco9U/sLL
qMR6IrCNONyxr0yoUaVoJXTjWkr8FkqYVebkmpYjgTDuvgiFXIBpe0E2S5UDfAuW
qRlz3rqcHvbzzkl1cwqrdlwsms/QmR7ZoGSYyPuVeUmcNlbMdte5MzMu0bT5E1Hj
I9U2DLI66FuMxB3ps7KLibS7x4Iumbu9pbPkkZ+fYI2LdDSA8lTnYLnjpih92z7M
vO7yUHXn0uYZx/T7tOSJbD4t+o0Zntywhx/kDI6b95VscduinpaaE7XWZevec5BV
fPhXyyMmUKfzqmoxSRaqEzTkNVv1rALyUDRiP/YiPv7PHVGze7y6ygE0f/3s5BT3
VWIXnj1b99M1NIfVkSob24einwkomoy5pwUQTJk+EkyF7VpuoSEinZ5vS6PGBPU3
82QC84BhulY6JkcWjYHkYFD0spk5lmRHyQ1xdIuAKYE8zZheO5OYcGvoYUK0QabK
/nKLp46ePPA8pcOyqOwQMm5oEm+jTHvwdbSqn911kA+jO9vS8fBIkrx6dSxOy3z4
XSq5iFLk7tvy+tdv5Q903m2BHTH60rf2mVr+wAyac2PRJtwLA3TtDT373eHNCrK8
9PKwDruD8N4glQSM50S+bznnqURhUT1CPOSJmJKC1iyUzrnhemZkRfFn46i/WWgo
f93FcpBhz4CUPFqG5CQRCRk+57xWtAy14EKn3s+AIlj8KwJ6CxrGmpVw1DpEQzkV
uRdRF8WZwi1kODyyR5DsQcuSuy7S4ey5HDSZJbzp+7xD9Cfu+LN7FbjUdJifwPgP
UQFq4mQGbXQJ2KmByMWEHdH2BG936qOKaoEE0tbwDo4XgctvSjj0kbZwP9pj3MfC
PReeLYHlY4f1vZhc3UxZASrMsqblmza+z2V4BGhYehlb25yl7L3GeofPqewM8PDH
5Et1o0/Ni6kIpzzgNKFyc409JmncyrLQv1O/cXsfBUmK0FWGjCb2ftaLxkcCQU8E
KrDDkACFh2i9tKP/zTBF5yRvnN6ZdQaPOLELdtcPyT4rr2XhsJwkpx95ZD0SIBhF
7woayP+p12K2wVuDquil8zsqeLyRGRtpTE7uulaXBV/8Y/lUDq4h0UXqQOFCCydS
TkaspwcAPoGJL1mA7qm+j/tROMpeS/r851R+7O4yfSLQpJgALKsP+irTZZT05VAX
ehkClrjJ/IN5RZ3omB1+nX2yETR4wuzlSW34WFYp39MCok4eR5Ob1T8aUj93TQS9
ncoF1CJ7W1FraFV+lYFzwabf3x3WBYXYeTfH+jJkV0FnEU0gAaPl/+ljwmp7qtj8
Vym2L0l+8fiqfqHGwREhVuDkP9zly7Ed0Cf9LEsCbVvDQhjMeryZjislxzMbjSQF
3OepAXwnUDwhmzcLV88vPrzhYqTviTL3ksilvNuV+6KQmP+KKWbIS9wTZXCTSlNd
j0vWdWicqH9+6B+oKHNZA3V7MH62PLLlmzNoWst0Sht7XuwkRH09G5oH09ARGshR
gfkS26a9caIQSPLRiCEWFfxiFcEcZKUn5GX7PbdSB/mjIEDXBPtCEH/gMZYlEHPc
ld/jhRigInQTBTlY/ckYJvRyO6yKVAgo9imcEIBtURy/4v0xwEcgsHpOXTKMToKj
zdK9ZTJIrgjySOq2EEEqdTa3f9W/OWxLHeLbHTO1u6YGsglNdT/vzht30X4tpvqh
Z1Q7abXzyxOwEWNZVTfWwFD/Lqui8y+VyzY9n1TPSzzvmVoB37ME6m3Z4iut/IwH
iQ5Igkxg7OIliAFVhQdjPnOENRn4e2khOkgiXITFyoWv9npQBHPVwYL2DDBjtWu6
/00kqrBFUsicxlmUOzWy1qDXDga1SjbJ6se5IJehddJxy4uou6Pf1xJ06OuUFvt6
BG4d853BGXoLWWsGBJcv6ZKhhy8MgWAQGE/JJKObXkr0/xeWUx0ZKEpsYzj/2rLs
sfEqS9mBdA66iseGdsAvNEfmEhhaub0bFMmuGMQHKNs=
`protect END_PROTECTED
