`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bv9F9XHlpeNrame71nxBI2LwrWHba6x9qSXEy9qbLNT8yaNdkEYhLmPqtyRVq7lL
ZyoA95+xQN9DvMpAtJ0vOaq35SgotsbLAcRDr490VOe5smPU7Nl24loCJYPZ/Oz9
F1JXog2bqYLCJL9Cr1ZYLSq7OYiUj0P5Mvwi+vuY2qGLq62wC/jf93Kg/kKztWEz
1IaAv0V6OLehphVemrn9WSQ5VIuNREDmJqti41j/n0OgngCebjRhnzWyz0TwYVHN
DmgtH9OqKI2XcZSUa8HGNUXdWX/NlXJ3FG6ml5Vb0RUK0o3CkmjnYf5rTtYQ7Wft
yONheYxnj1nKJoKzhovfuDP8hVlbjZR8kk2/LVEQ3vZaittscaru2ySxuKKDBtOy
ah/mH1axtQmZ9RHhlcXK4zSiZ4wXJjYCuLdfX5x1R4d7i8CsEKzsKFRp5bR1OJE3
8r2vJUPKrGsOgEXmfNAGkUqNZfQpafevw5+7VxM8Mf9/QHqX+Nn4PXJAJ68IXuxa
GVgBfjTAOVSHOjnN69vlhFDD0jYvP5QbTdQJaSlMDKPSzykhxkDinFdBcSBwdl1m
ilKGq3kisHBXOEcfxvZIRVB9yN86MwSXgvWBXN0AH6Cz4XVqDQb8CcCyQzkF+X8A
Vgpl+NY73aMOESHm24W05YtzfwGzGkTGodb6PL5o5tVqVPmuaoHscMwrn0fRRbiT
btE+P+16ZH0STmVwKJmO0Uyx6qz0VBaqgqlZO0RMF8DjDBf3NGV0bFMGTP9aMQZl
7nbi9GxBa/MNMOU5Dqq9oA==
`protect END_PROTECTED
