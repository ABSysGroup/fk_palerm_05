`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u5toZRt2ZQaz9OYhDms/IzrUpjCIItkgWnXP3DdI0rsi7nZ0tj7c+6zHdCToNHMu
JUPyF2bJNc/Oa7p+L018rdyByJz2rgFE0B0UnFAeIdqM/+kQkdB3tIPXMsYVx9w5
FXd3uEolv457WwTW4208GtQi5PSfjPaRamAZFLk2iaEGu7J9QpgojjdTfCKc4U2F
hH7Q9hswpHcExR00dDck5+BWPO/m7IG0dl1d+aPar2etdvX/NcFQQcY9HJgKgMMT
`protect END_PROTECTED
