`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hWc/Qg3tfL26/DqwdkdRk0eDGdIDwR8ZKOlQrIZFCznISund5i41WhYzMQoy416X
MbcwGEdVcPN4ZL6H6EZ8DM9dqEYmlPhzaIfSfPAZ1Q4cortobAuo7AiFPMtkTKe9
Lk8Lpib21JZsdEmvoUqQjpWWn1QUq7n5hKxJnYWMucHApRF1E7T/7tBDlYKBt3D8
O93yODOVUD8R5wsPhJ4GXPNv5x9oKgNpT5iHjM1WSBhUGwZYwB7GTTF4ee0YyeV4
1QXc025KraEDkUvL4dvCaFr8iHOFpz+Z2E2yERK27IjfXd4ueaVwqpvpSJXp2EbV
kdE32EDEl00LASDhmZyXJA==
`protect END_PROTECTED
