`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zdPjki/M20Cap26PRY8NXaerqF6iQMEs4qRp+Dr4ebWQB3GKYvbLX38VEhVlJVl9
XyaC4Zjbj1WSM5+/J8aG+xnJmp0DUBhytTfV6cj3uRMFVkC7YEMoLyJcqrSYJ1UM
+KHBJETk+a7e/IuIOEMcgX177g2lBJ9H17XO6bmaRvRlSRiyV6YYM6JLPPqyEZg0
jYW24a7k3kvUhd+1IkhunioR2C6JdfAcIFO5APVCfUBbM7Ny6K05trphg7KxTv8F
pfviBiJxCGykQkm8hPxDNEcQ0z8TCb0/9+wOd/nNljWXwwfFNyNVBgPUMymgWP/a
+Gsx+b/CWxgWLjFa9l2SrApglLDPOVJjTuwXIGOWz9lgMGdxqTYQs6Oe79gI0+QF
ZAztkcYzinPVZAurkPFEwP/lC4or5XR1lMZvcozjsuagvaeBJm6eqIBqBND52R5s
rv1nYTqKzu9HWzqmNyn7SOvujKBmL2JJgWj2xAoBOGeCkU3dVG8USDU7zTJwD1zr
GOwdf5wTZDy47vOY1GWCC5heT6kD1tO/OPqvIoBCeBsHMfqVrnaLJKH3N/bIlgYw
oyRxsQvMcTwZF7YcFG4+lD2xJ6fIczuwOP1zsnLW/rnU7wGGR0+L2ZVcJ4owBz8u
fKWsZJIfR6JBTyhLWKriyrjd+/oa2nzDAw+SaFrvkZY=
`protect END_PROTECTED
