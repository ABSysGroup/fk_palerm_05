`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p84DmJbO9ttuuDihzzCXpGj8aNKXDRPvkjkkT8T8FxWpJ/BMwgev5AoqKE9pyGDU
DMmfoH0vGdgkiwAGJneJhpzNiWkyYTxAp/rMzgtvNElNysp6ytBSmkiyN6rcww6K
NRxl9Nfb5PIrksOAyOqwMSsVfq6V5kVeDGHwR3cgWKJfFpHOGSq11Fb17w76x9Qk
ArbO/k89H8A3QwJJlHyQrMwyy/3zX9pxXAMvCf/LnkMwgPSpmNUyTy2fBSRGqa5M
HrdMwwFfAVvGsjNNyDWz6j/eYatd08vxbKIZ6TKcHmT0dTrhI1o97ZqdteIN57XL
loh9YC99ch2nChC6r8chFXNEqvKi9+zAiSfrJR5DEu5d211eErNiXBjzION2hXhh
7yxe6JTZZvzni75PMT6GsMabBT8Z99M3SbdQgYmXn+IsRZqF3zoYCnQEZBhz6u2/
Mbn4HqQMee9Na104Jlfx9JQblwjOq/+uSgV1513D3xhta2mBMm8ZB3adfTfYV3EF
fi8aUf4TFeMA/VW58k6RN7DmaDNqRULDcuuQoM76fKsgzrNHxXhXNCFhDDv0ko9W
K9fzKXTMcaqA9NbIvA4hZc1+P2L01b9YmpWfUe/5I6P3mAqAdBlBbrjS00/sqVRo
BxODymLJ9nnzqeJ+pGxXaVCgnkzX94SzNbwU1QxqVxTlo1VOJeLpkM37LP7lV5RG
6c3RpD+jhOW1Lb+W09gA6FKQSDcxo8wTC1uiazrmILzJPdgHd4a6rucL2wQTFu3g
c17sPNgzvB+lf7/2jAW1MyYQ0Uz+J2o6ggJ9vChVFLVD6xwJ3QMVBgQUquNFFwdY
xKJDBwugGZDGYspv/cvl7DrZhlCdsgXII4OPnCJYyGi5lbo0sOTpUM+lj7kVkF3K
b9/kaT5ZoSdeUnFt3nBhsKyNazMcCer6rKfck4zO0v0q44w1Z7ojsDT0GslLvYtJ
zwLjIhzqBgvg2uArQU1BlfPgoM6P0zUGcJ5zuxyLdnlgKbdb3uaNfRLW70UXpCbh
t9xQjg2Cv6urUqKsKI6y7kqND8sJmSDNG4pds3yLChuwtZOTysducqn08IJRkGKr
TyU1c6HohxsgxQqXUeJa3uFpq0YvM7u8f6/OFymu0R/7QwW6P4rBzvXIeMRjMS92
CK6u0kPfzB8BDT9MSEXem+VOWQEh+ZzOrWMYM88UUT0CWi+lxE6pAh7Dq/wecHMi
5iJ9MQy3WPoAQy2FW/AvqXle4hTH/oyVnBnAqtcCn9f9d6T0LBOKs3YMzYwLl75o
9e04A1tSq4v+MiqLEe+PhZ2NxeyeNK7uc79AUfRqa5nF6LitXKGcUV7zCQYTUQ8z
6v1ihEw6iGftFefrvWLoXa/iKA7leznG+rKCtKEXpHAAeKVbcpvlY5VtRxvRL4EC
9Naf0f6TWhm1pKWKLnkUpgfK30r3pD9yntSaMTrRT8hu7gdTJYbMkzcHnKtRrTor
57GnaG9v8J6irqKcyr1PPG/luDW9Qha7aaTo5Og9JZCOMKuoyHvSA5cBalhyZxBe
VEil/u6+MqZJSGjkyML1oJL+37J0OXmDDzlo2mR/01YcYRhOxFtNNKj+laUWBomq
1CAV8b7ajV+mLGfCnX73xDl1aW9FVqnbSBY+6rqELA36M6U4v8f4xWyWUzONoB+b
BR+jp0sOgaWL8DAVUrFf1G8sfYHQwAKzOA7LF/IU8nR9R5jz57MdWuf5mhDew5Pg
8+8JrFlTSmw31nQdRHLOEbxifbns6NL5G2jdtrMsoXqom9riOiEhHmnXJ2MumjDX
alpXImKN2ma8Ts+If0fXCwlkPkp8XWB9Tt9J9dyjycyFdpTBAZ6E8PNE/FXiTPsu
3ySSYjlIjfNTMOmFoDSjooeEmFpSm4i9aAWeFLu5C8uPKtCdVGNrr0ATDLpDkqIf
75fNVY0KZJZuiVdoaDjFWuXXDtlyARaKuNa/CnSVEyRaztFW0uz1EXSG8+Zmp0We
BTELt3FQh2F/rj+zXXKDUO8SFUAZGl6ptDfO/ZK2hTIDGkmosaaAGBXWgSEgwhoy
QJF1hHvTSpSqcHzLBvh8aQJdumeeCptMYaLPWQCb/zdQLMr2J3QNHKpElSDKseVt
xltX5VK0xbd26t9tUKcsTxqwib4//syMn/1/n5bGLKSsXJDbRp3YNvsLUi8f32yp
neMNVwCrXzxy5DLkOrPTKT3Kulen70ZyKbfLKOkNpxjdp50PlLcpSUsj6HH5ylv+
k3l+XY0oIneQz4BE5nTNFkk999jDrKxjeDsNPVTvSby4T+lMnLCktQrn7q9sEYw0
X0OnGJgPreXBYlv7sV/6ynjIYLQWE3FX5RqTfgPedqtluOxHFPhuBpw3zDa5fngV
t2O6MsutDYAbT+OsGX0NmdA/MzTeThZ/hJVjZ5Ny2L35H5QVxGuVrETBAyBL2+jC
zzTNu7QozA05vn70udeoqBKBftMFMoXVDFRJeFwu2aB+g8VMGKeNV35GV1Oara02
f3ZxeY+Q9nm2nrP5UEcx/nNnlGVGPxDNXqHYe2UJjw30FYDFNgEhZwmzUo4cS/IX
QCOhBao55ki7uN1b/aNr307giF6sxvfSu1NgFJLbDfdOmpKXpXEvcNXOyiq/JcYb
nauXZfUOpOxFc4SjDIe5hUSjglhaRuhelV210vta6Dq3Il0HlqikjELYDJKwbxnU
oX8/RcjwvaSMdB9byKmB4HdERWgZgwPfv4rXWg0CA6gMax/WoGuhUPSBfTMSnODE
+aFqR10YMSp6JE27nDc/iq6TyVamlOeNTxEK2nJXpoc/4USiu3jo1FEjSKwP8hpi
zq1JRZHWCjiovJNTvVZjnoTjwbNEAof4ki1yadocWoV8Fg69tV1OCUBbDU6oJRXK
gN3MEPpdLje7gcViSzvRkYke5h1NxbWj9BkoVFDX0DYoBlydV83TF9tryDkDSZ/P
xJ1xYp92Rod0G287nJIHquK9IpERCaTfvW2/WYlgapHq3QmnfXKtNSAXuHpLHcTX
NreuovFLRhDlP47xOGT+/hj2tllE2Nm9AEhlFFyWEn06H+AKErQE6wdE77IGyEFG
A2DlTL0ZQhS+xxg7P6NudpB7iKWbw878KTCrOFLWpNLSf27kWBgsRMPqgDfRy5eq
CqTgv+8r4d90iH0AYVwhSFRNyXIoBweBFwCqIYJJGyFq2vRh2dtWF5IGIBbXv3Nb
1boq86m3bGQ9zvrd9++SxlI4JRULj097lSWK6mb0yjlXxJCltHX1t0kns0M9Oth/
2erlKGEH5T6/T44FBN8kuRN/Exsp4XbDL6XEnzIZ7OEb2UIk5FbVNnfUS5hJfkcG
hpzl5AU58rMnd2fzv+NxLfj/lnby5rpPTBJr7C6LCSdoyKm4aSpR+plD57+Lc13l
K7rgSpjFPi56LyskNVZ8nuR5RutVXCGE0xSlcVOlwLOt6HGGxZLmrhgQUR+0CJNS
JhDq0iHX16OjMNEqWQacw6s5rOaCYCX5k9y0XrcLS+rubvbPLj6vsdvfv8h1is0E
7/Ux0ucpg7l+Uc/3GiDPiUy+NbcCYKJxoFbBpNUHDEhLou3rLU8JHyEdvBw6idYC
KD7E1E6PhYtYFIQeZOdcg4cs/KteHPzi2r2iSVTdXWTeGMgfF6uRzsBViQ4uvZm1
Gs9TReEfKOT6fQ7k4bSyfClHWNjAjQesiCSiSXo0cOWPoN1xHXrOcdObw1k8m7ot
O7NTTwC6QoJ8gF8c9khvrKH/2EY3liJ0lds8KGJTw8uvj0ZqyZCNUjfDZ5kks86+
3xUZqMP/8tBxCkl3WTg1q/cUuQ0HQomsooZUzZmDc5RIfDRu31PpXkhkoxQ5FE+C
lY2z1RbSJlsE/TaHbt8s3UrChusOKEj6YwT8C2+Hek0O/edVlkCR3NEKBNywIAYQ
ISxz9qjB8gAuQ9YtGUEAdbaQSirOX5xIBCdLOBaGTJav+W2SlgFwS0NRYXyGKvVd
RvxFK12hjX4SW6fIlXCZMrfILvZCalG8ObUuUeqDHa1XN58bSMq9AkNPQtg2zTrT
Ysce/Csigjo25hFr5oK6FqfakT19qIBuetxeKhsKypsf9WtoVfuYVp2YO7Atf11D
1Xw8nXXaEQNx8M/+NC1fCATQsOaok8AutN/4eRGz+3Ms0XNo2OcdC2CmNF60Bcxq
3KYJuGx0cwsbe5OSY/xU/awwBF60Dnp8fyQM+XLS2DL/GhTggCr/34adeci6xI7r
Z/qclCNxfexjoM1EeTXv5Dq803JClHbC1oiK03XcYfk8HmmLrA3KcjoaWR7KN4IM
xXDnrXNHTfJwUYUMeZ2eA0sq1H43hUb0A+TkbgWuVFIxTnl9RojA66nsDKwhc2FA
8InOdP2X16IR1H9FEq1KiTR0x6+OcZdtsZwSirKgqVa+PRgNHqv1buhGCf8MzC8t
dDCM2T2CGavmOrg4Fg+gqFytntCdjTcEhfNTbPwg7t6d0RSsQnfqS/vyH7L3s6eG
T3y+D7wvQFoPDp3XdKhPVVGy0tZgTHjZkVNaCRFvN7JJBReTnyX1ZiAmdO/olY85
/zIk6Elm3Ab0rihEhB9aTPrs/MxEk/qUBNZZdr8YUlJ/h0wGh5nWPE98wyNJURGV
npjyC/M+/1CKlKbu91INpC6wiYtKh6FVyeHitdNAdzdBv5iEi70ER3QJAAb5Ed+6
AjQ7Qzk7FJEw8u86rOIDk+pR1u/5VVZIDCeedrSFfu0zrE8o026Innf+BOPicAtR
+7Z+VElsGO2g8GWJlOkvv3HEBYgVG+DGH9MwcEL2FkIAmvZlta1dpGSDEzGBwGfc
xzI/RMHa+3UJoEbobBsbIwVgD0lWzw5O4Qec9DHGuWrxjHmmp4tukFiieHbyUIaI
nj5Gyl9huEwVA9IYV7jf/D/1vHRq6vpAIKgBd5nJGM1W/mob0o/b2rbC9WQlFOy2
rSm0RpnKzXOjUIDR4YGeq5CipZ9o5gZo5WN3l7RNNLm61AHbxyWL2Tg/DOTfLFUQ
fQRvVd4w3GnkqBSfz21RuhGzXmAIoyi8rnki8ObhEqJvW3tGWu/79iqURpS1WDHb
AHp/Il+wQRTKoTuCntnD9Suq9+lQTJl8V5FxNoiW2/IGyrbBhN1S3+u1T3zIcdRf
+h7pZNsJglistsiKqujd86lBOqVgDx56B++okv9jgjZAaA1PDrZOW5BLBQdPj8tX
bjwKofz0oPH711oGUDN9dE9iitH5+q+owgAVwySOMMlrDCfkYExE0gO6kKJyhZGW
lihvws9NO9BKHyJ/i4F19339xx92es8Os2YszWEziE+Obeuwda6WvPMNubTTfwvr
UXxLTGlOLe2r2ulvF/q0XZl/aQyt262v98m9gkFdg6ung3a6iG262QAhEKLpj+G2
`protect END_PROTECTED
