`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H/UvOPLHCUONzlgPECj/dOyIWW6U0E/SJ+CrLs47/1O3cGoSUaM+n0TsKcjIAD+R
aHvVplTWtXw9BuiRDjXljyj3/QDbdnM+6o69bH9s8pnanvvmd8PX4nWhMTmxe82E
MDvRUF6I0qT6FJ3WyBwv8fyBFLCgWvaLZ8NaFEwvDovL6b7WbYqI7fzQMtGkCldQ
wc0sdikknFmyxCYr8yX4FYbKaK9FEdBvpfqj487INPi8Pk/ZWM6DooIdkWz+BpHZ
s13B7mM32o8+bwpRZFjN7VhRUgOB5d+35VyyY5W/+Pf7b0ZrPaX8p0LXAcTBB5fT
bCSaYDDsuElwq8TBdn6myQ==
`protect END_PROTECTED
