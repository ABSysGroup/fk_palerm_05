`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UE04VFcEeoEX1J8PEO1fkOFoodxXbxxji7ubOpQaKys2nd+6ZA8PEDpXryY/OFZV
l8eiOZTeXI11v++Cb/OVi3UpGIFl3A1THq46V18P0QK25GelCE4j7jvcq3ISnJVb
bOFDVvVki5jfWwK9pDZsaxXgUKMuXwty2xZciXfy8fd8oxCdUXPTlXt4c1AjGZci
0uF19nx+uAuFiAR7TzwMZynXNc6Ju+HDkgdXnIfMwdytr1MjLksRcC4DgFbIhwJT
hemMwqijtH2dgujjSBJcnXO9PTdaZuxPTR7JNG9i4m1R+/+pxnANqdOGlIqR4v2U
wmr3HQTSo3rGgQf/Qr4XNQ==
`protect END_PROTECTED
