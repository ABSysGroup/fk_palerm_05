`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TU9S57MMVFvBNUaVdD3xsHrajObCaUVNIBeyFWPhiRvFDAmPNTaW3XSvTXKxsUfZ
IA/PmYqlYs6f+alyrl2jCDR+O/d7dUY99r02uXfUvuPlQmxWJnbawNIwLB3WW8Ew
84FI0st+lcT810I+0MPqi9lnCXQU8hqmJFD9my9YnejRTaWi7W02SmhHNzcLZT4/
VxjgeqVAi5HqKNp6lWNmIoV7Wf3kfbxKMcpnU4duT7joTFmDS36yFK86sIgmdja+
m0OagiXh5gAIHimNod3fSvozBK3nVAo7DVPjs8CiQi7K8qV0t4lsToJ6oc6vKkYP
zgJ2T9eiczZ1fIvyhkrhX0y3wTp7FQnvyMjXV1mo7zpQmiKkG8E6QYJpAvadRAvJ
qqPJfG/iTDpVo5ZrVrtGyTC/OKbIvj5hsGisV5xGTTtMf/L9neFQpUt2XGx4XfBJ
rKZbERBktdon0nnYWbo38XMzbfBYN3GugSs0H7LLKTPwYRGyn4mJLnFc8kwu6C5C
1Lg46OWcZlvlwPK52S3yoIQCjVCt/AokD/r/axP3e/Fb/Op/BgK9666/KLdkTiir
`protect END_PROTECTED
