`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fKq7ZiPrwXUJXcCq6cLPV5XNNfRueI+4ReKRj2EU4bHN83YA9ycmUjxRo5/lw1w3
ozj6oN0jPTV2oegi0oczRELdeJJfumt1VzhhXNT/URs4AZ+IO7ceFP57ltg9U7Op
SxTLyFhm+P+IQXm/6YdGqtbu4Al/ZSRqB5sMVZZzLCr+g9cynGnx05eDU8uRDukj
sAmvhUX8H7mzKl0xRTXAshcOcDyIJHjd90YShLunyWSTv8jVEyXiW4OmDG7oP87h
iy0f8HlEWjzEK4lwVyMzEQ==
`protect END_PROTECTED
