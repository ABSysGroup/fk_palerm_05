`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z1dSCZ6ro3GI1afZrlh09z49KQr4tQ9qiTkD+AtLTePswx4ta7PAC6aqT9sFapnm
Z2jPXhwA4w5wG5wdSSe6VAEpztDs7bRYKt8edPPXAWFT0Q7Ci7/Gr2i1rBz4i6Pf
as+be8xQvF4zCbGfBlYP3uCYEIEd3iAfcZKo7xFe3xCL2Az7F62sL0O7LGW59JmV
XAy/QfIkGQ8LeUryP6S49qZbAVRvt9XNP7hWXtU3IcytGM3rkvT9WVDQoXkVewWL
4y0ar+dK1egE3dLxZhlZLvWSPVjrDZCNV+o/0+gcwt6XdCOqdYAFwAEUf54jR/FB
DNgpdGoXjR+LDwF0xD5Ot0CkRJ1xgq0+/LI/bX5HfhF/PoQoVrCUhGr5qdwhCbEY
rrLqcXo0wxsg1dtHMnXAIeli41pc/5AN+Au7CIZC4iZ3RbQfV9kLyUj9+YQBFzNW
ua3Vj0OYACbpJIPUEEv9CQJOQePxldNk/rRJReMMXoVmeErJ3tYq7Eg0Ofr3QxZT
JjCEZyBH6XOvP+s5SPpmlJNdbd+ZK/0LK2VZMtuk5h1RZ6cmwU/RjniKLmte7wfW
bf0VI20QxNn3+P4/ba+62URjK9QzEMCxcftvwp/ExvGKyL25CGHAOOART6OvRSzb
dYn0Zizn0fIhbFqksw1cgWqS8RN2SJflMXXbUy9ieoMRRdXmI6LkrR60EuaU24X8
bs3z7oMXwsaYMe2aZGNfBAYZuVe+d4jggLmmcrL2Qtyf5RX025TfapT3C5royq/G
Aqs9VEv63hHK7wUp0O6SYw==
`protect END_PROTECTED
