`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zeVTfQAp5IDl++Wgbe97u+OAXqlWVYwYiLdsmQkcTUw0gK4XVtBojO8RBpeNODI5
7rsOCCsJJE+GdwJPHsD/L5Z8bzCPCV/MjV/R+P8ZvBRDeFcZ7NWI7HkV+i76qHIW
OIVqDTzXAI1o5/zXv52z+z1pcamS+D61+vj7BnEkYI/omPDe5E1Zfvg0EEjZwLR5
/LdiHzeTW3Oiy9I8G9As+d+3lwNiC8TV3/wdXsODJFGqWNWUUs8dgXNA2S0hsf5O
gSEN+d6k26qYc+3WzeTo/Y08QoOdC1cq7oMGHicIwC8Kkxr9+dOBInKiA665Jfat
bJdVc/20j8AyebMxAp9J+CEgzQG87xli2KfAnqU9WMUJ4aaj3knEphiAn23nMwtG
i6oKd+9/i4y6/synryMdVbMBXEnwMY27tcq2WhN3Ztt5vhgdT3Du/MJkqRyBhkAC
JFfwx2zCBgjhPhjHnIyDe1s+dTbb6FS5+nUyE1T8s/fk5J9nsKmS51WfCLKQcvX/
l17z4b6gqiijIVlI8+dPyRCjrDN4Qsd+rjHizU2KuaoyfwCpAhP3cPpQO+Ddv4RT
1GeJZuNwiB/HEahrLL+FLIWoe9YhB6/KKi0H2Vz2iaS4EOk2dwLM9n+9rtiUwwpM
jOPN4+0Czv8xr6vRmMBfd+KxLR8xcglVJTXnw/C97lF8D698CfHl2bRZF4nC7y2G
5xsWnM1zyroRR5TW679bE0IRGBjJr8iXWLm6iqb3aMGcEDG7Guo7L8xqlWpN1okG
W6tg8QZnP0ZEQY/ogNCNDbfUMyZ73d1OU5EsOLFIEkeShQFjDOcNOVZ1/tzT7gmi
MScM79LgOLiIYAqSCCOnV+Dlbkh8y/UH2WubWbxB/vjPeB4GY3+vI4Hs3WILGWE8
CgkPuAkd0Cy59DCU0U4uHtvgMWzorRqe4PXu/TWiXf+8sWweR1WHHPe16Z7W9uNf
`protect END_PROTECTED
