`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fcdRub1NyDUUJ0sjT6dwSaItK6IKM626pkfcpBAfeRiaYN+sVOqmDEG9H57eWkT8
j+fS6LotLtlMY++rVQ1Oq9U/N+O4BhuaLtw9nAU5Z/Um018ZHhFQOpdu1tZnT09y
u7o5uyXsuETPubV+A1U5ZTa6vAg1d9ki8ARIaDtzvVio0+V5RwW87ndBHGcWr4KE
KAIr1zICfmylD98KIhVPTq7i2EzjYrNfoMkaMSZDV0oxqDl14KRVm7ysfNBMY+5G
Be2o15rSghBXTpIRFx7Pvcjxg7t+PnKaQY0icuNDe78DT7KckcO7/YRnpaNPde3u
X3mq87ofD3a3irlyWaNpQ9hCgKBmNJgdEtejIyLtMw0k4SgGNDxdcrkDWe9v8zCj
vB/lI/MscU4Y6LT/RHC5Pl5I0ziHhzdyjZ36IqRFocHjRhqrdSmlPruz47BqMjC9
/9ij9g/XBfHRdM1LQ7RG3ItjnYCQBgqFR673CovHuzCKJ4eXmvhJs5sJQ35tmtIl
KMQDM4jbiVU504xyszXkJEaXaZ+OyZyfwAxUeKrZxenJzbjJ6E4XFOJm6xLo2y5j
pxFkRW16h+wCBj5V0Q4ObITsRc2z7xaXU85wheqvratHjCZ8I98fkFQSwQ8Rc01X
gKW9Z1V6m+zka3hrQZ914I/xJFU5lduAln2kmdFOG4tiADtFuWzy9GxV6fwsTAR6
nFJ0Zgioli+Ueqb6dCZ95O7Ophkosqqomdup0icrpwhyUZKiirTiDLu+ZtDWUUqq
6Uex/wND4g1oY+2qQAYX3Fowkp+PLIRGAiKtTWEIbiks5exdeQUVYEZsLCS6RbPP
bLrC1yEph3rdBBumq/8++fyt3KA89d97Ru/Svc7BLODsGWc8apJG7Fnqy/ghwObO
AUujMS62HA6+Mud+7qINi8bGkHUlUAUJrjzkb2QPScuFTCBG4crI9xykCxh0izeT
`protect END_PROTECTED
