`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dXp+ENbYexHS8t22vFb0MllQBNzuzOFKmxSeW+GRFO62t4bFtqYh2N5nJ6v/jFFv
VHJwisTCfJrij9oTCQmrDiu9spbhcBe9wT1P8LwjF0fd07y7nZswGOcIElOmCiZF
qSRlhoReVwdlhrIjj+TiS030o9CrAsjmbRpsANNafBXsIFXI+SETVZ7vz0ioZTns
YI7+xQc/m6aUGosGxW/OuWQ95TpUB0qNL2ZC/sNurL9xf9c3HovusNR+SCI4nXQb
PS9NI67fWggLTKOB0kBt5XkhdMAI7nN/qUthyY9y8AuoOwoGT9eTDYHy+MuKqEir
Mqly1V3jd1NdX0sR+83H4uO61nJJBoxUB/pr93f557I+/WCKcogM4W2rPM0Cv6DO
1+Nhmcbbom2OHnDeZfYciL5qxy4C7hkCJQpeUYpZTrUPK6kcS05gb90ERQRKAbcX
YobgB2fvy879wNK8pf2FJjGRd1K3JzAQ6//+KIz6a1s+neXf8eRW6NMYjC8O/t3O
FfZgJ8kLSLWTsw0k5e0qsX0KJRnIP3UoY5ohrqG4b2c5ugC3SRb+B7o9UYi3nEfb
G+kIi1vWJGlE4YxcSHWFlVZ1XzSAf+5Jeixi2C5ejXRwPbY9c7l+AEsez0tpI3XD
qYSgJOfBsEJO8j7jQt2+i8plGksyE+oL8CC0ft+Au+RiqiiKUwm7JH86l3fWUiMt
tSuEBjPaIcPhdc1t6x2ybcuYEGJefKMVv+oHLPvQfnB1uliUXz6YcO6Uplx0JGnJ
bj25/RKIO3ghPuqaAnQ4gaw3ERxpMFU/mf4DuynGUDbXQQSrAIlj/v4bYYhgtTQE
YMOKO4xTfK6mScHIBqH9sUn93qd/GhTBoU/izmeXxvVQpjQl0q1y7wP0dMcE+APz
95VMUtLZaHtjHHAhZU4GibL3qjmijf7CXhOcUDNGkKyARffkFREjXIQYZ50h9PbD
hpaIbjVx9uh3Gfvb5uzO2MOrXYgFaYHKY6fRi9ZEpitZZQy+GuBO5/ajuH9D41Kr
gRAYn8CSZK9MwKTeDgmYqTbwnBWR6ybot3L513X0JxJQM3kcv1qXDSZAT6PScHWO
6UuGPagLRJ3JkW6Gw2hY4yahIUZ3d86iPhgHppF7bYkD7zh5/91cwb+D4KObUM8g
gJPOxwDy9ALvwVPH5MZklwj+DO6z0hZa78XN2Upmrj5wLUlsT0WBj31nLbqzIlWy
4oWvn1+L9NgW1kUqF1avTqt1fq9RS2HkGQFGhRS2S1s4MfPRBwJa0+OVxzvwun+p
Td9PUKNHtD6AseuiROBpm54LicvsTOne/SXFH28ruh97Wm5CQLz2wn7FOCtHaaaw
CNby459mKsOmZ6iF2NHiErmaiTjjrE7hwRFTVzrMFAEfBFIUQlYklaoobxyhoS11
YjkFDOsKRrErhTuQh0knmUhKO8lLFd1Nmt0kdOIVgEx6bF8uKaBnsY6woFIoKn7b
Z4CA/dLUpRxmdcbYCYqet7lBmc8vBxcQ6P0sme6Gx4+Sqn6WXzSEa4f17E+GhGMO
IwGOlnnq2j9Xgmz5iD89qtVMLHh8uxurC/5YqzTJD/9k0SS8ntTF0GiDWE1Url+f
Moa8bCIwRWbAnllaEwIXreACs95V0VHWOBhTQaJUNrvO6uOH8bj0+66LFdOf0A9x
XtImx6xBUYanuHdtMYo5PLwrDCQFa8IUj6a1isCiEaIb0Zr9VPCVxDGHmhGgG7Q5
2MpCYhItqc84PzLiibdhwoWuKtbtQMIzupEM0d9hNJwpyd75WVDci+jZQn9h39N2
swDqSoa6BmAuloe3Pi8fjSwkll4urFJFUOB2Y/O1XojydI1LaMxPfZcuFbGC2ieU
z6+DyxHuPSL2jah4p/3SZ+ItVilqC1UeaLlJVl1Ilk6S86WzufMHSefHxXgh1J+6
WtQV3+Xtogqrp4ZKH4ZQviRHhJpDc7yfxS4QbKW6AGPy5DYTGxioBWwWQigbHyU4
1lWvjTaLm2lhrdxQ+fkhIz6g1tsY/zlzEM9G3L9bMvtdAFZIsitUbM2l/VhBT5n7
trMG0z8VVhyo/GwNGr3kjaKx/J2hjjgaxpgPDnEEup7T1KF13+ou9Ur686OBtoV5
MqxCLgXpqecddlIfMqD/KdyuUDRGiK7IXCpdBZFcDJRbwUQhMAvB8ghoFYyElrVr
TRE1E2xqD3BWPew1RYN6O3RA56W9dXzubdKYr57hZ6XrqSwuIuzjI5HucO54kyGm
7M7oHPk33k8Vn2XpW+HP5mdBbu38oAhKf+IrfX7OzmRSDxAwODukso9RS4hn6vtL
Dvn6RYgjNCuSfG0Yjf5QYtWi/dF14tw0yYy3t/5AbzRbRyeEx7BA79rZFZ81C9z0
YqjBzcMNG91DKmDXeOObU/kbH1shHJs9t4VIUiEa+Xtf7J/sYxFuMnaUbly6bdM5
gShYTll90UarxN6HQ3PHlb6D+Hxzv5lxdxysdJquy6fecNnFdlNFGvxNIYO2lqcI
oVG3VfDcl4vxkeGbk86WiZtV3DFWxdMLaCq5m3YAPXNhRauKXuhKcGM6H8Fzlz8O
ahaqsam7zYfJ6ckAYo1ZxCpVjfbL8cxW/24CFR4ybddV5rjGrLd8mulz53mugxil
df8Qz1bBZoTu1VNlzURi+BNc99cshyoRf+CnbW8TTkpUscY8HTi4DCd0egdApX2z
KyEfu/Bn22qosY9zIGiNECdH9KSRLp2NiS6FHMzjtphgf2L5EzaKeT5Q7M3Rz8Th
8TXMMs8VkmSyX7+fh/A2A0WlDgdjSix3DAyfY01ChuxqLjFKUjutU2p8gzT4yZdg
AxXgY5xxvjbGXxMHI9NAnCxDAHT7/QkAGynzTVT7Lw4L/y92Z4KfhjUuiiMUcN9/
`protect END_PROTECTED
