`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hzgbZeg47VJhBIliNdbxGIICynjWmyvD4GRae+EtkwDq1L39XPCCRLWZQhVPnZZD
JDVjCDw/kS53KvW/fU2vF3qB7pSP4sATCir7XyFz1VA5KOnDZNPvR+iN+NsOIFJs
KD+qeV4d7foNrz29OOQb+I7bp1LhVvTfJIpre2tqZx+Tc3ThqAFrup/TYJiRBHgb
Twi6jqNkN3qlO+MhOCDHWO+9CgsAAbN3fC7NPRLyfZM7Cp6S7ZZXF8OQRLodfVUE
7+2rUgRShRGDYpRu+rqV7War1bawU03ksfWIYzcWMKZolV36b75EB0DH+KcyRctd
1N5pVc1L9V6z/4C3fzBfJbt5UQYep1zZfpEW3ixfdxeiBo1kw6l8Jpp8MOm4faHU
NrSNGfhaZSG2bRGHd52KfYSUQeD51bajC1MHWzV+PKAXw9nLy2vBfrsvBhuc0AZb
zxOG2MTG9wp6DMXK9kxxR9poCZyO1rv5G7LozLPZlydK51Kf5I2R5GbI7MaVWc59
YSQxDSTSkOnGVjXav9F/WDykaNY/qPNCzAPkeRxQpCovLN0XiulBW2pjDlbGx0yR
MraWY1pjJM45EFNgmeJyuJ1ewpuGuT7YK8SDoKdtgf2rqUg7huhX8J7c9/+m9g+t
/7rL9vOZlY1Lcc7wjoVeUxK40Q+3yOtcmmzsp8yblpQyQIG3aQtBO8LoeXD4/wIF
3KssFVuTeaUl9qFXW54Vo0gz2hnq62lcDAhK+7XvnrMuzrmr84EbDV28Ur9w5DRb
EuzqUTZOU9yiW9pTiIXtTm1hIHNTRgXe7PkUTPAmZSZEaDkjfU+O0AH1L3/wZ+h1
JrtZGlzIwP1+lyDtXtyrIKg8/gabuDp5cjxvXfhmEmQME5pJrx6+fNgHbjgCS1XJ
swVyzWPAy+vJPpEwDli4EyOq+W2OpsIvC6skJfYHHMeyRmyYnhR2TIrsnPKisCiX
S7ovjFi3NMWvW55GFqSKmStlpRqBK6juD51iL5WVBcEkG/g+aqwFzIXOao+yA7Uh
mh5mdXz6IMe7GbAoTcI8Z+UBONcz3ZTntY8F+Q7HoZ84e3iaMmFyh8vepQ3GirIM
7NSSzq1gw0eaOGOlzyHhLnpb748ENojVRCfg9AWmFu/ENHJP5FFvgsoRI1TQwD7m
veOGmV+TxfQeHEIDMKVXWfJkpm2ZYTzdByQBHjktkVOyZTmrjjc+UESBabwVx/8j
Rt9wRqZsB8m9sCh5yMp6RieMpFq70FTEP0luK9O3qpHiCZwtV43ln/54AKMPOi3l
xGF8LElyq8XwzSIu7NcoPFuwtLFjNV8N378wrigZq48Qan9gCQXXkrvJJh+1M7CK
wk9fe0uh/LIDz7qCnzyZReTxAr8qxOakXKch4nTEwaYzXADt3IAMyWaDj8KYH0xQ
RDfH3QlAANEZIZHdiY4FAci00aJLCTgUuf+RbQO4fdr4/1voPBIC3e6+7IThyhSE
LVXSEA7T2ks0dbXYJXFJDatSdmYocEX4J8BJvU0VbczmA0QHwYdsAgCtAB40aFi6
fotKdv4zGujTMminWbE22OJaj8yQkQaEH2rtvpR1PRDZZXl+IgHIPwTtKB/xZPku
2vRSwBfsg0KEgcsGiIYbX5Pwy59k3VVRMgyAJ3v69iGJiBZl1NlogdrvVcj1ffAa
qbjqJux7Kkx/mLPEvn20HaDK0g4AX2m7EDh4+XgI4oCi8iNlughY9IkcOorlpBBX
XsmtUS8aoKPoSJh3v0noYFYlSuV7NCz0yUsDoORo9MP6xxz9LM9Zb2nGPg5nFltn
DGyHYvW6UM4ViTlqj6OsMhET7+BF/ZXoCGJqUUwSvRh1ACkpGZd/75qitSa0BCBo
zkey+P9MJPAB3+VjHDl8sJ7QwGT0HbVv4o7/HVyx2iY0SLjWrpd7C5six8uSVNbS
cKudPLCdoUGrTrkJg+HgymnV0vYgT8jLHs/BJhQ5LYP5XBtcPAbqeZAFViSsJXRd
TlTYncmMA/TCbi4e8bZrIYmuuGd0w+V97up38Cfe1/i86QA62uD0QCQovMfXXr+n
QRn8v8jO5+UL/P7682dLtUCFaHWKAvtw9FvfllGCUiV1F+N4KrEy3x992naTKAAO
`protect END_PROTECTED
