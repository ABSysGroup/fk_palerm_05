`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uRps8MW0bNif+DOZ/jAWciyMavX3t90uDH5eTNwWuHHDS8/ogHZAIOXU35uR0xoR
wA00CFDIwgQLLRQZsXrkoEFa1sYiF+A6Meyp+aoxiO+F74JVIqfV4SGNPmwdVvHF
EXgsWxqiRhefIMLdjYQ03ZDf3sZCgFC8D0es8GO81hulV3j/cBumuiwe/B1VboKB
G0Ht6A7GPpakAFLbziooereLYETuviHWx6Nf5+PKZV7bxvubTf8dD4yDrtP6ZF6W
ZOLWDh3XeYYN5p7v+nlEtgob3Npe2dDjIJ71F4/SJFu4mdrf+DBY+CX6GhUGdMHs
HkATuXYzplDSdK91T7aUXeh4N2kl7uZEAb3yucRuj+zTG5qu9RROwII2YiLV2uAF
LFiVc9M1UHHmJK1gDjXiPDUsWa5ulN+HONMo6TjkvawoLqSB8JBuxEWRszTR5DQQ
oWgdxe++Q2cMfMhdrEwHVZq8AcIabxEKPLSXyUJyDyF0cjqRjCJSq8ywKhvfmU/i
`protect END_PROTECTED
