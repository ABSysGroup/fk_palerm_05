`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
76BoygipJUokg9skTC/NBC0Kn29WMQHSzM5GEy8N74hQUYFAk9QksklDEd3KQ0LG
DlSZer4mB9rNiy2Or3LOeNgDG7dOS7AdL9iCuBMobdf6X6V/ET+inqk3LE6ZKwN+
OoMvU+Nb6FHF7/HpRelPvVKfObgaFr7Y4CbKKsGuAaWlyzeVh+Rldf55lrzjcXMV
64qSiFcwWG9Lx+7AUkC1M6kbKryzodYav3hysxOstGX0SH424vSe5I1AaacDEgBr
x+GNlq9vhW6bx6LGXzex2M7XTAamWPBPBBN/NNIeYQpcUceBF0oGK/NwK9+xEtOj
JkGfiY3WgW3i7Lqx8qFyMIUkwtAU2mbJmgadUVaz/aHX4/KGiWtPhdVU5Pt/eole
CkiDQofij4kT5o/jZcBH5pFqg9JzXbjswzsACeaOr1t5SJ/N39aZ8T13UK0AQkEU
RX0tgg4y5dEihxYTL5TvZq7a/nVUq8tNaeAKiWMnLvwAOHg+GDrnqIoMBwNdAmKN
hTZxlHoRMsB5AHOTYoB4JH8uN/yNyoPBFW3HDjBk9T7/UeYClit7jmIhbartv0Ob
`protect END_PROTECTED
