`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6daC2mijOX8axhNmZiYyvgRBQbBPsC6CQsMB7sfoB9l463Hj7DatakkjYBFqpmd9
JWmDaFuhTm8frP/2fBQHhk4+pKzdZgk4o8Nfky3veMc/DcQsx8A7hissOL5LT68J
FvnyPhy/lvnK/lxtXspKuO893N6MuFiNg0IuW1W0ZyRb7x21HLU+ByDhDGZwhSle
tvIX8ksJEwVeE+s3qDYAAJCw0Bcm9dh9KKmF49V6PitorvZgBOCBmKFPchwvuIMH
1Ge1hv/FvbHwxhgZFb2aIm+EvywgkVDhlV/Cl9gM1HxyNeI/Dr0/9Z+gWXHpCw4N
s+jYXYtPU77k7Q6dyfRZkA71n13V9cgi42+rekCZXzqjHFYBAoQc/S3QvluwD5RN
m0Glt3mA+W1D2UvtGhSh2sFW5+LR3+X5Bl7aD46EKe5O+At25+rl8K7miaLVkE9S
+n/7d93ZPs7vGPssTAcxE3qyrr5A/t89YP7atl2KrPj379T4IMmL1xuFzSoC9pWQ
jtK996rt/Y6xxA3IV48Q4QyiSHIMNqEfpEG19plO3POdHny3g/I17cYOuCsx96u3
kRvZ2oV4uI9n8EuureEDAvn4Nsri3VurEQ/U4tVMIBWmR/ZjSHPZ4mCgtpJj208u
Ih1eQ/hjxxIhiRLAEQI1c3KGc1ux4NVcLeLEvxJvuYqmqcK/Yc0K4o75/xL0OITf
zlv6A+xZFo3XkASheF+DU14mQG//KdVjPq02w8vCCxa0jiJnhYDFijT3d2NO5+hl
SHsp6ug8GWgEDHEWtI7ujrfQAVmsiKplTi5IQsCJ+ItcYONhYyLX8G13gT92uc0A
34897jsoO6ih1Da7ikhYsVVdSnZz9/k//lQSl9kewzCiTN5/3Uf4sLPVZnHpj2dd
nNpC6g/w0kne7f3GO6y8UvFG1wKfyQjZvAfDID7xUrtSeQ4ixAuaevTMFfIpWjvw
i6x2MtGf5fcR4NqKk+JZkcjm1ag2QNjA5oGQozzA6UH00cBRR4ir/PGPaapXWof7
rxZQxzAL87Y0L2COPBL+uEBg2YZZPNeJsiiUO/itM7knLyR9ewi3oLDLBf9xIIdj
aIoDAKvxONw3loTrCWb0xzOS7RleSoMo8sVU28JRpU1JCpG/MdU9hSgx9gUnFt1F
yIrvCSsIONIR0NHQ3+MNHTK5FP57Zt6XK5cGcSTTrZMnS3jAAlzrTKjXeAUTlGed
uQ1bOObmEhtuBWc0CnieGhh/HQtikMFsSaFlB8wnFcyHmgj6DQtxMQS/PNyAHS6q
`protect END_PROTECTED
