`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1GCplOONWHYDoQsK3jGmuMuCHrLBFAKR/RzYXD3yE7AC9aWTQkykxmKVBsxixX6j
CrBX9NZonCq0Qg5pkvQSogY1xNE7jdfTz2zbgZAYdPjdq1SFsOrSN+gLRWUVoEXw
UEde/Zqf+lrF0B2/7RGxfobB0RsbnsoZPGAGiulOxNGVleNpqaq3Qo/qVvlVVoDp
OLCJK3ScDJ8wdCD9lUtgEtj2kcTG7S+I5Ubk9qn7mI7yUHCygP/f1QQRZfncBxas
uzkRdgilC1eW+JmIdB09x6mjNMPzscddTVbBS4YozSX9YLhbTaJud01QBuxsU+lz
BTwpHpRXMLkk0MD6laGiz+MLezX8G451oaKrCHJmlFfaz6v6XdYD17h5lcsxa1cZ
UOQ8f7W9PrYmnHHGVHTG9D9F8pjElQieX9kv667Aw6syS3FL35VpfTa3NneUXE2M
Xluqu7thgkKv9JD9I0dbU1YFmO87soBTC6WXgIlzXF9Jlc6XOye+6jrFrZuit2jz
`protect END_PROTECTED
