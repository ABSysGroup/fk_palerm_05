`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b4rqEVOkFs9uoeZcV0LkIsfStAcYaee9Zefthw7gkApAxIlCEAjWYxOWNyin0TxU
x3N6p3vtSPjZh8qYv4VFSom0YOAhSUOghebEteJAGCwJ8hjlSkXE7Z1sJar915bD
hGiblAbsdC6x7woXgCG9hFZUC9daX+fSq5xiB1OpMRAASixxdyRpvcaSHRau7U6Y
Ue7dxaNP21JnEQFjx2JHc7zdG8ujMtwTQdv3+SKwMP72BY6i1qK+Vd90GFcXVX0/
pMrreaItVuQdOZ3MQiX/wJo4UGAANgd5RxEMtKcnuimtCiAknuYP5RCbeh01FgWn
O4NMC6FSbJ9Zw4G2LoS8Vw==
`protect END_PROTECTED
