`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mxvXR5vzxrXdJA0PVGgVIgRhTvOiHJvkGzNhuWFoFqydqQvE0TDvEz/7cy12XLUR
Ubo1h5PfxTKnjbuoY+bmPtdcnx0e++LMo3dDyAfXyal0GtmEP1xGzYuk7okvej5Z
1THbKqcVvMu/BoYATuEKTkRSOPRy12YMQxLEHB77HkYn9JH2frEMTDe4z/5xWwC3
GRI3BFTk5bUmwCmPeepfwdG8p6ldoEfvmo7U5FrU+mXBT4IZ0UKNalFtTNCUbBgD
Je/OPmjfgvSPydXJrrVzEggPZk/26eC/k3ujf+dRVF/Zv/Zn30izN27b1nSVCi0v
DP7ZAJuMs9ESh4KEQFYHW/UOlLysqpTJisxf38wgKs2TMEo2QORVvtX8rbH4F4ax
Og8Ho38sseRhmj9xAQwN6697LdWD9JgKoYiagu3bJUGUL95PjfcEU/iCQ+ABveDP
bkiAqvLAlJCjrXKRhI5zTw==
`protect END_PROTECTED
