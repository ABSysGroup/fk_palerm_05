`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GFimYAGQQuH8POsxpqduiahwNCSRQrcFktIlshgs/1K4BpfwIGnhZcA3j0VpbA9t
299dwag9imc51NPUNqGbr4LphVZ7i03nFk4s6rgSYOFfw8Iu88AqlQYCWdK3fY0D
NTT1lmAwZmLItN8DpfoAfVwToTd2kDGFegE3bMeRd8GbCXIR1frIlS5ug6TxsX6r
mO6PCCeiVx5Vr1bm0xnPLTIF8/5OKVeV08vhOcDuqqKvF5sJXAryuCHc/ew7+MbY
Ia5YcSaxUFbHYJrG4Q2N/sj7u3mX7dCB1FMeApr3IlcPPEuVoCHtLCNbFm6KlEP7
hw/Spg/0A4qmlCesaRIyiRDz0BhXr0veG8B0/0HkSG4qu4p6omyjTatC4qFPbIbs
tcHg112bXL1gNmKF0hTubMlUyG5Ofdp0DY6gUn85U0Y=
`protect END_PROTECTED
