`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iNu69Tlbus9Vt8WbRS4FzSzxpV84USv2sFTcKgBCnp9N6o3WjCajK76eClVCaKa6
EXlDqXfDCGXUrH2wwdH806QsMniuZDBQmkylFuAB3FPDLpJ7uGfiYzB8sb7KYJ+S
IHXIJfPUHudJ2z3KwGZucAnFAtCiSSmzyu+vFVQuixPvY4amzhoEXrGdCXG6BhDh
AAnOimETEI+M72N5RKToW7OnXVfk3T6kxEP4kB+ClTS4LbwGg+sYtSwUT+BF0n26
CqKO0Gd+74qvJE+dycgumf55uQL2SGzTRXHTg6/VX5yrE5kAoroHXBtoqa5jQGs+
0Xg5vzCio+CRrgB+9wXBLF5ytMAwohVgo5zr1BUDq4U=
`protect END_PROTECTED
