`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4PMfgECcq9y3LscccpM18jNwyB0wzb53qNgQ2/H3zU7r2tVj8mFEKomVpHFZCkoh
zYY62NwFVrJIc43fdgGX53N7cZ1en24aMag7Id5eeV7puADR/t/+AxmMHxbJkDg5
3adSr/YImc59GdB/6RMRR1vHbNkdDgYUP2yyoMC9/KB8ztwsbqEd2+AYy9eF1yOk
c1IKhmftALVg6yyZuMCs5xdo7xJPNMWBzkA7fr9FchQpScBGxdYfo9nIfBqTMS29
ZdAMJH+s2pzFFuIu6zT5NWzcU7iI7T7vPsGN9l+N8TbpEQ/Xs1NRYlWapADfbiJ+
THiTEZvL8+LzdoX4tmuovA==
`protect END_PROTECTED
