`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3t2q5YRhvVXBbM3Ek69GE6PlTMduMHSGIMRF4rTwSoxGCMYU8jm80lm/eviKBnfm
M57Y2d6ocDUjAqErrLK3Av7LgV+8RxB8yRrK8AVlgRlPeDmmK1borMSiczhS3a6o
DXgqt+cDybzwRHIobf8vjlTdEIsJak8i2VKq6bIW/VvGzPPGN23e8L10iljPDkcF
Z/KkUFHrYm/tbbYQByUhwtMfOnln+KUBaP6ElPUnKvvvnKodiPEiLc54Z3Z6aycu
9f15YBskYe4nefTBZTmUfpB3LFEUAtaCP4AK5+p1KzJDA2mXIHVl5Qu/Vt5jt4BI
56tkY/ZS3Vq6DoEbxioPyX8J4FwWEPoUxOgClZ0PpHW/4zRu57EgCOicZXjSNqKN
4AhMp29WFzJ0cqcThvBbUpYe0u1m1/XBAp1IIt/5vMvyZ1bC0ScYKgOY8ALMJFth
J4mj+4lYrDzc4tZWE/e2Yw==
`protect END_PROTECTED
