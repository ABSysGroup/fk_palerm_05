`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fv0CEBYjUng2+rUsmY96XTukO3XmF3tcGBoCryzKHVSp4Pod54+WoYmB4WfhB9kQ
4GZeRgTbMkQgdKgkVVhiXWNY27cqqgaWJw2IcyS6CS00+2bjABTWx3GuJ3FOkKTq
JmMkj5GlbvjVl9CcpXH4MCNrX/lksc/TMtsZTMJ+SvSTIyX6bvY/WINwWHEDrYSf
U+VGrHoDWNGHNXZzwFwMmBXzzTj/JHMO3/crkBSl4cs5TmcjbNDpf/aIx6vfc2Ox
NDX7NQ7EEcktakLGr4ucE4oNiiQPiJmZ4tvvYBH7eTy4hXh2J6MYthiWIHS5IA+E
ESZUs/VWmCENBvB6AJ+6FaUINGG8S3GQLT5hEfYTnSLVGhnJqCeFR9zdgLAvs1o3
GCO2tUzJPq/1KCCKmg7fGZ5Ehu8TG3/NEByXjYq7vLvh7byTSPZXlZdPLXqmVfxL
gArB+qEMwSKA0ODn+KPHqhWzDd1cTfYJ1iigyq9NN+EMm9Jq/ARUu7Bo97A1NW3b
Iw8KQRHF/Mo6XMkW45czXjm9vYKFJye/mJFg6lZ8/84hOR5UnDwrMKnVusTfyQmk
xzd80Bq7XyM//q09bQeY8n3VOz78ed8ZNLerMhWdZfkYF6tmzIwyNZD4FCfEh1/G
0IC+jOeBgi8wMAP2nCey8BTOgULAG2Y3bVV5F/p6YRPsnSueVjCewzEPAFCVfFp4
3KDpBJboZ/6u50jpP0DEsYZvp7+ddvsVNbIPlnENGYWaZDp8eFbikEOTOryX7ckG
1VOMgiLj4nTXjoimcLY79YZJE84GwhKzq9fjFceEVrOTBI5Or0/MEJInopxcRL+W
uenqSoMXcywIAYZB/4tBv3pX5Xi/xjJkpyo4HB4pZuyUYvqNES28NkWuYR1SedC5
e5WybHIqldzjJXmuLNvrr5hshnoHAO96mDuorJDfrDzh4JDww58GV4qFoi2kmI2A
IOFjFRdxENbGsKFk874nZGEqbDDs4M71jXGHrgNzbDvPYLxz1F0DWNHUTLgNLsMG
qKPzVvI9128XiSyta0k/DWssubK1QYfUJ9Vh/p8v6NnKR7xssvZoGinXpfUhGvjt
OmF9iVB2Gj49t13Yce5oj2nxTs6yLnJgDvT68o3H88poPd32E2rtTWcJkWnnAfWX
lgTJ5X81MmnCqNhc6lmhDAoCcFX9MvWWMqTEktQRb70I1yNxqLTym7kwYeVC31Yk
PaDebwBzSvHv8s4xmThPGqfNnqE+5b+Y0h7kG8MZwm6zieN/iQkWfMybjJdaiaV9
nSuBNjscSMwuRwqFq3GUSJERsVSYD25Es5Yl+3PdNGrChZ59b1on+Zl0lBkji9ov
WSLhuekTT41wMuRTrcGV8kpGWB+60JCLgLtXjywIq9mnVmRlpI6FyaGOiywH8jg4
MtMM8PGVI7Toa6HC12Wr5KhtywFH0M0lpDV9VFDSgs2jd7BLpnnt5EjY63jyMCnB
CK2Pq90Cz/dVo9l+pzEysn+S63DCvO8iukqdWCNq9O+q5KVbcQA61DcY5FrrwfE4
+oj31bqTRlOA4eBlJ5m3kjZ4Ss3foa1eledxxcTH2PAqIw2vxr08yL2gIkeAjjcz
YGaiMDo7dy9Tdg5/dwYBPcqrgnhEm58LSMNmwmPhaTlOFLm7MG1OjgPpVq5ZgWN3
Z8+abpjUVi4X4X0WntyAFEqNgjbC7b3mPomfcVuN1Y1aczXaTFb8Gg5Pftg05Wjg
o4S7bbyd2D34Kfqw4ZDDRxpliNavsoDOQpF+qtBGPmFiaAyJUHZSRPjMJ99GIIPx
L+V6e5xf6rs0MPfVVIgvgIwC1mSUX8LtK42SuMGmkuCYjTo/HahJ6DB6AXrVpQi+
gxaVJXpreNDNXmwxeeGtnxNuUxROQAOQTO24FoW13f+B6Nvk3t8ROxT9DO5K3vso
gPtiKuNKcdFo171lE5+oFZ0pLGDheoUg7Q7qahBQy51wzukrSV0PTNj5ubO1N1px
7lf10sPLu6UWE6jZ89D1DKa2SefIfpWMyKXYkO0O9RGT6mOBXDF6d8DTaYdg/EpQ
VauwJpCfKV07j5vGjzviFhW8ole84sPow9d5+0l+ad49FoADsaMCwGFGM9vih8vL
L3qqOynn18CWdTPs5wwJ/9drN84TRFOgACjpRjV2wccPIdJgKwz/Yt3Q/vhnWizm
vbRXzoYK/RXDYdohBb6bPa9J4XL45aw5wH6St84L+7XoH/n4p/5jLBBHu4zZq8xi
giSPg8bDXFHs7GEdNLKVr7AJUrbsxy1yrmrkHgK+ZnaZQD79zfrMu3c7Vygpe7aF
CYJyUPsGp4JYcilWIxhCvBY5qc/LDd33mXnFibLBeVLdPT0wRxdII/t3ykvaOpy2
YRRtJNj6Fo6fMWF40Jgb7DUzzjftkT48QTap4uKkfYUGeAVC1olXorxCsWX3IYDC
yXV58RI7XRDvcbdHmVHto48lHvUZZsz0GPuv7fz2JgF0mPlspLONxQXe+TsN2C3D
XlYf3BCoHg+Ehl6GpO1nrz96j62ciMoTaL7GwsGaLWYbNtkJg0ZJFoFfIW0fDuqP
aotJR/lRxsu+rOi4k9VfiuzlMpq0iJIJUzsvfMXQwkOaXRKImScq4VNKeAjaf8R6
9GcYmBrsDKaV8rLQjwqmDPoCEf1b+KY+oBvqgZggR4zJQe3shqzm1mHsfHxOJIzW
zuJJN08kY9ob4RQUv1Sc9WitIhQN4Rrqh0RTDycnj6lKr0AhW2XWx9APJsUE5m1A
S7/fCdy6Cg0MbwDZiJWkKWnY8aO0sTmLzXqV70ey4rSPkCfV2FVlCn82scsPI4zh
6/iB1kq/xURWPPHtAUKkcOx1WWbvDAGzTzl7R6k4yl4ZaCZAAH1snnBLOIf8a8QJ
LGLK8PGhiEnYxV2gfcc0ecQhpqqIUWFCCGcy7Kin/AndS+Oa9yfN/5f2BRKNhxqh
b3qZPuLgV3Z3Ouv5CusLlnobsUakN4vGhgltHOJgzkv3wCSWFEEFCTsroLIYziQC
CZ54YPECmZRLRJGzG6IzI50mbEWD+eTtMGf7ZaHauOOZnDLYKVO7d2qXWXmDdQYm
MyrVWzr/lcjwQOkS3Wnf5tmNnvRt7FGY7RAsxjP2hDotnmwy1FBCpFX/FLim0Sur
D7qvuNCamivciRYl9bE5wLRvH7Jk9ocCQcsO5TGw6nLeZotxvLjnhYoWLj81eKr4
ml9DqK8SzSWxJ6CWJWVKfMCUNODqyAo5pszv5u1KJmFmFYvx5y0lRO3gUfcAe3Wq
f3iX5NOCeCLF4J/OW097LQNrw6LVRPuPokk8514spykVPm1VolFYmehxuZyv1wk0
fzvOKSCa/hfhQpVQNytj96kxpYPiukO3emdU0LkFWkg+XcPEJMHUh+u5vt9tMtY8
VK3vtUpU200z4nmOrbQMQcbLIAVo12a9yNLBWKTrG+yZBurISlPOjMfBrpX/6lpg
hKKYnVZPutcQlIUebzsCiiT81dxZKk1Zqko3XR/XaZJGOx7Jdt5gGm5ICd2kd1Vy
I/UyGKhZIy4Am8VgbMfCxg4UwoxBhXaBvEv/dvxP8/3VpKtVQux1lUmxB5wkv5IZ
qjMNXSL+bi0IOHZgKH1EGl6sIa3m3N99hiuUE/CZwkOJlyn83e8fs70NWYBUPRy2
WcrUV2h0n8QwAQbDbSYPYE8muJZfFkNH7MKD+viPS/hnoTqNU7IAxOwO8oesTVaP
96fGgG3TQiQhAgIncSGCfwT9ffsKKTqc/zCsQdpWCjX/CNJWlvWjGO90/1IBlk9+
c+CxSHw4sD5CpkDzCyOTnVKdAsTjOLmqz3ES3X6yhFBXEExzDAn0Sh0gIxqx3k8m
8Jk9D3pY51m+RynvVQo4Z5AK/+1Nsbcy17xfbZC7IdtAUJKGuVsOH1HvOSFM8rRS
XqqIvbItlU56GU//UeT6dS0jOcvzQKGeU8TAxEoaiy+hut1YqEpGw6sxjYlVgy4q
/h6PhfBg8cKK/kIHTzNdoETgWenM/wIORzPUb1yt+ysy0KNVAHCz0LvYfW8hfN0T
8+rCAdUdzmZNLRMUNDwBy4M1Chzb7uqcQ5N0PcC2QkG0TqoftXBaOtu21iYVYH1x
N03PJjXNQ+056oeO5Fq4iKMB2JIaKir0UTITDtJyKSOKljPNjSa1m3n/Wt7EEtgd
UheT2A9g0qqmcbxJthjPlaFVhvP/Egv8KEQEHX6pCTM2k7m1OoAwPTMhK+ruTSRS
40cE1ap2UcSc+bcG2YsB2OaoDu9hmY6EOt4pcGrA/RmMkYFechvFhHFyNUcGBzRJ
va2bc6HvomeO9NFLDv33Zwt1VvkQmR+KxgG49hqnYXYCzadMNTZl8K5fQqEOIa1c
KkYy/jFoinTyupItntdTO2NySlGDCuPFdcjWEr5VLLtlFf7/Lw7WCXvPOoZVI+2G
wsqJUpI4IYKvRU2Wwp/1jQKtjAOJgSz5xU6tsmkAgOFEnu8w9YFKZnRWM2DxlFn9
KbFeRvfAJftb0+52bke0ZrJTLzustzs3t15c8Xzvhpr175lh1E7MP4GRpwjD4pQ3
4N8KFKIGHfL/zSwAgB8jq8gkJ0jiqJ/WdoUaJ284MRX9wAKTD7RzQa33Jrviohpc
fv/yg/p8W5MR199EDkhFVxILPUjTv/Wo1ozXExH5uUh+ind77bIAGIRWNconMXfE
3OPU0mxSGxOmyd7ucOL0l5I2uueO2ifjc9ahTFka+9T2W0XFjj3xoFUr8cw/ZyaC
R8BxXzK3yTj/ghJ688nxOYSbxbSblIwbPed1bHK1vxHa7xG33y4WaSKD6kGMt15j
5pJhmeEl2zN7yLCysHBgSO3s7Vb1s7bjO2uuHkgZa8M1Arp2ayghSM3wDDuurhXY
dk+o6ozRwdEyrn/jS23DF38agwPmYGkxJ97RbhRuGQ9wvnR6Jm0cPj4yhaXNDwkY
uF3k0xCvKfAA2aPGtuL7pl1TT5MhIL72WAzFNxILHVb4+A/tOPLIAIrcqp0A2LQC
NJM6HAl/LK5y3QkqjlN19HiInL3XtvJVuDGpLLx5VZ1cLMCPSJRfX08RHylIGM0T
OupPqWvHniL5lndU/jNOXzLEbE28eSxdxV8Ti5FCrKkHQSt8YvQz2CZfuIyeNMK+
CqzLu6EUdw5cj+UsUh2A7ySyvG56Nq/oyDx0788aGjM+QD/aMqbrlJB9Nb4JO+Ov
GoeC5RQRSLvPvBkyVqE0fUK6tqficO9aqcqO8vY2vVKqh0JbJIxlx2Jcg9KK5bzm
OfCMKOCkFWnSvmChXCAABGCfzHk/oqeKotorwNbgfyhG1Zll5qGNv6NQZ4fbIO33
KKzzoLg57ycv6yd2chZc9rwZTEGuFb5km98hDaELjjGfsqeqjG/FNq2MnKA23J+i
YPn4adBpxmXKEPMTxrgi1Q9LLV/dyTDpZbtPeuGs9hdt4Ixi2TM6hUEArn7ze2sK
byU/X0YKk3w3Qi60BzVckH7X9Bp0Tw9k1uO8MWFfZbJI9C/AqtOq5WxGQnJbG2Gt
h6gaSzPQanyKxIXjFriClKPDHCFMtMpK0Wo9wtnhOa74Gqq1NJcvWYqAHsmG4Al4
Vk8iWqlBXTmC3HuUhcqEKAK9bJn1cKuCDNvP+IT3P3hI5HOpctzFdCosjVnvu/bW
OK8WZ6plksKqUpWQETZh3FQ5OMPt2D38RQIDf+eKuf6eFcLGZ9G+APlAmjtGnepn
cGIyo4uQjK+/MBCgMLcgXFwWJNIBJlXreiRfSHRT7y2TQEqu/v6P6wXb+urDDcwY
2fzdZOdFG1ZLoJofZlakbyYcyESQu+uw7K28o33Wvqf25284yyPc98pHiO1obj06
e9CAIOkvi6vENeQFBmAxItNSXgI4slVpGoXi9/UePLsChWTHKw29BqYhYQwivxOu
+BGofrvI9PIDLnu5UZwdnUB9NcyOhi9IBkhplfujbESdPPmgvbXWR9FOKZD1o4xn
qLDDM1xfe6ZP+AYIGX3wQ2MFvp+V0f3X8aaQ4+N0FEY+A3enIc96SokSBvnCuAJa
LAyClViBkE4795PEcMqrUvDxedFGZwkDreIBPh5cEIraTuU4SIZz6iRNwgP6tR6C
DO1lA2Q3xupxdQDeRF92PiO0gZBjL99XljaNSjmPq94s9ypFldQkqZvkWzIpb8I9
Qzpxo5sPkfqSbwql/1NzeA97OZKYu7gMvEyJy4r2vZy97pnoOkfMjUu4g9mbxNcH
MH4MlBbTJLK7uEz9I7bjk8Kuy2Q6VNTLlUVRqhmdQIM8gLyP+M04B2dzShdk6Wo8
9AsdmPELBxl2DSw1ax4QIGrestc0XROkZ72jM9+YyRUlvgiN3fA2g8FY8bgs8fzm
fZiqSZ204cPBVfChqzUAhmYROyBV9xvw3w8MIUo20o60+ZeF7DI/Xted2nJPfMuu
Gquf+fjOEBpILRz1i2FHgMBzPuGeGPNuuFoKKdrjw9hJrVUqgLlKt0YvbVq7DMY3
v0WPgD36B9kt/q64/k82gY0Ylw4yrmpvcQJVGkwRj4TezCn32Y72nlQmWcKLfyeY
mg8vJXOaKzp3darh/7s6Vo2HwhaCT1oFEcsEeo0Zt37GTXdBRBGUniu+fG89VGNI
txpvUxPAiSON1vslHTy8i6f95ofYI7e17X7oaMintEwmpmvRk8u61fsUxviVfhhJ
Zd08RNjb/AiVx3cWB/v4amE4/JMDHHUNLXwJv7untjOg7mtSZcDWIHopa7/54fRr
JTPZzL5EQRMdgvyRkfQVwEoZs3bDOoIpj+yeGji+xBT1528gMC4cd9AJlqrzJIt0
JHKCB4WXS3vmEojRWnSYTPz76SoVQM01KGXcaubJqhYqps2TAdVHfFJANzVljL1T
220n+oFibqCU1iiuOwdn1vez9/RbzHw4qwuQEK429ZVe3b7BScuBADa8+7zxO9OZ
RdTImQT4hCvuoNImuBnTEpFdDD2LtLEhZA2aU8xgUd2gW9in9ss00ud3BzNZKr6H
xg+5KFXoIlHC9fDQL5H+RHQu1GNcjKYEq2XBgBZO/79AzBzfvBWRb5CAy/j5qSKk
nc+283nUpj8p+KxYoeUC55b3ZXLz6BtQrc38/CMZr47CSDWfxLpIkqi4Y0rf757G
XdeTcdlYBBsmy8EIs5H/nmBzjAda70zCeRYS6yjYJ3D9iNrNUsFr1/XlnhVhK8xY
oDUdn3u3NTLhY/WMPanSdNsbhti9bzA8KXJDf+ws10jCwhaeSdVkJ/FE/A+d2URr
elM7Pez5DFhUfjUXDiRXk77njqlvW1a5abKhZvZPCjCXU7f02ZEawiJoJbZk+1u5
Yfe9QIQtDkPSsByoEQ9L6vV7+C9OsPb7w3HSTKUhOgN4iz2PXdGJFpsjHQq+YTZ9
xkWQRtZOMnxi8n+zD7dzLU1/ccRwZvDzpQkAC7dDftPCkVu3vNgcUFsdnSdjXJmu
xa7CrKmfhGRYjN560tzT/3dDZD96ORtax81dn3kaUw17fVrKeoG5/WCuyjTV5gry
yfmirQsONqXoQJo/GTMnYktX0+5whWqVvs1VmB0Cv0xWP40T/LNSd9y7iU/0ZRZ3
H8R8XVj9l4y6Y1jSFVs0Ibbq2SgRYaedQQuvUaOuwcFtYJUhXiw+UgQSY2VAodak
aAeR5uBJFe/FRzCFMFYj3bHB8ujDppSdyQ6T0+HH7J/u+gigRQ6yolIPMDqoZnzl
MauPSqe5wOFqgrk/IH5GBh8vEiAVX3STgETxW/K6wryYtVK1eocfdfZATtWamlYk
lfVXFupKLqzxbzNMd4jZnEUtcexsNehXI7qLCvaT14mx/b95MYvmcGUiLgF+U9om
KpqZgk5Wvob2Q/UOm17TVj5mqrYNPKKwHxrR+c+tSOHYqH4+pwlzJxcgJ5bn6ejO
zYGdtKPPLRP3Wboc9Zt3zj5zRLF8VxBkEFSx9vkPw9NgA0CfyyI1PnKZ8yWPHLyC
fAXKc8mxP0GY+bVxmkzWssgLFcQHZ4IdsUuQCDs5DsCj01waJ/PqVM5zgmTQgIPF
TQeHZk8i44ZpBQO9tSWCmeaK3E2ornk6/aSJywNUxOJpWsaWQE3pJ423G4OV7qAj
FckzHelYR8etTo2mlNAVK7B7WqMYwRLYUkrjcVqICl/DxzdQV+DADudh/QtQRWff
Fl+60cu4NAS4aQucFcbJqCWMfF9UrMhW896oKUBSl6WKkBsF5ba95VfjHDPZ5chi
/DLV4prtdej+EvwbPBA6pta3jzqCECe6iMZaIKe14EjZXvDcZZmHqFgZrQrs+WlS
dDrvOgSxvDt8rDtv9xeF5JpcsdKYgvaRloXAfRPlhNvwMwF9P20hNiWqlzQJrhDc
oraeCNUZItiVlIrz9zXjmuFoePrmW6g5TixbMlPtIO3U5WyrknQpiAPFFYKcFPeJ
0uUS4nXGxIg1uexiQCW66Dlv69FO4Yl6o36Ham+ALIcMh9+efMNOk4c992/2Suno
3gwMFXRcy+OkUUwboqhhzgyYJO5pOXNROXtOgwnQjkgxwZfjKyk+XdRuJJNfUxYj
/05dNKy/BTyb4qAo2OzAM58kuDdKIy7dsuFgb4WKU/lva4ZPfiOz19CIZdKFKdMd
EEtk8DlQFx7DRhZBE6frrnIY9qcVcS0JubGhz81zPYUAZ7GwHCIj4jk1eIySM9y9
4XvMWZuDbneNGPjXKrxBrNbEJobyfrcRLU9K49H/mgQQo/YiIAmei7+lgiW1mOop
FU6rz5gpVNGLPrsf2rA6Lf930vYI6ojBNx3HsOSFN/d1bdKnYSrm+E9oaX4DgJCC
W7SN1ijhM5rR4Zscmc8FoGxHeuRUadPkR1SrWE74DyCvjwc2q/v6yUpHJJcUj5MT
8/Z2mxfRfH6jBYx8Etro5sawdKH0Qqh5e/C3HJcahH7RhvVEnmTtsVpGisrrcB7H
Yez1zwEpL5+/cowK223hdTj0UcFgGLbMLRujrZLYSnL7ZFGWtzPUH0/LAr+q1/Hp
eXhJ5aWdcOMk1XnUemSs4SyAUESqHRvGXAmwjskWF0rj4f111o8xTr+Y8Mrn9lCJ
yV+9Ms9p41P/mLZIw6o3FYVSYPSnj6XDBpVZl7FhQeNl1VrI06co2ykEtel8uNEl
JmQPQ9Y2QslGXX3JMcCqWYyrHMwc4FGTdY3RFMTOYC7KWmYq446+DG1VQBaGtpqh
a/zkj+Rc8If3zNkUSUvbaU7uN5YgHmm9b87jC3DP8veEB8WsFTJVhL6iqo/G2z7n
GXMTSkbNd2bYYv3a9U/uenMNFugblPI2k+k4KagdUG+Q1JuABf8RmEYZ/2rMRkag
7G/jB6fvrYcPhKJM+8MqYYhUeBIFFMxckTWpAF163wKnvjqlfkcyWtoHUsESfWcV
mCR9kkJuypntntSEdn2qCD4K4ClSKkFdgH0033/WHxf0Ingz77yUeiB4fc/v1lnQ
fUk9LEfEVDTgZSjQvid5+9O3qC/IUSSiZ7JpUfp3pITY8OwcScq0zJOsZcODwnYC
bcBcABvBiLduMR1aU9y2UulrO+F3jCjrBbPOaN4SwQZ82TYrTcS3AYdwI9H3lHHG
EOQ6TMnNQcSZvw0vD4/NB+OyX7W7WHV+ajS8hrbZUPcFTkNIB+Dzw2mJDUEHFLiG
qYV/QLj6uFQvroCJbrPmWVB6BnvbPmuEVpQS3NSnz3Yz1WZN1XDP5fti8h9e1EQ7
UlhLDrxLrj8lby1RZWUBA7l1gMRaqa5WR3Nud0jTbSqKqi5bn/QAH5kDanNXfLeP
9UrQdbjhoMW+Ib4qbYCP9SJwsyHa0Od+Sjh4undwlkV6jIW5bRjlUG+ohf3/Qc8D
eZzMRfkj4JOAF7Ci5wBW25IHcAskGoS/m61hVW+bGhNQm55rtKqGKGO+q4HY/4Ml
oLf1PH+PxFVzpK1L/wPyjsLGUVxF0kofoZXfKMNb/Np9mWBsFTNiT7OmVb3B3tn4
pbSwaJXxAUKJoi78DoLYX+N454+7ba2w0EA/Sx/i118KMuZqjELEDRmcXd8lmmAy
OurRAyJTQG+EvwWMazBCGHfaaxKgMcwbEpKj+Qb7CwU905CrNvnTkkEULm7rfY1r
5ZMe9BbhD4wOElJi+FP+GbR2kOlbrSe4C3URVDyt8AUXFWFDkBPePFXl7Uif8/lC
1gi0BuEXN23l2d/03e5509epLmhIAbKLU4aRiZ/lMBJIktYX+fOVS+GfHFnyeLLS
Ur2rc60vzat177Q5EOsknLE7TKbxv/R8/1xUTzQMnk9Egoi9ucA4ME/o9OSTBn5x
t03xH8TynXU9eVKVOP9PTu/q7XQksBdPza2qrWO8EGYRd+C69t9FmLECbJ3UsHcS
sa4Iv8GNv6CzIJtzlro6o92/xE0KarA6ozrWwIpg/ZOTgaLTabE2bBGn8rqHf1vf
RdylP2WDjRB78aFtkYquQQxEckYKI1LUfGEYDjfn9aJouPSdjdvneS8modzhfrI3
5D8yruUDdbfeLW6ybng2Zs7pIIWgcUkFE/3OTtjnZRi0zXhmwEYFBtl5X7WYD1TN
IfifA6euNfDmjgzPfcSF/Mrb9KIqrcG0BLI1UWdPdt/CZxc1VCDKlCCCU4xEjG8V
M6yvVWhe8crRYFja1ezkY1X6Dode/TQh8lGFiDnpy4Sh800cLCqKvWQ3nGpWCZGA
H4gr31lcOYZc/z6dhUL2e0h5Mw0p7k3CPC09BTCnDli3ThIxFdTlaa9AgdO2VXJ+
+CWi17mEMgoa2kdnu/chi+j0dfgwDChkWsp+4AdaX3EXzIRGWCG2+GDYZ32GP9Q+
ZVrKcELVUmCQPdGRTMHk4cQQawLNb4s/s15Cbf2yOMHZhkuuDmQpx4sMmcT/kzkr
9Bclq2YepAwGDmnBdI50EubHAVPuLLV90Xe52UMAy+9IyPqxj5QuGldPRAPDsLbv
t+c6O2AGZdS45rfg5YEs5EQzMYTIab71hNm/9UMujs7A4OkaQbqc1ag7p8UXjRvM
8OWvd8k6ZcY86qSJkYrQ4KNU3WYEtfTcMaA6oWyQ3Or2ClHNLqOZWVP8XiR/+twI
BYR089JToNC18/GqvcwCKhMgzKQjlFuSfmDElmmrVI4tj8NSUN0bG0UfEFoozzXv
YH0aLX7CueyMMssv+C+FMJ17zsOI9uOX/LdOGaURtW8je2xFbiBEMynfBMi+dBds
BZ2QooHEIlg5BFAGPmC+aQTCNIy4QHLzsf8u3M11SHZMYulDY8/meoAIAOds8F7Q
D3bzD+V6Yl+Y+q6F+RSzwLjWd6C1/+kpdbCeHL2i22CJVLOX+logAQCbLBYkbrGP
tKD0H6T8RX69cQQp+IDP2GS75XoBlpfDxWrLxFOctL0untmevn8wZLQFL36rIiO9
9Hyo1xMKcAk9n8Sv+w1nTmE3TcYaeOWnVopdJCpbS1DaTgz2287c0QXBUyhhGgrK
TKUYg6kq4CvEptrxxCH5jQXJYjoSOnc7aAhAAXl7ne/HA4CLHFumGTgA2bPmrnZY
FNHJguon2socmHMOKHQUSxyYBS3+fE2HRwrxZQG67Y8GBbREin9xKM9WNVzMYEFe
EYkgrLAlXcMhkoxziRSSrELItdQpySmo11Mo4UCyJ8pDkgv+x3nN4z5iJSmP+O8o
MiW8a52/zBKZaqx6Egl/k8i43m9B6RhCOogOTnHcCeAj4WNd7t6CZWWfb7n10+Eb
LHLmlvyGOW8ZCeC0x7nryzDFT65XxXOlo0BVrNyko4BI8W2pXnuEMb7iohuBrndq
RSh0sb77C6eMlTQxOnEPOPn2qNkLhNc3z49GJ3ymE8rS2RQa2pk2/EoLqx1hatDS
vU6JVWFhGNguQYkEw2sGXEv6lEj2vERzG9akx9GbCDPU1HKCCpBygAyLxTRYKCpk
44I9aDWwOZ5pdZMvq15HvMVllhdUXxp/QQE9qvJPjmSdI6ukj1+2EQckNOrHNGuM
OojWKEsVbPQ5sp05a2FftQkNYXPXRW5YtvaSDGmRNp5iMZ8UBVge04KYdYGbUa+J
+nYI/01DHaKvPJiqZ4afW/vCtZj1Q0FzpSsl1rdSppL9XVc+pRhLonASUh9oYet0
N7mL2Bb45c0putYcgqGeYiycQOqcelz5B7BhqpIf6TTcdrKGwiz4qJp1rryPnacS
d632HzAcu2TK03GZqMT5jxtif993onz6Wl3x3rL0VK4eOcYYgluDumzTZm7Fi92E
xxUEk70xSsKxZ/cEakyWH1d1qm/+SyF3e8SY6qA+eeh7Cj/DSRBO78xtU+9UUc5b
3SF7u54ChD0HegCIlM3HaBh/uNgruR7aYHC1HABWcJxZuVgfTgw2zt6zoylKYDws
1Ol14W2LlXVEWDC8vqijN3yO2zxT/W4qx8Ku2E8KPaHs//m/R609vjP1vQVdMYhw
AzXBjCMNKsyLkelnt31aUDh33Q2cAmFNXoNgPjwA8kkanWVIXv4wplgp8couOPVu
3C4NEXbmDlpQhhzCOnZnxfhmtuD1JZ9rZ8J26SufgO3nGnkNKs/Sys758ouAzFyl
7JUs9QWSdRRkbxfoAt4Tmn9c9/R3mL9MTc6eJyWDH7k+O1IqzB8SKbwuve3ihYmL
yQ6gHAYwVPbP9tdDiHwwULWhiFY2GEZsTswmZ6UthWCXqFC3f0l4Jvc6rRjcRcXL
u8lFztkdOUuvubxCOU4FxLymhKJXS4bCIwGx7+VM1dNpY73YS5RA7xzsPSDOVJrl
c1mjEW+pqfglW61+uRK78ZfaXxetqLiSeILnx5qGv+34G6+X94Z0wgQT/xTtcJZ4
BTLommRHj5hB2bpfb2E8aTq3kYV6pMyucmhsZtMAZPHFumqEJ004j6dTplAbEvxp
mY88K+jMZ3JJm6yVywB28PgVSqnAvm3oM5rVVbLlIlqSKhfT4e22arknrSRvfr2p
z7UMdYxwJgiwEINDmyGfDCddUQdRsHBEMZBTqcvSjBxWg7UUrYHffhoOwXDDKT9l
xi/E+A8GvVhW5nL67J5Ge4iV/0PZluA3nw1wjDxO33H8wx62fi8AYppeYBtAoPN/
6n5A5C3/fC0KFlBk76K8tnTv0lqMiYFo7ldgNjKthliHW26iX1SAElSlWNibDRh8
nC1AWO8bDhe3H08UBaWBB/VHrkOomVLkGr4UsDvWM1um6J7sucuaLGXDIFaFayO6
Te5cYfDHswgSp1U4JTCKAYLftMVNu866l1HRSev5s9yPa/g/+3ypbrH5/d832ojF
f7C5NUgAbUxm7CXXu/q6HmBi0ZwweSg1yF33++TlKsU41bVDA5EJv+cbUifr3vnP
LFxFeFTgTXBCmqRy3huzyEaODnhVYtKIjvivNpJoKE084SIATrr5ZDA4jRHseUK9
jCL3CpjjasgHaX+HHswvU86SFad5huZ1JQcVeUO8m5DnLdQSRO9+T8ZPwXu4LHlF
O8phupRBQxuE/IrUG8KFm/3X7vFOl+Wf6h5JLQUAuWh940n6NNYTwqJtNz0J8EtT
1ADf60t7T7aR2BuMl53QsdW6pO6Xl5SCEL+foUiRNVVSb4R0bQY9qas3zEN0tICg
tx7sdjNtNrIVZmayImkD0anO8b0xoQy7JwQwRG/topjK7k/Ah544NRpHvxAq4np9
U3rhkvcaVxA8qUcYFnDyw//RDok5n26hwogAj745AGbdE0bw9oZI43bgyhiveKNq
iPDTXKyiJVwVJCDlaX8ouceN8Vl+AhKMZ67tMIg+TVdSNntPi8m7LrLQdpjnoFHl
pMPsKBDPgmmkZ50PcmBbI817rnYbvT6GAkZZ/oWWhZIz9IBZ6jk4lxJu/tgBe0cO
+V39soJX0sDkFJ/d2noC/KeYm9Hx48CJfsEH9a6Hz2WHZdiItzobPnHVztC9D9Tt
VNNewYm64SmHb0QORervTaQPPhqm2/Jt3un73TfeWUu4gQKZbQGxqkD2SW5RW05G
OEKoJ5VZ+l2G4080TPoYUWM2mWwR+60C7tnWLXh+tVpC72AdtM+5cwpo6p3u65K2
gbVjSD21Fu5BPvKTP28bLEPmHRmq1W4qb0Q+v2VZiot8Qs47Cgdp6sDlNK6TsKem
4oRnBAdvoaiYR9JKUDxF9hh8qGt3M2ubjalf881RMw4TrBwczamkTzxJFh3GtNTr
EzAdWq3tq3pH3xB2vEoH4bzW1lJW4BaqF3jVeQai+9T9zCpujJTb7AbIPu+WERTp
jFGzTNIjga0R8rsn2lV7LszsyW36/eCnnkLDoDvX3UlYdxmDtPagqHKMw3r0HkPm
qnxiVUqY7p4S25VEc3yiJDXb9kcfUlfZwyW739fUhVLE1qI0AN/+DqUHKWsGNOM2
RcCt/R4gH3a/yvostsvOrCwDDb4dhR6jyuzb5+ZUL6RihJAZ2MNcacjIc47Tg/hz
+keT3njaBy55Gy/qzi0zbHO0BFPuS7pOwgEjocyB1oyo3k5+JjMQJHy1u2hhtfJF
/YD4x1myBfoh+wlr4Roov8jWHrQxS6iwghjfGCnyaUe4ARXy9VV/SCE8kqaLopNg
sF4R32JI9ID3X06UktMGsQTz67zFW0Gg6jAZTscj2EBuwh0LNz5yxR3l8SL0R/IS
OQVd+ki6mXAQL1I1Z1ZfoaolbZXO0cFxUy+N+4GeYX0KQR+Ce+Q5miSEaLt4t1Os
eDmYYbrdj5+JD/nmgEHZdMJRcfw6dCLcGGc4l1uxwEf2Hs86Y9wRfvgodanMHG+x
GXU5Cr7iXCGwXatlCBU8ddb3A6hc3M8HZaI/mZ3xJ0CrjOuGIfUYeKOjiaXQit29
q+f/53e1OML0iHuxOhBFYSKDM7y0hAvgXA5CrkwVEKuIXy2fU2/sNy+NZQnGbNhW
MKIhdZ3WNJ+/Jn9nlxDxcyg6Op6GzuwvcE2iHfZgZuBPUuiykIUL9N6QbFVooo9D
qWQA7gm11zoEX6SiVIhE7YgmIxn2mxvK7ZWSG/heC5HF0IL6V5XSYn5iJav455sZ
2h1Oz7oPtCRrCStROFKYB2gSP3W3lwbaPAxFGJYBQRYig28jRMJgLTj+lKzYIMqn
zYbAF10oc+BxssTWTR1IdQFNAqsGi4pZOWAfCJpu4WL2kyjdGmMnnkT5gdW0Rm0f
HK9FFl9nV59nTgpEOPiEpuKvow9ibIOGEL+xUkAZHqyeGlhhyoJIlIwdZMZnnt3Q
QaqaGnzAT47YRV0/1rumnmNbS1ZSv+JW4Y4x87HH2TLFuviQBZkbIv9gBfwXm10K
ujovxigmXHQIFJvh9LqYHT8V0oyoF6A2h+3ZnXomScU/2VjITDriFDoYd15uVoXa
UWSenEqo9R18SdPG7KYP9Fwew9v2ev9pEU5w8yXH+AM57we7odlm/+zncAT5aPcn
heBrve4BmgwaiOFcRjRpl8r9aZW2xuw+h6pw1zxfp93OYtY+lAaNkS2X6QyinKBQ
mKUD/nm8lL6u0t1gIZnQGjJAXVWhShgE09+YxET7eH5+E7fj8lOENz1RBQZVWl4M
iue2W5LKxCQOdfZRJJSZCFucY3A1ewYI0eX4ChbEsm9hmsKun74JT2b9fUrqNiy8
IJcBjb9+MqZOWNpExha95uu66I3VgfrxhuuqxxkM5RxNCFeGM/GDbuMxOouvTioT
KSSVKwahX19bL9Zyray10Swh68Vlo7V3P50SkzmPZQqsxvsRd2zb4k/gsFMQEBbb
5jitt1KdU/jfJhR2UR2oXMQxdSgYNeUd8a7AZrlut3EXv5wLZXspbT48KOH5gBd9
ECLoJCxA7LSVykSIcOluRIMT2feomeUE7V7bhm1oDsemJ+sKoCXMz9C53R8uxAvT
5Guq+Ft4VJSa82H2e9+sDKtZDHDnowaTjpmryTbrBgMaq4Rp/myqfy4nCtNIuDP4
rdtDXeKJiToozYu67kEtP/NvsurQwwC8zqYgxpfR/yL36ueS958AEo3BgyBIZjzw
NBFId4gqZ4MlAjV8WCHaHMKWGGs6TeyFdizeq8i/7f5rUjU6Bwgx6Zs7f+tJA7og
L1uJD0BRaL0luHtafecie8iNZ/v1MIrfJy8KNa628XOi8AojlhSduljYwohKXFEe
dwKknAKhpdgv2uF7TvAkjq2/N3YrAbuddEbLUZfFlbZt0hxlJFzibGgGLKC/+6YC
AAIgLHhTShzePZNQmknoZrAEpTn0rwY/RDatIfykjjs+OkA1rVuSVOgxZGVmszJ6
t5+OohtL4aRLNAX4BqSyD4f321gDs5yRmbnIJA0aeEsFMuxnJX9ojCAgSCTVZCPZ
PaPPpdH6S2w1x6vqwBgx73oBvmuaJbgdG+BZQbkaAVNUjX9sTArCUGJj9O0Ygury
CNrUn/QdhFqZ/mWxKmFGS5Zh1IEAMJUe1sjnXi0XrsQsaqsbygfDQKwLRe6bkEVv
3ko1aVCe71yDxRKEkXX4gcDVjdtNthAySxMhkQ/+4iDjcZZJ0B9yhssi7lusr4SD
q18MwPT70bSef/wjC7vTvpZLM/R3Wb+nieYxd/ByG/S3ViMP4VWYtZwZ63Bf0x9p
CWbeA7h1+MWfaNdSKzOlsWnkmxQS414/pRuOJGdpmP4eMqWraTVKdg5+eZMDw2jp
o3cwLGI4WxdvCHYQ6y1jBF8T+6qlYum4bwqugnnFCZEOW3AAIwC9XmZwdlbaAiWH
eQ+AJpVq7H0Hbj9Y0FMeO+kRfxU6orgcXkzkQGaOeQE7FEdCaIKda1ABQa+Gqp08
8MTEE10tBlUnWRw4trQyG5E3vVbLHIOlkSSBmSEBHjKZA7yASM9vLh2NQijq/8iL
U4jecCljq/Gd0OpI3MF+wsybiGoRbcNekObxyH3NEsEsmrkJxtjRuu6sfPmXENL9
9P4a/FRURaLMwF21GyTzv5/IodalUPwROVsxRHA56If7DVYhF6ka/CmgrxtY2eDM
XuJ8aFasQRCriB7j/3H3+ef0uIwiv2uDyR92VTvTqoCT1UKYL/7vqC4lyKgfooM5
5IPhw7bCTl6dGvH31YVP09CGMvTcBFfN/ZoHHgtmXqYCebmAXpOgSKJDEt/FKTjX
y9L3aJ1PXgVIt94YlYKw2wUITwT8qzonM/+IkEH+hxnFFn5yLa4lmfL2U4oqJkG9
Ih0uCtTRYFcon8K4/GeVBv2D7zKzmX6oqfhCQI2qtUalabJli40xzZA2j40dSXIm
dc0l7fIWFZmNdDsbWbLAH12AKGJ2ZYr1pPdhkmxQr6MHd4RDd2ZnT7Gq6sKE6BO2
VfYNyRlRoF7E2ajbyEk8APtnrfxAOkaE5cAZb3jrIAu5Cg3KcI9/udPSd3lxsqND
xV+p028RGfrjKpAZdIykTlJ4vixHsTIu0839x46f3TZZcMAfxVY3GYjSMTi0+4sL
l6T/GUbzfL4tlg3oAY/3ggZx/IrJcV8TUugEfGkxvGNDMf3iV3vL1wzpPFCscCmL
7FhuVqEnSDplMK+tKD/UbAx1WNNWsYjz/PAXIdX1/qF3MYF+1aXUZln+oDW2Pe/r
uAzQzZDvW86fm+7nFzQWmC3gNoq0CprMQ6vmOXYuKIqvWPG8vTD41vjoBEA0EVYA
D6e8O0Yz7KvPherr07GxmVulwTDtAMTfIMYKgD+0fe6U7nW+vMBVnb3gXp3aFO/9
xPGFD6tsDXLx2RNKISEHkZNjsA7AuVEUP+UDjjdw+Y6QYWod+IPZMgR6mfSq7kL4
3FNkoqxdr3B8m0a+aTkcJu9XQFJEtNGjt7y+tGWn2pPqkjYTqS+Pkkvm08my3NxC
3f0VE0ZVBaQ57Ecpyu3Z1b+bZm7uqWyMjINuD2mNr+26MYKaUcMb5X2KtRR20Muf
6hn5Dp1aMPUfHoyd0VcA+O2mUtoO/NPPZN+4GMYmzDYT6/oUFR625uR+KlbKhxZt
Zxh0+r+kChKzTFDPL4TYtoq9l/urYTl0I7vCLgMe+C79Gcz+beA9b9j3+oM9g/9M
cev6LpssrO9esub9Dtat6vgmA8sT/73TOXl0pu5HgcScsn1U3+NzEUJkjX6haUya
OAiweO+KwZOKkSmUrECQDRS1vNa1mMfxbDXmhXtCaU5EU7k6iLHUzW0pV0MG0uJF
SIZQhOX5sWRwq7F0Ozg9innRFaOpHWjBWhyxiG64YJ1FUkqMxcD9pmNoyoIqDCVn
cB5dEdstyyJEHAu8fObncY/W3CLep+CMePaYAAQHV8Ire+E+lUA0aYyrJ63SPo3Z
kKMDoOZXfzQWeLUr8agAClVWtUpmoISUzPB4dkmiwptxjGuaLfTb9fbk+uwvrR5P
5ScL1wYp4HYC9GhEY5rR7A384CSeBXTkumWR01+uhpns86y45XQ43ADnkjBOeqSA
ED0MmoxnTMF53l5kgd+6YOfwzuwkU8tTiW/ls2JJFbiRWIANh2OllO00/rMnOX6n
xkwoYe1T3K3Eoij2pnDeFoMQA5wR497QZpquVH8QJ284Fkwf1HuPfU+30LuutrTl
Dlft41lqXC30mG+WpVCd5e+Bi9YYXponqEMRktIepV4MCts0lVRt0JbtDgWDa1me
weMrSIFEukyl+qWzhXP5xAmlnlQwykA6QPPgh+GLcIMrscu8FRlUmg6LKHpKS2lE
A8vFkL+U//ks7xI+/kBcZx0+9tKqlkQTQL+Fjs2iKEe1PR6P2bKRXX6JJqEdYTJr
SQPP0R4OIEG3vVbJRDqaZtTFxLYxesdpJRIOUf1OnKf1jrDtvHuCJObbcMRGMB40
sjrj0KuDcBTn30xTNUqjGLohkUSUFU9CzFnurRsNil9DUUhsFJiK3Jvk30hJtciw
ZisWv7nt90IrsOyBEXp2p1wRJxX3cErvkV1IYL0Wde77ZJJRzIgpUcL3HkWyi8EC
Z+rjCpXV3TwTkLqW2FvF2Iy7H7/HrugtWBc41K1sBb6Wf/aBAWp4Wbm02u/Mu1vV
x8anWovif0BT035/r0mJ/tUc85DzulnqClQDxV5E9P7ApnhleIzf6S677Gu9rZOf
Jl9ydsnCNOBxGraynsX5PWTgtPM2mrovlxauBArmd2LDSpMvzHuGZN62VijcJnZe
Cp7syVmM/AdwEo8o1mERoveTXBZFD638IbwYJQoGwiiddkUF5rscxSdiSbT0IgSB
yKKdKHvsYOK93Ggzl0W8lwe/Ww7Zo4rfmHpeHZgsZexEbuqbklrcoq9Knf9aa5Gx
TuQc5zLWebkzggbPTO55M79UHqI9Vvbguor9iB4ct959yeKyS+ntZwvpcldbHl51
v4qxgOc9VYQb8S7gzlNbOd6wDUcUm1vh8YYpp7u13gOQJ4dA6zKrzFkSBYeHKuVF
65iCFwE9imYT12CWj0aRC/g1p4UNR8shhcg7wUzQxBwHywpDCU/44lhMCgGRJUj6
gjGuxBgiQUsGxvd0Qr2GRmJvugIqIA/SQoh2qCXn9jBXGVhrobJJjEgYM9YLMOaN
+dCeKuQRz7OxzDdG4wSBXnasii3Vph8zVDzxqCksbUkrckXZHEX1gbrsaPMmLK+n
FaonGF7JrHOE9yc6i1btXjRH+jrKCLZpZSahSxEC1HdV1vlozN93MR2o6v0FIhrG
9gaWGif10jjsSDSe9ks4Dwr2p9XajCzNGZEMQBLQYih1Gj2OI3YXW19sf2kvM33w
Gf3mZvQhDOmJ4495D7REIk9hfhVr/EYTGVtmFrCJpOmV/QzUDOPA+YzSffrulgYt
GL2ofa6giWl+I7ukvfTswXET8St2QqABCRqTbCYiL+OXE4WrGsBiaLqmNQdQBRKa
z0Tu2T1zkyUJ4y4dsWmdAMOriychYCfTzxFAjTGekYoAiob5BIr5XIl+8ksjfdAu
41yKEKbdxG8Xmf3w+ZRh4kqyN6UMQwfXwgX268x3daYh9C3Edz0dzyma4uVrt6LQ
UyDh/g/9E55QeXGappj0+mzvk9tNtxBn8NX5MbMIyD9dOoWWmqwt13XOmx+HMI5A
zAFgXP4GjCrd8US/ID2N8BLfEfdpveqUTi+RM6t2EQrm68EqxVcjrzzbxpf/g9vN
L7rxPjFr4KLm7pjxgTcAYl8VN4gRS3InzgZ54JHSBeq1lMjYUGwOz/uIKhHuA4KT
HJdG8iFQJSWmkf9njRCjqXCWGmFaCICFd1CjlqnV5xUmDRngnoqGWiMWl9LzwG/f
G1Sq2DHVIbjDakoMfWcGo43G/uoGfE+4wi8PhifhZAHx827eS3ukmnapohHPbsvr
tM36CB5nLTfEyjTL7xAvbROA7bq7xC8rECbmO9bDSVj4Js9Llhcmoq2foL5zziFr
OG3hAYPRdm285wB6F67xY/1kLHXkzrBsU9KU4Kcl9J0P0s2aqp6hApTTDKgCkINy
DS2WPvYzdYph4/+i3lAPSexjqQTtYApM7M8ni1Tr4QYIgo8eeGLjkiV/YWUw+Paw
+VWQY09RE8+4DiYVvVjPxEL6CQomSXy2E7CYHEjwWoWGEGULM2K5VWQapxZpr6Dk
hu181lgokaAgbBlzkXNZfvY9uXEUHJXlLB1Gz1RaLj+YVPRmm8lPWajwz5qvY+8l
gekCb/mBlKwkZF7TVRdJc8HRmJJc1TGnwvQMLpm29/ppNmc2GnthHqAiWZNa3J04
crQuc90O4DnUcul8s3h+yEviiLFS/WTt1T7JnuMi2Q8hDxwrQvAKl41zYvxugupW
JIrpFDCafrCfDFLxa+vtvOyscFSg0CXHzeJvpWo6F3B5d9vGXMIsdOODItiJj+5N
fcrk7Nv0racm9Wy8aopsr+FBerqqeBr3CCrs7Pm1jk4i+9SfX4iyHKjzI5CUAOqH
y5txuwmuWD9D0OIIXXeHBJHzpdeXuaCzT0uSDZp1ocrwxa+CQgedJV+nZ+pOAeKU
3hcOcRxnTdSLnFcFysbyBKsDBFrVaStIAmCOMEilfozoPqY0TOg9redDH6J8o+xX
noLUvg8g50ngXtoGAVIx1So1HuBhruAqcvikgnLBaIcxhGJLAfXMrb38B3/wlJQl
ZmYaLuXN687tezjbB0C6fOm4l7995MvsvWCxpzvTEyAuR1QBwfNLKiTvAsbRVS6r
5aPwJj3MhKSkDitIkWnYsSE6+E6yKz7Cotr5f5I65o8efWuMRlP25owMEmSFruMR
a7DhDa+SiR9jM1so85h4VAd+Pj6SMk3G/zUy3UHc6SimH+vvGjCaJLwXWwProezh
ryP99VIPD9lg3ohHv9m6lLtzXGdCkZ8hY/SeCQsWNwbclQsCL/NIJPqYP30/seoX
frxlwGE0WAXPvNm/i4BmiDsPgzUbra8dC8kCz0yZg7NPNLR7nsdQLV00MnxoZCeB
QZR/wH8Li47siGICPoxufrQo+KDxnWfaysrC4yIY1I4IR4EgGyQOHEO4XaqV5qUW
yywfsVfSFRR2j8deBQxbY13bzZushV0a0+ACEeP0bH4RKy433xQx904HOnjWAlDW
YyPe9buMek1nZFr3r+HU0kC97js0as4m3bz3e3kh8lp0ZJv4tmPDgSHaK3smoE5R
5Ww2+N32VmmcwcsA9racaHDzqg9RELlDaI7Jk5HTAxcEBCEYSE00dLOg1DxKEyAK
ZQO4eUQp8/eTFu065/ppJPVhn/JJmB+f+iAATReeiSKVoLoHn6XJWszsy81550Nx
iItzzKBcdSSj8ZqFMVPtffgHCXFC3e3bVb5wTrlVaazkODCC2rjm32sUrSwK+Uww
JocUMFtPDBvYxhupGda0Dh2nnt6Xhl4Chl5JKlVIy6qWyPmRysvC6hEEbegI0kdb
v+HNHvF0b70dcckOsPXD9r9UqcXW3ITTtuRlp1uZ/yyoCFUkhFWANTRhdfbk9JCa
lob+dju5zBebk+nj+jgF3nT6RQ9bhnu6iPoImLPj+bcNLM9lvXPx1i34dqZe66kQ
8w9ZygLwbVDqA861ZmCTKT3D+7HfuxO+B8RAlAYMVBXgFuevSbnrXNzdl0nOxo+2
SG6+tWe6COF8+m4i1JnxPZPvyP/8e7U1e5ktldhmLzvURLgSA51BQUUlB+CKbbpE
lIhTtLXhEGc7GSUwHrXAdl6tLo+LHRG7GudzZl3w5k4mFUildumes/IRImLUTypl
f/jJYDOO/D5gfZjABrOMLcAbkbrD8OJsrftvV1sxdczTL0xh1CQp9O9hCv8ViobE
jgn1aDsO/GEEOLqOayeJLxrMPotiO1NAf4WQNekx5gA+qHtKcsbSOqpzjpCOpAQ7
iStgkIPpznOkcmz4KXdNadd/LYNGqe/CmBfW+sdd6RUc13uza551QA14oZBAJaPI
tlv8UZ3Lv034ls6a8WVNfYY8VeyUZNgKdtE3k4gAYdvFJpgu9H/Os6AMeEcg8QpR
Xvry0DbOwSyhvTMhUJwHahIlX5Zv5sK23NynBqsTUnocr94jZbLMyCpgerIcBHPx
8qrbqbLRJdUeuuacJq3GkZERWdeKClgAw5NHBLlLykADMJWwMfm2wx3+9GaoLrs5
Zw/mtlipP+8684q7OCB7xs8wrh37vtuOEmT5QoLO6Qt1tG/2K6bbigB7PuixM5F8
CMunLXGhrVLvBRTRQ81XJDL6x8CgQu3e4KmM60G9XF7pToMGuz6XiBJeQ7Wv2Unn
s3eSjTxcU87eUR2FKK+5LCxQdJEAT34Evh878gNUHlMTsq50rtIqE1PUsGRoEFyh
qILbWztOsBATje1yz2B+pmEio20SMVX8CLZx5d7COR7aGRTTFNoP6gpryRUqOrty
X91236oJkpHaHfisAH6lGANLkV6ffGCV1DVM5LSmUf2hUOfvgK2n/UQoGgVamO8H
RLA4UyCATTTI2WzeEqolwqlKtgX36tmX1e+/BEBowzJvv2XZ8egM9AZDixqH5EVy
H6HKe0oFxjkDjWAMZZ8GqkAUwT401Dagwxif9mn4ARl63LNxmibdM24PG2oPsI+k
yNoEnKS9izqLZNPjUkxaZ4wwq37GMN+expaHCRhBOyXMnQg3s2m1oGsrLXxBvFD/
CtimluzeqBAsXLHS6KvuvJldoNIYODwzKyDM5a2M2AH6xLRjV/ngGSoGCWlDbf4Y
rLKPAFlcthsMp/N/sXRqnjAqIdRbfphohtgP66miFNou45d2PC92425OtEoCFYKm
ZQKSu34ifzGZBJ42XXqcLmn9OuSRiIpv7MW2fCpQ1oVyaypTS+K7BzjlPOSMUCzZ
VsfhV6I07uikMvLo8Juu0YyNxvrS65byjZruzTYBzqaO9hq7RWIWk9h5K/uD5erE
fhJHjBdPy1Pn1sxN6TICwmWVfWaMSC5IucF3gNGWTC9R10Wk7rY3ZNsWWQUPBCKx
098AzsZrQ/IR/sImQXuJVTRU0MXM0MRqdp3PXMC12wH7lwkIxtHxGxAl8hlBVGrq
xSkKno8+GX5B83ptdo48fgITQYTRYaoDn9LMidLZ1CrYdlSFYhaBivwBzGgyxhnh
7OIS8104grCzFa4u9hXieIiujMwM9omCV4sKuOt1VtagWkElfbaGpzKduMKA2kZ9
nXusymcDl8Cv0Bbga7DJFf6OidNkzxlTnNMJ/Z9er4D2oHrl2UMa/288VZEm5It6
MZiSIFDmO11bYrWO3FwNJxOfcHIvh4llKwGsEFW7hUAEof6QndQNn+bzdR/bQCXc
E+h8WcIXLrsKaoEB1T7EYRfLvAUULWH0sjb05Y+9pB2iby8xWYM6OYnSYU4Giw4P
yt1y9dGbVQdXrPiJ1ktT7ZbRyPCmFNDJoQ9YBB44jEE9R715Y9pYaqVASB/ewk5d
wCMPYVaqHtPgYlZNtNXyyKZxA3p7/8Ug0i+QK/5v0uPlxgWXM/5A2b0aDUcECZ/K
OKGmnk44f57VfKBhOd77ASLEdnd3lv5Tz4jcwmZgMMMvFiD4MDd0BZEKbCkzYIqd
090DjXQIcA+f+XSp8ufi/MCm5K4KzPqP5BDrqaGkvBkCasKpjL+4iAhs+baohKy6
EBo7Bx0zTp39cJj/j3RbuP4xBT0dT1VUhiTGmyfIPpDsoKLwAMIcV13zBWcYdJNs
6H5GDoPbURklnfEaJFZ+1gpuCZ+sXBxWdOEvVnHY06jzA/z4p+X/WsoXn/maXhQP
PrX+3wwh5zt268ezgy6Ggbyj9xezUlsvAoJuj2VV3v3p8c7wzRWEj4PaD+7dR3WB
dmFjS0TSmRK/BrtUIhpOndJKCLmMyOCn4U8E4y+ZD4fz22nS2Lm/M0DKB4qkU6M4
4i3ZmcqPVXS6rgdK8DkyTe+erdTAVkoVCJd9NAQYfoqCg4jVmorCxDyaB+k0GFf+
7omkebJTDX41TYnk0Stobzh+ypwZWPqzww82QyDHgNJTwffSZP7PspxL+e8B9+jD
taNkvvbq9EfhwCcdapFzEDhuD1M3WmoO03irHSd1FbhxS8RnrRTYV8oIssTKgxWe
+k2rvbZ+5KKpt03HFUh2RvzmZHykPxlWOJQMYbN524r8beXN6/LP4RMu1/oVd/kM
4LltFnfrnJWSLBtOmzC0tm0r2jzKswVaNfERIJWCGo8Y0mJdxVrVPmyihKpEvIw5
FOi6wa0uFAGKgLuGD8EQAv4SkRNshU5VPIKZIGcn2giHh+GRqahpeJvPbkbj3FMr
5fdKMpC0A+Y54cEy6R+GAwQ/qP/k/T0mbJEqVQItX5jyUhGVmMripaiW/TkgsXhi
JiRGVMDDD5NTvwrfmTmS/XVZZr2g3e2lGUgC5XMJFIeFbq9OaTJISxWiIEPbKvVg
StuSyD6au9/QzgTRtTAnL/lJXjxUyiCWelDFabEoMdZ4bFTEC+8puIpBFciqjqEc
+nJTIpG1FgPt0Jpr765sRvnL6foTvlLVW+K64DigGaNMV0E8WiZD6mNqsrkw2OHO
5O+eOkq/wir2p26NXJVFEnhsZlJcA9zfpMdjUpMx17mWDzh9YOB9aPdnu7SD0xC7
sKPNu6aghmfdgDcT+SW6jeVfCWkBaV+5BTFtPHMzqA8auqKp+XGn84MNqLV0mNAp
1mR21yf5TOyIN7mR309So5j+5Zs8FEuBD/9pq1FOnwITMfgNJ3BCgA31bGZ0KR7d
fcdY3dXf6cDI8p3jc5z1DSpGO0eI+T7DG7YdLaABPARhTrT4Uxv61+RPlLRlq7Fy
aWNX8FEoFJLTTFaWAEx6s5nxejEANSVu6nA467yop2Lhe/yxnQsfzYHCeuTfWhU6
cEQjoXoYf83KftnrCHf1b6zu/X34AP0U3TjpYh7ZPUpiS+4VpEldEQUtROCfHHoB
t8TvxpSHwLlfRIYDLQ6v/UvcQQTrNgd1N81rGf7xwRmjO4QhUoqWSiEfXIJu43K7
n5msq9ml0wMZej+WT06e+YxokKUTKuF4HCpQYvpT7fjeXFRn2ydAG54RZKA6Gy21
1GZxqS/kBrKFz4TYGAMxyLQi5oJUbXJ+g2LgFYfvfT8gMqc53dE9HLt8K9i4DMyl
2jtAaN2nb15bxjSzNSrCHJxsSnfBZh8gXeySgfLlEQUr2cZnwomwTgS6z6T+txck
9E0/ftPyHZ5Y+7nkYHkw5M8ukclxXlsq4aezVDaRo4SKTOGPkLKF0TbWbw68XRSF
fRi3M3gcKD6ngH5Qa1X0nuU5ZEdlJCvJgN0FVazS0O2Gj6TtZNaUGiEzzwM1jQwx
XG3pKcLfz+CWFlMSYqdizpGO6OnBMsnKjJdPy3j7W6L4oqHUFvkHfeMgKFeH4ep6
QXjQGUBuswhUDYCONEUqZf+8kX5dPrpIDUCBXWW63Dy2t3U95xBDukcPdX99M18a
ewPFAD1p7MNKppyLeMsAc3K2HrFclWvRsO3X3xcFFDfUYOho2+WdjeCbB8og9ydF
kPmlqPoUReJuu1sNV2L3JE74HkGkXmuanFdvI2omcVHhFqMCXu8U8R1eQrrRwlOA
FCcxkTQ+7+jWokz+ZsbXVfZl/g9ieZWfi8lLV3mMi9b8yX9OQAl7fcF6FLPd8CMn
jtQY1PM5zKhe3wwOVIYvZkCmiwKmYbPYCDXdjuDtaExyUFbpDocicoWAPykxszZ+
WUJk8nfGLjP93a/4WPzJxmInRO0GpeCRA/UPoMXX31PXzD0bLe9OOgvqCEz0uYkA
tS3DqzGzYlW469N7KAsa0w+JwmXiPVmzewCCwLap6ZdRDg5EZ2LDUS5jYv+2jOwA
Dr7hAGG2Oe9DGixQxxhhk3RcNt3qQA9VzUMRiwJXN8rQoIWnXQy/Pnw5w/6olqzl
2ot2sPDim+37JBFgTVWt2iLGvetgs49/6Z3JSor4DBUp8h/e/fFcYEtxklS+byzJ
TywfPrq1s1PJLYbEQA6SrBiPOkp0P0gQVu7fLtyqYC7+rnTsVTaT+Z5wG7LzhEbD
ZVLBYWCEmyiGCqlxCUpduQRckccxbyhkxS8wiGuKJoSvbbxKJJYBE4jnw5SGy/eu
4PuFLRTem2KzFWaBjfYhFm6nU1lDnzN/lnci5JC7rFhgS7vTff//g6yliE9Z1XT8
RZErbSsh3mOsoFtmeqaLJsjCepw/0+3gPaDqwXJ8yKsPurkYDPAUREgLanJzoQWo
JJN6bPW+1jvKdrLXmZOLXI+pXC52gsByTpZev/kKe1M++pAL5wUd5u1BIzbdKkEE
LxYoIZrKH/pXzqNNILzqU10HosIJxDcswYzudXGJ+9TClEAwCHIoHUoqa5eO7De6
otDIO1CPJhvqSMjA6sSuMOiOe4V7yMIuL98ZSo19kegbUGyWRnLn/iCuQ3xnFi1q
RLOGO7L2JP4rdqYcvN5hszsuEKJrupxI5kR/kmwGwP6x25esDSc2MhRisSoTuwMk
pFGXNo7i/hVOr2fJNWCRzECgfcKwEP0g38t91JD0PQdaE/cbzmVDY+cu7AMxIf3q
jQbfF751RbadmyGWxfp+v17WH8xYH4B+XKg4aM0H5jluPaUMYQobrzRQjzhI/uEm
X4+bDOyXVAce40NcMq7kWeTg0F3+DByDY9D5EyeLYLEzSQ+e5jWnDeCEYdgIgKXO
UbqA5/e3A8qzUrBK/DgndB3hiKQtMuP5v6f3JM/NNUy1cQxelrCWfrqauORor8dW
ObZH7DYfxakBSnv8G+dM/Yd7OC9+IQUlVmcizU768e/MtW9JDY7RrpB9Nnc9qpyu
GAYOe+0iUnLvvZTLx+cBLlUkMUXrNv6sFJ6lIQirGfjZ1dp91+ri5okHhNLxKt2x
0mpisy2mVTQq7hDgHNtl4T+aJhN88t7a6DVQP6kQh2CX7y5gN8idAFOT6dRxhzfj
gAwyVL/P6UfgRkpcyagM1VY8u+RqZh8huoUwJXqOCcuyp4LRhW4kC/u2XgNLfCSC
ScIsi+SZHY2fEBX3hlZpQEOktSDbw3JSs5l1AK/78Ba4fXeFpw7meI1XBhQkfCeV
/55Q7zo6giT2Wcfwp+qjPJYo+9JCTMrxVZB5jGmEftXKjzzV2WIwEogZsRaQeqSS
TS9FSxukBpSA0Xf8yM89ISwHF7Ql7iggBl8kE52uJTPIAElLRB033X0xvZYSqWAB
1Rd2x8nxrcnIIDjZlwYh1IkLeYSlTQ8igI+Kjcdmf5+lU4EK7uUDf+fIyXeyhm0B
/PnY79pf5Bd6fGAJeOfgJH5XW5KaLNlHJZJs3rJCZ9D0RmRpfcrqlN3ztBK16vWD
ngOVhZgQTtQZGHMFiujBFknze2y/5HJ7+WmIFMSAhRzkN9mTCqnlnPJxx6VDLBFc
noTwxBjZl2RhLayJoENaaMVINdCZYHecXjbX7PshLoPBNnwo+dTwHcPTu83WEIXe
1Ra3KeKhTs0QR2CNYG8CEFtmq+udU4nWrQrSyOxyJ3BhD3d8Om93/Zh1VUxH3rx0
g+T1vgrQ0NQE7MaxJQlz9U04spyPDngDVMmEYur/hHumenu2LQ5yCdktqHT87HoX
w5mH4fijnQNaBtV3oQz1Wunm0LRqIjN4/scFEP4KpBfMEqbkdGJNPi/3LezCmc6X
iF2Da5rp/oGYPV9KrR5mHAJkO+M+d9Gm86g2fxZCYF4weEcr5wrkQGfOlv+qygIW
JRrI/XFMDZtQMwAj+eBaU0UDmCFN2Una/VOyig2EG4qQJqoxGuMEqHBugzZORpYV
n2WMXtPEihzjV9UjDmP8rwgchSX8p2mzyJH/40lrIgPpbdhooYB8Kzhe2c9vP/MH
0GnOJ4WmgXvFQ2l0Z/nXsAf1WY5Q4b1FBMl7z5rJCexL0SDrqeR0kUf8B7rKqB7f
MjD0FaP90iQbvT2sbpuv3DU+uQi/geIXT523crBdN9rYC11O/UVFTPFPnWPGwg50
NWjNxc5vklcbHIepcGtefEiCHmEIMivmo9RC+E9inuKrbOPwxTqJ6zJb3hA1WO8y
i0q1HRH0myfQ/Zr3mHrYaUeWNN91jqC4E5sBcHUmZk2mli7DlwG2BwaSWGwoz1f/
u7umiNgh12OJokwOOxIX2XUD/hdFYuShT86HaX9oJkqVnNci3gpBEYDqZbw0kZlI
Gd7Q58tlIOv3cMFjTDAMEl4KTNkS+mknqBd/JS0KORSqm9qetgazjogmPTnYu3pe
5v60s1ANtIDSlAqWbqNJYo0xUcgAclbwXR4kN/TJO4rVV5uBwr5gTW2q3qggMku6
EMf0YQTaxdl91EL5TzbYuIru6PHk4UfZAM01UlG7yJqzJUSD9YYZUob3eNkFwUkn
jwEZNqoS8+BX3YfOTgC2XZSA6Xzxww4+SbSLrQFccMbHDwwxUMeamC3ly7mNHmE0
QJQv0k4OgNvyNl9Cj7mRTobs746q++BdSORj1qyAKg7XmxgjmxKx91wUJMN3gbyo
6AY7YJO9DAlDVx8asn9eCkrd5Dae1DSITcokKGwONDFeSjzZt+nprzWl4YBiuzO7
x08ixCtLkHgO196MkY9X+1RQymhOAC0eWsZD0Opk9JlSLJa2a4AQ6lY0KZstNjw8
bXeSWrYpnbG3STytycVl1LP55OuVw6LIUFretKAr7+mdU4zRQAHj5k+u7WXmlZed
uTYn68i/gc00BlmDWkyYPMKakLzj/mSwuFImriMyo9LlzvwkbfsI6XK/HJ45RCKN
I8uuhlnRjQRe+GyQpSoOgaM/sreLOp0g9xOK2s4AL38LWaS0WMjVB2MlPCH78Tvu
8rAEaxBDbs0QU35GBPdOso9A67BQ8FVWMFOI3/pGaEyIimwPcLBYfzWP843ixABm
kqrilOFgF642NZfDnWr215DTUgrc4Bk7eIJccTM95zTaaTri3CL1MPwlPjCNGDws
OWAbCqPHH1+PTNq3E0Z/S2NuKRBcIkKuMElf0Ah0LGomAJElYM/ZqO+uCoeuUxAa
PgtWVnXB+NiL15NDgmDorM+GA0/lyZAlrQx4+Avfhp+p5N1BaMqiBTt7WErDcQAM
0cO4t86/+LgB+am06Q7Duf3x9ccxD6BOESvqhN250nYxazGy8bmwuix4SDAULOtQ
2nbLf6w9Y4ujdAI2KXCTig7RQtjpO1I/ygq0EgJ6gRuxARgd5tiLkaadHhiy3Khf
TFRKeXXLqwzUBdAwthRIH6Sunjd453Fv/joExTCExSeH5WLXQSSRj2zvpRac+fnL
k+cFs8RKzdQDSBo0H/wdWf8ekO9NtQwjM3HFozkP1RIUPBkmtp/IANEZx2ETB380
iXM73lPZqJPm8pctrJgKbPwknDTBCeyojQwq7NnNWVc+P5Wikh3uQZhw/GP3xYR1
p1GGOoC0p8BSN4KjauU+LGPXLXSnM3Abd9Ynf+wdVEZ1XJy22t8U98KKbLA8YhCc
4PylpJeBEj0dg15RGR9zGnuiuiNF64Au0WMNKHevkW4hqWY3H13WmwqvEDSHZ6fR
pukWo97YQSRtZJhHqlr7VkcZuGenfTTkXyFH/x4UNEmXtZkvOgfx4IOjS2Tj5wyp
PJqE40pfzKzmHzIRs4+tnKEiN2MG4zjd2tnV13A9kgR+z8jOtXPzxu+2Ng8Jb80i
Xdidre5D4rikQ/2p5cK9PhqgG/ekXpbkxQdkog0INbBtE2a5mjNSGofL4O6GVVYf
5bHwm0h41wL/fQ0zo5bshMgAqzE3+hdqv5Q9vytkc5k=
`protect END_PROTECTED
