`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YcEtSS4dtPcmyfYmAoPmiDMC8HpRXfYaBPSs2E06yUEvuwnV7n89VdtuZRo0FARk
BYNsrmOiypKqUQzltofi2fZ+DQY4YdPKHJE5qsPPb/Lw+CNgkaOWQuUfPzBCyMRj
9BrTUdReJT4LvZQkN7DDMWE/yVDlDfA4tVdgA2IohaMd3s1shzmHe3P7sXwI/nke
pHEUZhSYyxLpMXHjVzeOAJeI0KSHB1eOejK8vMHRPlcnsLhBqlsEMPGLgTpDrKfv
e61LR9Pua+wagz1c506JNtVVJfy67adfR0aIY3oKE+wFP60W63lbWHVTv8DqNgog
J9aeC1ZxCBACl8X+eITS5X1645KcZgsVKEUzM7I9JTj6lIXztpX/0Xx8Yec9zBJ1
WNwmf7CrjfU4yaFvNfx7Doc6Qm+OnecrEJd3mWJDPpQ=
`protect END_PROTECTED
