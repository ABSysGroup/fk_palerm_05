`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ule5TEnVcWEFJmvGzFeJ+aBu2pYa4M3sxMmyqZrLgaozWpl4P/zszdK2d260i4+H
pJiJwDKs0ly+3wxdAvK5OLKWbbJCo4gchGqz9DUuU1gnM+Rkkb7OXB3IX6vVupdp
2s67CH2kyodQcnUUgaqnKUIcazL4VMxakiaNB1Cl9IbmpKfLubOQL8NQG9a68kof
m/dE5jGPzSaq5iZlhZdKnwV5c0Ha8+Jpl43W4RuSZPUri3CR0S9EtSPMbM9WekpL
HkWha8XqEJvEh3Aeu5VSLFjnUp3fLVd8oqOzIsmCJlDhIyCi2a9esPE8GDeGVOXs
Umpj7/nIhkMmSQGJzb9gvm9uKYz4+7nwemyyIHj1cOXaqB18VADgu0o5XyPEr8X5
`protect END_PROTECTED
