`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lb837hNED0k3ohdvl8jG/iugjKcB2Jh1qrle5fL7Vijt+neI0dYm4j+yc/t2REMD
P9/GqtbMiw4piuoe9FREfNij++yzz/Hq6QocjbmFJv7MVfug5LyVJJ+hNY4u9KdA
mGDv3EyMAXxdKbismjb482331uX5i8fZrl9oId99tMas7FgXGfw8YGKi0WjSB47o
azJGNShNjkhph/6flD2caNtSwv1+nZ23UDOpnT9+me3mEUaMg99v6o+hrWa9CNyC
zjFAAZUrzsxu2N2NOHoOXMsu+ti1CJareEhbIyVHmX4ygvab1T8m3zWa0EKM4QHI
yRAdPEAXjJlVrdkAEkLrUOUU9EInvGy3votpZg1iqCQJXYMHmwDhbbDAUXXhkqmp
QcTaY3jlc7Drgag+WSeGMgwvWs0nsjVjPo66SBpFpUR4+QUiN3fgoYQsjn7sK2Wl
9S1wxc2WJsSecqe1/BpnVA==
`protect END_PROTECTED
