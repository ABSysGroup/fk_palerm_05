`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GH9bGzOGwiSCO6iKZ9Vqt+9lxUoKsCBoHKUTqgwUBe0MrU7ziboSgMiN/yJxoDdG
VFbZrbGGGcZXG+uX4IUMXCibU/vZsd5K5gVEdGjw0zVzxP5kWTyKFlyJaI+4D6rl
hm79aOT16YIT5rXJtqWi/KrkCEFKajslEfnlS4LBPEexd3ucQWIQA40IGjyApkt8
OPlssAoBcVK2O0jtVUVCufI7PvgqhPCktk+jQ59HOh4snu6pEep4lYcRC5eMBw77
dTI2ituTXP/l63lDPXFtAsTtPZ4MPQO3wS8ytxsdvt8oI/S/Yk5gqs0dtdlwlX5I
1SL5yOAzmz5Tm7VvzPDJDofJqMk9qNArljFeATAi6dwwf2M2sKr5jGIpg7DcgnsW
ND2knS36/7F2sJxX+gC2lWg/lJp6OQbikdtK9HiH+aBmLD6WX4ZBY0ECs/gBh4yG
5yy7Vg6HWEjcmdcgqA7ow5tB5m4swEQ7T7PhSuAnGkWrMLExrLkOjU2CG+SFG+EF
adOFN9qBL0xU5wmJCdRvFUC0HMamgnq4RUqtREmHPutGerMoHHdBWpc+aNWK0Xha
DdEmwlrwEq4bQ69TDtHu7GGBGY5zIqzA8szKRTW6Jhm6yWGoU5ycd8B/UejsCEMn
sSnFY2rWu89u0Jw5pJTCtMSslwe3lPTUeLYci5mj0HsqXwFiwvY3fhlAmkhb6lFT
0JNBpZ+0F9Ix5nFZB1lnNvw9eBff0l5ea5oSLWhuGFvdtj82KVMdy9aLwTD4Udbv
p2RDzu3t/BGYSJo+i+AjHnxj3SA9HstL8ZFR25TQIHFnw9UnV3oGkzxxQT4cTv5S
d6wYT/tjruNxTj09qRqrYw==
`protect END_PROTECTED
