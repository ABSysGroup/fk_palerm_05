`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oI7w2Gknnwltj6bQ575GB8hxB8761RSuf8kgKoCancla2ogRmUwwcLzNfKNt3ZF3
zy4a1UFskE8zP9mNs18S5SGBmA+QDcv6hxjALUpX8wkanFoBmcT4TtHeKIojG/rK
14pMMVMd3Ig3wRfIA9nPLO2JHESNtSzhCl0t4mMlVpe41crrlJsdEJU4pSkZJjzl
U2tjXLta1LlSgVQt5/rJdk6f4cSumEYJzjqRLeJ0gYVxt7ZmF4PIngqDzsrfVfSV
ICs4mmgSF8i4Y3VKUeuatdh0sNpGIbVJRPAN3ax2by4S2g9GPoqreL5yCSylG9J+
7WdAfxgQbRy2CzlIwOCMknq5RLQtoLt9YXuQ/9b9SfkXlSpWybrWCvRk2C/T4muo
HFtyDRdoPFz+3QAfedW8puMzLvjhqD/09DKsg/Cepi8UKeEiMig3Q98P8s3FUd+H
4uHuxpI1TNha6Jv2+hGvfSqioPvOi31xumaAP/ppLJmqT5W+IcZM0YO/UKpmIq/Q
Ao4SHvraiKNb0Jz2sAIn5R1XR7CRnGFYzPEa9OhwjN3xt8jNeIlG9PIVQcZAj4Dy
`protect END_PROTECTED
