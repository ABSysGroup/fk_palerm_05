`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DxAZWXv6bNfANdPfBlSNFEaWCRJQ+F5W3hXEiC5oW2DyhOYGg01hx/6XAMyCOoAj
4NGGQvby2bMlxQl5ap1hdjlPmIpl3lrLm5m5us8mHpwMjnL7V+cqhT3StLTT2e9m
RvS+/MHPHYrChj2HQ2XQin8ANMuuTXcp4Y4oTXMpKr0WYs90gYa5iMugtKCXyyPC
Oqm28IFIJf4ZippC1AUPTnB/vGNo6wABgQJ2BLTlmDogDFESU09vmMJfvEJVgGsW
oinq0LRo95DRNQ3u6Fha3F7glXd0s6s0c67O5BMaJrW856lL3P3SoVtwvHb92Onu
OmcpbJl2uLzT0K7HTEJouTfCve3BJ8gkDxRy3scHWs3XXdfbFA/wEcoJ5S/y4osV
0ARWa/TW0zBTy+hefxS3+5vkFZkloTyY7r7zcygQERILeD4xbrxxHRwxP4GfvE6B
+SBEc4yPL8suv8tQHhG60ZXol4GFi5VlIN6d85qV1TsmHl6xO4wwGGoqEFadSm9V
yDdc1i+uQR5BEGHqnzM5RO4XqR8alViMVidWQRKZpRJpPhdvVtOUEmqVjrMeDLET
TCi+SrRh9c2jWu0nRH/7CvmMRzsjmu7N91KANHNemVgepZYeu1YCSQDUznkwqyiM
+TVcZKU3rghGuKYKHJR6kAL0CBxZIAYaU/M3ucHrjJII5SwPqnDJgMRByQDLL5Ni
C+B0VUooNCrOBttjk49+NXqE0JI8wvFUOkJrPmnF2Nl5tAPcDMguSL2yFGEjyXRU
SpuVvpb/Iu0Uezr0/7GkSw==
`protect END_PROTECTED
