`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MenOLwkh8eG4TAfhKLeVzFsEykZbc+z+QPbUdOOXNOlBRCUCcJ4HJ2k/iH7qwMri
N8phPZyivs672pjNcSyn7JRiKZoBgHNUM+QPOdrZi9VFsnBjWglJxCrXA9gJgUn9
ERbxFAePV/b9VbYRpX61J5UtcO0kpOmpa8dOSCOTatf3sbdFsfMMIdDOY5ebQwAS
Edyb/PXmgO8vTPlPvrOipgpSwXBgW9of6gwE+lEtQzimpWjna2nEV0CKj92OG34L
y4JSLgvqo7j+RCF0CONH7vc55uUgWU7JA7bdDkJHjTNDa7ivJ0C1MhYf/xNb2/PE
4Ii9TA8JrRSbfettAlXbzxhs9r/XmtwZjY3biSGxS3jyOUJq3OJWI0d67XHr77gv
EPhGP8STlwUbK7rUgHy7z6gl7bH9pnf3iBvKaRUCdtU5DKE3r4TVyVOnz0S6nGQl
E60g9uobfSrWijgnLMW4rQqJxw5iMu5tSdyir+8kmS5P9WiABUbGNfoo6pt3gpGS
3ixGEOgq3/aKXckFjZFfzPgYUBkyxtawFtdjDyJqjtt8W7zNb3PhpXUbKXJkTOAf
6LFKTvrfB224x0nK48wpSoli8XEqlaoAO4n1+L2MxVtt0EGWdUh4L7nh86ED7YK3
CtqgLtvrkPkefwey1KaFvd8FAmJT/c9rO4KVwI3SCK3WhvZEptS3oHJKUZF95TJL
/+B/V9CUQ7kt/HOwvflg3eZHZtIJrluyEgKHlVz309bUkn0zM/HnayJNEaountmC
IETFpJsJJIZ++l9IY9EfswOyLek1zLyLISAaCrDfjAx5imOhYK9dsQZVSran9nyI
`protect END_PROTECTED
