`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fIkQzo0HJX6qFrPZDSGbCc0iNWjHKyDTmZFr1qyLhCeGIkcIHQb9CKyntxKdmW2X
DkXTVXDHUFfikPwfmsVSqm5YQYq6KqbPJoFctK9DMEUsOTUfzOQKThN8LZ+cM0mL
U6vrtcvZCDY6+jVa+1cPCVU+js+tYGIwSBbnWcK96AWtbzrzMEfJ7oX5Lw6no8bx
HM33iccpOnE1DJqPcLMDT2HuFRi6dNXlok9unijd+kT93dr9gseWzo9m95aQq7ke
Gf1DPNkfCKHkZUXUq5xRoxwdGCtW0prC8B++oMoB/7jfMay/+CIEEyN/u+VBohJ5
O2+ig1iE8arTo4suLZx8r+7+VGjesHsqte0AnVLPK5HLcy7cEqnUpjR/o+P86oid
1wGiDWbqX4YZOLyBERJJ5WAPFbTKRf2SMAr38uRAsDLCfREg+A9zARUvtLctIBjv
`protect END_PROTECTED
