`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MtF1tzIqMVNcmO7+D2nwTt41OIAU0gT/8TeY/+pD2h/oAsG7uj38U5POfPOuLxd3
Tq9KfBuJ9/mihGYqM4SQG596ncvwZwTz04L+BiM08+NpKqr/o+Lgyc7f4PM+LuG3
MmBZRR7BIGBboWbEL+hf06KGMLl0IntHiHsj24s6tEYbfeLcbXts+M1np0xDbMdd
bbeBUx+bhC06XN69js/FxYH1GbHdlzR5WhJonkAEOGOOKWCEg8T+1eBktDHTHsEO
/g2BZYyRTOpvI1/qFgjRu9QA7gK/QEE+jU8OHSgmnqZQaOcJ8a/h8JGRmXjW64LU
SqFKOA6iCsAPPPQDdT9NncS4sPoOwET0JYSWVcl7RH0SSbDKboOX7/5ALT3b/CgV
s15yH/2qIYt2EN0nPthCkNQebozmIqWsJ/mArkIJgbvySn1hVr44aJlu2KEvXBge
SRv3PCU9MIEhTV1cpO+XmGCgcnVI5AZxhEpniZXe7z5YzTsm11jpxu7ppen0vOdt
`protect END_PROTECTED
