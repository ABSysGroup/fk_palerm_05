`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eDC7SnYKSbvkWeIuWv+8PFm3DZb6aggzMSXP6dWjnC7/wezib4/Pg7CKbczwHXFN
iKYeONBXFUWv+UYAVb4dfs4GWdlMQ3nJdiDE/zzO/IoiPclwsAHfGdz6WYiQIhi0
wPjnYIBMuLRM7jj3feE5BZP6iK3G08oPtQ/eTvWkordQ8U2I9vwsxiFOKllm68iI
lRkJj6lyYvccM/wZGxS9TNBOtimlmNgpnNYSJu387JwagUViXv1ywmEuZz+9AKvO
M9OaZakjgkQyAcjkOG5DKA==
`protect END_PROTECTED
