`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vu91o3uGIx2dgMYfAPOew2oUeYUAN4E6moVSLYPm0a11Mb+Zi2gUISDlKHPOVjL6
dwOx6K0U2vTNa9J4w/NjabP+0BZ/m1HcHf0Uw+cTa0g/TCFqGFVZq/7n24+hjfuR
f2Nr884W15N624sB4UghZsfprD9WYUcO4tl+sfL/Erto8xPaWvdO55mPVZPyVai2
qI0B8KwK7oMzEBsMYrIGqLUoKTyAr3Q03wMfuh+KKbRWd8xusG1SD3dDDg27NfOf
ZdSBBVIDhD5dcVD3OUH8vvzFLdOrnsyV+ej30OJc3wHSX9TRu6vA+DfPsVNrjE3x
dh+0Yhe2GHssPDky9f0oaPh+ZWeBu5ysFXxRRuckqiA+9aZf+PNWnwHjVHJ5upqk
OEOHe4GskDbkYpi/Sy6Cy4eznY362/WHYwVtaJB7b4TMb1oR6XIFKJDlEITDmAjr
xd/G4pwHHudAg56FkvRrHGmd2JJ5xDk/9SynhowcXkMofJOMA39YNe3LpieEL1By
MNNOK/rq2Cwtg0cBAW3xnn6JRnd8CFF9teZJEkrq0Y8bJFAS1YYO9g0spw9AOB55
Jo4Pqwx8LkvrFmDnivk6oPF/MFbPqg9DCO7IWjx4JcN0BK1Fbe2hWcB41eK0IK76
Zi3V8eI1xXwRFnJtziYJbUq67XMxtrPUDKRy8P13I39NiLFSEXKLr7HqI0MslYyc
6R3cQpjzdDNzAQ0NJdwiO+/AjQfPNUuKoyvmJxIUMgzt88we03WCJJ+ogryv0o5u
bhAO1bKdvSkaUIXkSF6bf3jCWZelejm1Jp9KAiNPT/pdgrmLvvEiDjHhYpVxUFai
2jNr+LUrSq8anKQSZMUuwvvlUm2pK1GR6WgA/covKEr6er+rkmMC+9EZJgF/Md3W
Aq6bthB3DnF6jIVSX8k2xiWosPgIdrnevMaNvXSxPbOkNPI6s/7IX7EKHZuT8kLe
gdfZRLTyItiMVAbZs9R/t/m9vqesqajJ944WH8jC29V43n8MRte3jR3fcOli5hwO
392eDsQbKJsnh0+CnazxZhYlOX6rsy/tfQGfGre4mrM6JRaqYaTN6vUYCUb5fH2F
2uBf2UQjScFqrITFAQGSOkn2zRbupGlg8vM9vqMd/Q1WBQzpi3NEh5Zdj4J6YT/D
Vm+rJAhtwFWuZ7VIsQXZTyp4TD4VH4nFzJAejREH2ern1Znaup8qJjxoHfPhUe9R
fWcsmxXULfzX5BFWrHSg/c+mVGmDeY/qnNgTCU1QOvGfNZdjU5/rPw2OI5M342nx
eqfZT18/hvTNunu4bd9BfZr2+K2aYuykwzZ2KGbgNotw9uUu1vzV6vZQnfmlDRpk
x3kwe79P8/2Xgg+2cJMgg5Y9jIx6AiFfniM3MoyRcJf2v3ncSpGbLA6qDXA/lPub
xS8HdWiY55QegNBVs5ApzrGQdFAKtvnKBIy5kBn3RXAGtypsDOhcUiKX2/8WbleF
xFPcXrWcJsrgtZaUsOGnQFBHZXeaCupToUdN5sP/VUHDhYfJH0fQfMyjNQTy6ye1
H7UjfbQBZAkqQ8ljORkvfgRjWFmPD5HUlqia4CyEhfzswFb/skuNBIcUPTNOJtrX
Y/WtEu6L7TToItkUT8euCgvMbHXE6vS+w9JibV5ci3JtJaT42TNav+ZeVihdzF5G
H5bcN4gMz9XAC4a6fPZtzFgEYperXg73gDbDCuEiw5QBYVYURLVrCnp9y2ke5qTO
e7KtSeH9xa965x/3+BEpsysMrohjpXfEzLRbzhyveakI8a6ybVXNo4WPr77otzqI
+jcri5aRKX15WSlp7g5wWyiE23HW0UY4U0TGcnCsLOmjVPm0eYT99sUOb8NQRN8s
Ue6pITsS9kJnkeSmzlaoXgEIMYfZGCiJ9XDBLU0jqQNRXFYR3E3Tk49uQ+6PmE/V
bAGJsHzE+gw2m6gmvKhSMre67oERYDEZc8/th+s6KZ41K3YOryNAAR5Uj2b1tLnL
28kNWheOTvR1i2RtBqHz+lZAOZQdnB4z1vNLW2Bf48KSVp3d+tXbAmrGX4Qc10KZ
lJOdaSP1LU+umm/KxqoOA+S4w/CzHN9jkgX43KPbtuuWOqB02lrLAkRUX7UaIQoF
VWemta0Q3MzHN6aoCbACTEDVm0Wb9pP9XHCayWCrfNQUqkvs8rWc1eL2C97djpP2
uLk2vfj8ODRCODvIhUUHy9mlpAEm4mZwqb1J3KJx76UG70+RkCMuctUJnMLhpFQ8
e+g/YqEAeVPhSIDYa7jiVuZG36fW8W6u2d8hv9L75lNeDbF9vvM9fKgJXZXDjzbZ
FyD9PrMrWHdREL2FAwT9IzVLyA9QNKj4OIGkp5BPI6GE5+q3ZyqvgwW+VS36TNEj
zSTO1FftGly/N6Q+GflDiBFKo96pplM60PR+CCqgW56/BHmS3EBS2rNDO78MOFMI
crf+7+OUs4HEHZgUpXUuwGXelTsVH3tR1fDeixF7KUV+oIEYXNX1cOxfRvDYsgXN
04EPUaJUXKkFDPpZGGBrsLCFa1rsw/dF+EEZ5WABv8DmKQj6CR4FqMBVCR6mxd13
yzhYhYIRhkuoz/ZN65HiDBUmWG5SP2Nexb2B0e9IzvJ6BGDCmvYQ0YsKjvMwZ3Ze
JUKrWsEFI8lct+oVdCXkcjyAhpEOWQN1uGFwCIPfbCU/gulqDz4glyOp6JmKcpNo
1swyllf23ULyVZomttd+QQl/QblEWS2LzJsZIGqNu5TdNW1sqU3jMgPnqtY1T6S1
CoRM6HbPVW0kkrqr2wns3eFGCu/DQMYiN5sj43BmU83QebBTeOyB9CGUtcJ6Hn15
3DeRUnxvCIeKsZ7C2TeOvTTfjoE3ncNojpiAX91y7njrBp9PBCFeBDyp7YJy/nP8
cMYEy/hdVonZa5RXzRYoDiDZUhXCmUr7xJwKFIObfVqFG5tY05teet5mWdY0ouUt
baUZFoGnQDYF2sQ2VtVdMdCev82vKLnaxWKiDyEO7iecyIrklGZfC9fuSQh0wyYZ
XcmZ/L88FUiSxswJaC0NWTk5DUXJBlFebBENX1LmsrPT+iCXfa04lXkFbsQuNvE3
5Gg9mf8Am2uQxcznez+iy+UqF7ZdpStbr/0JofXkVCezEu60L5vZeDWjf/cI9eLI
7px9mPWgmAnTPT7Z7X68HhqYQp5Tn6KKpUo4Gs11T1kPpSJdb3eeWsy1UqAjZ9qj
Xupi3VfzrBKML2bllFXHQsQ0n4AbWzlofWWo953nyLdn3i8r4ljehdBhUMps2ICx
/8Imunbu3wAcm4BkU+VHLu267zcEIV4g/ZwBKV1Ky6jr44VSel7azLh6wO1mWyxv
eNoq24a8IDd5FkcdXXWzuWzExYiLiCjr+edCbyLaUiZxLS/HencA7VDzok/kCpcG
ACWQFnmIVDm9iU1XVWXHlqAJ11wG3v3lpVcixOORV8XH6Vqgi0VoBE+JbM0J2Dr/
3osWYMa7fM80/aiIksZGqhqejZSOf/5cHSAxRU3woIlH68lKG8/fUhvyaQuTltXd
mduG3tFO5BWgCZg4NjX7K+XMq0gmoqm3ZLU/8psQqohMzkrkUMND7lpKAJietCQ4
u5vyry/MRyjXp6Wh7w7l+m+DYJA6vcLijMPXJ7fdDeSdiUWjVpU30T9y0mVYzMvW
DKPOn3jx2lPefFcy8PIV41DJyqcfuhYonGv4hjywbFt6rKZLGC/+WZ73wDXVcQTN
xvTDdL+1jg7nuNLSrp2nNpy+iFNx0Q1iMKlkOTLSNZIs9bjV6+IMXp/uu4ymCNji
uyjBsFyBP/t5yKeQPxvCKxM3yLKowtsILwK/cMPBOpH/RxrYdthf9c5XySBOIuR5
AlBsQaWtErN30RAp62jjV0SsowuBmnaUtguNmOiKiWBgrqTlQiKCVCrllLQNdzcF
tcNPRg3jS24/HozKSzadKTOMTHKMZrKiXakZmVDD1CpnOEavbMEuFudA9vFFlOX3
H8cRIJ4zz0OxbT9ZI5PIE4DRfdcVmQ4vCWOdlZJJMFpyLgI3WYpdMwys0t/LfRro
QC0GYPdx3y9S+5zMVlXUhAqa1RYSvYMoL5Ty+h7sD7FIz9o/CbELa1WBEB3iF6ry
dNRNc/9+2OJRUADu1wmDEdISJkyEVGlofuouXhOmpCVbtCGZqlcXF7SPHwnI3MTn
ZcCS8+8jLRKv22jlNEww+YwRBtxMm4YdoMVvLw//5CeSZfgQxuBAOKFAmLcqBwZK
FK+lEuJVQDaxV5BY0br7HaYKIQUOxZHKPWQyu/oAGk1l+rtptzPNljSaVLopBE50
YRL8CLJn4GxGpTWt9HawiVvzwbyyJ3eXoUbaZF34fQTvh1zZ47gSFPu938NgtHKy
uH+uXVbecBneeU1POmAuE8iCms65jC3S53KMAxcoNrgoUIeisgPsaRq7h1YlQwWB
S55ttEQANQB3LLGS9zhvrJmUbNXIT/IsoOKAuzTLKlcPjeUIwqVaOThy/8JxtVlF
HYsRSry//+fqLgegsVR9lhzgXe91EQvVUvq8JpLTkBMA0H9KIeigw4PxQAyupb5m
B5c6klIJhUKQTYxuEg9SqX2O+LAZcGJJa2ROaaHUBiFm+zZF2/+0EZ92sO8WOyWU
s9OcM5SGWNjQjYEM3nvfJoXHUJrQQ6adw8m2elJVI1nLB6vhv+n+b2zffXJ0sx3H
SlnSK0a8Ad2DFkXO/LzFTbPZFGN6nc3RJg3p6ll789AQorRAm7KFOyUz6PLg/ilw
soHonJ3YORqRvsAh3Zhad9OnBacAC3sQl3Q99X/1Hsfb9i8HbxB69Fz8rs6NoTCk
xmwYkhf85RL6d2xHiTS/RfbfYAuLIk+/SLcXceZa5e72WRkl8BnF4IB5eId1Oyf1
qk3AJnwN+o+cP0cJhSWZesq+h5vXhW+QOTTp4iwOPJRIGEhF+4STYLkxBPvYCNm6
hlghr6N9AstkpP/X5vAI4DLuEiJ0/M/6POwxShvk4BrMgcTSMjdHsA2gjp+EDzj6
AQI8qQrQ0CNXuoJD18cLx3Fhdw1JDGmQ/6fo/jXzq1QO0F/Teoudw8Hk2yFMIFq3
lJbOb5AFerZZ/NBfK6eod/pu+XL4qscOA7ix9LQMzUiauIWhdfXaIQrXhQ8KN2nG
LS7B2GDcYiFfeJZwpdP2wYfUjjQNSsYf9vPP7KZ1QmEJyeLWJQFNI+lN3CYUR9zj
mqCrs58g1KBPPOQ3YuRiMQ2mqjTwnMER8PXBXQbVuNPAgT8n0NRFvdD1fsBGCI6K
FN2gCU8Co0VO3kan8PnhTcc/c5iSoEdLEB8/nDJKFfmGfwB0oQxCcOf4jvaxTfMY
bjKXeRc7Vrr+j1v9jDAdSQ+5Ku5VcZEHYXmCXxwptJJs9Yn6j9NVOJVAI0c53l+y
Z1K4I6Fdo92lDnCG/ISdHHfRiBfWpP/XEbLnpmjtbvsyuw7VBHym+8pZlDHqhNEi
NCKh1i6na8Y8bMnkYXWH8KYulmjV5daY1USKVHnTkof8rBMBg+kDiKuTZ2KzOqtH
0Lca5KiqO9R9JRtl1y+EpuPCuLZ7xjjtFZPCr/x6otFwXiHGtpcgBCf8I+85MNbn
jvjVubs8S5DgasDZiRlkuGWGmHIhxfK6BTk58ycur+gSBplSTAIqlDp4sIHSUVlj
GtgCkXw93Dc0hqbGE1C93ZU64IUTrmuq6rFM+sgYPGqF8ZuqMm3xJP78V5osehXH
/LDCWXi1ol75bJlP0ipqrmtvSwS9Rqk9xk/+vldBrDuerVM1R8W5kHJ8GZGTRUg/
/rhhzf35BCeCcpliKk/hUM73z6LXhl/lvW3jZQofPI4CdK6gZLjlvYS8WiWBpnL4
mTRzmjgiVYo7yy9KC5Sw1O6HZo3x/Kb5j7jeSc0Nn7T8BatLjUi9Ht+HTBH359o8
5QY2vJqd1qKHEKX1NNM3KYsnxnsxF9N2gvueLh1DeUhohzoQLhoC1MuFq7Ao1VQR
v+Jv0r64/iXjrXrTWyY6VqVJCjgdpZu2iOtnewqe7dsEHlB2SO/WTDvR/C+UU6fY
zGC9ibT+gIFMzrgVFXtYUpzZUFUHg3oCj/eKTLDNw52O8ms3uuH0VDHcHXdtah91
cmMhN3hTwCj2a1aWQSMaHlzbZ59MTcFaMAEINVWtWB7F6Pohe351KORmQ/5y2uAc
zkw2aZQTm9INPiV6Z5XivAWmbT6iOg9nmFBU5Gls/9847VV0+jlvfwXyPJFJwR6m
l6wO55ych35PnMgYcbiQ6tnK/DoTk7ro2YYVdrS9/bObcNrJWrwnhjLyWo547fMp
kX76hxkQSVu53kJXjR606GxJcFi1HfWU9kIuLIwmFcylEDi359tMDIQvto6eImvv
iAnpEaNFT16G2iCRQMwojIXFcy2gqs9T+BT/SFkSKLaWAJcbXFqmncCc6lHL+c2p
i7fxgVl2qVw5Iw9kVfHatViraFnOOnM7/vUiMfiFbXl9bn0umsQm7N1PtubH4vHT
p1MM2Jnxhy//SYgrWOphpEXHgKlxZDQGfQbkiDgiYnrYHuaBqakrmXfo1i+0TSHE
ZawFNk0piR1K/aupZhbTKbGgbJUXLMkY6S9H0PfxWva6PewjXRD1O+t0LUw5Mk3Y
UR84J+d6eRts+v1Pj1FjwMdN5QuzrgXeTrZQ1RQz6u1UpZElpq7uhoPxEd1lJQcx
ndGu2poddEsuPNY7blDtNlkgti+qTJd8Hz8PibFUXeeKF1XaPT/86mo/Dixfuic/
pSazwYH88PNZnxBwdV5cdaeGsDGKVNkplD0gJBvZB72Hf2kA8h974Ayj8MUhkUy3
AUvPiUH9hu4G0cb6oNfM+ltNrE2TvcnO9zF9OBzhfeWh/jOj09Gz5jM+RBIOv/bM
S90v6Ia/fbIF8RIbwdhC+H548rjmsoRDqK3Gq6gypPJB5YzUI7yzyimOlSVxLHB8
2jnTm4zT8Q1UcN+fNLR6Y8wqOY7fBaDqbBPXRUJ1W91hegxbANdPjEgs16jx7tOu
zwlIZ3lCvnUg5lt7JtE2HKHjaEvx578AcAp+PMavyxPu21jDUxAaEAckKG7XBmms
Xo5rWIlIvJdwCmtjGOdJw4JZfcTXdPro9kGWY0CDnIoaQ/KKlUWeiqQdd9MXSJTd
SxYmSR4tk78QGyRizsY6/F7UtV7xE5uI3ERoxN5ou0BKWPvT21uN3VEe99setYFg
/98KuNDsSHWNIj1fQD7pCcs2myKI4AP4CRvPdtSa1wfKFvuDWzUn6NCkwfbqhsx0
XLioortLUvEkR1ybAzAFzLyN+5dgVn46BOLn7SGz5DVXOym1Scrn2NWZCeVt6Ffs
kE/G9SHnraCXpeh19vnWd3/2NNA2YrNsYKrOLE5nEnKM2eINmKRDCRau98KfpGMH
Tfrmsn3e1zp8kptj/wSIAZ9NSIsYfeJGXTzP12p9ucKp8HbqMPfZQRCDRFPI0XdC
CYpof7fO9w1Xka/wMV129Fv16MlhJlTt3AJmI9JyQjDX3Uj9xaHDDZl88RXVkElK
Sto3PqshED4b446xXqxu5qdkFXgkeqwpmmnb1LDgpHZ4FexM/C9WFNk2o+dadXad
8GkZ3pR7LRl0lKZILyMSBGhAvKv1HFhuhJpYZvcIWT+OlodAsLH3vBPxTTIYG0R/
IU22IkbJ86XXByF/WToLP62Hqteazno9LZUPBzIRroAW7Oj1DWuRau9JwYNjKLiR
+lFoIfGngvOmIk5bo7+dQ0g93gcOdMaLgYzJJ465WpqDB//HusBy1GZrHvfGlCqt
30XthzVm50LZzRNykZFxiMNjAWrg5oX0W5TSDikEyDzQY03Sr8fb77/4w+fuMBw+
FnivJG4b5Eiz+y3gmUZoBRvwTd2Qjd/Mmk8GiNNglcYNjhtXvbRLzIZmyia5EtHd
M7dMce61zbZPytECWXAdNuz8s+NkwoVZvNzFdjvBoccoDy7kWP0A/jKD5UVfu3Ve
kHUmgkBETsFaPN1hVKFdatVnESyC9pwgq39JoaYSw1m1ReBg4jjgpqFzApqy1xxh
1andsbaFkg4SduIVX6s54oxaNdevDvraWfOpCZFHzy7t+c0KCB0HmXXuBdfTEUGL
1nEGtuk5Bs9OciGZoRYo1OYFebRgL1jdPvgaJ6UKmQpkoFNXXzVXn0k5fYVZtrMs
hyeyaGkUqPR1Xzdv5L15dlrzmhlMTvwA/V37JXud8T7PHw46xwEOGpV0T1kkyELM
WRoT1cRspfsXOCuxqQSjuZmVSyuTKF86uw+QORKNhcHcLvoCfhJ8OnaEat1sIkwK
tHq3bIcEhoN8aacadJZCU315T7dGwZTBpXfY/9xbg+n4tVu9jMTlJKIcbp7HZvvL
+0ZCc6CPemBnQBpAXtsJa3IFlgCDIAy0kkRJeCw68QFkR0jmIEx8YOwPpdTNA0Ov
kTYIbBs4fdSoCcjvp9pNWJlSYYPwymAFVi13WZ0SDSdiGXzvAXrLbgfmKtWiwjuu
uX1rIkMMAh1gxNXrAh6FN5D6IAcPSwsziN4d+xXuhbAD+RkUWmjPBiELK+117dpx
eYKGUrYNATL+ATkpwe+U/7LxlqLf4J9xZ4QPPNF1vonOcxvNHuJBqVgSRCK7TrSz
xTUnOvgCsrUkba2vRLMeSFpWUYA9nAf1mvJj4z79hGN9MJmS9qYw7R/IpxpiF0EI
zlZFobnHPisqoEwyiK6HNWH8Jdj1gi6H0EZWdZLW5n3P4KPURnp/JUhzDRkuMnvM
k/vcPeKwqEdPJGsirOsQChAzedqUeqABqEblg5yXICHvuPEyuYwz1EYrfcwPxt0c
36/jj8LOsRX0qtQBBtVZHfGFLmwHb+uZY5o8p1Z1zTCvc1Pcfes2hyWDlvYT7JR5
KzKrxp7hVK+C7LTnjrqqZd2gxZvFsxT80oqDVtmiwjDOAPJ3q0zhdK7DZPsg8aTX
ImtUuwIClapo5UHkQ27JJUE5sh5tquw2VmR0429rVpSnqJOtmxplkloLSI+0qN6c
5aH36Kutgl8TKeqjNILpqD+HlBQP0g2ml626mlNzBNNmf8Tn3/E4MwGyGyRJyZVB
4v5qznLqnu2O/iq5KhSv02VsgSbVSoafaNfxzwG/yw+vcCEjlh2dTVsAfzHJzpXZ
UTyi2HO4gIaKD8/6xxoBzEqrBTSY6T8RiqzfLuKWGUvxDubS3ZumlWJNdyeQIgIn
deEXMl56JYzgPMEevXByE9HnqFOOOrBJL71fUBxjwPPPkscYBYpBAlT2jLfyUIVu
ZDhg+Ie7yGbM8fkJbrFqC39uOdrYA4DDlfXL686M32PHeeT07OhkhauAuJ5WjHlF
Xzdwk4Vzlac8nw2wPpPr1wFMyYNYAVF7n0a+wPHobb9Ggdpc+bC5IWNGdR+GiXtv
p1rtq9LNlGFxLD7x4OXAoWr2c9782KBDn9zeo0GD5j61aNJmFecbekZrbA6cRRLd
aEif3dX5xfvWgWitpn0dSsJU2924Q9C3aeGfcnE7yVZM66DLDrB9XovJ/lFriBiu
OJEjnh3ZHCOBr4rBDgjv9rtd8+Y4ouQQulyNEr6Rwy7GIsKkM0tc8C5JZfvmhKCq
sHJfn3TWL1rYOsqwnB6giMv8n62FJ4JfvKgeMykJbfODjiGT7J8gN4f8PvxhkAxZ
UDMlzv04cDhYZihmsfNLGMCWsLeHBDjeK9BC7uk23+1px/2QT7ULWp1AniwkLt8G
E9A/dHIjlmry39LQB2ET+9m3R+7SkPXI8OUptagc3lc8D+EpA39SkKPBvn6g9Wnj
TBfX8Kpr3x3i8IwdmX40bihlAg8mCubajQPBSgDuGMpdvp64SCfUg4fA2LGOLBPS
26otgcrFhjlQ5/qJmIxTduLyU3Ere+NLaCfgBq6KH4ilGpJdB4+ngzc4i8BHy5t2
A1NxYpBGyyvbPwrdaHErmGYAP7OMQQomEESo1l3b5t7O+S1AUvo+WgCa47SV9Zd5
YX2kQFMynvvntRRy3/qBzQAOjqnjeeIe9D7pSYamrzLCm5jmOZUlI3JdYtwWAW/v
oSXdhkFEf4dYKpG8gmn3ph2Vh8SPILfEeLzAgdegluUcuwsMiS1zCHQ/CRic2C0q
/KVjdO0IZ2t6ro7aq48V3s1dsaEtUuuxS0DT0n0YzhFyHZjohpw5gtEue3TM/ZSk
MmlA6pSpz+uyhoqAYV8sqRU8kgmNVv6fXpVOBHQRRAGYGGbAyiNgxIYuAfWB+Ub7
WIAm6JxQ/JPU8A6L6CQYNNTQeW9YvpjqnWjGo5jFYLxs//aQbkEulPk/3snNhh95
KqOEftDGY2bTY+m7r/wmuiobXQdwCp5dX7xbn2nM6s+pmzGdNbN3g8GyakNI8mXS
UrsEe62Ud8p4OFiqFkXhWFJMRsVTWGC8QE6U9jLwwXyQ28eeGqVhCuwIHSXpNztE
/Wuqr3Iop/DJjJDoDaEnXIVugYD5rpXRoreMxBvz+rCnOs+3E7ykk1C81UO69QT+
xb8QQIWGRTb4P76xEKxgaFH8jXvUVPIvbRjzUPDTGVNk98zLt8cYVKD8hzRhHfIC
SqTTiq1AhC1bSH/J7i36HZ9AuQBwNF3R2sQR09g1AkKEpF2FLK1+3y73gqFxf2To
K+zd86yA2PsY3TO9NK6+P9gN0MrxtWMgYgBMqXoxhZrKH3GVkJ09goHxvu2sb1Mi
GQQ+R0FfSsuB+V3MBbrCmyeBVs5ngnN8vx+aCv+iBW8YzcNXM2noVF4pGUVgD90i
M93JzsbSU/vIIPFtlKPqa/DzLEFc3Tj+eZqTKQcF51BAYzNWJk1SNEoDttApTu0L
ASR5sYqTp9zqgENouWYcoHVOkNgVij8p18GZIwP6AVUkpR5yFtl74B/VfuY1S4Py
ijP4rpd249qrx+7OASs/jxr715mm0t1atEBsl5KvjxGFJINMrXrK4V1bxPcnS8KA
ooRukAP5NBAelLLki9Fh+Zonm6+E4mB+0Scrfn1wEihXOk8vy5tGGZAOaDxcTAbU
K/EfeZsEcB5iE2aFYOyXa2CG+3B7dhivlCZDOqgbsZOIcHziqKkEX4C3rNcc8oyt
hFEyKG2/w+CMifhqRHg9edVTe2PhW4GY8aOdWLNmKYY2OXBdhvSKAK7w51A8ERQC
2rFzDIu7aWKMKy6BlAfk/kK8E4lnB1LqSniScqfKL4jL0zyLyaDX+JVNB6Rw16+8
9SKRcgMn2NvUw06QCPzqohHtw5N8SQTXE3SI8/M3x2uqrCtsq2YcQPokQpczGrVm
lTBERvFo+n+g1gbKSD3oVvJFs+fqdx4pisZW1xYW/3Zsv+1TKBM8DPovVuQvxvbp
M77Cm9Lc8BNt5KTiuriopkwAzx4ysdoKISzSkhqKJY8X05PEFHiTz1XEqus76m2h
Ewy8HW+QLhfhyvUz3xNopqvbBX79hfzpDbHBedgZgwKN1Tl9fg2PcyAQVlVyw3in
/cJIfoRlIB/YANpMRMfBALpFL/9N1UoN9m08RjThNK6uOubFNgq/LYJEVED/56cX
jQ7afdBt+J8I0reVkqrIt6bKnbcr9FDxehF3+5zHsRsQ79fqTk35p82yeh7/mEfi
seZg7vrI+tSbAtb104V1EmWJHNlf1v2chyXI/yFu12OzkpdKfKAQvyWWup2hqUnE
+wSsiFu/Ukd6Euh+VopXmg9LZQUb6yNO23tfWV7AsW8qmCJlcDueoveNgERcgnwB
UWkrvast+KZ6avJLcIWUEmiGt3dgjyVmGrMciCaREWv4+lmBeN2uOAIEAhHuWPHK
zazsIH5iewoefBxzauo6DK0vmGlQKp95yr2mlCte64dpdWMs19YqxseaN8TUnxqm
KCiMcymn2ixiiMVC7jHqUXasUvGTwiHFKjn8W4nQ+R7LQ865WsTbXnkmJMGi5cnz
LL3nfN9evKD8CjZFxlRPXIp5Rsjy6yuCpAj1iHXBbaW/KPBokHNh6t4pbY6Xj5SW
Z8OV0pDYjhQkRAi8Zg36sBnkSaUM7M8yp14BaaaFE8u1BMbP9ZfquVw6woh/lbFC
S9MlBhgqGV9zXOuENSDvom+u9ELHJzQqvl9Ntz8/yIUdpXhC4vvrxX1/VVVQhbRh
XJqUXq6AdqSWEBs5Nsqqv8KMUqiMn9iO/UyrsXW1nYbDWwqvTuIrG8PVR/WkoJhF
i896NO3EVEkcLFizy2K7JJoyNUkHspVbi59rOqaN/tUutewl7BPwVaykMZ1xOeat
EOyA33nMj8CdNNKVHLf+O/hgb7M1e8Os44O5BBcmMny93ScZZbRfuQFenybqxWdv
IqZk6uCLLteEKZ3Vqh7JlYaOeayMHqdl+ClsXd4CwSEwIZfkHF//ZU9ClknvSvGr
oc4hyaa4kwpf26dchJ1ckB5BPdr8LxWaufTyWpVGkHTeiK8uYhpNBw3k/kAzsJiC
v9VVDmByxLwfr5Oj+y9wjk1WrFgzx932QB8q8HJuwZMYHHAOil9aJ8g9a2ASXBY5
rgVwBCJx5SRD8IDG/dDeRlwuGaer/E9cgzchX3fvnyN5QSqh5PEW2r5GO6mNNx00
rB/WF+693AX/eLnmk0JpLIe9jR1YEhfb1oex6/6K0YE06veQ8ouLNzOtXpsps3PM
c6uyp9Oxg4AjYhmVYsdkDH7yRXxkR5+W7CCNDa2zPwbYdvn6Qp6m1anzRwrutO99
shVSrf1XQf8zYztMA4hx8JGMjZ81LenBGYKynmLmHKUeqwxoGSU7FBm5W5vAbb6n
CTptw8ABgqFo1PWT6cZJDF973J7WdtaHpw5GQ/8kNJ5BVA7dllZnjhayJuBNHrlC
K4bF8JANxWeXKevX9luyHxSPCQK30/GkgMMtIJbZ94TX4suLKsGh0xeiNAsq0Y9O
amEw4ggsDe098f+tMCL/ktmjf6sT50ZBmWXEGSs/BBOFxVI6d0z8geFhj9p4X3zg
luVUNiBAeFQMVknPzyo5bbvuZ7K67wfooBFrzxrdlZpdHxYltRSKISUv/NXh4BvA
s7WVwaBTjTfoih4b8uVZKoFnwFQgbhGnz/cNNlfvoh0gZ8PmUnE8oA0TZEIWB4tG
pXAXsSplUSerYfqozT/iTcwTg2YqBoHM8x235+cGg2TqfpWRQ2BcRP29sQbx8c2S
lV4+x2jheO/9t60NEOa0DTk4EsDMTJTNgWKhX7BBQInQjeeUtpYTwDFmfD/BETc2
4+StM0ie4jqs4GOjHE45bvpRe3DB/b4zQe4OouBvL4krt0lTptNej/kCEjJwu7Ql
N5FjQPUgPUCDSwutYKxy1I0nIEFOGYETPl+R6+pub+Ntwxutpsf96bGAqRTsqUvw
JA0qi2KNwS8qUpj8Yp1B+JirljNpOdpKcjWl7dwWws2dvQd+vNlSmDbw9rWN6DkD
6Yft4hirMnsnwTJ6JI0sGlKuwmblA1yB5vVnbxjaRTZUYqSR7HGU/nAfUdGXbveU
0+MWW6bhpWsXdLJl78/K6WLz+i4M/38IqfvfSDt+rHUgw8CjiVgXnWcnFzuuswAQ
kJLRKu5XkE3UDAUsUX7vmtifsoHeGAxP/4qzZdVWHH2UKOIN1b4OIcTHE0fkJsSI
Q8Yg50qgNUl1k/WxQzrtYnhnYn92ozLCuDWpEuZYCAuEqJt4vU/Aqe0qyYnLIt2o
X/5zBDEVyeU5/uoGlj6UjSoS6DuC0w+8XgW47CYj3MtjR/zYU+1szIiRlioVkeIA
G23z32n2m/CaBDIZcHWVXD/nK4okMjgWV5lc2MbjtJEgY598PRAsPudugUeceHTu
/LJT38tjiwvJUFoUhyBBqzdQhz+PZ9C3bU+pUcticVFcerLujGNXj9Ws7Q99skIG
bG41RhOTr0JuC2vDOLYNhjje2Y1xMIi+MGjhAg1K1xFDP1w2bUcffy/OJRXEyi3l
A1tqQfUhhS/VALf+e0MiUb1Xr9Oh0f/Crn703UePzzh8J60jMOaxkw/eA0OPFYCk
/n3EiuIzJvm6ogI3k1sm/o4iq0XLVnorwS6bz+dI7XVl+UiRrtKRMp7j5LwsgGwN
TmVB87/YFX/TEADkjioI3xST5ezKon+tUfAunEv4jlzGFWeMDmopSnZGMnPo2Shp
WYdBoBsOaS5uilbL1OLh9Ad/YB70g5TPsad7qbWxutSiM004TxCoun78rTi7YbPY
VxeY0NkPvTre0Pc8J9hs/5fTqazn+86K7FQaBuJIQC3ZP4AxwLnHCc8ue2oIo/yZ
wAlzpfCocILoA0ZsH8OIeQ7hoSjOhGnzHJNHxMDl2B4KR8gus/AKZQrEdHHLefSg
d+aoa6D6FB6Nd8WG7AdvhHGrFgy0GGbw/HFRIzRoMV9h7r99YxgZWSv0Pr9VmhvG
0EycU8z6jOav7Ouvzd6Hp+iYNMf4ucOydrUeInxAK8C+xy0M78OUNKSrIDqntvpR
rFdLeBeL7+9EBzcOhguCvYVRhpwTrDE39gWpuTpWPHYczYaj7q7pZE3wNw8VUo3O
lb5sosIH1/F2mB4l85z4YVyjSLJqDYSRQnbVidEdDd1l3SI92VQmp55Anxhhni4D
EmtJmOvos0iApipFB0fJZCjxCgzF4YrDQIPWVeg66eHtjeoPtDPsySGbBy4zuYY9
2k6VdtOVf109x4+wsLLamDbTnygy74XOSDnIO0IciRWfwY5QN6v3t+XcIcC4qlDb
XxDvyZzk8S1/M+QLXNNpLLtPa6F8uM5rLkB/lWG/6iAmyXvVL3alq/NJzweS3AiT
bkujRjVf2q+hCFK7qksLFrP9Kk7J+hs1njw19d3a5YCugV/JJ1B1gHMGaZhqgeK5
BP2O7L3Jx8WQVn8ixQtO3WKWCpHbPOJWZ0+O3VKa9/5UdvRbwQqgoIL1iIT/5iD3
2vWsDUjNoNMdsa8KhOYIaWI0GA3j4wf6rSSzxWmCy7UQzGKImu6DLeu6jun6kL9p
QVzKhzWdmpON4uvzaAkSe98fLMUdxgCRMneEhyI4TIWMmoB9ntHpdygELcCxLBAi
eYAXVF39D1MzfDDugIjRhzg/lDfR314rOVjqVmTHJZZKXz8TxLKZ5ztuIfGv4CqO
IH23yR8cUEsFBZ7Nj+rRQ3pWnCpteo5aKLmtkImgoIwjVrNTrmQn3lnYVQdDRLrz
9POFUsq/dlkIAtQKIjUnqqETlwoX5iDkixYg27t9y32o/Kf+32XS6kcaq26NahII
w2wXPDi6Rb3n0T2YpTBZ/Av865WMMjelcXEtOJEhQkUXo8KrsdX1D/RhqLNPHU8W
9pyw75ZJfYcYgPW8UtcdavSetBsreMLuAVkvj0Jc/89dRXPQfmaoSRSTJeGVT+tg
mL8qt/F+yXDnHNirb7j3pcSsi11jTSm/dAeM6QolLLxbDF8kiJlxzPl0PDBxI+6b
omW5PyzsXN7wlI1hMlj6NMPNfZKEv1ufl3fumC5vnp8Zi0TxmUqFMjFz+s3sMOE/
D+nX4M2f1qGjdZBdfS8BLgJCvTyiNJhLp5Nu0YVJLvoyS8clMyGT9Zzrfpdj8qOk
DMPGeDek2p338RLZDUfyT6XKDvkYWk3v/0kjQ34ekMxOuvHH1y5y1O9FNaeZgJRQ
cfVMgUy2+Dh7ZUPx/xXwxdFqnnWsLFyTiLo+kU6u44EjVUKZZckHPsR+TQMIm4Lp
ES8WWvwHEUFFD9wnfvMFreUmN0gP75V82egk8IFIJQMIA4FygVZNM0zgX+S9h9md
hDcOpZtA9q9K68+H/+SVAmSePTQFbsw1o3+tN6SccEVf9hg52l1KR/Ja49sFQdYf
rr9oQEMedjICdG2AMR6Wu1GbPDtIvzQEvMdG+fAEP768gPNBDznoNiKWTUbPtcFo
v1+qQlBNfBG80yHwlAAGRT8KlftWfaceJHfdMNcCINXRGB7HGmXB93zO8wPN4msb
jiA28+o0fJQ04vpODWrKwzH/cR8of22jFmT/K8gJCB7ANK4uugii8vBHpjvCGX1W
DaTB/nPKDAwjkeWx643mOQRKA3f+TETrT56/wW7jWPh/iGseRaKNtNfFiQTBJWFz
iafHzc3kA2uaCOCKZ8rJHSpGTD9qAIU+rQRLd1c/s+mzhrPnb+XKec5amtTvizKs
S0sDMNKIT4jsqq+3k+jW2T3DMfJT1jyI4hAzLHoQ32pK1x0p4NsNpe0JUP5nFLi5
AdQ6v6rkosrv/5B8TQdWxSfOMunzECc9mggXNsw7cLPG2eGp1ZJBk+LSD/XA96ax
NPfygp4Dl/ROCsvEZNzB1q7IX72dTk9Vn5khoEjABA1A7MqjK8NGzfWSQtPw1p6U
V1amatf1742oBV5/Aqx17+o02Lt3Dd9j2MRts+wviKcn+Ki/y0zu8sAiU23QInXl
9NF8xydikLUwgqTjqkP6wqHuLRjdfszqXKUY88olYYXId83J2P2NvRzbZw5OeX7W
sFz20x2zQM5TSZN7Aj3v7/ajMqvcih59r7QYHVLhiHx5RXJAWhVECyEvpOBO6G7Y
X4KrutIrkHy9FDxtfsRdaLo1jS10bF6fjjcd/NOYB8mvAMq9DJBih1y3KqC2Lk6o
b7K0G7GU0b1M3PkE2YoCeISZE6XGITgkTZC8FZff9CZc8jZ6mFVtU/yjQXkun+gA
JrF2txAA57Ote+kakWhgD6/fiL3hxX6A8Orhu5++MnkUUFJBa0kukSXAlYTdFUtn
AF+pvvmzHpPZoeIxw3wc8PgM16ySduDEHy2Mt7ux7vI5uhDFOr0+pJccNr6hXYxw
qFoXXH5qers+XTyl0YBD7LGZ2hKIWGcK7CDv1E5xE4WdbXOeVEOIMJfszM1o70zz
Rv/txHRQDM7S09EdOR5a2WEWkGYjMDMD1R9Tz4i9ya+jnUsUOAZMKr+aHfPcuDpU
HZB0lpUbZsB5OFgZPpS1tagdCfVqnxQ5+KDUMLFRG69f+yN59irfTaDOUNfCpjdD
+/JrFi5ro/jc6UdujjjQVeHryMOYb66fCRaIKcCNo80AEUw1UPxTpsJJ6Xh8anun
/iG9B8FduMtbdwyGdWEIHMuYRU83hpm+xMKz5L4GVdTsw00HJmBd3VdMa8wNjk4W
J4gbSFdXqSxk5M5hM9+cpQPLIrkWnv/X6J5RZlY4S/Bik3WzY7DeY4lQ1qY3m5oF
kVZuGvnDQIynLT7YzE61hBdbpNS6dnoOOa+eVUzghvNJovEDzaC5puQf6o1Xg3ll
k+ze2Ed6dYOP/v0g6LDdM3sr3vjIMWwU125pdhW5SFU4vDwjrnnQuGzqbNfnOaHa
LGU+9b0oqpuH/L4h4j6yWmTY34gw4ugz7+2LPNE0uaJIjcuxb9jJslYloiUeUHk7
pqgjN5kPFu/wjtXEIY+AVWFUYp+abjFA6tLqEzAbLMlsQphh/gNj2ZRQVhWwEXTi
nKYuh2mEsT128EVazoY6smhLIXT535VVMBneWSZihc3Mo3f4bDjgVhil+bmk0uce
vf9qz4RNvmRpps/fD8Jmv6PMvyxO3KlNPPJcwpxfYYg4dV5tVMNYPG1E0n2ZVQNY
4Ie0mbClyY98XIOcTpxN8CfHOLGib4fY0ZqeBtY7AINP1z64udvrmfvXZ3RD1pvF
zOSsBXJdEXm/bstcFEUqKOIa4rzIxYUk38gyTnT9xO1GYiMUUg4I9bwwJLZTComH
JSj2x9mSY4K22NMz9MA4m/ZNNnLgUJh4evC4r+MK5Rg/7ZE6Iu6oTOcpQxn5n9yc
jzPFed9j3V8BNdSxRMWE1LV2tBVPbzDemlWu0LGNMlBajL8BnwnWsBdu/k9WIFzw
b2xTGQYDhhkqcpQtOnyg1jLcAtG20k9xDL73NGg8a8L5YSYSusdn6zAXHEJcuS8o
B0o7j83bc+735B+PIUhlLRlEYg8gHj8x7u8dvRUij45kRB/nwZE50TYvo/4tw1F8
Fq4ypgYEfyTV5csAAswVvPlHBmGoAq51RIKAVq26ZcdvgCpWRJvKsdlOdpDprLGY
+Fsr4/kBWDl0eg8R6ZPIxkQPFmT//CGi2kMMoY1d/X/ms7isFEu8oHoTryyT1kKd
oUwkpOPcKPJfmc2P78uxYj6BLnwWhrVvps6oa+mSOiyjJnumWPcC809TLZObGjGX
YrQGkiM8oUknYSXGHqgNy5yJ/vKPaE1OfSdxJs5D0ioFj4Ow0idJ0rLGmyhNLcWG
sNd0H+6MCYl3iBPrHXyLtUEy86fuPplGvqDkpqwPvm0N/fqg0qz4tVN4UYw/X+KI
vlMsM5Z3pJVzkxqopj3+0PrgE7wdQtshDlsQRV5P9tjSAi9IL3sdOamYIUvGEWzH
GoLB4EarYDZfiSiFH14rVRbN0zIKv3Oyo6Pk+UE/KtsNmN8Ckn7zTTdBB9G+d9pi
0Km7kCbA+EoBEfSbTtcT0xGnj77nvnUpf099JTNTRf5p/gzrHee2wbNt4DXCpa7o
S/P5G3nX4MZOiyLgiWh+vxuW0vIcBi56j5QioP5qpDyUl0Q57pqq8PjooQk2cmuf
CigLik9yYYWzf+q74w+ui1REARHYPUl2XkX2P4NPFoIgjR6KcFyhHIQ1lb8tSOM6
3eJ18k+t/bYJ4YxEtIjDchzEuMCpmd1PxewJN4oRX3Z0gHwdu0/mKflspAD9p4p1
STjVBmlgqQQ59jhlXHVF0Co7Go8+BwMa3ygq9P+gmnEL4KxsuM41SFPLURo1ByuB
zm34Er6t649RIkeyeeCf1bnOniVjbvRkS6XlXrMn4puehQ7tbiJ7aA8uqSXtrFJz
wK3jTTVTzQ/ksfquLRTH90ua3zjurJRGFNv7zMBZRjtkUwxdYvfi4EluF4BD+0kj
q6RNiPsg9OTp6+fS++TyU5gQDk7Z1BeKVVPJchyqPhkmyg2BXdLIBem98D016RUp
GwLFjQP25qndEcrF4ZgQZ+U2h19YCrQ92OSsV4J8/i+n5HQNDCmDDDKEhiEe48dj
2b1NWxQnq0oArlrsMKjO1GNM4RqLYKrzsMzNeJhBG3KnMW6Mt9CEEBFzdi+Tqt5V
o/bjTnuJbsU9IDJyAgcKCmSye1MbMlaUSvyefauHaBf/SGdXYGJ8ddyIQsWQoQd6
64PHI1yXV15cC/FiDTkVa1yFBcW0iWH/kP3jb+IdCx2IaR1DpBb4N1hCu7h0EAKA
/9+6marP7AHOIV0h1dZ2AKSdcj7d8kpQRMQd7lmeKADBLvnL5n3O5usm2XorTzVu
rkh+uN3j5tZxqV6XRjb6aKKi78RQzR4rgXveUuCgJErCM8Xk+E4HlGV+GUZNitek
Euoy8/kNy6TstvHtVO2qzOQb7EOsUUgSzSXhu2RjdNLexT7B+60kjWlHCq6nKyxU
YJWiQRKFVfah1qkZ9SVnAQ==
`protect END_PROTECTED
