`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pg+3BzKsYenlbDqcV0Nn6SfV7kc8VmzSPiOAW2sjxMsliseTqKnZtZBeGlUHEbAU
W+SUWLzYgRMvRHOkUozzkhSfQsURK9/WLU5YQBnz+P3lYwDkzuCnkpnX/mkxXmak
Yet8OzQ9VnF/Ifs9tYmNqQ3XA0qra0injXd0yc+IgrnQm5fpdZComAOC3t6kM9ug
Mhx0BJSA4xlSR3urjs2+zbpGbu0IvUOoCQH9QYHAWbR6mXWqqb74en7xtQMxZN67
f8n/EZd7WT2dduxOx52DMIr1Sj4S5bL2vW7nrhv3uhQTI4vSemzWe7mPytjXgnm9
CALXfAwhquqZc9NJDa+mHyRq77FmT3gHh2C8ooHTnMyKzIGHt1i8OHlS1jVk1uZ+
24qlmlhZ1fFbS7d71+DuZcmLALL5HJzyMYvGCNGNSDY6mUFWDTg/0mCo9gILROZn
RawxnfUu3wdOeO0LGVblx29jELo7R9nB9E9KBmRjmZlM6UlYdimygwf7ML+FH4YO
823gx5guIB+In4TQepajX3OL7eMofG9Z8MN5CLHU896B3u4DBKn2RV+ZsjK+crGS
5yxSyJLf2RJs2qdcMRE62V6RQxnqC+esciDNFdyZkQjsyb+ZS7H7wkq8zD0v4XQm
bM5dm1OCNnyQsxgu8EkQE5K5Yc9XO7CVs80nHmk29v9dgRR3bTLTMU1k7qCpd6XZ
hrfoDW/SzxUo4mMN427rhq+BtueInIxZPdUri38q+Gm2qvJe8m5FXLB/zS4kMnf/
w752XN0w14rwJn7YlKbyNw==
`protect END_PROTECTED
