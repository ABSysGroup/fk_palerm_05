`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VfZZc6jYDHjESVM+biTmN54wU7+1yIZ0uLfX/nCWs68BRAlqDa5Gnm/7ldK1O7mo
g5pj8W0/b8Sgus3v21Wx/h1YlSLEK2k65T0F5x2986ymR2ENofxkZmp8PakFzFwb
6dvy5wnc97ELpu+tRJRpP1E0C3xSgXWd0A9mT01WWuEkSj/dZAbhwfCqlXSa5Zqk
LAEkxL0dS9b2T+AqN2VDtOLw5vAhS2nPWzgoRcgEqNgBEsKj5+WxmUMGIFYRAuV4
lQeWCuUS6RlByIaonjVKld6Ty+asZH+fvFgsiNWdV9K9xX0Qr61IyZzG2E1xdR2R
6re5qkrRdtY/Fyk1Xp7riNcAO2N+lmn0qhoU3jOW6tjx8YdZq8mX0pEBCwrAPPc8
DpzEZdEr0cHHORm3MQINuxrz1DXIrLz197K/ue/jvd8U9/DeJlQ4RRM/OTz84DBY
MvFC5uW7ycdy2ea4Tiqt3diSsw73xmRbDJuF0BRj0zi9HZNuxfePDFsciCGvz94F
TthnGYb3pWEBwtnUu5w0U39FqzszaeaV3zOXKM15xl/dgv0azOAiAWDVYxLvJ/ai
6BY+U/0PY515du6jPUB9JwkecYCbweBqDE8JY7JYRkXKbaP0kx3dYLArbbNT+Hbs
WsVQ0sBwVEo0R2FLIZPHQLSNHLQs4Tn+vXLYjJHZucjQCrBs5de/wnJpAZfPlznN
8lshi5nqSuwxYQWL4e76dqzaqa+LHVti1EUtj1IoLmv/E1YYpSgCYjNMx9MmAy2r
Z3XcO1I04NAa3Ysnwzvn4/SH/+887dOAwXWjsKKKrZTynyoEDhl0ugZ7mg7BjbvX
XgNbo3nebLQOJ9LXeO6bV+z/g5lFijlufrTlBeFo3xUMqB+wL5+jklz1SPbFyOIP
0Ek5LwxJplxWrh0eom8zdClixveH5/AOnlPQNXeh3uowxK2UeHxZyXlKxHzSH3va
`protect END_PROTECTED
