`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jRhzukU2dO452RfyHBw5gCNqLNGMDidzPrZkoVWGyAimS273cAxZ4g8T/curszmq
VCH3IUgIC1/gJLBpXDDLLV4tXG+NPgoI7vzPu4pDmAtrZeMcQ6F4gAq5ii56R2Bm
HyPjPec4uXLV6biumD0x0Cedytk21L2qW6I0cDeXWx3olK5cuUdabw7bpN0UhX8v
HWnBsEyIOuV6C6Qm3Wm7krwD43oV38vZbEsYomeUYc009h0Sy6XOxSt8nV7ekeWV
kUz9jB8AuMR/Q7VbjayuCq4DfdpMC7tvoHuidF4sVWlDnZrF6B62+BcWs8gBqYPP
x5aHz5MNM8CaUR2yf2MU4pdM4v45XFvIBNiuQACyfrFPG86qdmdV1x/Kskek4x+H
+07X0RyslOeF4gBxQD+OdbSMFEMbNO5muVO8oJd3Wt5b5HrHKtAFObLdeu7mSpwt
uGvmP+9+uHqjZfuB+DQP3IDXG5gvWLvxpotAvWwsPyEGdO6WFhhZUEetHWFzw7WV
2j7o1TrrKEt7GanGxXHRUrpDOGCoSf6g2whB2hSu0YHjpRyalqQIPwEHGb7/YRlr
PgEs/GXm3FGP/bR0S4JWCna9TzsrITieeIa31qSGqXnCX1fsid1zeKfFEyen4RwX
je+YJnRbBOJpAsaDSe1ccQ==
`protect END_PROTECTED
