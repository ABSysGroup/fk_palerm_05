`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GMRiO3DGsucUhfPx4PCVWG4eeo/2VMrOg4vlioXuY1J7qr6Z0Iuszd8V9rpuOf/X
QyLWfJLtweLGCsL8Jh+qfEk2iJ3FcwyrmrHkN5GL3wscQOBVQD95pfw8RrfTFpj0
Q4dNF2cpdpc8QCVAZBRKYLFKupk0xZgpB4XY89qx8oRJeMfZbw+x2YMyG2BUi2nT
Qh/8/xCuL0EJJxOXMej7CEWrHb/fCSYNkMyjdt+M3rTX/bzwrwav3HIZNNCFcdEO
TuSeDY78iJzq2eqL167QLd9NrDDOscWFTO7JQAt4il3Kv8tFOWeCBR5TsfuOj8WN
9D0xfRdK3zRQzMDrXk4Pwg==
`protect END_PROTECTED
