`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cI/E/v4164dVRE2QH84kC0g02xfVlp2T9tSB3mt69IVyI0GreL4Oy2Mj0yIm0uSD
KExC1tN0pR4diJYEIX9y0qTuiQsSXcnYBeb61IEKpBFuMMXnkp8NEhLYo77s382V
HO0otRlQmtDqYewHqs2+eZk54P27B1ttTJgd38/oqabG/EFenopyyAgeyKDrsH2e
MZYgm+A0xVrsvG8WNpnht9JxgfoIOt3th0KcxEUEOZ9r+A/zPiA1nqs7AW/tIGPE
QlNMCwq6+9msrPtxuQ51C9WXWGMiJundbxOON1TfssqBKl93PRkjQNI9cTho2OLy
7Ni4Xpvtfbh7M2ieyMd39pXcpB2ODOPUlfXrZy8F5vSrKhOx5Cl1PLGbkziPI2e2
YgQ9ziZg8IK3uSwhbwzc2C1fMZ4glWfmmc12dKRWRroz0M8EOR4yP90uhjc428an
qOPqRmiJKURaIxwwz/Uw0gphXGpsPWH4jxBUwmCaC+ZFpbs536SPHvVtQpKUWUOv
ISgWGAhIKXm4ITY3q6TczVOMGGc36OYqiyAbb31B38Y61TcltNZn2WR46bqyhDvo
toGVEhmM6EF9ArmmsPWZA3Ta6QW8edKryTNm026XdiT1C31RbK28heOvvIiWAvub
ydo9dHA0IMlh6Yy3nsh0X6xDrzk/QzQ/F1hjPQs251JQDP00y/PPLCo5gIDfOxA2
N6462ULBXLBl1cE2bzowIf7ZBncvMRTDvTQ9UzKTIxAr5JaVS2AzMFagCg315z43
EKTjEqZR+Q8U/UF2xkXo6kfCo5rh5K3E9y+CGYn2DJlql1mnxB8Bv7zz62pidO4c
OnvbOzs1CS3UR+VKKqE4oVhe9RiVnoABTTYGg2nY7OuIrGsE0gI5kJlB/lCYYGH0
vUy1EaFp1pOOcVfaxWNhUMT5YjNf+TvbYjYg+zPwvae1Sq+yHnCRYZA6u1FeIVwf
S/svfVAcG1jdSldOU6SzfzuefuBBDvzU5FGs2GIWDadvtMp/ugxs4PV3dTvB3qqF
2cV767GOV6fAW4PWPvZW5DUkr1nZWV5CpeuKIygDL5FjZ/wSrWfkKxEmdxDuws9o
c2ljy355ZFm4v4kp/MZl0wVMKmY1Z3ZwdSFyfTyhSFfTPDCGafATwiE/gFTn9fE5
LjLEM+hOCfhfD5Rswv2gLmTSbci0jITT0MY5Fu+9L4Y15F5hGp7GNMqiKhp93yJc
hXfdGWlY6pLcYwkFKQTXERyfvLpJXumX9CQIVKq8cojct9mbIUqSsYWbP6jsE8qM
`protect END_PROTECTED
