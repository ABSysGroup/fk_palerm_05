`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ie2/Z7STRWWLQoIle90TlwJ2+iddjrWS5vZk7Y7J3MsoGzG3qudA32hn9jhdRgae
+N59FSggR52ygV52ZCLGRNMR3RF8kG29RF+Vn/SP8AwtF/o8HrFBovKSXehz6/rb
QkzG1QqK6jo3Wvu3KdGeaB2zwLvD3Pb3sfAIWzCLn0hiW28Z6taW3SDxGoeCPJCi
o6DiFO/ej63hLC6LkbHA9G3EPk8hh3NAKnINGAgnzdOg8Cpf5zi0kKJex8rL30iC
tPnA/4E7AFpDgS6ATM/jgE9w2bY+59aWTuhmzGM3e9+TG6IRx4oDzNB7cLfF1X2Z
CP4789EU1031o1q6Zf/Kcsu7ECQK+LkJ2S9AjgDux2G3L/riArEbB6XHnn7k2ezB
DXShCLmAQ9qPqz+VSrqCVIJzJ74yJY5uO06c5EWUEaI/3KmSeHYqLC6Wf2wlO9IE
g9Z0tGuxpDQ7k4fpOORHnsQdlVDUssnJPuMip/btyrFJdGeBkGkhqOFZspDSd7LB
8mooDZp16ZMSclLjMl/vbSwN0itC1wrnUSib8987pAojThARsQA8mpnTPDyuchAs
OraexHDWavDlZnC7efLskWQq/+PbBfUgt18gpfcQEV3ESFjRAMIORYyRiR6hsrg3
m13+PNLlE9oV+6JhgZlFeHt9M54OfoOI/Hi+voRTanK06V75Zpj7Jtp7INv2/7P8
IQbJ96L528Bk3J8m4XoLY+kruzvKVmW6cI0DCmohEz9D+SNoC1mvqLxtWY9BZus/
AlARByxcoyA8Mp77N3B34ByrHT1RHraVbJiuKOAdsIU8ydeFIo4PwAnmV5oUupYV
2zKTg5NekvZcmxpN99KmsPOJjhb2mtd16ljTBquyDF51MIphth/RwvhlxsJAtVIm
8W8nrGcKRZEJZRBFbcuimbTZHElr5D3EzVMR7s5UWUvCHpN20J7zRAgSBsTAb/Ah
sjSSsShu/DpZ5lRZLqKm4WODsJ3iRD4LEJRI64BZrEn+j38U+N9pZUtYtBa9iNq4
/kSyVJDgf7bX1JBF+f/03bNPNLA3vXifHBIwPzH2OpL+f+0fK7pFGcRXfFhsE2L7
8fz82neuKD36Zz1YGiTwaW1RbZecg7ptg5tneSEIJxnoYqBg0QXmcByEAgNKY5Yf
nG1pp4tvkPLyv3Zji1uYpDCqPsAaL5BVnAzpEE5TCjY5OpAkQ7FHPOuJsj3RdkHM
nRX68cFAwo/i42LtjonMZK4qIkYfQ9vuOuIO44HEDrFbcCgLP9t4zMuFaOsVRLuP
sQQ15So3e3WzWp1AyuqPv4idJJmnlGU9ZyH+bL/Ylm9Df99ehKLZ/0BBSRMqfFdB
+S6oDhaPfcCK9Z7QVK7pYCpHV8ce1Kb18Y7VDEplC6D3N2dwyr1sXPDtdywgfJna
sgDTAKgrCZa9Jn9VJgXr8k0jB2AWChdR6/XwDQkkLcwjooDCttqUO6RAL88d5GjE
34lU147YG/C9sdHB3izGdQhyBkLMPcjfbgLs1z3jO++eM7qV2PDQ4BwYNAkwdf9W
WWEesV32oy7uMy8Ao3HCEqAGZLoMtoDDBNGk1fgos68+CULuCcGI9LBOQjDaOHNY
e1yWFifF1L51lqeRE3M+pupIOmv8MxeRGYi0Lu81fKUc73YVCD49f7i45tCma3CO
pyh2vGG6JYxL9IlQlss7q5rf7rfnm4kjHk13c/opmj21pncbB8BklnyJCk33yr1X
BQH3sRPTAgDHLI8heaxJsIP/aFENNTXriTMNV9TMJQmstM5tRK1KGuAM7HzIQVTk
pXRsLrPULKZJqnOMXsjlL1l5zGPvhnUOVB2zA3OyX3i4b7Is+PbHLq+OxHRI0Wgd
heVxbxgING0V89j8zk0dgQciujztjyxQbaSWjj/Ur/SOX79Oc1bN7jspm/B9F+H0
i74ZsTESoI9w4NmyFJ3KqtK6eC/vANR09VOfOAh2jslcK+9GOO5pVFxrdDIarpJC
mYeRsdLvN6wd0IQKECpV83PDJNkJNAA7GBjaLkB2xP5m63JzHVWgd46GvXO90ZMi
zgbwzhbNr3epeuGWyf8mRjn8Zd0220XbSBCxZ8G9T6dlbLj2bu9Tb8wrDtUf1pW9
TWc2Ld3f4f9HXvigjdJ3Xt/xgx/pnxEhVVGitNZLCpxxxnNTWC51m4S01mGsGOgW
sdHVmozfey4PB/eHzLYH7FljmzBMgEJPmQ6iU9YjXhLc3v7Wag/MuRFfufPuo0/G
iExFKsDmNWEYwhv0mssRhU4O2bQPLHUL44s+Tj45kjZqxoRTxjk2tyJT6cG3AzE7
gOS7ij9BSg/MgTmyfp7tILdUzI2MN2Pxvza/Qrdg1qKgW+1mKDdWnlqNO1kxZ/qL
JNeK6koQnjJ9sMKb8Db3gCEKjP545Ac360Vy0C3jxXhkhNVLl4GfZ9NLnGh6FyQB
tWdExk2fdKlKaihyNtHpN+3Ik3HiWnrB1S3fjVRoZH57sJihgtMpFB/mw0rjFoIN
O/sJH1EQSfp8EbZ/GPUprFXIPf72A6Cm+N64v+Nc0Gb6xkAH5zgkze7qrr8MHva9
bpn+GCF5amZ6A7uEPk9ebjUE1XlUWCGf39nksfllZT/neTAdabz0knnKfj7MG2Vd
tz6hFcjBZnnxqIbVZiku6GDNxTm9Mot0YpU017xoOzbn9TncqSrYmIZJaUwlrYoU
SG241f521bNdQRawV6aOOIAS9Zxdpe1hKqj+AtfLPMpvHDOvQ0ohaM82vt57jc3X
wUBN+7YfRegVcSCzuIo1vjzc5j3j2w+/w5Su/WFhVD55jI5qQNBioUa/jZJNuIfx
WGVNyX6XXs7SwCoqxWXBW2uimuqPCGaAyXeW6wMrlG7yC7MrOUzjzTSMXUmUn4f3
7d1T85GICRZBHkYAJBxtXsKI0rz2Oe0GsTN/U5fJtAOFKlJm6eGSzut9YGNPQ0Fz
pz+hbYLGFZrAZLXgqC+QIvsq3HvvP1Q9fNmSZSWdntkjrUiXCQaJ7RTXVE81S9on
9rEupeqPAAHmFOZB+U+vX2/RlCO5P60AeQN7iZIrxeQIWvV1xfMo+rh/kADR0n5W
aq+CDdI6ja+esAP5klHOzbTiVTjybhBaRK06fg0YllaebZAIYRwGcDEIp0fhZU6Y
tfI7kaRK/Ryy7Izqju7hyiLnkw7V+tglHlLW9bdfdY1MOMFsnAsmIinWEoVpmqs0
t1tYTqJeukzwF+pJcqkeFAArrwAiDo0A2PkakphqOzSkGAn8PlQAp1tzjbK7AtwC
Yt8ZoFYNQIO9q5MxGYpfvXRwajyXqUXAj3yAWrKzi97ZcJil/gJ9v0fhcy1ci29B
NdnesuDq0BDDYrA7BrZoBthioRKz5Sfv/zkP3WN9nuQPU/gbknXwr+abfgtZ2iiJ
BnhS5vulwNnW+lhc3hM9eKrnF8abwLlJUGmdo4IAQnC9a+sTQ56BpMo3hQZqqo6k
iMTeVrU2x+hr7p7+2PE/GxXapXfzc92t5cxC5KI7235Bk4nbtLal1IWQhbQjNfT+
tI+L5ORIXTvjMxJjb5V6R2Pc9xZqtOpANlIZYsahtISm5a2EV2ahssGjsYZTkDE+
9gHNZaAl2rrIbeRWmT4sa00K8sviQbBS8hMBez65pWXjmVHp1wY8/osDS4oBofao
9cE/m5k0iSCWYoCq67+Kzbrd9b8Rx0D11xAjgSvKjgpJ5dhOs8URgV31sdRQ0B3+
okUMmWWILx1CJvkMygIhKIgF4W20dC08wffFytaVo62r3LnPLExjH3AHkdNh7SE5
ZzG05sIddU6/V0BcOjS1uwCWHKAuc4ZA+vDx3+7ThUQi/aJnr+chQJlm05byqsfZ
mbsQnryZY+W4S+fx2RxsXt87DvtwQ18C372Jz/HhF3mZHiFCp6LXhHCNr4NKs1DK
4E+0cOPwjvBxPby/dcpbjPATayrT5DPUEmjakwj3NpLL3KTCzAwCF2Anloc5WWdZ
DRz3KRQJwyFFzudisTSS9s4avL8fNnAnZgEUGUq0jbinXgiyZu0R9oqbDxnNA8jM
EWOfWJMItp0TyjWyy0sF7OqKw34IHZcNs/b+efai8+RpdBesLeA7OSRjZMdnBBfa
K+0dIPSwdbrsOHj/FZ2WjBcS1gKtYQgX1yUa6/o00Ia30m7ObK2zHMOHmT8aVZfH
jvn0jd62ViKmxPCcj/0sBl6ZvsGDtywz54lKyi+9VJefRAQgWe0GbZH/Y3OO/cQz
lF768t1E2UwlRBeRTFx02f5yKUvykm7IDljsI1T88dGUSlggwKZr3rK14rtHfZQk
Lf206Jik3FWYOLx3x1f5Chxf+blwHJWk1iibaJvkhA67IZS0eUqiaY6WAi7PeaMw
Gj2QNGGeoK2SZppsarwWbyMjVOwTgZlOfdP++WxDJp+wyKjf3Mm3sSqAgOfkk8AI
n053AGVlDdr/WPLjLGDnS7tC6OC45S5QMeYu9nJ7HaNybZTkxxhC1oQt0q3mi1Yp
rSMV/zQ+l/Of2bELXCfH6SdNYsgm/QkXZkQOZ5YvFN/Wfp/cLLfmA5bMyqdgkL6r
c+wo99OxlROTrgY3fK8QkhmU7u7Lxxy02eIXFXzAiHcRKAVgDkdeffrAVpPd0exl
ANSOFi5uB6dUF5HpRRILKsTI9sodmCzuWveIGQta6fZbPVpPb99XTjt9t5Cp9VW/
CeP7ZqxVQpvT7aCo91s57GRh2rURlzwSOqtU4o59WSOSSBLh35qucRVHE21wGzMc
qk9Kly78QNESBllHW8aHOdr7wPH31KAXatcNnTHeXXSyt74PoQLCUjZ+z+8jFPcj
ph5hrxWaGtyu981FgDaOxKpDalOAHhyEI/qRg6978XWI2XXrlCan4ox/AjnZmbjE
G9kimSSXS0Jd2Fmq7YjbbJLW1VgQhqP7uU4bgaMkHGdHrI2xTvaT0EGW9VyQb0Rv
5sbQHnnEerqIQZKVJoV03w4QlI0xohRIySCyeZHFDH7yh2l1AvFUStGSSm23Sv8q
pguD6GXUD3QTAd2btWIdFz06CDyFL7364he+ESx3K2J2pUzHUuVA3N9+9YJMCDfo
YJ3o1xuFmRwBhCGdLxOjVaPjSLYvYbK4yNqnIa5fzgylQS9uvOGtCPLknAcqaHDM
plZwJc4Ae+QuF756aRd33WArSmEgf/z5tPfo8dWF8wiXdhfKZgJVSNwRX4NjVyiz
Mizfy2FscDiQQGXzTMSqTsBcIuK3hP7Nwu2tMxJtmL75jKNbnEB5kZVWthn4TX2A
q+WqUf4LHXjjJ6I8TCKPz6PYBl+UzmkpcDOIX/2v7MVm8fDZ/N2hAK63eVLc1Q/C
rNOp+Z8rBoghjMNuN8M/w/LhyUQGSoabfRkoYO90aIMwnDgsC1gJFjdeiocKrxke
6Uwg3BIdSxJd0g9UxowRAd1DR+0Vn/FPiT72/VWTBhnS1EnjASkfflGZG9I2dNp3
BGPNPmPij83JzMGKmlYdeUIylOOaojBBSPlN9p9EF7tJlYG13G2+Tb3moM9Bclpx
nnUc3G2Jv6govckpF2MUkismE/Sy37Fyal1VLE1Hhk0VHpGL9vZhv892fAh6a6LS
KFpIuKgdxy45+pc60Lt4LHHw/99uu95IAWKWPJc1bg/+ZnIu0O1WHmE5yUqtr24s
rt8pBXepfQfRxSgg9N//V+Rf6CDYFcAm+eeDO0zrFkp9QEz/z0/9e84Dd4CAxZd8
M2HpzK6jAIcVaLe0L0NcoRDLSLLGSP1+BKc5xYqT7x5R8uJflyyBEj63fkepA1MQ
gqkHfZXdKOUMvGBtR9A7pZRakT/853PKHEbwPkuX/J/tcZQVjHyd1ZBYuCLNVL9C
S4ovG8+XTxKsfhTtYeDYG3T7zo8N4CCEzUoMGgrYj7Z7hfZW/cTrekCNN8W4VfSa
ACd1QyFC6wZuMvWTp8QiKGYawuoV/dD3UsgwGbnHi38vVCSVdZmczljeIR+ASVXm
LrX+GmMerqjC1Y0f834BaFfAriVMDo7wqhk/LWBtV3FFdF03nAOd8qXMa8QjJAyC
ESw7N4G/uBKzks6YCgq4zL8CPELxCBUjc0MgkVpDoKRyJ43t1lQoRrBG1O0+ozIT
emdgG7qL6wQyntIvYkNYMDoC2zD/kCiG2Bx5U4PEeEgm96JM+8q/Itjq7un34E1Z
smld31ihV/5IjbriS04qMCgkIQbpyJPlczP721/Eqa8rlvXe+wtP/nit+SRbDexa
60RD1HnLPTsxw8+S3zwLCWUHR4mez9M12iH5BttBWVJUvU381EqouEzGMnzMtIZL
JP2p7u7EGh3K31WtQo57Y7SS0fI8W4ZkhLqwcU5WUc/Tuc7LYDE0vrbqGtqPCwCN
yhRHBpBZv1J4pR3vsf+kyRF7D8Aj+oKQBdic60e/DYvYwaoJM0jGoj5pmmIsPTSk
k90HC6l+FQjtNZaWNDQx5pTXbmN7zZOl17FIPDgw6qdGINb6iTWICZ1gDKfMwYvS
g4IPgFsdqi/KqbGygj8AfV0twaOJhn4Ncrd6h/ZBULtpOK+CuDAKvcKjSTPA1PlA
vXmKupdqtMw9f9MzO0Yb4SXJ8lydhU7CareBSBoTJiyigN7891mwfPpus+sanYQQ
eoiujrL5oCEdrXmvI47U9Dx2WfJgXRHfW2DtAUc9bsesHM7D1ASpXQOdjfU1rUHr
esN++crBVeZjV9kSxQBCLIawUhEOMt1qo0PRxFstIMvPKXj4KKhLdcGmwbtXX34K
YtiMmtYLX9+f0/pvAT4nLFqyGyfGVB7WYsVqjapVkEO7sAXLYO3Lxt50Bs6la4Iv
cypKqfyYmNCcLrItKp+eABZmsW8eDVEaV7Nu6FfbSVEouk9vWTY9En2otRU/pOgL
eAbdIU46/VZGCk96kwOeNscXvEHik1emzWx+ttUX8+/K46ATPzamtVqjK9xs2Yqn
8J6HOYGsGPEkSTJmqvKPhtMyAM0sV5J4/N5uorzcF6v1KGJoWM4rRJLNk/k2tHZg
aoN28XSaxkJbV1r7CR+RhYDcGIG/ayVZDqrnez8q8fKwjWOFvVl8/KVh4N4O8FbB
Qc8NF6PZVAyCddKfV1wtE71JPDUHDHPbQWn8YTrNsAifGXLjakK7dM4PFFGh/jPR
TiMrX6kmrZNB1DwLlyVyg9x2Rpr/vTXvygkVLxDPK+u6TVaOnkXA06Gosv8RpHjM
yJ7oxkGvbqDL/yEqRHKhhZ3qj6QJF2yGh9M45gVrEocLYEyzc1jeRM9nAGWURLU7
7XXCVFLodz0YbHgtfcMLC8qMEYDN2yGGW1b1e1JXpklZEJPntIhTG0OvMH4cT1WD
8/OKLWRP8PrylnwgpBMpa8K81Dup4p1prkFdrF4+wOoPexdxfWJa3IdzUDyb90+a
npjYQLxGslfXQfpyUw4pHqKvKReebBvVieI2OTKUFKsZRZHmx8BjZkDMr5ZTfBcD
e0nxVowm1NV1kIGIsEV6baN0lAZYm/wCO9QogZL9+5PHGZv0NfM+ghXYIskRFrHY
PBD02YkkMc9iwr91flm5+eEV6qgRtF04EIZ31nDX3qWE4jDKvrD1jUMMGe7m4R7f
KjMWgU8AwygDl2wEJs9t+slalUeyTB2qqULpVdD+Uud4owKPr1z8x3vm5aowAQCL
Ptx2JcR++amtjrks/UtK6TaSm7nONr0HfcC75jDXO7KHTb7tHJcEgwiaD++AJfqx
3AZ4Il1JikZwmMdcOdkM87psJdrKIk5B41wq3/wXqCymtzOdgjI4v8X5UgbsKAns
xeIoq8fYTTavcVNJEoHxyGwoiubIBeHJO/bKir/1XRHoxmELcJM/Tw3+XJIZ67Pj
+TRblrscZw6jVodqCZyHfT0hIJPkqwOiLad3MmSf/GE/Jp2xRvDdTyvgtkqKyDSv
AJGmOKB3xTElfxtP/zZm2E3Milz9CWPVJZo5CGKAM59nF9AS1+CgKHij21j1xikq
LqTzdscNrewlhdKIA/rIqJOCz6BTf8GqU2EsG6qT4YH0UAskAufYNBz154cZpSDb
zheW01AXyFPCih5qUf4HhbetByM1udv/QC1X7bcoUHOjQCcPWGMMfRFkRUokFLCU
41ikJxoSoZOnliUSNOjfsaF6B7oKGIG0daEJ84+/krhufbC0rk5bR/ht2zeiR8VH
M3DPxiidEvIdcxdFOJ3wOR801RLt9WLKuXWmIQq7tm3peLNVXSaz2CQ6BcHiqZm4
UBuFFc0sUPS++ZL3hokKhFsaSOJFl+fwZRvw3EuSdog5Tpn2mGGBCjGHOCkY+5YS
3r2aHd6hZ8RbITPjOlMUPk0HJkQ1Suja1CYrIfaBOhMqzIU6tbYpL71+KvNPbR6X
x+YtkTDUozXkxjhObfzVuwFkRM7p01hZU0DiX9ZnxVqY1GcsWFqpvji5yWLIWgir
QGw8PK3+2S0kn1t2JuyfR0K1kykOFnwMuft6+sn4bY2hGZLunk8/1gfcSUTVbYFw
st0eSA83jSEvQCG8Amk8Jk4nDKr0cUai8cLBZpH2fDyF2JGFOhNGQTEPP3lykHT2
PV2C3txRPhcY/sSgwuE98JsDdfUigrZPR1K4iZC8MQsE0iyeInDuBaSdCG3n3jQi
BcnTlF3jLKcTl2Jto/znKaoTP51gXuvCevDL2jEBhA1qHpkR58IvOxvjJaxESIyn
imxtsQpzZ1plNxfg5m3R4AkVhpC/IbANupA3l3BMdmso1K36VvjwEVB5gGjPPFWQ
BZLkZQQ1V/faNaoPsQTm/9xN5/A6NUZxIO4ExypAdx1IAWfke2dJ6XCnP3TV8rVb
FXpFbbBewdWuDdaqGIkTCCusTc6iyR4DAzzLI3qUIq6I27fU63ihLMcftz9Wb1P1
OrtQ7D+oZW+pIhiGEWyidlTB+9OZYLmKXvAB9gnIP+Fr6z2nEaCW3HgjiK3KH6d7
7EHmUxCacQFrAiJC9kDhhLaM4Ku8FSeZY63dPaNudGeWCEoL4iEFQYkbioVEaLWw
+wlZH2tNwd6b+gAY34dtLItlHTm8dv4lKmO8gYThqjGsrtAoK15aIZ+iWVMdLSkV
N/yZRi81j4NfcrT8X6apA7p3l/wnKAer7+OEA3L7M2K0cDMN3a6ejIaRBuv6k6SP
ucnZ4EeCsJZRu2qdbvfQXO/sP3DuDk82SznVoqmMD8RpjVZROUE52Lvej5Lrvfmw
0BkLhKZO7iFiAuGI1cNPONfK2OtdQP/0xbf36wOIqVnH87/MOVSAxCTtAbzxtp1n
8uZfvltcG+gCkfFgWs+ZWRYQx7Icq6GF42kVo5KxI9ad00zfeItEiNsBWjXgCsJZ
YXIOKEima+t1peZ6+PX419CTsa+awsPqFV3rnuVQmccTuKeB2VT0aUZmcEYqk4Dh
nOyjEnBj5tj40soLeqY2ZshxV0L+PvA3FOElZIj8PmQm0XTZR2v4OKaEK5XItYrP
ofa/cOJWGsLDKWSK2swD2dSY9aBilL4m63ve+9QWBCC9Vk0ffgUfdLfNd4vlUOPV
CRhRPBphmcw+uY5iis39OIH5c8HccfESgaW3LTVpdsUrSdrvA484RmLoFn0Dev7T
sMg0KShNUux2YQoAu8Z89wTwxqjuC+ljk4OPRkCRVG+m+JhJMIoYI824tUM1NExX
gb/VHWV8wwAlvDIXT2x4b5RYKUD6R8hX6lsG6AH3NBm/8KhIppFN9efMVhLx1fvf
brZU/sbxXrxXkcTvF0/DsXxi8umywl1QSW4jsObYXOYlis4bB8zwFaZxwF8DrPnz
tZtulJyq5ofPMn2aIqeZUnOpaaj9RKjnYelk8/KF6WhDIpqIuY/AXZWRiVfdhMkr
ezATX/VuaXyd+w7F/7gfy0IfX00sdvgHnIjeFid/VwdLQYufP+kWqWi5s0xY7JNP
aPj+ddHvjAEw/pVpcJMDpiLOjpBhVP74YmEaI2iqG3v8lbiT7s0UOpg7eCcs9GVo
9zXDKBF6+c68hModBPbo8wB2iZPzKrno70dO+/KKcshNN42ar7L3KUpLOXXQyzzT
cpTwNlMN07EGqtQDC2/rYMCKj/BGQ35pFiuHFhnKUIyYoAauan+cY7j0n+ttq534
OgrHIYWqCPBS/36Q4abCURxKUja6NGgt4WvPHN08VnzPGhlTKcn+5FiPN0I4I/9Q
ifvFo/dVgr9Aq2nNFSUSJAtdJxGgDV2hiEN+5rtTdFZKYbm0OrD0OT55x7HOJJxv
b5YhzcoXgthoeyUg3tVs7mimvNRJNac4F4qP63/hiGspPaqgWkBU31Pjqh9CKZpf
boXMLEYJfJtIMvx+1qag7WxR94XVmmd+2Z/3roVvQwyoMYKqaIUzGCwQpre/x1hZ
PTJdA/K47dfFt6lXQAt6uYPSjS/Yz2hN4kDjj0DhpS2lmzOlMfRuRSzCAjZpk+m2
l8NFC5+RYwo1teapQxz3g9uAdJ/RBeXo4AaSDr8EGHc6jtGeDzH2yLjYzR6MyU6+
aR3k3a7gj1kXhtCqf2J/isjzHAzC6ZpaZ08SjFPnmLpJZjTI/xt794T5GLRgRTmK
pfEsy5pldKRh2nXa7n7DCZfi8VL8OVy029H3gcQCUik3F0w1JOMVRcAHu1aoKqsW
h2Oi6VN9EyWJFDXCLgtUwxiZRRgEngxjG+kNDqEaJFGhVohUMNXz4B0L1ZSjFDJp
R8+YMpRHZQ62qhJshUal1cL6qudWCpX9gdEi0kXcjXIWcSJw4CtxAg6//I3NIKM8
z7luchbbqZWg9X6F5SJwZlXKFqrZSh1KkVmGkH/xegYOXGwIbqU60/2FbKq93vq+
qdV3xIXPjaibZJJ+FS4FuPWyuxpZDpzzU4WKI6wBX3QCds/nSUlye7XykMf+G4CJ
v+++yIpGvDXohlBbV43FsjLOzprIjlgNqdOiZTlQBhBmM3IpWFT+0WJhdAl0xafN
XofjTzJ5tYrz/ZiAfXjLMbTFWFNdM/HqaR+Wg5c8ppQ3r9NrmMvhXK6ZNGxDrA1E
HdgA4Xpwh7BntGQNgkbz9+d//S6EzpZXZtYgkc12m3osq0V8QkIBRcg7+xkVVMRh
OPjRrz+Fgd3L8t3Onl5KfLVzsBRu/XCXV8blM46aKYfzY1tOxC4g+XBlMK4UD7dT
paueAjv721augpoR8vClo/81snM6vfAwD//ofPjn3CxqxbX4VHRJkCMWKwNba2lO
pCIxM3N7YbJGCgNdcKsVNmRPB84tl9JCdsjmosO095AAsY0EkMRhMAdWByUn+r2g
brKVJb60HRkcE1TlIw4WnbK8miHlQ/6u2MnHIO1VDiHxcB1gPeZYko6hF9hRPYrD
9CAkqlr4zgL6+ZMnKbZPGGJjtnWy0g4w9a2toLKUn5zfW+534DYpvRwHi30yjnyF
hdQ6+YS593qgPFEBOLbYjfS5J+ZXKaaK/1s1kNarZwSrH+rduGjUDcERWRV5RU/2
4UC9vXMIp4I8zzBo1VBmfapaieAcVcAn+IEt1Tuf8/l/OFBaqxDhg8NIS6Fm0Tl5
Sn0Tae4oX9ZnF7QL5+ZjNqgCOvtA+MGvcccGjTUhGlDFpBpbiPf1EXmfNDf5m7/j
SdATRY3plBIOsOdj+N2xBMFDqdOE1YzArqGGOUqphmZTi3MFMMiYd3d+aRSi6FlN
g2oovV5Op0XhS+DqrUXLbHNLK1z0uXypUcXG2bQOhwkVyFm436dO+xAGQMeUL22N
x2nfWWu+Swnk7sXtt5AjB1/A2LeNqzqnOduOyhg1HHP7FkXGI27SngdAR7/3vmXo
kYXigBoDZHB1+A0RBi16HRB6Nt1c3YGvtsTi9ffD1kvJ2uEpmAtr7AM0J6d9GU36
Or3Zfu57/9ZfWksLYXyyM5i7TSkJjqpD7YBhNPnc40w6BolvhS6b4oZqZ1iCRXsp
oI9MNdg7HlOj/DXejKE2fJPvKAl2dzXGJaJpwJHV0M4oXzLluxV9wjRQ1dtz4Rds
frVVz61iIiLYFZXOSMg8vTcr7YYyPHzVKwRgi919nR08WgIlcp1ckqXl9jm1MWV6
Pm7DDpxAhSWtdLDzbspGiQHVXigfPLpJtQDXoBxiRud5xy6O1oguJjdGyN4ZgmIA
NsHVCt6UYs1nPc0uXeb/7rxuys2r74RXbP7zwtrDDwKxfdqlQOHnwrFKDcFWW87z
hra0Vh2PTmNt+oS4k+6vtWJ7RBpV/d+XpLicIyUetWtLeMmXE5EDBKYM3kUsAWQn
gXapoMhH05ZUvJCps8v3h7mwPBa6rTFSDu4Z7WqIBOE7luStGuRqKoE2oylOsd60
QFKQGmU/1KgYf4Ep2FBSZxxjY9vAClwBeNpfSGTAjn5pEzgmty6ReynrEhWRlmfU
ATdJo/zqTEnWLSyNQWVfY09qyd3ewFB6QLKyqZw1iANpe1o0NFkLkMpkJ+YzJnFx
0jVQZ20xLeRSVNkdoScXTBErUOgZNK9VgziXoeiRmdND5BDjf70+sos8oP4jfOXq
Z98Su/slFhGQ4NQt5nADBMBwOTdaEQSfjS+O7voY6A1zF3n7ppVy12KS+FXM+zeq
FeCdrYUA9B+Kh3GFRiiECCe7VsfD88WC3BT/eYrdktjIO3wxvb4SVlUuO9ivSnda
rpz+KRoF80weuSsrhGdrCkomtSJ5PETAvBELzfu65ZrH75IpDozgNLSMrakwooyg
UchO45Ln+v8in756YU4J4ZFQ0BJerqLdSxwv6ujBNcMm/WiHidUZFu2Aebh80X+u
Ea68fAkFK746TwSyy/AT+h++CTq8anSd8IfRjTugYQWZhLEQd2dFxW7A0RWgZHHL
rgpHXL3Q1VBkYO+xLImaHNTHSKQgzIhE42yG4DitP7qYFr08XUgQjB8rsRtAyPty
LdJcmxGb5Dd9+aAI6S6u4k2tuRyJE/jbAITp3sZvHRskGrBCtOfztDMGPxnPoVre
E7sMKVUVJ3FhSkU+d5BcSeEVQJSeStZ7aAxin7WtY6uXaOdYlctnAqxDGWqwOR8z
UTI0XlztMp0d4KGqAk2USga5nq27XbcpUlCeJvGe5uO3+Ru9U0oXDRuc7ucJ9GfR
AAPY/z0LGGHKnfM+z/q6oWGETB+7ITRATHA+UmgIJAmnbEcng4jqJkxJS2nF7bBQ
N+oA8YoEUlFW2HmskjjanwPz6jI+r2V60QMbG2b0cya8CJkqDJVOpYVJvt3IONr5
4b+usZrTEwMRoD8TVgY3RoBwwHAdbnlg5Wo/j/fmWRdLu96vJIbgjUl9icAIh+bO
fwlJlVCvuwOBSRPmqlm8Rv97tSNepVINP0Fx2fBihgvWU+Pk/FlQ4QqqI2JT5BlM
UhAhoxHTE5dL07Wqt+Nsy+YFhbYzxjgYhqLMAByBftiRXsRCdtAyUezIDs0y/OoK
6CrQKGz0Ni8K/kpbNLyi0I22/9dHxej3u+5zdFAK2Xismi3yOIcVrGsw+JTf3RlK
r8Zq+3/7F6Oq9Us5s3v7Ebln1lRVGnw3szhEVjb19IbL027sgpCl55gvFGmoVB6R
AKy7S0aFlzNwKJM/9Y6yoAia/Q2FjqBaPMk+KoNT/cNi9h/FvudjW/rsOyLPT+cI
cbxO6m3NlwKeDUAHcsOJ0QUM45U4ePdddxGm+gK4ttRj4vAp0nhgjVhVGNSs1cpB
0wco2kE/6BMT+D3NeXjgNsOn3YEksdsk/dRFEm+lJUDI2zg4CC2FHLCdfqMX9wSf
KkwXFtoXoiHDWkpH3As9L6LGWN8HcBoK/DdMebMB0AOPdGwOhORbtVdFz2Kn30tD
fIYEHIa99Y+jXVnWPbzu67OlEDR3aDHyhT3BS2+aksy47gxSPF4lPbzpdDdsppIc
602zo83y1bh22d/nWsNpIwoancdSU5BxkkMaldCG0zaFpZSIMROJ7Hw3HWGuIR3M
CraZNhyWwg5yLFbDPf7AYDbFOkoLQujZSqNg1mVOl70ERBFwXWIgneU/RiPsGIM5
x+8J57IWUFMzGa5n2zD8jodMLZk/OvdDJ0M0Bbqm/b9jUPk/YY6oVv/ZsnItVely
XnfigjCvBsZ+BAZn3C5c/OUa7YONECalEcU8H5/Ot6hCDUBvtXX3Qzb/wNhZA+rP
2aIaUSghH5hd+vkB9NubU+RyjhrGIsfLgHKbeYWBtz9RAhtX5uD8hMQZRUXxf+Ft
U5ZKnMLYD4AMj7JTaL0Kvnz6VY2YO3qG7elu7jvXNk335tOGqFvvEPbDl7gUAioq
ubBXjI7nRaofBV+twbFquMG0LziGd5PYBVzTZpiRQ2aTsNIlTK8kqmtdyXxzY03t
BGRRXREqt04dbGHZFoSWilTo7/kv/bb9wzpF9sHEJj9hAMICuUY3S117DviBMI2u
rRo8KEMS0GqM4m0VBLRX9f0bPB87uDGplkWD5pqSWsXLXHF4ncfZ4MTljVtAJ41b
dQfIpBk8jZgakBbVDXMjTl9mwJDyS4L+Z1Xr9pNbEVSpRxlSfIXNox4Bk0Ej3RxF
wZyGpKJrSphBAjY5x7QjfXaZl0Bnw1aYSLNcQQDKJpfGlR6n4u+soc5omhhp/1Zz
JR1Nqy21PLwZro2dTlSqV8y/tuE/QydKbSQvr6B8EQj5u0RdiI6DygRv2Ff+NP3t
LE8Y5JrnK1b2qr81dzEbhozTTpKwx0/eRfXMSeQ454SX88MO8BlXJmE3FbhgflW6
Tpoo29lef1b/NGFE14qysYzRXP+Eg7ZRIGCml6aTMedML/kJL+vjxPAkfXg8er/x
WHHFjB78j+D+H+RMO5QzHng5jWlmHvHUVqAsE+hxppSxCt35pbW0Rw4GupjZK5b7
/Q29CDABFuqn14XB8+oZUcQkyQNDQss0IyWUUNgqP7sAYlRTITFxk0x8CLwFbxLc
rWElKfxBuE1jAOVlKvWn1XaSPlpHCGqnbAjLpb5dnU2PKj/tCpft8nwKd7tPelXU
KKcjQqmOkP6N8z9tqfcyR0hrwjnhbuew2jFlM3SyCJ4n97KELqn4AWhZbpx8AyEP
pi8wDEEIa7c/1rX1yPBYSBVFIz2+YyPb7UDPTL+XEXPSRuIOhvTRTrJngC+nrYjD
WDJoe/hTTwhLfktaFbfB2pjJ1JRHRS+SBZ7XLpuVWx7nfmetlCBS0r6iRK9dhqMp
RGrw3b9mKdqSjsp6sSULb7SgtGXgcJa0qHnPkq2sKqzgUSk0rrrRWEZtIBemRHQS
vwh+8VLPTQ7KbDpjIF9/jIe6IpnydveLWSmRBXaH6ELsePZypM2ub1IAMkW0viTJ
ZxS5DihWbB0CcQI71Uui53r1SNtdnDLAFH6Wl+aZKH4EIFW3VT8hhGZBZk/rzC6x
bBCMfoyTQOSe5YK1u6aUitixAbEDLXqa9pu8cmQ/JkzG8S4sVXdwJkOU8eA1KCMS
5ZanxuKVZNYVx1oEVjY89OKL1gCa6FU5hwx0Ohlw3u4wgLlGYXB8rvH5/bo9xplr
Nw2yuh6AqbjUI4nx4kvI6qyOfa82UHh8SCiK2lc7Fw+winKnQsPvpqmL8PTkqIwY
wEzUOc4TX0ysfYHVYXejE5/4A8RYUwW1kIUfMBsRyDlSirc3RSVwBKsylJWoFxV4
vdmXewSrvlgxBdOCg+20mkNEZ8sL5cn4B1E4qJvufA+vgVkXReQ6pmhoyuJ4Ldq4
N/57ZoFEe7H7Uz4ODHCw+JIsHhIEMrqT86/2nDNxfBL6OKA361G+UmfPoSc+Iuau
cw+1KAbxnXIWaqt126q55VLJK2uoyG7t3HXMtdhIaWqKsKXwtW6UJe2odJoF46ZI
/UVD8xTCjzUj3xXD5/6oKLOhKr5w3K5BOU38YQSwBptAY56kbNbOAwIew4xH/saf
8BFGUx3yROytq2TcJqRo9wC00hgx7sMHyCiQ6Qv1j4HvVDp+BLbv3b1lyrvnRhIn
YBaenQj8GepJo7+cwh2pSWo//9Ae5+Y7UVvmyOQpo4rQgLPM+lpL5tYGDu66Dt6g
0RUHzhCA+o8LiadIACoKTPND7dT3bDRxBAcuYpDM1l02Kz2ghgoE0pBIc39lfTm2
8o4asfIvoGbToGpUPJC5Sy3Sr5vP7QMb4G7BL/X2+f96z0wIqTazCytgMjw8/vfm
9aX3FQUuAxdgxvew/d1V5nRgv2WoT0ndjrfblqP4JaUx88GZ1LiGFHBYBikYwCsT
EzSrUyGcH1rvIrrSt0cgXHRvx5I9rjgybZmvp2rnLuGGap4eirr45CyNW1nGqK7g
4/ZAuxwkOIX6KLqHupbAmHSZYDncDhXlSW3LSjJj8TTT7aUqw4G6uT7pfdIhUx1C
87JiQcouliUvk+MzcKDWbDLg6ffbPN905cUc/KgocMCKqyxYU724Lr5kwkuMVWbQ
kMJF/Uo0KVRLce0x6AlQvM7jlCWgEUjed7yQplyYCzFybyEcryBFWaMTcv8yF9C6
xj6+RZJiQ+2RRodIM15RDSAblhAWfJ3DBBUcO1LYfcyJcoHlCKhheeMsTIian8Ut
mZuTJU/klnUmz3eE8mtPcxuoOJE76EKXJJCLmiIEEbNmvNgqNmK6Vmvb0IF0Y1F1
BJMrfNmAFfbOJbiiFXgLOPnwV9oxhQFr9plfbkdI0D4rFoQ7sIeyZNK0YeHdKh5R
kIBXrEVzNSZCjdRXNS+WxU54DWS55jKOpaPM0RCkgYcSmwlX8h3jrrHtC9FNNKKV
l7q1/HSyrDQAACDJ9bFYZSU8pos3qrJPPksvaKw7eocj1EJqYBgS1Lzv1AF/4Ejp
gzKvqODbm1SmGN7ejb86qF/l5xhGQRqoxhgqI6jokJI230qorhkzMCvP/n/Xu+kD
eru1bsZKGXJos/GnJLl8noQk2X1NqDuvdx09blAvjCwIMf1dDWQl5cFrB8U2NXjx
BqvqUJsGDiD98n2/dhgRZE46kGezYdCu7+8pA7vjpFrduKDkF3X/xPEuNjee0HA7
/jJhcbg7d6zPlySWnz/8kbqnwTRaVzFfdRDKSHE9G72EnL5MnSN3Yp1IOIUehMYW
+GxjarQtZzc6VNmN+mVWGcsf8wM9eiPiqFqR4BhMmQLyPtMbcrwauhK7k80xQU9t
zFQOhMERWVQ9FdNfSruT5gFUsVEruB7w+Q0e4A9etAxEcrimT0vGNRIWMX3xlvUS
MeivBbXYhPxa5UR0apKa8KwpurlALrYEc+Uem5zGdplGZyy5sG1+BK4bxEnwkzI7
31gnLl1H4ZbGFg8kyezF2m66TlhWIo4Bmtg7s0Lu/0qcWJFtP/B0K2JiIjIax1FJ
g3X32wAN8KunnL8YNmbQwbrKRAXjAjVTGv4X7PGECiIAlOdhdlIqHxTsoevfZtwT
Sgc6yw8DgoaSCpjh3/zy+K96aHTt1iJCz9NZni0WhqHPWosXfSq1yYEGYnf7iq7b
863D4ChqasCO0zLrRB+s4/KttAqvYvNWpYIpiJ8dCPO6vbx8roQjwF6fCR7YD0EM
m7HO6v7QqtqiXtxhAVwf/5PVM/AhZ7FZN6EGat+NVr4kghFN6KsxilczGnIgLO3t
GjKwNJmPm77wSO6ktFcCxH1M7nkaFryqxVWMOZFPEwWhmNvZFBqvbVXLI7ZY5OXe
kl757eXauIDvsfeS5kaspRWxJ/KVDSktT5aoFu7uQfek8HrYhKf6WxAfPE2lye5o
sRms4m3sT1C6QzhernppocoJ6Qx/TOS0kh3fUuokkbkHjIAOcWIfYGSSzdQCjcz4
+E+NMN5k67aOkzGI1wmSsC1HLSWixZxItS39HqFef2rEPO0hH3red8BDo/FnQ7v1
LThRn4oNqMOF72kSZwDw6QuyBE44NdrvtV/GMHBvbW4IAkCG2uKb4Sq016dsYqzF
HJ1yQ66TR1vWoRIh7c3Mi861CzfVp9PpL1ad/He9IdL3Z29JBndsmjj2QmO/1K++
9fneaaetAsCO0b76XnQXku3eD3q8dbN4UZ5A4RD8eTHiobswHPM200KT6hXOZopV
NVPrEdbZDKa8Zck9SIE/LHFTF1jDFJ8FhAb6YhdMYW80OmZW2SCxwv8jb3Yk6bIO
Xw/DO5mO1x5m25mSt49GejF/tF9q5pmJXWS1i+CxOSj30bGMnjnQMQSwlIzer6wo
hHfne44kkco2PpeLy3Yvu4NYlGN0FdKy2OQUxbP2UW4WlmahW/rRBcR4X90s/0PJ
Gx9BIADa9R1i5X4fQKYooIOQAE3QDGoN+a9F28mUGg5V5MICIMdzD6uPJud3UuHx
csgleEl1wU7B9pSuH6plLagFO12sApiGG0wLmE4QVZb2QuCGnYMT1lUJnpmA/uAO
rbL+4iDFH1eqkj7AeHhJBW7CwyMClkJXdOkqvncjoM49YLxcMN7yzrZC5NowCZWN
n/FMocsJMWhs+FL2kzk/CzqoSJnYNQe5D3his3iuWsczNwS/fHM+BJLkma1Nxwsd
g9viZOoZpHzOWKp0dMq7wS7kVafpZd+rrmsOHYgjEx8myIvxOQYxj9X5M/5WFkWa
fec3nQFPr734IW/7HHSID8L77qwvRHZ/sijp0/Q+vlAirgaXwhyywsF0nIOi0e37
B1zo8lf8nAWIvI2fmqLjO9Pq03tR0ULasU1XfUqnEMfKR+l5iC+yD7+bTvYwAWC2
vQhBqyRZZpNo0/LI7VxAYifeQ7X0SuFaS1zLQNZXr6k0S8YK6W2W3hTCu3V+Op/C
dXTlID3WVn+rAJbQY/nbhU0lkAJ8nq27LWRfwbpBQllmzIVYG809j4pRlyKow9JY
Z8F3qM7kgXL9GWHNx+6A2aNpdn2PB2QHUGmcrE8N9HDJ+pFPVJ5eJm5as1xYKHFM
2MawExshnCe2PbfFNpmQKGaGwUOMpS5CiNFdXXH1lEX81/DuQGtONP59uV3gjs5K
8QM82yx1bMu+V6JTVpKVNk5NNQa+MNhrRnkPk74WRmfTpRyh0J0uZbpVR2HJo8aL
PX5dD4j6V/UvGTR8nv/D2lRfVnuaSheEdy/yzfmtl9KZEQOwmKPWkR5clPnFWpgn
rBEd1P4JCFU9TxqeV1CeUvhCbzz3n9BI0YaIr8ZVoaIs9IMR+Tk73PtQjQIdniyR
vaE5Q89Op+3DbSXCo5Chq/ASNNYdrPRlGOWYYTgn+H/je4s7uI6WAIE1AzIPkbtt
S/iw7qLVJLUIphoqVQ0pcZ4xZABYai0fzEZtRPytf0BpdSvqFUzxwtakW6MQUi+K
ZAeIpAAVmwTQaVfRPPvzZoRAZJWhXoHCLDgOV0dyZ9EGm6zUy6FPE74zAqPytDh1
BfElVnQjW9OFosinIZqFxQ6mBR96Bc8spQljEocJGv+wsXQBeqeikwGeoyDmJtlx
PFZkCB1oz0ibJU9E44o5P+79JMIciFnJBZKju2mW1BFcIj0l32/gRajNqYatE3ad
6UORYklrBTA74Ia2MGRu0ziUFQYtpYEumdOX08iOqW4xIcBodH/2crVBG6pd6O89
XL69gPQcWgDXU4b5cH2IZMZpwSUGxY6DNv2d9jfVvX4d1QQKtjAj7qug7Fm8jxa5
IdqR3eJVZljZH5f7NoR4cOSGg1O5VJHD13JcTvjX7ri68ceKfWo5jFdmdPZQGH5Z
paA2xT4J4dnZtwVi7M1rUdoZYIKskHygVItm/5rGCmc5euwAcfhwIRZX+tDqMtjj
vwZR0JxB0iXc7PtPPIjmh7QUJR+7iXAWjiJ7bgywx2Zq7y5FzywRVEPRSSa8U46R
dUaCz2nLaiEp6S/cLqET5+Yd1p/7bcZcBMCuRVi3CyV1XkHbRHkki9MedTGQL0Bx
anOFo3ZdYNw4BTyiLa50EW0Q2wIP9OGeBpOdR/SJiFZ0CucUvttryAy2LSkD+BhJ
Cs2D8h0iqxQuFg9uytoyGrl/BuzKQVKBT1BJBCBRQSFJ2pxPhx6q+spTTowaUqFc
0snxZEoyChhKPEFHlOCcYDozPeW0giCLflbatlB6mVnODRiCJ2D5i3tbeWdWY9P6
9OdbQ/uVshEPJFOVs3fII7t6NWRB49WxANZ0sy9I5wLZoU/I1y7VF18DVOfsPA1k
eGBcbxsVqZYXCHWmd7+0xxFk38nVHT5aoRHiiar3xGcv+Yb17KLiaxyhYCOyqo9r
h3p2tbGK9O+vdORmPO4Dkl78eJpyEUK7DU5eyxM0iRuEgQpP6piR5EzbNgdIxCmi
rao9AlCCNMCmxUWiODgl7MMZteI8cFuzkMR1Sj7JXuWGMvLp+H3zi20/JiZBv7ec
EMPa20qPN6ykSl0YgU0E8e7XYGOlmmGoPbLR3rqmmFBV6cRfQ0xrIkJCtm5DNJvc
Rxgqh9h+xNsag3kEiEYY0wxIulaYClHEX4gkPEgfJYtDtb/cp+M+HWVSO6slx4d7
LR75/+brI31zokh1+ZN8n/evVRdl3kPs2T41xAhlNJVFmudyB+F9UsMD+Jdo+wN1
SsTyCHSeFWgGeWdZNBf3qi3YdWIwpgTEgA+XVeXn+//sqC/XhnOnBLXJihxfCTXK
yuqP0cvkxYdQhWtyonppgV46Vp7U6+6Jnb2Wys+JnuBPN6rjwVxwn6EE57Ndyk+9
RnYbK/K73ynJ0VD0c56s66bvCQbqU9ElTRbSPJ1gmR0pCk1lUBsLMJp6S2sMU/se
gtVvVtITfaq8EzbiTM5u4Tnd0pQynHYjPgl/n2fg8sWZAH/vkuzG9DeFfhbIjAkL
RmDmqedfu0Qr3QSZwZ2D0iucXoo0e6jhnmtxwybtGrXJNbHn9TLc+qTfcReuF28m
JeeRYTY/U/z/ys8lfz24Et5ZEwEpZQQhlt3j0BwnMjXshnF0wHtlFJw3H5Myk34q
X3fE5EJBaai3fapeph03p8yWlLyAl387TImVI69pXPYD8+AHyUvpky8HABJG8c4l
qsbZLHLAwHtvdXdpFNCBF6+fMfs3kczTsaTVPezwvU4Axxm/AsdschGIe5zWbhIg
IU9bMm2mEE5tfz/C+0paVstbJoUry5J8BluddsbeaiiL10ms0978uNLY8LUo3n4P
N0I9Rft/Aubya4XCLhL6AQEKFodVsqLymk2ORow/mvdr4i7nioQuwQ5wr/hsMCBA
GwhPE0B+D6O8O51DZccHqCgdxZVTs7zrg9pENndrZMyVN9SEQvjMydzLMD+tZLgM
CVI0T/cuxwPclqykPR3c6hFBGUzuQWAljmp5VtN+X+tvVz42UBYw2iCCYpHYTRNz
qUHw9Tq7nEjyGj5s1NhY4IVM7RIclCGaDch+pZDu5w1VrxmAn/52XjSm2+Kv7JbE
hpy1YVbfc2rEhL4Rai3yv2pP4p0NAu4yNnR4RnibiIYsWDS0hWKGPHiaobccQUZo
qMb192bNj0kWxcl3o8XRNHsfPGi9TALeXvwJkPJgbVZHU+6RFZyopxVkdVyUGwGI
zRT+fk7UotYasp7+Kw5rI4XPEDkewOK+K0lGIp0CLV4qXejBttOFHUugksTvl2fN
py4OihRBYSEVVd7QaEzQVPOQ+PP20PebV4shd4zdmzmMrzyV9Nc0kAUeFbLSWVUj
ZUXTjvFM7MhpPIPkga68DAqJF3xsNmkODUaRXGwnehh59f5osb2LowzLcLUuJHNA
czP7Fg9Uuo3JTSkQeRxzwNTbjAKvVKiW0BkSl6pWg1Nle5RoA9y5/jyKxDYb/pT5
wiKcTtMvtTI7XfVALTIUai928HHakcXTIH3aboyhCxhhhRyYDNXUfPYWWi6XJpIq
sWD7MIqoAot8LjMCfQ1ZF/VPm/YfiqP1FMm6FEsX7kumBZ1Eo4+g0Vz4/lOIJm8/
5OiAc95VdPuV3ggozpfDzf3H9Fu2pxvVOR/EHBUzROLFtzokFj0Sm2y8pl7r6bCz
9LlqthkEG3MY4quRgIwhtnCaTtL1xizcl7n3N+PYCnXCfZkcHQa9RfJF3uCljeoP
QlU0+OYd2YMULg9VLaWVPS9Arg7fv14ZLh6Qx6eZ77CL+Xl1/YsAs92I5Dj1uoYy
Kd+o7Z9893qMPZZZZ0dm4WBmAB42Hp3CkTQJ9DcKuVU8WefIYRCRdYoADbmeFobK
m804OSqF6rK+zzonbEOSaVPnVGvE1hcfh4tS9hP8+S0gsLaImX/W1lODPdENkMoF
w55p47dhjb0YpMUH9hmw5Nhs1rPoB0IZpALj0/4+gH3AuYba4V0jVMVA47bneh86
FvASHg3H4z3ZoBqpthfSOwXek+VTVTLdZq5KXyqlZc+QcOHs7SJop5WK96NaCHN8
AyTiszmM4Orvufy0MhD3S2nO32cskKnc9MVMZs/WxvJlcgfr/hSaLjY/YIzYyJDQ
OtsRq+ZxYUm67iJQNidoCs/Bv072G0UH5piiq5+yRZfPeSaWU0mrsiKW0p4QkVZZ
rjCFABMazXycGtmAq3pz7Sxs5gsvd7D7iP9YSAHx1R4/f26Oyyj8New7pd6vUWSi
KlGfqCMTK//QqjO3afxTpObYosexbRAAjOlt1Ii6GTlM51wlnNFGHwzlWOsjsvL8
gN9K94wQ1oZj2Xvx1KSIyz5UAtawutynhq8YFLIfZ2RFch2uegRhdigr5GZVKCj2
WbL3e5fzKlFROtPHGRoGmCXOHpOCqDcgNKqgN5Hv2Yp/cUaXhu9QD9Eiu7lB8Ypb
UUabxac3JqtYtZCMGWeBphUy8GFCORZiwDBo6XqbMQVABM3CcbSTgZaHsE8hktXy
gEVKBGIB/obVFaWm2y99j5xUTJQ75TYQuqQRFgY7ujAB6xjxXitx3fKtV8as/l3R
ey1TPSKuvw4/z9rP/4HlmfKlXFuRskYVV+zyOAE/dQB5LUpX7NAgnMvFDCbfbCPe
DPTJ46aBLTaUph9E6WmEwCKB3SexNJLzMdOEveOzWnGwObtfTY9OIhUHX9U3ZhWu
g6//z3toEA/NvGPIrcp/IG5++GWMjohpelkcCdbgZrafnek6L/7FSr2K5BLYcpjk
eOHD4KJX4MhM3OoZM3fDO7yERKxbf54L46gBFq5PEozkjI9bBiGn/qTz7/Pmtv0w
kXGgMKy5mpuetlq9pHjmygR2RFY49D/W6Fa49kv5oQ4BrQW4CUlPtq/XBNRutj1D
tyDOZvqW/4RjV13eXyRn39dMJoq0KB9/n99JkMPpY2kZMSrZWP+3qi4PJD7S6+cF
P5d7rB91eMx/EAptq4FvIm03RRW57zmiPhv5kCs+yLC8sJgcDTcI8w9Yxg/v5hZ4
gAk9G7LlswUjT66Cgs2E+zSALTu2rLdITkvvaHjs9Hs/YZujJInr3ITEPHC/1izp
makxWs4tCXJ/MVtCZ+H4EdR4UM5hzMBWcyyS3phYu9qri7y/fszgS5KPcf+7vHzK
jWPQZP25tq7I2P9RAs2ChagaSbhedo02Pzfh+jbWUhEw8xxWD3kWAdjlOzhK4zUV
dFW2wdMbsFGAULy6SOYKY0HyCTfeH4G+ak34Z4xk9pCzLo1PJ8q2gQ9ZIJCPX5fp
Gb4Wdgnn4tJRy3hgoTWEZF2ePtAoyLxHVZaem3PAlvhrZq91W8XZSg09lIEKWm0Y
xrhK39t99/b1xLfKi8ndPlnGX3KikhhJJF//tOBE7zAycoKdTrMtrZpRhXBzVZtz
xT3pOVW1dr1emFj/V3mtHTuU8oZprtx5uB0ULLlhNXpUChUEX1OfXIu6jGQwcoEU
pmazWeY5stUuqVkLpFkMHAzp155I5I2Rxlh+z1n57z3Hb416Nzlf1bed3L7/kw5v
JS/RDKcH+4zLNQtWH/La2LAg6AbidBdKzz/Ktq5UDx30YZuwOtCguwRZx98JSl/N
BQolHsalLSs/GXd4fOmPOa+7dENFvcG6+nf+kYrvrOXbGzmU/qTiAYd9EU7dKvQH
02VESTkaGQIW4RHRIyCIctSVX6yKLn17Hp5maxP5YPZievMinI4cCQavaMGyY0pz
GuHY8X64M8oGR8HXJM4j7ObfGINQazA3nlH/5M1wHKQmEcWvgs8WRMHy0JdhoYW+
0Fh9++oEdQC+JRIMLxvQkSBu9rwH27Baq2W0mVYeGqL9DCLDOQle+5Ak6s+AGL3O
QoiW74F5JTEyZrFH+E/pYIAb6Mfydj5b5a+TJd9tLHLmtOK5O9blHZcDwAFbswz9
dhFQFbNyqU1gnGoczzAti8CKLuZIRnfVrZiqEgItOkaqrEYxNY/ZmHHLNrs33ie7
ff19e4qqzaqaDh92Efj8DVRan8RrA7qn2WM/F9dw2oYHpli+k4pinV8CK1Dletns
j07Moh4X904z5yEqICXqmqInfkjFzNK9Ij/IKbcDCITZEcFCa1lsYJKw7c0/9Dn7
0ek4fzZBBe0M2tGFmZSFU0dcHSig5v7b7NHx9MD8hehXYWXat5e4u7SztrvpLPj1
+eoZx/ZPpx+otORWYUz0a0XX9l+2DkP37DSqaUGWklCdlmMgV/glZpUUtmuRckh4
8XFdhHCplxvZcNirAdi1w3ZoXU3ibvTl/cSf0xvuLaP4ocbI3hfZcOLUC8abxu+x
eGoMcuyhdbssDv7q//sYk/BdxAbAEsmagPmnAuDmiBvUZcQpL0G1afATUlYEH2tU
0+4PIxlVYrPtORLzCfHtbG1EksUn/k1NHTdruRkB9gVQEBa8jBC6Yr4n9K6PQ/Sx
DrfzudIK7krjaKKjYQFf/DEm5Ond8COxI8Bl938XvkmkoVAr0DMr5t9oAua+rJQd
pTyjRyGhvSqvawSy3Qyg9rr5yNfGxaereSBNC5e9auTGHse8vQQUVihlkuaBMSBF
M00rTn83iLy0tr03JmUOTdn5rWm9BS099kdwvZ3C5HS+9mUyCGE1N9xZ2H0c4o3d
H/D3KSShDr4S2sCSxpXKmejHOCmP4HiEyZChNyAPippAEmdJ5m88d+TWmRI/E2xb
2LovaK/fuzn7X8QXFLyt3dXe7pbE7PPpwYkk174VoC70g8hpX3jDeoasDM5ZpA8e
rOgxPQZObQzN5n3x64q0sp+iTWhnThQ9wXwo6ySjM1U0ARxCenOaJRex9j5DmKbz
lAc9mjsJCVHfQFUYNfFJMnNLNx6gGv/4mQ+yViygjuZoAdv5Oi/5lRxVb4tjrc8l
DDVlPjwc24HfpinRAD/oZCDG44+5LNynruCvi5QbZq7n85MNBW9xnERkMLTeUAON
HodvvRaXD8WaffJ4ccoXlYDS/1R1FD9PTqzbbHL3YyF8NqYI1iBBaXLOV5SI3FbZ
SILoRDJD87+cbICa+aBx5k+g0/MuBg9BVclKJs/DwBm2i+7AhS6v0rl7ngJESoyx
0AzXYDGlMbyri8B7Zaq43ovAHuLXfWXq3kvjGVcebecu6XiHsDhxXJeA+JlS7533
N+cBnHsrXqwlXnbDjd9K2SEvfWcEWQd0jbHywJeeo2PyoCIoh7c0loxxnrTD5/JJ
uwKvQ2Rq1m6SSdrkexpfc6x7taciw++PF4njOm7mFmBDxxNxjCuaPlMfcC6H/9SI
D+/VT3kzSLsV/ZtKF6m6QumZnwyiJUiHk6vL4Q4tMtRIJ4YvaSB4PO3vwD29+rx6
kjF1rzH8ZJ+4Qi+M3U6XhwGLqROObhixs9f0XoonngC9f4ojEWAgcw0/GI1Pe0Gi
29OBroKeBULR0tZ3C7nsPMKLHVXic6qK5NnYAMJZibbvrjT2cHSIsilhOeltpd+V
37bUeph1w6prOGorCMkHp0+6W3j7KHXYuPb1FMfH4ZPlv0gCRdezlkaYM8IVs9D7
GltMM0rAcNr8Sq2nsceap0BHIuL7HhRiqeegomtfAkQVpEsV7b6pjxhueWJcwoi9
EKMbAn1qvR+o7H8gFvrs/zQJWuosW8gw2xoxm1j4DRIHrXpL5F1yC4d/JPX3H9U6
4KKSWn/KEeH1lK0PzQQ5cQnqG1wipwk8HCQ98S5jI5m0JFj03+m5KZ2FxoitXDUX
7MXoHqBeRlHy1wFmq6Bj5Aoe5bRB1FbgcNDYXiYJBczM3rseDxweUI3v+hy89nOz
DYrLMlqbj5ZTcGHNn0oMqaN0gEPQX/bKCZrALvkrYUaJd9WQ4IdQTlkcm+1FroMe
gd0fo0kXobo77TKGLbrF9Rz9lR/90yEB9zNaW1Ai1B+G0TUimhmItGLeiQb4qdUA
srw4W15wVqBGK+SKLthA7GVACWhyekRB7dPUGdU8txjZTVZefPaCUzUEJbPcpVKi
aC5B3rf30QGGwbQEW9LF2Rdxi3EyG3SVH6DML59Ib+dSdSiOfbwvj6QPUrYOQ0GQ
avQfCh3uD/GzCX2qGZlDv3EuX6okANOtB/MSCwK3ZpDIBHVBd63WXSlJZFfJsUTl
rK5DuJVSqqV+wLKEYqCEPfZK5993+UR0EVTqpiaiYmDF8gZITiyhxxhdmvOuKiu3
tXfjGKHUTjwSLO4QlO9cP2DQvOCgzgbTxEZuZFbWnfiBjg8MBpQ/DSg+cnC0e26n
SzpJqQQHWdQxHjOVk1EWw72cCw2Ri9d1PgF7aq+DbJwj8HfU/OQaa6RSYQ+5iBAk
xMee8+0YERYuFmIfohdX1xRcvmB28Yh5pquh+VgJSEgtbqze/oP5P+JmxRRbL0L3
ZEH06XPbWDZ6BJ01AIriz9hCKyJkxCI0OCn2NhXo4q8NF0F7eCihCgQmPKZYFcgC
rTFSR0206vVUQT32NhcdA9RMEk8QW7drfcI0kHWNvy7UQQiPa/sgqyU4mB5grFDJ
dNq+slkwb0YfH6ypTURGk8h/4mP9sbP0zWPlEcLuLyz12R+QNUSACRVYFZEIxwHN
Y1buCj6p8Lp1gWzEi1gK2rZeFdtz79pPJHw6r1drWSKZRcJFLzR+0TRT6SLysugJ
6iUYXF1GVyduBv5Qbp3Cb0thVxl4I59oZ5VRonzWnbww8uWb72n7V5IyoFEGJteU
EFGI3ttNXTEc8DZ2x32JN6uTypYWHwtJk4R/zk/RVQlpR3oz837AEnDrGJQozbS0
92Wwn7IJQ2jiPDXluPWX4tH2vI/EPz+AcNRHLDBMErZsCNrlBqMK1WpQlfuT2xuc
FBg5SyVg4BQEeH8SaYLcL3qRX3xUBAWc/Fm8NDHzqBwbG588Xes16fXNlqdnCUSt
l3lOXqGEWMidLMuv2iAuTiNlfq7y15ewCne02FRD2IEju5bmgACgOKyspOZHVlcV
mY+xxJvRRPxd842umtuI/THnW2LBwYhM3Mfh9luts7K9O0LxLJQTum4VGpTMawO9
CZEUdo3JLZ7ntEXExyAzsjmpGT3Ui4DgZzp8XA6eSSGREVsf0pZQsT5Rb/GH56XB
DP7rKYTVew/FxZBRaYoij66jB8Q10kt4c6pGyhO51fGbaXxuYhP5baebkPJZ52gS
pbiRk81D6X6YA8xUsEggxSPcNPZiUbpaB/AVkUnaqqFJorMb1bvblgc2mGdYQlVz
h2QohEqq8bilN9TGpH8bScqvodiG1ygu4evJ4+j8ttZMyQAWJEgPd5xEgVDwypM9
iyQJG8nd1i3HHLVM+q7UFVxFP5fWQvPhLLDeiq2xfxa1h+IeL+gXKTX3k2rs0OtB
eV5LFL4CrQEuPCToicU5CX3jx1/CAx5b2syhlbLUyPBZoq11e/frC8nULkE258e1
e5F8S7qtvJvf5aZ83jRAcvXyAr8CMOQN8hKOoUwgILEesoGoVCBGjJ/6fUQTq5cb
la3scYsLmpSZNCElxnNqyrPqZ9RAa051iKjFpirFNyRUfK4xQiUT0IOR8tJ3HxNY
7YeQnsBj8Tt0HwfOaSMI3T7E3vBMm2IgcvCeSbTuq5Qe/91uIRI8Vy3tKGKh6YYc
EE9prclU0AEwFZvQN1s0WYI+HrOPevA9CwlBSLdDN8OCVIEoeJT2LtaFQTDPmR9p
kag+z1zW8aRmrSs6MBMAXz5oNwfCGkH8CiSlxJ+3Tnoh3aB70kVZI7MGHcfsNeXT
Nonxev2NSm7XQTFxRk4GKmlUxh7zQdtWoPfN0tUxE+RPMqQ71gQWF7xn60Vts4Hz
j+GdiULe2IMpq6knpybHivyLGtH3zrVTfv+cKgZX5SFLH/OW0KAypOVTJOUm1C0R
tEc+In6Kdz7B14EIeN9PQ+ISmJ1wQhFKDy7mOJJcuWn7OksAHYL6k2a8KVq/cSjD
NxaaVIYMrSQF+DbRWidmt7J98sBr3We02t9IOTlKyJkOaY1LJZacM8/DDFeQzZsH
fQQZXxzdVV2lxBCVfsY6ky7mh9bGZBEQ3GzjwqmiNHcqHzE0M2CAFEL6pG7/nbra
gweGLUeo06oI8eo6PRSuMRJj54coA4KnfxcxOXZW9WAUTKRz7GTNYmaTZ4yJlKhf
TbLfcGeg5Jm+REZR8zndQYiv4Cm6+HearDyxxduOmitI1qJ53PxGAWR6I3KCYVpa
TbafhJAFR1Vma0472ebZcR+mGeM8eS8Ac2L4V3jGgxBpM7QkZW6lN11jWgryL+tX
yb/3qYKLUvNAZZRgDZIqqIP7GpIR5E5cQKaJMkkQHOUIks2UOxUfwmBjRJYAlwUp
+h3UyBC5t+JSFq4VahkWo5tyZG+OSKasIHusZStYGrPTdwZhmnV95wAnmfwmP5eg
yxWv5tH9th0UbwaL8d776XobF47/duNomp/OB5iGgAAanRdRfv2VbP8Y+xlUW/Xs
rzFAsBph/pNwXBDdJuh8807PnwN+5j/CN0ys0gDe7OMQW6b7tpmDO1JZEo7ws3ZM
zHxJ3lhjQ3mEj0c4LvKuozNdGCHGXKNG2+GqPGNWrb9ed2smJERPqEm/iT8gJIWY
/i21glT9MEL8IT754tw0XhuW/3FBGeRVT46mLaE+HzgFZZsOYYhTINUk3AQhELgE
llKaUYfbdAtg9tJVh0IjthJll/8wvZigUVXufYiLzl+phUFo+TeKeJ6NMTcFJbm2
Bq0IuI8kBchicRyjxnUl3GiC06IP+WfJm4prypzhQLnXGdG2nFhaOCw8hXfq5gZh
1GA8EXvDYIZTyypf0CaGdBog4pBBsOcKwfPMX8GTPJEmP8Kvl1XJH8jJanZm3Nps
ZRYd4mC+br0hRy24pvmPLzWs8K5fWVGvbSoLTucYNtf9RxMGuis4JZ9ltKs6vKAv
o7WJeVNP15dXx94cIOH7qgXjPo72jz83FmLPmCZBgmjgM7cZLVJWxMbXu7krbVU7
PuEZSsRD4Hg5e2UkgSwmaZPlYMkwUeUIZAL4l6biYy83JlXR6uA7scYGB9E+SaWh
mos2gcUJciNDm7Mpfcx04o/NgHMvdtqKsgLsucwgRbLIxYVZ8bQYfKM9tYGSvtij
izM3xLNgV9kljLyrThlk05Kahl0vpb+OtXGWnIwwuNZn89mxQS2uNmvuBgmhFx2h
0kwE2E1xDDu5keGJ2u8oln3r1xqNhXN5P2DC1eRu5OmKBA7KpI39X1nLQNUkCBjG
UMdN3pVs917wXmrBPuB8uV0Kvq7MO0g0DbGjTreJFueQatayWBHXJE7MdBjLH+BD
o0lXt8SQq0QbpOrM6/cVuVOZ0a6MElr7b915rIC6RvCeQxwDnjVM4l4Q3Ln2MIhI
yVk2TAdHIyuyIJFkemaQBY1w+F2MkCHaWWjz8B21o2seZT9RhqFKB6U1cXkcph4w
QNAsn/se+JeMslqoXyCRIhAsyCpoFjwH9s9nJubD3fkUFA+WeywTbKdwbsKiZ2Cs
ja2mN/xKVkSQb8PXpDty59xe7OnI7bqWFk2JW/HRrA4qremK9wnQDJKMXx526Plr
Pnwsf6eRV5IRzcENo0B1ErYgWk5bqZ2ogHXFtKeQLTxNkTmS4IniYVUNZwQNYXXM
mbTr7OqPtY38Ynbr8c0E/9mYndOzxu9TePZTMDZQAbZNabv4/7+RUjNkUOO5xHac
XS1qki2Gf0u8kEu6899UWbEDkPwVFDCasx57sMUariOMPUBErOtFbdLLpCUi/V1K
t71ZK+o6or2vXrCLpbNFpWuB9QlHVKQBgzAQauf5VOyhOvFZvy1bfKw8un7FGTfj
GtraVzZ+cBaW3E2IuYNgkjYqcncF+UVkUxoLunLkIdVJYp7tNGjAzXX4hd4V2ia1
bfsp79N0BDGILTuypwLnO/lv5JlpENETIn40N0kpRO4dRQju7eBVW6ZTQ7tzLacm
JsyT5yDV373pSkrCPgUrKNWvnpPkCTeSDquTQjuloWbBN9fi2iRBM2kblOwSLo21
fWq/vuK8gi0dLHgfpWaQfxzmNF29utUWrt0JqHOY72jLwYiFVVdfhfF0+n3NNtDn
VXlbsM5YoJM4qC6NlL7bQTSdOYetExzeQ/80IUXlVsAXecSzK0dXRCtf27isGGLe
viG5byNyirmLYlluUrSe0aSFVt8Fr6V+tV12J/0cqy+iRQljIO6cyRbpIM2mGlNB
+DCDDQexGzcFSObx8Zwzl7+9HflMLMLJAO7KYdquV345vV0i6au5zTAxCMCn5ELp
LdHVjEQl3dyfmxnZzLz7BKp2PYfjM+rLyGjMrWQ+d8GNrUAGRaK2/CExOZU4nHRF
ttoO6YQ70TIaSWeK+rrOUGQfGpG5IVjPMy4LcZIz30L5dXlZ5ew5BDBzh2gm5UbJ
EkFngdDhgPLkqKilALf8F3bwlDWYSXSYqJipkBm99Gc4Xs0ZBlEI7w+7IFVbCDdc
eb9y6CH22AB8EVH1QBbDrvF8OiP8+xX9N7ljq2Jfw3Fa6EVt/iL4v5LZCT5AaGCG
Ls48mRzLxPCzYt7AsKUp3TLGDUzL2pXsbljS3jXBD2/OX/ljMeH6DZysv22/+Y5I
YOx8rO3Z/afIChH4mI1zJpFWemEeLtK/gon/lkfU61hFkvraSW7vVZrqAaALNNwf
ml5UcTz5YTxqNNtdEqcJ+ItzzoohT64j02nsESuDs5m9ONwQJI9o8pkiTwrlrcss
33pVrEognVNs88Ore+2tBJqTEoOxMHgyyY6pt+mblNy9zy8EhxcWJE/RWHxNruuc
e9lPdVEGUmSD9G51+bG3tn+pbydtihJIslbYkohQm9kAFWadg//AwHM7ZlEMBy1J
y/XVNSgCr4b78n5atUw3h1oNdPslhXXi8zYEQidRFlgUCut/ruaXzbFUpCIwVV0h
90EfgxcVzCZCT862s/yqDyP//SMf6QSk+eGdgNyPuafM60V3veGNMRo2T+rN2ZzD
nwFHI91f7F87U3msQ2BDOgyV13h0zCZYOxuaezFUCObSCZhMCFAqBPhsbBYD04eb
caQX7e7I4jgj07Ev6ozjg4pv730IJ1hx28uvcjEzdn73YNg8nGEYZq+Lo5vscxoo
34U+5qapRPGl4UWrn2CZOc2TF0wYbTt0SiIqv+4YFa0fUPsuHug+y6YwX0ag7NZ5
6HSRouJhixvxa9JodsMIYTDjJmsCRP4wifnD/u9DEn+TyHw61ZH8irm6mkk8BFbl
hu/U1z+pDZBzc2ovQUGgDxvi2ly7QLaQWbsqiajppbmbUIhkYT4GNo6BWx3ssAas
ZcgXs4P2ddLXGS9ilpyZQFKp4uDDoivVTFkycchX+Kbohv479d3rwbSxsAwM//dT
iQ7rz0+GOb9DvIslcP3s/IWCQJvnAZVGALAtTkvohcvg5Zte27ERqqxaWJ6Adica
WIhmXvN5jyUFwzQTWcWOEG8kCnwne0EbRpLGnMVE7xUMqxejimXhl58EiuzX/GVq
KK5/GWEqcLbCG2smyJWcx9+e/NgM69zvqmaWLkezw6B62MwbK/lSpi31mrx6hKPf
2Y/5ykm81LUwSPCH4L6niEcRgKGf9BK3YEKpkAevXYIJic3lmxPCYgDp5ZUjHWo/
74JlwKv5+VMNxK7l2mUNFCxhT5+VBAFLljlxvqGnfe01xxZm6tq6/O2opy38ABUC
9qSy/KM3tcTYowN7CIugddvZNDloRP5ZngKmd8XsJJqv3FWQAkWcttEzY72IINiD
VqU5zAW8sXKuocMvSIwi8egGJM4cfn1Xfyern60lqZObYm446JX8zTTcAJ4FENRR
DpZ2YR5NeegFfqneYdxjtWRsnTtzv93UhxSfDA8BRtP8FOytnKriLA0tnpyH9Thc
qP+Oqfi2IleUrjvtV/keV25G29nIIR9h4sjL/2feVY+sIDrI3GZcmS4o2BKp6t4y
Z1qrBAe11UdWg3O5ZwXnb/LmqyRnJKVswcAZKhNptzFv7lhMCcrBwwAPhpaf7aPJ
MKZDi5z4WBE7ZG37JyD8Be4spL96/Dh6d8O7KBMGsXyiiZqHJKqoKc5ps09LYE9I
ZlPSQasjK2TZSfTyPSiNQ30KnqlcsMD8NiCaeEvIuYbBARYGygWS74KzvBVP1H72
QDKk10izbrBg/AKPvTLGrnUnWeyTjZwkqzu/CONj0oJHbP0EcmeGyj92HymmYOTS
kpu2QKwGekm2ynDNpltG41Q1AIfgXd54l25ZXn/R/8Td89HnSab030205hYdDujL
PCVmnOcX/ArdTPTsMdMBn8MqQhxbVCniytAJH69U5WHoBk8GSBuPQUIR/WNkvGdp
3j0LakkiupEdwcjlksfnqTQfta/7JfQZKjINuY2dlYPVuoF2emN6TMgiuy2KJOnz
tf9LKVEl3RUD0T3lABg3HMQY6x6naOSjnlu3iurgSUYLPN9TkGDGYppZ9xRkuJjP
eVN7bnJCrvy4pjTQqkuzToCmnweiOD5Nh4ol0aDrOew56AQkzH9EfFsts4ARdoC/
5r4eVC9kG5mdotZdsfGLwTe1oU9GLID0gp39EVz50YrVdeVSbkO1DDz4whVsvjS2
DA1/OqleMoa3R5psyTyNekLf/qb37k3zQrKsO2XTT3pRy70bDjW42/cBe+V2jW9y
5TCvZCtrJaoDZdlO81UlztP79VgWopfXSNA2K9QBDUOD41dL85KKec0v4QWCacsF
lV/ZAkpJXR8SQPHtkS5fGmhPn3V+kLOhBDC0YY+/0ltZfTBihGMKE0FwLgIeQen4
qDmNlH87nWc5pQSXYvc89WNpFGmsCTR9967uS3xz/qypKdIsTXyL/IQ5fhdNenKQ
M4+EjKj+tln9LxqmBMpzF3ZeJY2gE6nY+fgzSYKDVSMTyoM/59H8AwBtSZciDJux
K425dL+vnl11dw1dTBCLbXqIMgUg3OyMHcmMvz7mMRaLFth4BBXrzQsfCW94Q7NK
QqVgcRzjtnZFZaCRZNmNEgI4LkR5gZvjVapuxgPW7P9ThUGfmsEavEA5I1b5ClxN
u7ouwUdfZFivt5VfCweevvEAa4+WgrOHGl8m1ag2tCc3PFYkV7BZgCNxBhHCKYC7
vUPR7E0GCx/K+UrQHXknl3OY2FbagEsiog/xlm8833LxzP8XQdFHigMXuvvOx+tb
rhbjvuUf6463qRIms5C3gYXPunQS/8Sct+D1GfaX8gPUylKEaKg0Ax/Ukr8Ysco6
GwO9ND/nZlhwIM3nbp7N7eXZO6nxgnq1lQ0rsTJMFea4nbbDwLam6jpHK9lo/BL3
bs1xoVy2eaAA9OPB1nuIDsRS+qWwV5YLOl6LBDnIZJN0iOpENu4ZWLcIhe92fTkB
Js6btXgtJupMdq+ioB4R02fe9Hfn3F1CpB+G/+eeu5VDXj8ecw1dLwd0ApzIRUTl
7Dm5LP5x1sg/wR7Cq36DKGEYgYJqA+UGM7qswBctzyQ+5AX/2NpAWSynBA8YviIo
OIdpSRA0aCZiGxZzn3v63F9/7bxKzbuoyh4XDUekjZY6U9Uyzg5aZf0dWzpKMt1l
huspTh4aRWcztc1skJvfeVKM8NZnjyYHEqTWea65iWznLV3y6g+zZbXp8v/bKqFo
U+XsDwSCePyMOxCPEitV867pCtmAZ5AlGzkF362Y4Snh7NwackgZBQJ4e2HJfuWh
FLHAc/FB7j41g5TicUxdr8XHO1kXwXorkHaH2TzeSO3FN8rvY6wWVmmqH4wbAIG2
53vw6S+mp8fLj3DVee+QhnLvuqmhpHMm/GdDnMuxLYv70HoWuk4KVVv0zVnhZYb/
t5h3koUKEjLVEdgCfetWNBs7MjCNTMMrCLYYowshr+eA4B5NQF8K+2ha3728IsS1
xxoq31Kd2XvrJfrBicV/pkE4UbS6KmbNKs2RPF9mmuVrRrJdssCS0FEBfsQ6M1Hc
m2OtYAJK8GcPYFgl9QzxyFdc/o1PpmDx67+KqGf2Xt6hpoyhc16Uen1myk/MdyGw
MhUaisxWdKnpuJ9f5d0bGSlQnT/Y3e+O2jxA21S2GgtBXkMp6LoYRTRSuqmy/ZHn
TTusc3XUYs3n1bavWtblUY4xeaUeTN7mT68w7doqUif4MyaKl1JdVubqmzNe+E18
Tza+SMJmX1RDrdcH+Eai+2Hiozz9shXfiia0FQilTmxtY48GEPcWYkX/gB0NJ3c+
WW//uzjzEIeYJOmu5nuZfG6JGxhLIzVWUhLVXUhAJOz+iVix5FXCYrRoGZecJky2
obbZ+32HJQgwZ+SR5EL7E+8cQdQSzTOg80+3A9DJm862QcP2k0d6bSuP+kBju8s3
23T/55+1PubWT4ppc5yAW1JbmHKVzXXGYslQc594jyF98yzxwYTeEO5w09NF4At2
XSSGcKMeVSlFluIXFuCTOwhCRVGSs5AYXIhBPfQJWFwtvfRSRFb4SeXX9dq693HE
HRi2Qe60uv1tdG1dgkJCoHqsLmiOCrVW4ErKB1deZdgjLtMGY7mMuSS2TKKlE0aq
nmMX/oHIkIusUq4yLTkwm/Rg9M9haFRoRzIrRBG2s2ACfRMPdLXxZigbPTuhgrAn
5AEtb8ButG8ehEUgNTi/vEf8KB2MqWEGCSnXlo5MVSawb1iiYCBsKCcMIP2WHeJT
SVrm01NJn3XFWntxxSH1Hky5ZjMNElmd0YndpB25T27g5xbN0xSBivs/jEwK432L
NVRINfCK4dpvzcgMZ+A2amdPcOuc2Kell7nwYhukU0zbTXgKhSgQ0eFmrxyKryh/
PGDU/NJ7q5/D5zsihC81PKjnIPYandp4iSgd1+hrrZAbbQMqhi511F96FPHAl84Y
QBmgWCzNCJlkPGv6+f7pOspfVhODXltNmWZZE4nk4J9VMQO0936YGa1N2pKy7ywy
XjqlOALGbRYl6PxVaot212nrhlTYYWAkYJjEvw+kmrU50HS6mt7OgCvgADFc4zBq
yY33+d9xFVjQPbpLXDBND4M6JfDDoPAO257R67TNu5n72NEzldxcslT/wFMi/d51
p1MMCnf1dJUJGyYEzA7cmjFqUyJstVeh2sPpMw6Cqknl359zsWfTK31jDeFK5qYl
G3bOBO/EiJYV4m7PYHXm7Av+rF4hsxTBdjj7CkE2sL5Cb2ck06mprAl55gRVjkgN
GSoEJ0SLENc5cwMUXkjeuSa/vXnPduqVtyzvvDT+/OQ/Bqs8uOTam/roGotFPANC
ssacPaMsi3qqNH1t/0BjtHBlihDqlxOKQ5sjPWktJPF1cABtghEfMMXIdmEtp+JQ
6ObRuQvpVHKLzwnCnmt3eGaZ/WXvAm9ipUHQ9P8c+6eIM/ja0gW5XvPeh4PZ82mJ
VE7+In1Oqq7NgVHKjtHDd3Pds47oteVB1TuORPWEYawE77oB5ExON8vASTm7c7eI
VbHGzeH3zL/1Ax5CZkBxM7+7JKls2pd0Vv74wJDJJ6S9zVMKXizKBPOJc5nW9Rfw
BFfLhW6InwatjfkxHCY+ruQIlEBGTVr/VPyvLyIG9p1t3l1XSHHJudjwC8r5Qg5/
8JeZSQse/T2krJ0ZiTwo9c+nRA7T7E3HdKnam9uAwLCturcySDhcHfXV3il7kLPK
xscdVUxlpi1/PGNBIEz9Xf9QMIZhveKWji7Fk2gBqA3q6jt5inoePFIZBq5wtHsh
wmVc3OH+eqJv3XLv2vupuyhy4z1hdPW/CRjzHED4RSVVr3kDq+oOTjOTfLwmj9QA
/fnnjMzCZql1/KpmJPR+ymtqUjGpURBGFmLV1OqHcr1YQjWzfIA5mmxniCCcUWlO
PADflwiAKqyhdi284yuP8Yy934e/yCc6x7VpQrCNadGcMOKuHU0e/cnLMKFqn7Aq
WJPdDSX20j5QDLPrHKeMM8puJAyPoFnUKq6YQWaiMQ1jAK4pXHDQYgKFaDYh7vB9
mGuAdCP35Ay+s1Wy7Rf7er2u1nEgr4CZnhm8kYyG3aeF61TfFIRG8lH6LLUdS7Dy
3DeSfG4FGiKsnHNKnetwuIsXFXV02ioXElW6g2CJ6zDsAIOpoWL15HOwcEaACeOK
130MInp4EzC3jr5Ou7+jR8NnsfV780U2AJRxdTOgmrhT+XLJuCS7Lexub89Bwmtj
ouSHtG9UaP2K0SBbQXLEm6en2K/ipYaQcCOQZJO8x4ALRpnu1fFm8gk+nqhCYBFa
RQAxmQ7q6PFd8QXJbF4/EW1bS+Ro8TitVbpQvQRhPd7kXvYF+eoSaXyB2HhNcOZE
gkHYI1ZV27wEAM6zI2DFSeMIO5aW9KE9i4lFrnYiixZREzcqxWqCUYaepsEFeAhl
yxEoRSN1O64WmsmpozH/xG+BURHjF1FNgvwfu0qpVfJCJ+Wjq7abj3NzsX9j7SVx
fVagUi4ap1kCetCAd1Q2xdH6cj05Vgy8lgC4WAMtdm0Sq9YSNKzsAC66j9+dNYWr
iurPFrjP7zZdRiiHFh/0NT3CQRtPGcXB49K+fAXqNu3YUMqO7JdYy0IQo/lCIl38
J8c5EXuPd3C+CpoicJiJkUcLE4LP2tGHDbFXwq6L1+pSZjCE1JA0jPaehzRv0VaY
sSq6fkU/t1X93DSwMMOr9woPUQ6a1wnpVZW/VAYGwNqHfQoPNlMNt/ZW5/qkn+Ae
wuiCqm1dj/Zif+N9TXWCiVjKFV2vrGvE7430OZidCeIvjuLOltx0DfcdU9u/n8Kh
iXwOFiqpRpfEwgUcfvCIFoxp+vk5B7rYAe2uNJ+zBFH0op1Epyjkw/BijOcZkZlM
IFQy2wZTMIw+456dpfGvIQyvHs7IugUYVT6tyFfy0txSaNA9ChdBcND9KOpbPiPr
MJ+k2YpQFOPN6vbQS79xK04+mXecqHV8qFP2uaol7ezG4rWaWdJpPUmNkcYOUxza
vd9SGft1q90PfOlZcmO7VIPgr4wFUqaGKVzpjSYla6/7zPgSvcHQlxqI20U1Fna0
i3xjdI8vrRPf9qTkQCck3+fvPCbc/B3rMLrgzxWs2LYGBifZ8fpwlYGyJ7holdoI
MRk7jSA91Un/mqVxM3VADiNUHNxYyYNITXj95b1ppFZPqSXeVAwl0VUfIgAlRZL2
UbPRTaPYa0QjnvjF6PDB23jXnd/eR6/0r2L+ajwYPR8ShKKXoy9HTPMUfen540j8
w6jglaMeLItlY4v4hevhdQ923HZkwqWavHb8xEpYq0c29+2+tTW/mAymQBmInN40
Ys6OCYSYl7pemYguC179QRXye8mstSuKph23BNWj5lTAEweec3/Z8y6QYum4wsho
NLv4in44E9kSy9LPiE1H3Yct2zglioK5OnmxEOP+1SvmAZkfV77gkbRuscY4Ce7j
ITyKh4nq6qW5joL014kGJg/ckOywgNQZC17MLNy6RUhfcM3n8OkDsz4BC2y0P64J
sxmpwxT8XSE7YnAku0xhE11m04glapqXZxLlVm41TgQYIwcX36B5UJRDY2lQvGVA
+5oznjGIeKB1xC4SXbXUDrRojhD/m/Wr5WMU7G2XPqw//VF96kcUyjpRbGOEeXIx
U3VOtur2pQxabBwkjeW1RLseKGS+tThCEUwIacgtmo2sIdy6IFzdXEKdwdevuKfm
z5vPZ/nGfcWcZ3MEaWGb/ejIlHjcRoMOBAgbQEs3it7Aq9N7tQ/rylVa9or3lruU
gPrb7I9jB52fD4kltrc3+EcTnIfiEFRBYmZ5Sb7aK5hK14gVTAp7F+AWyt83gz7F
DlVF8z8cu+Yp+a0tLcm0UPXGrD5bZlzgMjtmGymdnzt16nIfJtzig99YyZzOZiIF
aialMlTc/0s8VuEyICIXg9CbdIljapyK7yT/uXxxLV9YCPzyvfA32WjA5ZHWx8jr
THekyIK8rxOvUrDsJLVl/2T3cifrFRAQ+ZzFMDqAeWicILL+Svouv7gBqGBVRdx9
lYCv8l5G33RvYQsrtEfSLhDBY33Pt2CnvQjMi2TY/tfm9hd03vxlv54nkPM5ec5Y
DHQ0G5pbh6cPiN0yqNyQF48xujEJhUapDLHmyTHGUY7bLIx8WHOTt/bGGrALTD4o
25DV5tVqKN8OqLIf0mPXS7DrZMozgDeRtPV+FZHnC2qYcS3mnOay91iIMdVAE3im
5wukMoLv2J0rFPzdPa/LTIxI0rIoD1wyGj3tfh2SXiaEE3auRJPjviDCdmlje+Gd
8GArZg3CzaiFyqJXlURMQhdqZBBGMX+QTggXBDA4nOhL7/6N7XtBU/HQnrWHklKU
LxH/m2+P+f6YTQHGbWIr98k9iVKS294BX8dG3RA9k5dHfG9zEVkPtcSQsiRmyUCY
dXb4lSmzA0dy//AIPrnVkYlwk1dOTWjRCyfhNmdsxupcsARvqjsnj8teXGpCsUwx
UCe3FO/dsR2ziSYThTkpIu8XakOc7OfBtwJSeIlxbKyI+eHobrym09/c/zkrCkVx
IPGFsnkMoTRrd2cDNqiamMCAQLKnos50LD9Pwrt6QoFhmSzOnOLRuxEpl6gGcfYW
YJLbR2PZOH6/lN6CclksFN61UpBb1o8piZduUgVNO9C3WsxDLRFy4htayUREpCwn
qG+O/BlZ0YXkE40/xt0IxpVNS/U6drJS3/6Oafk8GTNa7I3xOcKWrH2YFq2DuuXp
P3zy8srT/HGujJBEZy+xyEi++PYk1VBOPKV8XPTuchO6C7ujJ/BOLKHzFBzuIazw
3LyO/bGybjbsc1SOBzZJ3yL2vTIi9s2XbTcde8cIYLa21tItRMduHaBrs8qKM9+p
Jrq4pIl5zMkefD9IyY3rYIiIiEbnX8InvFcinn52LUdeHUEWdlheUq6B4gQThVeo
AJidhe32GWzZL4TbCdhrpbi4E3S6C/c2jkaMs6/B4ChLac4WsggwsnbDaaBqYRI9
9NlFauLnBNBOl6vA1U+3MtpL17eg/LbyHxmc191tL9AlvabvtZYUFgjenqL7zf/Z
aauXyVedanhlbcYms/M9ZbA08GeWluTqMOXsrxM1LTvt2SUWSas084Y23ALgXhMO
xy0us+iTHbG42COX43gVnf2bksMSReXh7xQLy0tJEbyWgeOg6QuwuPHSz6A89a96
aQ8auuiIQC4YYw2/174iEHccUvkAIGObQkb6OfbMo8IUXcLNIJOKVCefyzvaGMoF
DRpvpKb/XUUtvkIyG6LWOfNEs6AiwtX/lpVsWxVdQS7zk1sbXBlX16cPqUNF+chH
UIMk71N1n7bAkhz7hZ/ceaa9X2BWGtFx4WK8sD1nKNIJokkhV87f0Z8QAYGl2LWs
mv/h17Tl5+cjdpESP6jRwWDQ4IZ8D+uSAZm9QiX8IblJX4fGFPxootiQnfEHkI//
xgU7VOsEYxH1SPnSdlGZ8m+suywvw6p2I0ftzYU4/KcrMEwP7nu39rqVbBSaEJDZ
ju0RmtaUbiVXZboa+bZiTlY5MDC7+ArfQw+8FXUP/js6yr6DAdeimGFHm8RF2cKB
5k8TrN3azI+0Eq4xY6NLZefaY0JzbFunPYV/cOfuYuoz9J+ubhK33K0DwylL9kpj
KCmMwz9BcdjoAN8y9EB69j4Yb55qnj3hjQIFO+EpKbvr+xa8f7Fx8twqIO+qGnI/
xhraj2oa7QJ/osy7+KPX4Gxtj0izali+BqnrG/NP4pbmUcMhMoWH3RpsCxf9mW7p
g4XDXROYsO22fYKqJUImzAkgmquqOpk8OXkvpj7+pQwsIsj8R7wOZacuVdnDa8Fc
HxHeTfAEFmRC3lJpWFycUylMIuPb8dD3AZTC45dFyRaXSNsp66E5yGlJQ7XQfANI
oWZDa49eC9OW9v8/asEbredH2GN74dHOOF5oovcw1Pt9a7i6v71Br937NGngoUGV
PmNN55t6Eh/0pLrxX/HW9ZESRXiNZE31VnzrnaGmY4mgjiRvTx2bbxoble03kEy1
RH/EY8IFG7MmHD5BqPhr5sz8hp+peCnxCPm+9yO2zqPdXcfG+kLPqjEI/JwSM/xW
j59uyi8mTTxo1ao5T9CV/6birO4jIpvwelj/sqikUsmGl1hI92zIRgBKFm9WgOcM
kfLqKYanyKRLp7DeiiWMWhWfLXh1qP8bMzfqE6OXcNBxNW5AQBc4wgGVW7GwXbpR
QGyW30g0kTkB/4REmegpKNn3DickGTHTtTlx7jaUwwv8VT933gH8AtARdT1CS5h/
h8NXNnQ2qNldxgpj3df3+gLOeppzfmkMWgU3EymqCc8azDXyfQSZuCVpPSmtFbAV
Y+NgY2sgy5PGeqUWe2Pvg3FaZw7+D5GT7Fs96ZWWDjFyEueiRIyL64Vvup0jhxkS
V1qp4JDzJC2DFYbON31OIyxh9y9rA1nV58Gq9YUr63DZMIqw9EZkRAR+0g7b7kkE
3zXy9VyP2x4A9BDS0876OfOuBqeB3fz/4TA4ijkKj9KeXt8W8h93JkB6i6jBRugF
6jbEsSRI33NMFYKHaOYVfmIrnOUqasXBQy4AjVOPkTUaKW/trCzyXXbU7M5oNNmJ
//ru5AtooJlw24gof0N3BN8zxcWCXty/KHrcA7KX68RzJhZ4EpGaoIq8z9ciuVB2
yjG+OKgsBuc06jG4YWr9JQH1JnkqjWQjmByEfMs2cBhPA8gQbGrzlu1+6mBZA5PZ
AsEFTmVQuGOWc3WoxVwa5wCcv3iMRjSa+Sf3o3rTiQrhAi4gMtAl5BDAFyYXWN+N
vglZkBdyLoiuhTEYJ707WdBc3s6NZ2SRMWxmx0VLktkMKEYFxF88ESMsG2WzVIvy
XMget7pa5fSYbQTAOgLDf1XrqKhgqegDbWyWvFVRv4TNl/uMIsq1GUx7kCKVbDqX
BGFjtGff/xvaIr6HNz/C451mch7H/VpqG0dm90XTS9jyn7hU4cWFo/iweDz5o0P/
YPKMdbk9WBxt3LXa+SH69r10JpkRPunaYTiZ3XDbmf7kT2LaXAY9CDfg0rrXBrte
QrLosAiBqBlpQfqOqvhfx6zf78WFOmOLURiWnE02EO893Bwk1ejCAjJn/iWShyyk
Ux95piqo8mZtajCOaqFfzWkBV8DWD9Os1uBKiNgVeQ80XEsjoxouARZrcdi+2xL2
qKV860pJYiSxxvFByJgM+kYCJqfr9cFwCLVjenQ8IU9LkF55+yjJygKCv3a/7WX9
9NEM+nPOz3DV/+LUWz6zE/tnwOq2GSsBxPOshx6jZnf5heSH4jU5UVXhLqfiUseu
RmspEq4LK/PPlG2M0kMZu1XUSrzSCmYI9vTeN90eQNnNhW3oDcrE71Fg8F/E4+B4
xaYJQj6Hp/gypBP1JwtNk4Zqjb6rjMLTHxWp/kXURFefzd8hYS6UlAkkyi2nunKx
+hneSG73oCkBL3I1Ig59QoxvuRr8z9BqIdD1cySt53BglMgPiQHw3X7kjAdoeAgE
XRFd7a3GuNLxRU5DRMoxkvoqBk64IrVsu7Lcbwy0LMa2bYE+tIvjGhel4n87nb2R
FjJdb02Z0hqMXu3XmTRWcv3tPzwemtIHmDsIySU8TqnomW1kVZUjBqeK0AFYkqTw
u+/RzVXesC+VFkvYW1w6xpL9KY44ndpvQBfihQ9Zj7cAz/cFqbBeDgWjEEdv64Um
fheUjBexWgvulfrVcazAvenDFxutP2Ne8Ygstl1BMRKej8phqEOmwSppyJiXwB1l
KBBnJASh6+E/evAIOyCRDvtxJi7KF31RrvLTq7ecEDRtCAHbc9n463ax8Np07HoR
Fa4O/s1IBEJR9We80vPX2y9WmiPbojafDYE25Z9TlvsbHrJ/NZg/GHeT1ePlyD9Z
9WsjUlr0liiPeDQj/40WyKvXKZyXlMf5M7BErisguU56IW52IxYEXDVYuHqzxfX7
TJADE1kGD5U/uTeeAbYoxHOmqiMbd5H7OARbDhUn5YQwmZtOSZASC4Mh9nCaVmFC
VqA0zykkJlebtVX40fAsHrv2qIL7eJFVNJZAv3UzUXT3ygKIK5SnohnX9ilWNt65
fJVCE2hkbH7uPoX8XicHYvVYDNgtHb/wIqBCNk0lgT1iOWz9vhwlZ4gCk8nLM4kM
JZT0sR5IDVs2RapI/p7Ydq7ByxgliGTMFjMSj6lp2tvEq7n0XV4lL7rByoTy00v8
iEN9hckfH3wbRU0k/3L8NLYq0ZXIML+rJxGjBpCIyhqDtCfSzx9uOGAgIg5R8ZAg
crd02sHK4SpfY/ioCmM6JgBJCvF7zKOrenYNr10ZrS+1i9OBtXogwZb/5hwknFa+
RTfR5VdHPFLmsEeBQRgJuZ6LFP0yypcGipnZJ46q39sG7nPMkwmjhAGIQ5jWjSeU
9NZJdO1YqfJfHpZjiBuvqm5Inl9ZgmUo63bQL+dSt9IspIDhdan84WmVmfJwhbAY
+U6D8kGH5ZRm4Q9ELEerEUAiYJtuFf0xeqWzhs/4/ydLwp7llDp0R0agdz4vhpzQ
DhlKGa9B7F7/IEuTmps/gBtnQ/AYO9t52BTV9daBprPINsbjAZrtLQB3MvgnNwYo
LudD0hPMdA1pHCuuMjdSZBJUVw10+uJSnWOdvvo8ag9AecMMujQjgXruhLF+DgVq
uK0YosEN+woS1HpNa3pgwiX1JgX6Ntil9y+ILNghu/3VFeJ0E+6tKDOEgrj/+XYK
/k22fWsu1xSE5PWpzVQvYSXwpI5NHcyA3G1Y5g26c56t5rPBKke/tLin0RbT41Ky
3aKZOlGpfiHCqwV/uPdGQpYpnT9esn3dDlugElyqg8LV4UNCQO3YEowOQU+sbZrY
NbCKa9WLFWCrexmUeA2T6ORaxyBeC1K350Z5L7B9fAU5kvjMaZm9stLMbQUaRmaG
OqtQcLYqzcFl4yhVgfCfNX+db31D/ni/NVKE0LDkxTTQuRV97y/3/bh3FMQKrP6N
RKk/7hbmHdHkWVOgeCItzUJ3xfphsmFHfPebfEWiVNMAH1tDgJJbraw1zi3bw56b
KZ6oa55XzqKlztiArJ8uOsAcbcjEMaUvI5SIl9Ahiw8TSaFrcoWDozAcBQAAtOCg
/6WOY0lv6XzeFeIKXHK6jCcjjz3zZMnk0cNr4b1vVlyAcPeJW7QO2MNUVzUridTE
0yiIHWHh0ogHP9U87Q4sMbcxohvbLs4kNoXZnt2hDvvsZv9lMIRyUUzEWHEMEsN7
FyOOgAhsIVRzKNyZypoiK9oqV0VFGGqjBO93eKRSlpT1W7V4oSEJUkFXnw3ErGL6
ot0B4XK2+ebynxuvQeKj4v9h7dpopLEoBMzSjaxNxdmoMJlxXF0yQLVWKWbyqcYU
aBmZOqd/bIteqEXQv6YVuIHulkiLYy0lFHieVSbakzlJTcqHgoF55PrIKiQq+Afu
M6R4c/cgTkcNQRIcol79a/6CHNaq7tnQBbaCoOOpR+t8y3I5v2YjapmkZRWKig0m
t1295MZSJcahRs/ZEY8m7sorOY5RM8LYOWk7yDaHWlolVIsA3/Vpl0cbvA0zVjHR
tk4EX4qUYqN1y83T5FjMu4C/a8itYwHVxZfOyNRfd3e8UJ4vDYE2Q/bDaYsMaMmC
SJ9WJrpNJmhKC8Qdpntr2Z1ugfyP9wWArkK6amt3D1T1/NzJcUaYF5QHFSFRn59i
OagePQdDzaEPO1MuYrbE/jtqUIEUqNgkuwwfbca9qN4BZsc/KLKL2Jc0tGoK2jlD
vrTPM8HRksoCkDqIhBkSGXQ0dv0JcMyy1Blkvfq/DsDbVjMKXAdFpWQO7boUxKjQ
LxosXUELkA2rmWDGILkaeWifAnCrsAuTCMHNFuhzCfPwGzP187FVi2xYZh57aOly
Z2vIfw6KHZCa5MmO5ur+JJnAFe+h24mt2Y84pHFGDuavOGAYolhghkXxo1ZbXMyG
5UJGLf1tNyW87cW3JhhLTiJbl1Cd91x93qs6aUbdRybUxDmjDlDvj3LzqnPRKqLy
1e3ahueaoNhZ5ivGalynrSsoCuzfMpl9Vy4pA/51SGXIfMg046uULRxBzKP+2mIY
vUE7fr1nxcv1n9l/pOIMMs6vIXHCm4UhqULZJ6zUj+pj02OCgkVuQ6UvIa3dnd+z
AKtYlvz++Zr7g0TseFpkVb3Ufkzy2b0FPl+KIwqB2jJtR2T3dI6EbUMSsESwWWCc
fNyXwZMvVUGdODoRZmR12oWJhc3xfypy3esqJ1avUOgyfxpacr306hkOMA6bcTWc
X02lI6aRSdldHM4n1JZclFQeyL+SrP+ncCzC7rqMoIzOPAOxg3MLWq8xf14xCSI+
/zhhBgDCf6EwGYm3huc261G0W95kfp4FTvgn86X0cWySQ6rj1Gx+e+s2NP+YGHx6
R2aYatYBlznv2tHxTKXPWDzt1hema4+KlLaB1hKpbDb8k8p+9XPcEREdCO/f9tyo
0/9AJikccVsC0TtgkCIwR9UeTTX5xsU9cyNR/8sV1KBBM7jIWbq9qcprgD5BReX6
KmmFTHI9l2arS4V8z0bvcANIOhzQYTDSpDM5gk2L3Q0Ox8BK9kE4GZFElhQH4M6i
q1aRct/w5kR+H2wvX5xx8beiAQ+h7vqOXgT7L4/AYO1DGv7u5n1KEnKm3gcZlk+h
GwbdXy87D/Xf+VU5BA68nTQ7+LHCn2Xm+o+Inu6hl/SWVuNDOsH1+JJrGNdZCpLr
MbfE++aGgQMCY82KxyU6r3EAjiTJnkbbQuczoCE1gWkoT/9hligZaiFne+1qC3hp
TK16hammRBiA0YM4zKly2Zo5BuwHDf3Mt3eZKl6cJ0XkNVNgUwzIUW6XxScM2oNr
nwe6U1HfsXsTd25/jqMU3BXs3TriPof713AOoiqJftD36eX91MMfqRAOoyslrfxt
dklW3K4kOYlqNP2FGWPN2MuSJD5Dzfqe94sENy+BW1b1RKotzcgMIsXCozEP73cT
77YSEul7ZKxGz9DT7B+FL92kNMe5ykMw1WIZcS8lzl5RsG+qNg2L176XAiJhzYaN
O3FdTrUd6eJIG1zaB7bubl1srHwC/SrE3k7eKFRy/tOXRs+5+1s/yNzz6iQu6NFt
NwWIdIhIWoYZHfU+tIgZ2F089CZcwbDd3da4UI6NdY5fVmdMg64cCNXVZ+ce26sU
F+ChMADzI8lYvlREbcMyFqVDaSANqDgsZph16zePP8B7oqIQSDD58DSAXtUcoY9h
vVva3fhwEK148+h+SEh8vnTrETEqerqeTKB0Lo7KJ5iHfeYBH+EWfRMnZA5taHR6
a4nZ+cVGzum0bGKoMeQGFEYjq1vJhkLrDuVSfjTM0/KuQ7EuTwqdDwN8fRPnR0Ft
aR8B7LNBI8kh+C4Mc9o4hpEzDk0SKNFk+ucDU2qgrF/wnoYfzRJQll5+Aq1/T6Ev
eLxWy2vbFX2j2XtUydLwcxlxYG/+02jqesovP08dXavGZQ95MNyIf4wSvrUMKqiN
UvUJzGRSym2rLLtdLWWQs7dEJ7ZGEt3L7BMiULQokmNH6g9RM3eJZqfZfPhbdidH
uUiClvtmSN4H/MVs/vSVUCCF7SHEw+MK8Uvt+kRacWqBhWh03RNhadBd4hIyONsx
9M1/xEHlE3zfEVJYX0RSiaDvSgBmarMz4wHn9pAHuq7zLy3KTvnOiQxfT2iu4ZCX
bW4wTn5+Y7lNTfXpLB65s6JMNohv22cozmuA9T4GYOLZ1TmCGyASuh6p7/VyLf83
f5DSwBjQnztRXRdKayCXm1rZTfGSXQl6SK+UMQpic2RIMhCyTcPx/GUEeo0SqBua
cgLU7E+YcECKcEIc7xJjcIFmlLIWQroRZMpBGMfm/JE6doJbYwuJunHlTEDt2eNi
2Qz5btaan6PmYvmMApF0Sc/LXOsBWO+AAJUSGoX62DPjjbaQ0RC2H+ojMX+Eywi0
KsBHL9+UgWGdwRcQCgMVOMM5CF3E7V9CfYqYrQgKVSGB1TnIvmk4PMdWMESw6xB8
HlCGNaOV6rliNz/hQ24E6d/UBHuCgusz8MAotaWndEiY5+5iZHannXoaD4Z9HUZj
QeGE2ZeLRtZcXlXzCzHn09OhKkXdmBphxlHFF1slU3QK9L17SZluTpuBRluLXd+6
IBO1kgvQu9SMsu8Fu6bEN0IA1SIiBUMQyzXbzQ8HB6RMbbNVCCezPbpsKKVcKPGB
h6G4c+EggxbCVscsHf+u7HYHWVttHQtWk9FtSAcXdiPvUK+rCi8ZkX7cZa3zec5e
1FSWLDe1w1VcWN1GWKkXlk5IBQ3PAG47iE9JkRQQx0w51bZKiuLbBLkqthdIlNBO
oKEeaRfKCHA9fbCPN2Yeb8SSfagEVKWvyRaibJ1MB+PD+LljWACxDPki9gzCeu76
s96ZqgRO8dQ8rQn2Ko9baGKGUF4k9ld5aXKSN6YJeWZLn4Bj6D1oc02GHSOSluWk
grUZYogaZydMbBd28GhzA4oIWLgKHRb4IPl0KIQ33KwM1RimJ1rraOKPaSwvuXZY
9Ph4UOIgsSTzTaPU3QdlFP1X4PRCdcpKIIYtZmWKq5ZIB47b+DTYyfCnrb/V5+c7
A1tAl2yO+haGp58Tek9F4tbwWyLSZrf+mOXFM65J2kwe4djMESDoYHlCZ0en16t7
12F6dvasjPdCAqvjOjKK4Jgha2Hy5DoACPSlwW3Xlku63ipbl5SFoqdJQRKbWn4w
9XS9p39PONFjQH9bfr7brB1m4AeXh7i6l3VZod8RGu9dqJzI7nIkAZHjPjfedXyZ
HOCq2PQVwzMEwwGpwtTAC6KSr2cFRMj0AWfY94ODm/gwFKrM1w2p9vAxA1VBGu6B
nDqLADoWRMMl+7zUyhs3Zgwrd8Hb0MNk5zMkYHm5g5o5mqkBADwleXv94sm0L6zv
xMux+qW3PJwHNKT0Jn7ea7NSiXM+bKQa0RbWgUu2i1wBLKOxY5+r1yhFtlbiL11C
SL6gNmHvyWHbr5Myjz35MGAwL440wjeBam20aQ4QfdlcI6ffuE5dIjxLlFnAn/82
lWhtmmtV7LX3ilxTgRjD43S/HfJYbu4AwP0JU3PdKXTrMNafQ/zslgFQZBDjvMtm
wor0OG6taNi6gkLAkokFwus3Z8kjNScpOXwGtAE7ujBTcySfZeDcizkIL7VpWF8/
8ncczVwtQfKNmxTECcWkFahuXuK6M5WYsXgzAtx7kWL1dj8ZxsLIA5yC3kZjn9sI
23BR/hEv0tADk4bqLKSivzkzreep0+Y9pshy27SKrXFNx25ZbhjkHbFR9Effyqmb
f28uulVfoqOmuGBQ8wkXoxfkC1qY4smPOVEHguXR4aNczumIhRiFwHI4hmIdQfSF
TdSLyLPqh2hCGeEJOtIXAp4I84OCohTS6LA4tEky+ifMf9A7H5SUERzPmuo++tM6
Y3lp2TeDf+PexVKd0fnLQjXnpm1y1dtzSERygacmUHADFv/3oYpQUeFBOlUeDSmI
hVJ4DATMAMhcASAdQv86jqciaUJzd/xscUgbSFKIJ0G5DNYIx99v+EFHIr3ReAtk
oiRv3jK3tdJiDORGjf36vNH7zqOp6Os3s8LuA6vOla2JfQNEaESVa5Tcy8D6UJ38
A3D6jUckf0n7HZ1m/CuXFTT8qcghRCIEV7DDYWEwXPI6aBnW2SPPoYgXqgQJEdEq
I/9OG5vQrOd5aOyVRayLisXzqC9/wvJX05MwSkApyap9qn814d660UzpBZVDYXL7
qqlN0TdTp22A33VeGeX3JhCo0Sb21GfQ6l6ZCh1dLVEq62o4rXbfrCKL7wRvD8Wd
hbALMlEd/coIPdbl5HXcBSmMXzjoLkoZAEDod83PeCazeogVVcp2d4uuHwraNrFG
aMxMqdpk6G+nF6m5CyXA+y0kCPJAK7kgxObzXy8N1e6WI0dfk4AjoMyzoKjiJrTW
x6RJy9ZHhctvCbM96eO2OrjJCIpJsnaz+dEPnuXWvzf9bKNyLsmRWfWK+z07W8Rd
JcDBXtALdVDbYExXxdu4Rjvz2Jh/w6HcJZHSxwj+6DdJw7L5Dao70HCcupse3WBo
wksvOohwrkk/Eiouxt+W24RC2KMH5+3J2LiibqnLR57KzemmJ96RRy8ngSEINkva
CSQdn6lNQ3qJ1HrTop6W9+NGqWEJwAlFUxGx2kUp8g5tj/e/sp38fOnO80uQn5HI
PF0GYYlD39tiyDnuSymOvH8g03I7BDU1B1AryTno9Z3W+IjCaGpsbF1vKU+pYQj+
Ja8xpifp9feUboRtfrJh+9yX5RvOA2eFZBot0A/wK7f3F/4/TMpjpR8kGFMMeZ13
p8lBlaXbupAuDxYvNcG4/AyxUnsEWG1nS4z/Opf5WiDdsqIxI8xXStIi2qAUMLxl
nSOAEWlioPDvRuKFbAk10QnjwIjEKgdn+Ui6fl1hLGaynNneSJvdVFfHU+lZQpGp
5AnhkP/BfSyf6+vuGKw/VFJKnhXKo4BnLNasmJ7MF9XJESZOwlaPQ8wjagitY2pO
nAuZe27k7GzuBbP8m4Rf1lp8QegEtWwGk5l+lh+nExiQ/Kouegk5aiLZbpR9AOPp
ENqYyV+KYw6q2nYDV8MPnvA5BVnTXm9k7BaI+sisNqahzVAnkd96SIUUEFYUGYG1
QqIMmd+gX3xv3l4rJC5HjLiwYghuOlnAA+4HsQQNe4DcUbvwlk641T4lrLSHxE+7
p5pAMoVujyap8FSXmQOge9/hJqNA81zkdqo66jUE5Hryp4I1H5uBfN+YHt386euq
dSkrB3rNSmmG9JTmuQs+I5IhTIbQi/4s0PKlAH/FKzQ6qAno0Ds1xqLaHXNeHaPg
J5OSzVASk1d6EMnBsq6uAodARSUdezOHYoS6XMbMYMmqkKF6cE3qQnECmi/42CVd
sjkvoz3h5DKinDDVsy+DI4x+Fevr/Anxw/8xxF0TAMYOnUGDZJL94S4SKFN1YcHz
3iiwS9V6WWga9lSx95yrW76UQrtYfGALjFZNYWz/y6bKe0rhpEY7v7LYmkyKH9pH
yx8WPYgBbikZdMoqxBvMzxtgy0TK5Vdsh2QGTLojLSeK6Ua+vBwxND/AuuKbWAFJ
GUbR2Psb8/xIWR88tZLR3jGwp8PRcVePzjbK4xtyzRUrToer7ZV/1vcJjf1DAfKc
lssuA7ZcDoN11BlEgV6iCLPfKwRDSq0tKOSWgPnTbjGOmFbvE3wDQPFdDSh/1wv3
HU1pQkEyaULorzZemWGTeY/uloKcImcQOGQPs98qlKDz21kh/NSFqSACJKHfcYTv
ZNsmofOlIlxkUGC3TL7kwgGyDgU4oYEq1hT+iFJyZvlPmfbw8V2zb28KKAR2Jqin
bgGiPxAkrFw2UqjqZnzFx9E14N7NYrQArHg95i7TB9RtK87Ip0KSRSoN2YA616nV
mNRYDgz7j8sNQexdu+9ZUwOdJdQKPbqpvP1zcQEmCBbgjUS2gr1UWmwxuDCisprm
zRQ34M4mqFggEfpHMV5GHFKxEL+hVM9VhcOYq906QD7gerCFML5JH+vEm8mVp70Q
ZPIYtJORNOFuKIOalN5X7FXDoYZPAgnp7Dy5Eu5C6eO2Sed1DiWd9KgRSSuVI2Dc
RP8gkBln4ce9mc/d0UlKHxy0awkyL/E4uyOGMczQCKuohVrp/SXdCJ8q/ZeRg7wx
M+L7/+CdWMJECKX+WRKizw8YnAN0vTXKIZLFTbzYY5///NfqJlvkacwzCEEYeOG5
H2lUzic7/bzFaBQOHA2INHRntsjvpSQK3ZCK/Vy71c6a2x9fs4Be+gyo3v133pBH
UdGAeH/m48tYzAm1uHk4V+YRQ/FQ1paiGuRzTSHcwGdr+VCN/XhCihRHSIkCiUxr
BtwOUyjgLK4ZLlgONBWzaR48AFVv73KwmkLRnClPbAryGmjeENFJ9coiobJd34Wa
F3hw3KFEnZthX/vOsxoPidy6+TwdSqW+pqB+SZIk1RRyiaa2TE3lTeTZUki+r2Bl
6AQKP4k0XggQe0cIFKnmVQniONq+FpGBjyjDa7q06gL5UfUwZDWCy0DHzP+cAehc
jVlFHZqPIeNDOLOQp5eR7W6zJPNn7zmfUp2UNYEfDLplnL3LcpvQXtYn4TzulmTt
HBUgdI5kRBlo8InHIxtjTp7fyhv33YZ8CoRaKubErm3qr+a1Dm8rVTJljmnBlSmn
jjhjdk5d1TAez1I8n2NE8a2/qjGHyfUtlC1SFeiCqqHR5ptqb7qeAfdMQ7jQe5u/
whqp+ZOLkaAd9ZzaOclsSq/xCIAXIQSO++Sf39YyzcqyMGtsqFnIGNXYDsgAroTT
nRo7JNZpnzCagPQm3wK3WUBnZCd0Y2l3Ciht0tH9up7mRSQL71cmz0v5Rdp6FwKn
JynEq+8BJH/o4J5cgm4Z0mNoFHmZb2apKhu5lF+2iJBUvmlaJH3MYHHa8Jbw8PZN
7eDK+tmljErtnjbXgdpCBHqKH4HLx9r0a3XMF0LFy/hoDHleMZ7/7fyAVuNq07jQ
zf3l2ieaaIqvXAxgrsQ80+O0JpuoKQwwltD63NjI4Tb8hWZZXEeEFMgSetfDT/vs
g8YsR/yx6hHwSiX+FFzRMdS8thyhp/pC/AfVxBeODEdqHZibHCWlRQzJMXok2koz
1/i+ZK0yssDp+kCETq16aAWVjLNTBNphJey4ePqAzZ6xrYeglN5YQVPkUi3mEFg1
YE/15yg7v0O+jl0m2idX2mntdLVZGTT5bWdi0h7UKuWMEgBhjMVzEU/s23TCDni7
G1g7vEaQjAqV4C3LKswShfDRmy0xiwGjzqHM3Ve+QpWg6a9UZb3Ohj8PxdiTAJTe
eI8Mm+rLvx8zUkrO7dNB24Vg66aDozG1Mf0hYjDHELJSskjPPPCYhcIwLchU3+JA
o/zOBWYCXFtP3m/a9uVJBgwY2oXt4IYWkZbbbWQMhAWvND+paPSorairfgfUjuJo
fgr+JF61uHot5TepQV/uKU/0nHZmqqw3mQ77Uuq5QTOb4tGz13oJbNAQY7pbZpuC
yxTXcICXlSzxbagJL5EPcpLJVtg8MXBt2nOhiyTOxWlTIS/+r+PB4AJIBLGsHOH9
Bo2gHJ930IGh7EFIyBIghOuHhSo/UsrhdM2K1hVQ5vd65Z4vEgDQJz+ZF8ac81il
oRsqNjQ8ic6Wl2C0MYp9yjtVY/mEjNmdaHzd1TMDBgLHJiAPVpDDEU95fBRE3x/w
WO08y/Xt/r0KH4IXaiXmfkPFAgkokL6kvPOU1sXqA7svsF243aUosnvhmButTxUH
/sgybwUfNBowseicxkAexo54xvhepSnN1IzZREBjHpG6Z1yZ8zkAkgatkc75jKFJ
yZ/KRvT0ZdkgRgk/qxd8Jx1QGk6qZ2q/0MYhQEZvC3gnj6elFzxIRF8X1asSr876
8PVYCZCR1+UKwRjSjKu6vC80cfoTVmOt5kVWwFOWpaZmqiQE5pXmGHTDMAQnLDjj
VDYcbkEcHr9Yh1+4JJxFXeheO+Cn0m+cyBl8E4syxqMMyH2OkKXHGHdIpdzy5kTf
yk9P5O2TKiGrjxzCL/fo94yKTIeFSIiVQM7e4Y7hbrKyKjO2z177Ahjsj9eZS5Wq
q+wWmjTiVvFlmDKTf9qKMCgZYiNNn2/dvgSNfHoLNjrWs9ZkTLRW/YSWYEd6IOOx
SLI092t7mvSY6kkDTXfbWe0csDn4cEKJp8MhX/xaj4Wm5Yilq0LeGqPSu6tdQ4C9
KuWZSOqsRlNC1F7stBwLq9PInKibLIZXiZpANHoMFXC49GJrvrC6S5sGUKjngLGp
0QZxv4l3wOGevEFMhMhZKXAg6RGhpa04MlPze8ltvmsCYSS8Ty9HP6qLYjOlLSoH
if4VDVoFAWn5uvMqHHet7dHLU2ZPVIU1Y8MqAl5No4EzP9Qpai2aBnsVKD711a3Y
n1D4fgA4NhU+rZpXW+kryeFle27m6ZuFPdRU4sS0dGRxgiBRiAYTbV6gqnpaQg7u
ySXGs7IXIsqR5dQ9bb2XHn2UfbXqtMLTO8I/HXKnVTCB2iTUfrdXZhFcdFRDkSQ+
zJpqpi3+gNZJQMQ7pt9JO1VDEvan9asZqarX9OcEin8uc3DeO8x3BCb2anCjCZMX
1pma3WAymEiaX4Ila34OsLZebXOw3S9sskQ7zcEBwF5qq4r18UiZ77fscBFDDnKD
3BPtfxLE8x3p2Lxt9PGIz7Ak6+6lo1h+/pycGftUljLlA2GaMLbAvCX3TMiWGgxh
TWFgrjBjUcSWhIJKGhwlchp8k7gVURMCe8PwBTMTHrADqfkvMGtfSKotmfWRRJ6O
43RL3fUqzYyF+rYpRX+ULNafZRRMVV5FIKZaKdMCj0unSZuJiTJOW4DRKx+mTEh5
tg6kowC2jZb4fGfciTkACR3/L9CVJP/CsD6tTMXOoBnTmVe0TQ0D28MLdXOfcGef
xR87QN0KgWJDFSJqayog3RnlTUFqMSE75OEdhGeiJOKzN1h9SvMe8L4RarFHehSo
wNO8pT+HACgaP8zFD9d0rF2xmrcDT69dcQ4Z7P/IY6DmjzSJzQd21RCkxPSnv65u
+rF0JRMXM1vA8K+nl6e9bP0ZgWvZb7k+ncHskm+qUShWGxhMjEfPBXBoF0n3dRtJ
LNzdsM5zFmZFEvTYEzmRe3ssKYqvOQs/Ku6NR8/DGnTGvT3J96l7FOU0AzH2yh0K
y2fRmtU6jqFOTFTlSHi7g6tNDk6cEoxOqnOcWbKPalM9pLVv4xkDpz5stLew23LY
+WhgU9YGjuhNja3qsTUGo5JU2qppE+aU0kGv4CbM4O/qTwUAaJIfsr1oqyo34LuZ
wc4cNlIA5dHvuDa8CEzAbzEj6mfo6vl25fqpmgf54xpOu1CAEf3vpL04dt9fWi9P
8zI9sOkTQCn/qL+19/O92FJ/FcQX6PbBEiekiEZKe2bSk3cP4qeWXeEjIV9Y3vfr
1djB2VJkGVlFhRgjABjKR8LyD+As8IT9KXC55wbkYhsQzG2KxAVBxLdi3PKk70Gr
fNPKlOyK48v0U5Lj6KgtxYDDsQBCcwsTAG/oQWe0y894zi43yDzhpGoL6qNvCZmk
fuxPmxCTEmcO3ZpAIBxxYl+4olOcLTFgwKpmH96Ol1qKmZplve55y85ezrloHAed
yw5ffO83/skyPM6CV3u7j3BP1u7mLnPhGl6K6b4OnaueT2qvuhFkZ2nyBn7L72Wb
umlHq+OJMuTAHcGweLhC7vbdvyUmRBB/+7QmyO1to5vFbj3ccs3Xn8blL66KRNl7
yaw+rL9/KHDvbmkjGD9hMbnAB5iZMaK/RgbG0pg1hK/vLFrsfH2MOHriWodId4xT
4qhnrTdSEIAh/EDY0pA2sPIKdmnI/3JFP2iGvCfHFJGPC1SSYm0wjV77yRR6v1C7
xf08dQnaYS4Pb6zDRrE3mt87SvGxTr2BS7ZXUFiWbQA+89mR5UiBrhknDEpnR93Q
mvwfeaJUE0EksF8nJEkd/Th1kK3GEj4pYyFmG1J36N1TKWaVWGPRgPGU4OyjJvLW
raJZvPQnjzKzHFYQKmHqUygGkUjWS1UKJbt58Dn4MUMO8pFxbY0n31EStY5rZQM6
7DSEnc7Jt3sMf8UDdqDBcwz2KdHs34nwnO0lrLRBg4Nd7go1SH4Gq2qVaII4VK4m
rqMu0UEJ9xrgxszd2rDUg10EQm7W2ySmW/oJk9XoeOLlK635hzdzuCPGkBzTMPsa
d8TJNyglOZy3BqWjt46V1rc3Fiac0Gvldx9YBNQakBPWZ6iibCDrtaXc970ETq+7
IsvSCzO5OoXSSo7+MHtuefAfwmyDTr8CLiT3Zcf4X0C/SkXhR+fKUAClQwhz682K
Y4YGoKm4iyhq7GbTeZxWwgbk7XDd5Se4bFetjVreLnM1aBVO9Jl8PARxecV19xx+
/brv6jkAsyn5Pxf0klr1BQY9Jz4nVNYfRatxRUxg25OJA0ebHkNtH4QGSk+IskS4
C6vvWzM3VQeEzHWY02DjknsZ7TdfsM5jU0obIsXPrbKCvibUn9aI76dA0V7sDMAI
BoQvkypEb7KP4w+VFwdrigQg8aqmiJrYVXb9B64Ra0+fxggOnmKH8OlBtYjtXBxm
nBxEcpmOAdIPFfUH84LddgCqoT3yhiBbSYtDS4McyJZUeP2AzYLeXCVgEPoUPkq6
8rOv+d3L4T65IGvy4VRhkva+LnROVvE6ZBKLqB3XFMwHWw5qwKb4ZRx/SlFIi/W7
yz+WPCQq6WynreJ5N++V2Bo+c2SbktZfn0LH64ZNjHMvI5WYhHIEpKDeq71W4t4V
C24U0pZiPICPbbUG+pYyOshpn2usS1m5UE1FoXOV4Uu8Mkg9g/IHlbkSKrTMa/PM
K3TvUxC1aQAbX1r4skpGKYxpv2DfihVfYC4uKiCvVgNzFwg7P+EN0wcvD7C3H3jS
zz7DBvuXF/0CxEKlnfoDjhxltrFpjPvKJ9Uv+6SXuZ4KiDuMdR8gnQDsP1xSfMV9
hc41jU1hDUKH1/ueVwQmWLgIUQzv/dmGxWbxiuMTMhmLqAUNP2VqWe+wsoTtxMOt
AniFsOP4TXuOdC3NZZnt/oZHZrlNSq9NVFRROiySiV33hgD1ZED+sPsfmvxWj+h2
yXqOSEIHnSoR33ZOZ7J4idLn5VUAshI3sqLN9Bg3ZfvzTCDpqT9qCBmoTxnJZZG2
mWtSLhf2kvfLt4n9EF5ZEDpcM4dwMIDMtiFNh/+k158/sAGKGv/Qc54qyzKg4ljY
qMzuq6lux9cWeFxFcz8GGvNjeP3WZLRuXfz/vECQ00b55kwCXH3J0ADK30vPPUx0
qumjH3jcxyXQhwdHUaGMK3dA9AkND93tHsC4/3a83jGO0y3wkuYSgNodXsp0U6GS
Cl9IpKzFR2ytMedjh3RdlrO/IYb5qvKUIjtWOy6E7Wvefu07va24GjD/JhqYfXdt
3+Uuk/KbiXm2ADWaNjruoXbwbSuPDiA9ZUM4hv9nv3csvqvdfWdN2q0V3Ws5RBZA
fIf/gxh+kOuWRymGMhZPW6U5WsV7F+7orrUUw8MyHpKLLT/B8cwZSsPh+cIxvzh+
FGmtCkO078/uANJ+O4WTDejofj2aPgv0irs9pPjUFKgLXWzsJC/Hz4KehKWtxDJN
BNxicLUl6TI14B9iZufhgmTSFjfD0M7YHFARXneNdMbT9WpWMXbIPGgiiF6XmfwE
uyU5u5CLJdEi4gtsKMi0PS//98m1glC8ZYzg3gQxCAuoVr0G7MOmh28lQOPTutIY
OyEheva/2Rp4lYUpjy6kr66cLVCg/m/iCDq7ni13O043KI4i0AkcPZQO//acOD1E
NNJtfhq1XvuW8+P/M46QQUI8kjRvTspBaOskiF8q/MYLYmfz+6rsQkU4hjjvwckG
1oAPofSoDFpZc4wvB2Rf+zfaYLsq5ElryXqEHOZIHRMxD/81DX/YdxiaRsNyJd1p
t1H+uCx8h4Sc2m3qzswUD1p88Q+YU9SY35fa9iv0eL9TbfDT8oP7mGbZYFaRJpWD
UivcnfcsiyHYEmJOsrkhYYyZFwpQ7nkdwkAFgDnJroA5MuvXq/SQEGZgD07/4EI7
+GITyT8OtIjWOjLPTyLjn25EcLSbhUKhtD682U7DA2bkGjcmww2kOsos+049yLpA
YRUwsiitwp0ey0dYdDXCU02VeQ1ReSkcA3u64b7WWVt2/3wJuTKtkO7aDDM3baB/
gYM1COpX7MFgRpaoa9hRfPW2uy8t+zL6t3r8YFR3OZ8vbe0tyMTzU9otbDJYrv46
wYyUrXqlvr0Q6qXiIt23eB9dKO7CMJqSFuW4OM8QcQRZfC0sZ1aVXiRppxbiA84r
ClEeUBbvO4+/QszdTvfRmWNsKstEXsWRIXEK2vam8UXX8iHhT7ecKXd1gDBaLz5Q
hmyMrpBWPs+1el65bC68rX1z7Z0PEJFKGqKs6tuHQJiHtkzq5bMdLE9yy7Bo6PFs
q2M4NEvG51UfgyZ5fq3aafLRAGrf0Moqvyqo2Ocn+VQi8QBmSzRkXcRADH8hKTVm
p17DhD1a+yX/kMh0KnvVbHmYyVixXaBqMjDkuCqt9bY8uWeMU8urPT6NNh2S/uag
YomkKNBxVg/9M9U33RXjp4uQX0ra43g7zXBt8ukuN84Lb7SB/6KfyLC5ZLuQyDkI
pz2ccqJGepyHDOjfmYzD6+090Wqv0iHuqvQln0McsjVtBpDgGapC8Ol8ZP5gsNAa
2PZxsUky6eW5mqYcMPcRsuXi/IVTG0/tt5raD5KgppJDkTnT+CuJUwx9Z8Rkm5On
PwYyj7BJtEm3KlaGxx+HJxTk56wI2t9UPQbPUk8QklkfLWfC98+PqxAUASllbPO5
gmuESIVPWQUPt0fMfGuDJE+7i0FoNV2BPZu+H8YkDJDzbzh1ce0piqkEBvwEyDNV
XQyuvWl0kLp2widOOkAafTFCxPj+pj0ZSWbiXfFxs9KaXvZ7gHUyHsrZ+Qv/jrBj
5ZFoBmbylTpbHWjMRqg3g5bp8M+qbpwCXRKTWvPh2MH0FTcQi0XEimz7vEDfoTNw
fKqIkxwe7wLEkmn14Ym4qFrZKcW+volXGZo11cwyXSRgAqVGH9eaWwzZulAz3BT/
vMtwTaPsDYfjg5P2t9imw7qcwOwe4OEyw81blJVTOqU9221CZT3OoJ/QO5Rp7pgT
PRHA/WYgHSGIi9KB7YyYWZatIyPAvdpgAY0yTlk6Rtcn9Y5w4yZlHy2k7jzLUibg
8jVv6Qk3Y4YsNN5G4t8KeobvSjyIljxBYkPdQEz1ICi0EXLIBK4OlJM+1EMMBE4X
SNU3bk94q/AfOgvgRgnNVOVYFkCXgkVjZXXK6nkXEZuonntx48U/us+6XCpwIqK5
nRHHLjBjUT87y6VIsTN6ON1VdKf2KaLaTTN54enNiTT/yzERrVO2f89HtZ5y/Kah
4UgGHuJzyT6aiZvkRwwz9FrSHAjKecasY+ZftWGsG0oxWkE2TAwZLeTH9eITvvox
a+cI7MFc87XQyyLqeiUbyToi4bzccQBbW/o1DVMf/G+8Kmz0FdO/PzjypElx5Tgb
htbj7xk4sUACmzuHhPoU7gL+5HTfFGt6xHl0zhw6j7m2xgtAgNgsnxWFp2JBwr6O
OCuAetzSObnlrD6lidGn3jTHGdlXq84nM2fx6KESvtE2Be7HSxIKTFbfVusiaY47
t+lv0PMeVEFj9Dinfgn8ZskKmJhx3Ln6y4RR+fdj3abvDsyk5ZlmCzcZJQ59zL3I
SY9FR2UvZ4v9Pl21iUdy2Sv14rk9GpJy/tyx0oW4EBb0sNSYC0k7HOx8KA+rIWQh
LwK1a9qyiuzNJjGOpxjoOLT5785KOlJdbxGfKDEY/X3I5eeFySgBHAmjTEC9vTtQ
v1LvSqHldaSkZLmuepjiO+c8WTm051tsc1yvBevC6a+ECVOkrtMrD0N8NRMsnUvM
VCEzVwGCjXYYvlHd3Xaiz5WRjMaOiTsgHr65m/8g9wRKt1I4tB9Jrt6vK3IzpAOv
IplPm0QnlINffsvOFK49kUDsrPMh/IeeKTV0LbozhWwou4v5Dl8ln9mLwcxlv8yr
BbkLXmh6pUqc9mtBxjSD/sAGiN53HOfwfr2QeZksIj9KAZc9ZFEE+ohaLEKwr9o4
epWx6WAZ+JwEkdezJ9l/fJ8Q9YH4Vc5SzUucfr9SQtiow9sDSH7m3Qs/oQapWgnf
t2y7n1mPgpDwLf4tBZMpYGt+Dk7XxlgOu8jM3pqFSqK7aNXXgJ9ZtqqsgJgC1z6f
nqKjAWRQr83Yv4JI5bvND41HKetgFt4slTw6w7UqZkQqcLdxEeBLqRG+40Pnbhai
C1/+BRMXixbxvPo+tmmQFRe+m7u8Rvt53IosXsF5wB2LstPFMtH6aGNe+EifrU6Z
c0HLoefxDLX3ASsuI2OgSvAl+Dmbp7/qPY1giy/Y3iz9xdDF7Ox35V3LJ5bFGDgX
4lDK+Sf9piKAt10LOXD8ARPa7FVnT3HE0m6BRft+g637kzm1XsrxX5FWOhguTfB4
gW7kC5ik+Uw8U/UzpUxDEjNFc06ovzdHQ/Oc7U+sDBc3tYaxRrC5pdugpQBN4YCI
bkZB8kD3kzZtOUJyVvkHoPVWYZENmafl0iNAc7fnf+VtwOEYiKprsp6I2+UkTYAd
5bNE52aFH9SgEmjLe/8DgkXrGAjALzEIxqcgJl3RHtWC1Nzq+Jw8ihmac+NhjXTR
5xfinFmxrO+PPc1g/Vv6pM+1rh2SCF84qT4SSsp+Zax75XEAV5xofPqgb0KnHNA/
s+cGltuTc75dUS1f6T6d8KUYJTdhw82tfi9QRlxauyEEKanCwLaVad0gyKIrl83+
kiiHTKrNSV1OaTGTT+cvJ+UqrUEY2qWP0i06iA3OxDNAXkdWzXjgSB/4WPamEScK
yEOunBg5kynohISce5HPDSeQNQQhQaY7WoQZ7OP67wrIL6ZP8Re1zT7wQuqDfP32
RuI4yaAbfeoriq4eoqsaTgeHYpQZAYTA3066o7tZEqluCDvy34b34B3AmbaPpEoR
dLUJ6/nCgsh+pi8NRA5+rYk4xe0oUfM+XNZ4kS5oQVETfSIrmNSDmdNIYAzdrFsB
9wr4pWY7H1A/UHGpCLllweQ5LZJ3eHnxKQT8VSYQQOL2hnKxgfxeHM1Sk0lDmHF+
ASDw55CUhKQs7yw2geTHQIHwtYa6MUk8zoKw3UB6wR+ju9z/fyLa6W4GODrjUEPR
iwemxsFjvh60STWBVJXZPBo5+QnllR+MrsrAfIO+O9ZCnTgSV83cmybKGOcB5RR5
gm9z+1WDSc5I8qWpqQvONPLXpRJhRPkNpIB0T3xuTFGSet/HKbUony8Zal6gKKHO
JI3CRpnIk7U3EjBY9+xw/zBMJ/ol4Cb5NEt+EKV6JoklTR6/fBCXcDVGsikwV5sj
hbOJlPFpFW2Ewobsh6goWuLkYFw8ACyImxo9rCJDTCsXyXbNgyY4T0P/2LfvRgyJ
kPOZ9HK2bmRSCs02wR9dEe/EYvz8qJ8d3sz/szyYmaQTUarjzz39Aq2IZn+TBry+
AhQwUEMMOqucLOl8wjS2I/EgZGE4UdT3OnGtxTQeDkeiDH+xjdKzix5saaG8fVDQ
9CHoRNYIi3wOXfq1KYJUXcPFwLInAEjFxPEKOuPooRcNIiOdkr3m1qFP8LpzcB55
GbOPSMQv+4n4PBiPMvrihvwkkRXouAzdHBXUo/kv3vjkVt4Irod3EAW8AAle5qNV
BGSD09n1rzWVdmqRdV4JgHolTtfgdvRcQV5QWjwT+t1tfBhrKnnZxepCb8ZNryGL
pnjtFt+a8SLUZ/UqRWMqrZbt0ZzqbX8vSGKI7bJ+8Iah7UTCTIK/YH6eX07MJJ/y
+M6Ta3QF3PCPWPRJriY382yB3v1a2r4QYRhxe5MfSQceXiqTuwLFS8D3JbZ3hJJA
2IGPEr5tXRDOE81r8tM6Zr1YNXadhZ2kXHe9Kv3c7yYqxikPni6dmgDAjKDJyBo/
SNFf68XPKJ3NmEby1YtLM9Tw1hK40oLd434Dwpe3YJsv6BmPFl0R44vxBdpAJToK
6xzOk6+Y2xgxNgTzL1oCwwWAbNtnGmPMTFubBnHkUg7sNcIYkOpjh+enlVL/E7ZQ
hB+3hm7T/n2v1pDUX3UUBv2VnINv4gtpOsjh1Gne6os+uPxYVvaGVScm+Gh9NsbJ
FZ1GlOCgl/0FghFvlX47TQlzAhjP2M6E0rHRlDVRfjeWxv5lcQgkfrhl62E251wR
8waraqRsDO5ElLjfggom9GgqJo9zENm/l1jm2yDvcIs1I54XXCoaEBV9ulIfBsYm
Tzw6pGZhV5LlA5UeM99FE0zTDLPqvurGlePBYNMxiTbpaNDWrrC6kak67T+G5NNu
h/1JgwOw0CqvP0x7RJptUTbJX40ARfHihZsbe8pw4LEF6wXjNdaOOAlHX3OOfNOh
IH4EqYg+d49C5B4eurbgC2tY1brPJwuyMoBRIwdQU1l2tzquF38JG6DjAFHtpUQ/
Z8ivcCxwLrjMSrxTwZeVJHQRUzEaZyFrBzcWUc/dPxeZJuL6TaWIOAu+MREVUUvs
L7tdOi4ahbX9Ow1739meA1A1T94yV3Fw9Nqb3AFWCELc399enuLbR+CYrSG8viMn
9RLqSfP26mfWAdf4W1NVkBq7y9QzekmU03Nwi1fa+OXiiWWlgK4Rmi9iU389WbBX
G14NXPwsMVDatiE+/62UpR1ZWfkSLcwOxQ/uHd9GQL33YANpU2LOJM2de9e5B5Rc
vbim1Hbni9bzqE6+iw0ylEYBG31LBJ/SipLpzSBz8BYZg8i11BK9Y8tM1rowPu1B
wkrsy1y8N2eeRZJ2qUO8E+bOMjMBUtDHuJubO+9oKalJMj2xEcxhd0c+MizWGOtc
WboA/d/PhaK7NR65ZezntdQ7YaI9+290b7q6BNR+PnG8yBmzvpVrY2gkBx59zbqc
R2x8QoO82zUmKc9tZZCegVbcsZ2e8eoiMo8EvLQFTvd73woA6GCUTux8iO17ecD+
hSwndu8EUGkBLa1Bbka76kvPpRiv8WrKnfuJhwH3ZlwLltHkpgkO9NWjsCYBLTdb
Er9rQMuOlJ9bitOo+ptd6yCuOe7G3lm+wwLWbvm+H3inmFa643yP/8KVwz0gzXkp
i6IhaEZaaxQC27F+9/Sd0YqqIM/P2R8794RLK+0ugWpsMVELSYBEb+qDlTH8c3LF
qWBJqc4DH5/XF8gC5TKze1PrG0ttRsvt1nXJci+lCJz+/ToLRezlY8eG4Hj33Kpg
Z3/nFRordOdAhZaZb1aOPBvS6bPeQ43JItWII/kcw3LsTBU+pkKUA2JM50lHUWKd
h12bHT/Ah8F1/x94Rh8KUwgzKkj5FCA3QFZvWV9WDLDl84B61N1Zs9+Rf2OU9AUa
AbhTwyGybLL0N0+Mdj/Gd8OjfluNqh+PCeD5IB9kriMxmFftwvN+mgVXGK3ylqlv
7uPl/9wC8BeZr5LMl0FJpa94+CCfKBIUd3uUYbbU6f8c5b6Kik1FVcWlQ9ZjdiIb
mfIejBHWAZrTQ5CMwDV9L2k/Jzd14OB1MQQr4WPfnbEcfaFJUrI2OFIo7EI4AWaG
lp02UVTWGpS3aqAhk7c+CAyAyrzJ7EqOG1LTCQc1oYQkX31yGrZk9YLQpsCnoQZY
Tb9UeBT0PKNHR8XIuxSmTi5/V5n3Rnasuuq+sv++WihTJgOG36M/3egE9O5KVIEw
czB2zpUzp7as/MySQgjZ5tVuT5nDyT9+W+ZJ3pnteDBaoyLp2SUXu70vTyC3aXUR
J4rBOd8CeN+hW3jLw6m6A4GCCPz3fuYz0NVp4eE7V8G68tCOAH39Qo31lRyTrW47
cTB/4w+Z0uPNgxaOSUApH1+vZWMt7ohWQ2V4KreQ3H3JW0QpJUGCQa0nsjvkxdLT
nO3NEgbqlfis1xjjej8YqXDz9s2TeW6izlnHf3xScD7lgJKsZRIT8j5M+ixNLtSF
Ks0H+WGR26fFKXzsl9/vd1//sGmuT3IEi7SlA4gWDX/wnUH/CYYIvLVxceIDRho+
9Jg95sCAyGttTTJL5v0gfMV1vtodf22BNDJ0su8Mo8cnbl+s4ug7fEP7v43Xr6Tx
Kb37+VYYIMBx+P3mEjgMZ5IA/2BGdMNhTB9+kv2hnJcnYCaDGullcTl30nvNld8T
2JD1VwpzYhTcRvjXfbwVXcFoyTTYjV8R9AfeE92nWxF9ZYhRU1hokEEY/RdsAr4y
gQ+FzijEsHbE7cCvOnF5Mqnlkf4o1A7PqgtItDMTFJpKkH141cn4L8idZ4dhZ3DD
sFNazpwBimQO9o/x7HFv0ll1s/SYqODYcg4+kcShRxymAFgBlwTc8s++rh7DN0tb
RpfegrBqSKbJSTZ5XWwL4cx9d0TRH1DqE8m/77goGLhSwpw/U+Q6W/16+SI1ipOL
kUyIDd/SrJW0c7QjPBrEXKk3tDdMIhs7rCSLV7fPOW1Fzw2SkMAZcP/74F4iSvVG
EzpA4TF5ildADyxg0sNzUL5Qautsu1fhc8VRFu1nTIljyqmvPBFfyH6EKwYpfco1
fwKCbg7x6mY/85+mn/zJxC/1cqG2yBA3ra/NeCTkvmIavfo/Tt7OF1ImRSpeEgqJ
c9BRq568GyBqGrQiFGINatmPr7GEzLSr+NZETWk1xXgM+2c62yJFNM7B9GoLpE0W
YvGe6QK/FpdMuBYgjEJNHO1HpaP3+dSOsaD0ufZwlGt4wKlLjEpLFPJVcUPi0+wZ
RYdDzpnyDxqtT1rnXdtR+19oeEWMg3s6a6uAugjyFpLZQSNBpUm0w7aWW8vrM626
/B8AmrvRc3tB8KDLORV6+dTPFhn4ilCAJDZc4fRB7G1ijM2mIyEpzVDMJKPmG7KA
P1ueriskH35qRDsiIvgZ6yy+izSvLviu5joZiK4o4iK6AlSRwrV5i24LPBKCtTCr
OHw9IldqNuuuSVrev0AjMEq//dJ5gffNCXgj/p2ToQ2STJCP6OCuZ7RRq0nMROAG
WaF1RSvUeNV/dS2hdtein+CLJgaPk9w90uu92AgX1czWJEaLPIR6GBMvjQ+c1hYv
SCTesfEJtvycOhvNLYUug3CnrYNMgXPETXrd85LT+kfCum4mmABrRhhKTUC5TPFv
YIzi4pdcwIC7A9mOqV0rcQow+ljz9NEy3hgaLPbFnMpyvKvZAF+ZglgBnzKgKnng
pFKY9N6ANAu7MX46PPE5QLPV7SPZUbg0uyQWvAAsjmtCC/svadXd/JpRlp3e3Hd/
Kp38j49vu3cfkkT3bMyLWQMHNn5qzmpJIVLE9mz11AwfyhFMW32rM8a/KApVagKz
32GDWx6h6hwsxNjNEfm3Q6QcbtWUThu6Qmyi46n9U4rxNACoflPwWOAkwqONwd2t
6m1ELToPtCh+M9dEw88Vkpyj+d502GGjDy9fqHdsWVT2eiGVWBHzFhPFZQwCINlG
1B9gN+MCbpH3m3TuvWKUF9vp4I8kBas/QMIX55DbhqV3w2U2h1H2DQIAt2NEYrp2
WP8uLzWdXxDCRXmLkFP5d4EUoRiaRhevhNYWvsMBd099nB6Q9dqwlgFPAxe/3igj
1mBFY/IpPAc+dM0IsPLrrhr3bVFjwdVVKJgEAmQEN51lOlXkAOwViSPyU96QEtcL
vqtuvWnNnxhEbnLDdkEICleugcD0f65Ns/ZmsV7lsWkXhce62LIbuPggru53FLgS
pufSl0QnJkl+jl6FhCtH2J4eY72qaJw+9YPK1EhnAVkgmluYLnscaN5nppZnQcKk
qarRX5okewfEOAqiPdT1zBHFpTIiUZq6X4HtV3PP2HSODGWv1K9SERPJRqQ+ShE+
+9KUj19nnNLJEWnCMxfxJS3LDZuz5nMHn01UPZO3Es8DTVLWv0sXxjWDj8c6WtPO
5c+09E/w9d8Qrck9dLFuUxNFcncTGipKPX2x3hizz4JuAN8ZqSu1Ui0USHcbLllz
0FfErYXiV/wuzbEXtM2oxhTEzhhA+QDR9wPTcXyaV0PgXy3Kixt/rUTTLPvRTJEc
zvx6guzqnmi3wzfFSSDk75U0T9oSRtWautWSF2jzHH2Z9e91UDhzRK85vq8uQKcU
i2b0OrNEyUBGs3PrtTbC4SREnY3NrbiKx0AchExejhCkCGGpzYgBrhn1DZver1i5
5B5TBkwKH2nfFAuWauQMQjl1hEec2q96VsKDpus2AHn9llPQCWyLTf9pdiSbL7ff
FPpRpWHl4nAUf6HjQtiOMUC2SAWq64PRfKfQcPh7daGAv9yxjWQmb/N2/MXoyHXP
hihf1uBXYXVVjQOIGMat1Iw9BPS2lYK5LuTvJqrMOT8VgcbOb3+sPItyn7fbSqfw
LvZSMuDzhhWidVFval076jTb/abxrumw6W0h8VVLmKZ6JJJEiTJKLAhBqhulIfij
YvFwnWgvCWKXB6uMhqMNVkIE/EwaSXSqwYaEWvuZ20OT+/kZdXRheL7E7RmtdxY4
yLFS8S7SOkYn/TrPSnQDqkpZvkB1fwc6OEfJfsaAuk1t+d3EDg1CBlemNSoG1rLP
xshjwCXElaY4IRYZ3mymEt/nESU0Hp+LBGb4t/JRATnG/zZH2RCYKpwoPcToBhBt
CjqFeSM0oxLJHG7a5E5YUxYdJtDbxvd6F1C5kvyeg7CYKlxlYInuFH8gi9B8LLuc
TbaGscJIXusRQdqdL3BlRCxootTvePCeZVJQ4P8+iW2GccfU6K21xLcKXU937Wvv
YbH0RWPqv7zvvjDxYmCqCXRk0SxFErQ8P3L68jS/djXCnag/tugkW98MDZjCXgbu
VfB3dzUG6S6M9K0aawmJyCG/T+Vm0TuQr8XSL9EoYDDZRgWq9RHrAm4UJ1qJGsyv
79IuW4LHOS75sA5KF8QjFFOirDb9og8jqToX/eFM+GPTXwCWdHeGf++qJ6tVBa8A
ba6AWhTf6vAJTQAf0kAc8CqdVlkczb+UIhpAoq98jO/VcwNFDwBi+5LV3npCRUyi
eqE/zNTRAVW1/3GaPGw1oC05kZB8TmpyPs8Wesww3NyVq7O1MjkO2oS3nuQRNymW
y6uipwbaTlgnnHk6luNE5bMO0Kv7qzYAHsxcy6wBLnA3w+B501UXV8093jMVk0QH
UpAPuywuY3RTt8cvfEptYP98CIRmy95LExAwdr6fWXnvqYVW1u0UPXlR71KgErsr
gel8sPqSf5d9M0CiNgYtpakgrbbuOfmvVEWGJZ41Nnr3ty3mmQsQmo3IZhcGReYr
Q5CN4ooahegbL+wiUrtKtjq0oDOdsti6p/QiuN86Fx9vG0zBs0/1U+UnYCCPwKUe
gSNeDvJEPXT8J2d316MwAOgEQKZn2XpGWKh3VDZQxenDl/B6Ze17KOZLwPwMofPO
rJ1PXctvzbgz2WU9Fbp7sf8CZLb/xeB2w7WbX6pmzR9j5t5L0bNUc51bce4wGv3L
y707aHtQhgvILOM1l5692sxkxAKRimv7Y1qdDhPFi1isDdPcx4RMfM9RTPbyICHO
vkGdGJLmM0fKPK7cTJOjM9QxPbOPmSchUIXccIGrvKsMMNamQJEilbWFDHKaq7jd
ILSG+845DOEZHC+m0mPnR73aB3CUXepy9eDUBqV/Ey6O96vB9fn8svfTOCScHWtz
sEcto4D8qmFn4UpXCnNV4dRIcrpxyUaDW9cHS3fEfhbEApu4fTn8VGGWKF13mKRK
8AQud2VPK8DOeuLXAxZkPxvuB2jPrp9w4XMbPOMcior31kItVu8eeuP/IXbMk8rV
xFiQ9+9FDNlgMP3ULx7MuE/jVKOoGlk4Jcsg2qFQ7HGtg37EasyGxVWhH8k0SOhy
Er5AYiNVklmWPeVjH6CYZHhyAq4/tr5K67gL/0WMVZlYdATRBEgTi1M1borK9SQZ
82YqkgVcBY0K7UgAfEipy+tX915botkP3duzOxs2K2uaO3kRqPh9uwOB4pYZp6ds
14Vgb4gMOeTV72DbWnffPjwVjRScADamBP+T1N3JC0CQrcCxsQZKUPj+qCUp6Oml
Rco0UGXVIFrVX8eYyZKqqy8Kd5417/u+lLTp3Jzb51aMtZL2wapLdNHk9xrvoPif
LgaKeU2wId2Rjy/zTaZdxZrmLJQyla9Xxeqm7ASSC1EEPAzwKPV4tfvc2wHmKJUz
9h9+VGzmAy1ESM1ki+gFax9FTT/XQ6c4NG8NxzbY0mYMc5hJyIbi51JLE1SMB4oy
J6PNa9jUeSskiy0T6gOLWylD/UDeONCJNSVxJWP89CMLqSL5ZxO2D9EWNTAXrUWM
xsQdMvhfhiEDcizsa7AgKltpfF7QyIs3ckxQil3meIUzveo8NZEFXcYWTMqCT9/6
/vN9gAcE8EB+jZu4lQhyJuYxz1eCIJHh0uIhhbN2HN1bEgWWZ7kC3YNUCd4hPdr/
lDlBxwu/028zxfbBjs7hezh/07I/0GrvczzwsWByDjaGXaij1Wot4/O2x4iHZ7LW
Ajxy0XlVtTiRwoer22xeXoX6Y4hxakXHX5iDd7EvH16tls3DR87/TGqTFpJo0Uh2
b8Qki2etzJUKv6Kxl6vjPQbjFsiLXRBpXPh4neHXdQxHoLA0JtF591QOhyAbUO4E
3UeIlfyArZJGTLdf4cWn6sGcMkvWH/yHQd9+kcQUms06ijf196XDv+P1w4fx0PtI
CO8gIcWKi3m6bRfQ2ZaQzss0QQZ74VTzcZE94S6rqgkWfZw1HjogRREZpvS9N+q6
MzEY3jVDueMmtHc3CeF6FL+Z/698Z/TsTkWTJCd1vgRQnzqfIbcmh+SaFo3o/llp
GH6tghTegP/A8N7C8yn6YdLqhl2spcSmT37MAv4QjNpbGUqKIJB045cNxwfZBDcX
NaPIqOvHcVZPES36qFsX1CpT8tMq4ImkcLtbB0bNxSVF24GEziMpV7wE/s2Z7fKf
kFo4Z2L/X9KdGEbYL84Wj+Y0WFBWeUL+4vZOlcg88Aqi+2yrNKnpznhOJSazLajx
pAdasEWbP6oS3Zumnlr//1VGbCTIBbhHvmYuw4LfJQxAXr+Ae8jYdKXIf1EoXcYh
mCoz4yZVty17dXOMxwGv1LTWHSt+zrqixZlGwUn1qFxDcIhx3nvvI8CRgv4GrcDf
myfr9gFE46u7uspbpFgr0z1KtGHtsVlbAHRaZVGteLceI4mOseOXcCa5tyiHLFsM
ec0NjKWhADhkcyrZvQqp6yKmkPLvFhU5C9redjt8RHy8IKtquGz10kQCqGkPbvbf
QFsbNnPSY695WNYwiCyoIqkN+sjl+Qkx2WVjzWTfO3JPQcfcJ6EVjOTyQ31eI9wq
DAtrgYzd1m57Us8RVw0ifoc/LiwQmiUdQZnNuwgxkcsTs/n7Vy6z0HIrtnyGKHyF
+lZvSI68LPnTLvDIhWfxBiot8lvGCZJMsmCzVD78H8rtS4guENj97PQNGIGUvxkW
bC/BMP3pafZ8e8BVNJvtwHFHiukqJS8S8TDiIY/flf/aWj79KdTsLG02hEV7xeo1
O0N19GSivK1P7sAq3NHn5K87ZhIbV+hMTmdfn7LKMz1GEXqqdGjIcsSBkk+Patxi
kSHp/LNerWNSzYME4SzoOAhs3oT0zrdwZ9zUicTObDb0KF+VLqUHBoBn4O/iwzi7
kSWPjadGpKoSlemAAGTGfI7dKNWzKDqOiXpYflIRXUKjC5iRzIZcOs9BCdaG5PQU
tWJVmb8IXrHZNJBSRk17BP37pbGbHhufOMFY3Mu+zs5b24+sDERDAv/BocACkKBZ
JzNnP20OfOexBpeOdXXMDMm11Lx4taZStr2tl7Sx7Ng8swDwP4FcILDaN/NGETmI
193xzvlcVAm08OYI8caVXoF5T0t/N1FjzC7MlXTiYo0C9LMOpK5OJI8ONSDBvVw2
ZXw1TvRHe+dovBzXGd9hUXQ4pUe6I3WFeT6Nnxuwfb1Wi8wM/F4aHuzaMdmdGMxG
Q4X5G2WvUIGKQxUZ7VHUsaGQi9cIbLe+MD70EFMXpW0XTC4btEb/jvrUqAraApkV
Qk3awobOx4Ly1svfqm+eS30VjcRX/PKxyw2Es9bgONOE0f3RsBp+8f5kR3vlcL79
4iw3e3/koLlf5tDclwlbPg22mmr5E1R4H9a+vbx4q4VAynVWxXyWMD6358IJZx77
pEo8iKE0XBTNAEsJhUAPfTKc1DkvUBLzvSIJ3kg6hhtCLoM16gZRw7fiSNdzUcnm
MsecOr4LHyVuXe9v9GheOTpwbkASJx3a4NzmvfoyqXTDVLdDXbva4/gwBtyaNHBH
0G+VerIsxexBNSFv0SuSGa/4A/uE1gO7A1QRZ28jqCNrP/iVH2At4NlHO1Kgqb4J
TxlyjOgx4bp8aQt/wTixhVx9GPHHXX3gElkO/SEYf6qjyn0kUHVfJlwPdy7i29kN
qn4EmQTXekJOeHnYqAMqul24xXVBYlSXyKzvTzn7qxkmaO9IAQ0JqiSMUX2MiJcV
HRKZQGhF3REwBF0cHzEoHTk8RRKTeihKcU/S52ee6V0wxohjheNkHlraQxmo8jxC
o1sULtwH24iT3XUXukyScD3x2v5X53HoEEZzlEH50CjkFlE8jl9BTqiPPwlLHjpL
xD2SvnLP7f/PfTEozhAC4I19u7eE2V+FpoyKhk9pi922B+rtIHTXVo2+eRWyBicf
NHjr9Uj5Ohrc+5gl5SZ/nJvC2z+8nxEcJ3B+woUxJ72/b6VmtV0rC6pPsxxPFjDi
KVAfmdoI2tfNa+NGiVaJteQxMP2piSe0JwAkaHBqC0kc0hJJMNcdN9/ruI7HgqXv
JUU9S3ZN89D/B4jcyO0cRaRVtfOPvpjaXKeyUjEEoYOKTwfPbeSxmthy6O8fa4Sm
cmJqJjnHWqwHWwuwmyD0b60W3Su0mA0JvprC1g7IeFEwvkZqxJ0qKIP3IytA0wOc
ugFIhM23rl0vFPUnzdgWHbSKkUPL2jP+ZkSvFD3Ic7N6lzJBHNtVgunm3rTUJM1+
87kx/IBZuXHQ2PNt03F5CAu8Wh5ELraEtm1ME155zMq58CPp8eRGomE2m4xgFLKA
be4n9Z9jNqidNMYOAdO+UqRfUMWUtOk8RylyweDX2os2YkY/fhHNc091CMEj+LRm
8H/Qg7DdMJZms7lfG2FsuxXOD/o+LAoLUL9ZMn+pmimoBAw+VuzBCaOrkCxqVmmr
k727Lab/RlNT1jydlLOQM4S5OXyfnbyNU/vn4LpW3w3e5OllhygtvbyQ4+QkRK2C
LR+gwMxTxOPT7I7K91OZLwdO7cOw9y88L43PypuuARlm0k0O8+CGn0pccwaKaN85
FYnUB9Fi+VfIvq+pf49DU4WoAmMBiMKH2zAPbSFeftU=
`protect END_PROTECTED
