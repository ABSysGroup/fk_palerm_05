`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YP96R8yJfdOECjJjxnwC1wSu3tkHgVV4A43Sw4G6PCkttWl7p56k8NfxaXQ2xKhn
eTr7q7eimV6Zeq8zRmHJAR5xgVIAWiRmH5k75FDPPoOwU91EtZpUvYMn07jUWySf
5waaA69Mc62Hv9+3VtGGgMcPgSbP4oEOdY7uHljCRwhNJLihbYYRrVH0cGJHK0jR
i5c0kFQzI9dQAAVlAj3oXiWmw7URHa98UvDQGD+5MM3QSR53BrxpgER9mfe+ArhB
665YpdDKexwRNSI6+rw2TkhCiW2fqIUdhciZgCOdIAcNfOlrlLVgEUgi0cRmdae7
Iau7xw2PJRxGzO/XK3VJUDg52MyP0OD16RmvT/qeFAC2t9QllmJ2YnwiwO4vS8PQ
cgqYzHmrhcl2NEirbBSMs1Qe8Nd9SkJBhpFllxcBqb5LS9AUpzqDvPKnfqrlDE69
FPJePHT/8k2qiKnHauX8MBjgS8CS79QpPTM79OGYK+kgZCRXqComPf2IIjOOI61n
TfKCtWT1qtgJlhaZZCemjUEVBjAFFQNHux5XOF0HwXQLhUH7D7p7YHBqurxz3wnO
LGiHemByT7rB5WKI62zc8CkDi8RUnjKKDNhhQv63iUGgKWhbF8GI4HYStougUcoh
FwPyb24Hed00NbpcwLdQnCH+qrnXG+LHo+c7HfPLrhqvU0vRweu+785chsHTGSXN
PFMr9hrrXyBFn2TGmvEI7naRB2bhwPFItiN5zju0azfiInwsW+plukLv8XXiuwNR
yE81kHIrfbfOmxbYdKzAbdZL6+Z4bYEX8b9fDORapl+zWKSy8ujfr5fvi4bwNhA+
nUfLcsROb9jkpw1jMP3/GQlULOSUACU7rc2eSEEwrdPdVqm7MevJY7BfeaDq/6zh
HqPly5lM0b1JiX/SpPQjdze5Z2lQUwVjh4gLo6yAmUR6C6XvCdx7p1sYViM5zzNt
`protect END_PROTECTED
