`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eBi/gMcb52ck2JtvUDNhF3o4wWN2PyUczJuCtxJvm9hSf0ihw4VnZ3/rRgU/SW4M
L/ePZYEB0LMTMVoGOaY/iLopIAV+xyk3+1gvEIGUs1cCQ3uHobDDIwna0C8jK9+Z
kS0ICqzzhx5CbljxC6HX3rhB95QA0sOSQRkGbcnlF6FUpigbBHHRzcc9JON8GvEj
wsQjVOn+7ixr8dwco0qYPyTeoezILSgxZAA2nlF/ygLeW3kDRc4jVTfxd1Ybx03F
RpVEmEab1M1bPpTJz8Rql6NGPmANd+EOtnCFRzva+iG1MelwMECV82saC7SLVnl5
EOAPcQRJRQoehDLBn1Kx4A==
`protect END_PROTECTED
