`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wtl4yyasblLKhFbn3E9boc2aUuE41hdIR72AG3lIQ6b7bq4az9R8Q/Cd6c7MQ3dE
AR8NLH5Vle3xTNQC14548q6BJHlrB/higZoAic8UfFsAPeMnpQ0nIMfCqdWtKHJn
rLgsQ+ZaqdCQYb6+v3P89d9ubr1c2AzCYBg/tHJ0lcr1XDxXizH+2nvxuBJueVee
MszKcOg5FVLaqE2wHcIY70n290VG3oCxwXDhMKQnMidD+ZPDdhKhLTdwxs7hSv2y
aap9kElsN6vfdP6x845PKii1xmPgUb5436ZwPtFdyhEnHmBWzm3RR07Hsi+0eBhY
YWj8cq7PTM+422Ii83ohd5YwvkCkqTeRQ5L5Lnsd7bRjr03g8QYl4QQdDXbCzRYz
i1AvSK2RtHU3CwlN3ynwM7ygZJ8uNPMXrphqbPgjV1KBs4s9NO3OVcdBV7eLAz+h
`protect END_PROTECTED
