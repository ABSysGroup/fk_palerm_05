`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ggm9knm3azNlHAxNmV9/V7ugYPiona3In8NzH7QfPjz2Css7aKkmEBut7HOw0wWQ
NJajs/pc2F5N29I+amPIv15wK/mCQeBUUx42LbhRdsIffw+okxZX5ZLICCZf4afi
ppl+yY0EfZm3jVCy0VlOJf/ZXUM0x5ETCh+9Vt9XhwGEdlgtnl10Oz/9hxUvSucK
s2KyDLAr1s7rr8loRgAanC6kC70ebEx90eTRkMqkGr5UzZJvO/ZBht0u5Z9OnMrf
LSRZxobZUr2f2AehLEqQzrHTaB/LMSnuJihxvdr5ETlIFjCR5sB+OdYN9KjVPGrX
XveepbjFRKSmNVtoZBTspg==
`protect END_PROTECTED
