`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3glkxrR71T8yfBKpmSIeneBMuTrxsGbJ5DOhEavU6KDHs0E/gfeus+d/Hwh3ouID
c3sMxZjvd3uEs+DEM4sjjL+MsmydNsqIsM2MNlj0ZJdmTaJJpKqrxaKuNGLR0DOG
3p7SfXvOJL0nZUZP2Fbm8e9/ckQsQ/MefHSMqZueiWypmLZgVg71aa48k0HqzA96
Ml+6ZBg3KFMfCAB5abSNHWBxjvs7Ca7plxMINKWIm+9TaCuzqOtX5DZfkFfBo/RL
EroVRrki6AqRgWtcKFrfKQ==
`protect END_PROTECTED
