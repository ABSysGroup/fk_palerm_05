`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
umSZPEDxSheoKd4bcSxMkH3TLs5idPBsfqDynLSQn21h/tadsOoFfQclvSTkLaDw
UoQnP2xhKHxb3rDJ6RCRD9y+S655bCAundVK/xpMlCd5/yK5h3s4YM+bBS9an+Cb
lUx7Q730NHQaWZyjafUQ9NwJmA9R8eJUJqexoI2FXxH+oDMX8i0q+QABECeOI8jq
SUV6H5lPYp5AvNUm4MSbJ9GM+FfB1X6xmIjMq5dpFEz0Zq9Y4XQGmBQ388kVrNta
RnurZMXAOHDyg5jdMHu7M3SFPTsKmdee4SB1oyECliAG8H9CVshUIvRyUAznSUhw
mmbtxDI2iiKwm+UO6bpjUg==
`protect END_PROTECTED
