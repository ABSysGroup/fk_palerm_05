`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Gc6O/nu/1f7tg6EG+3fVltjdBaosV7miItgZVJGQOVVP/kW9XR5Zh8DICvNQqlZ
Bd8JUE+jMeHMD4/MKD2bp4MVCQEOrsRcsMoGkMiewCjidAZWrORv+Qi4Ml1OqaL8
K4dUWjaEDaN50I1EwPdW2/zEQBVHHCqcHMESx2JO8KDEIkcJPkf9gXOTTCSdvnh+
qOJJb43cL5IdYg2DoPrepFqDAhJUeadTBTBUHqWTOLsj1KT618lCZcZLcVfkCmdY
l30OJBRNlmjTrBz7735Po0lQ/vy2y4zsqMaQoViC7AU=
`protect END_PROTECTED
