`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rjGa4Tfizes0pQSGfAotbjiCGcVTb/c2aLJmrMPveJZYaLW9d8n4u84xQTYMHBqL
MvYRf2kOe7tHNiEX6+jRXapAV0nj73Wa8PKrgFGD8zw0fxY7NLIhXfcUNne0vtTm
UBdTx67IFY+C26dwlQQ8h0rv6iBW9K3ZrAa7NMXsB/0bAYG3qkaD/zxeeuUKqxwC
DflZm52ypcnOL4mgJ85UBwaUcM/PwyZMCyA/WxKW65UP987Pax0zaVYmVUi6KPDZ
BY0VAXEInfpkM2cF+9ylYb1Ze7vhYDcoSa2InqJILFeCBto2jO8S/8+zuV37j8jM
LltMnFKdVnmLoIVLsrCJyRXqCZddeakYxLlW8sY38c5qCUhB9MgSZBvSFCRuPe+n
iE1B+uTC9FbjJRgmG7ig9g==
`protect END_PROTECTED
