`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SVLuyfJVccCWLX60iN7Yf17ZeVcN4d5ryZJWnv1RHh2XSjbHqyD2EaBT6nUm4mrU
tshRaxSyagh+if3EhZvaOWoxjCddxeLCFOBDmS6hji94Z+OGgfihtqaXR6cMKCJE
g1JhcQuh2Uk17TQHZguJk32+EVnb5VD4FPLVmLnk04zmQWg4mkfbrjaBudGYktjJ
CDMNITkglnelnL7a2FtAl+pRjxFcjzz7CyPebGGzPqpwIlDPm2oCJ7FxC8d34xY3
fP4pz8yo5pbFEwPn0Ncwpsgn0i7OveuyOT5MTscsjB2IqlA6aBQOnXGdmQr79umJ
ZUgkDORCgnDQQFBiAXUYGc4Fn3NLvrmCBsKxOd9qy7Xt9FQ7nMTOOGfsApVfkDBn
5xKwFko1iQTyxuEIfOFarWb2YufmaMNQP2AI4olvZEI=
`protect END_PROTECTED
