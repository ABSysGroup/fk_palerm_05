`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p+SJ6q5a5EBcQB8aLybZUo3MwAailCZ6CNoxwd/4tB17N7zWjCHy0crk2jV8HAea
7thOllyWo5wLEcqY8fA5uW/V3U9Kvk+NM+LKr0Sx9QB7MQkoJ3+3K1SBudMLCNvW
VoRxwwW1WYrHJJC/u0qaeg2CVnljVUmcPUW9LosAn1YAdz1HW/ArURm5owHJe9vt
FEvBDqSu2vgHa0lFzq1+W4l/06YoEyFlT2FJzT/BXunkioh0IztphD68G9b9IWKP
PRtycxGTT1BLv+adZyR50YM+lE+N4o5JkL5YM8U5dmcxl+3k03RZzWn8BHcygoBr
w8tUbw5kpkfdWqYzqG6A71+HOOKfrPKlvleNUSiVVVOPSDpWtZ9oidebhFLIlevc
E7eZ14QbQMQDN2fKnXTu+mVkdSNecdGdrbbNNKLaGUzEby/nINd4bxYcZULhhM05
HpvLxcBfWFJIZXovaIkBCwPrgRPyEVn4VhHmL6lfw7PLrCMqjYqaq8MId7Wb2zUY
xztMVQLIu6rwJjnSfCDM9Br6b31SoYtzW1wxSubJsdlddwkjnLfREZSj+vwDmJx0
Az8cYnVBoQsopiwHgHGkNlR1VqqjMtsbjlWmxumPZyPD1+nkOJjVbQWk1ljF5qWg
vpa8E2cvwuv3N/DgH6KA8kYfBaafdvaeNJuWExNK0xbjid7xS9rzsQEqrK8mWQCR
yOtOtjJlxMdfpSUtnziFnn5uQeaMZlbObunyeXIhXnGxxMiFSJL1r2KYcR/+NUUE
GITsSFBqRzRyHBSh8vhSl5Z6atDd3S7cf+Ljz45tvmrrMOzcWkg8Yf/GayG1RGXJ
LjGguhwvr5L7Tl7/Fmyg4I89opkZfDy+FK+geOS3xfL8xpjJivJiJ6Z0DAJ3CQdp
Lf6SMg8R4/GauM70IciUlJdHntm8nof+zZtxXoFln57sj9KcsDzWYeaBJDplj5ym
PVdaPb6z3Jo+mIPtzG+MJRU4PK0mqB56YzAMJ8DvKNRQOMFOvV9OxL9y/yhqkxFA
Xo2cj3aE7SfHwOjfPAtdt1MyxYWgnaYufr0Zgr7s7+LlfyR+OJAnZAZobmQ8MEOA
l3xDjOrgj2oEUzYxR3t7m/JK1/MdAmF/uxhndgaFXCQkQCFkf19yl4kZsNecCWdF
HnyIzx02YgJEh4+hlDqtr3OMACPRiWHaTwuswjBqhU4gUCqmDd5ogydulhL+2Ngw
5yp4Yv7KOEdOot34GnicNfLsIt4471UDg7V066OUMQ3KtC/Z45gt8V+lHnDFJMPI
QmR0TlJxiyYcyVOabPIOhfoQZZYyOm/0uxL86KhauH46BvrdN7gwXhUKU0Ai7qmi
b9NOMbdDHN8JlLnCJMZitz5qbGqDSDkAwTutXqROV3JvitN8oU2QKcePuSaFxcgd
+1jXGvaCqyU6FLDpVLX6yUhZMYCG7RzOEExHxXOztdhsJshueKAA/rch/iFn/H/G
2NoANXQ2HdR7tJ3i9qZmgid1CeyhCszL9tsGXDFgiEES7NgcZ4x/S4tfEEi58cgg
wXMt7J0FvX847b52ax7rPzJIZ8VAyH01oUms7oyckiRFwjX+zPe9t5pAceu97KrE
MdigspuMmD8O5lOE0b4lurqVvms2Tk1H+83uEiNXTowoKar+oDKx0nUsFUTSuwwb
B6hDBnRpEkZZojWKA2IUQhx7cLiz69ddQe1nz3obdjEyUfAJcfJ8IFWGf47ihQYh
XPl+xQGlPfgFbmRq+WUUkULhp7pGD4yxPnyu76AgLXcLOmrsIn3DCshVK8HYlQxT
9YiISO5he0kzzeOuzZVCUkPZB0p0t6ze1AF0vTpNBBo5mzwV4U55P5Py/yeOQ+oP
f2N1NX0dba0LeaQMtsolhQmoOIZvChoxVfJ2lmOMSgbIZo3y/KznTAyTKaYZU74F
`protect END_PROTECTED
