`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XWHCMYRl6MLwzqiP409Oxh0CGEOfQN5cGrqG3sEVHFh22sYxYbTmtNH5FgFzraFt
yhgiX8lac2gjUVU+HCPw/jnrab8sMEdAZh6fV7SNTKxYhOzipKyVb+hv+kfuqDIZ
AuF8bCLUFxpjFSwjMA+W2ohtMK3JLk90zbUNMHEP5kE8oPtP1B4CkIgUUuf1mGlf
BH93UIeUOmVWgEDBa5CmMS6hKcFyftwQS0dnsOVuOaM8ZOMtPRtU75fFYj6vtDNv
L8zXT2ZqBFlaJ27/sDb6KdfponCVUh+vcCbXI3MBeZyKh4ZRAvf65AhJdWYCSMtd
KdH4VUn88KlafLdHAA07yNzow88phLbSBwmaNx8I6dyEsaHnA1OJq0rMR3UgXNad
wmJtN9XGQWGQXZSMiYHORlX1NThjpDHXtux8qPIjwFft+FwW1ja49sRcA/QOqasD
RBJfZbijGWF1w4otRJu0EwWUyR7D0pj6jG8tG1AKmNXvjK85krEu+sxHssjXIEDT
r02RPTbCr1A3BZumZl9yNIGJVDJamDVj2VeeK/mgHCH3MPFXzPQwzv+1+VQS8AJ0
4euC9TQ9suLdFFqYmF9XsuJ3LJFbiinLm8L89HMfBtOnUIIX0j2HvzuGCX5dmunp
03DqeYp1uQHUFSxXG2luuxu0pf/Mb7TJMZHjwvvaRGEHg1lfCr8sZ7F/vZB1bcAb
veUPMfs5ELyrjOOdu1ub5PjUAOlLBglQ+A+5SBoR7odfOYx0hwjnuDkSwDNuwbAT
xXxZ3UGwURNia4eGFjtGNyqdUA/52aCcZ6c97Mla7wZ06VQj7guo9CQ0fNR3B4cn
48dULeIFoBtZW7tnXmXHMOhDkYB2aDvmmlrvlKUlUxHN6mTiDAEEn7nq9XTf41WW
HVKRAcvnotnIPhbv8LsgvyC529xhQAfu1glxCCHUvWJktAM90JYYGim7sdehmZGO
W4rV+N6KHvdYnSXYZo5otg9zRbJta+B6GPudd5OOG3Z/rxKOOqSR+PLY/Lm/kMMa
YPCbugg7yGQeK1PcJOrN7BOe87bFhQGuUrJJYqjw9kPns3EHcSTsLfH8ov6SKcLz
J+AbchB2mhcGtg3TrE4WIrPuTBQaoUzHL2cb8bI+6ZFtl8Zw87mRw+wrnJ5+s2Mp
YysrWID2t2MGJLw6//IcrVzzLYRDKDWNJ5oVlUANkJROrIVRCxcWwTQ+yBXk5I8i
AyE3IpI8bn6nkgRa2X3oz4mQVmwqRVL8XsGOReJFGcTbTZ1tNGSLoF0HZ0Xs2gMA
46T00kWRthjcIbHa5nI5cw+bTUjVx48xAbBPjPrnD5mUBqhVWi4sXRwz7jOqx81/
eqdegxH4U8PCVZbAb949CprVvmCMD/GuTnuwNgqzki+osTakhEJGjEiUII/gIgY8
nOdXdeyRk5SMNqGACE8PSAfKvqZZLSCSIwb/9ZLPg9B0m9DuTo0vv8wz1SKAaQ50
n/YNRF+0Hd1N6WTbDoNIGpSwtat4w/pwAYUtG39LnSW1tWHVD0st1dnTwGjNp0oA
qP/ALPnRjldhvKgvHgG57T2B7gDRzbsU+s3MfKQeXs/yvDFvfK7Zy0g4Gw0aNhPm
s/jsv81fBEKFzSI1rjUvK51veG9SOGV39XbIWCk1NkXA1+rLGbaSNBj6jQWq6Oow
BIdBKtlgm1aV6/piguLvVH0Xe19TBNSdF65lOWCU5Rdsx7YymLlUZGVFobGEkjQu
CnoiRV7R1cLLAmzmxlo0fKwbDaEj57u85a9ZRi84zpkhRW9mu/HaLPiEPgGWOWL3
gb0ZrmKaLbQZIThxF0UP11nbEEI11sYj1dd7uedOw+EopyVDLVyHKd6T23mlCpqc
F7xKlO8P/XcPAlgehAzrvS/0nCvRqNAxyGs7KJL+4RZOa/ENO3ivpHQFOBiJ5u7p
65KQGYwL+ez6JWGUpKMM8mjnqB0/f9EKSXnJxCZoFBhO+JtUSOtWEey3cmksjKNu
VkTwR+tINr78fJR3+rh43HQM+Zpf+huQF5eyAX797d7LKkL5ZXXcLgdZZypUyR6y
lFDO1gE24Wl/HFpmCzf3dB9xn+h7M82YZOrVQ4vn0k4/4mC/1nexb9e8T64twcA0
lAGtnAgSGUkSjyAOXgw5FPi1TZldUhbK8/rs57KZscVxPCg/dsiB9tAuH+y7xBOA
GBpm82S07lg3XeJ1Cl7hP64DtZhgsOgnHOZ6rPSIYOBkMtmn+tpVG3QHb+IykTfp
aBnivfsEShEh160CZtAcl6WDucBuldawkAVj/f2gqtWOGGFouHGKso2kC8RpYrAV
JrU8E3LuFhnT1Jxj3ouLCBNfpE+03DOs4Xq0EXeR5LJnapRcCY61RgBGxMQSq9qX
89Ft+Rfxkp+qSiHgnG8HYtyl4BDPL8mbn4kQcX6gDkr/ud46TFlYig01Qk1leQtV
j7g/Wr/0wqeXChMoU9QTJwTkQ4FrH+9bG6XMbwxmLSUBsuJPM98U/2mUEkD4oPVr
s/mL8E07lxUsk1AcoeTgJVYGJ7rUomJORwhUMW0wrOXkENSwiLGDBHFfQWfiy3mn
h+t2SKbcOPkqzvfz1WZ/OkBOVG8FGFFXh8UE+33kAWFbGebvgNrNaInODNNBME78
1bMh1yghyXNxZbJpAzP3ohDJ8I4kc34MNj/vjaMHaaq4Detc008YnJZJLXj7fiFL
5aBXpZezo7Z2lJkR2kkfUjqgFkrg6yiGIfiUWr93N4xoLfHbh9WqDTBhxSHOG0sT
znCVgF4DaYRH7eVYcSmXkHL4UAzDr6nixBWJ2yIusCbNBkCm4CJlnF2VUpeaf9W/
XaGDcDQb87ftLv3uQrCVT965Kz0lHSv+ZlUtibT3mhIvESEqVE3sjvjF8EA5AxSN
iuzhqiw6yPLlPS0JPzmZMWAHJcM9bG7oJ/pi+Y5NxxPHoElElwqE0APNDckh2B5X
DQCNS2a3LNY3BGCT+4GXJRANzEi7pQS3zqmFrN7rdLmbenpe6/VMamM46a5BZ+n8
8xeUe2kbLihYHobZKo3o8ULp/NjyB8NUjEK2Q4Zp9oaqAGQyMy8OJ+AzbHk8jFbL
xftpIaYZ3aPwqp2uxlcRJZK5aevdJth01z6K1B6uPY1xiHyb49GvNuIguP8eK0Ua
svhPxZ78+vVuNo3NNSaHj2RacrZTbQ15+MG2FAOTg3wfnRISn7WYtxiuDvRBIsTp
OxLloHxDoTw8WfLXqL6mVr6/+nnFXllusSMoDXvDS/IwyeqzO8n3UW+Ar02y+fjS
uAgde71GuXUPv3LPQEWk/1ZVn5kFsFfcVe5mTt5TSpDoIpvDsovaDIfU4rLUL1js
P3mjPvE742pS8LWUGjkaPLPqu5fik760PryZctlgV29orNaGbVVTC583STJS822a
/T+zOjjdianw8ZFpEWwWFKITpgH0SsLlapUj5pm9P/X+IWg+qQzrUJ5b8bF+DWdK
KVBuXO6d+aUXFz1Fm5UFpGT9HFzFpKsqRzQr9brdjO1mzBHZSmh8gdolR9NXigkG
edykZOR3ouqxry8LOfSOYXfGoBDriU5zY0Jckzxct4OE3cYkfg82XJJxkDHxjLl8
23dRq/YtFggQ0A/Biuv0yp1m2BvEqC0LSkfAMABX0M50eW9XwsnW0Wg1fQrBhrbb
ZmWCJptU8MH35fRvq8TP2cFAkp7W540p6TgFEtDWksQ=
`protect END_PROTECTED
