`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tHfmWhJfFSGQvEf9A5DO80ddrp5u7fUuNtqLEuuvn155XBjvlaOsBz57eiHCk3yp
ogp1bBhtcRE9Xf3RcH7MPYZVGokvnOPiEbtZshaNOPbJSeEnZ3f02WwZIa/OIGxG
6HoA9mNYbqq64Ekh51VAFzSou7w/ECeZ8GErZzgVoj7D+/Bk6IJhCEmyIAcCzWy3
urChhDwod1YzZv3TCATEAK4hJD5TrolnjOjtdgOqj/570ewo29wnzFC001o8+g80
zdvioK0A2w/Gd99+t4Kwqn2SmKzW0VJu7VlmC+IVfbe8P3Nf4iQSFibd38xqV7iV
mWeGTC5eRz6/sdXa2olf8nWCiaCiZ+GqLkGbFiGDaGTLrtaFTz6bwfRVTaGF40X2
dJ+Uazbm9ia/4z3iH0a2uC7pdjWa+1d5yKAcvWwOKu7QWaTkKkiig/VeIekL1EWv
0kldp5Fgs2kb7MY8fleyhO9b6MMinnWCzDhc3upd7MeuhxYlzLXuuyl6LDaoviiv
atrqgsuVxjQwxSFtLvxL31TYcZKRCC6QXsikx1u3zsJxWMhTlPO/DZjpGfzDQJU9
jPoe2wosuec1M5ayBjgSaW6QHvlUnZL65dyunupP2kcJGHRcZcyp2fJpG1p+JQyj
PwhUEUi8ZkdxIa19+vQpimlDomeFaJnGOJwD6jsWPEzu+3kbYk9UendQUYgZ+A0C
z5VQZUuO+b9vTi0Jv2Vn4DJ/ZX6NsBK8wG7YGNQBxgw=
`protect END_PROTECTED
