`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FDxfF8SgGR4zBUYbcYndymcXjr7Ie70frW0rHgguk5TCG0NXuvZuZGfkXoGB4mtR
se4JV58tFeJsDMZ6a1yjDaUXiSr1wv2cUZP+ZcQ1sJExqfpyeSavd9kD6CEHDEry
Hat2ivhNDO6vKCYJknNVPP+RI0t0YzP+mZfkeRFITL/D88ZaRaoFEAe26gCG4X0J
sdDeDgHmwGTRE5JfHpz4VTJIR8+FUtHpJIX1sWVYDye5hR6SXKIMeUru2fttQisz
8tN8+XsmbNlRlp3oGekViIOUxAyiWF3RhvWmUKhNfhmXf93xiiWnj5A1YFhvOKbi
mS39/KL+HzDxSwnfqr27fH55ijmLpk4MVjmvrCNSPOX+7T/eUoE2sMIqinkvHOhz
aaSRNyyzU8ou0bPCPj6ZKEGWzM7eyrmYxLOEwXvti3BPZKX8aPOa5XDK8UU7J83+
mLIIwUqpIdjG0lR6FahDKHSiubjKcZUZl1931HKK5FTjFZTuGH+Nxpy7lhoD2x5I
Up3EXd2rUq8CIpB68SgqL4VFiKBipfX5ATw/mrFJOWWA4laDmMP9z4P4Umi05UIm
eB6YIqJTzUMXZVtwXBfe5ASwZzH+keD6xst/zk1bW8WmnRZZXbPeAHspJ1aI5TyS
svRPayal96cgQAF27rZjUwUjL4aHBDvMWS6I09+H0FWKca2Ja/+caeai1cQdHe4C
QoJPulXP7zF8oY21d7tcoXQfX7unCqTtFjli4TuyUR0g5PywhgC9sFLAoQwn61eN
eBgxDvJF7zHyD9SMCSSUP8LSbV4AnpFPhW6I3Oae+B9jTQ1jAygAxpQjG1YOCPE/
BmMeHN9j02UECvlPcmeNvdq2rn9UEjkQwJOPj7sf8R9RzwxDNFG7SftmNPo24CEK
4STKiCbKWRbGgYVrv/xspfBJJ85G8VubkDnoISouCv2zMVEpvqAT6tB/er3mXqmL
2ENU0vm7nf+QjbtNUm6PIs8FuGnQhDGX+NCkMHYFlFsoHWQcaNk3BPQzhEn6oENE
1+7FYWaclgFsigY7u57Y4M/TqtTh1TYWP+reCOxaito3kI9rImH9oSx+wPDtBMsO
OvYahHTZzp+FHe6Z+9xoPad14NFFidV79SlbL6DvdsmdfWiXdptHQpPCzs9LN9AR
rzTdQnbWize48WDp0v+hTIYsnpWl6utDSRV9M18bA/zXLbEUmn7hUp4n8+8eOjlX
1XCDhmBbKe4CEb5D22v1/9tG0ch1U5sfdqFbuypQW+4ZVlVlNGsRByp89BROY4j3
WyTNofMYrnsIdFhSNJqOboLCwr1PLkRoJ5H6OOmf+0uAY00uSCfntRaBGP/Lyp2x
8m2GOBnijBzbwvUg1/YHppaJ+TPnBHxK8Ds+EyEhjfkDptebaAvWXe3AHaEYBLyO
wPVRDUzcdocAACFar0/cv8yz15Kr3wfRAT4rqtn6W1FGmE/5lMXHHt7IB3xNrkk1
DkH/pqrj36cnhF0RqNWMRe5dCNCMACS5p7jQwUVLPIu0QNTxpQrle1rwH1fLuIAI
efHOj1+WhVaouHZTZGwBQm35I73oQNctbSdkat9hwlVvyQrlIxVTpnvmUCSa8y/o
FycbVGOP6GSXTvn+0JKzT1aYf8LPj80yjADt4P+eggBz7z9NFa4vVuKnX6fsieLi
7DSxOhh7miHr5eAuEzQydePfhzzxEHEPicl9AA5pm2ES+IBn7MgzyadFkv75qCmN
JZEwhL2/iXPAukNaEKBWqMpA71gcDqcX7wrFhuLndJJ3eyZk3Hl47MCHlK6JQh7j
cR5EyScx89rKvqzEGBtnc/9r5VwysMM/kSdKg3/uvp+MtZ6IEw4wSVb3bwUESaaB
rRXbKMfnEa9j7uBJmkWrZhdWscMFRWjcK/cct8HRBIvn2E261qzQ/vogOC1/ejiq
O9I0/rv//+F5uR5KGbeyMyhNGshwW9THPLuSM5MKDRN3ojDBWfdcZT+ESErRpbvR
vNxaLLh1h9IAIaK31WSSY0Q5DBpAGEzr2vs1OaHZ90IZmK+sP/BAVgLo1LAWdtog
jTrsRwLCsdFurj52NXKyvg0Z7LvyLroY7puuVgidID95yfTQpDSF0OvjqnRtnn19
8ieeIVHQG4FGYHQyLXppahSpLbZEzeO/FFYm06LU1jfG78gf/+IWsm9tzebArXR7
NyWbIlDjyh/ndUDiGTY8k3I59rdn6rCPpsCNDCAA2KSEmCaA2+G73qsTsZ5QpD7n
MwbDMKUBPWW9E4oniQM8fJx77l4NRV+XJ7WgmZpuSz9RdFiYP6Cuj76hl3t+UzWD
A362Qugt6EM9XSKPUxcnI2GvPhxOe84AWHp9QZ9fv/8uiyirHTdxYCV+te/Zns//
Amlpbuh2u7VoP6ZdXxUNxiClFwJQb5xZLUkzXMEcd8usdkkRfueXSluT66R2Zt7s
LzO/xgTuy4ZVS810ZSDTMdXRkVUCr3l037TYIbHkMw64QzAjTwLmEdXcVjieb3Mn
+udmSpv5gXXfcgyDIvPP8HvUMgQfiCps8gQEKL/r8OyUMUP/YP22JSnTPFBDi7ko
7QXs+eUExu5Ho9FZhXR7OwOqAbItJoG+5gvF53p0ROSyW5r0LHQ8rTug7Znvq7NY
2rQ6+6QSq7eGw1ad2fr9S9aAq4GMocIYs1oXwz9JYsNEA+AsROKnyHK99jUB2mXM
HBYPVTV9OwbPo26y5H180HbK9ZWnuBqfYFIlPZ6ui1Q=
`protect END_PROTECTED
