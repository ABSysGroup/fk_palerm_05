`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yYaFDB7tEjpIH7il2F9RV8E28/gqLwAT0bk+c5TFeEqifyJyS5RiGJjlLQ7CJxmZ
fYJlGQElGBZm3AcCE4g/hPQVUWgQEpKmNnoDPN1b0VsW4NxI82vnREXioCVS/u9C
O+lpEMFsi60MCuv6a3xpThciApmXFZYcYkZ+Fk0Uv5n5+DFAwQKPjq3bj9gG6mWj
2iPpCfjJ2sCGayvstIEnLEHNps6hmgSrAm1lewX9FN+6gGuXzSEm5C9I7zSrFD0u
qxw0BxnpKr6WMLfIQACnElkvxFd6pg1faWRC9z0T561rVu2U91pOij7fajvwfh6S
Kxc7VYKwyuIrGaf993+zqhZe2jBRhJkSzn5AzkKshDgNF+Au7ifzVkhopOn146pP
Izi+jlmlwoyYzApspvbo/Xlt0uOkgzlEHUvuAWOjN6D3kI6eVx62Cg8Diu7fCChu
wI3IQSfLmKKBG1qoDwZswkUUjcEvQMDNl09nmbK6aUM8kQJglZylq7g7Yoqu48i/
S/ZTttfzUvmXOLsOgpjIh7Nhylhd4vC7yH7Tab/Qr99c7Pq1usuF0a9jogHPsTbU
Cmu2oMokkIPZ8tNPdqDdQIphUxfJkAfQgQWbIPP+uSY=
`protect END_PROTECTED
