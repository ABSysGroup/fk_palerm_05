`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7aIBm6HxpWMsWPT9PIEX2voYB3i1caki55vMTYoZBhKmi6WmeYEh6wsqY0aRow94
Xrm+htDCZVnuR6z+DU6vpIfFsMRKCYOCh2O8Vj7TT9xVnzIpGves1FOjsYahogo1
HWF4N7NFTZp0vg6n5iw+QQAeeTbW2MyVAj9IPbF5+AA21iuF5EynDVh7feUV+Sl5
jFjFOPAqDsQip5lh2bOc1PHrr0sLKXkPF5Kqlz+Q8+NAHEBV+ZA0HQla186FMibg
E+unL04HUbYV0x+MZK1QqVI9gPWLkC/K19BEsXELGrSikjgIfp1YIOIsf+RomzSq
fmCl7rH1K73tjoy5KBkakJzG83nS1Xb3mB3gk3kxAah7ZPbDtu2DqHjOfhisv1hD
OPrEXZpszONIf9kaU5OW8MTsxtDSszoMi1K5OwgjmzUkaF2W1RURyNnm3X9n+ULf
0LU9gAWC85bJWxZAVUavEkWZ5hKjKpz2sMURIdYsT4pB8RRhdFb5lMU3hwScpaPp
Z5KcWSWvEKuoHRuLVw8W2+mXicXuZC1TiIUbB0XLazK6Ve4PA0rdvQwa5xTawNx0
wjNLnADsdDpwGqTVYJdNRw==
`protect END_PROTECTED
