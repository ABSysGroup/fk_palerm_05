`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ISQW0XJloVQTgK9+n3soK5ONVpZME6mOOMon1LF0Qi0KXUCiq6ocq3HLFTr9Yq6J
lCXapasnXTEz15ZN4lLmNhwCio+kQGHI77XRro42e1wx634wOt7qJwRJrMyVZoHT
BjwpWONzHnYhNgBjJK08NGhgf8omnxiR4ZrqlDcJsfeLr+/PsbuK1e8Uqu5NEpn4
OD40QE31q3gq90WbEsOW7fGA1SXeaXogF4ArJ6saklMAiuxGNTPDXtz+ms2+bulx
yQDQC+Fks4wjUPo3ZtruqtTj6kdr0wUHQZ3L8pHUH28PD/+psIj9AAOJReOtOPp8
WrnRKCpXaUYeUYBw9IDo5AJL2kPwOiyZMlal3kdAQJnxdGmn0427lLW/9zQ/tc/t
XcxcHKSstGaqN4NTyqQh2nhxzYXfRePCAZA1RPCy+4MfFtrqBL2cEkqhzswCaeQM
Xsqi4LlohjLqGQt9Ct9JJYXZdfN3N98DiU3lcLIBw41tAH2gSDdLzymf7qj8kbe8
MgWH8Lu9rgVj3neoJbIWNyhbfu28W8umsoYKpo+inPGMYVvy0LSInLlos1OLOQwW
DthM6BK9jXg3kVjBPu/fCiEEbXREyXs1Uw6nHH+8/yk1VQ38nitfQTf4g5M9+TLa
3vLPCLNVboC4NZQq4shxNollCo5RHf1Bcak0JESzl80MQIuCVROOAsmggV2lhzcV
CV9D3xzY1A+/aOZxxX16cHbZypPaobPIbhc2kzeH0nbVUOHzQ0RBB9NPBt2h1h/b
jEQsds5ODit22fY24GtFxo1Rnd49vofvuiMAhTzcq6YILbwrXE+cE6mu48sRyiEL
F3YKjjaj/3bu2EGzkbmtEif03QmrH2V1tmef+XOho2uXLeuK/17DGW1DsgB4a/TS
gtkFm4zjdJsE1PjN5DyWAcuDH54l0Wjr3gJh1V4hgXpbOYrhYo3dXR05FRFTi06k
YZPpMIFTSphtpmaWsZX+oe0aG3WtJRU1fu/JEanJ/wvVmVEC0UJ0D/QcU6g/IICy
5i1mbZ2kNKwAiPPU+F6bxVj8Ek0HMO8TRwfkFxMMJ7YpVOL3o8S08w8gbcPGtdBM
um46c127bmc90UgPgXZ4kkEPoZtV9PcUmPvZfbPWOjOFVW6oDqDjEGHt3mfzmMEq
7UIWJgK8gzwX94E9LqUj4/4uKYSqgZ/T+OdNDWPHfq0MP4PuyE7uQX/37hjjwg+l
z27e9t1yBai/D0uxhM22ii4p/LqKNAnDvHTDFa7AWJ4CbPDLmcXVEWIfY0LT82K+
3ZzU+T/fv9YbPI5TI9OEzzdAmhpgEmMS5G37eoWuqonvxQp18oViiOC4InVi0dXs
cCdxEDEqIMoslJDyOadD3fzkVsdQuQwD0BInHIuoFzbcNOk/LwfZoQznLc2gwMPK
+WnRBBPIDAHtm0h87eNw0XtOQEx4yUSk3P/RA6OqWkkOH+RWkkjFcWOLgIHLly+k
Wox7zL2KZCBtKiHwkYe7FvUgIChuMXqQf8FgbE4qm94ruNihlfhHvX28V9dLlnFq
quH5Cas7o+OlWDIzUR2BZgUQE5VV5BpRvs/HZTyjvK2pvX/PNwOZrQkqg+HsyDa9
oXkcRL0vzd3O1LqeeDvI0wQLQpXkfJkjjXmB/S3xQhnZRrd/ZSUXBgOGWyxJx0x2
vDvt1nlj+PamONwbKNMN0QLObqj+ui2Pr6xZnP7fA8HixTZ0Y+2nF6A4h0CLgLgG
BWLE8xCErcH5CMgI6Q/iaB3Qm+gnufJEEI05b9Pbd3hq9Aj1lizIEk6xMhsekY22
oonpf7K+BvVpzaNDjR9e8ONT8SB56FF/JhvbN2U4PU9TX686z/lvIins4falp+VR
EVBW0uhv+PFXGl0CgruktyJCYfTBojB5g/CpAPFh5vK7EGUile0UZVoTUfmSKwqh
i1H6x9ulvlDcPnVditjnMmDXqdBDT7LhqOJBuY4LyFvd+MePnrwOmnUvLoPnlZLo
68lrYME4MckjQd/MPQ80qNEILEZq99fOS6ZW/TS91i4kGYOMTKy1hTgv+ZAHS3Db
Zc9buCshCxRCMe2TwV2LY8fxc+Ucr6ym8H4rUQygNG1JTdBqcxiN8IilEnA5NBDy
aHVsBu1GuAh41U3gQrDi1X1QuPWtXku9KlSE/4KqMq7UxodsJLa6OubNLjOfLATE
2lxxwnZO6I1d4FG6LRTSoLKe0rqbc+WBdYer/IGKhs9VQtGDE3FW+76h1njy1kVd
b/x4yQU4UabfigJXl0EswvIUIpHVL74jj8xo7sqRmsCDyAHT14JYer2hAs6YFBwF
sFw0ShT71MDh2BTt2YCIVIXP7EUkmRKtjJK5luwnXSBfTQqiR9Wf1oJ5oyYFpRU9
OX3L0u9ZPHdV2cXec2DEnse9UmtWK6xIM81dDBu/xnWKl6t2BJWwufk2+WsMiZjg
F6yf6gAHAm7uWuKE/vQ1tZiFAaCx5+6h6kaqDKsGSwrqt5eSaaO9YTsVxNUW/p/y
DFywBzVD6sEW+dtbmObsXQi64IXICTZndv1yyZMKAssiddeMsnyop4SCiX3OLpsb
bzQCFvB+La4T5M4Wy4Glc8BFe5s2lzQDp3P87XF84p+Oe+SjQPyCMbKRpFBuQr5V
Ywfu2LzWG9VPmXkQTn65CMAiVEkJMlsASP/E0eIJX4OpqBzRHPxE+XNN+51Ya1M5
7OKzyqMHAHvTnxusRjCneTZGO1jfliyZPlcJqGaIQWutXp9MBRKKp2utjmanDFC0
TB5sKq13fdvf/Il95yy+wT1R4nyJLJYP/A/EZ+D9u5nz6McMYiGPtazkLVpn6Mr8
f8RIXdTxEp3ZI+POx7diaKwbyJp5bzllGZt4kb+sCJtbtwM8LbXMF8uSEhha+cxQ
5RMw5xyYwCwNplDcBPF05cmMN4mCfi6k0lWs/HfIUFRQTBLOjyoaJu7pwmy+/0BM
nUbDCo4UE+ACq8s3oNWrHx1UJaTQDJGErB3tdvhTy1EdEtn8rECvpGmCEgZUjVKe
4NEDBD9AERYnwPHwrRJ/SXAkzswmxwzuxt/maoF815N4y64sLEU0Hg//4Xw5Tqir
FdGOG95QvpjjDKKCQyVsvVeGGtyxhAjvrA/qTKr2MPbDUafiUHRhb51JqBt2LBRA
BSsU9JMlRzXBIuYUGwNab+N8C4iBbNbrE+6U3KdK77TRvK0MrGKPRL7Fck5KTyc+
GYNiiYfX2J7C3E5385xWj8oQE4JEAGxGXWXmsEZUITZXv+bP07ZLFl5oO8P0di0h
ZfyUdR/iNMkKMlKyQOBJPDFUPpPmfaQ+XBX/BiUpQXqRohfTd0SifEpUCEhqpssv
kF/JoiLckFN9JITFWfZZ9V1cA5v+r1XxJLQPVTDsn4JzmphUoJDcqBYieGh2Sq0a
C8VFNnekJkPf0aLOFyqYBcoXUtyef8Mno5SmLnkXqsXPb2EXbs/yZbHpa09+kaki
LsTaKToTBqOoMOQO+MeGdSBzpxquWqVGmXkO/yqQC/kyiBuQjSj28DsxeGnYP9Ds
3rndHw9CqwRAMI0bpLqgkRfzZR7zw/lFPDGSyPcsT1pw9UT+w6TkzIouumoxsKN1
637gG0IlCBInytaw5Z3kLDJdSPg9ZbefmkAFf3aKMg6LMy1FFVuGL9WP7b6Fdem2
ajVlGUCh3ICyvERAr3a8YrS+WI7sTwSudRJ4chSAjywTcKkGze6JgMLKwzsjSmDV
yHcJexIhu/8PxZ6DRoyOUuqxUBuOGghgVFGpicHJt9gHQNiVCqSivLyREFWjcxuP
9/AhU+uzqd091VAW/AwguqKVgYNG/FlxQFI3gh4AOqa1KvJfkf2Skufwd8qF7Ape
Vu/88ujhZs3IwxGJQaMf9Oy/5Qag5cTDpJdvFFR9F6CGjT1oKvPyPfmxkhowQEdW
24weBdZ9bJLCJCIWKtdypQ2N2YYFRSrR27YnWPnUK/e9eIBQtT8og8LCke7TJzXa
VEVsD4btUtfdyClDXC1flRB3HimQhMdJN1ysA60kQgY4fEIVMFkqJ1UxD9ziFJy9
3YHGsJlvS1hhraRATLEYil8ovivTeEtAV5Z1IcixL9bIXros4vXrLZowWlw5dzJB
znWp3h4V7b5ny2kGmTWcBAG7bDOIQBEwIKFCyrgvbKAh9RVxE+g7VeXeHSkTleP9
oO+Evv8kiRHGHdPcYo2RUGd5WxDtypfFOmhbt4CofWadIdhEbsXxEsHfcf0q9kUR
V7+6lrYvgOM2O9adcD0mKfftrkrv7+L0okwDKoBoxi12uAxkDMVjUn1upPHoipzI
`protect END_PROTECTED
