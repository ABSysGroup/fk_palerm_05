`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ev9lFWlCI9vVlTBckKN0mLO1ZoWygcr5l9NVsljOmbVifrAawM8Pmm9vYJTQSs24
KvCTSRgnP6nMPuna+23JlbAbvCHn5vGU3NYip55M81S9IEEw4KAfDXMSkCxojoYz
QZU8Pq+Ianwi7G0CXJQq9FnPZgpXXJHOnEgQj9rz6fMVEWEL/rj8bISIRD+nGjlr
lACtTz1ukA2QshCvnD3ZOGxoMg7EfK3Yf7bSkeqmIDxxLhLHsgDpTcAKshObR1+3
aK5Y2r2/+u00hSrs9i2Hq5NCMMOVW/bGtuupGKmau3WOv5y0Yu6XX3jvlR5Qu37u
WDvpIgNxaHhjQ1UMtfrwTXiO8iX3nFU9SQNU9an3v/VnseA1sXi+JvbM9Vqu1/Wi
RHABytupo+/T+NP4ihVvy3Fdjl+GAuzCBLa2WE6hy0Ar4Kkx9+d34da2JRuupuSB
ruNZN5fCtfr83iSsXI128F2KnZ7F/QzhXHV1KpWNGb46IS8vj89kEKhra6CGN7VG
FgSXy7HDmEZ2Uk1gFobEbEgdNGWZQqwr+rhnX+8k2pebZfcUu8XOKy0+vH/nrFjL
XTXUqSdSNXfjhSx5b3YGd1PNQrwyoUjmmGVlrfoH2i5jYm/osn6QIQE6ViDGKrsA
TVQMgk0NajzIJhlWVzVAv5uu0rcwKwyMhcpYPPFOquHKl5vACU5bDawt+qX4p+Ph
PiKq8s8BOtdNjSWALussIinKjuVbxUzSA4bv8d2ywNMUJsBPd0IBeGUMfC2pzGJD
bZnzG0vApVcbL1w1IyXOYlcoGtzVsVIocrnmeBMmr02gTKy06zDRqRax2z/OXHsl
/xj/qF/DigbFiEVhL2ACyNMuJM887LQ8GVDktUX7IZsQxop5bL+G0OmWaU8bYrTy
WL726BP00Fq3B2qFCOUiVA==
`protect END_PROTECTED
