`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xnST6UFbxS8xo73dqDR1v05R/4A1IN5zsql3rUkUIGs8BcleTGM5I83OlFXcSavt
y6nj3Cdz0zs1My3nxfbT+m6MglVotPehCuCnA2u7rKvsU1sN6LJwpLH04TYElN0X
tsJMu0ZZmCSbKmkHBbEnYf2/mVa4FU8Hf2qmnLc5z1n8uJbuQr2A+2H2ONOAnb69
CmY7SaDHHf7cgY5zjSW9DULJbml/XxgFPHj/4IkkxvhZtrUOyHE9SVlgyvnd1hrY
Bhd2QMtOKbqjKVRmXi7MKxHJ1WaEDEb1sZcqIoyYkH5kqz43T9WVww52wDLEkCDT
tdB5yMFRTTZz7YTOVVOYUbdVTjk+o1KaXIRNfPE7OnIzxvziz9aTV9T0AmK29gdO
22dDTigGHb1SP/uL+KACO0VD4o50vJAo+7OEw9nsdpZJqpN4lfeuKjp1c6UeMbE6
xigUiqgBOVVRiFjrn7XRlA==
`protect END_PROTECTED
