`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zb9R5Ho3d4cxRuvm5GuHduD8kAO7YeeOEDceUNePe2ritw/V+2hOfTrlU3QDTqlZ
CksXTFk9n7wSeuF5y4YJi7xmK4n3xggyC9Ay7tw8tRwOqF+c2uxmJtiILLCrnLFE
ewB2P2vEXgKLW9r0rikbhj0/CzuVX+CgBo04ZrV8yYu85Ms0YvkvX7rKSSFzt/c9
kV8bULwaj3B5Y2YzyjcIzQEC2iSwMJYyTzmU8F5ELC1Fsk+LsUs9buBg+AwzqWby
GmeUVq5tlmNjcoIXAj1mejhPEuQdemSMCk3ADa52qWLCQMXC+/u9U9xAk0EhF84G
FnzIapLMqOX2RnjdeotQrnKbmkdz4XicTFQWZmBZIDNnSUq2eogZpeaun6MZqtad
NJeiQMpcv5rcMUnVZeOAtZqmKryVdB6IKfFDPidQ6W+2RJGSg98QXvrzdVouFoJ8
arAAtMP6cYcqd92Gb0NnNNDEuFaOdAbUaDFoe/Js1JaXClvpqbuq5/kCMH2IhTyW
rLP/kYMQu0XPh8YHy9pnVRB2iwtUHAk+AZlB+FTlfttxCvgEsrNZ+6fw6ZrRa8xq
Tt4oebZZvZUrvyT0ZExhcMmt0a78akEYLIhuy/LlqMvSBienHt98NRZ6LL7U24CU
pKof/tmnio4UaK4lVnc1KwlzIDCn8gaeMErtxJtk8Rvid+kT3+zW5zDFV7CJ2G3/
JtWYyWQEOSinDxHrI+kn5YFjTuystnFRfSY1NRzqcIrpLNAkNv0GQfd+kwlmJDuP
Bxd5MhFTYPqBgglw0oBjsDkPKEx5rOLUipP5n67+0lk5X9Qj+ihaj5rgFXXeWcrj
qrckZOv20WOk2HAghpirymBvirxUdZHrDbTozQK+FPijrBNyGT/bwid5VUcoPsPG
GS3x4kKVS/kLxhj8n+RQKi+0jzfu32jcsXwr0cu5lkNqvWZMFSxajlcht9+8eEMP
XreV4hR5pYojP8uQ7joIYHSa6sroMVYcYlsgoEqO4CpDkqSNirHJiGSa3bWQNFbJ
qMXyLIpQtr0sa1lvjUi7rwvjepN+kPGX9s6CY0okpfgdHLoEIxTe37+DX9q2HfVN
qEkzobpxZy8ZuWPSMY1oXohUK4BgrsU91awIYzPbwGXHMwDy1APH5GfAyTXBjkEH
jKzz167k27Hv1lalw0ZNHXhPAC5oXG2thZXu+sYEEzHPRDejrsBMLPNmse2Zu9SY
DIxL53aM8bdyLX73dQNgOXet0pyhz5+ga2StS3bZIVdgZdxHJ1VRwimgy5yej43V
qhhdOX7wQZ+HFD68N7TVR7C+j1TQlgbOU+BIdot5XaJ6D8Qg+gTj2+Z8xUpUb1Mx
cO588zJQzfkF3s6oKVnS0usNG7/obDGCVLiLISP7eNCsfUhT2MqxQ9+ZP20qClgJ
87kyvEtqYUErcP5SqTNBQMP3gyFYzngJRRj4hTK4u93X7GiGK9W+ZHUM9gsw2xid
N0udbSCN9qTdgAC0AWqiujBatfpkyuZCkzAGxy4IKLfyqIvmU9dRbU8AZR0Y7GgU
8PJor6bUqSjUbPnejGLEQUwDAuElvYQxJd1Ou9cPGYDD8eUwZV4RpOcpXRdRLjgj
lk9gyT6iDO8/zvLUtd5wtgyur6CKvo5Zn5SAD+aOcC+w7RHyZyWknfg+/Jv2u5nu
uWPVSV+3Zw7aegdNV9TfGfR643LjCTHxyzi6+oiog6s8p570PuDhPv0mdniIa8fQ
U4HJkgDX2ZakwjG0kxkrCSYSYKFo4MguyCHHAJPG/wta6KUspfG9EGm5jCJGEBOB
v+xK8BRXb7wN9uY014F8ss6veNOJkJ+8ZssTrS/BNXaU0QankngBjiVvTAejFjF9
sG4/QiKkG8mE1lbgRhAhmX5OGh9xN5k2t8JB7q9uvfAHTF531bnW5yGykZvVkVOH
nJ7A8RLxxY/6iABF8PMCEyTZOg+ab6hyV2eDe482QGgp8UsptPJShTXVDInCdkmn
BlO5SQwhjQcpJ3FAtMKxq/HRy922P+nnORwNJB4d2LgFLPaxPNNHS3WJCvtxM7od
Znc7OUDuskle5Y5UTnKolgLaPQLsleDtWGdZZX7O0vFbwq+H5bjur8br2BdbIAj2
P32A4q/bTsPvJnAwqfk2Nf9755WgI3cqGxYXCGecQ6ax5tBRkk+0vGgQ5q2zcTjy
p6vnliQ2eTB/50pgcRsYdQp9zRs7GKzbTlO4ExB189nGhLQD7KmZB0B8YYbOH0pe
bCqTCefMqUMl1PaydJ6253DjqTDFDLdxHm3gmh+0wlPUM16dAsOuUCagGQjUaHnd
9LlZvg0SIPJjQJdnYY8lKS26qYcyo4EZAg1WkujSIyLyvM7dSxKe4t93X92r/Eax
CDowGhn+vB3jWmlpW2XlXe6LiLTL8VvgKp1mBeaWI4kffWO1ugrmeSPv5vPctEvo
nZju7kX1N80rmM9PdAonhDYzYOAasknlEbMxp6fweGlTBa033ZGJT0JF/W7kfJY6
VOldpY+m4AxHhqIuOGolVTb5bpwhHL1EyvBPRoPf+HmaDiHensBDNuHaMKtm//mr
Dt1rqahSfMs46kUtUKajWvlx/lGjHf+v86ShhyQ+xjkjORGF7jZg1MhWVEEsP9jC
3usWfmypiP2W0D/q6HGid2QV3yhwQKvdEQnADotG3KuRWvOSVDpr/DmKq42tZdo7
Be66atwLaKV1vCrbSWJf0h9op5hivM8UOK4wZPJVhZFuMSt4AwfGAsCoG3ip8WAQ
p+8DOPUCq2e4ChwK3fy4IlS70IsgAsMtW2DItoKpS+D3Vl/ho7FIpidqPycoVWp7
qsxD5K33FBpjUJfacG/AnxYXFO+NRXNvT34oYT6sg48fQT65IcIZX/GamCVWtU1t
vPqZVmwTYJ5xndPWn7/bsQwj7uISGtSpJR8lRiA5cRrLqjEUobI1afbTnPPI6RXU
qW9Lej9oPP4I8mpJqHQucfHWsKBGs00NXe3aoeD5fGoHB2L8WwjO5JFkiwjgCaNx
cI+IWj8vHISxgotJ+WqPa9lbyhfVn8ooPy0xWgEVfPXo7VpDISXJDHM0ygi3F2aR
SYf1sZZXrkTXFigDVgUFlKKYE9kXRUEcHlloaAtLrTjBb1C5VGI0OzkLOoEQONyc
xTeYZ81TSuaSQFrxXzhjJTyyA9QpxQabOVv9UYMa3Db2QseQw2vYFIi2FD/1XwG7
XZ3K5HHvJljzCqpKUAur/AaUfW+C2OsbP9w5wezf4dScrIWyIwXi2UOaD2z6QVli
oKmyxJQKE+fshris3JbYKM5zurPizmwMY23knsnzHLAyJ2uu8iv6Sn2TYdjTgIWJ
TEZkl3f7Lfhqb9dSlN2sVUYXgYUT088nRnOHYjj/R8TO9yIOjmMi4solkUkReEOx
q2KJUvbUTO+7cY6Jy4lDF0hlg/0rrNhc1+r/obBmRND1BscKRRgOYGLPslSIQ2nR
xGlSrBNesdnoZDO9TjP/bOIn1MDYuVn9RSQt8Av28XC74DkWjLOYQ+0ZCvOl0S1k
F7y5nmgGqnSKsEcOO9ieNG7PmBvO8OrVh2pD0EOAmaNfMOARmP23fPHUx5a+vH27
RESZOSb6ZvQLIz+9l8r+DnDZXXEF+iRl+aK6FH1Y5cjCBHpCATwUL/on+5Iz7nkE
7Ibf/wabd9unu+U+bHz6IfWKxiHA3mMaVXOP90SvhOiC0yBESoaP6mE2Wb2s9qUu
qIDrk/WqZxtOLplsR5gfp3RtuNRerUoPzQpEonW31Z7R3JnNnJFoUkqnjBSBaPch
dRpW2SudeFptABfBqT7cZX+OVN4r+lM+QaWJSvmevjkNQ9+19c7E7roKY7lC3YHJ
KZPS0AOmU0Yu2dzYtdAiDSeT+WB/21/XMopzHMi+KTV2n6KzZAJ0PpDweF+ll7e9
X+Nd0++mROjeYd1CPmBPusXQFh8+EEWhT2hkHPIbWcqKRPKLu/Mbzx0MarzDOo6P
e76qwSVMLbkVY5eHM/MONWphycrC8ZVA8pz9oKG00357hH2n9BtNyVpnOh0gzyDN
pFKYDnHuNmYObMUNz50QuEIo5VX24N80ErPADRdDIb6kOWLpBm8JRrhX70vtvch+
VCUtEX1vuY9DKL9BlC7VWLACNNnvDvNEJjNgORRMoPWn3lQLD913+BPzNZDXYr/o
WUQmfFXshi9maUYhycLsovuu54t0aQwtlLfa0JslbnAu8QcbmEbWn5FHHWwGMjxt
5tYDRPfvr2fcXZlOJ4hCTagIZUPJ+0OO93GMgM9AiFNrFY36RFwy1xEN4Vc1bBND
xcn45pExzr7e5QMgi0Kl4sxM0k/vYfAiV3Fi4E22pG2kcRoggP7KnMjP0rBV+cYe
DaTbTqpDb68duc17ksNUgzqD6z7Qszu+HDdaVBcQ+S7NpaDwfAJICmdyJfiZGA7g
fH7WzD5Em8HPBiWXFxM0siYn+ahm/+9y3UH7Jonhz0+wFAARfLjGnu815d9ASb/3
A/my2ygWwQ9ywWbk253I8p/eGDSuVDvq5kCmncdKep8wF3aF1C36bH77qEj9ieuI
ZdcGlmlDpd/nYCHgHJX5K60FhCy2acPul9ztxx7RQcxJzP4sdsdwoQYD3N6u6p6L
1u+O6acyc8E3ehCmBmTcCQgfxG369CZNJOTOaDrRS1dHnI+EpXiGPQdd2x9WlCHg
p81RxPdKO8aHN66WwrRRzz6WTfGY7wJwwmpJkxp5rcIzboGHIsifkOwYFNFP0ptM
LlpkSvM56v+rMA5v40fQDLQ6pMfhPxxtnVsQyHwaGuBrPeBfbXNeqzZKQP2YQB7+
043pajUN/MheeU+q3aUFKSHfsuk+kYOAE89bmavI+FWQ8zVLVHMxUXB5k12CcsKZ
/TcdLSvRttYgY/qJjc8/9ZDrN3dAL09byg5Iikh08lc=
`protect END_PROTECTED
