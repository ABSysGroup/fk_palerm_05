`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kBKlrhK2/IicXuytk5/nR+VOOMKagR11jStCk5YqTBixnTPfqSw4D/jBk01OJee6
hc85SPgR+W9JTyTCVlYF6xf7J0oil+vjU4V+kIrd+XoS0zLwk156ufSiefqH4Sev
kwURoedICCM9QsTKhWPS3/gals+quW4nL3xQX5YfTknoBO1ubNdqOLTY2O5vFuPB
LuVbAvHY624avYRjYaATVa2up2LWx2I0rPy/jqqA+VL3nKqvsoVvCe2ntlUh2coV
Th+TAG99RFDGUcMObdLg3wsh0e0LIEtJtLd8nm9GCat9X+aQVQZy0chvgTTWRAGO
dTwrlKioKixF6ESHXmGeJoSrnWylayAWuMCMzV4tiaocAGNY7UlUL/lenLhRYpdi
cGOvZGC21quvpbxqvh4o80/+1Lk2sy1BqwNt3hGN4fGbGR8TN4+5e+lUsdbAZNjY
cuM7ji7+QEUmDxCrwcpRs0Iq3Q4+M9nShEmNe4ayaZPdbG5bDJdz8sFdxyMClfZg
+13SCPTNhhfMVlKZ8zbYqPiu4CuDctW1sx/XsadcHBCdx286VonZRGkCKNEHujBq
sqkzglzqHD+8EcLk473mKhPWnRiwrx7MyZBw9bXhBAQ=
`protect END_PROTECTED
