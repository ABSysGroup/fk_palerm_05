`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jzjFpWT0rb+ZBlgnr1JqfPApfnWH0IvJr73POcQ48PVjNPXpDu4xwLlTJni+CDWc
fzyOca5XusytlFGvvK4Xw5/BzV0ny4WRD9oQwwTs2FYjuYOfYBksQmFqRaCUJgq1
AIUd7Hpp/DvYt32/6d/pGUgLf3bNtwY4BiCsS0fJ/etLHRSRztuqjYmdkRbD3Ny7
ZSopjkpDdjmoex4mP/nY1ZAz265ouXesbM2cOJuWP18ePE/yhugoYex5SwtJu8SL
cOiiB5VxAmoYPd1hZQ3sZd4P306ggn34NWRYwbGFmUmhjC60HgSk79rRmdoUPSI7
Dzl19kftObP3IAKHZghx4dH2KuOh+htGsBEoLh6nrQqhuJkChfD+y2BFiB7N4Res
Ve/DPf4Obr+h5swaIihCB0umysXZHyVaCor/VtJ4T/L5fDWv8yloFc9h1Y60mBl6
`protect END_PROTECTED
