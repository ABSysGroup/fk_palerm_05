`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p/xMjyhsf5JKTaXY9d5mvVjtyvdNo06X/BJ8BPZ5DEiU9x5e1nn2k+YgnC1veEgh
y4lSo/9F52jhHZT2ZQYTdqLCilZJXVTg1Q9Lzoc+F5Ep5vsy6E3/z4/HtcYBqoP8
2Y6qBEmLq1XTj4i+VUEf+ib8yt9hcQCWJnI6qLnCfX9Nd+OI+ZMgiUsTq17HmbOi
eXB5yJsPsZOJhqXYJiVPZG6GNgXCtR4aw13yBwM6M2V+fu3EY0qbT4JA6QWcHRoA
uBvjXmUg9B239fu52/WuWBtfHpNjJHJxVbX8tJCBwipMAKo3iAgd1vXtSGn+b6Ap
TTeo4xfdYswlFt0anHNirupd+0xMNMOmbaWlDcmXImqdZvBRpD5gozXGB5/rn+ng
ITBIWhViDq9Wg9DgTKDktR9E4uwUcMZpNDGgr78blXgTpe3QlNzzpVa8XV6V7/Oi
F/Db6h3BSUVYmSiNO8WSPcvZUldvfjGr2SOscYYvLepKzKov836yOjy7Ij3ZyVhk
`protect END_PROTECTED
