`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tzNimt3nUsJjlF/YQny5ij+vcP7d3wbUIKYn/jZQqBVl0lHAOU/9Y9WaI8kgti56
YtjiIKUv9JAnIPAmEKeY0D6ehJPT8JTcQjLu472YB9m6uyAUaNmtj5spIQu4kgAo
Ogq2x/UtQv9qDVizLT/jbEaWiWUaJa+GsPLvJOFaizxCt0Tm953LTG46MnrpAyhS
73TdIjHz2RVMKW8eM6TJLwXXXbVUKBIqQmr/PGdRd9CnCjmm/UjzeIQAzDCwgBRG
tMS0BuJ1NlBVw2Y0Mg4sPZqh1D3mZ1lbms972DpmgW0XBi+ivvTSC0huszT0hbAh
xWkWVvUMxd27PRMl43Bk14hxEQM11oWG/nJzpZhylCiNDTT+rRb79mb/blNsR8xL
P/yY6r/qgNXVZwMNsROqiP8mf7qIKef2LglTIPPMPIhGzemXwFl3sgjIHAsY18wo
cEQph7LBrvESazelKuyJg2uJrjVVIA+oHlUjRdN4Lbw=
`protect END_PROTECTED
