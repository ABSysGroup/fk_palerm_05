`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y1kG+HQz23htCm3ZkkZ6ygU7sUhhYt3ZzM67XDHNkZPi8jT4CFcTdTSHpT5kUkcS
ny1y3s3lo7eS7zmJDYVNRnvNpD8lhXXEDQV35PeRYXVEbwjKH5H6ZIH/ZSDcGOiF
VgJULWH+si7euJdBOlnz2D0uTEsol9eNOFAP5Gv3y2oEFsEV2QiU6NZjfNUXiRM5
JXDJQV+xdhulWQ+xM8Qz2E5fyG27YNNDR+looeOHppFJFLPQoc44etd8cTMsIVsX
6MI0Wvp9FPjqISdJxHFnkOJkG5DC6W0SSt7uKJz32hdMjJIYMNKlV9K9CUeTsEwK
34Q0GnZHW2lAezy4jpvLXg==
`protect END_PROTECTED
