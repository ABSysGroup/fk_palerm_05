`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mr8xRrI68OjEAdW4HJbhQtDHgyQQjRQugoy+rv29gfthMcZ6cFovFSKH69n+nAQo
/YiyiK7Be+aFY3DAY9ArYBkiaH52soLSduNQrWIOXNJFrtwLBpfU4Rxi+0TLbGje
r7Ubg29EOpGTcJltYcGZu27p3SU+JryIL+B6KTFWgkubhkEeR2BlXbYOx3Zg1n5w
F0KbQk4Bv9fjuuxpYadTzxgK3FmdA5MvIs1gCp3h5/edBT44zIHPwNP3wNd3qA2O
1W8nJEgxKYHEYsy2I07HjrEYtmMPdr8/7D2XdjKGjlFAp0qq3rnxooOOLhuAK+Sw
wEKLwMbkjNJyMDKy8/qMyv6UYvlhbPAFFuWHWyT1gCXsYM5NtFCXuNxxR/VvrqXi
`protect END_PROTECTED
