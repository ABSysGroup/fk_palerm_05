`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EHWe3qvsxf2jkraUWtVTYbrDCgCR4nw4eig44pbsrFHCbYyi3WJmAOkQe2KG0lky
FZ6wwfqkFiQGX9YdCLGGSXFSW6QCqQws9+n5Hmad2tA8XXagV3cASj2Z7UUsCdgW
tMUEYMj3rxg/7E26anFOdQgejxsdHB4rfxHnFybF3itJHyO+4Mu/oav8jNqNs5r0
2g3+SF2v48nVvYnTtupP69tbUaaQOrxREAHOAkvlo9Jw1W/6zhBS+TeC2EzsAKfD
XDVZ1rc9Z5mYYbN73fz8bZOJGFAIAq+WI91sMcx4wdXk1G1p3aKmTGBwd2DIPKqd
wmrxfcTxkrF2eEd9dzZiFy8qKBzDlcqnt6iPnhwPx/mPB1LIFQJvp5h8sBHgNtf8
rt0b3sW4Ls0oYLvz2Z4mXe//QklTz92KkzfSeb6t+jzEsn8q0SZ/mxbRmvXPJn8u
6HtT0kvEbAmO9GcyVl0VrlMqViMsI6fKCMgy3z06X92MehZRxcsMbZVIDR2v1oNG
WwA/uN8O5m8kGoDbPXuprSA/2K2byvPlsZlP4FKAPibFDZRU2mQ1ZFAnUgMPgpXN
pLQUhU5rS+Sm5eK2K5ik5p76TePu72EqVBAvaWz3SrA8yYWJ2tYqeriSkKXuiZqJ
RH8nQ3N2sWIcjQdOBS2L8EFX5J3qGJa7ZODdPvEctkXlzWDz5CiDvkt5kX89TVwR
lYlzBNzZqOXNFBzfLOR+K5rUmP2yi4yVCQ7CQVr3jZn4bfIEopjSKwY093ajOFvh
wwwGlXmvAEESZIeOviHql3lbv4BX4Qt7VabXTAJrFKySllRhgDsRn1gmAI5j68Rz
v6/vdIqMexXaxr6AK5OE7WQQwkwQGIBy6z3nihcsL0tQBOBcZAH8wlQzP3Jv9wqW
WzfWtZU2QFK32OmbOc1I3DpoR2wW8m0K4eC000N6BqpGvhDItqXdL2unZbHSlNRS
oOliXQoiQf81vZUZvBQIIg2HoSlHfyhnllEEIYRw7AbMH+6s85ZzeytuQPsVTMD+
tAFfx0qpLvrXmG7SRwY6LTr2p8eB2SS970TJUPTBHEUpCsROvT4VMDlHO3esyhYo
qraUfQGlTFVbwTtN41yqYtRnWJGf/cQZ4MSM8mopkp9CuvmYCzPc4fw5JkRaNGwF
n1JcZiIajs1NOouUYGh534NAGjnKllLzzm8v92SoLE8yEiZhU6OKdF/3ixjV4nkD
wX1IbQekMr2+ptvdUMES0yLhYAC13DJsUNnimvneQ2pmLysh1xfbMEqrKs3jxb/b
+9WAOTjZ/KBawpYLjfItnBbGZ3mBzZu0N1a/TaBs93iiik7luyTVZIgfsS/kovLp
bk3bZb1x5QZ423w89Dphqw==
`protect END_PROTECTED
