`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ClkfMveg9GnifNI8gNWzX3/5XMgYkTaCcZ37UBBO3HWxfdkWRokd7xm60XLCKiw3
KTt8l2nyTg1imm8LtN6KshmeeAtMn2OFutHHKSPjsxzR4lM/xn56H1MthPYG10uA
cegYOUimv4tPU992yxMKN3ctJsXig0QFQfcZbo/YU8YPnchPnN8RXX6qxEu+LazP
KDrtv3vfgJ78hXxPkGZ+w1fUP5ioJef5MQsM7cYValwSW16Avc+b5kET5SvE3Hoc
Q1vWJstby9vH3BZ0nV149E5/H1FZooxwUcQ0HADUnOB6sJb4zqC44TN9zHopAhgS
udiJiH16RJ69Z3KswpF5wBiB/oq4saEKh65ZBoViUBzxuVd5VMdGjCtOFaGblxYG
GoXrzyiPea/IN9W3NVblCQD+Yzc6htShGFJ5UzMbXDE=
`protect END_PROTECTED
