`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
clM0o+pFDDfWOvANCFEyFy0Gqv1YKeg69RTetBAToiexR6j7deHmcYUfdXMWok9L
a+eNubqKSMVvHOjMHA+DjtvUTMSRbEgeRJhKTkzzwMMIJVBMfC29qUGVHE3yDjbg
v2bZO2Uo2n3dCUDn16jRvWX0ecAhWIJAKLGiy/QGh9E3XKGC8vTA+wtlpyHF/PQ9
/RHxmBTOfDUqz7sOMO0oabGmX+Dji6qu620a9a13OsBdBQdk8Q25HykvWQkaILAf
Ea58+4DgZiSm51c5lt5l/SLOrbMI9GyqsL1iD82eE0rHCh87Syr0LyDCWRP/NLcc
ah5pJN4FqYYXeQ9sZAUgbuKE0RLErACASaJpG4CuXMm1XjaIomV749ASxXJ/7CUB
en+neAy5CxDbpzhCVYVUfKc5KwPjaaAEDw22iX94j36QZCCCPMNJfjbvsYsEC9Xh
R7sqsfIUlEBLV5VjQlOETrTZ/T5Qmv/82mJrOQyaamewxHIxqjdPLTxb+fXxSeqQ
ZqExK3yo1QRgMjvrUWoYew==
`protect END_PROTECTED
