`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yuyB+wHpwXsXg1wK6p3EBqjsRnzJM6lRQQTUJtbtNsYLyAKGGqTY7c27A1c4MghM
jjOmYY2+rnGW3JJWeXdwO7cB21fPoLWtgTr0cExhF5BcVYJGes4Ms54qXlLelPqX
6KqyvbIZ3rKxNWC1idfl9MdE6fNGhxO2Tft/RvD0tE6U3nBFyQmHv9/NkY2YyKWN
y5PPwLOTkmQqJQYaqznbmYW3jsarCUSwTo3/gCJ0xkyCRVEB4yQWj6kcx4KVZO6m
Ldg9pszmIyCYWeI1aym9ArhzdDgV93MmMFk8AbTqiI6J3UVNbg9m8FmBt48URZrQ
YEDQAjB6e9KYysZBW86SBCgpmHBnMXwv8gWMFpSmqtes/eBajksAd2jRAslZNyJ7
eRSDmn49NAKg5xEv7J3m58fzCTVYkNQCcNf0+W4opcoXG1Ch8j/yxj8FbNMShv1Z
ZCyhgnMlQB9CpAB90n1Yw2Z4Ql+VYN5UH+ZGxvCGMjIuInhtmmAHrMHA1H4uJVFd
9eXTwV639SqHVJRaWVD0vMISNPvUhpOw/LFenFBgp7eFViSB+ZcokIE2KqsE7ItC
Awa6o7pIdZd59Qhts5mgKna67acbRfg2mD5CMOVi0JRJOa5vjpmX5uJgXc6KqvcV
WE3RhiE3l7ho3GcVvv7PucN/V6g69Zu+w/YUjVDgQ30dBMf7+ICBxIWRoFA/sgUw
0fNIkXvWRDcKd/KWvlBdoGW2SN3NeFc+uOBBxR1s4CF5OMQTh6K4XywBDNjwfu7d
giWk3ieVeromR3dJ/xaC9ps2dQCzMo5f89zCoCeTLkAgH6xhLgH/0l0FvTbytpcE
TjueHTjYRjuCwwZClRi+c/RZNCErbgWIMzXODcnI1HJ8l+Bo9uiCtKFCcLbmUL/G
+hxHUpnxVjVZvHvdTWRsm/omE2Z3o42Yvho13/GdppyTgPck+yXeLoNuu3zaZ1Um
hkkwLBY3bazaYlDBx7MMP+DjbYVoBwKDfZlPdfWHE/odj0eWsjrHOsCohEana+19
ZfwsmIOfBI9/RnHc0Uq/wxJJWyVnG3i8fl25DuZ1zm7sXy5aW2cEev2+Jc7sJszi
zvGNa7cGGrJflcgeU/3JhXLd3NoTYgqwKItRQhyryFXBXk/mTWQPygQHRGrah8PP
3g8mePLHcpEONJg3q8iVAwAyu8XduPSQh7I+5EJOJEgK2TSu5rOvYeRLWdueIOiu
tnz8Uhwhaf/Q/t/VtzZUSFFGlaECgw8/qPjCTOlSIINfADkOF3FLYsLbaISQTMym
emNIdnPDX71jWmmNItw5dxxuenKzAcsYMZ0UtRhabzE1Kv06AUTgWsvNHWnu+LWS
u3dtx8UYZ5JJIhtmO93VFSRGmCk38uoZl68MQHKfhQbFglBknIW9nhloz5vbISoD
6KF+lLS/yl967B8EeRfGetsn1AWKkFTvNAI+3bE76cPzlYHKlM92bKWo0SOZFnxR
6q8ikySMtcJuEqzTxomEK6qHFsC7n8PBm0aJBFtTYy6u8Y5yh2mOd/eBuAGrBwGe
t0MBeistPZv+Zb6sy0Jk+eVUeQgiK/yRRNToYE0jcrqw1RrcJjF91BLd3dlrgH+I
KyuDHmVIyG+TpicqqGgyDU/EKNZsb2qVWB/Mve/TjWEwUJDW+aU3yujatWynhMs5
/9Ge+a6Z0ZdK9wIz8IxihQE1nHjdVtqX6NV7mv+IEol9Xrk4xDPtpwdYtlMk+7Uu
CGhMIj6LzKj879fbE30x9w==
`protect END_PROTECTED
