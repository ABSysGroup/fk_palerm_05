`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MTfxaHoXJT8Qhb7QAUn176HuoCNsD+hJEKH+MmnKUsk098Jg1LiDcrsvvrd/OEBZ
bGGjIYAf/jZRDVhJV2e/Tm4rjjqaZ6tkS0WHfwAO4bAGptJKjSJMfasOhb2b5I4O
TjCu2TXTy7XkN57TufrhjLW6vE8TSeFJMLJbnmXgaGFAUxu9qCMjcOPw/BCmQz82
DlZ7wNhdugV593taxn6bFTcjYG0NWBolCyfSyJpKVsKjFQxSxno10HdnRFbj6pCj
D2YCz4D47AGfGwkJS6z57XrYUTzn7u9iEP0OPjoZgWME9Kz53aY8CCjP4dUE+qo7
RY2TxWsr7HuvFwDqYxFfByJCuntbgJMVmDZQ01wwVgWt2slSb83mTSwAoku1Ayoa
Bdd+haO9DGr48PcSR/ETH45Pi4MyqRon4FbJqHjYOe79XFmBUPy5j7sEM3W2sQV2
COLnxRQ1RNBt9kJm73vIjVC1Zazj23SphSLhFqdSK5yzsbql3yxpWCumOTA1CcmG
CSUrwVtMT6S4IEAGprGMjnfpSo8/oyjxwzHDyPtqWMZhVspSnh1yu6GUzmMXca1w
pxcixQGFTdxjY/5i1y0g6uovueoXpZ1Yep0sdHPXTEDzQXPsm5NvclU4C2B3ENkf
Af5nwOMiFjRkIkrhmYrwA130kyNZDuZ56h2LoHu08VMRZizWa1TKEu9Aha1e2c9A
wjN0H8Kt+qkuYqb+RuYvmmVV1M2TUy2VX5MnlTLgn3euvv69aLskhxhatUGA5l78
0uoXDHlZCenvyZAju2Kwz89PZEDPwyIN2hv7srWTtmgbLuNYfKoTb6L6cfuY95RT
qJUBS72vV7H4mNwt6Qwv/Q/1caqCDghp1dZ4f5U36ebSSlJrFneKr/XpLRjoPGnq
0SrJKnbMBnNpLS8j0nLQbmWxdExfQfLEiVggx4NiMcd7xkcV3BTDthzevkbWkLAv
BFwbUkfCLzCev0IQPzgBwxMQqUHbizHW7KDW6tjug2D1yYSIg89s4h3sv9m9X4Nl
bwh7S9ABPJ8Cl8uuqKjovQ==
`protect END_PROTECTED
