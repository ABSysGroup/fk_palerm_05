`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6+rUGVu/HXe5rn6cP61oE7j7z1gCO4Eq4q07oLaOEabwGefKT3SJ+SuM0uI0ky8e
ZNsEwkAywX1wpZxzOasc3xv5cNstzfvuq/kzLbemSfa43w4ZFawcqW7RSHdeHT0t
IJNoZv6ARDKRlWJxymICKa8ywHG1ngBB0V+kXIM25LOsHzF+QwKjXhREcZQbCHLq
aljvR7m5pdMxgbdR47vb+LCbQQ8I8eg069/VAPFuhqMh5SHo15eM5QsTYVTgDtAT
RTcsQeuFd1+58+gvfnIriumLO8FzjwVJvfu+3erwxaYXZgCPvRgmOR0Lm8cDa7p/
UQxbwasWPvmHKGHWuScb9I/dkSMBeeJE2opf2AlUSb3uguTnRMxthRr8ktoLu9Gx
ZtbmSAe7Cnj1La/X9yqNN1Z3939/9Lsfz5qKoW4o+NJ9rEf9llTlleRMq/+inuaE
bv6G19iGi11d55hVNMyFir0f16JjVnV2DpusoayTszayLU9XvbliOoVMRmEp5Fg6
oCbULqTdgAtdfdGTHx+rysNTygHKnB8lvGHizuq696QvkPKOIBrkbasWNRQDtSPq
MDQ6n3QToc/ITVUBoDOGff9nBEFPxV4qVDknN/Z+dyQQrSHU5bmQzpNrhIYutMwl
wSqiwhPWdlm8JPhLAuTRKJNAEJUehtbNs54cqntgxxiXdBPtRVdbJqf4sVUOG9PD
Bpw41/OP44Bx2zCeL4aQmJ4LD6vDJW6yC3RsTClXM7ooHlevLsL7aeILcMdGx7NP
jsvbA+49YvU70rA9CUWzNhDr/Kqjle9hs1ENuK3AKTejDTKKXpubng/Odk7tl3+g
k4T1QXv+K1XScqXG29SS0++LDTxrz4i6qGy6FdwnjWFUo4P7PiO/vIuPmlCEwIid
0AdWZi6gDZESYd7RDhpEAMMOAgvQ72aVQiHi7y9TDwQjaiwz4RkFqZ35cChbFGGc
`protect END_PROTECTED
