`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QYofPl6bUpgSX4kXS1ys3ALnIMwnga/NaqIREW797GLm7a9BrKUyQzoCPgh9tjBH
nHWGeehQeRik00HQYZX/lJhgE8H+kloUNO1U2zoe85jaGKrmQgrUiSclDzBHSc04
WpaguSd9Z6ibaip+ZN65Dog0e4YqKCQkD5pT7uyrJnY5hFkwBuZ53RBcbzK6vZ2w
npIyYc5cWJf2WiQsJjcMBuvNDTzdsjyj2KScfj1EuOGG4P8g6x0rfchgT1cU64Ma
dNNd+2celPDYQgAcU7wq7rHbH8H9HBo94wkBhBKKpqwkf1Ty8VacHy/TOz16Rxpi
rKuA1cINVvsq9R6snz9Q1K+b0B8aw+8W83UYtBmXA0ECdl8JGAei0ZWgQhMR4uB1
oGUbfG1L8d0UO3NPvp9s/QF5lsks3lY06Btzj+dtLuyBzX90Z2KdVexlBQEd5AWb
oBEUXR0ZsYbidVXwF2JpiGOiEG0RjXl2WcXXUSJdt0jbT9BSWDjW6Ijp8JM9aOsj
QUW/d6Fz7WClxYHYbOLZvU0GPLJyMB67WjJVJiUlg69JxLOj5hYgEDhS8QoKXIj3
W93Ju0+GdyerRNBvBvHvgDNToWwvSuB9arxh0hTaNIdAzTILKvyyO8Sn5tG2ehil
PRUhs3l6SL0HdXpKirLrlk87LuGnQ512W50EAWg5uT7Z/UQzZmKaGSXqP6HNZoc5
veOlk4MbzzfCGGYBrn4qpYH4nZGWhtY4LPjEhqfnvq4Nwh8ikaz6LCmAo/mfeoO5
smxOUHs7/lbeiV+mzr4hoP4ocm5HeIliwN2tPlGdLayenlldi6TLApHxEl5uNDl/
PhHGV5ZzCT+9tAq+s0ljvlDuwmXq3Z+wG1BKX/Jol3cT1J2m0j88cz9qGIP5wLsP
YPd18k2kLIRtdqg196hBa967nL5UNhWOb1IrYbRmZGsEuJTSrvJiTxwC8KY85OBL
LjfY23qZ//CCwwR2ABIWf5mo4tSBrrDXs5urCYLD7+CEK9ub3uPdd3fl2sEwYVrg
b1Y6RPlV8GwXpx/YW6QoHjBEIko85oU4ksWW1g9Ymtswr590/pLASrMGCOfDxbcG
bgXEDfL1p3e1FGoJsLi9gAXqWSTDf8cix4iaQFK5A7Kv3hhicWCrgUD/r3yuEYdB
loQVlylyMaTXL4ySUW0PpBdX0j3jJENn0uB7kJZQdJPRihlOAzCpcVoyYS8huieE
HMJPesb2Dx2o/2aEOKdRbVGKP3nhg5CeaDgxPxtOaI4cryz4kBlh/fjK3cKGH4ya
JQM5kNBENIG7qToBUgy4k/yzWWO0AIfYf/OR5lKgrRWhFFghKSXm22ni7QbfquDh
75vcpXWwe5zIn4e4PgH+1KQQWphaugrMmOZgsc4fVa17UB0awq9wz4oDll7vpgV8
hDyh/IZ3yGVVXPB2K84YqegsemFFYW7Dh/M29wCvTEZVzBDSXZcc1kGm4ej5vqm5
Z9D1l3kDWi5aCuGPKb4c4vG3nxBjxLa4UfyxkkN/5LJYYIowK/gwUGjBAobC1eA0
UBJuLtJuek7iAMiqXv5eQxemTMaLGAO/bwLbLVCLPZ9WV3UKI8CkdIHy1JSFfHD5
4CrUxMLh/iP/uu/slQreFw14vCR3AO3EiqaK3ocrhHLFrmUxs0BcMECgNiP3WeE0
//fBd7l/q+S1xk2YeucXU8ioefp7BhlTQ1ETB63Bm5aSfbFn4VuegTCUfIbmv5yL
0jpfhp/IXNNLMNA1Aufga7LpZXRPmFKiwWFEuZUggHUbTP+rGXMajd57pmro2Ncd
S6m2ydVcnyJbZ4TFP1izegqsTv2FUP9YMJ022/zrHaGM9QMu/c328XkKBPyLdvH0
Bi70bmXs84t2ZWIh2nP2LzDUL/MG5iWFVRDd3INuN9cGW2rfQFCLfkcMsz/0dS3V
0HfkVFQgDhMX1l4DSzu+kQf5+EiJndL4gLIg+kg4kthLkBckYJtaHPfDdtmAptZo
VrSsjLFZI4ennveDtMq8YM3wHOQMSUic+imGU/1FpRRxAhD/TJ1TQKza16bcYlMz
VbxuRstxjO7AcKs15z9+CLTMpm3ugjgavE15oZEtVAs=
`protect END_PROTECTED
