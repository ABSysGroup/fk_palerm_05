`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lC8lgrOEUbD5GG1YdVu2sinRhJFUJl1nT66Yc3RAW0Jwwn9XH4/F8+FC9DFs0Kpi
Eenl+f6O4PqKVqaS3DbvY9SYvFGJgu+BRnxg4TlJ5KWJMfTOh3IgjqR5ALQcEDpr
hUHCpO+deC6HPtL+TRPhDevFgQ/51ftn63/7XyqDibpgeGKDdgiMcvhn0H1O8yPx
iO+YBqEkSSy3BZ+aiefGH9b4/wpAXhbkLDCje2zjLEhbXXPoK0ibr0WtU9OIYNEV
qZqT53wqtrI2hBIa9g/mtHc3LFsmWDshgxtuIKI6qAULJf4p62ZRGQqO+ANpkz5J
TRfUq7SPFNIXa0QYS1OenqF9/qYxPNYZ16FGE6InCl1U7bL6t3yc68Nl56+SwR5V
lCBcBULIqYIfk4xJbShm0uTiq++OonV41qC4Pe4fEqpP9v6x1weYGZcyhNc6Q7r2
wCvZU0eHHZTOKrRbPEyICQ==
`protect END_PROTECTED
