`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/iE3bakD3w09z4OlCw2xzrmgdbOE1N94rLnfDe3mZs4r6m73fu0yRaQu51p8fTaM
zpAKHrRLTVnfDCnqIegpeTeARdcoGHRovUtWMC8mKVI/5KmuIoJC9Eo19VpTgr4I
y1Pf7BotilRB/LbxbD7jlCF3mOXZ9hkt2FUEVVOyVT1YDZ9aBUilaR7vhPgP2BaJ
m/1hbDK2yuOY+ecZ6KUvJIi8DhEUG847B5x0YJcnzvj3z8SuzrJTreBDPvVorrrw
URc8vGUWJ/4QdnJWseV7MWCRju0ZQZa5f+GAbP5RfjeQ505DS4bJfxp2KWUhAy5D
TKWZTuNgnS2VsQSdr3nb8w==
`protect END_PROTECTED
