`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7vVl3g0vIqx2CUytVewlmR3bTTDVnz0sLiWZBp99oz3Q26PeHXLFS9feRyQGYytS
Gp+1GRnOopV3HKSR17McJZPc6uUywhtMMSjQkb4Q9Q4aAxxIcb1zQjZZ4iBvh3dy
658fTH73cx1Q+fltl3bh1QpFmEqJNczDnWhsO/8GDvrdQSUoM2eex7l3MXVPZjFK
S5GB2jgdarjWpY6XG6j0InA7Yq3N1yhoSe/oBJUkZXqTVdPqQ7KLKUD95ZHR1095
L9860nIBRTGCkVjAxEgJqbKGdc2AGJRV1ivIneWxkHoEDU/uiHRUB9Ia15Y40Yyd
tU24XRhre8M+/e4aKMYtZA4kN+MFujUpNXiB9ZubgHetHlA1RPD0PZzZSCmOMEIW
KzYKsnvNm2/4tcGHlWbbIzn+doRuPF3kgwXSNicGW/PRafI/SkM394axWoK0hhqY
`protect END_PROTECTED
