`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pIQjWAc7FxLEYv71ilCxByUwxvTfD4szUI69f/4ti8eduY+PAMPei5MINBiX71zG
7Q+lstJ7mDMAgP+ctQV1PnTbnNkGodKs1iHTB04TtcYSHWiFq0TbpJyFsELphANf
m2v67nWINsaBPnmsZ9Huhgw07F5eva2W8y4mpc5+JHRTCUY/D7ebRMvBXvo09zsX
AOa6UCKg/FFCngeZjqH1Cy0K4lqaNQoBUQJmL2YEXHo4g4GXwVuCLbGRvpigUE+D
dptCAiGT4mNV+d1i4ghsI4FzazUoTKgZc5TymITLH20eiwn2ts8JW4Crh+YQAA94
cv9OhW8Cl+2nc5LTJ0LAeLFPa7JSZALzjPzMpDevJn67+n6XUqnvcpL45qY8ROB7
oeuQTdHFpgG8MBcZlrdNqNWXIsS8B0N9YXFPlvDzoq2pVUcMrUidTx7uzXIhJRQq
iO5QUc5sgGcRbdIcieDpsXjUXKfNDCJx4chE4dWBJTdpUxCJabZGqvXzzG7hVhk4
`protect END_PROTECTED
