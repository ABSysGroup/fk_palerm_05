`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0WBJHpoklrV4F4YPJZDiNzG4C9FFiM0bXgY6yuRl2Hz219eG8VDdwG573kcqbE3N
mBPXQkB0L+hQv1EO/qCiO55S9GF8WKaieWOZndAxKzM1iQItjA+NBOEkyXAl9CHV
RmDwwMQ5YlOxZmdKDm+rC5LUjSuhYLO5r/4VH+En32FO279sa2U/0FlkJCm2EtoZ
66JCQ68xKq9mei3tCycTgacJtdiyyP1t5FMDa00jE2dYRuCWmMklPUKDr5VyTeLO
VIQRh22fEDrw7r5lSZaGdpMjgrXMM0UKrGeQuLUaEgdOjAOOGY/JXMimMg59mnnb
iakgH/btVn93WOoW6PkqUW/zzuRVMI0EngSIHmeo4cUKrUA81wuQF83+gY7zEzfp
9rCrmydRa43xT0fGE7RxpkceSzSfNjPXZOiIRESSswhRefyGFpKkadE7SI1LEr2z
7cRqVsPZXEbuFo3xBeyE90OiwnAZPN8w5ZmNwGcSOUp7dadhtZUqQvlBIa23KhUY
2w+kniFKRYYh/YGN7lurCS5zbaZrKexI1Xzel/RM0WNzAosVDUflTK7iP8EJ6g+4
aZ7WfNyntCc7CG4F89GvY+XZ+ADLN2h7q9RnkL97fcPSSgxex8WFlMmLfQ7cXt3v
C5t2/wGaejkW+0gjgUiNfsihsQPdddeh2OtRxLXPB5Wr2I5UQFp/KldS4350PXqD
k4LJ3khM6H6w5PKmUBHKlEn3CovvicbI2CDlLqUi1e8rroP+04CM25dSxsHtccB5
AYgaz+k9orlrVGVmwjt6H10vmbReT7FJwv9MZm93MbVKwufvQocickQkM61YhgYz
K05Ju4hRtRj/tMpmYgODDjghd03zxoradHiNdlG1mpg+0bd8k/xq4anXaeSTCd+m
ngRHug7OYnfFMvFfngPJJTvLgTIzkOWThZeBsGl31AXYESYKnDi7vHrfmmJKGl2V
uvO8D6snuPlMskShVlqbd6WcOgg6p5/i0GPLZIwx6mORu9YMX7YVYqvcKx4JFWVm
0kEU7qpznDz98Cjb4/Jj8YgBcfCbtwgPyRQOgbYXuAWd53Se+RuybMhTadUy2AxW
kRnM2pOIMW6cOfBlttiNCSPQdDTo5rF+N11HG4m6XZtYMChq50RI0fN1HoUv0HZ+
DR8tfFJeurleL4LqyXY0/qbKFWIfMHb4+cFFYdNFI1ALM1RtQmsI5rqk9wfGYVR9
yBvPSJeKTq7jS9OAQbmDsEzGrc6kjZ7LdneoKHQB6jjIRFDBeeVoTRMGHuttco9v
xUGuHWclEKpGnBhHYEG6GpI7gTVnhJUFBSIM9+wlKDg=
`protect END_PROTECTED
