`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N4bdTKe5qoB9H+lubSTpJhB0bW8cMOBiDr2cnIyDn7Td4i1x+92fB9+ne45+nocU
yie9gLdIKEuqL4XolYGUbn+VuJPSDK/Q5MeS6Yh4rHurGz/S4tnFbrvoJN0VDB4v
h8hp3BmYRRy2YHz2gRlXv1GKYAABxBpGdPUMZnsjJWaG2ETHc3kc4crFYv/BzrXy
3ycy7SStbN6s1XzAknYHPRA0zX5/kQy+NW/X9s3Z55VDeOtwe/hY/3FU+/EuSRn8
usAuCWuK9s8IZ+aYWKOaImkC8nh3De8BgbU6uSOvI7n+oMXVvilCPIyeH5611lQb
Bf5nuXqLgHGr06gfdS1zuUrbSOxjS15jXs0PZH/ZMYHq5fSewA4lMt3LEl5UtXGn
yE7QkPD7B3/53AniM58jH8bi+2ljUnW67ZiNc6m8VElnfUOaj3rPSGfkpcOxSAYU
WNUKfihQVGz5Slg4oa7jLn08QjbXEdu+4dnx0b9a5EfM77tL+H+uu21lJqhPnchz
1hNXlHqOueQ0QRv25HXrmG8uHr+GrHf48LRjFI5KO/dSCskuWd/oJE2tFFAQFobC
01xlVenLuftrmUubkq81kgvbsjR6vAK1HCxKxR9PMR2KN8CBpxINX39umPzBWXDJ
2j9v3PKI4hcwrgLUAavDBUwep43BNuoquAeq/iArUSEcN+I1+ZV2QgBKxl8jgMm1
zOgBONR6tQWnmBQ0rr+9jLVSw5sXaiPg8cJBP1EsAzptMqNAF3Jcgw4HaWlXw12p
8M2Vkicwu2k4gwgQTDED/hxchMSFI7KNA96whyTklnL15DqxPL0uRD15h1AqgB2Z
trVzvoMqVZfTLOZ1vVwckhWU00+rKVNfEPAhe2a+nTVaqzS9x2IikWbyEAZrK93g
7Xbo8E/WjKpnS4YBBaEayJyLOT//doq6zTeCeLEw2a2XIi7Jo8rOYbbFPJXmX/PE
CJG5iyceVxOltsubGIBlDy/xJ7zS++cQkAzluSl8Mav9wrBDhV6PapnpWweB3HYx
m5/r4j5V3vaa8d9iZVSFPdOK41j6I53zPFcdWZ+r3hpYg/GS+oEZWRsMrAeV9oz5
prxCrC1PYQtbKZUBIJuR71fyz0yOmGBaqBYcZUKGwP/9rF03EyXMpMoAp5qWuIWz
dL/hcwDi4zZNTpVkPhuWv4ddcFA908oj//2Q5VfDlCspWa1gUiyeEb9drX8gmTNq
aXAQQzfOSBjRiXky78fMcFZ1W6wL2XaXp3nNzjjcBmKfJL6+OJBwPlqv8SN1/+LA
20U6y9ugBhu+e0/V5+R4bsTZczPHOiIj8/om+aG3mkQdRccC5ZzOnQsdTR6AdKTt
WK6lara6jnFUBjp6fNdGZRPBZgzXJaY3l5djRH2rtP3KKu9dpQnruznor2UCwvRS
60TmgL4jEVSTWo/sKUWyUe4kdv9iV9J7gffeFWNCQhnlOM0EAx49cQRBtTQG0lwe
HlsjjT8IT1BBMIaiGEMBAj3mYHkN44ekC6YRUaq2CJFFyYmnNrZc1J2zqXYwr/eC
ZwLB0+0eq8gYyu1Gq7FgLO0kN4g1vkf3NJBQGM9L+U2/ZpTeDKloUiwjNS1Q5yLS
yYlyjHN09iJnG69wvgbmukmKUOl18t80/8dUsb1+pDsubFNPen+GCU9LxxhXnZ+1
4vWNP4LRVlNGuvHT7n+NW+yuwJM95/cINi4jWdVbuIthkgyJTjgajwpyUDpCKytA
dquhNcVgQXLWaOJnGQot49BFyZCfb19FdKI43YHo8qgrNt6/XVOIJ9lfvZ12iIGN
Ap69wa/7dO8d0KnezlOfZPgtx46qCibEEYe4XoxamMuClpvdV6A0RktKfFahKNHE
DLg6aCWVXFSkIcNarOK5l2dsl8LlNBuaXWo66Oczh2WD6sW70cYHD/4QtwcDCs8O
+AqrBwNE5onOg4nKyrOGolvS45YJSx3MBkQq8J+dCNS9knb2fnwk50ZDUPDtKZzo
d7s3rHlMXXhdYkLlxTf7mrXBfuEUeJno6F4CvgaEiaF3FO47hMAj/6AaIsT0ZvEr
z6Itc7HUu+XM2ZPrt0OsUAS4qo2pwKClC3UTHXh1DOlKQeqZMJTKt7JK+r/YrvB7
QQXPOzcfERrREPO7ybZdNzMTOYLprubmsCk2qQjlACePzEI8bfZ/rsqYOzWtM21a
QRQLwwvatwz2JdUfgjtH7ad9ra8uDKfqEWoiqcsxR5M/9GxnRX2gloKpBNeYhRxA
Ge5KipH2rUJXarz7kAGfY/XFJNISXSwa1j0AYPXTAKCVtaPwg5vZd2qUBsDcjKqP
5DUAsH4Pr+TUSCJvK2OO/vsaTFUKDjcv6hka8i1OZsVmBoWBYYA2moVYRyOm9Cn8
`protect END_PROTECTED
