`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ANSPu+6QtYIw/xL/ri7puNPyNa3iLhO7qXFdQhXF75xNlPdrdgjpEszUrD+ixG8L
ku6VG0yZlgr6zcFVL6wPl5Es1cqhzqsC1klBI6kh6KZowq1refKMj2J7gJzzdSxy
8+H2HRpfuPi+4wdkxXIA6xHGzAfrm3MvXvzJeFBtS2+DpW2TcoNeF/ankrkkuSEX
7CHs+51Cqhq6zkD/IzklXZNcqnFVE9g7EOApx3J/wprthPaVg4wk384Z+lVSHNHP
8FmrzzZx0p56OwSc2lFKjw==
`protect END_PROTECTED
