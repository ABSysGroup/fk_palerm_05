`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3lxrf3kkmSQXWeKRamekFIkMBYMjpUVjqEMUDv006tHXPWb+uI66dIKOixZ16Q+W
+BFI4vgNtzV4fxx7IM4Lx7qYrqGr47qdye0h2nMV0WJ9I3e3uB+7aR8PYR+PYxdR
LqZQ94FwV0aw19EYpNNQM33Qw7VoEn98U0BuIZlvtDLIOsvhtLaTRmsS5wlg38wh
3cwYsovZQEVlQPc81H/lRKHEP2PM6y+FW0IbObXf79tPz1EvJMDwE3bK8WC2yrr9
sZogaLdQDKs1Buj694JniyUcP8Ojy91t7Tc6dMcXNWvUatAVebcQJ1xBOAksC0bZ
FpS6lWt3Kwt5lGRu2HhKeQ46yhbDC5LZ4yDUk9ECfFk2LPDNxM5rJD7wdIkxW5w/
`protect END_PROTECTED
