`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/3WiYyO8hOl/T7kSYKksNWDGEzDfWVt00keNfrxlqn8hX9mJgea/C31kg12dP9Pk
I7lQ5JZhcqXN/qrvl0kos4/IrM0hXL5y/RtimoAYnzw9BHUu2Wv+eG+QePjmfd9T
4umtKkSAkj04tYvGFM4TIQV9yd1NQfY7pxw4d3oWbd+QJc39iYrUFL1sMzgmEhPZ
/9YX7xKCFNuccY0fpyXGFzzFXihk0hvE3qVXNwlUtfpv2q+sj/hOTEZZdkLDIXPI
L7QFi4TuOY/bFgx1apYHL4oSamqyefECdKr6OQZx+Wzcmy/qW2lB/z8G2ceaN5P0
531hQxrRzF/vRQ3bqcINWK7WPRSOvbrDJQcibEMkOBZWPXKAgfE3NJYuiMkSorA4
eSwHUnOSjANwCzO89d86jGWJ2fkR3pA5O23udxLqUHE=
`protect END_PROTECTED
