`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zjIpzb5an4oUfSnQNZWeYGX9ZgFpV+lPOedSgbi5O1BTT4kpAJeCHVd41jQrYj7/
5N6XNsqfsbSHmjWB2KVI/ayUEbvRF4wQsC/DxcSSCeX1gT1WJZD5c9Y3EEYtEl+i
53EeLM3/q/Zull8ouIo7+l6MxX+1kZBBkbJeWuy6cA2DQm0nUOEeVn7uo7h/Bdax
8Fv7iXKm/FcgThOZ4oLR72xP9rfxhCKnZXnYHg7OXU35FsTYnxj0rcsCAwmt8YMa
RnV1HPJ0KPH34ITb0vSu5H/07DRKWK4cdY4YRYIeXQx11py/k1g7ww3jw4dj+5v/
LOIcKWVdu94FV6LRytymRea86hrHT9M8sOANF2ePDJonm5Z/xkOTU4m+jugdLKUR
f3LRv+z9q9NVVK8D+QmkAHKn+r9i0gpQbLCg1R459R9UE3MxdgR0avQQpK/Zz6Nh
`protect END_PROTECTED
