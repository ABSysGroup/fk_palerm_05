`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nES+PX+kkr20kuH0xpor138e3XmbOjNTolU50yTrxv2yj3r5Pjc9QDEfZ5r83Pj6
y/wPRLvZUUu1KyGfq0Q5bHlaKHny9jeqFxDem2jG3em382cBo3X3sxw/AENnm2iT
O+Ia2YFcPQGr4vp95k3WzeNKRxf52J2TbJCGN3vXHztM8sEwGzNxuGsf4NzRRbfN
fwXl0k8nofodmysb7qT8QYKA1jQEuBObL4eCwpXxq13wGerMU7G3T66qS+EKNDPt
RCnw25szgAzm+BDt1OuMjuLfbqI2TBCu3Tl7IHAnsv9KIlpg055oYxWBIlOGf0ZT
yxO8E1ylsY3euEGxlaiDbZj6RoUiHYitCNAO5OUlBMHva0WJ1unEg3oWgznga+nL
LDMuvSA/CgVLCGQD4I/8gyJenOCA4V6S5xHkHhWrK98=
`protect END_PROTECTED
