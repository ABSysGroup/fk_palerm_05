`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pT52MhVl2b5nu/tksQFPPc7VdC27a8y45Q4ywCMxoMORr7aK1+aQJlMYZ9LPjlL0
/IyyLMWktlvg6e5JSjnvapbrhRCWDVjukTwHZkB77WyLtKfhVTPFfbfjQ9MX0/td
Idb/5MT7uM/1rNOGctf6A7BzxnSGuiiEyVTjRPcGpdKipRgk/KClPvUM1J0diFEL
MK0HeadRvilJ7/ysNLwy56gVoIZp3L9pMlv8Auv/AGAcDTGel1GdzpilEm4ld6dD
/bAWjcxV8W3+9ciHU+Ys7I/b8fPFPCk5wmfUUpdJmU/293ZTGV8HUGFQzLvimetu
hEZTTucZIJM7yOHO95cj27KhM/6jQnVK4GoLOdeIWh0odSLhKUMC+gNcjInD1cDk
`protect END_PROTECTED
