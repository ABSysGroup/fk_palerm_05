`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0SMFU/5tBERsOWFfeq9Wc3IWmG3bOx27F6o+aBVEZuhwhWvGgZm/0qLeuqLl7DMz
LYw2+biBRTNRLGKqDWJfNWJ8XjAkNrqUMJmpw+aEI2gSUoACSY6C9myEhUcoCPu9
miCrz9J7v1YsKJzj4mnemP39UD1OjDBJZ/mexXGGu5U28oSQF2/gbcPYx065A7oV
s02ryIUog3sLLTsrMaEIzQjoPhyaRWnihPp6jtT5KgkGJj2ibAnFzcnM7Z4RQxot
FPUzBuvFxS5tgLRvWtNr+c81IvQ1plC4Yck6tO1yHUHRRrcqZZFGEsbnoPt+eUHF
bMrv3rsf8JPXOBtzqcq6nee8A/cR6ZeWQHTEOD5KDaNCvpYns82+7R+llOzdnkVq
/5f1mZMem5IRmcBXbuxdHlE9uz/5OOeyyBwhzG7a2jhLTkhNTaaLhOID4hjbsV5g
NyvQMvOPNCcWnWgTEO9K4WTr+IuHh9DQIELDJk7ZXk9iVw8z23Zmc7AnD57+1vGa
2Pntm78cdMxgNU18jddnJU8RemwjSKvwmRCF/AphZRfGbGh62n+JgW83nDaEvlA4
UIbmxdGap7WRffXbxIsyTyMQfptaAQeQJftX6QEWl5AOW+dJ7leCcag2Wtvh7tju
EwoXg+4mU9VQGpwpcQahMDVQKCuPp9b4UlqRf9hr0X00B5mQ3S91SWQwAjbh6iwk
5g4DlX+iupf1nCv01n6a27japQQ3czqn6su+/28IT5BKzAh2Yw81DRY9HC9p77L9
1ZN0qJCT0svW6+pt2TU7lZhktQYNmHxN8FQTs2R//iw0n5JK51FpFF9QH/O4Ef9j
e1ghrgvnp+AOg7sw5M32qGzy9JBSPuCmHegJnaUb9TPgp1s1dxmRMtZ7W/i6Cg/y
wU5rJEJbgRtF34p8+nQ3eYkHUREsAgXIsJBMtZTm+Eqvo2nTS4EKFQIxf91RDIar
wki9oGro4R0yAWA+y2vg3eXxldJkfVdG3jx8QWrJTLQvL6AEa4LFpMkTkMA7ZCPv
`protect END_PROTECTED
