`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0zHfNkpq+AUI8jY0gi6M6+q8o6Xrt1bjeqNjKtVsT76ulx+1wM/Hci/x5Qd4TpVy
yEV3ERK1D6bMjZyki9CH0QJX5sMxyzSoTmNdbXhQLVX+aBCQY1nQngWzB+Yl0KPZ
ZP64RXX2a+7j5SGQN/1K5eHjB9jmhUDkxKJ+ErNCg7VUtSX3WrMHdPtQ3uuMu7BH
P9uQnu5Y70JC0m0lI94dSBE3dcsKuK54JghfAPvnHauwLjXN/eynsaKtEnGU1oei
ULEspGqS5dVnOWfheKJnUD8Hi6ZO4WlyoLl10FsesiYha+bnzni7t+7LkHA4FQ3Q
zXag+fzfKMU9xsJ8xTtrwjHnsSLmhNDaOxYlP53BVWnlXhsx3p9egphGUvbbDgrk
Jn4+Qkp0ENwrvW02W1ZyjvsBOGVqliV90WDzRNYWHSn+Cd4kYZf+cEDGMN8TBYg0
Zl7dqcwn2LMRCI9sZdiybxdqLVGE+BK7psq0H942+O7qLAvdEcYQ2QW4SUbFOjCv
1XrocSWfi/XqFWoNfRJAKS7L8HA3OEHE3dx79GqhvlFZCYd0nREnr2nYBBMSTK3M
fY5q0DWHFt/ag4dYi4eHtWPrP6GfwFinHF658pOumkX7Rwjn23L5DgTg+vzRbs7a
Msju3ka6qZR1eHWJYG+B3Y8meuTrn4ACQWU2NBmduurK7rik4LWM5GjsthYx9BgP
ABosBPL7QTbAGVUt5ZzPZmp4a9HUudy7mnePcUuO/kBBsXExWYYF09SgcwHZV7UG
J194tlQKqMgmsPUmb8uv4EgpLgAozD9lAX/vj1IkYcJLz6xVnN4UmmskX2K2FHkG
e3esXTYOaV+9Dqi50pVCbJiy0zk8qi6WiVrPCa3nXj/BwEp/9+Hs2aQY12BtpfSF
4AQeBUE8nBIU6rtxxf0coxpX18ag9W8tFfucqqJ/UZAaROdybl7XJ2MRTascbYUU
g6gm3f1ohK4Lj++OG0M6/lEpend3vzUz1PYRZ5pnWATgMrVzTl3oi8PpiyR/F/Ep
1THK1dGpIHqGrxhgIjFARX+EL4GJem0HTm7K91Af1BEwWYOvM2AeAvwvNEzeAkvQ
dBiYJSCRLLpyzTTiKQCycTvfMftjSpjFx99A1yhLd1o=
`protect END_PROTECTED
