`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/t/ItZoLPfBwwg4aDPzs7qTO6eS2NN2QXc0LxWZmeRWp8edHm515HPw5z/qOSIec
G/TYnypkqgXpJvdNnRW2sXlZLcSZMRopN/ivzqLm1KUGSn8naywhncqkXR3mUEjv
yQruO82iepRG+gZQf/olHiR4Inkk1NZmevlGD8AqAb34YsaNUf1zUPrgWtpjhKYc
O5WQTJ3rshx66o2JDBU3FpVidN7xjSVTaZrNPnnBBkrZcDWPoMAACdBazfNRsUUI
frKcmv7MayQsRht2gSlz29fAEkTYlySZc/B1oVvvlvqISL3IqFyjPDHyQkkhh2+5
YfW23+JsZqfZ/LcAHVIMTiKThq1+tLkSSyK0oFKWJbXL0JVlA8oR3PuihJpCZrHE
ZL5aY0X/NbhqYM0JL+V3iGFcBvwXJh0BGzRUkEncQsm5zPeKmpYBKgLLDTN4xiLy
vbsxTW+6/Qkl8jFxUgNSz9kKUQkrIBtK3Dw4KMLaMvqcabwnde1AMAnBHLzsu4aU
B0H3oWh5i29ekPJLECaI9HLd6mziukSIJuZrrkHhIqVQa3O9mNi1z6FANPRbBleX
K7hqqJ84tMKlvB5ZdqOQwdsXpqSVLgWy4WxWE6FzJuZp1S5elLjL6t7eLGJl+Q1z
ubkE2SMe11KifaBAx2Izxt+qiKU5kfHLtmrxz5pLGCg0leh/sZz8VoQQkUXLj2OJ
L9MtPAXJcqCMh+hMEZDhTT1zRJoO3Nutjbxo9ogVnPpiWPENfKUwo/pY1dF0koj3
7YXTBWgvMg5ZG381KP9T2vmuhYYcFdM3JIW6zChtDHU01mgAFKCmdRxT2qgMKLOn
uthKxGerk8rAmxY6nmgaJW6iF+oRLlmm/oSqgu4TjNbaFGqI+JZfNOAyZ8bHdU84
ZVDCG+mVnxPbNNiZm7kKTpbSEgRCCesW3jhBwPD7WA0qs7aGVcIWBISJk51kCAfW
ZDfS32zJvFfEV6UbW61gV9xRAq6xiZ6DK5FVGR5+L4wdwfcDwj65pMDwk5+FED1e
H1hLQxGavuhvDjaRcofHLnkIgbd8fUGt3F893JhtWWkDKfN8v9J5BrricmAFlTRb
CbDNtXO38zRzuJ2scCv+X30S/63Vmg2wIM0M0LFEtsniN4TgXdfKwkSnLh+mpGek
ZXW84bdvp6be5RHiEEMC/n4bC+FQN1bzAya1CjEVS8pWAN+rnOkTp9kvcE5RSoX4
nijOpJR8SoqmyLtKqgc32rsBopceoOdgzqUfBZpzLYshK/R+lk0HYpat1vfhnMLz
iyx7h0tJ09hIMWFBgkPg3MpE2GiVSurI753UDEmtnw6VQ0LCBgj6BPMbLEDK3l/T
4ADfsR0pkUarDc/BnfUDAAUrqgM5BkaUMJVvoyAW1Lg=
`protect END_PROTECTED
