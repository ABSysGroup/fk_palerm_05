`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
474qRtswEq1v+zmzTMpwSojQnEuD4S0Lr9A4AQdoDAgYKpLvvZfY8CWsh+IVnS1M
uUae5S7UdIHThZLotCtKtW4cekneDEcT8lLRRwKlGOCl0/b4tcR/lF8kKLcR9FnE
E5deut3HWgGBCaSCD/pNdfrMnFhl4Eygfo6uFd/PcRItf4o0FoDHKwSGrmzN/pU8
pEaLi+DNL2zwGnwiSd5IWQ9Tiym14ZDYZgxfEpS71BkjDM4DxYdq7LsPTUA4BhkD
TD0esRCTgdM39H8zZcvJ+sQ5DvDYtSHeoliWLqdKhMaa1lYcrnKbFH4KAhh6h27M
HzsKLGaY7C9DB89+W6do80mAnvV8yiTXx+nuempQsCZv/C1DAxA1P8D/Rhikd3ku
L4RXeprX7VmNOBciS6ddWbF/bhWlqyMe1xk9at5r20y2vRpBqPpcObD6PNba35Us
9/Fe+2uJvPUlZbD4tq7N5nTTyUhcY8jT2wfIo74v/SNgQM2OWIi1PxJc/5VCrF4M
A0pef9wizKvc2lluyRgtkqGnZevRS3Qd1NWb2xiwvEl27YBxFA9rRuLR8zG9HOjY
W/7WPyAtCxOjo8fJEP7uCkUMisgirQahO+4bxgPi/2ta6aa9L4rKerKVNVJ593Nm
iInD/pkaMZk9mJfZp46G2Elqb9/TUky3vtnt4grgincrEugkk3BPTjKSx2DsPeY+
EVyYPw8zQD+c/eU4OvhkPoPtdUJKOFaE8bMXx3600nKqGUB0OXh1Ry3FiDxFKW3y
pn6jTXxKuqTEiY9SLKP8JtvAJA9qRjko5Uozd/54ZiJOr+OApW9hgNT2UhCQZ93l
`protect END_PROTECTED
