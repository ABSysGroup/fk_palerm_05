`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lCdrVOhMRbAMfZjQfDTHDY8dXY4N9ZOn0iRQv8UDOTcmAQdcUgpwDph8bzE29Z4J
62qoDtkmBkkir9GGS6ncGwpOyUspBhX6JeATyNt/2Y461CRF2wd96eUZVwLPENN3
tsFnvsIMSKgC7yHjT2S81tXMmqFF6f4heW5gdH862mB3p9Bj+hs5/M8YII7wdJh5
lrKYjJM6okmpa/rnffBONHwj8ceYcHXi6hhw2sdxwG2nw8eQLuKz+82l+P3iS+pu
KUr4tlmSdKDgqtYnzaC5mDBSSdfXIqUON1SODcfluhaXn+D8CG48t+8Iz9Df+Mem
5la6J6lvOfzpFhfC9SKwpff8ZPxaYEI4rQdy4Y1aZmMu78WZcOGHo0HoG2m+mW38
eEz1vQ4w0EKsBKRjFneJooQsdMah6r6hOP++7lCsJuIRwkadCmu3I3bhRt92fX4T
iAZjeh3Q8DaED/5Z6930Nttz8X2wR4xd42Bc86jPqwiaVcKwk0abNuGkVE00Sq30
2WbN2osKdadv0cbLnYSEJUmKXwCSIFKIo0PpzrxM1+tNY/rzPSevM76PBWHE2A03
mTO59aQ52WaXUMML3vGOy2gyXQj1XD3j6UfqH4qk4lOJYffOsxoyMVM2kVMlSaCF
ykXe+v2yuwCNb+xmx5esP8YUmJ036iTKBbUkd2eyW8e1N0cNqUM/VV4IJwLO0KmU
nFX+PTPgP+gPefwoYt1bLYIWPhuwLPeoFp6Zx5S2gS8Gg7oztZv4orCxB/aVeGT8
frYTBAPEeyhFsfzxkP9hNLSs7ZvkBdRJ4f+xxXGwO1g=
`protect END_PROTECTED
