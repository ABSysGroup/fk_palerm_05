`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5AuKFt8M4FGRlHybG8i6JFKpI+CXMplpvfxXEsgZRYWJ3hLh7PeG7IWZBhKSEGRF
A1ik4GQQKzcsJAxKVTE3g5VWAH67af3yDH9k/k8G6P1Z0TfsSKI+k3CkeuM35p2E
ImyxxwoPE2nQ2kjO1fz9y7STcHWUHiPtrHKqPojmBnCKcAudUMcC0pUa7gRdQNSP
Xn0BSF3CqKembrY9LD4aWS0+2J8NXW3oAzx53K2H8Uq4u/ierQINbSlsE4JjWmDN
VIeCibGwoL8FR+8dYSz2gVhQAY6Qhu/Un3AB5SjX8n+a/dNkNds6yd7iqQXLuudi
0fLus/Fp02jpcGDtzBLXg8mJF6ImhCrWv++qmuFNitW3ZGUjLtel/D6fq1h9H+XE
epgpbkewNIQBsyltfRaasewM9P6hvUV1lKCGLwzWpOg=
`protect END_PROTECTED
