`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RGOodsutqnHL8BwvKCz3Quts4qHQWMO6r4W/zRhCFPntbi2sehb50yGc0izSdU+A
qTnlGf6OQ1Tu+fOHgzbuxeq58BphzShyjxHgVEbLPfcPj773mdBRlVwcQpn/JTH7
UhcY7rYZm6E9GZZ2sSTHT6RlLVdbnoQEsa+IArtdCzdHi5cBFzBqr1LXu5HFUv0d
h/BqEIkPPdQamCCBptcdTbmsZTjATouqnyftoBegA3r6Y21Ns0Kd4vSCIwqXqFe0
SdFHLONQD0Nk37f+j35gJ8FR8UkTacRkaVF1EjgsjlCNivXsZwmVQbfZoDI0NiWa
9GBjoFxvY6rFZXwOHvvzkQwdfkImsbjt9Cgm2z03yEZF/2CMqacD/XrbZIu+l9GL
0p2EBJ7evkMVMmFAUHoIojAP8NIl1dPW8c1xF3w+ixU=
`protect END_PROTECTED
