`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jf7Rqnme8q9T8uBe9NQwpXmIM0RNhpPeHFqLsLznkeR9N+zb27xAo1xehhwcsUhW
3Tzzy3J0OiGrNcJeCTrwj21CeyDsIJMabO1sD+IkRL2heTV9VSHvKW5ym8//oczZ
i5RVtgfG/PDnu3Lj+xAZaaDPsRVpRe6opJXbuu/vV0KCaoDPI9iKJTiMUkjl0Z2r
NCJx/OrSzV0yb+7Ojb5ynV7L3v1tFZJ/JHDyr7qHGa3ZCNgzW3c57gHLFNdzHfNF
udMUrVtwf3/vVcQgGI1XgJRCkObVMYL6lEYX9Y2+I3qRWFnBCmvFV2nbzYgA0ZU1
7pqbhvCz6J742fOaRDiuYTIGfUH/yWiXgH1ZxybhlfFCDR1qKvlVGPbnD0ZoFRLD
L9f1eF4tAO0XhdiHGDv0Gmbq8r34+7W56oqJHedz4hkNX9C00m0TGx4+FTsd0Brt
kCx6u5h9I2/MA+gxLIKmVwKuwJ6ZNjE5YV8Nbt3mE7crDX5n2nUYNfrtGE9kbf7b
CXW6VzJmXNhvxnJKmrZ4UV4jEYt3ZHGGl+w1ctKfYyc=
`protect END_PROTECTED
