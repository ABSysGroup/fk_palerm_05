`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oxq2V8fxvT0ZJ53dX4KF5+KIush423Wti7ob1MPdCcSNN7LSlRK5iVqTri+2SZ+j
TIzRC09qyf9WvorBoL+VOcW1Qf4kZiD6szBdFH0sjEMmdPfrd5MxhhAVg/GcY54g
WRChbuRp9+oDEJwYhMwVqqwELqWCmsUoLvY+3g+DWtM1vBbUZW5HPSrkz/SI5GSH
vkVky8/OVZr+wRF4On/KQnUDRf2Mba3QYM2rC1ZEXALpEIB7pKW3TcVK0ngtVR/7
dFbXoyu8CGk5q0LKqv1rUoRTUJfsrrJZ+k1lb2mfLVlDFYgG0AVZXSzEncOMCOhH
8rPdcNCjAC2eE9BSZVVknA==
`protect END_PROTECTED
