`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cJbiAoFEBQSU1KNAe1ePSp1B+HTpFfBdIymvrg78HNGFxB4VhRzKuG4kVGeYqZtX
Duo5NihnVJ4Jym0yfYbzo2BzVuiQn1eJSdVYuqALFmdrCLQtZ3lHTBC2lPoXfK5p
OO4hGjhhRwAB8HFSIRwpfkhDGx4mH70GkbKFIO1Jqbp3ZF+aS5tfKcVRArtz9jLe
RYY0tWWcZSNE6U8J8pv/rIZiXKxJsgNHB+5oGB58qNJRHSu3gP29fyHcnL6ntYyd
0Ogdu4u3d+dmtEj8SAcLnQ==
`protect END_PROTECTED
