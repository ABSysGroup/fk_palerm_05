`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fEwM+IygQs1O3kfhvca497PRQydGrRFNGNupcv0VF0/XeNnjvRRYu3qls4925/A8
V7PPaV3GpeBuYtJyYHnPtgy6zjbHbpDId8QBG5tV1dzYkJeWx1GhEjlMx1tQxpOA
ZvoRVOma9gZx2Y+q6xDLA0GkazTTUnyRp30cpbCbR7f4jo/JGQ+jNLKJA01QtX2T
Gjae7OIhcTNattFl8zLUabj6EM2ACPdulvpDQvz3p6gWjjZvypSKaYt1aGciQb4h
4ZaiC0bSB2J2/ecJASpYMUHlTFf937uXQHvnolHqjOJTSjeLL825S8mW9hXBchav
qwuUJLoQqW7+ZAjEFDOuObKLbd+/rUwj5BsUiZs2JQCuUbjE22aULJz8tYrAlyxQ
nItQnZHADgY6DflIGssyKxhjNBgzirjFq4taIgl8LrJPuN0r4ThFM43M17K48HIQ
OmOkDtSlXVOitbCJJ7ZDKe0kmgxCWJgam+5PhllTEDOGFbWHHcUD0FuuMwF/9T+J
tEHPVf+Ai+s3Sx9n8+H/UXyZJGctWZBZqr8cl7aUdFOUL38om1rPcwRPfeutKB4y
fzepwpGwq/9mtZ5lsWfT07cKF6M+3MYoYKrj5cnUo1MWiCpu09rBfdb2wzawvvGm
IqKYMrouH/t4r+2n+tY3WOmK9vMk8vQhv9Hd+IqRNbQEJdsPN05tqG8XiCkWasr4
LT4+44iMk5y4cQY3txTWqJVA61jv8PTVQRds4bTXdnaiKoD1rgy0T2L1cioE2CPH
EmaWAU0Xv9Oi3y2QlRXrlCYas6lqjWh0u6ePM254AR5mxi2WRAe9EDn0ja2wSuyE
kjBf1gw7KbRndGB6hEqv4Cdxb7oXbAyxbnTYlIo3Uq1KJU0BFlvw7a3YuXJxuF6A
mnh9oBSDu72umOfKKvLmWKSIajQmxRge0cdZCcmmoN+buGM9ApsLO+sRjLpJ33TZ
+H7zf86qKmLVpMv2rIEhp53/z+v2sqU4AdFgX5Y+anG7L5KbyDz65TbZZ1K88PV4
ERyWGSLJvjQ30OcuwvOCwYTOSGSEYgYZYw7sUyHBLWH4wj+66puJogGms5xzGht3
dXKf9TGQOTv1Q6eirF3Qc9bcjVUw2jxyMXVT/JjzV9TuZVx2rJYsQcdFxmeKFaiC
7wRIwLUtLmEMw/PYQ1rvpVLV7as5oz68rkMGJi70KehwBmf+7jr7R6QMHn+6DJdl
uJyCG7RF6vNYJMwZPXr+e8fUuHyZ/nii5ppCJykBBtTYUHJI7+YDs/qOaTQef+uL
kDEAfqFA4G/PdO9YEXLG0b7qxAZj+xT0C5vTXICWQ697zZROzySjTV2EkKhd4BGN
WoovcdzHaFHF5EIjKDMGv1TcT/zuk9Zuwuhph+mVROPQ04uRPBqEAPku4zQ+Y/Jl
iBSL3XtIdq7uTkjQQnLQXGvpQl1LMmkieYO6EK403s3B+7A5+aipKRyvyCjLScrA
0NmeCadxJl9nJvoF29fwmCeJho7M7hIp4XJLKtQfrMU9L+EDAjnB9sB6LW+E87zp
l7QmTCvbdvly2cApPlWUtGMyL5Nvjy9NvvADIUDkmgjO5H+1BeVazVmSHmazSjPr
yqRIw4NVhid0t0mgJnQ8nmxC1Rmf/XowrwUxXSvQPPHK2or30+179zo+HxH0VwMr
Za65FvEiotqUo19nyJ/xtoHlqeSoc/lRRz+KbUzkyNqmJiuWgd8M0yr8y85r5azo
XmsK97Q5uDtZPbRWx29GZB7CTvGo4wNDD+f8nl0gX9X4QQXpEh0wUKi9KVQ0vxNB
o0lSffRNFkGuUbZEV2y7hIf2LN6KkLiJG3TZwkSWkbEzCFnA7DEg/KZXuheOrkSU
HHrVaQAI6slPmOooLW2j0wetZCLCJ3aZ6ndxf4ENsds60ZLKTaDxDaZOUKSn+wHc
itAbgV3zFaPoIAL9kgd6OifiMYCPvSDNl0FcFMhbXfown4yvRHbQgMtMQAoHDUxy
AY1OjFSutm8OoRpa55CwKvkrAo6u5qK1JtSqJCEKDF8CjSNxzBDf1wI2IJFGf1Go
SYbGnh8u/FIGq7pSbxOF1LhXxJoEVQ5UiZ5OsbjH/YVjtSBuiHaZfNcRao3U7Q2u
+F8YHQzDegzkBlYkWcVUJoXgJcz3SguRxCARC+Q842BkDwi7oyK/HYfvvPaTyZQ8
AirTS0n8/jdAhwPBFnYkUotno4LunWbaqqNeiN6YpIyHDVHm3rBP04BRkmo6PLGN
sxoFqPIVWLTLNXG6jWQz+XJB4sEzOL9hh/eeCs4o0dpIVHc9cyBFSbZdhIJx0Xf/
08ltwFFZJi9qqSuCh60CMvnn/srL9ckFkX5z6IrGaS2RpsbOyD6p2YuqyB5tKdWT
Q53unYNi359SnlQ0wRYweXAIYa2UT5y86YhN4qyyXPzXX6zTluok4OK/ElmVdBNy
bZQ0OMIOOSKi1fryQjAin7bqZbQgM17lxIuEO7qnWsNoFtBeUnOkqxJHGdE9F1OJ
cuOv7c3J5o/RIolMhLZE/VJeCJPRom7EPRyMdFtoUy0tbjBfq01kJ43CbDbj7djH
ue3twxRH5oS3IdIeUvWRVkQ/dK95ZF1ukmlcNyZfx10bbpgBnDzlw7Hg8uHSQVI3
yfaXLQl4TdJnY7LcAgPms2IdF5mKfRgnyDEHuKkuiYbVVoSzQe5dIWYrS8cL9LHx
b/wKViFs/HOoatJ1Q/LD4PKIPhGxUjHTkuFsE+L3juK0//uqnowZTMIXlDDH+Bqu
1VNZ7lTI2wM+KBPCArN6w4UCujX5whMi6GxcarIWlF0FJ3WtW7Vy5mIxz4kLtPv7
YP7H4lJx8bBcDrfPsLtHNfzRkvWNN7gkSVdTRYQnSjQumQLAk0UFkZL1eLi/YFdA
CjdP0GigtA3K3E8fa/b9ur10zFyrGNAX40TdDnwmNpTAH4xzT1yLcEKPCGUJSiqU
nOP0bKtmvlgAaJiYwW0kZUndM105KfQRSIOxIqmiaYHzZWKRh3OlwViza4oBcpDx
ZIqNeM9F7XxomJuuIWPBFfPNhdnXTVg/aUnvX0PTXwLWA2Vic3vAkuSLKUoMRxhz
iEioezHa8MW0Am+e/qH2dxZdxKO8gaogQCxTAKrO/AXhoZ3x7iPmGAH9nLsCG0i7
tM6uWReBJY4SvKwowzgoDmN8XIyXoiaizhXLhFqqJ8qZ0BSpIq+Bz8OU+rn9tP5Z
gGcA5nEb2FlaQ6AQnWg6XHeGBsLfacY0uMCKGx85jCRNCykSuvYOa6n6FpsizSPB
sMWOL/DzSjqdquOaSBpnWA==
`protect END_PROTECTED
