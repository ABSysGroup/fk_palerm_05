`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uBnpiVNwZsiSlsyZIUWsIv1K9lH39uPX5ziuIfNmRVL14e9h5qpjYjpFpply5zMR
Q6GQ1Dw1ZN7kpNIApr0MBR4Ej4YS2z8P4JFA3q0SkKvZqslDpP/zjp00ai44uOjd
HbRWAnfzLXywxXhltSuEASWTSg4Z3NPr7pGPcEWbTYpoQ6jbWsWJjn4WoQWWGKfK
+OiEYOnEDbpTbUUhWdFhPytAqYMEfEn9ArPDyfZ3GJGThuNwBbtHVz50PV6elXew
n5dGuHxvdv9HcvKNXmUjC+PhqmBtSQd9kFCGGftQcSOyeW0ufKgo2ZCiIt6Q2LlB
iXZk0tyE5Y9g41WZrdsFUNHFwF0LIhn5qLL8KkTLJRo=
`protect END_PROTECTED
