`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mP7uDzRqiG0gY5al7x66NyjiZsox3WYYh+dZHNURjtVtxgBnMnQSdfawNvbCXiNs
RQnw4gCy9YcE8gnL3GbSfuVUEaxjqEiRKfO2RQcZronGIiNV3PEyRxjsa0rKvrKm
1f0STbpaVF28rMpKI+9pFSh7YlUT2qDhxETry7B9BaQkb9eXZ8gpQ8qD5qMHTwwA
tH3peOO0mj9VCSntrUxD222lULBftgWT2arGZYGE5niyWvngVU6+mZ8iQH2TwZaG
iT+RkrTS9L9ZUVSS1sBwoO8zDuwWTj3iYKlJG9Sua4bhv2t2ZbiSlMvw6xsu+MDj
rCY98oeLCwkyOtKn2fT6gFoAUi8znZDCGxN7IF5fQwNUzdz7XqBPDUQF1rsnNHQY
Phj7ZqP/OVxFFNnU+MWq6D//0vG3xnSFAui0MhblUO3vm2thbea5jR4Y2dWgdqc1
1+CZNebheIcZWd4BR5CM/JFrcwsE/vjHpRXZzEnTZkz9/zRxhK7Mr0EbS7+CoGDt
hLaJfDQSP+qbd6WlDGYbskHORMiSGXV2108+TJrEQt8BVzriE6WdH/KreLZOaZTg
dtnAQijC4/U/ilxlaUlLZw==
`protect END_PROTECTED
