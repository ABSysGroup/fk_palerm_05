`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OEAwZHC8dxPbgo3J8ApSfgg5sAFN9aMLoYeqaOZWmzih5L5QxotkFD6Uz6J+d2sM
FXnNbNSifCW/txmCN9Q4ophEYJjVxfhO+2BiR0JQc/WI+Cg1Db5Uadr70XIMnK5+
4+fQFvXlOnJrqR6/xdZyHJWynDpSe2u5I176Vd2kyDlNKhUQsmOlP9Axf4oDAG/2
wY7Zt9q6bYxQ2xt4Yx2UrdPbeY+Mvj2EvdILjIRP/QEJ5vFLD+Fbg2M8c0f3teJ2
bNsyH2v1yQz7BshXA14ioMFVNTmWB2QJO/PHjbGn65ITIXvx3qxVZuFGodY86VXg
G102p7aqac85x6Bgfg7Qc4ugeQhOsA5Nu9aS9A84LTs0DWc+P+CV4tvyZignDFjt
NDvSkz6PSX1Zd+t5QUIG+Q==
`protect END_PROTECTED
