`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Evz5EbrtEnFQG/lku6mOrRJtg/RVC70OXhZ2dzRMCZTbNHsacdVop1vSH2fFCqmA
QYpMEQTLoqvhR8+hL3aoKAVpEVaxR2sZwqXtKRqL7c1JURmISYOsQgKomTQ/3FE/
zk0yANMHEjXJiEaJ09GYoGXsFaMu9mF1ZBQ9/g7bFjLyOjQfdSMPBdcKQ7zBt31Q
eAMubmuFnFXiRgf6S42S4SzA7N3edJN7vnEM8//0js2+UqM8+FsvYmaq7HLqTz8N
shb9x5WrKEPE3/gGwrHaMee7OYBpMAyutzeuWathYwA9MXi0slNQ9iQLs350sRTn
uw8grXJpDrH2xT4lOleELzhhfVqQ6UJ6Qox7hlS01oVqYPmSuvnHUmmqB/jPYcHq
uPFzR5Mo/5tdRokK62+YyAUVS7zu0dAZSZaFDI9rn4/WoxM0wt5Ub7kEhyM9cRap
2fSp7b9sYhPxCLkm3nfnve3lokjzH+pKmKFi/G/54JY=
`protect END_PROTECTED
