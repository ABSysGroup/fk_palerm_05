`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
06ZWR8eOQV4Di8kS+uXndUwbC6hADNCb2MH1e6Lg15tDZgxlSQM49eGfKjoxF5nC
VfikfK8eA2LBa8O0eTmkhcwp77LTRm5tSARUSouhIQqDmPDz00TcZctTJjCp83GZ
w808GSueKR0e/TJCfgh6nLxzrDBdPUHmPUUdUzYMN9lWd2RdzNN/u5oCRA/yH4Sj
fpAKlkGHFA80BwpzBF3s6y+3vURQ1cCN4OaYxRwTvM3IU5RaZ/sdsqLjV4uoyyvZ
aON09CVhFx4KIgA57CTJKpvn/wpcczNmOQ+RvEBlKTk74YaXGM1jonjSc7iz2Aro
cGFOav3eNkiTsOjlE0qSHhsSIhVP6B5B+C8/OIFI/18q0t8iBF7njGppcHthwW1N
OAncleya4vCT4DdZon/Fg2PFCKaCg9MMgnpeyor9paY9ytbfRQWNef4HXbKGp9CE
xo/Sgm/5IFV8EY5WGnj/CNFeSLL0sJmexQ+iTzakp6AG5iwlSsRCgizqVJxg2N7e
I/anZ0GVXrpA5Kg4A6whzJyn/LIHKDNL/ZYB/ecr8Bn/FcmZO5AvC9eVC6pkJ49I
/iMmKK9JuyjleplTe/EwTw==
`protect END_PROTECTED
