`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6FJtzq979atz9LshM2zS1po2CAeTvli+wYCJd8oPUoEolUPtpqyqHDxHhXJXKuhR
oKXibzIXIihc8wzrYRoE6sG2ho3+6uE3fs1VBgI/f/Ksv/edBsCOXAH9yxMaHyYR
7uTm7Dt4Evv1x7gBwpi1FpZ4i8NUoNbx2jENXBSwEuc28hLU1Pq+0X+tF5CGV76u
+dIt6xBm0z6Mg0DAsJQuJM2ZbYJgPPZnl22PXH3ZVzlmd0q5IaW5QrJCFUblas9O
lSochPAYL3aFfHFBT4MaFvBPJQwBN3azv+QbYjVaB6EaQFs3ThPlWzE0oJiHtW9d
uHnhmgKFgCct3Lh9dMUE/JztoCUV2CjDAITK31GjbBB3Zpg7lAEXjKV0wUygIwAT
L2UEHwCBCzsFbFHgb2TY7n9SlpLUFAqY1eWGwlVwk0XDK03pKAPRSJOzjwD7xsQu
MI+3Rd9ML91RnvcSXTiTTmn3S6Cv0uJl3YvKV08oJw4RrX1UCks383nd1T5CPG/X
7HGTNsSnKoO/G2olkhro9b24mmTelGItxnBg62eKlQATK7jP7oIDt5IWM9ei9UYV
hT4kHkoDoEI/kUhHj+To0yi6+rArfhjIX3zTqyHgY4LVna4kjNlooIngsh1CLyfS
CGPYl7hCP+QjD5IP8mBLvTIlMgdyTOuvZRcn/+/wJFM=
`protect END_PROTECTED
