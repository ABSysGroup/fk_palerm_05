`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YKEJT2cWQ0JG810Z59cYeL9GZ56wV82AAPpQhB5XqiP2CRYGjF0Kx7WIUk2BL7MK
UfOX1IHaFp+RwPttKnEFeGDqcMCkgNGMrUVvvP8xa/IBrlT5O6GfFt4W+qUPkrsP
jIEk+xoT280xV4QVvjY+F+WEIVlhChucWRR2H1tv1GwTPxjlD5HgtE+NOBVAYrun
sfkhd/HLOIm2fYzDghzZLcpS8axahfI6n4OWHQNQ0Hnev/HQQ/gXeD81khdiHCwZ
eQEXXui/K0GwnThm0xLN1Cfdltyxht2ge8s874Oe1xe8iCpH6se50oCGz3TOJ5o1
WY4bGHqnqllccYsFzQM1c2/KHy5qWoACIatkIWCK/En0WdGALcMbUzI6KQ9jP8VS
3TnK4AJtwPo3W3rqDU2mm3aFElZWaTx4lyDwq+l8TXn3mYlzzfgmBWuJMFjJ4Ucq
0AnR5vI8KjKhkP1PI/JV++Pk+rkiBhjU1r3kwItwDFdk5N0/PpmjzK9gqHHHOPcM
tcNO299dECX+CSkQdUPJcuHWrA0cub+zDTZgT82UeHEax+91FMQ839vRf5p3uckI
K3NRXNq5nAG0Yns+T3IXvr25fMKYlzBxkF805zTx/oPl5YTXKWAVkKldsvqmKjwW
eN4enA0vfdk8WkqlELQUnLnpUJQEBtHYDZ8DXBgJPggTD8ND7X/oplHZuBWqYh1J
KxDxWQAJ81ySuyQ7De1RCA==
`protect END_PROTECTED
