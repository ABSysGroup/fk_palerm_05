`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HxGlJkQE7Yu1vUienrYKJ6BevfowjddrmVKWsk9+8DbfrIHGGOmMUCGVotQVnz/m
fOu83i1nVHGJF+ahf9T8Z5G5MTK83THgkAzC62sfXYVUpbVdHInPku/orGtefzWv
orJS9d4o86oY4zNRoCtACBRYCOvqzXvaGI08djtwDxZBow26L5CGoo39YbRCVrgE
CPAIYnyF2DWKEoY39pULbnJG2tGOuzH9Q47XJIv2oz8nCa3xPvNRBhaPw4o3xe8h
kB0i+UccIAUlV290Ca//PZ/mRz3eHHKfzYyrNjf88+ADkw82+eVEJlLdSESGRWSY
8/yfUDkbIVy94P7Achh3RddKHe+GqANmzvQ8DxqQ/7HbPwtJfjBydWKx/8byo8zM
4dSnp4JZDLADb9YkjSZD1wb9d4RuZCEOok8jBU7bKAsMAw1ovbxn7uAC+uukoS8b
35XIhVjsUMj2C+GnVy8bZh8ScdSm+w+AmIEJcnziQIyywOXzaSp5NVKm/GEM+FVF
zapg9hTA/cvvFOwp5Bqae/THSDpxQ81fTX6bZDxiyw/V4NGoTXEz7tKlBBd+PYrj
XAnMX7HcXNsydfGvFPs9IlJ8OnxixgWUKdgLmL6rnVKB4uQePf+FFLt4GrXzzm2P
n19F9Yku1CTSVR67STJaAg==
`protect END_PROTECTED
