`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z7g6hnlmJ4iMZUFvA2Nd5BlhWPOOQKoPbcooVnsMUiKQPjw2CI+gK2lQmmec10VV
hYtkBSD7bJZBW77f+FQcXytURDGhmtty9/SNwJfUJd+lcJukQ+bj9FKwSwvf1vy8
yXbv+IEQ19UV41FpfhZqU2KHPyq9tnqw4zqBsBCWOjAD2dzr25AO547RaK4Q5Hzs
by8FZNxOPu1l3zc1YX6EJYvLdreJUUSQ+kQ6w9AWFhAFztH3lwrd61PBBp6NnCGX
KEjWEM4FTNp9drU+9lmshKcbXCYmvE1PybRGRPb0UnIFeERdxnYAkiaq4XMtZYyz
cimu3by0/lYbffih1pe/UDaNC+JoyrYfXTyqeokS6tDh3rcK2SQSVDbhoXqfpEi3
QgL+zDcSN8JBmqBa4HtltAluQTNpK8EmqYWskFczVer6XZOPwzS8aHhohlrX73xl
Y+UvYbKjLFrodJEAVIaXoDH2Aip3axeBBhjPBbkj0XwDMqV1s5oFjDUPQXKsi0NZ
pCiNnScMUtiRpa5y72ZVf6JBJEJtakJotShrmetLRpIAkcOsu2WD770+HRqYYwHK
EYFcDMM702HmsL3mk99+P3H1D622Fk+IEyPcbpzqoLujuS9aSLtd+lsb/umpHxb4
wPDdc1F4lTfdy5Y0b1Htho8pZYiQMkshJNIWAK3enSLbwKQgtiA2gco2mtnQgrX7
n2+7jhMtWgsPi6WyUXNfqOpHruRhgaR4jOlptkEei9UveP3CSIyFzX5lI9Ebe92Z
LXgQ84tB+8YxKE2ZBaQAcT403YsI6FZHkEUohUgPp8Wuf9juEdoOMwTfME9+zeJA
mV5JT8bZGfCHiA1XJAYyaZThTEjYyM5MhGO35BWju1elx3quyck4QKr2fSzzDr14
yAnwE92seSyWjzAQmdURgqp0D5CfXkTajBFHczJ/sGzSHNs9H0IPUz0S3QKK4nfP
gbEAnJE9AhoBtpbce6UGFfBUWp0LHVNTu4+cKzEDhPvkDrgJAAAIldAMOWZVoimy
Q7D8IDeawLskvLbVM6yjH82o3ePI+P8QL0QpaI/7nF9gwEcHf2AtzrRq0cs6kQkL
VBySfvjk8OzrsnAsKF/Z3lEiFhq7xVQPpGZHUo5sE/LWIErADXm5kFnhl8ZpM3az
HePbw/iyIrcNaHc/Iv7r0j6PcEVbguvZcR44DwL6nwtL1Cpy/s9ZtN6OHyYOVZ3G
HN6pTv1DcBmOlds4hK+8+wzchAGWbV2+Aqbh6/hHijqPHvDn6u5hvR9r+2+E7Lmz
qkYNU9n38j3n2ki/VuDybH2M3GVsVTmYfailoHk4FowFH0Z+sWogi1IixaDs09mk
NRP6fc9EK91iFWmBYTHIFeVlfy5mLrux6Sqg+oreSLg4fgWJN4OEr07PRTYO6R27
cf52RUvBrLbQB3w91NxMth+kxzb/Oe4EZrlj/jJ8ELsMFYxH2K6mKxA801Yc5WML
+ybmycuUwpWpWwpzexlAl7uRnGOZbDsbA7jwGlIIejN5CCf9OMIMp7sXymgUm1hC
KTR++lWY3zoBhjHAqUsHAamnS6soojaj6PMuEIUxP7SFZLvrAIVl5vnbHIX7gOFS
apyQ5gCxd6VJb2xfsjOPODdHGYQk1b2j5X/TYqTWDFIFRoQM+EZMSnIvm40uJteL
Lf9QXyyUJ7Q3xZ/pxlTZAcPmDgvl773MDiW+fLN7YdB4AG1KSzZwXEoIVZvuCv+s
dIW36flJ6/Xauok9GUFvfSn4Gmqvdz8i4uniPyevzAIEmia8UUMyDwCkm38P76/M
85Weu095AneO6g0p1afoonEFq0x5A9lIwnf4Je5sVCd+PY6dpMf6lq8ZcUbGoQ1B
Ze5kPe3d7HbuS2KqNLfYUFsHcVi42OuZIkaCOj2x3kjMF9pjsjcMWyUQ3lVJJdtu
pK2nKpti32mUXrh77SfNmXaBHHu/MTy95Ew6BDK4DID/cfwx6C7Rw1L1jGHg/jBJ
erw3ET3Ut47VfJ19Mtvaj4s9t+dwwdcezSAljeu+yTLr5bmp6WXzxABzc8WXc1uc
cOLbrGIMPMhi7QYvU91hM4noNswv8xly/C+W2nBaKPK3Ul0362dMxADlo+DWyeae
TxBtqQFHUYxYUnPoiFOnXBMrpetZIquUb2SAVBkaMQ3T6q5LTsTKqiargbCYmWwd
Wvfc5aJc+HbdQBYlWoUuI1qINDYsI2JVx+//gLFVUCGiXA1qti7q82Ou8Gah5NH1
TZ+R4NghT6T0Gkqh3/g59HKm+Xq99a2HdT4dIzGiZVRjH1b0JEbY8KBFl/ornl8X
`protect END_PROTECTED
