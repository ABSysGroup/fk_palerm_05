`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L/aArDUfGryLct1t99plQmVts+jl1/lsgh+zQRygW5R9YZuxz69hJMT7MfMvHK+2
fSSB9AYiICvv0+e55Mdg1jU0bQV5v6PGr1uVKXXqqUPAVhzBnVaCe9LNM7QOuaFE
KjTZnpbg9T+HF1PF45NKK0lSDVRu/iSjHs8hnxM5ctaB812j3vk3r7of6V+2zd/R
ol2X7tZ/oN2Qs+jUijTws3VNMUVgMnEkTurBVPX3oMnO1/qUnoEdQTgpeVkyTcDK
ahc9Wk6ihAzwSdOD8WEXzPEO8q6LJS+zXkPfYabPoNx8DhCSWxVOzMiol6lHPvnZ
WqV53LBFP0WLzmnXYK6+6thFisqGTLd17n+LvJtgE52FoTkZTQcN+5GE/1/CLxvf
7cJiGL862xT7p08WFMbf2PPUiDIEslxYnSt4iY2HXZpT/us7RotzLsp+LrnJhpQG
XyG3LpF3jSs+cMXz3xDEUw==
`protect END_PROTECTED
