`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E4dBFjk2/PyZHe+L+XDytsFSDRxLIdW9BhrWgCWLyP8JX9MzFDl88eBm2S5zHr+l
gAp2XfBBknIzATrxL/Zfw1cya9IRWZg4AJ7HWCvG+a7E02ldzcgUbFn4zUp0vv0p
ehzYea2dXa9W612PGqalD0Rd/7RovYnP9RiCInMq2AC5n5cEcxkwCDMIRZVhA9hA
JyjkiVS6TziLY1820rJmT1qPwGB/o2FfVUbBoD3KBq/64P1/mlXsgvPYoyJDEb6T
wEkwYMMqJen5OgfY/BlU0Lhgv3unCdELT05wNQ8gxF5X14G0YgIWiINZR73pfKeo
MAdXOMziwY4wHTOamQbElarXA3+klKRsXjIPX9AMWHaBgd7U52Oxak4VW/WlcXjx
YvEaSKHRuelPGZOiOW04UlN7dwO7r0FkFYU5CpFBRRwEmVAq3ZkDtcmtG/u6mAtg
CES3GIEDknVxL3nrQzVNxpuXQ/tnF9SclllgUfHSAUPRrb/LcMJ+ACutpmyKJdyp
soep6ChR8nUB76crJjkBb3ZoMAgvXAkswYwEfEEwqEMTBjxClKF/47Nv338bR8R/
IrtHEwj0RvXwBy8jfSwyULsBIx2tpeRBxznFLcenJjIsCMFocTVMmfMb5aVzDrMC
kXR3xJG5flbWoA8TFrHg6NhHCWwAZDtmrmTbTAAr/4zQxgPg85o8Ls8qqkTO2E7i
CPQ2MmeTogXSWm1/kiiWl+lI1RFw+jI2Sxa7D8g+Tmq2cC4JyNYISi6NJUdHgnal
8L9MJ8jflwHq8XrH/V3mLJIUHtoYD0gLdmh1GaZQQmhOH8Eq+SF7EF0piqk3qm7q
5zgcJ8uwX3vRE0K4hlyPdWfkq/NypGV8kGfjvZa4vX4ZiQMyDxe2ug0Q1Kmr5rFF
UYNmT/ZATb8GjOqm9qLUUmDpi/BOUW+p+pG74dErux4yuowvgD+85hfONDFYRfF8
KMvzkmclyssroWhZOwyza0SVLS3fh/I2yYegfyz3JN9nYpvxzdF/h+cu4MXnA524
qOlgwqhFToNfV8X4a8xibYHrKOT2XBMVtT+GOFSLTpvXj0ILGAiEbd19QgB2/U72
cRV6aFQF5y7Hx0D2nAksMD4iMRxeVJfKPt7ks2PwLZef9Ji8TrHbwUor3qIHVXd/
m4iWP0qhgg9a7HtO82HVMM4/ZNjbC2Eku819yPo1kH+U68OgO2hXsnyVZyxnpuGf
RMaN4YytD/iZDCnnpiv1JVHfr4yCcG/8x46m+qp5rm7VdWBfkgBW+cD+ImNu8Iak
/QzdKu/JD5juAZ0uss7j1LLt2qaT3fnJnwgCvqAzTCzMWY2esp1RFOlxv+UlmUXw
MZ5tcmCLqTdICX7EoxXkKOK55SthL83yhMg2rm3i5wI7rmXHtvHAVS114dNa7Nky
AKUJ8wvlI5cql1OvJhxbDCMy2Esq3KZ7ifzP/gp5icFSOj8GMVub/jhfrQZvl7QN
15u3nnRKJToAg7uqv9dFJWnWk2szg43PRuECuI95CCg=
`protect END_PROTECTED
