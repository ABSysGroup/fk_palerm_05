`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WHDmHS7l5q0jviL0tVG8czWrvzOfQKDjAmLQxFyDMFWTYSUManCpZs6/aCDi4eVc
yn31D0O+hYAvad5PjEFZXQg/AMSm8a3yXVz1zywkXJNjHyz/ZErXyZwukIf8wqJ7
ZMcDY6tRp3ln6PA+PYLWzkunjthR1tLE45UkZ/UmJuTmua8t6rn/jrjPQDeVG/Q4
80t+3VFUj4XFWRyIA7MUe7bJ3EUXCD9qDEGdWRotLR3v9UlyKJx8kc1M6XDQnmlR
lnVImYfXLoPuvG8ZKh7bUnuMur0QEdwi+qcFd+mhAYbS4PxgrSsYZwDTd2Fo+Mdz
4KusvYxJi+afH7qpDTHp5jDzGdq8PFUwCDWG2ReAoaFZOsTj50RPjHx/FtB62dDy
YQaKo5Ja6voB2+N5TluyJkTbISpJUA8fu8fsBz1LN6k2ZxFZ406tm2myogyh2b32
E0quUxSkiff7fO/ef9XDQnlorUxCwlaW0nuVGobfsO7y4rEZSwl6Qp5zU07qE6lo
`protect END_PROTECTED
