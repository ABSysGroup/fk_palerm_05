`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cqW8UgeM64Yd8fpV9V7e48R4+PjD3O94sug1xlnnEALUc0xVn2+BMqHVxefWIthE
7NmUFkBd9XixKJLjUDVqeUz2aEjeIkIkMTXd9s02DzNb0Gigf+3UEtLOzNg38I4l
2DoMffJ8Vyk8OyTY8lfIH6wOELsYlkG/nwzuVTsEzRiGaY8Ix/uMpS9O1sygAtR2
GQcvPPudnbsy6ZGeBW6HNZ9F9HNSZKGNqOH1UP0qcJNGxnWyZbUDC4LCyIbc1eDj
umBKVxiUtUPNIbZuk8tUWsie1fFb52SlyAFOxvf9cGh8xsrB/vi6dz0kpsp7xu0T
ovqMCQNuVWNfh84BYqe1+4ppaZqOd22ibs0pOjcZkevM5ox34DzqPyp6K6o3N+s/
I8JWO968jKZgO1m0DEryLXY62Qzulbf8Bsvzas37fcTpOtwWcaqGMOImBnyidC3J
q0uP8L9DM/dWFXHpVpFzVP5qxrLHcXkctta7N2nrHUO0NMdMSql/scdBrABKSZPE
iz2WQZPs0LBqImTj56LQbzANIZXF+eNNC0CxCyg6OHM7nutSki3VJ8tN6DRySowm
3ohK4We7CZP34L2kXyxRHfzcLo+bF+jy76lxsMiJpg6XDQncwf0EScrllBYdQLCx
+Mf8/u+46YpMb3ksJFL8slQM6ftfs8s4m40WVFTNHSM=
`protect END_PROTECTED
