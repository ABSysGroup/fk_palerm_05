`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fQGSRpvkQ3pHSnbCMi/QfIPeXKnDrIq7Bc2jfLCpJNBWq7+RyiywY8n2FssCavcY
CmAcxBYP3AqEPKu7bn2Z/L9b0e+R56mCY6T+nEH4ysFmI6v2P424s0bL2VASa0Qz
hAXYJXp8hA7EKtR3lkNhIGg+HW2Gnw1mXDRmBKuvsFFI49Hn8irEUBWtrPKSUVRR
m06k3aEhwO9mfydpGRyUJoK3ihU5yYkBfH19aYkGN+pRXiY3WypRQ+1preKDBS44
SpvCanNtG5cYBeyXnMLmcpwTCYvJjiTLyk/+nHTXnrCAppA55Quk+7RtjyYKhXvE
wyEdiDyaUsR8v7n8hKD42jb6yqTqHOWbpcIY1i8iWbUZFUCpM0zRHKDh1Klhp6BY
G9w+xb2IP4Uq3M/sUdGBuRDkBOVxg8KhuPXR1CD7XxcTca/2CuAOSMzXOJBfDuYW
1h4pfELB3JJ7zluTlW3tXMSAZc21UtzJoZxMs8lmfPWKIay2cYVwLu9y5VVTI2k0
qOn0tbmzXr2Gpxs4a8ijQ64jmqAa8vNXCy4pXTf+JTG1e3ZTOq4S7UoosDC1JHpB
rR6a+VDcU8lX64UOmA7Bbp7HemY0KMDJFO7HAb3EZmb4yl/KYjykhi1kuouG+uNN
ZConemM5LIgSRe9YGqz6KK1EWQdWzglpxMsu7UaOclbEXgO+IJ/9Z2vJXgVHkARJ
wULZpwD/DG8kUknD4Y3GOg==
`protect END_PROTECTED
