`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qaSHAvcMligXP11UsgRvXQRqtkOFo9R8JA22xGnqAZe2D7zSgw/GDaLccxTWWLc+
MdBwYBppd1OuvzMQch4Bze9dVbAmFn8AOuGK3Yak8HE2ogMwWOk4QFNQIW8ztfWU
W8AOGHQsn87cUO4sm81QHlOFF4jFNkdWOfIWhpU5ay6/9GRQpIBN0H0mnoqf4spD
sRvjJjIeGVzb0zQF0hudzmq+cY4fJoLNX3/rrW4tWdsMMYSq+tkkEQyfT/GT4icy
JtLEeMqqcr4F0r+bnzUuUMCaIdTmIc2ltvf/b81Yjm9JRe3/csSBAdT53Pd1s/Im
rioeL2rWEYdC12Do7rpMICkbF5GeWNcYD0d/uYc0ZxcBILEEj7zMBrPtxvL+/om2
cgpd8V7OaPlSysHI3pbmj9ADdeJp06benc5ZYIbgCCU=
`protect END_PROTECTED
