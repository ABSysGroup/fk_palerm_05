`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xLGFwmx3nXkAAbjBbxPgJAj62lUnjDYX8ipZ4qRNUBlH3jBde1+NqwJTwrVSgyHa
OU82p1FXlajTWcuoiaSszbX34AK+T/x2d1Wa+FufCe2udnvl0QPQZuCKbae7nib9
9rJ8acBJpWT1or7FCbepbeKtnahgBxBSUeihhHBm1SPkWafUljKh2/Y2tTKJzy5V
bFiQHL9q6HjSNz56Ja3FsIkcQUnHjSQEILKgazIVuic/nUMfu8AW4XZP5Can7UII
IzcWmKniBLETCKe7Bl4HPHX4xNR6gLg/0OHq7qqYh9mf3aVA0BvVpiKiisIata03
36bgjzE9xDhOoUuSaegWCXGh9HPRHApJ0E1UFAtWz2Omga2X46WOzSOqS3U3khnc
cIqymKqPt8wXAH4LeRTnqZmjiU/2gQ8y6MD762B4n0eHFEFnUTWZVtqWX2dTEYiW
JsfP6dzcvKEpTlKWm3Tl0DBegjwN9jZq3mAqNmM1XYz+RTqW9QoZ3CebZZP0fX7E
NnOdvT28usNOzy03Jx+L1m7yLWLi1V4kLYuTHe/KYCovFa0jdSWD2rEk0EzeLsx+
Lm0Q6si9xvNZT5ol7aXqKF86h2d3Nisnr3XlVcy1oLi/e07Cg0uT3OpXP5hoTel2
IuAKG7J/tNLQd0Wlzb8es1XeY1Eb+BZNR564r93e7KDOELZu7KJAmR5tFxKtmKMj
MIcO0tS5yk4Bt4nE2yLlha49Yf4JcVi6vq87HR9KYb4CJ7TtI/3IP0E+VmjAoIOs
AHKIr/4VCyloVGBks0+TUsftBzlroABOazdatacvFlkmlEtf5XbCWllnzv1lw6hc
cgVZG2/qJyAroYj87pk0tlQKuWiYxsZRlWzFjAbuzTC6hjlrQDjI/u4O4TlxF+Ef
pTsLZR3DKa6gZJDQ0Actu3zyp6deJ18XbzllgCjGc52cUmgY8d3w6iqDaYuMlGgq
1y8u+vv/nhLNwWskf369ays7+fj5v53xjQZP9M6oA8kJwyVJ63xxl8Yef7D0V3Jp
s6fjKt8PwKcl+g+S3CA3mG9I3YatH/GB1ygzKCbXV2dSBHvwvchOj3MQutkvGrIg
Ct8vMCCLuDqugSwO/2T31qKXNgzU8MM269BrpH2OMtGbLBdszewnsGYUEfZjGCOk
wQtl5Rrz2y4I5i3tkMFw29HaCIrqXr1guo0+5357PXZEx6v1YG/eQxh0bN78xSn8
FTrU1PU//OLwJYituaVRjwpb/oQ6rQ0mRLKyK9L4OC+uo5Ac+49KekfN93sCTLmq
HcsecUKgbeAiTUGFSz3M9V5X9gVXt612b+qft7JS40hDZn+vpfZbSCk+KWxQk0Fx
Xy8Dx8VONN1kXrjOxsghp+XvZlPa9RCdSr73N+mQU5/k9kS+wXn00mWDoTCpaRa8
Jh/Do8SpKFEG2IYB5JGed2Vs6jK4g8k5fkYZB30GZLtKJW8wArdyAqzHoCUcHK10
tbU0Tif8Lu0USVFRCTjWTQ10wdlvaURuq5yMl1kZokZOhT/OxhvI673pUnpT0EJh
iDDa+cg4fy1VeAbSuWEqRCWW54vM/H8/IoXaFD8Nd5Ha9T5cMn+iCl9Q38K4NCjU
euVLWXenVAQzL3HE9mWfV2Q406bMXIsmXBSD3WBnyKUrUCe8mR6+yOdY9xhEmFwc
sqRefZYncfz44WQjGHLc/avJUfdsaUujgnaMzQDOv8Sw8O/4oGOViXkVPyWtR9b9
WVewI/OwAuaRIaJqsXg90xfoXj2gTDMLmfD8PRzAPiVK09UdemPFAcIyYSC8cJWY
UbylqdoUWBv7gv23gzPrwBICKFXQhoghjjqtznMA721pgG3bPx9gmhRjSmO1m5QE
cLxOha22YBMXgfcJ/5ttCLogvbT8j64U6tc00t8oT0FDOqMZ+WFJi3hpqODqkCLx
XIW8gjrDADE6rE7uM7h8s3pxs2V0+IWsD6Sr9Fr6i+l4gPfgIVH5fE/DLqlEStOK
6C/ykW3IRbegXmdfcn7FZ6easumE6pnT3wXLtVh2YdGrXL8ngWZMDBOdW8ri66ok
DqEc6poQi00KLHyz0dCSVHeeC4syAZ+si4bit6W+fD/tmJ7EsRcxoBSP4Fxi2xwQ
UyXTBJGBm4eyJiESTwz7UKr3sx1TM2Rgdv0+LUzMbO3rs8CInSo2RdlNkkVi/3tw
eziJdWbDC9iJdrssdyVZ49i7ypKSogrUeFUzm8UtX4rfc5yQghmPUlZ6jl6TAMox
gJ0K+uRKdEWw+IEZ64+yO1LICDulJ9iKpJ1crzfg2YAti3jDmcP5Ko9z94ddD4Cx
hQf4VQTEXxwPWKc0wNoH/8w3zM2UczF3O5s35x6ePF1v9+Ao6AvOHq79Cnpogp3d
6WAOKcRgZH5m7bcYpI6Eiv1+NojA+3y8B9bndl0Scu9SAxVct38ehdgZsIL1x/9p
U2LphUTUifIENLavn577It5XorzWkJMOVdO/+qXkI44YzkHd1t9oKyGB7d5k7nq9
kIRz8OWtazrWSKnbJod8hyJEg9W/l/ML12QdUTLvrrn4M4N0aWyANKXGhhoVGos6
lJLfZfd95lIhXIAAhabLT0/yQqkRnY5hY4ric9mojmVaxIktib/G1wGPVIP7t9a9
iOu93ymwlObUDcaOCfRhbh30Yk2HGJsR4Vtktme6KfWc6nlWRtMOnCHC7UYC7bAB
U/hooFCVdGgZNADF7OJFNINm52Pc4PX4xdgKy02fUboUdvyUrxyE5QVbpHdHjb6d
Rj9YafwhCEb5vBtV93CdeWBllxl4lSE1M6MmS/u9wr/ivvMjwsMpGb/WdLApXJz+
2rRrctzY4VLyIbbmwoX9PdKB5NcY6myR8Qk9ojHZJ6S5KO6+81aHKIO+EPhBC1Pw
pJ1vVDJHmUFpfqPzR2X30xDmSdSpE8a+XdcCrQe8DeDQ06s2jhpiTLa8HRbADr7r
x0xdTKjVUfBSNYVa2TGbmxMPIRrP75c/Z6VlFTN8exD+w1BfAZRXtw/GQx5bg+47
4P4fuLuzf1ChIVqnjJhwTQs54N9XwS1BJS0z1OscLAneO2hra3vc6Z64WxCU2Wsg
BK5SMmQGhfws+h2Y7M4gkmZAeJtqKifLQ97kRC79+0dJ8/9IoyWzFXZ9rtt1Or5J
UGKx5sWcx4e/wIoL/YI+PrRmqU1vtk4Rqu4EtMgicNtNPzTY40/mdAQFgIijHen5
cJuflYBTzCmFZwLrGVhvMNGW0GeDBNN56c81+g+e5e6/4EcQVDLBxSsZrhFH9qWQ
j32XD+TJuNY26BiSWuAIdigC2rTmaZzv/FQb8iejm8dgMaBPqkA6Ju3izv4HfE5z
UJYHBSUkxFHNAXsdqzE/A7Q/YRFdMsByvKmJCHBOoLe9xD7lW7KnAVJmjxVfxz8J
TKDpD+1/d37wVhdS8191S1EBU19Tpm8/OXV/uDR6Lez211l/FmocbBG9kKn2yUyK
3Vs8Ey2UyGGsm/bzcN0VG15Hfe6PBOUJERFm07VTkP6/Pwr4jLSodDjWJjODI44U
YhyyVhZu4SYe6jozT8V+RVDFRc3OCNCOWAiC2pwdOhgC6i4eu6dBBDtEiDG9dQOj
xvSI/3sE+e5hAVL/2MMVYSWxE7KE+psyCKZ7J/ticFMy/5q1Ik8wbUTzMXzRjpsm
VXTwTREe9WFOTSIoETPUhnAC6PU2jMpOKJsS2gd4D9qvqmGOtu7kbL3qyVM3yvRt
lghqFKbrntbLpD8GCKio3wgM5m0VZUgI5JMcvqO4OmnexUtCgtdrt++KY2MnUNT8
MZJ8FSVuGOt0a0Eyb48qe8TwHh55wTtydee/tTTVHk672UQb09WGm2lkYwShCu0W
AVNtyZ4o4rQmsuUdXvI2AvTTAMwOqL8mmuqWCDsXYp8lR6WY7u0m5z7a3UeyE3dh
z4pSjmT7DlK2vqxTam49HbaeDIhbcLdYu6ZmvZxOUSyLuqGS9qkr4q8zw5X8napp
v5OUIp643YTNuFtAYxo6S+VSeQeZChYQYIR0uLjpMhBntj8x6kRkuqngmN9VxLnS
FHWOUVDxkxzgoX57ochxWltEvwpInsMvF0Ob/xEBMCbMVSSrmap2j+oKCM3ao3OX
MXHYJMjPc5mTbCg3Nnljy1AfRDCR8M3t/gvPKpnuowmy8VCqBp8HpQ5c6eJsJp7V
QYhzDTzm5cW+oDwGlKeKEiQqL+iDc5aPBUEI817EzO2EflJOfp4Sn5/dt6RllM4o
vZGR/XkMvULZcG6tjLerqGjw9AhrfWaWJrG8P2Eubz/MpiaI9vykvX9hjH+kXJA4
9IWGOeNGbMToh3lAU6/FbXegeyT0UQcJMMC/qPB0xzr0U844p4FGtVWCX8JNNnF7
6pqQ2K8cniB9+6DTzZESJ7Gj0wzmmIcLWmZuJEm3paiMcTVQRJYQOEr4YLBCWCx3
psKUosnaWEbOmS7WtFcJehTXD67CMPafjsijSVh+BWPkKr+8Xmbk3uRTCeJW5XU5
Og/4CsbPsIMfjsg39YiIc6DFq466Hl47et98TI/DCAyl5OcsmzFbaatKislUH+TG
rph86RZD+Y9EWDQeDg8d2LYYvQmmp7+ERamMbK5l2LL5EkQ2s2tRVEEdf4HSZq+q
Nl3QQxHehabqFMZdGKpru0Oks84SM5j03AHOZ3R09pjgXf2uKVXEYPc76stS8j5+
MAAijKshFzdyAwHppDkooIVO2geTKbeR3S97rnHziymU+wIrYJ95mX15tPTtHwcj
ie42cvLoaoelUYcuR4hk9gMvSD8NTOskpTzs3l+UAk4tZoYvYpbXDuaC3JMQO5w4
pU2Po8Gh7spHukC3hqjBGKPKFtptb+r2dEhFvlwKYIZ2JRtiSsaPDcFn3hapklBv
Fmi2hrO7MXzbMfhL29fmDwKWSPMkr0PbyRPGWD1Iz5I3PbzyYInNZc+P/3xCm9WT
KE37OW9uy8I78zcT4S2+4XFY8Mwwd9mtD/ll4MRg5tFAZo9nyqFUPFCUqdGT+GJD
70Q6E3RaksljmApESt4rNVYooWQYvmT5TrhM4yypDCQt3i0laSlGSFdTFLgUo08Q
OLYr/AJE9nJbD6B+E0zPkw==
`protect END_PROTECTED
