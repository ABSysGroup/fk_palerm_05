`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rxg5IQvL1mArIKDOer5aoTFb8z0Z+ZjBRi6cOpT4HvHrONibj9LB2uyFtBLf1LRx
9LVav74zMyze/fxC5dbBaxQdwtJlQhIrlnPVShe54XvTq8ICyoHpY3R0DZyX3F4R
p+wfXGvSZrKieq+ggRumDdTPkxhADAUppzYH28MxCLOZ9e2zIggWFIKcDBSr8otY
dIFdYQyPAKACjDTHYP+Ai7p+FeuLX3OWirDW0f7lS2znO/iwmXn/3oUMdaYlomtP
FF9h9ak5ZuvBDGFhv37riJi/0JIHbfG97XJ9GX1KUcyR808Cd4EynnIXd/5jOOIQ
0W7fwzvmPuCbMnvRDKf7wZj/7RXirIPmFbUjfjZf2+xzypkj275Q7azjOvwQwjrM
`protect END_PROTECTED
