`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
14k0WQvihLfgm6Et2+YRgg5wIUDAq9biohMywt5zrM4phAF68lyFv4TASDxsJw9A
P6JuppHAs8ZGOiqhWcIWEeg9QI5/XHJUp/Bw7nRdqutjNyl6pmq6+c7sfz2vbyTR
7XSwDnonUOR0Zca/PkBPeTzuoqYNeNL+mHw8bZgI7EwMk0OiuHLz5vW7P5JAhGOq
dMWudlEN+tDToFwWRWzL55ZSJtvkvp/sPfV76/MTwWGD4KQqAEiNi6YPJMMa+nWM
6leO+gHiacWlgm5GR/u4dPhhb1zqf2s55EEulTOBJYQbKf+q9P0XKOR33cuCFDeA
ouUMI2vl1RJ82jo1LfZ19V2O8+QIAN4ZMk/MgQR4Uwynsc5+NS7kJAcWyP7vP6Sg
j+gjyL0szP9Tk5Iz7Juhotqf1GmCHNZZQdom/BROjYqmCuYKQAlSCI4XOXzLpINr
k8es5jxB/n2FmiAR38ClBVGMMg+0HNliJjz548gtafOozb4qaL5y0+nJx5DDRLHK
CyH9sLc5MaHAiqGw0uBHmAfeO45qTrdEWj2xxuLTdXKBYeA0qM87aqaYm0IKF8+s
TJ2bUVqkXkCaLHafgXh03Mnv69B40PaujOIaNqbVq5e0bD3HH3j5FZhrNp6IqSpx
UZYbzeJP40v1HnYyA/LIBXJjL8MmTi8f59NLNfQ9VF2H5bgG3jdFK/f2Vdar1GST
UZKk3OCZA8aaw9LFyAQzJyj5m2BesiLt54vrdUpqaNdWSzuxD+UBvEdfxkl/Phsz
AvoVUGho+S3iyjIO+pm0H1H0gR6ZjdRMokp/SFKhCSaWeh4Vxkxt9ZsE7+yP9Qc5
VlQARQeFsXTySshjdroILNgCDMyIr88qBat/XjoVUzvMJTtK7UigQ7TC5ImvOq5r
HRXH5YvH2HIvRByxIJAZB7yj6X/kYlykqfhZn8B5IXBRr/eAIM4vo3+9dMMeUHLy
GHRkQV/h/KCpWDbMrwBPhei7dtp8I2/hKrpmtoLZip7Mf9Pe2BVg8/UiSAirt8/T
+I0bItpEH3YAU4wRtbGHLUrjy9bpFI3qYVp6nMjMMC/pn0WwzVXXaEYWuqkAFt57
T0KxVG50IO2hrC1NvdRZME37tqWHUh9QDRxojMMEfsUQSF0siC+jPmA8ogJ2ZARR
82Teg9/aQtgmlyZ0XVwvtUITpmddGaV4IUp+Ppxe0Ui7opRy3aJg2prWsdE3+bmX
QRazPclijNYiC+7vjsu5JTa3nb53xYau8YnO6eFJKDQsCrSITVNbrYKXESGDz77B
08yd4uCJnNZlMH/fSV3Edx0H636OqW/w4b1eNUE3O5sSV5JwW5Vk7DF5llGXNzpH
nAdpvc5Qk97p4lr8T31d+ikZwuwXc4T2Yloo92NlaSXzP27ZuhFOfkzBxFYFj/5s
TClkbLxcRIYGtnvZ0IRwXKlGLq4MSB2CisDic1HfYcTBr7V84g4wVB6/zIbXqyRL
Eo88zepbmQ1wiq4SYajuvh/l8AOc+ofc6oqCXvLolfAlKnykdNzCLTMqWNkxLeLx
gT1zoDRrjXww7jfZwy0vU9X9VJlhYh/dFyIEFB59QX6kh1FLE5mO/k0o71HjCVPY
CxXdHwdLjRaDcuBaLgbDQ6Ai0XbyCiTDR+GcxNOy7SyJYfwVJ7PeJlQR1Wc1YF9E
iGY4Nhutl1krlBpkbNOrJJ1IMK9Q1rFo+h08sOwERgJCgwrOcjZMW61ADKXiaxXA
7PiXqh37lK1cRsfwLmJNZa69sRx9y70Lnn6jimr8qSdSMUnvM2lhQf6iwb9vFwUL
Pik5mtNlUEkoTODQdf3V0gIeItQn4LAYc4dnEJwPabl7lISK6c5bBs2ztVzYFd/A
DCwKvoB9pVS4guSCQpPC4A1eNmDkMRh0G38BU2qlAllJ7BlgiEv7OmLUMspzBvr/
xim47V1hqA4VdZBx1RtZXgFNeYzxQHadGMgKj3lqs8CKxax0NgIQ9Jf15nhDIVYB
RHGo6IPWPlI23cEcQPYiFImbLDSw6wUxu+f2NHcAGZOzh56yTa/U9MN7XNdCX4ac
e9VnXShfAUNDSCw4s3f19t0RPyGSOxTBE8xusPVDD+pvOhlRoZCDqMo+gXkLcVr6
PBx6R7Sryk1bACax4aNvqZnDxvUtaJHmZyYNwv6y6M+mTRjifxyTqBHAUWERqz3I
WylNnfalGhMls1eVm7Ytx8WwGVIr3BLrlZjJKQM/3/96cyroD79ZE+Br/y1Zcj86
3N8WpavmZmbDWkOp1OHSBgbA4C65bNGDYmsOF6gmu3NmqdeIe14hoZWTHaHT1OIJ
BERhZT03TGeqvy8mm+2V9ImrWrd1ZAYm2pKnlSn0Lftm7Ai1RDUFWfoIkkuI3mIS
4Qr+gkI0cLj6qLsdeHSn7RoH5yUSydTz2lLefWFfua/fktVrmWUVSHwVscjvOoeb
FysmMTMCUpiuDXzZN7icRabVl1BDVX9YTaEDbdYq+IbNKBhUOFkktn9o9OqyLs5D
Q7FeYobjv9F9lshS07PuhH4EyF3XMXWllYICmnDTaJR42ccNKnuR+InkXKrIJ2tU
7TvKUPcVQ4CedMAk2L6LLtcLTuWwIdv0htR8FgfZJzOMunVeMmgLZeptg+4KfyFQ
WATkdIeZuQTO3Kkpu1BWL6H3lyhnYEUQ/KmHSRvD5ejGDDLZPOwnOulDcHnq2yZl
UeRCSa00nUm26FcpG7u9WmRPyHPjJq+CmCsN4zpZri96ouaIEUwo+Z0Ac0vEGgrP
yfB5oHmoEHJNhJSpDZ30qZS3u1NdCtNPR+suInSdKzrx+AzLvQSRLKXYE/wjTpMa
tSEvS7zE+Y0aG/5PRK2TaT0Fepojjktl2OcLpXhdNKeyCVpkf5SdKzgxf+i3yYCa
PVoRf3PSe8N/ExdYt+om76vgMD79ascuN3Hhux40HiHT9u3jSxEgfGPrTKQbr1vS
WlogZDMw+t0O/aw0efJsV3gszUMaiksT2zrsjZZWDkS+ZCl2cQar0X8lcZyjfKyV
3PqOsbbFCtyFToGFatV5NNTo4vLg61Gg9CvBUd4sQXcckylmSTFCwcJtvh8sRFH+
S/+5iw5LpRs18tAvlR7DEYqPn4UrANBrvysp+Ee1jB38Q/IzPdBNt1YufbPMhD+c
hPCZZavgfXW0YOwEsJD7UVHlJ46RqnloDYPd301IeEt1IX5FsBVaeOgUdNcf2S6Z
xdRB435vCMPjIu11fiDyiE4lE35cipKvnjm9ZHLcr6XqYFD4i6DutfRBYZdBWWHg
IOvaofNDENB0CprolIUUDYgwpAZSS92vAT4UVXz/jVVDzTK9b2xbW3jVe09AsVEu
rUAvNj0FZldDCtb20wKjkVDeH0+c9H5KOOGC0EZ+V2kQ2pxHm2JFeC/CJRQG+8ih
rLyJBnmv1x2QKXug5V+KoGpnkliTzhpDqR7KU4cBzcRi4WhKvhPlIUArAWWlq2FY
VOCPr9WYmZyXMhAfVJXotl4qTihJCFlyEAwGOgT+dqL2Ah/fNmDIdXuQAyw8eove
Rep5F7X71YBQxbWSNgLCby+btQ2NHppBHFPb4akxZlIJX/sgD6XN+++90ifaGMNi
r7oNq/zL9FHWkoMwCP33PyhbK5FWPzztklC0RLPy959DNUVpPn5zEmdXmYY9TpjW
/lGWdbftEOZiE1Sll1E5JbILbJnA6HhkQcFzMc/Q7oLBRqlK7u7366DU2C34j/AY
fXqRk3noSgt/svNf5M/RBMwe1/uPjtT+leuasEQU7dhpWXh2MRDBSLP9QxOWjmTe
siLd/TQCJ0UQQi834/r2cw==
`protect END_PROTECTED
