`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OwQCYuWf5uOvcvkCugHKnRPJ9oc1rPFogTHzHCB6FyLcXJrhbn24b6TY1qOcefno
aYRokl0gqYRL1zrEMdZhiNRq8ed4Q42IPtn4EuinAgqht7xQEkEibX+xtVbBo/8A
iFTVUBNPkerFDEH2Y0iLJlbJnpEvZHMula7L7p5mTK12FwKo+Zj8PB9iFBTat/WJ
LN9UYoVcoQoEggJkZeSntOfo/Zku9rvuPEFh818o1TJdNYqLVtD4uxFu+ni9w5qn
WuYPNuVp8zToAr5FeFuIAzEQc1YqWizEm6kCrpp4tCNVum3hIdXKjovH0WJ29WC9
vRv4IVUqiSwrdAldfgcJkA==
`protect END_PROTECTED
