`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OvK9KbPQTn7Nv/ixzDukPX6+fvpbedsottKNMi7RSqWdsoQ8lUfI63K211q0EAzp
vuDIA+y7/zRpMkglCzKwHrhn9YCCvZ7vitjMb5YtqcR63Ufu+B0d7O/G9KnmQWyk
uQSoNODjI7YmVpPhbhXTpkZSKsnjH9791ULQ8iZcczlMate2ZeOsb6P8a8zigxRO
Amn/V5SH2gAMxtz2JoycZA012pSwrOXDA815d4rLJAJCYaUeeLh67/hhWoup/5zy
fIitIuU57GSkPT97ihzxSMchCze9R0UFcc9jF8OlI1ds1Yl9HU38fI5RMwt6n5JD
eQvnvGifZDyzybArzsaipw==
`protect END_PROTECTED
