`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w0eJFYm92WxJq9O3KNgErSPmsQ2331sTF0+rkcjCQqWYQ9HVM6Hf5RgDyExPuhRp
a0um5mshw74niPpJlG54quWJSpSXCzIXApWBlhD2knucQtn77tWaFWoxGd7Cf3eM
ZWe6C/FsWcb4kMC7aVC7b5XazSGZfKIBLP71ReJzB6TNCi8jLaSkhx24G8sbrej+
Kxvzyx0eR5jl7AwslaGDY/QwYiRJj16sbGSMBvsPktEXsqXvAVaBT/MscnawVkob
eLhdEtqFP+86va1CZcBqAA==
`protect END_PROTECTED
