`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QnA5s+vXC6OygTO26dgURROh/VmdJL8Jc7XH24HhJ3zfGBgWGuRFR82cWy1NzbZG
B3s9yyheM8epGNqiR74wovifK6nLAZgwLGBmH28yL/nbN2mxa0xzX3OgU1f1hSD4
1+9KxuOHqbUv7fqS0W3gQTfC2FF9E+tBT8b5O313fLcba0Gdap+B6OxnOt0GzW85
Ys81JUMGhnWM7oM+Z4fYGPY+8O0cZkhB7+O3W25NBNRsE6NnSjQz9cVKtkw/cXAI
YHKKpTfCfAqQIj4TlcZl8+T51QsnBuE/HpnhpO/cLodnULTb8UhRCzQp1fi5s3v3
Mg5GhyXbYEq0DYAlStfabFEWVZulP/lwfir2JrlnpkU1a5i9aGvGYC09TJ6udBhf
jy13t5lGwQzK5nK0vY0ZMhVX6SWYmrzt9TfIop5HkBKEACXihQzptWbLJWHbmkFG
t53iGcTB4ODw0QZiyx/e8bvKWhdL6yOdYkql2y7+1fBK7YUrYA0RS/sXtMpuEn06
JZy3TbVoAWDev8qkOfNQRRLXJ7Xddwta40AUdCtqECrFVvWbwzgkhyvELkBYJ+cF
eGZ+pT39LxyetmROafcbTZzZWAqPNeJ9BYsoHcHGAUT/5C3mbbOae48U8Tyl6OB+
K3eaCK+F4Ob4UklkD7X2vG+keiA6Uj65o3bDM5R1xfCqh6023CSBRPE5Ca7Xu4Lv
cbPJo2tvDrJ63A5aSllzEOTFp3qms3EhOSdN3gPfw2t7lXf2ElsGq/X0LuGSRNIW
jSSj6tze8oLTSqYXBxii6A+2d8jNo5xiN7qUuT9F4HxZNUt98oUwVhGH0q9FoLAk
Z7QDrquUFe3XWptS7wjOVGog56KIrtUfqXfcSs3VfBwJfHDm1t83mPW8drPf2VWP
HkiPngeW1TqP4z4MspQ+2ANBuaTIcguLJhqbaklKJ33B9TxI9BDvwGvIlJevHiHY
`protect END_PROTECTED
