`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DlJ1oaYdKqWr3pjV6LC1Qe/WAw/4UjZvIKOMq5QKlw6ueG5kXB+T9hzFWAxT1kFD
bkl1NZ3OYDqKXGr2ywevEE70+RTyE6oyuh0+SAGHVFnnX3e3CINeNM55ra25qtEq
y9qlOHG55V9zm+Ux55NFDHfytemDRjoZYy3dNJ9Ld4ExxbiXGPnB7ltoCokn57Cm
2prItNYDo65q8WYmiSEW/LvpZYdYJBthODOaQWp6Qen9VyoxSF6+9lpDQKgg1qMp
lfDix3qTxPxRHeU2easC5pILw68Cb6oyL1PWs4iZOjgmAPZlRyYMfdCFLPkIoHQm
XuQRIK96NJakuw21Ru+c4Ky8r2xj1S2FtJfy6GopPp2U+TMFbmz3vwBYlJemsvOh
G2ar1BT9Uis/KKgnK6bnGZ8zjFeM1t4tDqfYgnK45OrtHbg2Lcf7yG64VH5oDh86
sQmAsCUNmFVL89I+0c3RcST4fcBv26yVCmXhc/hbfyTpnIdrFgNuS73/6hejK1Ss
TrimQicJRmfTjBC2G4Ads6pM4kJ0yyJGkwcSLh9EnO6P+4M3tCV+0nWMIK0A3G1/
nnu8HJ5dtIaJp8sujM5bsJpPUZeSaKTRIevDtKaU26KqOqVY0Bup6ZbS7BI2G2Dl
RssSWkHh+0Suu9tb27wW9rrMNwjXfiotP+vhglK0dh0DGJ5eGQ13tTTquU7q4t0u
5MfnlDuh+Hduew/MzrVOnFSaPtOpkWVOzJ3V5Xi6Y1i8iWk8S1Xse24TDfWcguzN
TXCg3ORh0rphtLH+9nMrvHhSd7eHXzLiyEN7SAEZtlBL30toQGxuaKTHHJzH6X2c
low0vs5jL2gWFfYnZkNaa5uWZH9czUHdGW8ZY5rUv1ec+BbsZhuUxkoPTvOqFqQD
zOeZ/WxKnmMT/a/vJ3niW/ml3qyfndx+zef//y6+XJKPxt7uKia5dMqHpUky/mW4
QVXb+Q3JCMPX6K7XyOcaJ8m17o4/T0D+QVKMheRcrpAYJK0YHAYwg8CV8vS2qpm0
8SQ8UKgQG49g66uF9OzzBEMwPTelCfnxJvV9zPJVDUwoZqcekS9pEsDcKhNScYZF
/j/aVueDDLC74MVT7dvWnzwY8+74jRrYFjsmJLeSIDQaSqBBPc+A5E0XjYFnakkr
jyBtZni14XxigmjU6hgMwTdGzljQ1r9RAtaNTKbAeO7xuU5b3mT6nyL4Fbxc5GAz
sezKRM+Fr4QCJrGy+PwXGtWETUNphMp4iC8ZFAg8sUT/JT/KBIQ63V0FIeob0+uM
kftlhrtExMS1mZ2F9bE1VUFjmlCMoNJIMzyeJnA8yh4wty4VFLlg0NqthW+aOHgI
1kgKS7ggSyjyldHOLpavXgh+BAaDDzJS1M/lZ9RjDYPKImi2vLzswF7bt1KovOfn
NIZtRtaNra8Jx76dJbRzlY/5x4pCFIgFSoRTvsBjbYEbSE/CV7TPJxhB3uqOlTPe
XYXYQNcNyolN0xHYo2tOVBG4eeR8kpXttkxyq9Xn3zrWxZBCG8RW0E5APnrxgC//
HpymKxfPNOAmdk48T7A0YpgB8d6PBN6rWasoJi7wyPDLUKqOY+MIVoYPuTV9corN
cVIdnx7LMOAo7PcUXJq8xz+blZ7K7sUuaxfUQ7y68Ig+7oYG3iXzD+MqAP+FjXVZ
OnkDwXVQ+zT4NJSduoT7QJb9fnWlpEZKmFMkoBmXP8wWB2ob8rg8myfx1TgyHUCx
szvCBDMV02Xw8btlxVDFy7ounu69mQbHKVicnBHctYY2W+vdE4TQJeM7HyEa6Nf3
m7H7yylI4sKzwJyK0ivWkHSifi8SEZWGi5nnzgBBnfnrEq1pYUx2vUSzA8U05xub
3e3n/Il5dPvohuZOIMwSZ3Xf5xHyWryZsW13TLPmD5xC2piBYs2ly+G6QNN7Lbpk
97rYrfczSwdIniYu2TviRtPQBNUeM7gYJcjympzIOTr0iYx3H2Ia05OuYxcyRGQu
B/YX562VtPxDu3pFJa0hEqD3yggcKLSkPjT4DvVJJhlQl816QhPBVgLp//szQ1qs
jcSDtW+u9/vro4mw7v/kbnmoCxP3QxvsCQ7nZp+ypVizzV0vt7kL4PmcGEeN7RzY
oK50SwgRn0Jp6CKahP94czTVJQDcJBmW5cnk+cim0ih4TTObPCjDk+GQTuIfTFsh
nVAizd5w3UZOILLvw1hEZ6GPa/bOkDHHZDttDq8j4Ekd9MdnrU9lY+gF3ZaDFeqZ
kjFOuXiaQVP1lVgXHpNkBQ7k/aeZ61v+NHS0/+IHnd3A+nUABXd/uVR7ga5BrQzQ
2XJ2A45l+GLhQa/BHm3Vk1rQ6hAzCj0yd78n3cBMR6nDpRaKXE+R5L/TrwTbqcn3
J9JdzdE/NsxcutRbhsfFzldcDeDbS5lFql/BXht9ZtJ1G47m2oNJPPqtTQUZ1bIM
j5Zqil4P88xsm1FaEDstgJHO/TLdJOS3IkJHZqZcxOW48lHYBqUq/PIAGYCszWHp
51FAm8KctS/dVeMHgJtthk8QP7SlKTbW+tcFvxljbNDmGqgF96Yjs0V6oD3wmGE5
kKKlhCkevTCZV/XNglw+s/EPKZtbzyz4IJRGtITTQttn5JVZPIcX4zYOqwdW8QzS
Gwb7wa5zTSsL1pWQExzid++SwW0JdMkOO8cfNayW9KgZy9py7nap1pa5BWIiIOKY
VJGkeW8OR9eu+zur93FMuSzdRQ/aHOTPTxZi6g+gRU7iWtFjGKhEbU/QyIfwGVhG
zC3y5TbOR6YylVOkcrA93/oQt77sccPKFZFoGZ5E2APYkf/tRUbcr1etbl/LUsfZ
berD06/v/Svqsoxp0fn7e3F39k4Btei3tqTkVSuYhQt34idcv88mEdXA30Wu5PLr
Z6yV/kWBXaau6QVqW++dio44pBGIdnoW0xsbEFwkDbBpoAx+9hoSvrSaopYWsiQY
1sf/kl+BurF6z97Ge+CHG5KYLGD6211VJavESfuNiJiZ8rHAqzuMoHcR3p8w/na7
4JDEZ610vlHAMCh55EGX3TiJIE4Godgz+GG6Vf9BvZCIbDRuj2Rc4/YZAQ40UQjH
ybA+z9OChAzqSQlNFJlouJF1Ug4xukqN2VdZbyDYH4Bbsxu7FBaQ36yWUsHwcO2y
EidWgBWwKl6Te3OpOCRibGuqlf/+76bCcE2HRjC8EdiMuWpw8oBCuTpLYhFvlb77
dK1G1VDYJ1RmkiwrOufD5F9ArhljY/PRq7YTlaYWLhUiZT81B6C2VawZv9uTRU5q
OsnxVOe0VTW7oZ9mziLgi7g5aKDhjAelsHpcFnUZ579e3ouYAai+uyDqHnHhj7Ap
Bq07khuWqieIKU6Nau5IXRc/sY0XjuGS59PN1UNw9txQMo9qDfcaLEL83849X4K/
gHD0YZ6yhwnjUxVXtA56Qdd2nIO3l7o/9IEmYXr/kwvKI0S6kQSKyNxDFc0pV2tp
qVZZo6XlDfLp77NB+k3Bf/Oog56ok5alo1Sqmw5w2OYlrFBEoKM4V5x1JLW2Mi9W
JS4ciFjHvl2V1qZxAX1UfVBVAaxdHx8ksM3eP00UA2MZuZEWu3+ustV/Kb3ALsz0
5hZ4P7mZ4mRnhLb03J470ZpKvDz8GYOfS6e0LC1FH+hv6eOYIlA5BlyGwKiGBOMf
FFiO8GLT8BaiEytHo4JhDN0uQzQZI3l/sBkleJ+IncFRO9/pYfm5KJl/R4KReV8r
+rb/ixaViZZFtCE7SYnWIqxh22Xjbji0mWoCIq3lZ2UgIvKJWmA+1c1hVgrKG2du
ZMj6Sr0Ikm1Axt3IkQ+OFg2HLhjvEwFopP9ylzz9VW73sESLIemmiC5I9FysyUe5
LoruEtg/kWGdkshtvXZ5G0wdwFmUmiWsra8ZW+cxFgFyoyxolQCjg5sYpj+auFcR
9T+HQA5/ZCBU5cucm1acts/OODt9teOXTjlh+rZiqmDx/KT/ZqJ30N4kGc17jRUt
P4Z+96XGS+mXez1ZPOFNMWbnYmOm2M2XfjSI8J98AXWuOoZ3lacxWEyV+tyUm+KZ
p6yfcBOgPEyxXJLh2yn2MDrtABKbWrLG7HG5BjIG5YnHH+/B9EntBnBEZ8+vf+UG
qOEttDaB1XlYlgTXDtER4TwidfEPT+54Z0XINQRw3S6bZYM6YN8pFFYNSgvX9eeF
zJCMnw9TvgXYu6gOpvvrdkk37d/6e9dtszp1PZOY0pLcdPANSlnawH0naCCMLNYs
GZX1lTeQfGwcKvpnSm2Bc76jCXShV2L6gIanaWoq8k13SvJ+KGH96nYA4PD10JwX
dEik++3hYi1X9s8YTLKtAFZ9d4KvJUE3TXO9nxm9dXzV9de+pS6Xfi0oWPMYeanx
FCTLXeJxspepPHygMAHWCgzt984YLYJqVOioAI+c6jL+kvBj1rizMriLDMKMFddp
4dgyU4qVLusiK/SLHrSWvKnoUZo1txfPNuQ4KyUOMpGdEvZMty/yxjByEY/5c0kE
iKvT0zrQWK3XebqLrjEcn0XXwVz5HiR8UfEL0R0cytPDH1yU5VgyUkRabWoJ1mt0
/Lc5cmAC7vqIKW0Oj0LKG+1ZQyUCJo77xuRjTGX3IgjLejhcXrN2hq7o/irqH8ou
Jpo4jP1htFpOzQrBDLeteiuyGvEwf7cVfsnQoT/nEA1dYgIGfPY5SEVGExDMxjdw
xdnQBvP9Oi8xb25F6g53gF7txpLDHhYB3UTRoCOTpA5eYqnv+VHr/pdvxX2LJnDL
vYFW4UK+OemTPtHagW2KbsMfO8BK+DnAVMHEom2cLKjU+YvwEoRT96qX20M+CzKT
x1BFA6PAMNaFmOvaYYDNyA/+t8kGYRZIFpJ93QMouAymSHuBhT3tzviTEkvWoO9H
KH45vaZ+dQWIWI/9UnxvBrs+9yjE6w1GvtwT+VhvW51ft1q9Ids8KbL5VSH/LjaA
4g1EHllaDMALOTKBb527gCr9kbTKNcfA+sOJ6smrzpmIIh5ckiZAGJJ/6+ldNowu
QJJVmpxBb5+fLsmQRGow8QmZzpo6qsG8on9LAqA8KKxvltHcF14QcGYmQdRf59FL
qFkQPo6329gm4UsHP0CZbPbGDFA2OF9NPbL6cNB69q+FGEMJZ0/pVJADSkUgQDog
gX7iXiIrAfs3mRNObAQt+GrTiHACgdaSphaS/smo/6BuJtoY25+KPNohLQjy6Umq
3CawOoOEM2tufNFaH3LBSyAgkyOrmNgaQ/ZtnqtRN/YIa3XWpO1Ge2neC3kIhOyC
ry+OsNZ6UhbrN5JfvC5mr8/dLPcVKcUjvZ2m2fAiFgOnLA+Y3a0VIzX7RCz/licF
VZc7jAeEfPt/k77vcl93Uh2W21ckybQzXSREnCVub7VYx2WfMztRHb1zMx0l4Olm
KC9ygKKx9YaJoiWogt8pwnrsVef/Aop/3pcj4zvwA7BZlAR16usdg40dC1I3iv+E
S6RCx40fEYLpfRFz0NFnl/sAwWJDs8Tu31ws9ZMb9fcrKRLP9aoiotUZEOnHhiW0
mfneFkrn/dl6u66x/L/RVzmNxYXIUkasvzJdnzD/iuGFmpBdUYDdSMwUVqBpb/ul
ePWB7EfWm4NQOCNWbqu6OgJWRTxdotm2jpgbC+/mUcDUlNTOup4UEN8RD1/tcKyW
i+FSimhHJ90nrLD15UJeNzFfDZqrbAp3/JJBhL3N0XZp8tDvzZIJVESEN7dbVjE9
CLHj6lmciM2FJH8scMEqZzMMFMLSztFNOd9q2DRyoD2JksHwglriopS7ThrJFf24
3rSfw04D0G1S1GARMfPkZZhEtO1B2pqWv6T53MjxDKYKn3ep0iW0e62KudpZIxT/
UOI/TWXNTVrSTRCCqVGC2+7hwwXZLuN9zKcrUiZa9doqv27XH1t3BKcH2TO+Fj2n
RgP6uisaSJDWrnkpFHaDNJ7kBnWRZ0YF1CANkKDeL6IMGUVSwBZB+jFZwtVIfsYF
TEtcBI4bejZYfSMyqLfgNdpMSHOKYEKRPxdSoR2aXKLFyBEIsWsTYoy/U0uCIMl/
LfhUtmkmXRRXrjYb6+LlrtPBAgYIGar7Ui1UGTapVSt6r3rGuhjim01PtMRfetLC
2tLpR4NCOi2X4yLFCMyEyCJ8eUyvfrxy+Zy7CSEeAlQjBHLFPYv4IF+N4W53TEVh
NTJDEs9ZGHkWoWpYx0QizeHycGdnbY/p9BJumPh3+ov7aQZDa0etKBYo/4YXjHpK
Ue8scgK6+K67WXwC542fiQlfkR81MH5KiJAd67hYoD75jNxUl71oj59C8bg38eSU
p0nyL3c4eYTt6jctSacxjp24vC+yA/jLMgcrgs4cQJCu2upCS7/RZIryLGlEvsMp
M7szPx0ixf7GZE0w9kE0XanKn3RvAI42u3+fMrMU8jcr+8BKQ49Wg/BlHQ6DSNmc
PjHztkfv7PXP5SDvOybB4khHIGbPeIjMSSUL0EGKG17dZnhu/MF+mm65qi6emOkl
WPywSFpVRrbr/zYMsUL3RnU1ciuqN0XnP1xsUBuXHA6XhX+Ho/+tOchS3h2PY15i
Ab4kaAJb9kSgxAWdTzqcPOXrj2O/mf4dV7NcpdmvadmDxIwvAgoM61JGaUQ0a9uN
V8I42DTegCMIac51WAOrffnN1RBqAF3YkJYBCQYCt+/I28v4MRZFRKEBBx2OUqS6
DmwXkWSwVM1iJOZdL6G63PTpVUZMrXCXaxqucDVqctcG1wH4O7P4p4wGUH/V2tqT
mUkG+PR/t8w9YAKLik+5l/kd1qJJWmXqw6PAMBtZphmZSso4bwY1+rmMQG2ooCDX
By+fN9VfFaa+4yL7LkTuIhsaern6buuV3qqrJPx6icAU3MkU4jCCuSmB//r0p/lj
LjeRZtFARCD6ceCvwkszU8L8qCYq+wFo6djiGD/geuA3uuOKnlwFua7Opy1NZBkF
fdLJ6+mjQ6vTIeUs6C95JMJmRY+ZEEfbXF9rMmKpjkfjvkQ50fJDAtbFyN/ufUu0
dKLABychfuB8ELQn83WZxEpsfXRRTu/p6AYnVLn1yogE5JnAH4OPBrzOyJnyjP5o
VBFvJ9ApCyOrXfhtFEMKwP655JkIaJ7S7H3fzQ83SciuatEmKlNUAONYN9R5vRZ1
rUm614ssJ4vi14ZvxL0aRDUnit3TvWybl0OMCN17lzQsrE3PWyrbXbIB+8mP5w5c
Yku7ez1jaaNYz1jWL9saxVdZJb4VG2LGeBC7sW8Idp4E1s3B13r0L1xeIJBHfiTE
QA3FykIBMt+OBbZ/iOwNmLc8yN/x4uvz0w6UkyDstyrWtW7VbFP4Q8IydbUifSQY
WqmTYBW9WoRteaphEyCkLBnE5XgTTnMcXzxwbfQouvbskOHqQckIOrzm6jvzlm7X
Zy4H7GXy74HZ8Am6skbcGOVNPr8Ht7UEMcMh4anQDrlKxnqscOR/k9BOHCsn4Uxd
8s2dB1+kWobkr9YJV/LhJwdQpigJ6kpGJMPbfNAnGf7WYPVPvAHGkCtGpqzmHH46
A6mZM0INHe4pqffoQQqYAHLOWrZApL5FGym9H8u9QFPOYPs/2DYEnVcp1zGTVVSa
pM2DwztNiCQhUQFuAUZP7HFb9PlQkkmaG+EMoZy9lgpU+vIfQ9Jps3Tx36oRYn81
gv3VifEiLimCfWh2FnINrU496NFyJVZ77E+Wk+Z+8i+LaeSYjOBjCUXXk+ioaS4q
VreB0BIAm1WnGlJdXUO7xWwmWPsvj84/hyx0l6bY9CDuFX6eqyycYrLvJP0+UrVr
QdATJ4ThS7POkW3s7VLyjKaAFBgjxgYVrQDY+PX1dzsFV9abLnkBED++viOG8hl3
SJB1Kprhr1MYTROuYGXolgvc4kbsYOByLF4utO6Bm2fS9M/wySx00G9MltPUPghQ
4apNqyp9gOWd8/3waGvReLKJ9KDPG81itMdrKQg318O5feCMTN54WGGbr+uYzSIs
2z5qmfPL/kP3+An6lYiqZj0uC+NjJ4fwI1Z/20ZeadDzlPIsm7ZkDJmlAdpujdQA
jTAB2Zy7BMyq+gr26IqzgL9yjSuPUMtoPraZuqzz/FAGuMlhULEWSSmuzJy53yOy
qyDJmxcMbYH4ssVryHkyoN7zosDgRzIN8gNu+/9JDhxf4usUIivnAMfEFsGZqrUh
VCLxKTNhTFGLqTllbiOBjoMZ1t96BGeZxV9mu+LgMwbk1Q53spOXIJ9oypqwjBzz
UzVibIC83ZJPGNudqAPJG1O+ohUaGBoYqib7TsBLRdRs3Pzit2BY97C7V2xoP+hK
8rg/d20ygTYgS3J8W2068/6rfdYY83ejxf0hpW5xV3sB3jUuZDzMDxZ9ln/FrAdh
8mywCwSDwKUHkm64Bbo4RjAFSL9dhGq9yD8IH7rP9GcXWxRYsptZKcmU4iAA+/Vm
zIhhb7hhNdunWthtB1rsq6VahxVKWGPfaupDxwrG89/eY2z5t5md0eLSeoVMd6p1
wuly5Qp7ymHM7KcGwMcsPLfS5GM6VSwms+M0J3ox05GOj/+Ob0Iu+jrgKqH5/ldp
H/rx5ZAfKOPpwHwINTpC6KdFZSXivFvIE7Cw1AUWL/HzJy4B+Fq1n39Q/wXiXvNi
La4VF6fLQ0nZLTVoUeByAZTFNImYdDUPYdL3+1pcyFt7jlBWHJQOR2Z4GDKZr/BF
ovi1Zbzsvo1JAXTaNRieU5hbijEFoxSSGm6iHyASqqwxImgD8OUP1a16mskGNPN7
d8mBO4A3/op1F8zkulE0nCQaTl9XezUahdYCTFUmfgVxIr8vhP8BEjbQ/RgKatMd
HpGhNObjZd1Lx8SvaMslK5rPn7+1yLHJRH1JZOv64UcuZjWzfopA+U9Z/A9Dg7KM
5KinxBRLz1uN/F9JUEbV9TN8RMlUGyTyooBdyL+O2P6P6tVdQf5YtKAwkw7bLAbn
MjOKSvt0cjvKKIJkWfuhfiBRFIaHphHBo7vYKGwggmoukBK8MHdit2wfvMjt2pjM
sasE7cJZ3n96TUgFWX+5RuWm8gz5cX5CJEQpzAGj27X1gtmAyxygKfu3tVaIgKGR
U6F0zR9MxcLUjnZ033tRXC6/cM8DQdUs0IF4kf+BJ8zvq9b80//wDowK/YE1Y/4h
MxGQpN2BVIztDpB5RUD9m7RDEeoWoYzwO0wRk2ozaBvUBzzqp+qkcnzG+yoZBkzj
S2Vqmm0StL6iGqAscp+hvs7PMxot7oDx55RC7jlzXvZUCFBL+D6orXRuP6TfR6pi
tCBWrjc01kMrhbGNnQic/CtCfWrxRaILg0CZAxc+VZ9o2xYknpnP0B8j0KvfI24z
RLYKSp5HLRaHkH5D7PDv15AbnORF8oOUv0tt7eiXVhFUsQKYQmur7XvjoYRHGkQ4
KJK4IH5mBkuLcniPqTS+QB3F4rr6dQczYHlqc5Ox1218mGWSBguMC/iqYunxcoTe
uTpyCu4pOdcPcxT5vaIc/8LzmSwhCWHxe0dKC7QQJdZA8MRHwLuvN0FoK2Jb633W
J/dd7WjB4E6iKwPF3mrlw9ooft1nUB7PPEogpXX0s2CmEJEXqgKNvcdDuU5YuLk6
AW4591qDo+fbOcI5pO+Qfny47z6ygwpL0rOw1Ag9jp6LpfYJEIVzU2S9b72n0Smr
Haxd0BGa6xoS8VzPiqeW8Y41XsqrDMgKDMXNW6juGMH+8Hkle08azfosxSp+Yis1
T6iN6sP72sOB/euHrBtYPDaJl4Yb3QPQPGTN1JMpgYOTwJnxvwntttpneVNxPXep
CnfMucxOOKJmKBTMoJjIo++VASDQffZl/b79byrgpPEMPAugOlrFH2TvOlX99XSe
FetaBRQ1jKwrMo2tdRraMZou5PHVe0ELs/gUVzIH3lb9CX/KQIiQlL5e5lLCKVqI
MBrZRruWwqXz7IXy9Pc5laRXWK8e9mygK//Ucgi6iTtSfyIcaS7sBVDidia5HlNS
R3mOs5p3pUOaDLfTLae2sheTwjOZEyh9hCA/WplffFQw4MhX8hgdCZSnhELpJ4Qp
qVFTudJg4L3oECXttTKJ7DxD+kcETjjVjD/MX8ejcBcmskx4WS8FR72v8A+IiaYR
U2pZMA3k3/XHmWOniozEhCtWMRoYd+cG+Lz9CSQN59xBEPH1BG3l8SytQuJH6HFr
5JcMKeASEeFotbR6uII4xqI1Kxy4rXM6xTqp/a9FeaeR+imM0iXNnhlPQbxyXLX6
BwOx/Z76CO19sFXX9Lup6Gztx0oBb7eLFI/6/a30vNKTpCaanoplZMjCOSMxv/pk
NdDb2kdsYq7l6Z5QQz2ktTJ1lPI37Ded3wCpUi0jrM14WFeEPWjavHCDg9p60q3m
gKbkP9NgrZR2HdCP2cYFPYeIamASS5XgfewBdejkIRYOipgIV75SQNfvxPFbmDGQ
NG1tKtSfB/rXOmYfuGXJtQyqnv8QpGkUvovNNfROVDI+Ks+zn3BHNbsMxhyuDM1Y
49B3q40pnPFum/DXv5hj3uMEJMflC46JPBeTzhxFwoM7dYGA0XiMCKydpXKpLW6T
lX5VORiLk6+GRkqB9YZmw/g2BWhNXj4YDK0syg0u6cgx4THceipoHEL5Kraz+3Y3
PAzmAh707JzBOS8NYB6nEfPg1uij+JVeo5nxnOuUbUUuL6YANFIHPUIg2R9RwNNj
o+bm/MHr4kPcfcwWVT8+FCnfg7Oe5rCfKZhf2liI5PEmEbF5ripE3S/qGNMwzdVI
pqcPma98JL42b9p/jpiG6HN8pCONgjwrYXgVGb0UH9v2Tg0nmj2L/6gl7lNItwYY
Ketem0lDIqxQzUgMiVyD+3PDK7RNL7IUxOw5a6EhuRR9rCQOY7aW+SVPNi0XFNR1
u3Pd83e0AS15fLdy9dNjnhVfM0Nvl45+Pe/fN+5Esla7OxctGsZN1MP+AQl/3vqD
KzbqayE0QvsYaPWrph8mdvENFrWADPdcUpUzmU7RX4dO4xZTc2mPATjTSguMw88d
o8fpZHvKiIy8UWov4TFllwRb1bGy9yMXMWUHhvdBcS7SMQQjFKJ+Cb2Zr3UZ1JQt
l3TeOgHfXVJwMp2w99WXKg709pgNLq98hBDTwxJcAG4CpLbxd2yavsTxi+YGU2rg
qIAgXL9/Roegx5BQVrWrrGkEdcju8vvV/Vg8NouE2IiC3YNyH2zKlLFEAJzH2T+Q
+tIy41RjKt6C7epISlAbmUxjUGruJzWP6u+WxF9+1CCILUD5LHoVIwlf9Qwd6BGd
9bJz5HWP5bJxsg/D8IHpf5V6n0mKjZaY7X1E95dWU8IiD/2sRkm3D0y7qZUW3aIj
q1V4in8YH0kZ3RLlotJZzym86CCO8CQDtWtEBmVTpAIsqy9ptps7djL7VO00cE+/
defzs5SK07n57Ndr8QpJb/jbOkw4wBXq0mfuBqDOcCJKqCvzMYj3EqiivydDRl4/
rTthN/0ZblK4WohyYS4AapmxjKq8HJFIB57BT9Z4roJcw7LTOJNfPtN9JiyxWhRT
87pRe6VHnVjXkUaFbesks+lw9Tq2fBH67mJycG3LR1/XErOmBqY642JzgRrf9cq2
iesV7E+IgS9K3qZyUQuaezbUQBXPNYRNN/niWFSJjLq1K85CdYEC8WsbhfkV43iY
84UZyg5ll/qYacFKHkz9ssOByBlCZlhtW97VqFwfNlx5c+dJ8HT9HElLbmdfg6Jm
ebbMETorIlQ0jE7H6fVeE0YoU4qtkUdcSdZD/jjZuBGsQHjuD/4yXSp9wvBOf7Of
P5DoDV7hh2cUaS/puuBe0qqOk4U7xJFMtB1AsuYWH/MjCw/n2FyJ2jH2Is7qmqIB
SOktgUP2WnTbNhD8ua2kz2cvBJq+ll6aie+5MjWyeEOQ5EOFuw8g7byYFsC4fPE1
hILaYck0v295p9rXdr9HGueVN8pL1b2f+wLcHrM5AsL0mI7l8TNY9IprPXodlPyK
23u4imT81+5xluvE+BU8aE7ffSKUjku4shmjfNGIestYP7vO9rv8ydiQ9VucrTxD
fSV2gCrZB2Q4paiByqPCvcLuHE0cJ1+QqVZj1T3PK0bZPZoYRkaMXbzJl6JFSgnH
rDbmiNGX0/6pSCkAUgBSsRlGHaQ4KQounjtkO7xTsxAAXs9umyHzhf+380nsBECF
ckPC2FLMgeLWHfT26ZsO9B+D2LKHsWHSVM97hHzNSC051KqLqd+xGGbJJas8/r5Y
G1fmW4l+CtoDbafxP0dd6Q==
`protect END_PROTECTED
