`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hVwhZko/3iwRThizJjIP/u7XMtCNpC4SiVOJOWtdvTVZvI+VEGfp1sCpBCNOwVQG
9OhhkaIN1ftIDWiCfT/snzmdLohT6FNa69gFAHY/bHIfPMcTcPwNcdmt1ku3Hv4l
vQE93qTBChhR3ZLBcsycn1Smyex11/PJEZop8gwtky8SIIkrSkfy6ktfMtJm+PPA
LC412uWIY2w/o3ul/ct1N9c4dOc37bhOzq06hxpeSAd4/kOP4LKwKqZBLaa9e8ZQ
yfgJ9wv7xOKBDF4CID74a2BaIR9TCfpDzZ2p3xOL3LCY3NKjnBre0Wc8tuaQdp+l
uOT8RS7Hb95diAMXZ10k9kCl2WD+AaFGpIX6lbUYPBmLtJNUJNi2dISwYSzwInYu
FUmnLpbFvsV20ygVZAnr1c45osnQbmIwTXEzB7TXrw8=
`protect END_PROTECTED
