`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ayXW3TrXAGamTNPz0G/sNGGYYQTG/z8cDx2WKHIU0oUmBoQq3BRRJLq3o1Sji/G
EXBXyvkW/y3J38BhynrcIZspxTV2wIGb5mo00B8SqLsvBCBaJJ07QEDPXCStSXlJ
Perpye9zqNT69P2rXr3yyc4q59khFwDl6/bBiyqUpQtvweHzkOCnBjnzWHiza0v/
F/5js6dHNl8/Z+vcQJuJg2LVTbEK/0nSlOg9IciHFj7tZk6d+WbPn8udhZrLyFgJ
2HHrpciHPmkeJyDxqzJsIvZfAdKq2NFPCHVJS+zQ9UHR8wrnIAEdqk1WAapMcHS6
oJV7vCfkKNLwIeyKew6Daqjs9UvQCJcNjvH2eO1fuYA5HIw5QMgG6DKdCKLt1Nzv
HFBnSfr6LKYp52hCGNY3zoz60ic7IW8uYSUOdgnEzFGmrt5dhdGMoEAda3oe++zy
HkY/0a3Q7kjL6uilvBvSz9n0Ddk3GptNsfXnVR20VwUjXJK5A8rqn1q1Eb6u6ArP
crKlE0dtCAN55+hiYcjYyzg3u5mocIRnjESEFeXJkvNfduQHQUVKsZidMyJzcikp
tdt4SoSzYD4B0imMtVIFb6vBG32Z/U5cJPnkgXZUt50fHVpdfasFK2O6dHy6Zxrc
1fOuW8s7zI7ZEaUOMUPbsesC68QZhbIOYdk+G4SsVfFLsVGiMY/UwHazEgvrUsHh
h3i++DmuBlH0I5m0kiB/c0nzBmjWau4LvDRGTRMg4i8cun7OGexNciGHrL36SCm1
XoOeILcKhDcVvpBc2e/4ZMIh6h+4qJ/jVTSofQHEVLGsDxfgcz3fAzrAdel8fQdO
lewoa9ebrT1ZOvhqWk/3YxoFDEonSD3PFwklStfwImhPC1SYzld9HhIKq8Cg0BAK
ZFttfw9EtNtxsYDDuJT3uBL64WuTt9NXtrmmiybk8BnXdMgQ1/7ZEjCvKXDvhspu
aSZIuL+1T7eQ77KOotJ+NihQ+oWnLrQJJid6MD4HBV9AJvIURecGMVokuv6dNy+q
YQLh1ozFeCcKwiUQhaXwk/j6CcSGDMRZ1j81TbWurRrzkwP3PeL18KGpeys68UN0
l/AQU1cGanUUGD4Lbr5ZwiBjPG4rENHAap+aEa3Zv7y3iCwGnUonHJeBA7R8fX2Z
Wt+emIUgsr7fQbS3/TpT0GnX+xNLH1xRCF4BIidG2y4o3DW62cZGQmPlYtfGqEei
uO+/9hNZWMo1TnvqVyAflFUlrYLutJ5mlzWduD5/6dqVlLMV+l+7q9xLSZ/LeFra
KoBcAq1o05IxSuBcTKdevsNNVdNpWbNDoMhCy6ZwrmTPVXXfmuds95yULk5EMswr
cfGv8sQ/Go/RN+tAMCv2u6Gjxbq/fifxGhJ87sTlfVeIDx6M3SWL+U8UAc/1uWPj
CgFco391+IAiND2YM6H37ir5msAgZkS7qgp/sanZzwLmNfFTQcROVfBrOcG+GZOx
Af0Yim0DI6QsjPznJnrrvJ6iGe8QRzgo3n5lT/U+92UYVMfDS+yMQg1orOiLhsuX
CDweowF8tfSmQcszwNnobY+PQWbPlyxswa9GSfrkLjkVXNfcWYZvYm7el6ywPWWo
eHT1fZBPi1rXdEIeaOPAp8yGhERPyHEPxfHPpdL79TyHJCB6Pofpcw2B5xKaLKZB
syabiqM8Co4A7Hsn2QZcf17MS6/R55FO9nZwGkTxcD8Ql4L3rXCwEOkTM6WWta2C
Z62l7KiG7Iarpp6g+o+DNn8b0heOYB4NPertacC8rioJlPDUAYS4hafGJ1lKrogZ
RLvnAaaaw99bZXS2KTS5n2OK2Pc0AG7FhAns9VT6zpcFXALJj/NCCwSkjAnjRTIe
UTbzw5GiyF3zDaConerIQ3nDk3VZdmrABenXYCz7JxZyIsizb7/ZUovCxyKMD3C3
Eo0MZ+OYiHswAE8k7ZfsImly/ih7F74rP6KBhTLFGbayw6Jp9ZVSnRC/4tvWUccB
Bg6QUoFl6diQqp44b4BeeoPDa5HRGFB091SOjtkQzADZp5qJ3E2w4WI+/aO5SOb/
V5IRcCEaKebVTBmLMo5paNJu38t2CvuoN8LlTDuQNIqzjmoovrS4edSFgexkVWyL
sXJYVDDo9vne5vv6DiQ2SQp6iJlQOcLK+ac0UaArCN7rNZC5pXnOBevZfKuqVqKT
GWH25pXrd9PQIBPHqXobDoR9QiGCKpyQYj66GDmCfH09ss2GyM1FMzX/StjjnQJ5
o8Fmgr6YjliBZhtTZmnxSFLQzuYyT5JHxXr4EwA4ixBgm+E6iPuLxWO1BCJolZHL
416/BhdEK5LRLn2iKgy+e8OH0D17sUzPdU2K5fHYgKzE32se6iv/4Rsu9lklNyfC
pJmdMGFRixn8wPjOqTuBxdFu2YCASErD4S7+dKiB4BgZI2XlFZ+ufAp3PtidoFbL
2UeBoBoriUIGW1BpGYyzATEn8LvZtdSZPgN6Zc2rUPxzbcJ5lldS50hkFbEBBj31
qDlSBYTsZUDBhylebZRYPJW7RxPo44DwrZp7HVC2J/rZXQCuMzvNvu/CENnKmtqN
CtUGlI71h/NC9Cw8czdnNCUMLeucdDDToJDV9xNjOnlZSwgcqQNOfkwTiy3HmZLp
lNSug+nPLIlfb/aOFd1R51kBRdFPPXxNVL82sMnCwlgSnUIlpGJhroubo6r0eUZ9
ZLIlVyHa4qCJM5XRkmMUK1q/i4X+x58spaJzOISG5S1XgE54GpH6XHUAmL3SbCAu
NjotvdfRYb//FPFSW7XPSD4pN02Z3gohrLF8zJZcSia6nIODrs2vNIYCRRTfmDnd
l3bdXdL4V4ss9e8IGf5ed3cJR3a/Z6g19aPgTXLQRIiq6rX0nE0XEAMm0aCMp4om
/xATfWB9mXkz5WJuD40FWUXuleVQsoA0tcfzQtK8C1Dm2zZcJAYmQUJ+QymWMQ1M
PDvdeMiVjI8TXob7+rF24xROOzHGavRYzA5Q3Ojdon0JIOt1PXEJ0TKlL9KqBdDH
t2JyBMjR6bZ/HdV8N/47vQdsdzBKggrGf8WYQXAPXk7GRW+x6bw93pf276JzDrRu
qAcpMRdv0yim2GTUqm6IyaLbwyxSTAqlpaNeMyuygPDNur4OFbzAvpA+7YBj8+gE
HSEOp5HRYipJAcmsNNbHqmjjFFV30ZHJITqeggum0AFxHFCToDOkAthfk2C1xaPO
nY0zB18eDB1yaY8qBFZNlVpa8xrdnfviLsAW8RZfuVoh0zaAkt0HqTG9ORXGgvzm
CLs53RjfZHeC+TnENfYUP/sFrLpldUt/AzZylV2wK/Aq47UlAeKThwkpFK+7xprN
CdWkP5J6TY2/nY9zR/6JC6lKJ2DeZ8ZS6ytmKdgAEmhXjUDogCXbaFj96IjLtrca
jCP2PzCl4X/jL5WocOQme1dxmpytHPrKgb9yhVRckqoxqfTCU7MjqNhhccK7HPmb
IDuHPkf983aGExYFw30pEivKE5Uv2KV7Qe429SqTYKpGaOYoxuO6Z9WIrF2TUFxr
XJAZKTPgPiS+KOaoy8Ku98rOALrpQAC+QcvwbvWol1qFdnhdWKadD49Wgp9sC4i1
eaLA7J88oyyL0mSguRnMoLAyyB5LkfOSzsJoR/zK8y7bVqMuu62+77z49nyCiMSZ
QCi77UtWqJiWu09FDuLbtBAscVihiROsdo7Ki62Y9GJHNm5ztz1xk5Au3yM9NipJ
Ogjj689sMNjfOWBbEKODoLwRXf9vvkZMKRL3vgtZLnxVlCJR4ceupyZpeLYQF7cb
QAjVVsbp+WRsnaonKgv/JVQWqXSu5e5YDH554GMipTDwVu1jhVZ9IxJzFmHTrFRk
MN4RVZDnlrlbTM7iMIT0Qtx6vTfQlVbEfnu/BFrrnKrTfGcFTWghdbPL76Vq3Tk/
OF1ILa7KHi4xSHyUiDx+6h4MH8Z/eFDLMQT+o0Zl9uZx85wEDn2DBzocO8qsGm2/
rz0PuUFRH+N1hOijxwyMZmfZI6k3E+btOak7wAR4EdysXzUYfOJeQGugKQasUI3W
iCvmHTEmMxYFvlI0qFhzai6QVGt7aVBTYfQ2ewJuwYqI2Y6mfuDhodNkiNyuGERY
eUfCvPSYy/158efgdxl1HwuNCCyvuXDRx5yYl4W3D2HCC/69M/e5pytg+L4HziBx
2COn2Ro0ukA2C3rNQcxuMVcyNeGFRzCPnPcBk9F7o/AqPfdefTJNyGTpqkuv7Lwf
uIdQxvKmL3NHUk9oRFrGpxS0ySdVenufeWHLsi3wFbtDQg6FCKQwXdI0IGHBaNNN
CloA1+hoAZ3KtlmOXtysTeAIcL0GzrjUlV0RoGWTMIQgne2KrgmUjVBcP1GIr9Mz
qtnH7R3P8/EFCLwR8yIhaNwLmRJEhkp3h9UzM1SSdEOitClryreZnJGPDWropG7w
RZg/kYwULsUnSMCcWmxsU8InICU7D/2zYkw3QmPqsD2PMrunaUFIaVVYmNKA50wx
OqTdaKV8ZuDIAC0Qg3cW+pIxx58Bq2MJYn+s2CngUq2/tD8xlkJVvyDyJIGnnMYS
CnDQd5BwiskeT1JAU0AnhCfivFl3Tbg8S+y3L+W25rYwtfgS8plHOC2s7iQ/OWvG
WQndidInJwVzBiNGC5nSH4Tm/iXXdewhF4DxyzSc1klsOjIpB8igQTv59i0YCSG+
pN0Qn6Ie0UbcEyuIKnebq7POVFyJCCjY3Zz7C+/duMJUqRVUwXDZxPAqujgOadSv
ccxlQTE/R6XRuamrkfwk4Kdf1PZS3YrXskasc+T54fesua+vftrYZuw+S105peye
ZlrtZCOPcFYz0h5KRtfZlP2cPAt8Rh+7kvqs0tmNamqMcSXhLRVfMFj9ihW/aAOO
vMDZT9wbfHpV4fSrCzrBg//XFElrpT1YCVYTidcIKl3wVeUtDoI1Z3/vMShVQDhP
FtAZyYhXQqTIavv5djYg0jMqPVrMOVy+vKiaPuLzCR5nJxXb/IIP/zSw/cebo/ap
CgbbV0PefJiCL8jIFWDFO1YxCwNCXc1OdPCY8dFZTYoIEmzpc6Xg+8+SqhhMIkvS
cOaGb5lt1OFMnBeNMpKxanRJPFurYcm0fqVnPztDYLgmBw2kv8sOw2SXl0jqxH8B
Drkp1y7+D2swphBf6ekTJfEGjHlxyTopqHTNcYtEP7+5tGxDX0rgI29Y6MSVstE3
rhN3S1HED08ylUFfYsl/bDayzDa0r2dvw8zsp1SKh1v2/irgJfBwHLJhJG0tALI4
T7RK1SxFWIuuebNmioz/8NjoKq1vieLi03iSgpUmws0xmXxTOcuUsblehH/xjcEF
FuEGNV9owufWR3oR8pz7KRSAtxLSadjNa2lbIRiFpgqIlUmDJfpb6/36AhrNSyAh
+M/7ok3kObJ1TPMml4kcf7sF0ZPYn/JQPguz1mMl/J3Aa90Y4Tw5DU+fNwzJDRBb
iv0ZhRNpiZkD/MT4LmZ0qutbtp5QgisAeDQu4yNyBLYjUk4oQ/jpG6HzsTXz6hFD
/GsF62mBAMMXhtDMzkrafXRS1b+pt/Witego2gI28GW0GaQzQWAE1YTbtnrLAuAV
dN1zDhlKgH+uxW2d/em45gRvJOeRct0GegA+BeVL0TDaHNDi/gjHzpcm73RtA9D3
CBe0UqWQv0DbwpjNYmBd82ImyabfR2BeA3WT1WcflNkw6dYkdH+LBXFZ4khNmP9s
wBSJ7ahC697RPeGCEY6gBthea16gl8u8C48qkcFSiwfFYICZISYQQsMaOn1Xqz7B
CRksDhlbttyrt9GXQNkQRRlqaB9kBMpV/2EEa/jTe//9/Rm9xWG01gNVLtJCk3ON
2+hjbU7Ug7lskhC5Q6eLlm6x+i69hmkQIxE1vMvU1JCCvFcNeEYAtNcprUDuz5Wx
LICQ4WiRQtwhAjIa7Kb6PDhj9ndGiFmUKP8D/fDgHGzXBeT8DYBKKgWOpFmahyRg
TWV5b4/vMPOPfnw2G8TJkKx1II5tMIWu33cNV6log7Jsj6pBi0a3XG8A1EH6scpQ
C1ov+E07p3Il8iQhYU6JyS484skdOxqHfPIFbfFMlubQU0xxs5NNPa2teuQl79IB
+WqES06o+3v9bggXv69+BD8aj9YD6Jl2Wpufv9av9B/F+34zWpj0RzkLDi43MGqA
rFK/l0K+DXH3PQVd7IQ7fRmdiS640/OPmojdzN9NB+noUQ0yBfhEtuxGXyqVuFHQ
5wvXnEY45ZVP8gTt3yXXPtDyy0MLoIESWWkCFne+PAYsL2Kvfbym/IIzh5/0fRhg
7fgYAgNoArpf3jypDPEPNRYiy+EE23A/MsxgFQueTJZ3BH2cLKeUePVMP53N11+m
IvvSZqlYCvLWDPxHbns51miJLYQ83UL1k4MrMpzgQd9JK0Cvyz/BC4dFnN7JjzMY
h4CUoFYM56V3kL0aW/7BolNCgsy6+FcxW3yznfxmCMf9e2mbwgzhH4lWd7TmbIWS
7BRuZH1eMSRFjaODzxf9qVj+/cdJf7CkvpT0jKCFX2POJxzGFoPPOdQ6hBKfCHMh
KwZI8WpFdAFv8yLuMNU1Rv4riQbO5FLobGcolHIbZ3A3eGu2UrScFdPY3BEGoRAh
wxxPhSiGJ4TyKGvkD+mvuMI0U2iTHb0M46p6YK4i7F/odfNOcEg1Jcl0cCP0IjeO
4XZAjXNAxT+Mp0sYaMqeJUMn29M0baCkxTiVpVUHtDlFUhDw6IDLVgbc3+yO3MhR
o7y9c9KRuelIooHd5KPnParuFE1PFkoyhicJug0mkKWj/Td3jCL1l3xkAfUeoQ4Y
LlyOHBlIwDbiCfIz+Yqskz+Qc9OBq6pUjQ07tCUxJLeJEqpJh0Mrg/ftINEYj66/
s4hRkfM/W7U3He+WZ/CBqj+FZfRapxkGtk61QrtMUl2NITbHqSMJSd98o9aGcvkx
QaLMoP4VpE6uTc2GCcZ95OVD7Cq0QXe8AUgnlwV0j+P/s9zpy8qj3Ygkzb2uOt70
gmJPelwwdFGa3MJ1TrOjWu/Jnu87PRQuhACiPOvbbRGBL6ckh7XykHF72qO0Kg3T
rTEsKMW8GDhJngbfY4QPH48EDAMVFUFsPLAgfUqXxfsXyjpM3M2l0dyodDuskShu
jt+vPtXb34cgwL0gpV8JfMHFmwGwWlauCUWnSkzGiqdW2Ug+piVW7rVcDir8EF85
g0upjQvOsmSPQxWOf8wkJAk7Kb5Gvd13aALCfH8unhIE4Mgl4DiMFB7nA0MbhOzw
koYtvxxcwq12VB79W+QfVQ==
`protect END_PROTECTED
