`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1urUSu0I+pNgjmLiRYYyv/grUUCtssxTFTN4FLo8L1uZVZm9SdxiRgus5VWJrMS6
6BUWaP0IdR+HqSS4bDJbo1aNpAHBunDSRzkU1Mi8Sq5PQjnzeZXZRtcISQwK1c4S
hOfS+xdXpvtoFLnaBuJgxJMY7HN+iY0pR0dpqFzwIsmJnJu1vNZ4Ypt1rVvPHSY6
ZnWv7LA5fV8PUIIxv3/z9iBdLWc9WtR04iwhzbqxoBqqHoY2wgLTbdnsFYTMB/VC
fLcCdQS8Hhm8tipZjktvVS1AYTX7oPOrRNRMwQRuUh9qHOqkCVV6210BCo+zNjx+
Ug/7JGYI5N1sT7gJiHJQIPXcZif5h3WPEL6DdA4g6kCxfrlDFaTdMwd8DUKbpKG1
B+yhdEUg4itiDp40dA6cmgry0Zffi15uzTDn+a3T3qi+xbrQmgnZkEkIC8fnpmDt
7xaOdvR6GbAboHkWiTvugZYQM3Eg3cplSXNBtoaLU9cAjR6OBxuXK7tN99khvkzu
lgM/4FENunevwTICiRcMjw8N0Hg78e4M/fcL1tR+hUueXlXOjrTEgiasz2I3DXWD
PsWzMdqD0Wpv5IRyhyKBSndma6YC7GXVfbk2V9Fo5oqrnwj/rEeoPx6r5JwT4oDj
t1RLf9iEmgz7De6dZysO8zfG9gFMMKONGmWf+KEGuT3iPHW9td7jpz96glCC16yb
3+5A9QXMQR3Z511EDd6F/14orjZAaCU/GcG2ynQU6d8o0op0uEGuM+EFegmMCXH6
GkG9tklG8cUdpxjfwkTLQ3Pm5BxFbLjtJOy6UHrygo+UB3ljm45LccrD1CdFRaJm
sEuKRJzg3CLPunEsdrj8zdt6Y70URE24JHBEaRE2rxbip66+bXVorQvWCFVv4S2f
cWcm1At6oxBdMDMur9yQRFku9vEiGqJBoTMnqv1lOtNsJe5D/CTlZlXH6pZSUmh7
RtCe3Y2RFKTY5hgNBaonzXi4eHpua9lk2tP05Y3uREoBGI6BtzhWFceUGSLSGGSw
6rnhLvZo3Ml7Y0K1OZ/XytFSLdYTOQGCO4qWKhy5qKX20kh0HPEsXfCrLrXLihem
eO23lIfY9o+JRUCFKBfemGm0VupzfmkAeMIDmsAyCTm3mebEHmAksK+6DC99AcIR
GNJz9uCXW+58G7P7U8+xFKX2A10/NBbA6J8rx0vlkfF2NIanQ/WkrmpSD2yzWoQT
WIoVwwoFYaaF4swbKne2/9pqF49jzsv3oLol9bvSKh5cQQ2FlAQPUMivMti73xNT
Wv3bDQFRMhygnR78cd40T9dismG2z1MslGrG1vHKgCuZUwCGSX20pb30IvN/bJly
iieRUMdQ1eiODqXOhHolcA==
`protect END_PROTECTED
