`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lZBPui0sdaMoPa0szTSZNHB9lLPoedXze0OYsjP6/oJycOPMk6f5BsZJSiVbnMhf
blHEQu7Mj/5cakUHolbTbE/JynvtNcpET9OfFUFDz5xf+L7L1+2oljqbwwOFWiHx
95CDm3pxTDlKnfXOw9QjycaY70ffqCz6C3zqCjtlrj4zqipFNPm5NNiRLvMWwcio
fN6Ec2ZuMj75TaOpApVJKMuYBLnVf/a5thytAFon3FA1AV6h/SBYO9G2Reswjh8B
YvkdvStxWAGW8hgCWYZLvJHLPx928q+ZsCFReqlyuvWPBFQv35fS8c6VZQu0FiTU
NHlxBvfKBd3PJr7vgo0yejPVr6JBAxiWFrjaXzcsJkzISzeYIWjq43j9Xji5x1vm
DSMXDcEtrCJJ0/SJG7YZnSzb84iDs2HtR2AwD+T7isEev5zvWMY3XsDK831FiM5B
QRKDpEsu+t6gEQvn1qaTpIQbJOYOeJJv2ug+UaUE6h858kHCMvBUD+Nwrepdg4We
n+Lxe/TbitiblshEVDSBB79eOy5wkRAtr7M7R0lsZosJuJ+yzQahNKY3biBcr9GF
T+5AZJtjJOcRJ6zbXwE1jr/3f6A5iC3SkIl1eWewnQkT9PYwzq96NcBI2gB+7uRO
wPieCrW0U9ZuWzzfPVOlq4KjUND7XHRkpTCufQAeiWYq6B2LWCvedt2Qe6kSVZyz
XBTZCoX4aWodNkNZwflKbfHXZqqnJ9HfwrYqFwKRaDTi83wzlVknJI0MSDS7Mf8O
46oK94CUxnyx4LHPaz4IvUytzbsCKrn7B/XLYGBoZpDYcuQB4gT9xBhBprwqIgEt
rAbUpbL0BmY8k63WV2alUTI6I9cJJbsCDCJe69FG7vZ2Dm9nNsFF4yNdWthq7aG9
udZkvojes3vbhl7PF4dd5pkeEq8rxIIrLNzSkb4AYncQsdPlBIbyerfT7Wy2PDRa
CRhXuZslYm9f5YWrOFSIeC+MlNdBUvUlAq2WogYGunn2I/j/HMRxWAtlx2gnZS/a
RCPoWWshktQCH1rte0KSSTNNftA7WnCGg9iivQ39JJ8d3WsLVhX8z4UGijAulEGN
P9HblcHbBoUKjocaICOdNPhaaVRwO+SeBdgy1cNf5z21SZRc22D/tOPmZNJYtzG3
F3wgrK9xmANX602K4zS8ORcGJRQReKoF0ZOw9Hw1JRu/X5sj1Yc01uNNs4auzZvi
4h4tij36wb8LgWWl5KXeIhzQghf1xiyd9CDLrSDfIGkUtxx+W5q6ciXJ4CDB92cr
x481hzZwFjY3DYrtXcrZsZgkrYUfNDO0A2e39mrVJjIRPbsLBcoGZAdX2efnJP7S
yj7SOBBxxVgmZLymdYEOUGiGUHUlHi4ytcs7qUYZBaU0gynAL1ny+PIzh8TUYE9T
bmTUPPNl9BZfc25XnBkp6D+VqkCOZiGIUrZPfF7OSf69FoFpe4nPkxnL9d8TnTxi
jI9ewLSikpfB3eSnhc87Fp7X0YR3fsf9i416QJlgHit/WAVG4PgP+9HaVL4bKSpL
g09XmWIwHXN5lsFea6sUiWtM5VhSkkJNBGq6KRFek3SUUaBe/qgJ0wznllxIZkeL
YQii8oY4pz09cny7+hNKGUb5BuoMFDhlF+dZW+qugzgmjOuLhqvcMMC4tzyM5t8X
oaf3cfIdopKMdYM0LhdntyQwV9qzCp0VZukN2bbNtx8bhLIiBqOXMXpB0n1eZEPw
qsVP3BB3s+CXAer0kaOTtVTHAjjcKR3EdbL/CQjZ7pAFkq9cKPP4IkhHsGEAgMYx
EEfoWzCXa/eJfprJZ5UrC3U/jDmHqbaqt/4aQVrqxRnAQlmzAbHS3IWjhv29hitY
mR+szLmuH6ta/zreDcklLvVmtpbC/bkBvYQxZ3D9WttABIpXx8Z3nbmdco2x4jcU
ZVS1EylPoKc0JP2iXD51M72cuyi8L3+i2AVshp9d4dMeXyRHLblFQK7FsyfMiB19
8+OUue9kbYwQTF5MRJUgUThZKB1HcvPxFRehaJMNxgnhqJQOzmigmWt69jgfDdH1
7U+coNcJkovlBO6dzfquLowuBIk0btHxHlUyRWh8kL/lYasgcBsI0uvVNqPshIdB
b3Kk+ttBwj6hV42JsA2aSBR4YFK5dMURvs5PR6vzwzqt/vnWesoGH+SlPZz9kFYq
hH76x3FYKpzUk4hDbqcaTYb2jGOiITMDFIIgxJzDwUKiabhgndbSrSZFuFZIbh6E
411Ga2/gWQ//y/8CR2O80Zes+7pVbENNXCVIOgxwbsJrgTJA2bc3BPUJv/vp4THZ
4gTE+ECfIey/XRB60PLe0fwD1JOkQjHYo0O4AT1pTVeiqlnPGZFsqoK876675wtX
Ng8F434SzxlAmJpPWPHpqlXsDFfKuWarbiPkZMoR52BWCtbD1RzG31MwegZUOLeJ
0Z4TyWbK4QddV+jwgHCEnzrTYby5rCps99Sp+c+lNwIEzxijR1vllA0ZFw/zlfHu
viOYTJkTMf4ikPdUak+yKmzK1k/MlxyWRDD6hrmjAlJkqKtdvU6IXzyzREYnN0rc
LRStO4b6y7y/ylNFtSq6fo6Tg1qEinZBSZmJsz6rU0koIeRCPUixzzVHW/bNOS3h
EFDLGumpile9k5Jp7uHayonGw7osjLGsnBuBQMgwmZ0mzwL2oHjww6TDJFnLe0tm
RC1CaLCiv2WIhGW6vbjogbF0gsfCrLQlb0tCSELr+MdN/cOd+xlSqj+//3+Hg8FT
1MpmpU/baY4XetwQEhVyVHMsV5hov2cepJQzRbjbY5p6iDMegzsEfR0z7Uc4sKP7
4NiIi0S5eCG0oQiYKVosTYD9m4Q6ywfHAQizPFG33qiR/mh68EUtKc5mloSVDyIr
pvg5G80Ex7O466IR0BuvQPahpkDUtWvpTiK+1xCKV0ezljNi5g8DZ2VBqzzg6K+i
7nQiROFjlP66Dk8CfLQpgbk6NXFzetqftlmW97Nm7mSrOiHuvvmDr1vlYYPGyC3b
sWI7d5D5S/raMiS+0sIhh0AO2ZuZumBCasN5rfwWw1NeZ+VsG1y70OM9mEm3qZj5
WWfM9GrrmovF0Gx7M+88PUoxUGDHUhArp+hbNWR5iBn4rL/+fnE34zravzXcfKBp
R1jMPstZ1uZk2S19rMUPMaAX2uwiXoy/tMkZezbea560StasFKjOdBfDvxxjNvor
L5sKowG8o9Bjw9Wy8ceXXYj6G63H1Pfk/O9BCNWutcXDE/DGNVrJZlPdSPjWV445
wYoKlVzi5LeIe4TzFbAW1MGbFkevT2IBY1JpHKFVRqVpyUxAPzfY2evmAGtwdDGZ
0IJZ/LC9fTrxxpvevc0+aCaAF3GFMh+pW/j0R741qTQ+zrwtROu7Ljv9+yiXmRrk
k2pV0fI9lXi92TSQ/m8ZIwTZK0+pONof1w0qtauHAjpM03HuQWHBOoaKDZj5cq1/
aG+KvfpY/+ujCTIhMUwep3o6xGdyqlSAo3iZlUDpOg5gfAE3vgToVOca96yG+zYd
/aKRJdnT8yYnPJt371Xwg8E0lVC9LxRsgpiLPPQmn7pzPMLoaKxxjV3hlEUs985Z
yjBm1NybWY7CW6+um6mlZy/z0u+na8D8w67w2ZVh+vFKhxwKGfXPeMal/Klx/DKc
+luuUunk4kTgkW6U/rJ0LtlXD0uVgFE9aQKRNZ9493heg7tc1lwr49cxBgdOvQXU
Xwra5CHx8YGlSo3PFMmz8XThZvK6KBp6fYT1/7K2JYexulhq1KtRjMgHAHFodzVo
8vkoq5bL4KzC9KUDNJ+IYHBNbT1eNQGoI5GnMjHROH5CRsXp3cnl2FEsiIMTHN5r
UVTRReLF/G01aSdmHtSH5AwZxO+1wWkEhPcxBm73hrcIg2+0egZuMYJd7VTpYuhN
ofLPDl38X+9QEoqy88PgXgrOJXcwJsjiCBecjG13uHHcREHWvHoZZc2x4tJFKZy8
ib1k/CX1TGHZV1k4a3OkWy1XyknaeGKBbBV81l27BeRM9aacx0HbrJpoPba2KaKp
lr1rvvY2m44Z/H3A4FfGTKVHHPnko12BioQf/6jUWj4Azb1nBt5XHLUAbp/mvTJR
KCpZa1OhMXs00f+tGdPEGB/qUrJcf7beeIZjaL6m5uQPJPoJ3O2aqk/Cck+HNGNP
fXuyXZg+l+BqGSZZjFc0JrZFg+z69UoBUbazJhzsCzCKUjyc2zqVhWhpIMc5DLki
XQkOcH3rg6CTn5/vgeqpe+kB3qdEIEpJZUmYGmzVMXneseybglFRXP1opQS+6TA4
LDMTk7mFAHXc+wlPZfPzcCT2/jm1G45hkZa5wIl+5ZC62xaXh32kLT3VxJIgH223
K0inCgb2WxZQIGy/4mft8TcCscLxxfTUqTlDuWbOeb4+3Hb89ZYJBBzG7f1TGqH5
tcVM78egRxsvWfhGkqm0ryCanbZMLk0nAGErhjtCmdwopWW2v7+G1KzW1Ndu68GV
2+HWkUC2WCWOX46kPrFIc6i3xqfj9GieVlvl2OX4R2TnFeioxSZnIZn/tv/p6iaW
tyLLJKwrxTL2ChD1Ue9SgK4tvo0VJhN2rhTkOCr+DSHkEnpDX/kLLKiKugfcmK4X
WCId+MGUsMFATU+h0MPJQxc8lAj6jLPsvrdI4SliQVOOjOlMOGdR5Oyqb9dgDzcc
C4lry/Ix38EAMCSabLuYT4WiRUvbJGSX0W7c2ehzo4zvr79SzNfRbm5IJdDIGolN
caf5+1fdG22Rr/NRhXU+XK9TIA8LzWs3MvIzykOKtSwrJ54I3/zaZQQ8YrzMJOu2
/NwJSV8P0bFP5nmsMiBmP//Qbe0hiNO5GyijWZbODOAi7/3AqexWWiwqjxnX6pZd
viPD9YSi1KjnLu/J8k+4FgolWIuUzkuxeQTayLsL+3R9cjSkQLH720TNC03kQ56D
iFJYa+8BOeRZ5z/7uFHz8yC7Ke66IOkccSY6AA6djPF0mlnbtG+ag56JW9Du9Co/
IT2jQrXXQFityB+B6YENqAS/NPtOTn5sl4SQFssQobkoIWUqRsTjBoH8SaEeg8YZ
SnFbPwNUY11K0Gv7AEaB50WdRSZWeaGwkXCez53czg7cb4C14E8sAqF6x4/7u+hv
dysC13szN1d/W2TS4ES4lJjDKXAT6j30KvsUsE7wL0BCBQhnyCwwEMHethi6UXCO
0bcDaQrhmhECD1p3SBgqmTsqJU/Ib22p6LiibY0s+nZrHw35vv2JxBDMSbBsPHQ7
I05Jgz/2ZpGqQmOOf9FFROLXF2HvAQ8P61JvVL3RYJ9Q2L87G6Dl6txX5vgEX9Vq
scLuyttNdSJcoYWdQPiHlzBSBt7uFcFSn1c25z57XaIL3TcaHHyp9qYmm8Ztuy67
ehPuN0C0pDc11rvdTf9gMHfloeK0T/r9jE6HgY9Rhe13aE5p6GHILaT0NlAtckzp
oY+0RuCF9oSa1eKnmYDCEKLfWQTa6u7wnvAWin/3AL71L9dttCwOUABjxMBUNYeb
onl0/8Fieuwu6XJST5EyJl/ogSzNaT59fl5GE2320lhtJezgaoIU0wO+fMVOS3yZ
4WIwOdaZN1OqRaHsJl4VFihPVt35FdWnmeoc6DGtZEruj+AuWI038i99RQJlhf4t
jmreRa+etDY7a7B3RcWelLVLDfGaN15Ii+t4tQVAdEj/memhwYpuNRNiqabSfqVT
lRp1JjqKqin8e2oJ1X22+lyfQHZ8ZG73u2Pmfjz5f3ti8h69+G/+4qvZbNTOZsmn
S1y0ecrfvO8RcWxcz3gGP3XADK69M47BOixEHuFYPMy6RK3K0kadcqZ6pCZbNHt5
1V/x47Ge1tGrvZ39bU/CeTqvbHdqYVz05IGml83CRZjhnek3hHjPFVukrSUptqDh
VBn5tRXwZfYaNYlq3Lcf6GaujSae+OFiK/GfWxVw56AjSSipcvtSDCmhjta1aeFU
geLY0ZTmmkQETt1zu9il3g1tzFN+t3bkse2YS94HfUXNcfNXe4g3CQBRB5xa5zgr
1Svi79LWb1umaiehLk0z4mSIoQKhTbYvTUv4oslFsS8QvpVkxJ/CO8dcPZGvxFf5
cT++q36xL10bZPgxqYc6a7TDhvBK5k7ZQ36GYPywlJ5nd6RCl9ZnXYSZ5XT4vgyY
6HHdLcsZHDP2B8bDEo5OLmk8qheS7dRBNU6tW7oFiDEAvlC5U0yZ8OOZP/2LozTY
5Jx3N3xwAO1s8/v8Zpo5j3uxvlLjH3II0QoEoyfINPaZ6NVCwWE2wokPjNcupVjV
vniHmbKUivu9pbK95pOaRauU/WeW1VAfnvbnAx08yeu9KD39knqzyCvu0a8BpzLt
UIF3bl5GyJJZvwiCP1Y6y75dq2N9BGPuoYR3swks9hmDkRjPygdqXMze6hvNTnk7
e43UMAb7LwbdEu7nD6XnqGZNt9ramRHFn83+v5n4wHckSNU8m9NfbqMTy8z3dDTK
UeZmqgW42BwhLqkw6QrXyXi3cVKB99vyaJfn7I0VokHzqjsNY6RLcJrDCpPP+YTw
OKBHG5xfphYRABmZqhWnhTQYleMZd4+ZoR/8h2TPCuxCTIj7jtvK2xMnynVO9QoQ
M8llrI1FjC3Jl6ibaaNxslCMFXSP6TyeuqbK5DSVzNUhzg5M7loRyloAgK3Nq6To
YbcADXxtgDiqDe6OTDBVmzprY+cDZiLcOmsreA3aYjZCW4hhYyTlMjP4OjRqXeDq
t8seC/bTRR6+8DM2J1oRA7qFtIv+RZ2tA3TgyAjkp5tOZp8Q0zt1Bv96giWzXkS0
IkJM8Hb1D9eRwoh3ZOZSiLJ6hNqQ/FJNer23gPRzTCW8uxttvjn+W8dhnWWHxpHC
7Tq1bCtcdqzpAZw7KkvoXGo+h8JLcqDDbtyeUauZ3O+dLN+fhfvxD7BCRcMXupMX
/Z3tccBy+8fIYvohME40I90ZlND2T2HN0CO/ZeKEKX8PUrlI9TtmvNEkHKzkGc3J
`protect END_PROTECTED
