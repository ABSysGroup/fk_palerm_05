`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W1uOts9cyfUd98Pkn8FQEflFSvwvDmybxWX9W+s6zUmw0KMXkeyHtZg50DfciZx2
TAkLrx59m6+3bSzzY/F+Skni+5OdJaIt57qXH/Ek6Yx1KdGliG3uo8W4Gs36Gqyj
qjy++FLTRpsOxoWFbFJu7/mowo2UVUTyKxS8AvrqzJ+I6vPl8oOOBWc1jqoiIpVw
ET7RqqC2gwdJ49IW0oiMd5Fa2MWl9QdnLEDILjDUbgqWsOBGOqBoajV1wmDyJDgv
UwLplupgjXsXdX0vYMGp6uEX5rrMm9RjMv1Auyq6b6UfV8Tvyb+C4iCmcMhOGc9J
FME2Us8imsBx02CzwdwKAhUWKxsCsLht6tHEMBoJ5S1bqblw8tFUX6d2I5QvXY8f
`protect END_PROTECTED
