`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lAURGPrIDx3F0daLU1Gl9CUwh6RX4Hehby0uibIALBzZ7NRX29oOQt/vFbWT+SQH
oZCwB7uwRdXfFnCRuLu/u96S36fqMCwtya4reD8UTC4TMjHeMM/uIdqYUM1Le2Fc
pKJrp6OosbnhxzcrgovYTHqeBKQaVpa78LiGax4MuE3Iw0D1Bh4m3yieZ4O7ACdo
D5YYRVnIQSzn7MZSaAytkyvcQXDFGYFHnAIhn2fS7PS3Wlem+vIeUqC9C65Ch2Jd
Ma2AemRHFoVEYuxtZqGskK0TZeh+Wv3hHkRhyOluKZmxZjGGZ8CFQgT1SWnPNuor
MxlNzq7k3W1r9jPfonTwFYlffIWA8JEOS2FP+gMNfoCN3BwBxJXEHVnfD0YgT7gf
K5Z2fJT6QPF3ft9U2gToKghivq8i+y6P9kF7wugHpa0p9fQYIzlw4Q7fV1AWf4ri
1RVY6HK2BMYkCiOTirgzvH4ztJ055oM3oyojA1ScstlqGUsHm96us+Ive4eurlj6
09Kikl7JBG59ND6+M968Fq0KBWCUQU+mVxhGBrSy5LCdWfoeP+zmMauFiQ+U27f/
vRtdp6hfTU/lAbAYIue9cxZ0vRjCbgW/0AJdViz1GBU=
`protect END_PROTECTED
