`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GZzUWIUP3XiFNC9TRDMF4S7pJwd/Qnuth6rOorms6afWTpa/7WsMnl102RgOcGpq
2JCWSRfCH4KtFGKQY9CK9/smd70tVXaKUt7bgjpC4PzM0Hjoo+o6BV5g/1tVdcA4
/P7t1KMSGYN5chEoiK0i+1lOV/U8cZ3Vch8gPezyx6pRf0yaFF/w0rFc4mu9Stvi
2sHI+f4vIRAViO3Hly77UbOLVcWyNjABf+Ti5GkMoaXqSzn5yP5U8PVUlnqv7nuN
IKxIUozTwy9BRGzVaCydVsoZg1hCyH02PJuKmJ/3N5O6P92STNSFaJ8hsaCuSCJW
mEgUoo3rh6DHrMkgb7euRVhp6ng4TXmeX+gI5RO7nLj1/wOiAZpjFDZ+Wrv7bOhn
DpHYnxDV9g6jv54EyUgNdk6a2L2EDm2qfR/XQwq87EEcXN+WPp2DwZIiJpw9Zdmg
Jvv+8Yd+IFkOcnz5W9xVDbZpbMuoTBds/jdycgex5T51Guq+yICEOeYZNtednYqd
hNRW9LHmDz1x6Zl2h8wmsZdmudeoOj63Za8bPSSN3nc70Gq1TXyGmX2yKfQp/zTx
/Ud/lhAQIHACd8LAAFWc5PWNf/Do0VM5o966NS4IaiQamnvFETHsN9RgsIQosECW
CtPCA9P+0+VjWvNgS4WGd4aje3RpHH68B0Mlm9LVGBljdap6nOHdNI3iaW4olGSo
utWNABs2/aKiUFLudHjDXgQWdW989P2JBGe/sUHF7pJSEBYvezXpK0/DNdpdQRbo
/G1/Be4XcKsImlGp9mR7q0c9jhImks11dS5XhfV1Hk1MLn2rOOL54fNvK1XGTuVO
TRuetIWeuFlKG0oadabQejU3RctaC9USYBFjD++//ou3+Jvn04YIXa7N9lAg3EQQ
LYi6aCOlmLxUz0VK0y1R3sQ+NoFt7ZEq4zwpCLM1ybBsyYK03yub5KJ1DBJUvyJ8
LYw09k/EvG6UUZCI4eZ09pGLudeE7U8+rvSKemoMWTE/3dCul81ClumgpmoyGG5i
tm50zXc1tmNVAl7DnPh8wdpG+LCBnSM81zgpoubKh1lmDAS8AQwKz+ir7CILG718
FZ3Bvso2C32yO4b2zqFkbVj0Cn/zAJsYMD75uhdoYECwcpjLBACxmqKytN8lm/Iw
5DXL/DuPUZwKFRR2HshDSt+t+UomGmmpnYZlrzGYxRR5l9T87S31QN88M0+AxnBc
AMoO7f5x9ZcarrVlDRGhg2YmZld+aHB9xtsZpz0oibydIZeoub2PR1JZxgGPOq8Z
/1nAD5qgb7uftUSZYdQfIiI4DtvCcK4FG4GQpa3vAxu7YWRYPRpLKUO03awwChPO
ws1dkih2Qbiv67dOYCOr/f5fN8d2FXF0gGBJZ48zEcHWBRNWAfzoXOPlbdg5YRgr
3JJb6KhL9qkFhiKv5LiBSFRFRVR/ubc3GmdrCQjZm1rh/hQUEg9xfh6vKmBMZSND
19v/PJRWlyRMSqy1z7CYE+nV6FYUslrwa34FxPLy+tvHYntMEfHylYnAiL3Ls2nC
rFacZD9muRVAM6W0wX41I9+XHWlMy1FoVWucLK+hzG4TpK8ufpNr+MEKjBpjM8tf
TA4a6GLmbfL3t1qPydZWyMu+bMhunCMZyEIaCHSpljDJbq+WMatvo/qHJxtnHMf6
Kn0Xty6zNfiDWWZT5nfF5hu79ZxGjd987njGrI1uiMZpxRGXmdgXB313B1EKyM4B
/sh8ZnFMuNikqpGY5LGV8HPFDQlcV1BFsdiFlX7imCvU1iGGIDcRJ8tajO9csYtb
dntCNSq+RqMhmfceKLoHK7LWiGnVUIcV9mvVgI/UAtmaa5JKVeh/hajgcXlP/hXR
CnWYB2zU6ODfXH+3dD5W854ox2c+wqvaEvrtK7qgE4YBWDF21PuCUdmeLDUEFN+y
kT9DN6TLdvTGK/gPzwEPfI9LKCEzOg8gP8Xz4WCatg/uYGe4210QNn/nKONikTQj
Yxuq3McfyOHOFX4UunHmtRVKzA6zl00502i4AVX29dS84C385Ft/Bw3yEVujhp5T
rJmg4IKReQ9VdGuoEoN/xv+rRpSx4IImVQ1+ZDHuFwVDzMRIZEryjFhSKoonLNGw
rbl+D5HArlRHLYhNS4QfRBm6qT2diTQxXfuWvFvLitnkkb5Wt56UpYqemm+rkH8R
zMHMJ9f3Gn6wKGg1DmmAFb/aEqkn/V/cQUI+u38IWW17kUNW2gBy1084RQjd3Nsz
MCncAOutvuE09FouOiAjpjYOrBGgCQFhnu6lBQe5U55iqf1slvjrJKYk0OcVRHuX
QULUbWKLDlwMOrn0fHzDtGMxT7a/o7BJdw1vaWunD29HHM6HKi8zj3xmdMgnJdEo
EgF7KRtIVgutxt7j5v4YoPHnzZMh5Q1Puu0TFzz2KKb6OV68Eb5Ny/5UCquNCzoI
cxliELZJxZg6g+1oCB0sA3yJwOHiZy1F/9DGevWaW/MaHDfMs00IF3cRCoWRw8yL
QA/+xsBTtYkZqrPFIUUQEZqQZwach4a5R6N9FolZSYVQNKZx4kLDc09F+slWb/11
TQTEcHDqg3WQUaXlSi31VAR05Sfm6kHWXkDQJszK4NTokaFhBJxjIB4CRsrLnxZh
TGDslbwcPIJ80L/rcT/f/x168iKAO7auPKDa+gT9JlnraxMRSe64fq3TBCRBZYoa
VOkNv+rJQba7tiEFwUHfzp+J4R5UjVnxSG4VK20UB09fIFRox1I3FdQDoBlP3PAN
6hQaA8MMNiPAyfPnHSCQg/r07u/oym50N9H8wEKvlZESFyzMEHkCXT9S0Dy0EjC+
ahRYADOV7AMWbgu9/p4KSbjyrCPf2182cZSJ5MPSW08NDPbyczSZK2KK15jXPgWm
+6oP5eA09g9bdCNUc1paviBnJBMiQF6+guhiWE7Q89YYIWzVNEYy5swuFXFJB8KL
ID0yJjbQY1ZjNOCo5PsK5NOfKoTFY/4xOlhsAbDcJ7GvAjVB71HuPDmqjo44/j0a
x2dpxNhWAVpi/okUt6kUyC4iNPufV+c2CLgVsOD3JV5R0TfREgM7toG3xlEQIWaw
SWwX5sD81+3a0pYc1+1/t6LZtIoRNNNk2XOAkOSnHJ9Z1/jgJh4vxfdUWdXvAf/P
iIyhuKstR/3Tqr5tBSMYv5QSKGZrsXIy5NcTQSaQVTDGgqq+eucOfGCCfKIt5Wdp
k7ABy1queR5lv6a0peOnytTybIb9aYmH9V8U7IptDW88vKxfvZsKEH/55CjXd8tn
UkOCBZxDnR7AAzzJT4wq1yQoJV4GWroPK0iga6wXCVZ07KzlurH2Oj0RHosB5AQ8
zqcb26Aeb/KDLtK2OsJdCLUsM6Pt1vvduOQrLqNzQtYMQb1Q9L8wEvWKmKViD122
pd6Yrg/j5dxxtkzyFxt4IkUSoTmcHSh7gtTZ/VFJ+MpAFwuULRXjvZcs3eIvMtHl
e5wPng4R3jWyASe/3ZfW6wkx/AcJWw81vaT0a+bYgsLX6mOWpxlBden5TwaWDwBu
jsZZDB04jnnzbc7q5pz2gg2FLNx4RpX+OqkQ6b5tev+u7jUriI2nqRpVPqLRAKKm
cAXGWncZYrSx1CoFclyIeSObNNuadtT/8d7AbEhkEOlSNoWfp2AesAmrCWJPpY+H
p21Vybmd734x24gdpo3h+owuZQHj5r7hj+L8E6U79eqWr/JHphhcZdJC72h/CwVh
YnPOZjy/Bxizemrghj6TzPMQYaQ3ABHLV36yFYMkqP2+EsOm7qwYqtl1GGg8dx0P
EzofDrODI2Qmm/4AW370MQcronLseOgEWlFqvAu6mquZ7+NDyAdJtEZRdXL6oL9v
Kw8rMkpkzBgRcDP8z+E7C5QaxbCm1x1isPjDA4Ymx+apWYmHXhH4akblT7YP5cju
D2PG2VsGZzr8h7bZgHuqYHJGZldohvEx68hhtiuoyROGXAXPNvRXPKch6VesA6r7
azhcs2bNeS6LHojUFhapYZDojgaVnrBIt9KTKDQt0W7U5v5/qSpPFLpk0o4JbNN/
gNhyan68KH85P+vXuVt0NRyU7Xes5j0oAPbIm3Dr6VNVM7Q95ICAHSlwueX3ImpP
Ckd5kl18pcapOr4yWqw5MN544Ph8RzGI9kmE4NJzCJR251psf6t2n4OhJqykov9o
rEhFEFyBxjaPdFwZW3aRLLhkwmlHOFCxAPZXmBFLdcKBY1745iv98JArNBOhgu2m
AyofYTzT2LVPKoXT2SJ541nId2okDEq9xzHWo0s3msOayp98faUv5P60zPukfNsj
BEO9qWFwq11u+f6nZFLxDp0L8dtONUTHz87WdSu/2JnjnIvx30e3L/QSoXqCK82K
i8oUXde9Apb+Px7d8IneexbYOX6nLkWJ4igUFrRe+Bx+DHa57KD1BRlKVQgbhrdG
LHd6I0vdJC2FIOq4kuf+KvuaX7+jBSRw/GSgkpn2M731EPIZ709+XFr2uaTijM8R
2MSmaBjgZbGu37eV6HUC2HkazS5ty3q60C+hb8Ld5ZHN2OIFWw+/vvY47wscE2t2
FtlJ/X9HN15YQgswVeHMKYJEbTzfsi8UPM/5AJUP5TkHDPk5cvzfkLwRVlZB2d9p
H4uZFcneL1A/dR9mAwF0SubtPKEu0s03dIyP2cY2C1y3kwCtVFQZKsQDQ89uVkgG
oE586n4OlOk4ll95rQAke9oMm25jB+hO8tf4Bcs136ZdUutsf7R2K8F0CBS0LWDq
m9WDIITf2RNNbn8hwJ1ACnTySSO1XmD8UeyYKw1/B6kzjkjmb/CzBeOY51rWyH4r
IGMGwPWmDM9/H71B3T8lN6PFlhmAJGCXca/8ayvyXEHLof3g6x0kgApxWQNxaTsV
RZkz2rmFbj/PoajVNDCSZxeJEh97SUoHs3w5CqXUVRWs70Q58wFue7L0uwkcXTgS
xz9vwWT0kO0qnCwWR7l/mSDMnVqFTRmB9Jp8gaJmYTXR+mdkVYwBSOOXXBjuxEJc
8Cd1sE/ZVwh3dGXOc5eR6HEb9lTbcckHwsiQzbYUgOF/Wb4Ucmpjbc6EdodU7WUv
llKHLnRVJ10Z6Qq5OO8RF9KSEyz2/4z3tjmi9eIRQntv8BDDnKNUn5FtmleFDRuv
MoQic9v56j3B6Zxu8rkmO95mzQzRMmebXCQpP9QIHuFm9q3uIZ1G0TZIwt9z4BIC
2Z9dtdvpW97W/57jyv9PQ5vgRVT6d030lVTPkCO207TPdwLfl069Ks+9KX0OR/nI
E2/QmwqnUQ2uo8WNSaUvim1zXHVKqErtKDJW1haN/Od4/dlhPlqCUsOFWO1BnCNO
rlkspxxJMHFaFo0e3hLBXvHsY0zBH3RnlG7Tj9Wt2H7TVCkKl1ISXF++VVuOyy8b
x9gdmKe9l5Wjg/K8wv8cGWKzBjH+fS597E+fdu3BpZbtP7z8YdGkaq2MV7U0/w+j
rTXWFL6ADlpjR9G2a9qMD5cuRMMPt7Ym8ZxhKiWzhQOLloeWvX3oO3UpEirAvmKP
PUQKVrqGk2MzhkMAFUS6G6mRbvsgwNXSLjTPPyIP5kwY9KMc+AhhIJcxStvWMwD/
3+na66Qzb1DpyHn4tV5NITRxyJ8033O9QbkcjkIcFMEKQA4IutfMbeKcQzKQmdzX
caE47iUp3hGC3e9bmM8fwRRQ7/gTQcQ+KMzfrzuT80npvZYDZdzaAu6MXuQOQFB+
`protect END_PROTECTED
