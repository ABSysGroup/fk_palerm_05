`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YWnpxgO3FQo0cFPS+VHyiyRNGbQnTA47cKLM9hQmVSI5f690fqJSe0jMHx27wq/m
auQaKUmglZhldOG8qQ8nspea2NdRKzXwvgu6BvR5+XWX0nc/v6tKeal5r2TAvpUY
61YO3gdxaWSmVZwE5L+oHYOmL2RDXuq9IgRSLkRvG+rR0geWaAQt/3kRSGZdOu0u
LRb5zh4tvFdKehqAek8DsTQuO0cnUJimEFTpI4cr6paP08S9y1yEoj1f25hMfHfi
mMmSXKd7grfGX/hR9uYS4v4K9DEenMeCnhN4Z7/XDShIf/zmvnM27oci6T5K3atc
pQlLxbi2tNUF1J1HWAd8iU0IsFbTt4f0Mem+kyvVoZ0tK7KMcIK8R8gt1eeqRm+u
HN/X9sgo1tTlAqPYdI82Qte07J6EVQ+EZLcrG95/wZmrlGYAeE4A6ljIQDU8cvn+
JgTHCYjU7UAlyM8GmygNaxoQVgnpHj/rGGcOA0Pzr8PH+f5uTvn6NT9yMQ2k8e6l
NtUvBPmSyNLp3bNgVZpmMO+/ZPMNUvY4MQZ6ZPlvZYz5KBxDMvJGVEFzNz578hCw
3W3OCHwhPtkSEtEL5pXJFWxLVDsI+r8HGT0a/wUG4zm9BT3KsWBdvnUoz4hPuaEh
XLN7O7DUdhx2xvasbI6OJAD1obOtV9Wdx1m5zuN108We7pE0E3wTVoVXdSUyFn8P
V0JJ1QI28MdJYwNzb6kV78EkoKP8CDlZ4FbCEvrxtajVZfvXpmX52U6GbFQp/C6s
BUOzxeoENrv1FN9hRhiwbkbqpqlX6yky//qLZ15oefqPtJNW78OT2S3tA5FkMUW6
qrvJpGTn6TOMWDA6nytaRxtidPi4EvkQI+m9uLQRKq7VphSz9KA217gdh/+ZSWwF
5Z1kQDAyroxqiaU/sKpyL4tNmtewHNISNe/+fiuKqEp6t4GcfMGd+TVBcTeJm0Sw
M79kMsxNTxvPM0ft/VjROf7juegsqKgX5poMy3NSh9m6I1t7w+Q73ISik26K4khT
jbi0MuGgiGfRQyUTq0qWAgX/vpRHOpjY0+3pt1bjibJ/K6WTZVQW/ySD0iE4iOYT
en4nIuU2iqpfwSEBi2xi8xuFkim3fnB8fgy8o4KaVUtiUITdjvKW2StEMgOx43A5
/Kg+kcPOthVk4RvRwlynwemqJ1ifQdX88aNz5tUK98G2mBbbvzu9zytOH6yfnZak
ZEnum8sxabJh3kvAON3rT7v2SlzN0AOzIKNg0hY5qA1QJ5lV5jKlcmBHb4UaWl5e
5H9qD9+Wxel4JC8hgpctqU2sk0XgGYtK/KL/e8yP/N3Z2XU+/Jd2H5WMXUrpANof
+D9DHj9B7uYGLn86MjCU8PnuSyKLd8TxqRF0LHh1lLD9E5PudY0RykqyFm7cqCrp
DPJPCj7J+nztB4y1l1UsLDJ+2T68DgBC7rCJrAru45sKRur71BpVE9DmYSx2OTRz
MoIl8qFIHeX6bXYk6M0XqDjP30jqnhB3F5NRnCoKEANU/eXFBjlSn8ZqX4JXPBzy
fTdt/M2eoHVa6j2gQi234fZ6sMgEuQESIthL8GfzaKU2+GT+cB+4mETsZ4momcgf
vpsuR0o//CAsjlcolPwDkUBAzGR9W8LSu2u7qhD86JR0fad0hnoHX5E6ReP9/Z1J
XsF3/A6cB+O7RWS2xZPQoIR7LkurJtQFOsU8io2acacVGrlFepXE1h4vo6yGBxlM
CjWppCpRtQZeVlU/bNhLee+2V7jku4pVmVQtkfnlBzcynnMlTJzSf8Di0uCGzA9m
dmn8qVk1Tdk0XNAlX9aXtF8t6/52mLFuXWnBjW7tFmLiuDs1gd5+sN944s6HqfSz
IGbXFvSNGBOZXdnNI+PTTEsv40xO4wvCOdb4CqVqcOn2h7qe+bMoLamRceooysJQ
NfjGdi5lajQ+N4zSTYUGsFPt/m5WGSf3jPnnvT3uEleEGzi2w0+C/jmVqOqaESuF
QFvFP3zPHTMGZduwc68kQfVRYKQEpPv4AgAVrQ6T6t0uPMpiubHhhBEs4obh5ps7
0xzGu0nujarogLf3iURSydpG41D0r6p0Jplve4yqm2t+LrCtgiyrh58tKncDWiEz
kqpx0sJ4G3XLlAaRMnTxnY/n5hI1GFkBmDXD4/kbPZewvupS2mC732hK4ozRTYPc
x6ZUyIkNsoJs1QzINhJCmMAc2hppYG1fD+ZP+0sVOAvpIgB1asu3crwR6LhWFUIY
Eq8qRthyKM/19mj+bd3VVQSnfIrG8lf1dwIN1zX33CiUSjLyaU8dfZi7NGJ5Z1ED
UoGkbItI0F0UkcYI9HY3q+fVL4yOHX7QsCRd2YojxCNvfSfcVt+gZydvFAoYTSah
A/AvvEOujkN73ScKX7L1P5M6p8yvJ1xHj9JxBreZDMnmRUTEyOclKI/5h2Wh0+4k
ZsaF9mQ+GUa1ujvG6KeVE9Sq14agqEltHVXRf6P/Pg+lM2jQjcmIP0wZBzcxyjEG
hIduypcIjBIOnxAc/7tPV0jrksnoC8VUqf0MGArblKjhYSSNXvXm21D0FJ56962M
DTjZbHVQsrweXq6fT6GON8+642+fO3KC7xdNLj7Oco0h9822HTFaTIPncMsRAtsj
OnnoUrc+c5Nxzb4FVd9iW2qOuQYt/PIbEmz0CZYUh+onOtmLWrAVW7EyyDqAe6Rt
aShUtt41bx+fzxEDDZsgXuXHSQuoO2lPS/12FrrALCQF66S38PMmzZXInr3on12Q
ylYueaVamwznBpIU93WhJSMYUiRUZ8m0pn6rlU9ndead36Io0mfnL/JVWy6jTW1e
Y5DKi57IF/5cckbkXbD4Cj+DFjCwCAOzmMyS/R14NuK3QHjCH3iYfNbw5mjn6Rxv
hJ+XOrWYCdHx25RYhd6HBTt/Y65cYpVKBrFHcjQHND+rfVh66wuy8vZo9LCB3CK6
iDI4vADUgWDw2knTAHWzadjyl8HAzO74o+trC8z6wRu8J3WHcJ5bSB1PkcpGkmF3
uRPWgqlfp35kQOcVCI39LYH8tsVgy8U7Q5CFmlW7Xb+28JgmsxRg7hugAJvcaxvD
Ddo3pN6JiznVCjEyrjB8z8P590XFdObAsJbXJW1oTDOYDtjQaELXcdXNwvu16mOl
QbEXrm7sZySITquxtF+AgeoNMEOZgBN/Abos0N+HwhEHocgeLE5GZW9UKJs8XSN0
gDMXHIjPTde2uThkT+PVvhgWtKWsSrT66rpbvm4u6PFbGmlpJE7NDUShrf/gLLe7
N/4NJKEWUybedLpFg3X4XyC0pyR43ZwnosCls9DTg6faK+qx9Ga1+NLo4M8mrFTl
5NaCFNGceybMJvOE12MwaWiKxXwxBZ6zHc8U4bRCfaf3EHfhLp2JoJdCtT8dfftm
yPhMWfe/lapvNgG1cDIDWV/EO9lLKzud6Tb/tu7m3ADvaYEq3uEV167VcDDCZ4Xj
tUKy333DYs9j6hrBtcM3EDWY0EQEylGqG/ZsswTotuuDrc8sDRijX6v04MdgIyIR
ISa3RoYnTHf8IzzA+w8U7zrhaU8lckvXAXzWaGKn/mflXLzoMExG0LtKH9Qv9Yl5
VbyTTOBXPuuEDxgqWeUkisJfSchgPcLrk5v3VxR/6tH1TO2YA5/vgufrcBSHCXDB
MBCJ7CdguOyW+vjvdKOWlKG/AbY8aFu3wLKVn5/9ZQHhWgR6OIjTuf8Q8ZF9u2g4
I15uNDLggexIiXFTvv86upuZLxcfWG1J6xTdiGSsRhW6lpZJJNJcprBNCxG5jO9M
XsW57NdVtr1BQE48wtuH/OXVbg3T/WoN1D20FYvCk9mmyh8hUeRhJkNtPDM6WE7k
1QDR5quZXdlcCwic4OTjFJhzYU9JvOMCKiSnBvAypuDriU00QZMUQlG1X7uc5Ktm
oowuag5Q6IZUDKK/7jOVGvCjs/dHkZKs1chP6m9GUCh/5QJ4PpnWhJ/MX/74ynDu
xuyo3lgSXKCIe0oAU3X8wVIs15oAaaJt94pac3uQoTqlqtJNFcR/EvDNXPM693LP
S9E+TaztGzHSrYHVy6gBCTpx1vOq852I9Xogsm8KRsMJ5WMUNDlL1qV/f70RF4lK
cmsFmpdDtozxjqp4nvothQ20deNRSG/hqSt75LCg4q8HVS+pGNXBvqPwnZlXBH9N
lODnMLZ54JK4cxC0+Wl1lVf44Snv4T8ZBn7dfBngEXiBI13OPz/of3bfKs3MtXYa
vmRm2OHgx6D4CO+hQQL/36RaeapDwfrWbtYh8S/X5Fyxf1M+IdOc9b1Z+nXCSPBN
p6Xk0vwKUdyTCibA/FFY3UGHW9MqnVFASZlwofUCrRP+tN7VvYgs8acquS+03Wco
Y1zDSDDntaNPuEz8YcU5x8vWtEZSm/kpMOFWK2QvhocexTbdc7VgbzvZA0agZp2a
z2bRqOsaccfzm3+PZJaRho19tq0qDgEWtwqzskps2EdEYRB6LZHvZbQU9nPrsi07
mH5Ymbn+nLHqp5cR/X5m9y41DDF0JkwzASzgSAiZA/HOGPXR4+7tngcAUV+opM5r
mTMTvTOlMPoMsQH2aDo9uoBPqH2x44Occ0y+jWiBWY/iK3fY2dX/nXZ8RB7dz6cc
QZCsibsd8+lrHX3ylPcP7sbNtf3eTdw0WKYb1CXg3KAGvb+sg4yEMRSy+hTbqZJk
R+beJ7SlHOuh4iGbbz6ONCaaqiX/35hzgvdtFw9tZGvQeWMpGWvWtgVazvPhcuqt
568E2YxmCNS6m1fGwpu8S7QFkdo8BR+zS8jbR5vCU3QwVaAJy70ttDUvy6/aGXjt
2ARlAIsmQfzLwseZn8Qy3zhLS7A0ujU1PXW7lAk1CwabrChkyGzb0+h+7G0d9Z72
buFIQzqKT59vwiVpYAPpmA0zGMOs4Y/0iBeVZmKGy+wjx3+zyQqkXejgSyQri11f
bDg1o102kBep6PsgJz7gWiX6Rqk2p5WfJ9wcz/KKKQhc5lafjy7SBLAhYdPB+rp2
zjg+Xh9SSFRspDzCbpoM0BVr6iPs9MVbbBb2d5MTFgP6hK+GcdtZ39tpGQM5Kq1Q
iLRKKPkNpBG/afXnj+Lkg4PqJphmu8jMrqwRp3S9IA/vLPhnCzweFb6n7cBhBTsH
xhYaf0UWnrhZggRmIV1psJqvT5FPl02SzQiYs8hEe2RjZxPPDx358PPHgPPwIqqL
54v41HICNPusZzhnB5D39yPT5vjv9km31/UDRPpvs+8b4jNRfR7Q5uatdVXrzjv6
DE3IAlX9hf8fZxRQzVT6blZ1y572ZaqFPge5VM/1rZ6KUJlzIXsg6q75Rbd6EMxe
MUmmvWQ7X0FfXBGoK585zwIZHrlrJUuSWWrPmLi38tSqipQpI9DEYHzQ/FsR2EJk
WudhxxHP8plnItioP8yGSYcOM2WmZqB9V0ZLgM1tjf8LkYmmYoAbGmvq61QeZGg2
aO5i0f2pPLltfW0zCPg7rp2O0A86CWqe1VczWpswwX5iojkPO5hjCMTy8naxYpcF
7cu2N67C/hIe+t/TheJoe3HN6JsNXOAE41//OAplUEeSpBnK4KjHPt7YUK3XNFTf
IEkW9CzAE+j5oLOMvqrvto35WxFy1gY4uY0XP9uVQyvqw3IC4J/JFq7+QI3btoxR
c0uqWiLzX1Ox4KRGWavF3x25ZXwa4CVZzyowB/7cGrwur2xy4RewE/1sgqxU9W3c
FDwqKZDsDkJ7J+MHSQHy0HXP/comi0jRr7abxpzLPs6hSSR7mA6cfhLTCjKbowHS
SAnH5GQy8AoVnBsiSOMZRNCSavJmjCdGrTR4Q68Z45SKocZsgHrZYfORe6kB6iJi
0gZn4Ex8XLyHrDaeFp/2VeDytJ50gG5jCjo+R/P7afkccuhGmazpG0o5e64YgFqA
BEFB2IhcyGr7/Fp33lVVw+J1D88P8RZuyl+xgITdJqxQeKEXn8J1Y0NMDJd1q7i0
cJ3lnNLp7jRb9zE1Uv5MbSDSerTsFNnGbpv9MRjnbT02ValZ1QqQC4+vFAG5bpk6
LPWhYcqX663RTZ4JEXdiv+P4VX2K0fYerKVwX3fcrDlZGHiyyixzMLpxzS5y5g8Y
gb+GzXmw3vJ4x6rLQkVT3EUBtiOsaUXNFqfUPDCPZPfkM6rro81XM3V/sejhg1AK
rbskbAUtSjJko7c82OuYq3RpN8vSDI6c/qTnJc3rU7Kmgk5jTgMAj0UgdrJXOuBx
KVXA0A4yUT13VBFPdHVGp/8CLNcomKqXQhdaJr29p+odcjKsWrd35Z5UYAMbmAgU
R1CuLtuCGrLAP/Wug5NMwJPoU/5MpXqT9fUxVeb0NAhN48bbQNx59HpdUsiQDd2Z
Nh5iIiHxYTj3LHniW7I6Zbr86ALAytlpNJ/wheqG9051em8dwxTFjRixJjz3Ac69
2/rTK7UaK9lbCtux7M0KSSmrSJfhslJUILzmNflMrBynHx0cNOYdFwg3RMI81Go3
tGyzH/Fh4q+w70dBa4eAPV5xyLBbXk06zXOhzeQwgP9UneLVN+s78FpC508QHY7K
KjYo2huZ/6kMX8+OottkxEH25itIXIQ9PHvVaiUVOJdpCXXiFRUr4Bp9KU5KIyoT
0JcP0qZIkM+4yJrqzrfXR3d8H5hxSNNEp+mw6ymCAcBiKKGiYssD+Khn5/aNTk0E
0rX/5OEkB/3Hz1IypWYmWUCyq53ojMeyNrt2Vsxtz+ekcK6mQlhszsUqjUXJ+X59
a4CuxE0gMaYn/D79PPsuftdCjmsvlzK3cVV4hf7K8ipOgJIAdXGs+8Al3aS5GVBP
hJiSrpEnxNtAuexocQvSDrL9C1ah5RlqtYIURM5EUQeWzbGCX8YMwcmVQrmJlR2V
1ewHrKqY7yv51vPxotrDkSSEVJgqF4yvadok10uYLB0RhWWgqldLGMDrMt62kTcN
PFa1Mn29QrWWFC5igBaV4EqofLRvhkmSowXce4SdSNG/1MpAZb7b6GTgQQNAiZU9
+qWW4W4/1AXisQ9I2s+GjI9AuYVkAuB8iFkEf4/FDGofOnTxSd0nrWHAM9I42Otu
lVctmrAuzvxEciYxhHfLdIfQerkgx1+2zc1udxPzgsL644Nfw7MQRviHl0GVYkuk
h9DwKzWWyQFbqGpjYm9hSLulk2/bfrf3rWYspY3G2lggyrqTKgaIV2HJ8a1USYbb
R4UJlxmNbdXlI9hlgeEg+cnKFHtksNUIvGuJgnNPHgnfyZEUlFhF578e+3VjUeHU
pDhUKuYAVTd0OVSaBUpzK+PuiqMIACqZhSp0ghrjSdlxmtrEZfal43RdNzACD/Id
vglaLOdl9EHr6tUgw2oK6oIncs399CYQoJ+dkFYgzdzo87NFqYCqexrE1JuGR2Sz
rvzGzO9eeGnJfcL3IsUvCY4advjGnKqdunbK40z++FMulXc78fhV/kk1C/uUYQgN
Fd1DiiI/Gv9nwn1lgHZe5pSNwhTVkttPCWgPe3rJ46NU1XEU5ovX2lyf6IIUOaKM
F0WE0pmwD+N4uRa3kFGvCLnMVpLjuMjDxHz2hoQqX3xvB3iS2XOzJ5hKvirFe5/4
hfgVQXh9/EZkzwhgRA6fLRa6wejPAbtbGUiIZQ9Q9F9XXH5VcFzvF7GZKEc4EWsP
Dp3ffb2XBi8qkBk/yqGtc7TulH1AcD1SeB/w7SQ3GdLpcf+iNmIbRQ3Iq6BG80sW
39ShUzKD2IsvZ0NVfHeI/wA4oW99WKRgrbVjkCOXA0vQ/zIsgd1vRivJTenolgDb
78OQKlau/yKux/SSW7Jgueq5PZbeF7dh/QlobJL9fGMzgCtAdaCUMc5dTz7gug0W
kc9FolfrkXlc6W3ubmumK5u/DLZcjb2aT6SnyZp9XQT3M1c/rsuH61l1uzrXqI1a
1mfcGTZHVVodvqDuWhTcHw/nS+GJ0Fb8ZrOZ0PecNpat0o4NVgWITijIs3etpBY5
pyojgWI3un04z0cv+47lPDcaDAwwtKdU7WDgP3OKC8XvjFkod7YAOPwV7022rL4k
NCGoSA9ZTdfs4D8hJ1v5NJJNHC7602Q4aDGDM5UcYeI3FxGMGuEVehaPazahFr77
OpcikwnwUP12vr/Nt5zplAL3pfGNdBTXQJEiXs5nh+Y=
`protect END_PROTECTED
