`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tlFUYesblrZ4UJaXo9nA5PRE1pZYyZNkrEdA9mefxBMevhNrGlyX2sS2NZA0iiAo
7wmhZOErzwPKFFCEijS09DWjbb9jlQHWm9n7Q28M/M+UduT5Tq1l7pvsqUYkLe0A
sT59tV1cw/AfHRuqGDYq59gWES0wujSKC1Q/Zfi+kMdB+G8pNwgSGxr3ZpgPct98
cBsgoFd7lvtbMg7goOZhvkroyanSbd2FY4ubd0BMKZ5SphwvHsX5Xdy5Kpd7n4mE
dGN6Yv2wEhIezYx5GiB/KXYf7rZVwTVnwsj65+DIyNJvLepUF3+I0H4dJsZnqPsH
CNlU6EUuZDCTxquyFi+Bl4joGdWJPe38LnWO+MvnEo+ugskeoTMWIF280GiqpWRN
jT/S2+gEVE+bwymMoyGY5A==
`protect END_PROTECTED
