`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KNOjBPW9d3BHUc6vZx9QgK5o93JEc4yXry1MAAzMHXuKqis1QxdaS1UVJ6tal+MF
+YrV4MJqowSQx9adeSHJAQ64bmVaA1/UtFzJpZmnMKzgCu7iqKLTgRAkxPdDQEw+
RQAML4IbzVuDw9qOfd31OgykwAeiuFI3lfByGU+AwXyZNusOJu/WuCATGfwqJOdA
XnK5GutOcnpvPNzoiPLqNB/QwoB7V6ybRbA8Ohz2PmAsjjDfklZtoILRNOSKxX2O
j1BFPB6hUzVx2lDIQMHa35H4/a4BIGJOCMFkUUYNGwu47LIthyk9LUZ4MpvX56Nh
CsPMQp70BoCATHR5X1wjvkRMYYLtCSEiEms79XQuPT7K1PDHXvn3xbKVTG+HoK/L
o+7+MZSW4K/P0Z5QJH8RR4B/xxJ1pVRL6u/2M1z5GU9Kk4Sf1mWn29fWagsxsHNW
sMPcry9/OeYkjUIT9ztfXGx1BSd4yzCVK+KsClM6FMs8NR9h1BKI7WFkUzG/8F8W
jRrGEiC0scuF+KDX2OoAynR7TuQ2Ls3pdxUZsEaPP1xx2pUzf6rqVvwaLq0JZfbR
kjdxMtleEnb3PQL0LXTOMCxmgaRpUcaa3tLExf95MSd2BnFOTy9jlVY25whUdROO
G31lWOr7p2I1WmgUGX+PEM0QlT9hxsj+1WaBhyU56BRHiJEdq4ViDie8FfYZ969u
v8QCBujMg+46y8d19YO1s6yBxjxpm59c/NPkSO75VpkADcriB+xqBxd9ez+WvkMt
7Nn61tw3nLHRw4IzkUPyZnd8iJr5dy19WZ4EIz0fgMSmK7nkDaciy7Ew2RDoF+IE
mTzMRoktL+KxpTmUdTYu9KRIvx3gWoxTuz1yTUgAlk2YOLpUfQHQIfALrbM3jPw2
xaxL9z8AXQmbe4MKKSU4OpXiU8Qy42+86dJrmMf8Lwtq4dmE+aTY6XHpiyUe/u2W
ifnVV7G5EHDr8Jn8eXGYtSPEzdJVq8qWsJUF2hFLtK4BqRb8FtPxVocUlB+uqteD
RRyvT64aFikk6KV5PuKC3er0zsyj2nffZ4gZ/5hUqUJyHn4Y2pK1py6IRg8nfu66
8wlRKjJxOo1suMAxN8mLD0AGInBF89Z/6A7p4GjkiLWbFvzw+uqm3G4BxbQUMiVn
JWilxdy/OoAK/P+xz5Oc42OSc7Tlkml9Qx2BFTb1lryJCLlE2pt8Vp0Fhy302YXb
qoISSOIUYTNkRlrbVX6ap2q3REvX8whhmRc7jVGS9Q+Io5XjtizR7E3y7CCHzQjg
pmaWKzlSCTfkKMmChK1biJKa30LKpLNBjaea5h3PMjBzC7bi8PH8s2H1qLQo/m8I
mUcAxXFX6aAlU+d21QEeq2pUjxdrLP4VnijfTNbe3ERQWO8VOKBCJI4BWLsI2nxt
W1g1jHCL3ONINd0uNT7q1UE9wsciPIUk2fzyC0gWDaDMfWM6JkSvVTtjoJvkW0as
GqwZZ1rJSt3FYdo8+9upzMWwapQJfAbdPUVCtWgNzjOaibwH1gIla64moSHncvfR
phhk/q+vy/RPuAPiGdjXkHM2XT64bO8XovG1epXXvuubLy7X9uiwUYppcTE4BSxk
mNIH6HxuL8tjEzGWSVWTUH7tLm89lt85s5Dth3fZnCS+Rbk8QNhm98TpVG+wNNF8
ea5p/1XchpYv/Is1HJfMO6S2kpTm9jv4/j6fJWJCIhLY0Yo67mpOgAYmEVQb5yCW
vkJFM5JVxaNUJe0UbTb2SJKMYk9bHb7mabgnGhPMPT/kRJx9diP9h5mcBlbtCABO
i2t9shacJjdzNoFxoa7n5jTQP9fe2+zg4I6JzJWjrnZoJWr6J6aPny2wcG9lWbKw
hweb2epTbMnAKySffVevSboqc3j7383VUPBlLgWIxW6H5pJ4HfOb3ypHeoGMswep
OP8ooi81yBzHF72feRtZ85dfzomlq0+lR0gC2+YgLkbq2W+lPe4zx+PxK00MY8ER
UqmMGsMdI/A1XjDszAreAvn9mImYywrowt5AauIFOiK4x8e46CNYoBunPQkSK6Oz
ArXWa6JYvQzWelz7ZQO+f9mT8I+9EDfKOKdNhJ2sQQYapNanspvjzBbLuvEHOroX
DdCpNTrazqlNDlw0hbIWCLSuOjDWX0ubPfbK9lUeqS5QJjYCjafmt1K5RrqezwET
3/ZKKkt++bP3LYHck5wacnOu149dN8utRGO+mQrJ11FGTSMEC12aFg23ghiKbDXG
cIiRW16TYwv8kd7HxTiyl9HVUm/zik/GFumjivMZQ1F/9cWF41Dh/WdAneQT0C+/
9Uxub8S+Ky18AprJyhXvev3Bts65fiC6XCEMyspEfgYBP7rVi6tmCIcsKirKbb8M
rUIhobXOL7G69t+sNHLzGvkEJatWiwdsViLYDSaS6Xlqi46cIU7A9W80g57sysuW
rZpFv3i5Ba8WsSz32hP+5nws31PNorUiFXV93xY1LHjLCZcCZSem9teLXGBCqBjn
hI+Boowmxrxjsz5lV/cBsIGMknPMx9n0QuSjcDqGq5E9Xy7Bs8+dM5hkmYxMa982
/rVItEwZtnm254gWmhnaHPkD5bKxQs+9SStHSydjQsBPQHYxKuf+mWE7Cw096FGE
/xrC9U/Zkfb/50oLcqS5gySJnvXqtCVbm9tvwE2y2aMdpmIP0zQV0McIaG09aMK4
Cnb4cLNbJYRavUrvgly0IQA2+EgVZG7Ifroei3wAE0FQn7DrW4Im4IN+oLolDD0a
jLq18i/b4XhwImpdevAL9TNiGa9yBf3or2xVyFx16WDAdgjV0OB+M6md2Rjz9z72
kd4VrX0vmL9STkj8yc2PKHCRwg9EEM9U9K02cWv7NVfWJbtwi9m7Aq9s8ITe/pMB
tygvBP30WaP88gaRSiHrPSsF4uH+4vGb71GEYNjjr5dpUd4SQa0jRSmQFvPK0/+d
dqg3lTGseP3AHlKx0y++GzAollPKQcTve/iQw9UktLB9IGH0aXdloLvkE3WNCjJy
aT3pr/FSJFdQZU42fXCGTGIKjuaxirUjGHVS0gGPWssH8JxAT39D93tzbjlUO9A5
LUzDkKNN8SwkHaaCqAIWiglePe0v2ZJWkiulCJ5fKoIJxyHYHKPIYt0PXatGChZj
SkaV8KjBq7SvBnqs1YX6U2/UrE1qg8Hi1iiKoS4GtcHhk1nUiNi2xTNeWz0Jr3NJ
VbL2htqOQ1l9lguT+EJ9ooCXncHCnpEeaFJM9nviD/l8NDTQ+7tuyMlSOc8iOF++
XyOzUfsuRDSaZq4/Q8HrCyxkgc7FIF1+MTuXO2zkoq7GZTQ1y5BS/S+HAsFQVKTP
Ax0vComQClE4sm5nnEiBTvReON9N0YvC69q2WnWCN1PVo/Swj+TeXRVEQGMaxO8v
rOr0isTzjLeJGnFaPz3CdA9ebbsVw/6BGn/XGuM5LW1FtJi5BKT0FYD2JMyV3ZcP
xARE7H2U8UBUJOnp1ElZSArUjTffeNr/wS8NkanddfYFF0z54cL5YGjvQ9kJ4h80
qrDcmvyB0eqIGc4LNrQNezeHS4P4rOW+o6F58+rHAj7GjE/cVH+iF7AJ9Jc8lUNU
UA23A52FfxcSaN2KqsSiSo3vv2yXB4G2iewrICm+3rO84IuLsMOz2SF1+quT6ZLG
muoOAtyN/jOlgBRsWunNvtnQX9fVzT1+jSAsh6k2HglDNYCJbyWu8Qn+mCGBruQE
11LcRJPxq+/+MGLrJfkuuKtq6FNyk6CTF0eSgoGa/R5b5fQmRuZNK/snm74UAeEc
cx3CD5mtWhRiebr0mffpd3vjLL+0glo8otIlqetazt6yY5AhbF866eFm6YuXuPsG
NnFxBcMr0aZYr93uu/sD2aev5Bs+NjGHnLHhYNdvmDw/vsMM1z9lHpNUkCSKemyO
y7u6Fx3Y1unZ+21FP7+z/q6rg6i2vAlI5RTGaOEKW4/lpLHw6o2klI7HAf0WLKd2
GIjPCTJpd0VjNcaa0/4/y2pi8A2iap3Y/ozysy5TY56So0O6oCyX7RBX0Z+EMXuf
6tmW4lsANPuMc3q0UQOT/IvHJYnHEQkrMKMevFFVVbO4/oP9j4wG7lREwvEe/sXs
hxY0zInwCdMi3BxPSNsGoCgrHB6DiEikTiPaYDHveBtAMscbAqIOFdrOP3CnX3qj
YAQKNr+Es7ii8O26UJbW9IxsFn6fsGDKlYKG547IpPYPPTbOgA7ssRqPDR/YxJni
/F0TmxXo2lIAVfiGaNEOTufptLrbvrGKoqaRUH3SYxpsewF5mPB7OAANLATIN022
UyVz6mc8rL1YY5d8aY9bY6mwZZ0GCBUrHH9TLDh61ERce0BUEE23+AXfn5NUaLzJ
r/M0w3EcI9ms2Ub0hC5L8iHuK3DazSR4fOLlBqflhrIpUZ9qGy9oMvOusqQOKfuR
XJOROtTEAq29FLkVFj3tPN7bn5pwFHwC6c2+tS993Tn41GfpJmoe5ejwwaZBVIWv
SETRcn2CWUN4qxFRWuZaiq2rgoBHhVS1P7QkmX3Jgb/83vZVh4T5a/8o5ZwE50fQ
19GTsWvCLV4lTp+r3SodKCrRkKR9+NiIet6ydHpf8TB7iBfW/hund+5wb3uoaoGt
IfSTp6eUv8uVFjfPkcO/+DYloSqbGPD2TYsYJBxhsMlLdopk7jArpr4gOKa28XWo
3fakVMWmN/PP7+oUS631lJopG0a/THUBm5163YJQzKKY3odVm/H/in2mNchhygrB
UjRbCccWRDenenZcKLdfaOsQPD4vrVadvGUXVm66CGnBL3ayDb0a6hNZx/uleEn3
jih5dKwEQDVlBgFDVbx39IxAvuoRC5z5f8bTbrnefDB4U0Lckmqqr+c8TsfVEALu
nsGKK+P3U+JPSrTUGGwfTuvWpKmcQnvotxXIEFao+YJ3PoQE67GGPipXlezZ2QPT
7j+fiU62BxM11jAB/LEXqWl0/D5sufsfrDUo/FVj2oGWRfwyTJfuc4oWxE7wGUfJ
jsKMpnEFpmiMmGa8pIGCPOfHX1esGMftgiDCDs5OST0MlRvQpJTM2Xgloax3Ngjm
w7x2yNz92FCn1I5tUkIml5QA5DXaGTpKjyEOMwW6k6QqswFbT7YDToALycz8GPCn
eryweZ9e/JthI7vi0CkRdr+xSmza8prnpCq+weXAHXOCQw6CUajk/Z9+8eriRXVV
wnT+qQYFjOhtcdmf3laenD+NRamRg0LF+qTiKDxFYYp9ABeXx9Jh2thm9VgUzVJ9
xBFhea3ZCo72mrWMb7Zt9pRG3xGoCy3tbOw3adLpdYRB6htnVUqqg/AG9W+dPyXo
cyPPjK73gltxh0dwZP8i1DWElXu9U08+FakGuHQmEWlvrHrMjCahHaeB6CpiK8Zi
gbWbq5WJwCNw2iicF51HH1Czy/4PApkl3a2Wv8+Yqw9vPGqUngl9gKl5Y3IpOo25
tVJMA976JhQuKPMRCupBO3WivIO5zb8vdN8r38HXRTs5C1orOjK2kOkoZyO82BQY
usYbvT97qVBnXAWiefrDz0doC00b5pgrJq7quTFUsglTDhQTI11FybsflS90f0lG
8acJaox3Lq649WYowvX+Q2nCtFWMPoMrRZ1OpLYq2h+D3VZLy9StScyifKsypLlh
DxyoVN156dOYtOhMqPQAHMFP8SAXXTeQzKGVoPyJnQVZ54lzjo2Oh3JuZgGVjlVh
s69MBWgLPwSJSGNVw4QkrsxUlta/uiTH2aTug6S86R/h86NIXvfIijXKf8UInQaQ
lPZPueDPVWzwi4SCylWwLzb0Rn2dGZ8g/zxNMtW5ifaF8U073FAOylcP3T1f9wpi
Fze5mNBakRwbgxlkZey+6k94YSTDcGKqlCY5GCmjrrHJYrGwvfbxrdsurh2ae1HQ
u3wHIVWNPO+eAzVxBM8dRJBWPBix1cOe3zajGH4Ymuols377VQy3HpHHwg9Dkst+
9GTsKB3bWAf9OZ/3mC7Cm4rjLsoxpCL6B9pX2AK88kzGmIE0m60NY1J5PiSuv3Zv
IraTRyuC2qn4OoXuUq2bTrNt8SkcbFzSt6BqaVZUGkKoiXd0t/HPGCcvsjV68Kw/
MscGd7MvtTcEh6u/371qyf3Ag0AsFDhv9tUuP0nYjj7mNk6HqOVCnDOyqmV9mnRi
lVVrAZfwBcOwAcMhS9yjqDJQmfazxrbVt5EooHS/2mqjzzyg83kmAxENmT9kwamY
lnCzap0IdjbP2mHcRODB9h7eXOkNUIpE/2gvkNPnrpFncyDWngqoHzTZAbmzYxjN
4IF4u9A7l0ep1vNjGn51q/XT0qWZsxR87dGKiLYjOPSf3HdUNgcHA+diCcRDn/2c
+FpGXiCaxELqTvz8gPHI+dQZTtSRDTMsQQvl39tBrwBNgGYC+vTyiQnKw0JZKiVg
i4LCkY/EJGX1dVn34PMbl3cK9n+SzHTfuVpBArEmEz+q3FnExCmFpb27uHiXUyBI
RpCohqTR2U14bSn9vThMf94Gu6CSWOlz6PqKa3F0sJVj+8ZexZJPcC8v4A3f1Qh5
F3aa5MD6DZBueqtdYlBvQz7CqZdF4Yavhj+5s7uM1IyGGETYwY1HrhdHBs4wjYvm
2T8ni2fElNs7G/ZLihbzq5VuQb3vSkDEzDGn0ASJqNGxzaMtch9Q8wz9jB5XwnFw
isORtqWMUY5vxw/9OFRfGEuKMME+ZEc1WM5L/bB0lChjYRbn5esgK+3tJN+cV+bY
f7Eum1ysFOlpt6r/1vSiseu9Q1K7xypLakE8lg5F0HICdmanirtFB18aJsRseeTk
0Y5YGZgOniJxybMDIBj1/a4kA04rNsPQK6r2LrrN96AgyqB0f75SBCoHCNH5PUJH
3Jc7q3mgH2/bdK93zYjFA1WDW44NSY+3cZ1eVlgHcNcoJvQ6k5jD26zvP1gcgEsa
Z/snP5a+wk4gzMvmFTnXvDAFbKwz5BpUxkgLrL1llS+RQ819rRzYQtz/PnQGp90V
X1RYvZTxQ8DHe83IZPMnrsZDkef6Lzt0TJYjVdHSPE/Vcji6o2LbgBdH1rgTySe6
+l5+5s20WfZC8nIdPLR+Uz7vdvOi9LzqVsbFdg1F9qhMW8rKDSmdN69Q6SiP/EDC
w65Izvg6YzctM8eguHjC4E/xgvkP5PXmXoYovXFEC7Wtq8CYL+dKnGA6P/Auly8c
h+3LRwxdY9m75Mq+7xJEMJsrLaUD7N+Om1GJm29kj8I8cahYCdawehHdLBBF5dSu
SH0+vveSuhEg2fNR6jrZNGPpK5cnr5YT4ZlhE/lOYVJtcU5Gn4yXLvSvbRDIL/3A
TA6yZOQjgTuXsZ7PcAZ6jiY7/KGwFN4GyDJiY7zWOJsZgC6WIHA+jN/bW60Zx73J
XS4HZi/EfMjc7c54tOJNUposyFNpYypFL7HoAXCNDNyvrTE5211wmDPQDOkXiag0
4Zhm9qwz/vDJCf9oeoW0LWLeyu9rxFwFvo6aRcXxBRZ/LGS7XOlYciLek7GofmD/
U4akjWvv5m9MeFYCNwrnmh18LW05eWxkhWKX00/tnJ7UWdhgIamoI+443y7vT2jO
RlU3WD/aVqByt4iuQJ6Jm8fZ8JEva1mXKhXrFQyOa+/YwofXuQlE+H26b0oBOsf+
h2T6KgZ+2NruyvmcnLTcWi1ruF9w3Rrb937jvyJynTaxroo+EqC+7Vym3oFL5sEK
aWH6SMa8tyten5C3Q6wzvoZ+bbCSg/eEGhk5hf7iWwqtVXYw7hd+eCpozxAAmmxf
HXOADMK5dx9iLKMSkdJ1dhF2GjZU62QwVjZHPmUfa6DjkGHzg0iqSMhxU+RoSPgq
2tN5YIjmXqxE1KaLX8exewpi0m740t/rllY0vaC/VBJUO9RNUrle4HNn2MHEts0v
4uKvRmMjapAH8V3pLhpva7xcHgUcu91ekVq6W5tmSEYWjyX3/me9lYy895RYa3om
K3q7O8d0LGLubg15v/RO3ZKlFOyGBCzN60N17FlSTtzQHoVTGBRm7xNPKVKLEyjl
/1IWZyEavgRrK5OY04xoZbJdOMMEzF/qKDERN0Y1mo7KdtoM+eQ1OKxgcPeHi8AV
AbkOGYp2MXv5xIoG+RJkplEUCEOXjs/4BLs4BBZ9IBMGvOBHYrem7zJ0Co4WsfzP
aAYcQ5yMy4PKVY33aCyFxkEWzhJcBY3zxpu11l61o6BoditH242pXfLwl7bryDlo
VwbpEK1H7qidKn6sGykXtM8km5PBw3LALAeXTkAapVCitfjLi+vvWFrIQUWi63L7
gCOC3XLyjUrXeuZ6FSyd2xImW2S7ANgDrxuO4OOqPs0G45KXn3lboqd0CkYl386l
ncE98oTqUQCPvyghopRKpEfVdBhmJVItLXJ9s0821t4=
`protect END_PROTECTED
