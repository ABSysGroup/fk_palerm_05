`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3KP5fh7+1dAHS+QX4EzzQvjcJtBNsCMsupDP7w6C8WmAbXnhCNL4D5VmJAa0rFT4
ImPtIa3rQ7XHMefb3Qqep0WHxeKCIrtTDL4AqYy3jLFNNGy0dL3rZk0SE4aI1tPP
QXhzcP3Sa/mjRj9BEjc5jnQiaGZrCaLHN7wyhX1k7txpYYdRHHdn+1KjM38hUq5z
+2qc0N3IdGP9avgOjyb4mqD8oRomEijRq//na1RZUaPqpCgYQAnCvqHQ1lSyNndQ
FA19euKn0C3gmTm8zO9UKsVMgiEW49NHNN/+Kua4yCYJy8inWWXqm+eL7wC7wQJs
dMw7ClkyVtk4NuQTtM90eO0Dh6UjRChGdX5rL8Jxrn6ee6DeKSFWoP1cEFtU5d19
OgSwKeoDRQxJdU7tkgFK3rm0c9t6/HbY7PIaqbYDvelGx4M8g5Wdo4OYKRTqDgdQ
fv7ct/xDh6PgaJE8EkI93Mm45guaF4Vpt87D5F0zm3HMRFRZqYP5TMQSzTU+Ih5i
Bd8F+1wf0BEA6KfypAS5ItompjJtu6C2LqBiL9ZekEW6zn+F41MgsgxRTGZffoH8
mubcwGIzlYXabTYYdJiZx438oepzNPRf59K19LzOK7tBzggMICgTyDMfoUSPdPPI
YFa4y4CB2w3VjuMvqVjxJ3ZELSzBVgQby7DJSkFip3CCBwQ+JXDxcO7CTb7nizqg
tpXdZyThkLzDdgjfCbhsNT8uVKSNmTYkYm9JxmFPg2UkUVKFBgYZbD3u9of0FMJa
PfbjikNAyp6sPgw1HcAqlCNgqlzJm06Ox7O1sUY1uTZnrZnXE0SyZyWr1cUFrPVC
V1eoEbt3Zfxmip74UayQLV9329NE9uni8mPvYEFQsAR9UW8QjyOdulOGavxoPHoe
NQWvkzqDAaod1LUEdRTTXL/VTpT9VQQRZOe/qBCafG4BjCynRyu3kASGQnddNCN3
nh/Uh8xun99uiaXQpZWUBAMcnggTmJpFZwgZ/1aJ+dPxUgw7ylnkzwU1RitGjeIE
3IcPQ8qdNni6nYJdKSrbZg3ALWuGXKMf6NStY7kXniELKpzNAI/WwWGfMFjpG6CR
HXFiqiFVs7KJJEQvVFDZHqx+S+NmRq3jPaBC/oQA3GSfUXJiJe89clvJWiyWlvdS
QjT89K0mAVpomJ0nD69AqQf8PMMXFYtmCFlM9UO6CD3ZgBwmm36GFyw5TpKbT7px
HhevS5fvbPXJ1v17U3eV37cshYyTyhEIPTdjcnMnPJo/90CDAnj676/uRUkr04pO
T5sXkqLZKTjBKc4mOK3mH1IQqdCIIk83ltOED01hWPmsIv1roP1IFkxMw+xzlkZh
O2pzqUUi12t7NFguG2e0DaglMYdFKx6qoeDVy3tBewXKVEwE2FXC70bIWeNrjfdf
msn694sjbyHyhIW60Jtw29dxZYUtLIgYJ8lBqoWiOBXEqBZ8oSraECltZ4jZktbj
sSm1p4Yod/V1vz0CFXn89fgodHNF44XEjuPTQW+U5WpyE9fNrPAR/OuNLp7mMJ6c
50149MWtVlaEA7egq0E90+F4xfcuhQtO0qjUzPS5YDJW5U5e3jQsOutRJ44IFMlG
J8NN9fkUdD/f+Y91Bx4asfpoCF3UM6qnLPI7fio10hR6dKHN2vCGqQckHBa4/oN+
l2syFCDzJEVN02pCkPt05Q==
`protect END_PROTECTED
