`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fhNb/jxjmPnGQLEhWrYm2kd3+SHbu9tbKQLrV2MmPuHmz16yw2RaBz73B4YbO3LE
H15ac79Ds2aBUm+FbMH0pO2w8p6dtfn7y0iV/CMnD5T44VLQZHuYqf+5uocjJmuJ
5ImKgq/k+p4zL6jG2j42foUmXoOErOoGWM+idC79/nz2ypujvelXtMNqfD4lLJWy
UNIkwiTx6QdMohnPfymra7tGu66+OSn4sKm2ahdSYymaw2C0II2lM1WxG5+OqA+c
mLN3dPpwDLtMCTJ8o8lN5W6JaTAU19tO3nflgnruVRpb+xr45frFLgI9KINcCj87
ShahUcbBwou1igzFvBH9VGzQkJcxWKPlGNbXJZNpuDbCoJHehAY9Nzuk+G2Wwdaw
9BVoCi/jI61nDxY8PJSmyEwBQWTeOaInSg/OPiXQAtZRPQB+PUjmAUNjZjBOyxci
aPKUzAcPhgj87aJ6ZWC41YTd4FHnKZe5XtJBUh03cnGNcu29JM6i7E384fqrRB3D
`protect END_PROTECTED
