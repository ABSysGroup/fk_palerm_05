`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sqqki7w0oPbRcCOhOnorBtmAxKAyneMP9uU5AUuMB82LiYYChiZXtu87DRmi1svL
edNSfU1fZ87XLfL1SmiM1uNSzUW9TEc9wWT7wXUwLWZp6SrOAc+bGyzjbxpcFnqt
tgBTkNciutxmELSvdkJGIaOh3FKJbjEN27ZVqY5Gf4OqHoOrfWKn36qR36IpaSXf
BzRFRQAosm/q898wkB0weBgIqN9oMm6OfUdcQiWVUwG2KXdPsU1tTeC0BmiUpXeD
88HPOeCnY2iuk5Ota9FjXLZrlIfwl4DYzCpcwTCubAY6OWbzCEaD3TGHBGq8YFTU
s0YuygQS+9wObwYPjeNfeAP9+Z67hAgovrhcqx+tAjIyRlmQE5+p0PWuV2274DJM
CBVa62BsNZ2Ak5DRDZSrDLWywOhxIC7awnSJF5lsaK4CcgAAuysV/k7OmP3xW0SP
6k45KfNb1kMWkr0S7P/NJWZ1XlRlaMrDVe0DSAz0pBVU6XzUF8DqoADwtWWo4wQ3
UPIXhfOz/VEWPbyVCGF0Ut6N7jRBvLCdB+5gjTFMnPi1WxSxDmQUrw2Kj0T0vXZv
`protect END_PROTECTED
