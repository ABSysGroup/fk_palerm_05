`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p04Lq1xrAIxErJQl/bZV1aMwglfysMMBoIK2xUJM8AWakIFd+DfrG0ivGFrESQuT
NQAEfkgJFhYS46JjCGPuXOAGu2Sh0Ir6XFcIS46q/DBl2SjGIlNAH7GqvX1Lm1E8
xcXapokkfhMeQdrD96H1IWNnzcpLQ7GwAFPLbvrajepLOmBHwawGED4f+D1rVhWS
4htCtj1K10t4qCqkNBl7Nlx3Y75ARXAS/QjJ0ts/OZsUIyvV/3njEONX8GXzDtyg
Gifro6Vp32xZSkRTv669kwLWAfrpc2FPCR9Hv9ynRfEOUBLuMs+JbPoZH23bw+h3
hx/edQKN2wmat5ppqCG9NdpwlnSw5tc/a/XLxGZ8T3or4mErLnnT14Ya42tBnkdG
+0H/CzIRzXS99BVAzCCfB186TCWlanwjE9R9e6Wbo+wZ+uNNEeG3p8prLGLP0KGf
xip/qP5Xp1EaidYYjT1nCO4CzUUF8bDJThHgqGqVsGGQuqGY8rF7BkJWJawC9Bye
4XzHcP8d7AbhTRzE7DUexd54nf8PvaUR6wQ7rpbqFSP+UvqVY8yGMiyyEtpMfTE8
mYF4fLcR1K0/CE7ew0lOUmh4qFksHwr4M1wD+cmzrwDJBWYJxLOQETrKq2RKgzFW
1r694nWlgYxKDmMjDn+lEOb7vcWYeQOGk7tihYDAN6XxaxH+SHhP02VQwlSVRo9Z
yHAo3sKeiwhV3abFF8AR58mVlY4J9r8ZQEUND1lpYvgPPtEIQfnmFFx1T6YL0O8n
gzZnf+yD+FYRfLtMh4DrmNz/o3ZsC47n0yYjGI+5ZhImvKye1DPsh1SzMAri3Da6
ODnGmvZ/CSBt5CDx9Cbt2p4Xx6dXtAj115Juy1SS4LwOulsxOVM6hVLVO+8XzPMa
5jFNf/1iqlobt7Z0YHeXpqWmF8pwrd0VNDDPlBWq/NE4tMl1EwLlm1vc5Omj5hZG
g3prtDZXuEaweMnSNL7uiLm9BwFPkd4lgQeP/B6zFZjJx4/6pbYUzs2mqSwLsj8i
4/Vg8EGIDw+1uUmRhpJQPK7cIcwc2Cv0FzLEgnOzWfdprizkmGksy6Ed1S9OhLfn
iW2AndHfGS1686YLyjapGbv0wzRLQRFDLYJRHMKIVapytoGWhuuvydIflh6xYXL0
6mkWS2MtDESknTwNuygcFpPTOiE17yak+n7Ili62tYk6uSsAXLYtRj4OX23Ge5D/
c0SnS/eHGOdqx4x3GcNpcwbq0l1hu4P4tgoQNCxJQDAlFiBb1GWBkzaIlXTvAViL
fBSsYb0Xx11Ui9KMayNBJFVMxvG115AyqoRW6hac97jdXxGVY4h3oZ2LC6U7DnOq
vEYcPSEmBH+Ro3de+cX/O/uEg84UTvFD83UPKOA/DSYoGZEuDBx0aOMGntMhM1Mw
pJdVCcrXRWemvpFixHyskDCMSn2/xrOqV3SP6Y+NFGReCPFNQ58VqqRCl6Nve5x3
0UtJwnQBfNXcoKjZPTXgPZ59lk6qWYmJTs1EZUj9prggU8oIRKFrX0BsIg9Emxud
2vjLu0Nszh2MxE8NzWRo7m+wxQ8kwaNaPVCmSxV9lzfzyRI7BLILf/czOZTUSVN2
DGJezkPbZkw3mTZSnMGt21vEp6WL4U2UUUZfH/RqMONvXaj3NnLL409MirSRMux0
9uzgcgHNz6uCLpR7JDWFCEkXq4knnFDCNX6UUo045CcJxohVA9Ef0SzVbaiJ7kTS
kKuIo1aLurwFafPno5v4rOiQREApnolSNeZv+8izHDLkSuOgBUhl0pkrVhLNGSmN
uyCy07VYpvQ+SIQIneLuLFiLLZ9zJpUAql1s2+8u2u4=
`protect END_PROTECTED
