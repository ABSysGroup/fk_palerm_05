`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uV2NvdbGLSy2b4uD9UotizHkKLxAVSm3upYjc5KpmvcE7CE+K1F9V6Zg2NZ7E04W
NkEoogZggsnvvYqow/rp8l3zmUT6VOhm/CYikeUblUJXkKKLE8WOYwU1Dxla0DYm
Cc9v23Ir5PsBgkWgXyBFpqgz+Qhd+8Ovc8RhJIRxy4c5YkOm819tRppFXNNRHiKS
kY21nn97sByFmniVqjsXJAg85qExUnx6udbV0rW76tQnoMJDhgs1DRcy321vLCE3
lE3UAz5IFOpP1I4yyqzxeWLkptU79/2mNPbgXpF6h6BzK2kykjGNdNCnTti4gLH8
dGRtYdfObp8cT76Ujxh4g35WHcUBnapWDujfJeJCxcMtEG3w+2qMkAGAnEB3RxgS
j7p9u38zZ8tha8ZyTLg9QCgD0AAm0jXQdAdD0wm+6QtG1gfq+B6XROhpfb4RfXZZ
1k8MBbTMfkhA+T3Iqw8OsvkQBaB8HzRCUaBnKKhslGcXGR2bdpLjiSQDMPMw/S16
gd4Zw5lXDX0Uztr141juVoqnx/3wsG9XYmydA8d9TJaHMIfabtd12CzPDJ5PGDBL
ikKzdduuhL4h+4beM3boCGAmjjJhH4vVBgoMg/KlB62aiiRrJ/FsIy+fNic1Yzaj
7l4kQlpvYTZI6CNcuPe2cCXdg8bjyhRtajebeynqAZKqG/4OJpvdDTfvkVlr5S2x
WoCRhkM0NOJpepCtvI9q30qBtJhCu7WtgTLTOSdiaJTOok0ki/fQOSD9jCTwpQhG
bcS7Iov76CrE75JlxNcbFeQ/rMVCVB22i6uDjJirYpVEV+kXCZBijrtcjjHqMYCm
QZiRZ/lANxK7U79aF5J4ziZY8/U360HL5dunRChOr9YkUER+avJc9zJYhUSOcLTy
uR2DjaiRMEC0LNWfnouruQ==
`protect END_PROTECTED
