`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oGl47Tc+e+KHoR1q/pUlanXLgbmrm3voC8+wT9RZm0sDW4tOKW7qPyxzIY2hN1Pi
6NFJx+LyQuE4xt/re6J6KvzeWYqr6vkBTFIg724tqQ8K49fiMPFXkwzNGlmVIvtZ
vpTYcfZkAKuXnVp7qYuKQzNZXZgfPA0QhYO/6oXH2vZ4N9RFdJ+lk2Fs0SRad/QR
Iu5qvv873EPqge7Yzv1ilnEiWZDQevtcBjnHJiWFhDoIHeFTcuWSjsRFjEjkI08t
eFfAKZywEjt96D24G/sv8JG9DAu1Vjd+N+1xz8CdfEvPIa6seekNr7eS9FU12IYa
aO2VmZgAg6VpeocM8uXJoXT+QlA9S3XpJf04f+qxlk4jchuA4eBghEjVtivwmKzo
YmzYl5BvgbEj2s5+V/xc/S/XG9vB2wfva+QWOIn3tuQFTEKUCU2HsV1YujBFeGaF
NJx6ze0Fs2QzNWE2PCLfS4G2tIRIsLoM+mdqmhkUX3wIguE1ol/7ZjjOB5FcRUNK
f/zv6CST+zpSeYXyZjlzQPbhKiUaYFDKkPZYqK3u4wA0h+Ky6o7yJ8J4vT1euTut
SE2uH2ZnMamq+7V1v+cffmI3W49AsJtZ9Y8geCRRlnzb7EWsSGgF4t08wycY7QeA
vCKfpm5MYqvZ+5BqjMALeTbRwIUeKKpWj0UJa5Wl1iMS5FxbhEBoUeaDbSEo+6fQ
dmDyFhcuL7HnT16wl6xlsaDOEhjDyCpVb58uwfULcxkmPGL/tvAyENfG7q//354k
tHRhctvESf4v1xWy3BBKE8yse430vtwdXuBmPRd6LtE5kYrOA1H0hWPtbr05sc4N
`protect END_PROTECTED
