`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x4Nn1QyMKSD2KEChUGPH368wN5acSz8Vs958V06SPYgK8sdHXtEV0qaecZ1M/xnF
5W8NxjMzJ5ri8kbBczPnqaYjrloO3w7ZfKGzR9h9inOJ9BsRkATuxKIohj6yuG1S
39HjqArt5UGdD1wfMoKeWw1BkNiitJGTgoPA1NkRtZgdoy4kOxkeGByJwQtWMepy
ukp7lIucN4V+gkNJflVEut9+7mUjzc0vFN7QVSAOmsqEsHq+nbTM+wC0F3NEnyhL
Yt9XLlWxYB7U5iOHhEqYICLa57VJ03Xm9j7xbYTQcBBVZ26R9YJI7QgcWz676Iq6
b+1scg+KV3Fsr+7uVlV8YJKQTQ0pGrMmD3Yo+Hfe2baeehDFzeOLiPqXnfCiv93T
ZnxgZqGoMjgty2ob5qqje5fBlyUp8TTQ80B2zAsrHaVIISXK2jWo3RS60KK3s2kh
Eq1I/zimloUq0IJd8XUHIKhwSNEkJKiW5ZenvIjyyq5PMg8hyaELHQQLaCvhqOPw
Rj4e664zUGKuj6+bfIfvfvPmi1Cnu6L2+Lgm42JypFvUx8TrA9oOPch94pjRTI7o
+r+P/KtUnnHk0laLycIORRVjFC23a9YEdZ6JfFvbcNGf3asN+62fUfO9g+Ms3dBI
pkHYI6qajUGsU08H9HjTvD0GxNX2aW/j/XIbocWuTPxp1dQOhsh/0wQ0Vz5PCui2
weAnigSYkuneVVbsFzLY1wZMEz2pWbk9+Im9FRjh48ix22TcuycqpVu9zvLCLxPc
C8JhuvQ6IWI/ZdOMCSFdL5YCsGyp8NkW7OAt6VSK+dIoGjQlOLEdpC+99oEIim6L
`protect END_PROTECTED
