`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uxe3abKzQQXnJDyvClIr3tte/Q6wYp10Os+wLIo6aqT6KaoXNtu0ZzFDtbWKwnT3
BDGnySQKAMRdb3yQHMyFIGhHcK/112Wg8jD6fhQUsYoi28030/AEfe+j2uWeZ96P
pLpS+YI67juSn4t73J9lPIf16f3KFYgtdM2tAfyD7xIizfAKICywUioNmF8HMN2C
lj7ZbkQio/+rZoO5KiGzcUn+ULJ0CaE97YCliH2Vvy2GP7KnBS20I1bpYLmlNJ24
bqPB93AfcyOo2eC7UpAGeOF/5ZltfSiw6VrCI15Z8fWXJHTJnr5yM4uxQUuBfzZY
Eq/hJfAtktMwzAdlQyO455gWr/jPW3P51D9q6LTMgI7OpIOsLsF3DT1U1B+gbtVO
pbITNYSCdNsFfkj68IfeJ6jJXOSm3wnNvgSB+dFXS9XQlewxcEV/uvYYGENRGDdi
jfM3KTkAQfcqrbrvBPKjg3lEOMJBVEAgu1xxfbVi/Xk=
`protect END_PROTECTED
