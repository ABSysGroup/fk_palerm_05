`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1UuSqCryfOPgV/P6IXSZaQZ4dCw1M4liYgCGfEIF62TTEOSeB4MUmxN0O0p1d0TI
ss46Pml+vFti/fp78M++4SoSrCTzfwBH9heKI/lzoL2ZwtZ8vF8BZIVAJuZDlxr+
j8KlbOYpkjD2lcfBXNXIv4OFctAB7XnvWMzfdfbwrAxrAzXaLpch5Ue4gI8YTvID
kyUoEQTHG20XJDhYTr/YJPJqM6lfCiafCVC2jb1XirRjzI8QJPNRTYNcOBDV0H1a
E9VGGDITr13l5weWo4DOc59046H4CiCqRHNKwFYzsNcawq+Kyt8uZJBkrkm1cBxw
zF3rfaFBO5eGa/v0S01G0OP/ZgKZvPeeKbum4uxdtWdV2ZFg7pGexLrHQYp8cd1W
BdxIsrQODKWKddI2e1cLs1fSky0KunRNPJ7o+4lD+gzO9PpxlARRYa3uDLFPEI3d
S7SIeSNxdeSWgue7D8snkWBYevj1kDq4M6p2E9YkTgAjprMO32n/mNN0CqRLtTQL
Op4wyISYitG0+r4emFkISnu4GSbytAdYmRSwsF/ZcSfQV357MIg2c7jxlBq730Jl
fiYPfgmefP+oWv1KWnuhuqXwAoMSj76y+pUruYJoUBQ=
`protect END_PROTECTED
