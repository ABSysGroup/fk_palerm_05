`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UnvSqMuEnYkjQUjOVE5NUQ3maQI4q5NbNpn+RIOe5TVv/2RR9j5GWHn1lquJDryZ
Rpf8pD22VwGbDlkHQ9UbIyj93CMCJa0XBLfJAtHf/p0vBNJz+jxfyj1B/YIsFxik
ouCPopkZm9xZgkeHfCT4GmKRuS8UF723h8NI8dpg5QUARCmq7AOnprHEJFot2248
OsJFS7c8vPNdUA8fkz5rakunkuXmd0K8mXMeSAsGvn+pqt6hDK3hplXc8hA8IBL4
9ldmplFiOBh4CE5Lioe3W88xOXi0HJw6T6bqwo/o4Lg83nyQ15VPGCeC6hQn5MeM
KAyh/Y4ETXS5lGnZbASJz0jhEl5I60zEaI11jPEMBoBxe95HRqe6cF3xifeBQITC
/6TfkrfVXI8aVN13+t3j6HAUFXCI6BfhYinJRhr4INGEgIb/ltjagiE3czgbGOTD
1bjj/uA5UFwnyxAI4uOLcVcsRYPQ2cAAfYkM1CaRs1NAJpFNHHI6b1mhNaVG0Xpa
yrTiHEFghgqQO8NxU5lwLlCbiaWWvNTzU2LKL3mLvzChcAeECE7alcIN4iOdb7Jf
+eQb4QOTd+1B1o9lfWo/4RSUvj3VFOotHhgLBRfiXvEyjGIEDWYbQOsRoMqV3++y
V4ljtJPjvstsM8gTi7MOZJxF5J7FfKKiexorHmUs6SY=
`protect END_PROTECTED
