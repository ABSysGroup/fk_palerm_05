`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZpheKpMbrvlpt/FmrYN17nDonaLnhzitQW8s+T19nGQMFC3imsbnlsyg+6IQDBu/
0kA92MLujtREmSx93X3aYMzg3uqvYAVdNs0t0GAUvJGdiU5rJeCkqh3UCnbxSkr2
8Q1Nqdc9ZtBzreDbRJ5YEjfU0ihkDiTWyOpPt1qzHLe9/NcgLDTYm54ZFXdoX+Rc
X/By/NiWxPN8FviJ35pXOqdvlmB1deX2BxR00XbJEKrXmevOOVr5USrxDsWmDywH
E8e65khRkNUtKMpSK7scYK53svmVldOfja56tZzOX496VYRe62M4XxEvMgr2TbYa
5I/35fnxPbQyBbBkXCG6WGmrASHGf83YBZb3tPXgmc5TF12I/OjERrxdlD6besdJ
LTTeW9Ztmfn7WnoFeYsGDNLmFOt+SkGKNz2Te3/WmxgrdccckvUBLWFoyIjrfwz2
xKCu7w+R9swGNdKWjBWPn32KegTeaBT34qqk189iA9eJGe0wAgIW50Z5sJQjSAtE
AfO6f86G4fC2FQJRN3HLZKQyLMbQU6RPfOqSe+j7orpXWSmSOnPQYEF4RPWW/CKH
nfkAxljqGBiqaKXKu7pI0Vo2hoW7ynfZbc+rYKgYaZ9G3+38tE/Jhlj2844gSj2Z
hEEwF2ivnhYULRFcY9lE3quHZ3Q4cgTb4ehuBOfklhLrvMl7/tRtV8EoauGrMi4e
rZ3Sivc1FR5pNO5NF6L9Sqda4Q7zfcJvBSQycwSXP1vvAtdwF2pGAAY0MIv05TqU
NrFjOJ/zuyMExzivn9ctM0fdfFU1Ee9pqcc0fWgmnqI9y6YtMCUgCJlWKIYGr+5J
47BINN22edCDDRDJuKCxEc599MI3+RqRBhnBepKFBSrf3hIhAW7zevtFoGP8EujZ
zyCdQqIE7iMZQv85c52VxMeDTqzGGzBCx8/3jPuUlWVsgCFsG1yPBvm8nvKZlmD9
uhtsHTRUzOETjAeUXafemIegaTlwQ1ev5DLP/R1a14Ex0UceR0PFquCANFK6Oshe
fywt7/JXv//MmT4tzm9a0Q==
`protect END_PROTECTED
