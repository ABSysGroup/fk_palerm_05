`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vBtHDPWYrh4V8aaPVD7wInoMfNgZ6UnCGP/YEcXqiJlqtGhm0+EvlD2djAOYYRsg
miSL9CUdiXnwRnMTJH14ckE/SWEhHhMNQEpeYXfeF+sQVIeQ93FID6RZ8tn+SJr6
EdU1NJ+KBdeGAbYhUur4eHEM9Ok9dLQOI/P6ZNtMYzTzB8MPiZ1g6fCGQLSXTZCe
DPWoEeTe9aM/O/Qo7I9SGjKMv553r451XDvgpLQbRhGWZNECCNHskJ0dmlGDQ8Yq
fmmh/LJdPdvPtz9lkXOyKY36/1OnWQqqbRIDlnUTa5Uo+68rbBl1cK/HmL6ZbCnS
Eds55ITDhMQ6ktHsbUzJBVIaD5MC9Zegrg4xjrl1Zujp5HUJ3DOvDdBQkDIwcOcF
dviQr53uggjmesAuhfVSZ58gZOdxPgVaqRGpgWPx3mk6eItIBz0K+KXr4sdiHuBQ
4k/3WJzAt89R2S5LCY1OCtHeRU+YzSzjyp/95BQHZzRao3077zr35URl7ea+xZr8
VnJIatdoZM78729Oz84/MDTY1jdjlh93gML7qgjderE3muMDgoLbjjqVye4eQMkB
Tzd5KwlKBk/l8FJhbGG3mzTsHr+7CqXby56Tp8btG1VTIC2hKdca3AQAW/vfwput
3uej7jtrtO5Vaoe9u/ZvetB6odjsIh87EluvdF7IM1tDyjk0FXYOln2/IinekjRr
4ipo+bsSqjibrFTdsbI2n7u8KwPjSaq7YYLlURS/1njXuXLWAWTaZ6x6gc1IjnCU
70xmznJJ8vN7bTPF9eQmgewzaAdR39HDW1EHR6V0Znx/NZYU36wmiL0OggBdZEHx
pT1M7HW3cPtgeuKlDgKng757xm18l7oEu5pvkadwAzrdozelV7MflP1sK6ZVfnP/
g9lpp7vUKoHIW1rP4w/5ROqDWEroQROlul3xflXrJO+XUYtIbecCvr2gyxrozdlz
Xo44a1QGfaT3UZd0Gw0h6C6C6CJu97Yu609M2+0ikJCHWTxs0KizrZ2AYYXNd6ec
3n/jfIJbSFks/HDyb+8G1yT8KacB7M3v8TU7JziRg+u7xKR4H7/qZ8TS3ArcO7q4
DhdAJfSObfwXX4W2GxiHBglNFN3m3uQGCsJRybBLWYIw26UOLgLnpsbbiNifuOKw
o17q21RC551GroXRpGEa/DG8SpR7cDDjtU0Y/a0z1vQ8iaWrQtbDtMP70CF0O3dJ
mfucbduOYdCc2fXrKq+o6tpLoANdR/IhdIfIgB7DPpb9ILqrc4z1KZgOXehyklwH
8IOBvtAa3sKOyFJK0BqrhuJBXEVIdhra8svChMuwvR7KL3xTd7AL5/Mpj6W0YItt
iS+tDrfpWLcJdp0b27hJkKAoywbvJA3+5RGtY1NR992dtQW8eEb2tYhx2dxmF+M6
Lp+Im13BEN+JVnf9iP/t4CcN70hCrwnRMTB+pDnmK/Gn8GuBkV6wPaQwvDCTEQyX
jCz8EBhE7b9M9GjjRyIWlQFNM1Vl1u38Vs8YwCYw0k/1amQQWbmn3BDoGUP//ENg
GqfUf+bN5g3RUB7GTdBVpCv0H15mwiQSYfpVpHebF2iYOzcPURlHJ2pdJAp18hpF
FiPWZL45kWoWtJWX+ay800wvpSBN2REeCsYvz7gMYDUBxS4za5G06X+Iy7jAv+Kb
npOYdbSqAR5wJwXxEvYsL7SD1GDdgLGiD9hoKnD/TxNB5Ht5tFuy27Ypa7Yn3G6f
NMRzkSDRrpCLYFfVBB6EAVVOSn6unjVwCkqy6WQf0Rj8lB/E5fD7g8Gkl+qF8gvO
TYHvHuX320xwTCd0qXrjKCxEj/HWS1BpQ2xTRCXltYg4zHF3UziLqrTfO9s9FgxM
zcD9Tb1ahF7aAp3nlbj4cCwkE4Layynd9VtW/k6qC4JSJ7PODO3Wh6fs30GGbdAP
/6rfTRlqj55wI4ncPfqO0/X5oMHGygyMrj3IeW/9eSpdiOz49+nzM/ZnMI2kMoeI
sKTFHvpm6hmjWma00jLVTotDZ2pL1X4KOGp+CGyIJ02jcz47e4Z+oOXWLrYgx+gO
0QduEAKbAcnnUGHQR0GKCLng/6KTJO3ka6TfG+O3cLe0LuJ76o+TQ8F94JBzQiq9
GFzpYFumSY+5dlrydX4VvGr1YGHpeUjhhPmXvyti+31aiQQEPpc2cZQLIdp+m4Cp
Yq7NdMXu1aXG1Hpm5/pNTepw0JuFBAGIdoQNbWHcSTDmLWMtqukLwSebdfqBvj5y
Z6tWJ0Sppvvk0D/gBTdxARVfRjCP42ed7U50svM40QikliTckNcvbvTqwpMbEFnr
TIbzfMp5R8QwAQ9pmd6YmXMQsc2b8OOihfUsIJ416JTUUi+9g/axPEPe2AMiEzq3
IwAnyVMQyqSl2xWC93Fr/Vc46zJmX3K3TZrtmqXLy4c6fKDMO0inmGegCFxXk7KJ
lCAnw8YHHhOrvb1uRSuliDklRmtRCjvUPHhcDWptjmDAUJoyLRiNPEayLDng+p0j
7w8SyXQi/nCRvUX8tdkFh09Bw4Xz+AG/5YBO60VMbBh8bH8uMQA69t/NBbFPmM8q
605vDZxZOHVYTLa2y5jy9g1RjBLjX0OazPDkKylWZDh0AOt193PApYIKm5CbUQmx
YKJDIwkO8mympqwcMul+1i8+hI7OMYP3sh6yaIFnuMLX4c8/ZbtUA2y+CdCEKTIM
JryYK7cmq3kzdNo10ItNy/28rf0fitTFJQ8fW7SjD+A5I3wukHwvVadDxMVObxSP
4KxZwyYUtaSkMNutbys3Vd5B/EwAB7RuUNLB1oQpI8Ej+u8POy4o2gHBHdPQbRF/
RlQ2xBqvQLFzhAP3VC5TjHla/WwbQcjJis8O+msfD8ZLOuwr0I1LGLhHMhWqsd4s
PCnd2VtVXeGmcex6xwp4T+RKBH1yT3WruXSibq+lP30OeoGjPq2KJZ49fr1jKjXp
ns3kSDzQinhLL6ho3PyElqZLY7S723eD019JFOjLHVH/rlQYaDG11V3CRhW4m0iB
tZHYXIUG+WKk+MaJX6KV+P+iqmz4REuNzOhdI2QKEJqCX9ymu4eHH8k1XxxdTGdI
Mh4T/+ChW/laqjbzAeew05iIRVH7iOwSS2AqhkR9Z2pej9lSADgGRZ/fHt81MG4a
qyIJzlJsZk2oaTfhlmfvvU5h03T1d742/f0sNlz798/qH8n5C9s3xGOICnJOxQzR
5HbViTV9xiaZ8lN3R/AxccUypOZn10Qbvn8fY0M2oH2edhTQFPGZPGdkHqqErC9K
ftxxYHb58qt/cm1pg6Moej4xSGjSpSYS/Gx+pXfg033TLwa9Aqx3k0lN+aXdB/wr
kG0FxiO6w5AccFXTvElI/YUT29x0XVzPM2T7f1wIG8iIxF0X8tQMZO/DptuUP9W4
BzVPq5xbL92DNdFCkWhZRmmVxYhxZhp3eaxZhcDXyw4jBFI/H9bXRcvSPIbCYJtS
D8MbhvxrLwmJIgi7eptfMTVkc3hT6nklOcG3A8K15PMRIRHiceRIlHoNpQAUBTEr
SOlrXBA8inWW7TW00Pr8X+djxgaGP8XbinUW6oaoYnji8LLBxeFn8yuLfs4f20p2
yFasuxvndJ2VUVZ5qnk8F1xH9vBwXyjJ3jrXzXy2HuWrFGF/yZejx95AmQIM1uuR
NePDWx07lbZd8kLomTg+brn2ubng1T7NjyE/y6lNtuzSdY8gvEyTIaft+ZGiccUK
waw1Wnr5jjNck7ixW1XaJOcoWMG5g2LUEFGdkRTbbV0xX7Fm3m8Zq0eHvpWAPJp0
DoSUxlcp/5WX/qNeDyU402czZjB2p4nYhZf/1GBppM8wZ2H1n+/33untJcFNyLYt
EnLmUoBe67aLn4bDoHhLfPAW/4pzxix4jw5J7fYV0oMICWAZJsO91NrZ4dfKG7eq
7/3KwI4FNgy7kqj1mmKcPnInFlFceHHEeejYhY0fIyq/sT3d//cLQiSngSmhcPON
+0sEhgKtjbBgIrHr9b19sGeCnb2VM8wknY0/nV3pJv+picLTp0RLmJjaN8RpFnc/
aFMsECz/obwSUqjeNCSe6Wr2F8xIHQIVqlvFjLgokoNJExNOLmcd62AUo0NQkx2E
3CQ/k3+Yg8A9qzFb0Y+ffb99KiEXUXNi7+C1/WE2REDy1XeJlKq8K+cpJRUkFwO+
+dVTJTYS/Wdp/kIOwTTGRU7MeV/y7GNTMG9nLiP1cBAON20yCm4Ks1ubYkgMDUsG
5w0Hgy+Dcg34aKduqB1gJEtYtKZjnEuG+R3eZ5Eu9bwg27gebXYsjLyPG3LzRk1/
7v8E+6kI3urwsTXXEF8UNPS8iT1T+5zAMdNmMZ+FXMjkGhVPAvBQ0FYKNkV227D1
0H5uekjY+cBJ/dKZfJ6LAVThqrqA10PVBO5R+IYYe6PvgqSxGknE4TIq+tMN+Vbf
nk5596RvNfc1YsQ81YrImYJtoH1+AlqqhmeL+fQzEdx6ZYzfb6om5HdImYLogJ52
RNkI0kAlwsX21J7VdHAMGD2/jciqITZc7A0dWLMWMc43f4ZWFaTftyZs36T/SmPg
/ip9XGhS3cPhhYeEU7vPfXKJ+dPTTfJxOUbKd9Jw6GW7ELgkhzFkdJjpgVxJg5rW
kOz3MJ/BbaisPvNygy5aeASkPth922c+XJUG4VE614SUtc+3GV/h8goqgbtMlJy1
H1DBCRk7FWS4ISEabu/uYEy4W8HD0bHgqgRbxOzVuFV7l4XYJoBSBdDp1S8yRK33
PteEzyA71selBPdTzhPJfmQBM3GDQg7FyEXUEPre3JmRZz3oX5+S/0a39xaHBdVc
iVBqDRrZqtb95RTJsr3McHyRUUoGKuCtOaPzvCF9MtCZqf9d2MMmVsfkibW9zL/x
k9pe9yJdsYF+QlvigqwWONU8+esrPWyEcesGTXo/sV35Bpf9IZA3JmERXFNjRQFt
X+Q5ssA9Zg/gNiWHcPJf7D03kKy5xJ9tr/EmGgXuQ+VsD4Zd0DKv+DEKVs1u3vQe
Aq9uJmQaBIvRrW/nsHFKBZ7GZtheRGPy9966YzeA666FeVued/kTIhQyUxlx176I
m2My1X7lETplAsYgvr1VIPhf4vqqcLxzUnyIGscxy0qr+G6TZt1Piy4DSsKk0w6i
z/Lwdn5ep4euhWKKz2sAl4GXoU+uCnaaid3f3pQ1pzz2AuKtoH1hh+F0YWNpqq7D
6AQer1l2CKO9DBax5uO3yFgavgK82U1NY/x6NpahJ1BC0dDcIlrDYoIiBnTJb2xP
jO+5CtUVzdDLrjnRCu5QgEkPZAhQnDG1Qq62hFDdbTs08WGdNs2bKpKOyKZ/alZ9
glaYYyHHhR4D5k7ka6leQri/nf6uFuy69dqtKLJ+dIOUn+NqkWqt0I0qO47fpo/M
S0oFCNdw9fVDgABpBlaDGO0MrVcroXRum45R0wnv54giDbj92AkoUCkWpGumCy7W
9ReVrbXsndCvFQnL9YIagdxldAaMiWdvtv6LjpUz7F4wxtmhAHTeKMKwA2nBu80s
ldwVac6M7P4C0ZHc0rYrXzelm78tfDSwB9lvT4T8/g0w4V4+8PKEK688PydWIhlG
el3jsYM36r0vaHfUsjlYd0Iz9bKVbVCnDqo6QZhcKyiIUksTVuYxeDhYURicgaMG
pDQQANmi6iiUqInaf5UMokv593dJ+FInnhx2k7x3cII93d2z5rN5mGJqPSCb1O2a
tjNFifA7MbYB9xUjmiQuC1vJ2vVPsa7WMRzYhgadpxxDttdAgPd4FMXu7zNrhPhf
2KWgix48HDs++MZ4EktRvDEhf2eAtsSyH5JF10+fylxXTpVZxdUhZ/QSUx+eDjJh
spf5lHofAcw02MA3QzsX4CbqZpmgp9v44+Av+ZrJm7q6aYMIhfk3uWZB+aIg+lIb
CMXoKeOj22yttIaxRI3gDcQtHL9myhxJ0d6XWzxA0XevjopP1TEPxgosxRxKQ2EC
`protect END_PROTECTED
