`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EFP70d/rHUVA4KQKvv/j7qPhJ4NZXmnNHjnJgHs7VLpN3p4LWj9rW3964hYiaq6D
ZlCn6MF3QwqKHGWTY2rjM93iJ3ETR9MBZRw0fpYzE/6G6uIC0V4lpPx4kako/hyn
45Y0/WrkjMCIcZJ3DGrPx8wQZ/MAa88/eTaj0J689SiZxEe/yV3bCgzurcoplyrB
7bTrf4/8hgjVWX6pFuwK0cttrwngTEuTyTbBBqiDM62FJfM2FOblF1voqa/jZCdh
EihUNKiDNtleKC6NXctuFQ==
`protect END_PROTECTED
