`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aoZd2wMH81oAIrtJtYcP8Y2akX/vts8kpLXLDnUplKCZPHrC/iI7N4W6iuFfnBlA
YvvnjZ3euygTfE3/53O4ykVti6MHtbXzRNXr9QcS+y1mp5pE/RP+dyeYS/2nsKAu
lpGWHuSlnXctnRhv02v9RAZTK0itPWibtT5UeDC0bqOfApunmyA3RsToDoHLo1Si
7tpjCXIBjhx+s/8UcTEdAx1ZeifQKu4TR5rFT+du76TurIoknlJfnRYA1dNI9l2S
9O4ug5p4dOb89eflpb7TzjPTAZ9odpg36SSXZoUsCTC8Iv1XDLj5tOHJM2BkNOoG
`protect END_PROTECTED
