`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CiBALOrtkoHzlMPlbnBlaM81OiTOB9iEYg7xtkxOcTt1309WLDbibjTVpAa91HGk
DXTxrrOuzni6S1jqycBLLgzBMRG1BUQQa2IYBtjxJLUj4x0uYbgzROm8le1y776n
SKSV+pCNqbQTwjFtyWgF9QX0DEgt4j7rs+V/S/CNG0Y9eL/BfK8Spg+zxXo8xEon
MiTe8wyxjySp4RbUrXXMT8jJPgDDtSB+b0/4szIHnBOml3/CF7Opcvnbl7YIqdFf
mPpmgRMTc1mrlqYfUu7WJw==
`protect END_PROTECTED
