`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
43fM34c2GXTschg6fWeghGPtorz4joGaj/5w7uX1+OelwwkGoNy3kPAjPyYu8Mal
jsCa0k1qtTWu6uqymovZ+NcDDtjZd5/E7C37ufWJwC2tHV+ILqVw5box1I4XlzXV
PaHBam5kelOW4gkb4RE72+PZ6Wc/3PKA6VX4WOZS9Rvg+zOyct9p91KxGShBEhuD
Z1DBLC/jUMg98SHKkeMN4JXu0p663ypLLYYULHkJjJTd0AMq65+v9+yFz2nwnfe6
pudsx85iTC7LoqpNFlgiWTuUhIL815SAjJxIYdEf6FWOC8EeSlRqvI4kL5pfRIbX
ZYrLURNcCrOaLu6xqxs8ChAkzPMXKq1lOBTAKJ6SpjHqHFWk1X1J2OfqaNr/zK/M
MMRwOXLkOH+GqzQiIqaqmfLmGpLlFclzRwvbCeqovioqBA642Si6rKYQj5nCQ1kX
Sk3/Ac2vi6G4Vf4pvsSbZAHdvRZeGyn/GszCxZeNzrz1opPoIzXZoIUr/hl0e9s9
h3kFgUBQefS47DoKolZsBCCwQCzL+VHLYHN9ev4jnw5pj1CwS7zyk3WmNl5QJsSc
ihj0ughykfcyfbz6u2Eb+kbJoFzrsBS/avQ8qITXIlUztSazVTx24tUzU78PTQCV
hpzLRrJBiD0fUjv6f2ljm8xqsJKL8VdjBFYVPt/miT+bQlVb8lFhak00yo/9qnEG
r+f2bIc9OqQzp3SYgimQLoeH7W80AWhSv29ZX1T4Vcp5LmmBHzKsCkEuQmOkBMp5
KrDHbkuwnm6oR/bMZ6gUUkHd32Z7YPfCmoj/wZtLu6QGnmUgv1EXhzVfg+QCRXzk
26yWkfjFrx3KuT5QK562xw==
`protect END_PROTECTED
