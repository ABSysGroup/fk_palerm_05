`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PZS8BVm/SRx4M5n6DI2/vyJQ0QQcxoUH+XoL50xECuZB4oNLPR0ui60H/RfUeBFu
b8hXPl1hvWGhv9j24zIBG4uoVt49r/ixAa606tkN6nil3TgPHO9/NNMlMMe+PiD2
B2B2uRO8LJHsbuvcCEb8YOB/CG8E45WEr11JIfp87s+tsJtiLsVnSfotObFM1LvU
xRS1GavzVuaa5fyiyFDTjct+4NnjAGSsdYtwqNftGGrfVssmUK7ZRDDkYmYUcdg7
svt4iAo5CBDXV5PBoWqSV077HT1CXp0vHsswj2z9Ly0wvwvj1mqsVVRmeDJiArPC
m4mV1u1O91LjtoWoRJZdkCGGLxk9bVFzwTeIxMETbksRUwtCNbGek6yNWQkh+ia6
+S75VLtqLfIuwPw+l7e7CNDpT9euS8nO4EVCaxOE83P2Oc2xQlU5FHX6SJSi2lG7
PZ4YsIetwKkvOP0POlbmUPjV9hM8slEaeRVxFqlI4agAl3qe34+uHMeJknGrKL+C
S/5qMCGIVzXpeue3jLd6ab0mVLGrlx8V4qk4SCTdUB7+vUEB/+guigfwMQ+LggBt
yAzG159VaCk1a8z17HhJy9iL7LlgWZ3q16H3DgcsFbY=
`protect END_PROTECTED
