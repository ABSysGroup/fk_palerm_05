`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AFfSQoIz5G40wtyCYEH9EWSBBRw8ABqfxM4Lx1Uy3T10aOPmVaC2IGYdtxy4oc2y
QOl0qcrOlxBveXsyO9PCshs9CEtNhjnM/cmf0W3IjgxMOnAHkRBGJW7jiCjVjE7+
fxsTRDEzelzSTom7/hTNUGFztSIFnxCZ7Xy9b2yms2Psg81BR70Tda6+HqZy3q6f
rKp/X950ecYlzAoYfjOFEjOqo9+Ol4W9YOTagl/3G3NIBZcPqH0S/wCSxDY7xttP
`protect END_PROTECTED
