`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z5fyCbYvdOJ7pVE4OA3FfLX00FUGCyHO9YzwDbhMXas5P6deX0rTSiEoRJl72O7L
Q2wb9o8+p9beMPgGQ6ducaxx6zmC3xAT7ILHyQDEr6nOkqYyO0XH250FYZH3Eae/
JL3BPfwoisyYBBUco/VvPcNGHkUIO6l/D7qlv5BwJrZ4omOT4yWDYPAP3I/if2nj
n11t1FdWVqv06uKMnUH5R/OV2Sdpq5PguRakE+b9E2X0wq1mf4mOSJd2U7M70BDi
7h4UUiTvrmhZ7uHj+NIaqKSRqbVc8K0XJxg98MQOzWn8xXYKxSnAke4iCVidmdll
AYyHUQK4Y6rDX+06asdoA8fbIg71TjuRvhtVmM8gWhOu6W8wTqKW96pPQtb4QDtq
L17gSRumErCNNSpIVaU4+IHs8g8U0FOk0dAsiTTtJ7jYd25Fev6A6/fw6qmO2bUn
`protect END_PROTECTED
