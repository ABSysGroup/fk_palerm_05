`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IpPfjmB2UFGRNP0/14wlCtzxS5FGvw+dT2ASxBGXCFuKLxWGXui+nTVCXfCKJnm6
5WMWzAPDAn+LOu05zuT3TZXPwoHUPLFfdAV7wJSe29ve9cRLXM64saw5j7R5Em5/
35Qp6YNquzjYlFhU3adJyVBpYWZYBiICo9/nKs6RYmax1ktekvwMBqJlyhlqhEes
RD1jV1aSlhzRFHVGrFTVR1ok6MaOo6hP3rxNyP2ELAOLHbHajD23m2UqcDoq8zPe
u56ycAMdwJSWo780bzahw5K1Ah4ECAVbrfHjt9WwfuIVO+px+S4T8DwyKfuMuxAs
XqvSs6YfWYpJQgzQZFJdcW6+WP1ELYlGd1uluFDKkWGD6/bd8QTphnJoNmqKD1PA
6F3Clkjshpw9RvVsDCc4UNk98jlbm5TqvZe30NoCeaY=
`protect END_PROTECTED
