`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eFZqAL9DSKx5xtlmQbATPDgXE4g0C/ajKalgJQDr+DYbCO2pvj5AdotxqCBM62Ao
Y2ii9mThmllvAS5CrSFksqViVKkqN9C2WSa60F8w6OnCrUQNQfuosblp54MwBiEZ
vgO/MFMHjAcQgKZsYEiYvUvH2JlAAeC5tZJF+93ZmORLQvRnUhuhQv+C2Ku8VaZS
iSrrRQHAHqGqPwiSSYZ4TnCG6UxIEKhEd3WmnZXcG2ao+QVqSQEeXyptH3O/ZMXJ
Rkcpgo1dDDjUWRdde9nDnUnQZzArNZy2CDBAiNNf/+4+pIB2ijo2iY7JBkMQklnq
zHH91cRToeXFi8/0lmekeqSpetHoZwhICeJdoMTiO1EuKd/6zR3fD1t3C1VinhMg
ahRs0FCXXyrTPQfQzJ17RwzZafTHLyHagEgom4WrsGXDTIriH97a8aNSJYXXB8EN
9M+dX0qX8Oa0yBU0nEyjOlXZNrOL4UM9Bc+lpSL9myRJcC249HzyoC/eC5q4j7hP
BstDwOGca6xC+fOgBjUcrjDrd2klAkLD2DorbFoXs6Ni77rkxSmLIlaDvoqOKtxx
1fSzceveqgGPaXRVHib3HWMpc/K7F+Z7pCM9irAVMJ1NJfQ3Rt43DibRwd/MdRMX
wrCUeuYfwhFZEA9O1+cZQoCYxWUs4ONaen5aeCfLdno=
`protect END_PROTECTED
