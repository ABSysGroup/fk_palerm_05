`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yHc6dJyJw2kkODPLnMPYCfegYXVLV7el9mTml+bRQw91UAXxMpLAI+gSy3nJ/oSU
SMwLWg205z1mE4xck8RlGX2OhIN0jjDZ3LmudWo7bMuFDsUCPoZhJZ1CRJNnLyd3
U4/vkm6swz0Z9EH0EOsJBjIBnfJ2Adr97JqjJzNZ88lMbSXDCZ7I3SJVGBNoS4qa
sd4eBE/lSBd0X3WDQ5dy34zjZmBORiUdwpS785j81RVmaTHqt6DvT9RVXbPEfArj
jXKleLv+9OwADBaLgDu6HJzvQ+bbR23GeS0rXNvjGOq5PvtPHJUfgt++vCjNbCpl
bNAMom70gWn0jNOhFsYyxtDipx71slI6Ifv6arErzYju1yfKz6cX5bsmi45+l8yt
bCkt0JJXZsjfdPDDBBK+JwIL5FMwF5Mk7rauW8DCUpTKe7atm7D9bE2fzaaZwEVq
6CVYsmPQaOaXHVnxbP8QTeEZx7RjgcqXB9wb0ULjzhbtBKesePUDut7HhsdYhL6V
2FGmAZDYT2VrmMUDrEZ+VtkCD2oX0iRMzok/p7MpJpqMhrmVM31Xgon6Z2fQeYqw
0I9g/gT98ZM8dFC2+UHQOD0qYHQPY2HMAsIj1aSbaeiVRYzPopdZYBmX45dyePOh
VK9YX1C4pNV1QBBDx1/wiZHX8zoqrH8ez/oe6DbjGIK+G+3ugDVtMs6RvQkE09JT
O/lSaftlh0gm9i0RnCkxI+E7zu7aPgBXHMMZp/5U0wB8+doNfwIH/lhy2l1etCUm
TNNsVTjVNMYTJ/pZCRiwag==
`protect END_PROTECTED
