`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ReUz6LtvLYxSU1H3rIpPUsEFkhO1wUdCzmg0+gHkxTYURvqFdhD7mhoz6V9PkBqZ
hLPAVCq+niz+v/iElUQ/lW03oye8FHuLPJnUwz12l6vjbV0y2fxJkci2Mk4kEIoV
TuyleZ7iqbd8ROWMeWqLiwFC4/F3T1bVV5cAPU0AuvMNxFyesrGSkPo/98GniVQz
Oo9h4328kPIyoiuIXUkCn9xhjrkyJU4gD7G73mJKfO+ReFTbcFWf01O5W4Wr6u6y
gjqRCTSQ7+i4H8uPqhoI786wkPlaNo1SKGbnGMlQ9mew8ZkqNXCZtMcWjUL+Zbbh
ARxzKsniPd+81RjntSS0MeiLe/GXwq1IfBeW5qZhIzQ+zaD/wCHnMh2RDdPU6M/a
/kqgr8VOT+tNVxp0bztSfYbE1/d8/zNwJBlsb6nbuiU=
`protect END_PROTECTED
