`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vhzvy+DVGR++L63/42UYPVW2iarlK5TNLs+zANxLmtxQAscvyePW9e9anSKW1XHd
dFD9zG8HQGwDiYAF1tnQzJy0CzCNQA12l9ti0TLe3oKdlUXcPhTcZQgPvSmSsPh4
V2FEvVo1Iq+mNWLga0Muk3Fsy2P86CdflXilLrqoJx5Ff8XSFJ2AefPSh6My9DBx
52iEjNV+JvkBQAfo+KrupeaB6i5gOJjmnukKwTewSz/SZtamN2GTwzXuLNQXC5KD
jidhFsT1K64Hu+oWYPunoVpkNDfjJQdFERwJYBWRB5X8TQcK0GmjVcwum4MJI2s5
kfmjicFzXtoJ9f+WaGAyvA==
`protect END_PROTECTED
