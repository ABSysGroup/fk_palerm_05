`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a0slTcaqbXsXr7dgYzzEz+Phafm36l+gCqZJzTwKSbBj/XdTWWWwvbaMIGw0pnOZ
7P8HI1JynbAoRqweMDRyVVQson/MkM5yyZ8eJpb9Tac5xRqPNWGjczLYpRDY05p7
xZnzBXejfM7nf8Pm29cnKOvWI2TUTe8Jf+qmzx5/eadDe0eLl9KXL6iacO6Bf6ur
41XR8vSQ6wI7DENAKaQL0kfhUeJFO6sFcXclbvlBtwcdqIyXi9b0W+Dyv7j5OmLj
z/UjM/t38RuQYsCGoxywJ4VKNRBM8Jn2f53ql1rO0UjTx6ygQ9WgEPGayYmCS4Iu
dxlwyG6BHA7RSAEx0mZnhw==
`protect END_PROTECTED
