`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7jUsGOCBJ2mBV74mKZXC1OWHgmVWLD2i22osZhFMm5e7pcTgzh0U5wePM+KARgQd
5WBV5lieqom0GJlk/3xDBZse01F8MBhgV9UCOQHGAm6dt9mbI1hlY/iuWbShM201
/cJx0dOxg1Y/TLVSSfbxa8cb1ZakMjL5Tys5U8D3BEGWTSjFvLmh/nFvQ1mYnYs5
yZIJ6U0OHpSjuoEuoVVbpTOP5zBUqb4aX4bhWfRQDInvXL56IZ/PgpwrPauYTjN9
6NWgcD2Th4ZnodBV650+hkn7Y4gWS0msMyUuzZ6QDlc+AuRZ8Lx86gbvN3x01Ekc
ApU6tEW+rSPrZq1ioVyHlNnc5QTSLQ68U/DHhjo1vPXs12G3DKkVGjcrlxF9FkV+
rya9NF2gmqD6zWYvVatUg0M9vdz0671w1iOm8Qgd1aw5oMGruKnEetVCpaV0RRdQ
9UAYiCrHY6K+FeidO2EplCAf2zb2OdlSlw1MeuKSfOcpxzlZZVGgs/cGJlru08AC
KTd7ENXG/22jseXjpCrhEA==
`protect END_PROTECTED
